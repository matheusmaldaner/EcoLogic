library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(2559 downto 0);
    signal layer1_outputs: std_logic_vector(2559 downto 0);
    signal layer2_outputs: std_logic_vector(2559 downto 0);
    signal layer3_outputs: std_logic_vector(2559 downto 0);
    signal layer4_outputs: std_logic_vector(2559 downto 0);
    signal layer5_outputs: std_logic_vector(2559 downto 0);
    signal layer6_outputs: std_logic_vector(2559 downto 0);
    signal layer7_outputs: std_logic_vector(2559 downto 0);
    signal layer8_outputs: std_logic_vector(2559 downto 0);

begin
    layer0_outputs(0) <= 1'b0;
    layer0_outputs(1) <= not b or a;
    layer0_outputs(2) <= 1'b1;
    layer0_outputs(3) <= a xor b;
    layer0_outputs(4) <= not (a or b);
    layer0_outputs(5) <= a xor b;
    layer0_outputs(6) <= b;
    layer0_outputs(7) <= not a;
    layer0_outputs(8) <= a;
    layer0_outputs(9) <= a or b;
    layer0_outputs(10) <= not b;
    layer0_outputs(11) <= not (a xor b);
    layer0_outputs(12) <= not (a and b);
    layer0_outputs(13) <= not b;
    layer0_outputs(14) <= not (a or b);
    layer0_outputs(15) <= not a;
    layer0_outputs(16) <= 1'b0;
    layer0_outputs(17) <= a;
    layer0_outputs(18) <= a;
    layer0_outputs(19) <= a and b;
    layer0_outputs(20) <= b and not a;
    layer0_outputs(21) <= not (a or b);
    layer0_outputs(22) <= not b;
    layer0_outputs(23) <= 1'b1;
    layer0_outputs(24) <= a and b;
    layer0_outputs(25) <= a;
    layer0_outputs(26) <= not b or a;
    layer0_outputs(27) <= b;
    layer0_outputs(28) <= not a;
    layer0_outputs(29) <= a and not b;
    layer0_outputs(30) <= a and not b;
    layer0_outputs(31) <= a;
    layer0_outputs(32) <= not a;
    layer0_outputs(33) <= a and b;
    layer0_outputs(34) <= b and not a;
    layer0_outputs(35) <= b and not a;
    layer0_outputs(36) <= b;
    layer0_outputs(37) <= 1'b1;
    layer0_outputs(38) <= a xor b;
    layer0_outputs(39) <= not b;
    layer0_outputs(40) <= not a;
    layer0_outputs(41) <= not a;
    layer0_outputs(42) <= not (a and b);
    layer0_outputs(43) <= not a or b;
    layer0_outputs(44) <= not a or b;
    layer0_outputs(45) <= not b;
    layer0_outputs(46) <= not a;
    layer0_outputs(47) <= not (a and b);
    layer0_outputs(48) <= not b or a;
    layer0_outputs(49) <= 1'b1;
    layer0_outputs(50) <= not (a and b);
    layer0_outputs(51) <= b;
    layer0_outputs(52) <= not b or a;
    layer0_outputs(53) <= b;
    layer0_outputs(54) <= not b or a;
    layer0_outputs(55) <= a and not b;
    layer0_outputs(56) <= a and not b;
    layer0_outputs(57) <= b;
    layer0_outputs(58) <= b;
    layer0_outputs(59) <= b;
    layer0_outputs(60) <= a;
    layer0_outputs(61) <= 1'b0;
    layer0_outputs(62) <= 1'b1;
    layer0_outputs(63) <= not a;
    layer0_outputs(64) <= b;
    layer0_outputs(65) <= a and b;
    layer0_outputs(66) <= 1'b0;
    layer0_outputs(67) <= not a or b;
    layer0_outputs(68) <= a;
    layer0_outputs(69) <= a or b;
    layer0_outputs(70) <= not (a or b);
    layer0_outputs(71) <= a;
    layer0_outputs(72) <= a and b;
    layer0_outputs(73) <= a and b;
    layer0_outputs(74) <= 1'b1;
    layer0_outputs(75) <= a and not b;
    layer0_outputs(76) <= b;
    layer0_outputs(77) <= a;
    layer0_outputs(78) <= not (a or b);
    layer0_outputs(79) <= not b;
    layer0_outputs(80) <= a or b;
    layer0_outputs(81) <= 1'b1;
    layer0_outputs(82) <= not a;
    layer0_outputs(83) <= b and not a;
    layer0_outputs(84) <= not a;
    layer0_outputs(85) <= b and not a;
    layer0_outputs(86) <= a;
    layer0_outputs(87) <= not (a and b);
    layer0_outputs(88) <= not b or a;
    layer0_outputs(89) <= 1'b0;
    layer0_outputs(90) <= b;
    layer0_outputs(91) <= a;
    layer0_outputs(92) <= b;
    layer0_outputs(93) <= a or b;
    layer0_outputs(94) <= not b;
    layer0_outputs(95) <= not a or b;
    layer0_outputs(96) <= a and b;
    layer0_outputs(97) <= b;
    layer0_outputs(98) <= b;
    layer0_outputs(99) <= b;
    layer0_outputs(100) <= not a or b;
    layer0_outputs(101) <= a and b;
    layer0_outputs(102) <= not (a xor b);
    layer0_outputs(103) <= 1'b1;
    layer0_outputs(104) <= not a or b;
    layer0_outputs(105) <= not (a and b);
    layer0_outputs(106) <= not a;
    layer0_outputs(107) <= not a or b;
    layer0_outputs(108) <= not a;
    layer0_outputs(109) <= not (a and b);
    layer0_outputs(110) <= not a;
    layer0_outputs(111) <= not b;
    layer0_outputs(112) <= not (a or b);
    layer0_outputs(113) <= not b;
    layer0_outputs(114) <= not (a or b);
    layer0_outputs(115) <= not a or b;
    layer0_outputs(116) <= not (a or b);
    layer0_outputs(117) <= not (a or b);
    layer0_outputs(118) <= 1'b1;
    layer0_outputs(119) <= 1'b0;
    layer0_outputs(120) <= a xor b;
    layer0_outputs(121) <= a or b;
    layer0_outputs(122) <= a;
    layer0_outputs(123) <= not (a or b);
    layer0_outputs(124) <= 1'b0;
    layer0_outputs(125) <= not a;
    layer0_outputs(126) <= not (a xor b);
    layer0_outputs(127) <= b and not a;
    layer0_outputs(128) <= a and not b;
    layer0_outputs(129) <= a xor b;
    layer0_outputs(130) <= a;
    layer0_outputs(131) <= a;
    layer0_outputs(132) <= not (a and b);
    layer0_outputs(133) <= not a or b;
    layer0_outputs(134) <= not (a xor b);
    layer0_outputs(135) <= a or b;
    layer0_outputs(136) <= not (a and b);
    layer0_outputs(137) <= b;
    layer0_outputs(138) <= not b;
    layer0_outputs(139) <= not a;
    layer0_outputs(140) <= a;
    layer0_outputs(141) <= not (a and b);
    layer0_outputs(142) <= not a;
    layer0_outputs(143) <= not a or b;
    layer0_outputs(144) <= 1'b1;
    layer0_outputs(145) <= a and not b;
    layer0_outputs(146) <= not a;
    layer0_outputs(147) <= not a;
    layer0_outputs(148) <= 1'b1;
    layer0_outputs(149) <= a and b;
    layer0_outputs(150) <= not b;
    layer0_outputs(151) <= not a or b;
    layer0_outputs(152) <= 1'b0;
    layer0_outputs(153) <= a and not b;
    layer0_outputs(154) <= not a or b;
    layer0_outputs(155) <= 1'b0;
    layer0_outputs(156) <= a and b;
    layer0_outputs(157) <= a;
    layer0_outputs(158) <= a xor b;
    layer0_outputs(159) <= not a;
    layer0_outputs(160) <= 1'b0;
    layer0_outputs(161) <= a and b;
    layer0_outputs(162) <= a and not b;
    layer0_outputs(163) <= not b;
    layer0_outputs(164) <= b;
    layer0_outputs(165) <= not (a xor b);
    layer0_outputs(166) <= not b;
    layer0_outputs(167) <= not b or a;
    layer0_outputs(168) <= not (a or b);
    layer0_outputs(169) <= not (a xor b);
    layer0_outputs(170) <= not (a or b);
    layer0_outputs(171) <= not a or b;
    layer0_outputs(172) <= not b or a;
    layer0_outputs(173) <= 1'b1;
    layer0_outputs(174) <= 1'b1;
    layer0_outputs(175) <= not b;
    layer0_outputs(176) <= a and b;
    layer0_outputs(177) <= 1'b0;
    layer0_outputs(178) <= 1'b1;
    layer0_outputs(179) <= a and not b;
    layer0_outputs(180) <= a or b;
    layer0_outputs(181) <= not b or a;
    layer0_outputs(182) <= not b or a;
    layer0_outputs(183) <= not (a and b);
    layer0_outputs(184) <= not (a and b);
    layer0_outputs(185) <= not b;
    layer0_outputs(186) <= not (a or b);
    layer0_outputs(187) <= b and not a;
    layer0_outputs(188) <= 1'b1;
    layer0_outputs(189) <= a;
    layer0_outputs(190) <= not b or a;
    layer0_outputs(191) <= a and not b;
    layer0_outputs(192) <= not (a and b);
    layer0_outputs(193) <= a xor b;
    layer0_outputs(194) <= a;
    layer0_outputs(195) <= a xor b;
    layer0_outputs(196) <= 1'b1;
    layer0_outputs(197) <= not a or b;
    layer0_outputs(198) <= a and not b;
    layer0_outputs(199) <= a or b;
    layer0_outputs(200) <= not (a and b);
    layer0_outputs(201) <= 1'b0;
    layer0_outputs(202) <= a;
    layer0_outputs(203) <= not a;
    layer0_outputs(204) <= not a;
    layer0_outputs(205) <= a;
    layer0_outputs(206) <= b;
    layer0_outputs(207) <= not a;
    layer0_outputs(208) <= not b or a;
    layer0_outputs(209) <= not (a xor b);
    layer0_outputs(210) <= b;
    layer0_outputs(211) <= a or b;
    layer0_outputs(212) <= not (a or b);
    layer0_outputs(213) <= 1'b0;
    layer0_outputs(214) <= not (a and b);
    layer0_outputs(215) <= not (a or b);
    layer0_outputs(216) <= a xor b;
    layer0_outputs(217) <= a;
    layer0_outputs(218) <= a and not b;
    layer0_outputs(219) <= a and b;
    layer0_outputs(220) <= 1'b0;
    layer0_outputs(221) <= a;
    layer0_outputs(222) <= not b or a;
    layer0_outputs(223) <= a or b;
    layer0_outputs(224) <= 1'b0;
    layer0_outputs(225) <= b and not a;
    layer0_outputs(226) <= b;
    layer0_outputs(227) <= a;
    layer0_outputs(228) <= 1'b0;
    layer0_outputs(229) <= not a;
    layer0_outputs(230) <= not a or b;
    layer0_outputs(231) <= not a or b;
    layer0_outputs(232) <= 1'b0;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= b and not a;
    layer0_outputs(235) <= a;
    layer0_outputs(236) <= a;
    layer0_outputs(237) <= a or b;
    layer0_outputs(238) <= not b;
    layer0_outputs(239) <= not b;
    layer0_outputs(240) <= not b or a;
    layer0_outputs(241) <= not (a or b);
    layer0_outputs(242) <= not (a or b);
    layer0_outputs(243) <= a or b;
    layer0_outputs(244) <= 1'b1;
    layer0_outputs(245) <= a or b;
    layer0_outputs(246) <= 1'b1;
    layer0_outputs(247) <= not (a or b);
    layer0_outputs(248) <= not a;
    layer0_outputs(249) <= not b or a;
    layer0_outputs(250) <= not b;
    layer0_outputs(251) <= a;
    layer0_outputs(252) <= 1'b1;
    layer0_outputs(253) <= a;
    layer0_outputs(254) <= b;
    layer0_outputs(255) <= a and b;
    layer0_outputs(256) <= 1'b0;
    layer0_outputs(257) <= a xor b;
    layer0_outputs(258) <= not a or b;
    layer0_outputs(259) <= b;
    layer0_outputs(260) <= not a or b;
    layer0_outputs(261) <= 1'b0;
    layer0_outputs(262) <= 1'b0;
    layer0_outputs(263) <= a or b;
    layer0_outputs(264) <= not a or b;
    layer0_outputs(265) <= 1'b1;
    layer0_outputs(266) <= not b or a;
    layer0_outputs(267) <= not b;
    layer0_outputs(268) <= b and not a;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= b and not a;
    layer0_outputs(271) <= not a;
    layer0_outputs(272) <= a xor b;
    layer0_outputs(273) <= a xor b;
    layer0_outputs(274) <= not (a xor b);
    layer0_outputs(275) <= 1'b1;
    layer0_outputs(276) <= not b or a;
    layer0_outputs(277) <= a and not b;
    layer0_outputs(278) <= a;
    layer0_outputs(279) <= not (a or b);
    layer0_outputs(280) <= 1'b1;
    layer0_outputs(281) <= 1'b0;
    layer0_outputs(282) <= b;
    layer0_outputs(283) <= 1'b1;
    layer0_outputs(284) <= 1'b0;
    layer0_outputs(285) <= not a or b;
    layer0_outputs(286) <= not (a xor b);
    layer0_outputs(287) <= not b;
    layer0_outputs(288) <= 1'b1;
    layer0_outputs(289) <= not a;
    layer0_outputs(290) <= a;
    layer0_outputs(291) <= not a;
    layer0_outputs(292) <= b;
    layer0_outputs(293) <= 1'b1;
    layer0_outputs(294) <= 1'b0;
    layer0_outputs(295) <= not (a xor b);
    layer0_outputs(296) <= not a;
    layer0_outputs(297) <= not a or b;
    layer0_outputs(298) <= not b or a;
    layer0_outputs(299) <= a and not b;
    layer0_outputs(300) <= a and not b;
    layer0_outputs(301) <= not a;
    layer0_outputs(302) <= b;
    layer0_outputs(303) <= a xor b;
    layer0_outputs(304) <= a and b;
    layer0_outputs(305) <= not b;
    layer0_outputs(306) <= not a;
    layer0_outputs(307) <= b;
    layer0_outputs(308) <= 1'b0;
    layer0_outputs(309) <= a or b;
    layer0_outputs(310) <= not (a or b);
    layer0_outputs(311) <= a;
    layer0_outputs(312) <= a and b;
    layer0_outputs(313) <= not a;
    layer0_outputs(314) <= not (a and b);
    layer0_outputs(315) <= a and b;
    layer0_outputs(316) <= not a;
    layer0_outputs(317) <= not b;
    layer0_outputs(318) <= a xor b;
    layer0_outputs(319) <= a xor b;
    layer0_outputs(320) <= a and not b;
    layer0_outputs(321) <= not a;
    layer0_outputs(322) <= 1'b1;
    layer0_outputs(323) <= not (a xor b);
    layer0_outputs(324) <= b;
    layer0_outputs(325) <= a xor b;
    layer0_outputs(326) <= not a or b;
    layer0_outputs(327) <= not b;
    layer0_outputs(328) <= a and b;
    layer0_outputs(329) <= not (a xor b);
    layer0_outputs(330) <= a and b;
    layer0_outputs(331) <= not (a or b);
    layer0_outputs(332) <= not a or b;
    layer0_outputs(333) <= not b;
    layer0_outputs(334) <= not a;
    layer0_outputs(335) <= a;
    layer0_outputs(336) <= not a;
    layer0_outputs(337) <= a and b;
    layer0_outputs(338) <= not (a or b);
    layer0_outputs(339) <= 1'b1;
    layer0_outputs(340) <= 1'b1;
    layer0_outputs(341) <= 1'b1;
    layer0_outputs(342) <= 1'b1;
    layer0_outputs(343) <= not a or b;
    layer0_outputs(344) <= not a or b;
    layer0_outputs(345) <= not b;
    layer0_outputs(346) <= a;
    layer0_outputs(347) <= b;
    layer0_outputs(348) <= not a or b;
    layer0_outputs(349) <= 1'b1;
    layer0_outputs(350) <= 1'b1;
    layer0_outputs(351) <= a;
    layer0_outputs(352) <= 1'b1;
    layer0_outputs(353) <= b and not a;
    layer0_outputs(354) <= b;
    layer0_outputs(355) <= not a or b;
    layer0_outputs(356) <= not (a xor b);
    layer0_outputs(357) <= not (a xor b);
    layer0_outputs(358) <= not (a or b);
    layer0_outputs(359) <= a and b;
    layer0_outputs(360) <= b;
    layer0_outputs(361) <= 1'b1;
    layer0_outputs(362) <= 1'b1;
    layer0_outputs(363) <= a or b;
    layer0_outputs(364) <= 1'b1;
    layer0_outputs(365) <= a and not b;
    layer0_outputs(366) <= not (a or b);
    layer0_outputs(367) <= a;
    layer0_outputs(368) <= not (a and b);
    layer0_outputs(369) <= not b;
    layer0_outputs(370) <= a and b;
    layer0_outputs(371) <= not (a or b);
    layer0_outputs(372) <= 1'b0;
    layer0_outputs(373) <= not b or a;
    layer0_outputs(374) <= 1'b0;
    layer0_outputs(375) <= not a;
    layer0_outputs(376) <= a and b;
    layer0_outputs(377) <= b and not a;
    layer0_outputs(378) <= not a;
    layer0_outputs(379) <= a xor b;
    layer0_outputs(380) <= a or b;
    layer0_outputs(381) <= 1'b0;
    layer0_outputs(382) <= a xor b;
    layer0_outputs(383) <= not a;
    layer0_outputs(384) <= b;
    layer0_outputs(385) <= a;
    layer0_outputs(386) <= 1'b0;
    layer0_outputs(387) <= not a or b;
    layer0_outputs(388) <= a or b;
    layer0_outputs(389) <= a and b;
    layer0_outputs(390) <= a;
    layer0_outputs(391) <= not b or a;
    layer0_outputs(392) <= a and not b;
    layer0_outputs(393) <= not (a or b);
    layer0_outputs(394) <= not (a xor b);
    layer0_outputs(395) <= b;
    layer0_outputs(396) <= a;
    layer0_outputs(397) <= not b or a;
    layer0_outputs(398) <= a and b;
    layer0_outputs(399) <= 1'b0;
    layer0_outputs(400) <= not (a and b);
    layer0_outputs(401) <= b;
    layer0_outputs(402) <= a;
    layer0_outputs(403) <= b;
    layer0_outputs(404) <= a and not b;
    layer0_outputs(405) <= not a or b;
    layer0_outputs(406) <= 1'b1;
    layer0_outputs(407) <= b and not a;
    layer0_outputs(408) <= b;
    layer0_outputs(409) <= a or b;
    layer0_outputs(410) <= not (a and b);
    layer0_outputs(411) <= a;
    layer0_outputs(412) <= not a;
    layer0_outputs(413) <= 1'b1;
    layer0_outputs(414) <= not b;
    layer0_outputs(415) <= a and b;
    layer0_outputs(416) <= not b;
    layer0_outputs(417) <= not b;
    layer0_outputs(418) <= a;
    layer0_outputs(419) <= a and b;
    layer0_outputs(420) <= a and not b;
    layer0_outputs(421) <= a and b;
    layer0_outputs(422) <= a xor b;
    layer0_outputs(423) <= not a;
    layer0_outputs(424) <= a or b;
    layer0_outputs(425) <= 1'b0;
    layer0_outputs(426) <= b and not a;
    layer0_outputs(427) <= a;
    layer0_outputs(428) <= b and not a;
    layer0_outputs(429) <= a xor b;
    layer0_outputs(430) <= b and not a;
    layer0_outputs(431) <= not (a and b);
    layer0_outputs(432) <= not a or b;
    layer0_outputs(433) <= b;
    layer0_outputs(434) <= not (a or b);
    layer0_outputs(435) <= not a or b;
    layer0_outputs(436) <= not (a or b);
    layer0_outputs(437) <= a and b;
    layer0_outputs(438) <= b and not a;
    layer0_outputs(439) <= b and not a;
    layer0_outputs(440) <= 1'b0;
    layer0_outputs(441) <= not (a or b);
    layer0_outputs(442) <= not b;
    layer0_outputs(443) <= not (a and b);
    layer0_outputs(444) <= a or b;
    layer0_outputs(445) <= b;
    layer0_outputs(446) <= not b or a;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= a;
    layer0_outputs(449) <= not a;
    layer0_outputs(450) <= not a;
    layer0_outputs(451) <= not b or a;
    layer0_outputs(452) <= b;
    layer0_outputs(453) <= not (a or b);
    layer0_outputs(454) <= b and not a;
    layer0_outputs(455) <= not (a or b);
    layer0_outputs(456) <= b and not a;
    layer0_outputs(457) <= not (a xor b);
    layer0_outputs(458) <= not a or b;
    layer0_outputs(459) <= a;
    layer0_outputs(460) <= a and b;
    layer0_outputs(461) <= a and b;
    layer0_outputs(462) <= b;
    layer0_outputs(463) <= b;
    layer0_outputs(464) <= b;
    layer0_outputs(465) <= a or b;
    layer0_outputs(466) <= b and not a;
    layer0_outputs(467) <= not b;
    layer0_outputs(468) <= b and not a;
    layer0_outputs(469) <= b;
    layer0_outputs(470) <= not a;
    layer0_outputs(471) <= a or b;
    layer0_outputs(472) <= not (a or b);
    layer0_outputs(473) <= not a or b;
    layer0_outputs(474) <= not (a xor b);
    layer0_outputs(475) <= not a;
    layer0_outputs(476) <= not (a or b);
    layer0_outputs(477) <= not b;
    layer0_outputs(478) <= not (a and b);
    layer0_outputs(479) <= not a;
    layer0_outputs(480) <= 1'b0;
    layer0_outputs(481) <= not b or a;
    layer0_outputs(482) <= a xor b;
    layer0_outputs(483) <= 1'b1;
    layer0_outputs(484) <= 1'b0;
    layer0_outputs(485) <= b;
    layer0_outputs(486) <= b;
    layer0_outputs(487) <= not (a and b);
    layer0_outputs(488) <= not (a xor b);
    layer0_outputs(489) <= a or b;
    layer0_outputs(490) <= 1'b0;
    layer0_outputs(491) <= not (a xor b);
    layer0_outputs(492) <= b;
    layer0_outputs(493) <= a and b;
    layer0_outputs(494) <= not (a xor b);
    layer0_outputs(495) <= a or b;
    layer0_outputs(496) <= not (a or b);
    layer0_outputs(497) <= a or b;
    layer0_outputs(498) <= not (a xor b);
    layer0_outputs(499) <= b and not a;
    layer0_outputs(500) <= not a;
    layer0_outputs(501) <= 1'b1;
    layer0_outputs(502) <= b and not a;
    layer0_outputs(503) <= not (a or b);
    layer0_outputs(504) <= a or b;
    layer0_outputs(505) <= a and not b;
    layer0_outputs(506) <= b and not a;
    layer0_outputs(507) <= 1'b0;
    layer0_outputs(508) <= not (a xor b);
    layer0_outputs(509) <= not a or b;
    layer0_outputs(510) <= not b;
    layer0_outputs(511) <= 1'b0;
    layer0_outputs(512) <= b and not a;
    layer0_outputs(513) <= 1'b0;
    layer0_outputs(514) <= 1'b0;
    layer0_outputs(515) <= 1'b0;
    layer0_outputs(516) <= 1'b0;
    layer0_outputs(517) <= a and b;
    layer0_outputs(518) <= not b or a;
    layer0_outputs(519) <= b;
    layer0_outputs(520) <= not b or a;
    layer0_outputs(521) <= not (a or b);
    layer0_outputs(522) <= 1'b0;
    layer0_outputs(523) <= not a or b;
    layer0_outputs(524) <= not a or b;
    layer0_outputs(525) <= not a or b;
    layer0_outputs(526) <= not (a or b);
    layer0_outputs(527) <= not (a xor b);
    layer0_outputs(528) <= a and not b;
    layer0_outputs(529) <= a and not b;
    layer0_outputs(530) <= not b;
    layer0_outputs(531) <= not (a and b);
    layer0_outputs(532) <= not (a and b);
    layer0_outputs(533) <= 1'b1;
    layer0_outputs(534) <= a or b;
    layer0_outputs(535) <= a and b;
    layer0_outputs(536) <= a;
    layer0_outputs(537) <= a and b;
    layer0_outputs(538) <= a or b;
    layer0_outputs(539) <= not b;
    layer0_outputs(540) <= a and not b;
    layer0_outputs(541) <= a xor b;
    layer0_outputs(542) <= a and b;
    layer0_outputs(543) <= not a;
    layer0_outputs(544) <= not b or a;
    layer0_outputs(545) <= 1'b0;
    layer0_outputs(546) <= not a;
    layer0_outputs(547) <= not b or a;
    layer0_outputs(548) <= 1'b0;
    layer0_outputs(549) <= a and not b;
    layer0_outputs(550) <= 1'b0;
    layer0_outputs(551) <= 1'b1;
    layer0_outputs(552) <= b;
    layer0_outputs(553) <= 1'b0;
    layer0_outputs(554) <= 1'b1;
    layer0_outputs(555) <= not a or b;
    layer0_outputs(556) <= a or b;
    layer0_outputs(557) <= not a or b;
    layer0_outputs(558) <= not a or b;
    layer0_outputs(559) <= a or b;
    layer0_outputs(560) <= 1'b0;
    layer0_outputs(561) <= 1'b1;
    layer0_outputs(562) <= not (a or b);
    layer0_outputs(563) <= 1'b1;
    layer0_outputs(564) <= 1'b0;
    layer0_outputs(565) <= not a;
    layer0_outputs(566) <= a and b;
    layer0_outputs(567) <= 1'b0;
    layer0_outputs(568) <= 1'b0;
    layer0_outputs(569) <= not a;
    layer0_outputs(570) <= a and not b;
    layer0_outputs(571) <= not (a or b);
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= a and b;
    layer0_outputs(574) <= a;
    layer0_outputs(575) <= not b or a;
    layer0_outputs(576) <= b and not a;
    layer0_outputs(577) <= a and b;
    layer0_outputs(578) <= a or b;
    layer0_outputs(579) <= not (a and b);
    layer0_outputs(580) <= not (a and b);
    layer0_outputs(581) <= not b;
    layer0_outputs(582) <= not (a xor b);
    layer0_outputs(583) <= b and not a;
    layer0_outputs(584) <= 1'b1;
    layer0_outputs(585) <= a xor b;
    layer0_outputs(586) <= 1'b1;
    layer0_outputs(587) <= 1'b0;
    layer0_outputs(588) <= a;
    layer0_outputs(589) <= a or b;
    layer0_outputs(590) <= a or b;
    layer0_outputs(591) <= 1'b0;
    layer0_outputs(592) <= a;
    layer0_outputs(593) <= b and not a;
    layer0_outputs(594) <= a or b;
    layer0_outputs(595) <= a and b;
    layer0_outputs(596) <= b and not a;
    layer0_outputs(597) <= b and not a;
    layer0_outputs(598) <= a or b;
    layer0_outputs(599) <= not (a xor b);
    layer0_outputs(600) <= 1'b0;
    layer0_outputs(601) <= not a;
    layer0_outputs(602) <= 1'b0;
    layer0_outputs(603) <= not (a or b);
    layer0_outputs(604) <= 1'b1;
    layer0_outputs(605) <= 1'b1;
    layer0_outputs(606) <= a and not b;
    layer0_outputs(607) <= a and b;
    layer0_outputs(608) <= 1'b1;
    layer0_outputs(609) <= 1'b0;
    layer0_outputs(610) <= not a or b;
    layer0_outputs(611) <= not b;
    layer0_outputs(612) <= not (a or b);
    layer0_outputs(613) <= b and not a;
    layer0_outputs(614) <= a and b;
    layer0_outputs(615) <= 1'b0;
    layer0_outputs(616) <= a;
    layer0_outputs(617) <= b and not a;
    layer0_outputs(618) <= not (a or b);
    layer0_outputs(619) <= not b or a;
    layer0_outputs(620) <= not b;
    layer0_outputs(621) <= 1'b1;
    layer0_outputs(622) <= not a or b;
    layer0_outputs(623) <= 1'b1;
    layer0_outputs(624) <= b;
    layer0_outputs(625) <= b and not a;
    layer0_outputs(626) <= not a;
    layer0_outputs(627) <= b and not a;
    layer0_outputs(628) <= 1'b0;
    layer0_outputs(629) <= a or b;
    layer0_outputs(630) <= 1'b1;
    layer0_outputs(631) <= not a;
    layer0_outputs(632) <= a xor b;
    layer0_outputs(633) <= not a;
    layer0_outputs(634) <= not (a xor b);
    layer0_outputs(635) <= not (a and b);
    layer0_outputs(636) <= not a or b;
    layer0_outputs(637) <= b;
    layer0_outputs(638) <= not (a or b);
    layer0_outputs(639) <= 1'b1;
    layer0_outputs(640) <= not a or b;
    layer0_outputs(641) <= not (a or b);
    layer0_outputs(642) <= a or b;
    layer0_outputs(643) <= a xor b;
    layer0_outputs(644) <= a and b;
    layer0_outputs(645) <= not b;
    layer0_outputs(646) <= a and b;
    layer0_outputs(647) <= a or b;
    layer0_outputs(648) <= not a;
    layer0_outputs(649) <= not (a xor b);
    layer0_outputs(650) <= not b or a;
    layer0_outputs(651) <= a and b;
    layer0_outputs(652) <= not a;
    layer0_outputs(653) <= 1'b0;
    layer0_outputs(654) <= not a or b;
    layer0_outputs(655) <= a and b;
    layer0_outputs(656) <= a and b;
    layer0_outputs(657) <= not (a and b);
    layer0_outputs(658) <= not a;
    layer0_outputs(659) <= a or b;
    layer0_outputs(660) <= not a or b;
    layer0_outputs(661) <= a or b;
    layer0_outputs(662) <= 1'b1;
    layer0_outputs(663) <= not a;
    layer0_outputs(664) <= 1'b0;
    layer0_outputs(665) <= a and b;
    layer0_outputs(666) <= not (a and b);
    layer0_outputs(667) <= not a;
    layer0_outputs(668) <= not b;
    layer0_outputs(669) <= not (a or b);
    layer0_outputs(670) <= 1'b0;
    layer0_outputs(671) <= not a or b;
    layer0_outputs(672) <= 1'b0;
    layer0_outputs(673) <= not b or a;
    layer0_outputs(674) <= 1'b1;
    layer0_outputs(675) <= a and b;
    layer0_outputs(676) <= not a or b;
    layer0_outputs(677) <= 1'b0;
    layer0_outputs(678) <= not b or a;
    layer0_outputs(679) <= a;
    layer0_outputs(680) <= b;
    layer0_outputs(681) <= not a or b;
    layer0_outputs(682) <= 1'b0;
    layer0_outputs(683) <= a and b;
    layer0_outputs(684) <= not b;
    layer0_outputs(685) <= a or b;
    layer0_outputs(686) <= 1'b0;
    layer0_outputs(687) <= a and b;
    layer0_outputs(688) <= 1'b1;
    layer0_outputs(689) <= not a;
    layer0_outputs(690) <= not b;
    layer0_outputs(691) <= a and b;
    layer0_outputs(692) <= a or b;
    layer0_outputs(693) <= 1'b0;
    layer0_outputs(694) <= 1'b1;
    layer0_outputs(695) <= 1'b1;
    layer0_outputs(696) <= a and not b;
    layer0_outputs(697) <= b and not a;
    layer0_outputs(698) <= 1'b1;
    layer0_outputs(699) <= not (a and b);
    layer0_outputs(700) <= 1'b0;
    layer0_outputs(701) <= not a or b;
    layer0_outputs(702) <= 1'b1;
    layer0_outputs(703) <= 1'b1;
    layer0_outputs(704) <= not (a and b);
    layer0_outputs(705) <= a;
    layer0_outputs(706) <= not (a xor b);
    layer0_outputs(707) <= 1'b0;
    layer0_outputs(708) <= 1'b1;
    layer0_outputs(709) <= a or b;
    layer0_outputs(710) <= 1'b0;
    layer0_outputs(711) <= b and not a;
    layer0_outputs(712) <= not (a or b);
    layer0_outputs(713) <= not a;
    layer0_outputs(714) <= a xor b;
    layer0_outputs(715) <= a and b;
    layer0_outputs(716) <= 1'b1;
    layer0_outputs(717) <= 1'b0;
    layer0_outputs(718) <= not b;
    layer0_outputs(719) <= not b or a;
    layer0_outputs(720) <= not (a or b);
    layer0_outputs(721) <= 1'b0;
    layer0_outputs(722) <= a;
    layer0_outputs(723) <= a;
    layer0_outputs(724) <= 1'b1;
    layer0_outputs(725) <= a;
    layer0_outputs(726) <= a or b;
    layer0_outputs(727) <= 1'b1;
    layer0_outputs(728) <= b and not a;
    layer0_outputs(729) <= not (a or b);
    layer0_outputs(730) <= not a;
    layer0_outputs(731) <= a;
    layer0_outputs(732) <= a xor b;
    layer0_outputs(733) <= not a or b;
    layer0_outputs(734) <= a and b;
    layer0_outputs(735) <= b and not a;
    layer0_outputs(736) <= not b;
    layer0_outputs(737) <= a or b;
    layer0_outputs(738) <= not b or a;
    layer0_outputs(739) <= not (a or b);
    layer0_outputs(740) <= 1'b1;
    layer0_outputs(741) <= not a;
    layer0_outputs(742) <= not a or b;
    layer0_outputs(743) <= a;
    layer0_outputs(744) <= 1'b0;
    layer0_outputs(745) <= a xor b;
    layer0_outputs(746) <= b;
    layer0_outputs(747) <= not (a xor b);
    layer0_outputs(748) <= not a;
    layer0_outputs(749) <= not a;
    layer0_outputs(750) <= not b or a;
    layer0_outputs(751) <= not b;
    layer0_outputs(752) <= b;
    layer0_outputs(753) <= not a;
    layer0_outputs(754) <= not (a or b);
    layer0_outputs(755) <= not a;
    layer0_outputs(756) <= a and not b;
    layer0_outputs(757) <= b;
    layer0_outputs(758) <= not b;
    layer0_outputs(759) <= not b or a;
    layer0_outputs(760) <= not b;
    layer0_outputs(761) <= not a or b;
    layer0_outputs(762) <= not (a and b);
    layer0_outputs(763) <= not (a or b);
    layer0_outputs(764) <= a and b;
    layer0_outputs(765) <= a;
    layer0_outputs(766) <= 1'b0;
    layer0_outputs(767) <= not b or a;
    layer0_outputs(768) <= a and b;
    layer0_outputs(769) <= b and not a;
    layer0_outputs(770) <= not (a xor b);
    layer0_outputs(771) <= not b or a;
    layer0_outputs(772) <= 1'b0;
    layer0_outputs(773) <= not b;
    layer0_outputs(774) <= a;
    layer0_outputs(775) <= not a;
    layer0_outputs(776) <= b and not a;
    layer0_outputs(777) <= b and not a;
    layer0_outputs(778) <= 1'b0;
    layer0_outputs(779) <= not a;
    layer0_outputs(780) <= a;
    layer0_outputs(781) <= a;
    layer0_outputs(782) <= not b;
    layer0_outputs(783) <= 1'b1;
    layer0_outputs(784) <= b;
    layer0_outputs(785) <= not a;
    layer0_outputs(786) <= 1'b1;
    layer0_outputs(787) <= 1'b1;
    layer0_outputs(788) <= not a;
    layer0_outputs(789) <= 1'b1;
    layer0_outputs(790) <= a and not b;
    layer0_outputs(791) <= 1'b0;
    layer0_outputs(792) <= a and not b;
    layer0_outputs(793) <= a or b;
    layer0_outputs(794) <= b and not a;
    layer0_outputs(795) <= a;
    layer0_outputs(796) <= not (a xor b);
    layer0_outputs(797) <= a or b;
    layer0_outputs(798) <= not b or a;
    layer0_outputs(799) <= a;
    layer0_outputs(800) <= a and b;
    layer0_outputs(801) <= a or b;
    layer0_outputs(802) <= not a or b;
    layer0_outputs(803) <= not (a xor b);
    layer0_outputs(804) <= 1'b0;
    layer0_outputs(805) <= a;
    layer0_outputs(806) <= a;
    layer0_outputs(807) <= 1'b0;
    layer0_outputs(808) <= not (a or b);
    layer0_outputs(809) <= not b or a;
    layer0_outputs(810) <= a or b;
    layer0_outputs(811) <= b;
    layer0_outputs(812) <= not (a or b);
    layer0_outputs(813) <= 1'b1;
    layer0_outputs(814) <= a and b;
    layer0_outputs(815) <= not a or b;
    layer0_outputs(816) <= 1'b1;
    layer0_outputs(817) <= 1'b0;
    layer0_outputs(818) <= 1'b1;
    layer0_outputs(819) <= b;
    layer0_outputs(820) <= b;
    layer0_outputs(821) <= b;
    layer0_outputs(822) <= a;
    layer0_outputs(823) <= a xor b;
    layer0_outputs(824) <= not b;
    layer0_outputs(825) <= a or b;
    layer0_outputs(826) <= 1'b1;
    layer0_outputs(827) <= a or b;
    layer0_outputs(828) <= a or b;
    layer0_outputs(829) <= 1'b1;
    layer0_outputs(830) <= not b or a;
    layer0_outputs(831) <= a or b;
    layer0_outputs(832) <= a and b;
    layer0_outputs(833) <= not (a or b);
    layer0_outputs(834) <= not (a or b);
    layer0_outputs(835) <= 1'b0;
    layer0_outputs(836) <= not (a and b);
    layer0_outputs(837) <= not (a and b);
    layer0_outputs(838) <= a and not b;
    layer0_outputs(839) <= not b;
    layer0_outputs(840) <= not b;
    layer0_outputs(841) <= a and not b;
    layer0_outputs(842) <= a xor b;
    layer0_outputs(843) <= 1'b0;
    layer0_outputs(844) <= b;
    layer0_outputs(845) <= a and b;
    layer0_outputs(846) <= not b;
    layer0_outputs(847) <= 1'b0;
    layer0_outputs(848) <= not b;
    layer0_outputs(849) <= not (a or b);
    layer0_outputs(850) <= not (a and b);
    layer0_outputs(851) <= not b;
    layer0_outputs(852) <= not a or b;
    layer0_outputs(853) <= 1'b1;
    layer0_outputs(854) <= not a;
    layer0_outputs(855) <= not b or a;
    layer0_outputs(856) <= a xor b;
    layer0_outputs(857) <= not b;
    layer0_outputs(858) <= a and not b;
    layer0_outputs(859) <= b;
    layer0_outputs(860) <= a xor b;
    layer0_outputs(861) <= 1'b0;
    layer0_outputs(862) <= 1'b0;
    layer0_outputs(863) <= b and not a;
    layer0_outputs(864) <= not a;
    layer0_outputs(865) <= 1'b1;
    layer0_outputs(866) <= not (a or b);
    layer0_outputs(867) <= not a;
    layer0_outputs(868) <= 1'b0;
    layer0_outputs(869) <= not b or a;
    layer0_outputs(870) <= 1'b0;
    layer0_outputs(871) <= 1'b0;
    layer0_outputs(872) <= a;
    layer0_outputs(873) <= 1'b1;
    layer0_outputs(874) <= not (a or b);
    layer0_outputs(875) <= not a;
    layer0_outputs(876) <= 1'b1;
    layer0_outputs(877) <= a and not b;
    layer0_outputs(878) <= a or b;
    layer0_outputs(879) <= not a;
    layer0_outputs(880) <= not a;
    layer0_outputs(881) <= not b or a;
    layer0_outputs(882) <= not b;
    layer0_outputs(883) <= not a or b;
    layer0_outputs(884) <= not b or a;
    layer0_outputs(885) <= not b or a;
    layer0_outputs(886) <= not (a or b);
    layer0_outputs(887) <= 1'b1;
    layer0_outputs(888) <= not a;
    layer0_outputs(889) <= a and b;
    layer0_outputs(890) <= a and b;
    layer0_outputs(891) <= a;
    layer0_outputs(892) <= 1'b0;
    layer0_outputs(893) <= 1'b1;
    layer0_outputs(894) <= not (a or b);
    layer0_outputs(895) <= not a;
    layer0_outputs(896) <= b;
    layer0_outputs(897) <= a and b;
    layer0_outputs(898) <= b;
    layer0_outputs(899) <= a;
    layer0_outputs(900) <= a or b;
    layer0_outputs(901) <= not (a or b);
    layer0_outputs(902) <= not (a or b);
    layer0_outputs(903) <= b and not a;
    layer0_outputs(904) <= b;
    layer0_outputs(905) <= a;
    layer0_outputs(906) <= not b;
    layer0_outputs(907) <= a and b;
    layer0_outputs(908) <= a xor b;
    layer0_outputs(909) <= not (a and b);
    layer0_outputs(910) <= 1'b1;
    layer0_outputs(911) <= a and b;
    layer0_outputs(912) <= a and b;
    layer0_outputs(913) <= 1'b0;
    layer0_outputs(914) <= 1'b0;
    layer0_outputs(915) <= not b;
    layer0_outputs(916) <= b;
    layer0_outputs(917) <= 1'b1;
    layer0_outputs(918) <= 1'b1;
    layer0_outputs(919) <= b;
    layer0_outputs(920) <= not (a xor b);
    layer0_outputs(921) <= not a or b;
    layer0_outputs(922) <= not (a xor b);
    layer0_outputs(923) <= not b;
    layer0_outputs(924) <= a;
    layer0_outputs(925) <= a and not b;
    layer0_outputs(926) <= not b or a;
    layer0_outputs(927) <= not b or a;
    layer0_outputs(928) <= not (a or b);
    layer0_outputs(929) <= not (a and b);
    layer0_outputs(930) <= not (a xor b);
    layer0_outputs(931) <= not b or a;
    layer0_outputs(932) <= b;
    layer0_outputs(933) <= 1'b0;
    layer0_outputs(934) <= not b or a;
    layer0_outputs(935) <= not b or a;
    layer0_outputs(936) <= b and not a;
    layer0_outputs(937) <= b;
    layer0_outputs(938) <= not a;
    layer0_outputs(939) <= a;
    layer0_outputs(940) <= a or b;
    layer0_outputs(941) <= b;
    layer0_outputs(942) <= not (a and b);
    layer0_outputs(943) <= 1'b1;
    layer0_outputs(944) <= not (a and b);
    layer0_outputs(945) <= a;
    layer0_outputs(946) <= 1'b0;
    layer0_outputs(947) <= a xor b;
    layer0_outputs(948) <= 1'b1;
    layer0_outputs(949) <= not (a or b);
    layer0_outputs(950) <= a or b;
    layer0_outputs(951) <= not a or b;
    layer0_outputs(952) <= a or b;
    layer0_outputs(953) <= not (a and b);
    layer0_outputs(954) <= not a;
    layer0_outputs(955) <= a or b;
    layer0_outputs(956) <= 1'b1;
    layer0_outputs(957) <= b and not a;
    layer0_outputs(958) <= not a or b;
    layer0_outputs(959) <= not (a and b);
    layer0_outputs(960) <= 1'b1;
    layer0_outputs(961) <= not a or b;
    layer0_outputs(962) <= 1'b0;
    layer0_outputs(963) <= b and not a;
    layer0_outputs(964) <= a xor b;
    layer0_outputs(965) <= not (a or b);
    layer0_outputs(966) <= not (a and b);
    layer0_outputs(967) <= a xor b;
    layer0_outputs(968) <= not b or a;
    layer0_outputs(969) <= b;
    layer0_outputs(970) <= 1'b0;
    layer0_outputs(971) <= not a;
    layer0_outputs(972) <= not b or a;
    layer0_outputs(973) <= not (a or b);
    layer0_outputs(974) <= a or b;
    layer0_outputs(975) <= a and not b;
    layer0_outputs(976) <= a and b;
    layer0_outputs(977) <= b and not a;
    layer0_outputs(978) <= a and b;
    layer0_outputs(979) <= not (a xor b);
    layer0_outputs(980) <= not (a xor b);
    layer0_outputs(981) <= a and not b;
    layer0_outputs(982) <= not (a and b);
    layer0_outputs(983) <= a or b;
    layer0_outputs(984) <= not b or a;
    layer0_outputs(985) <= not (a or b);
    layer0_outputs(986) <= not (a or b);
    layer0_outputs(987) <= a and b;
    layer0_outputs(988) <= not (a and b);
    layer0_outputs(989) <= a and not b;
    layer0_outputs(990) <= not (a and b);
    layer0_outputs(991) <= a or b;
    layer0_outputs(992) <= a xor b;
    layer0_outputs(993) <= not b or a;
    layer0_outputs(994) <= b and not a;
    layer0_outputs(995) <= 1'b1;
    layer0_outputs(996) <= 1'b1;
    layer0_outputs(997) <= b and not a;
    layer0_outputs(998) <= a;
    layer0_outputs(999) <= 1'b1;
    layer0_outputs(1000) <= 1'b1;
    layer0_outputs(1001) <= not a;
    layer0_outputs(1002) <= 1'b0;
    layer0_outputs(1003) <= not a;
    layer0_outputs(1004) <= b;
    layer0_outputs(1005) <= not a or b;
    layer0_outputs(1006) <= a and b;
    layer0_outputs(1007) <= 1'b0;
    layer0_outputs(1008) <= b;
    layer0_outputs(1009) <= not (a xor b);
    layer0_outputs(1010) <= not (a and b);
    layer0_outputs(1011) <= a and b;
    layer0_outputs(1012) <= a or b;
    layer0_outputs(1013) <= b and not a;
    layer0_outputs(1014) <= b;
    layer0_outputs(1015) <= b;
    layer0_outputs(1016) <= a;
    layer0_outputs(1017) <= b and not a;
    layer0_outputs(1018) <= not a;
    layer0_outputs(1019) <= b;
    layer0_outputs(1020) <= not (a or b);
    layer0_outputs(1021) <= not (a or b);
    layer0_outputs(1022) <= a and not b;
    layer0_outputs(1023) <= not (a or b);
    layer0_outputs(1024) <= 1'b1;
    layer0_outputs(1025) <= a and b;
    layer0_outputs(1026) <= not (a and b);
    layer0_outputs(1027) <= not a;
    layer0_outputs(1028) <= 1'b1;
    layer0_outputs(1029) <= a;
    layer0_outputs(1030) <= 1'b0;
    layer0_outputs(1031) <= b;
    layer0_outputs(1032) <= not (a and b);
    layer0_outputs(1033) <= 1'b1;
    layer0_outputs(1034) <= not (a or b);
    layer0_outputs(1035) <= a xor b;
    layer0_outputs(1036) <= not (a and b);
    layer0_outputs(1037) <= b;
    layer0_outputs(1038) <= not (a xor b);
    layer0_outputs(1039) <= a and not b;
    layer0_outputs(1040) <= a or b;
    layer0_outputs(1041) <= a;
    layer0_outputs(1042) <= b and not a;
    layer0_outputs(1043) <= b;
    layer0_outputs(1044) <= not (a or b);
    layer0_outputs(1045) <= not b;
    layer0_outputs(1046) <= not a;
    layer0_outputs(1047) <= 1'b0;
    layer0_outputs(1048) <= a and not b;
    layer0_outputs(1049) <= 1'b1;
    layer0_outputs(1050) <= b and not a;
    layer0_outputs(1051) <= not b;
    layer0_outputs(1052) <= not b;
    layer0_outputs(1053) <= not (a and b);
    layer0_outputs(1054) <= not a or b;
    layer0_outputs(1055) <= not (a or b);
    layer0_outputs(1056) <= a and b;
    layer0_outputs(1057) <= b;
    layer0_outputs(1058) <= a xor b;
    layer0_outputs(1059) <= not b;
    layer0_outputs(1060) <= b and not a;
    layer0_outputs(1061) <= not b;
    layer0_outputs(1062) <= b and not a;
    layer0_outputs(1063) <= a and b;
    layer0_outputs(1064) <= a and not b;
    layer0_outputs(1065) <= not (a and b);
    layer0_outputs(1066) <= not a;
    layer0_outputs(1067) <= a or b;
    layer0_outputs(1068) <= not (a and b);
    layer0_outputs(1069) <= b;
    layer0_outputs(1070) <= 1'b1;
    layer0_outputs(1071) <= b;
    layer0_outputs(1072) <= not (a and b);
    layer0_outputs(1073) <= not b;
    layer0_outputs(1074) <= a or b;
    layer0_outputs(1075) <= b;
    layer0_outputs(1076) <= b and not a;
    layer0_outputs(1077) <= not a or b;
    layer0_outputs(1078) <= not a;
    layer0_outputs(1079) <= a xor b;
    layer0_outputs(1080) <= not (a xor b);
    layer0_outputs(1081) <= a and not b;
    layer0_outputs(1082) <= not b or a;
    layer0_outputs(1083) <= not a;
    layer0_outputs(1084) <= not a;
    layer0_outputs(1085) <= not (a or b);
    layer0_outputs(1086) <= 1'b1;
    layer0_outputs(1087) <= 1'b1;
    layer0_outputs(1088) <= a and b;
    layer0_outputs(1089) <= b;
    layer0_outputs(1090) <= 1'b1;
    layer0_outputs(1091) <= a and b;
    layer0_outputs(1092) <= 1'b1;
    layer0_outputs(1093) <= a and not b;
    layer0_outputs(1094) <= 1'b0;
    layer0_outputs(1095) <= 1'b0;
    layer0_outputs(1096) <= a xor b;
    layer0_outputs(1097) <= not a;
    layer0_outputs(1098) <= 1'b1;
    layer0_outputs(1099) <= 1'b1;
    layer0_outputs(1100) <= 1'b1;
    layer0_outputs(1101) <= not (a and b);
    layer0_outputs(1102) <= a or b;
    layer0_outputs(1103) <= not (a xor b);
    layer0_outputs(1104) <= not a;
    layer0_outputs(1105) <= not a;
    layer0_outputs(1106) <= 1'b1;
    layer0_outputs(1107) <= a xor b;
    layer0_outputs(1108) <= a or b;
    layer0_outputs(1109) <= not (a and b);
    layer0_outputs(1110) <= not (a and b);
    layer0_outputs(1111) <= b;
    layer0_outputs(1112) <= not b or a;
    layer0_outputs(1113) <= a and not b;
    layer0_outputs(1114) <= not b;
    layer0_outputs(1115) <= b;
    layer0_outputs(1116) <= 1'b0;
    layer0_outputs(1117) <= b and not a;
    layer0_outputs(1118) <= b and not a;
    layer0_outputs(1119) <= 1'b0;
    layer0_outputs(1120) <= not (a xor b);
    layer0_outputs(1121) <= not (a xor b);
    layer0_outputs(1122) <= not a;
    layer0_outputs(1123) <= not (a xor b);
    layer0_outputs(1124) <= not b or a;
    layer0_outputs(1125) <= a or b;
    layer0_outputs(1126) <= b;
    layer0_outputs(1127) <= not a or b;
    layer0_outputs(1128) <= not (a or b);
    layer0_outputs(1129) <= 1'b1;
    layer0_outputs(1130) <= not b;
    layer0_outputs(1131) <= not (a or b);
    layer0_outputs(1132) <= 1'b1;
    layer0_outputs(1133) <= not (a and b);
    layer0_outputs(1134) <= not (a or b);
    layer0_outputs(1135) <= not b;
    layer0_outputs(1136) <= not a or b;
    layer0_outputs(1137) <= 1'b0;
    layer0_outputs(1138) <= b and not a;
    layer0_outputs(1139) <= 1'b0;
    layer0_outputs(1140) <= b;
    layer0_outputs(1141) <= not a;
    layer0_outputs(1142) <= b;
    layer0_outputs(1143) <= not (a and b);
    layer0_outputs(1144) <= not (a xor b);
    layer0_outputs(1145) <= not (a xor b);
    layer0_outputs(1146) <= a and not b;
    layer0_outputs(1147) <= not (a and b);
    layer0_outputs(1148) <= a;
    layer0_outputs(1149) <= not (a or b);
    layer0_outputs(1150) <= 1'b1;
    layer0_outputs(1151) <= not b;
    layer0_outputs(1152) <= not a or b;
    layer0_outputs(1153) <= not (a and b);
    layer0_outputs(1154) <= b and not a;
    layer0_outputs(1155) <= not (a or b);
    layer0_outputs(1156) <= not b;
    layer0_outputs(1157) <= a;
    layer0_outputs(1158) <= a;
    layer0_outputs(1159) <= not (a and b);
    layer0_outputs(1160) <= a and b;
    layer0_outputs(1161) <= not a;
    layer0_outputs(1162) <= not a;
    layer0_outputs(1163) <= 1'b0;
    layer0_outputs(1164) <= a;
    layer0_outputs(1165) <= 1'b0;
    layer0_outputs(1166) <= 1'b1;
    layer0_outputs(1167) <= a and not b;
    layer0_outputs(1168) <= not a;
    layer0_outputs(1169) <= a;
    layer0_outputs(1170) <= a;
    layer0_outputs(1171) <= b and not a;
    layer0_outputs(1172) <= 1'b1;
    layer0_outputs(1173) <= 1'b1;
    layer0_outputs(1174) <= 1'b0;
    layer0_outputs(1175) <= a or b;
    layer0_outputs(1176) <= a and not b;
    layer0_outputs(1177) <= not (a or b);
    layer0_outputs(1178) <= not a;
    layer0_outputs(1179) <= a;
    layer0_outputs(1180) <= 1'b1;
    layer0_outputs(1181) <= not (a xor b);
    layer0_outputs(1182) <= a;
    layer0_outputs(1183) <= a xor b;
    layer0_outputs(1184) <= not (a and b);
    layer0_outputs(1185) <= b and not a;
    layer0_outputs(1186) <= 1'b1;
    layer0_outputs(1187) <= 1'b1;
    layer0_outputs(1188) <= 1'b0;
    layer0_outputs(1189) <= not (a xor b);
    layer0_outputs(1190) <= 1'b0;
    layer0_outputs(1191) <= a and b;
    layer0_outputs(1192) <= not (a xor b);
    layer0_outputs(1193) <= not (a and b);
    layer0_outputs(1194) <= not (a or b);
    layer0_outputs(1195) <= 1'b0;
    layer0_outputs(1196) <= a;
    layer0_outputs(1197) <= not a;
    layer0_outputs(1198) <= not (a or b);
    layer0_outputs(1199) <= 1'b1;
    layer0_outputs(1200) <= a or b;
    layer0_outputs(1201) <= 1'b0;
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= not b;
    layer0_outputs(1204) <= not b or a;
    layer0_outputs(1205) <= a or b;
    layer0_outputs(1206) <= a;
    layer0_outputs(1207) <= not a;
    layer0_outputs(1208) <= a;
    layer0_outputs(1209) <= a or b;
    layer0_outputs(1210) <= a xor b;
    layer0_outputs(1211) <= 1'b1;
    layer0_outputs(1212) <= not b;
    layer0_outputs(1213) <= a;
    layer0_outputs(1214) <= b and not a;
    layer0_outputs(1215) <= not a or b;
    layer0_outputs(1216) <= a;
    layer0_outputs(1217) <= 1'b1;
    layer0_outputs(1218) <= b;
    layer0_outputs(1219) <= a;
    layer0_outputs(1220) <= not (a xor b);
    layer0_outputs(1221) <= a and not b;
    layer0_outputs(1222) <= b;
    layer0_outputs(1223) <= a;
    layer0_outputs(1224) <= 1'b1;
    layer0_outputs(1225) <= not a;
    layer0_outputs(1226) <= a;
    layer0_outputs(1227) <= not (a or b);
    layer0_outputs(1228) <= not a;
    layer0_outputs(1229) <= b;
    layer0_outputs(1230) <= a;
    layer0_outputs(1231) <= a;
    layer0_outputs(1232) <= 1'b1;
    layer0_outputs(1233) <= not b or a;
    layer0_outputs(1234) <= b;
    layer0_outputs(1235) <= 1'b0;
    layer0_outputs(1236) <= not b or a;
    layer0_outputs(1237) <= 1'b1;
    layer0_outputs(1238) <= not b;
    layer0_outputs(1239) <= 1'b1;
    layer0_outputs(1240) <= not b;
    layer0_outputs(1241) <= not (a and b);
    layer0_outputs(1242) <= not b;
    layer0_outputs(1243) <= 1'b1;
    layer0_outputs(1244) <= a and b;
    layer0_outputs(1245) <= b and not a;
    layer0_outputs(1246) <= not a or b;
    layer0_outputs(1247) <= 1'b1;
    layer0_outputs(1248) <= a or b;
    layer0_outputs(1249) <= b;
    layer0_outputs(1250) <= 1'b1;
    layer0_outputs(1251) <= a and not b;
    layer0_outputs(1252) <= 1'b0;
    layer0_outputs(1253) <= b;
    layer0_outputs(1254) <= b;
    layer0_outputs(1255) <= not b;
    layer0_outputs(1256) <= 1'b1;
    layer0_outputs(1257) <= a xor b;
    layer0_outputs(1258) <= b and not a;
    layer0_outputs(1259) <= not b or a;
    layer0_outputs(1260) <= not (a or b);
    layer0_outputs(1261) <= not a;
    layer0_outputs(1262) <= b;
    layer0_outputs(1263) <= a;
    layer0_outputs(1264) <= a and b;
    layer0_outputs(1265) <= not a or b;
    layer0_outputs(1266) <= 1'b0;
    layer0_outputs(1267) <= b;
    layer0_outputs(1268) <= 1'b1;
    layer0_outputs(1269) <= not (a or b);
    layer0_outputs(1270) <= a and b;
    layer0_outputs(1271) <= not a;
    layer0_outputs(1272) <= not (a xor b);
    layer0_outputs(1273) <= b and not a;
    layer0_outputs(1274) <= 1'b0;
    layer0_outputs(1275) <= not b;
    layer0_outputs(1276) <= b;
    layer0_outputs(1277) <= a;
    layer0_outputs(1278) <= not b or a;
    layer0_outputs(1279) <= a and not b;
    layer0_outputs(1280) <= a or b;
    layer0_outputs(1281) <= a or b;
    layer0_outputs(1282) <= not a;
    layer0_outputs(1283) <= 1'b0;
    layer0_outputs(1284) <= b and not a;
    layer0_outputs(1285) <= not (a or b);
    layer0_outputs(1286) <= a and b;
    layer0_outputs(1287) <= 1'b1;
    layer0_outputs(1288) <= b;
    layer0_outputs(1289) <= not a or b;
    layer0_outputs(1290) <= not b;
    layer0_outputs(1291) <= not a;
    layer0_outputs(1292) <= a and not b;
    layer0_outputs(1293) <= not b or a;
    layer0_outputs(1294) <= not (a or b);
    layer0_outputs(1295) <= not a;
    layer0_outputs(1296) <= 1'b1;
    layer0_outputs(1297) <= not a or b;
    layer0_outputs(1298) <= a xor b;
    layer0_outputs(1299) <= a;
    layer0_outputs(1300) <= a;
    layer0_outputs(1301) <= not a or b;
    layer0_outputs(1302) <= a xor b;
    layer0_outputs(1303) <= b and not a;
    layer0_outputs(1304) <= not b;
    layer0_outputs(1305) <= not a;
    layer0_outputs(1306) <= a and not b;
    layer0_outputs(1307) <= b;
    layer0_outputs(1308) <= a xor b;
    layer0_outputs(1309) <= b and not a;
    layer0_outputs(1310) <= not b;
    layer0_outputs(1311) <= a and b;
    layer0_outputs(1312) <= b and not a;
    layer0_outputs(1313) <= not (a and b);
    layer0_outputs(1314) <= not (a or b);
    layer0_outputs(1315) <= not a or b;
    layer0_outputs(1316) <= not b or a;
    layer0_outputs(1317) <= not a;
    layer0_outputs(1318) <= b;
    layer0_outputs(1319) <= not (a or b);
    layer0_outputs(1320) <= not a;
    layer0_outputs(1321) <= a and not b;
    layer0_outputs(1322) <= 1'b1;
    layer0_outputs(1323) <= a or b;
    layer0_outputs(1324) <= a and b;
    layer0_outputs(1325) <= not a or b;
    layer0_outputs(1326) <= b and not a;
    layer0_outputs(1327) <= a;
    layer0_outputs(1328) <= not a;
    layer0_outputs(1329) <= a and b;
    layer0_outputs(1330) <= not b or a;
    layer0_outputs(1331) <= not (a or b);
    layer0_outputs(1332) <= not (a or b);
    layer0_outputs(1333) <= 1'b1;
    layer0_outputs(1334) <= not (a xor b);
    layer0_outputs(1335) <= b;
    layer0_outputs(1336) <= not b;
    layer0_outputs(1337) <= b;
    layer0_outputs(1338) <= 1'b0;
    layer0_outputs(1339) <= b and not a;
    layer0_outputs(1340) <= a and b;
    layer0_outputs(1341) <= not a;
    layer0_outputs(1342) <= not b;
    layer0_outputs(1343) <= b;
    layer0_outputs(1344) <= not a;
    layer0_outputs(1345) <= a and b;
    layer0_outputs(1346) <= not (a xor b);
    layer0_outputs(1347) <= not (a or b);
    layer0_outputs(1348) <= not a;
    layer0_outputs(1349) <= not a;
    layer0_outputs(1350) <= not a;
    layer0_outputs(1351) <= b;
    layer0_outputs(1352) <= a and b;
    layer0_outputs(1353) <= 1'b1;
    layer0_outputs(1354) <= a and not b;
    layer0_outputs(1355) <= 1'b1;
    layer0_outputs(1356) <= b;
    layer0_outputs(1357) <= not b or a;
    layer0_outputs(1358) <= not b;
    layer0_outputs(1359) <= b and not a;
    layer0_outputs(1360) <= b and not a;
    layer0_outputs(1361) <= not (a and b);
    layer0_outputs(1362) <= a;
    layer0_outputs(1363) <= 1'b1;
    layer0_outputs(1364) <= b;
    layer0_outputs(1365) <= a;
    layer0_outputs(1366) <= not a;
    layer0_outputs(1367) <= not (a or b);
    layer0_outputs(1368) <= 1'b1;
    layer0_outputs(1369) <= 1'b1;
    layer0_outputs(1370) <= b and not a;
    layer0_outputs(1371) <= not b or a;
    layer0_outputs(1372) <= not a;
    layer0_outputs(1373) <= not a;
    layer0_outputs(1374) <= not (a or b);
    layer0_outputs(1375) <= a;
    layer0_outputs(1376) <= a xor b;
    layer0_outputs(1377) <= not a;
    layer0_outputs(1378) <= not (a or b);
    layer0_outputs(1379) <= a;
    layer0_outputs(1380) <= 1'b1;
    layer0_outputs(1381) <= not b or a;
    layer0_outputs(1382) <= not b or a;
    layer0_outputs(1383) <= not (a and b);
    layer0_outputs(1384) <= 1'b1;
    layer0_outputs(1385) <= not a;
    layer0_outputs(1386) <= not (a xor b);
    layer0_outputs(1387) <= not a;
    layer0_outputs(1388) <= not (a and b);
    layer0_outputs(1389) <= a and not b;
    layer0_outputs(1390) <= not (a or b);
    layer0_outputs(1391) <= a;
    layer0_outputs(1392) <= not b or a;
    layer0_outputs(1393) <= not a;
    layer0_outputs(1394) <= 1'b0;
    layer0_outputs(1395) <= a and not b;
    layer0_outputs(1396) <= 1'b0;
    layer0_outputs(1397) <= not (a xor b);
    layer0_outputs(1398) <= not (a or b);
    layer0_outputs(1399) <= 1'b1;
    layer0_outputs(1400) <= not (a xor b);
    layer0_outputs(1401) <= 1'b0;
    layer0_outputs(1402) <= a;
    layer0_outputs(1403) <= not a or b;
    layer0_outputs(1404) <= a or b;
    layer0_outputs(1405) <= 1'b1;
    layer0_outputs(1406) <= a xor b;
    layer0_outputs(1407) <= a and not b;
    layer0_outputs(1408) <= 1'b1;
    layer0_outputs(1409) <= not (a or b);
    layer0_outputs(1410) <= not a or b;
    layer0_outputs(1411) <= b and not a;
    layer0_outputs(1412) <= a;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= b;
    layer0_outputs(1415) <= not (a or b);
    layer0_outputs(1416) <= a and not b;
    layer0_outputs(1417) <= a;
    layer0_outputs(1418) <= a and b;
    layer0_outputs(1419) <= not b or a;
    layer0_outputs(1420) <= not b or a;
    layer0_outputs(1421) <= a;
    layer0_outputs(1422) <= b;
    layer0_outputs(1423) <= 1'b1;
    layer0_outputs(1424) <= 1'b0;
    layer0_outputs(1425) <= a;
    layer0_outputs(1426) <= b and not a;
    layer0_outputs(1427) <= a or b;
    layer0_outputs(1428) <= a or b;
    layer0_outputs(1429) <= b;
    layer0_outputs(1430) <= a xor b;
    layer0_outputs(1431) <= not (a xor b);
    layer0_outputs(1432) <= 1'b0;
    layer0_outputs(1433) <= not b;
    layer0_outputs(1434) <= not a or b;
    layer0_outputs(1435) <= b;
    layer0_outputs(1436) <= not (a or b);
    layer0_outputs(1437) <= not b;
    layer0_outputs(1438) <= not (a or b);
    layer0_outputs(1439) <= not a;
    layer0_outputs(1440) <= a and not b;
    layer0_outputs(1441) <= a and b;
    layer0_outputs(1442) <= not a or b;
    layer0_outputs(1443) <= a or b;
    layer0_outputs(1444) <= a xor b;
    layer0_outputs(1445) <= b and not a;
    layer0_outputs(1446) <= a;
    layer0_outputs(1447) <= a;
    layer0_outputs(1448) <= a;
    layer0_outputs(1449) <= not a;
    layer0_outputs(1450) <= not a;
    layer0_outputs(1451) <= 1'b0;
    layer0_outputs(1452) <= b;
    layer0_outputs(1453) <= not (a and b);
    layer0_outputs(1454) <= 1'b0;
    layer0_outputs(1455) <= a and b;
    layer0_outputs(1456) <= a and b;
    layer0_outputs(1457) <= b;
    layer0_outputs(1458) <= a or b;
    layer0_outputs(1459) <= a and not b;
    layer0_outputs(1460) <= a or b;
    layer0_outputs(1461) <= 1'b1;
    layer0_outputs(1462) <= a and not b;
    layer0_outputs(1463) <= not a or b;
    layer0_outputs(1464) <= not b;
    layer0_outputs(1465) <= b;
    layer0_outputs(1466) <= 1'b0;
    layer0_outputs(1467) <= not (a and b);
    layer0_outputs(1468) <= not (a and b);
    layer0_outputs(1469) <= not b;
    layer0_outputs(1470) <= not a;
    layer0_outputs(1471) <= a xor b;
    layer0_outputs(1472) <= a or b;
    layer0_outputs(1473) <= a xor b;
    layer0_outputs(1474) <= a and not b;
    layer0_outputs(1475) <= 1'b0;
    layer0_outputs(1476) <= 1'b1;
    layer0_outputs(1477) <= not b or a;
    layer0_outputs(1478) <= 1'b1;
    layer0_outputs(1479) <= 1'b0;
    layer0_outputs(1480) <= not a;
    layer0_outputs(1481) <= not b or a;
    layer0_outputs(1482) <= not a;
    layer0_outputs(1483) <= b;
    layer0_outputs(1484) <= not a;
    layer0_outputs(1485) <= a or b;
    layer0_outputs(1486) <= a or b;
    layer0_outputs(1487) <= not (a and b);
    layer0_outputs(1488) <= a;
    layer0_outputs(1489) <= 1'b1;
    layer0_outputs(1490) <= not a;
    layer0_outputs(1491) <= not a;
    layer0_outputs(1492) <= 1'b1;
    layer0_outputs(1493) <= 1'b1;
    layer0_outputs(1494) <= not a;
    layer0_outputs(1495) <= a xor b;
    layer0_outputs(1496) <= b;
    layer0_outputs(1497) <= a;
    layer0_outputs(1498) <= 1'b0;
    layer0_outputs(1499) <= a and b;
    layer0_outputs(1500) <= 1'b0;
    layer0_outputs(1501) <= not b;
    layer0_outputs(1502) <= not (a or b);
    layer0_outputs(1503) <= not (a and b);
    layer0_outputs(1504) <= a and not b;
    layer0_outputs(1505) <= a and b;
    layer0_outputs(1506) <= 1'b0;
    layer0_outputs(1507) <= not a;
    layer0_outputs(1508) <= a;
    layer0_outputs(1509) <= not (a and b);
    layer0_outputs(1510) <= not (a and b);
    layer0_outputs(1511) <= 1'b0;
    layer0_outputs(1512) <= a xor b;
    layer0_outputs(1513) <= 1'b0;
    layer0_outputs(1514) <= b;
    layer0_outputs(1515) <= not b or a;
    layer0_outputs(1516) <= not b;
    layer0_outputs(1517) <= a;
    layer0_outputs(1518) <= a;
    layer0_outputs(1519) <= 1'b0;
    layer0_outputs(1520) <= 1'b1;
    layer0_outputs(1521) <= b;
    layer0_outputs(1522) <= a or b;
    layer0_outputs(1523) <= not a;
    layer0_outputs(1524) <= not (a or b);
    layer0_outputs(1525) <= not a;
    layer0_outputs(1526) <= a or b;
    layer0_outputs(1527) <= not b;
    layer0_outputs(1528) <= 1'b0;
    layer0_outputs(1529) <= 1'b0;
    layer0_outputs(1530) <= not a or b;
    layer0_outputs(1531) <= 1'b0;
    layer0_outputs(1532) <= b;
    layer0_outputs(1533) <= not b or a;
    layer0_outputs(1534) <= not b;
    layer0_outputs(1535) <= not b;
    layer0_outputs(1536) <= not a;
    layer0_outputs(1537) <= a;
    layer0_outputs(1538) <= not (a xor b);
    layer0_outputs(1539) <= not (a or b);
    layer0_outputs(1540) <= 1'b0;
    layer0_outputs(1541) <= a and not b;
    layer0_outputs(1542) <= 1'b0;
    layer0_outputs(1543) <= not a or b;
    layer0_outputs(1544) <= b and not a;
    layer0_outputs(1545) <= 1'b0;
    layer0_outputs(1546) <= not (a xor b);
    layer0_outputs(1547) <= a and b;
    layer0_outputs(1548) <= not a;
    layer0_outputs(1549) <= b and not a;
    layer0_outputs(1550) <= a and not b;
    layer0_outputs(1551) <= a;
    layer0_outputs(1552) <= not a;
    layer0_outputs(1553) <= 1'b0;
    layer0_outputs(1554) <= a and not b;
    layer0_outputs(1555) <= b and not a;
    layer0_outputs(1556) <= b and not a;
    layer0_outputs(1557) <= not b or a;
    layer0_outputs(1558) <= a and b;
    layer0_outputs(1559) <= not a or b;
    layer0_outputs(1560) <= not b;
    layer0_outputs(1561) <= b;
    layer0_outputs(1562) <= b and not a;
    layer0_outputs(1563) <= not (a or b);
    layer0_outputs(1564) <= a;
    layer0_outputs(1565) <= not b or a;
    layer0_outputs(1566) <= b and not a;
    layer0_outputs(1567) <= 1'b0;
    layer0_outputs(1568) <= b;
    layer0_outputs(1569) <= not (a and b);
    layer0_outputs(1570) <= a or b;
    layer0_outputs(1571) <= a or b;
    layer0_outputs(1572) <= 1'b1;
    layer0_outputs(1573) <= 1'b1;
    layer0_outputs(1574) <= not b or a;
    layer0_outputs(1575) <= not a;
    layer0_outputs(1576) <= b and not a;
    layer0_outputs(1577) <= b;
    layer0_outputs(1578) <= not b or a;
    layer0_outputs(1579) <= not (a or b);
    layer0_outputs(1580) <= b;
    layer0_outputs(1581) <= a;
    layer0_outputs(1582) <= not (a and b);
    layer0_outputs(1583) <= a or b;
    layer0_outputs(1584) <= not (a xor b);
    layer0_outputs(1585) <= 1'b0;
    layer0_outputs(1586) <= not b;
    layer0_outputs(1587) <= b and not a;
    layer0_outputs(1588) <= 1'b0;
    layer0_outputs(1589) <= a or b;
    layer0_outputs(1590) <= b and not a;
    layer0_outputs(1591) <= a and not b;
    layer0_outputs(1592) <= a and not b;
    layer0_outputs(1593) <= a;
    layer0_outputs(1594) <= not a;
    layer0_outputs(1595) <= b;
    layer0_outputs(1596) <= not a or b;
    layer0_outputs(1597) <= not b or a;
    layer0_outputs(1598) <= not (a xor b);
    layer0_outputs(1599) <= not (a and b);
    layer0_outputs(1600) <= not b;
    layer0_outputs(1601) <= b;
    layer0_outputs(1602) <= a or b;
    layer0_outputs(1603) <= b;
    layer0_outputs(1604) <= a or b;
    layer0_outputs(1605) <= 1'b0;
    layer0_outputs(1606) <= a or b;
    layer0_outputs(1607) <= 1'b0;
    layer0_outputs(1608) <= not (a xor b);
    layer0_outputs(1609) <= a xor b;
    layer0_outputs(1610) <= not (a xor b);
    layer0_outputs(1611) <= a xor b;
    layer0_outputs(1612) <= not (a xor b);
    layer0_outputs(1613) <= a xor b;
    layer0_outputs(1614) <= a and b;
    layer0_outputs(1615) <= 1'b1;
    layer0_outputs(1616) <= not a;
    layer0_outputs(1617) <= a and b;
    layer0_outputs(1618) <= b;
    layer0_outputs(1619) <= 1'b1;
    layer0_outputs(1620) <= not b or a;
    layer0_outputs(1621) <= not b;
    layer0_outputs(1622) <= not (a and b);
    layer0_outputs(1623) <= a;
    layer0_outputs(1624) <= b and not a;
    layer0_outputs(1625) <= not b or a;
    layer0_outputs(1626) <= a;
    layer0_outputs(1627) <= not (a and b);
    layer0_outputs(1628) <= a;
    layer0_outputs(1629) <= not a;
    layer0_outputs(1630) <= 1'b0;
    layer0_outputs(1631) <= not b;
    layer0_outputs(1632) <= b;
    layer0_outputs(1633) <= 1'b0;
    layer0_outputs(1634) <= b and not a;
    layer0_outputs(1635) <= not b or a;
    layer0_outputs(1636) <= b and not a;
    layer0_outputs(1637) <= a or b;
    layer0_outputs(1638) <= b;
    layer0_outputs(1639) <= a;
    layer0_outputs(1640) <= not a;
    layer0_outputs(1641) <= not b or a;
    layer0_outputs(1642) <= b and not a;
    layer0_outputs(1643) <= 1'b0;
    layer0_outputs(1644) <= b;
    layer0_outputs(1645) <= not b or a;
    layer0_outputs(1646) <= a or b;
    layer0_outputs(1647) <= a and b;
    layer0_outputs(1648) <= a and b;
    layer0_outputs(1649) <= not (a xor b);
    layer0_outputs(1650) <= a xor b;
    layer0_outputs(1651) <= a and not b;
    layer0_outputs(1652) <= 1'b0;
    layer0_outputs(1653) <= b;
    layer0_outputs(1654) <= not (a or b);
    layer0_outputs(1655) <= not (a or b);
    layer0_outputs(1656) <= not b;
    layer0_outputs(1657) <= b;
    layer0_outputs(1658) <= not b or a;
    layer0_outputs(1659) <= b;
    layer0_outputs(1660) <= 1'b0;
    layer0_outputs(1661) <= a;
    layer0_outputs(1662) <= not (a xor b);
    layer0_outputs(1663) <= not b or a;
    layer0_outputs(1664) <= a and not b;
    layer0_outputs(1665) <= 1'b1;
    layer0_outputs(1666) <= not b;
    layer0_outputs(1667) <= not a or b;
    layer0_outputs(1668) <= 1'b1;
    layer0_outputs(1669) <= a;
    layer0_outputs(1670) <= not (a xor b);
    layer0_outputs(1671) <= a and b;
    layer0_outputs(1672) <= 1'b1;
    layer0_outputs(1673) <= a xor b;
    layer0_outputs(1674) <= not (a or b);
    layer0_outputs(1675) <= not b or a;
    layer0_outputs(1676) <= a;
    layer0_outputs(1677) <= b;
    layer0_outputs(1678) <= b;
    layer0_outputs(1679) <= a;
    layer0_outputs(1680) <= 1'b1;
    layer0_outputs(1681) <= 1'b0;
    layer0_outputs(1682) <= a;
    layer0_outputs(1683) <= b;
    layer0_outputs(1684) <= a and b;
    layer0_outputs(1685) <= a and b;
    layer0_outputs(1686) <= not b;
    layer0_outputs(1687) <= a and b;
    layer0_outputs(1688) <= a and not b;
    layer0_outputs(1689) <= 1'b0;
    layer0_outputs(1690) <= not b or a;
    layer0_outputs(1691) <= 1'b1;
    layer0_outputs(1692) <= 1'b1;
    layer0_outputs(1693) <= not b;
    layer0_outputs(1694) <= a xor b;
    layer0_outputs(1695) <= not (a or b);
    layer0_outputs(1696) <= a or b;
    layer0_outputs(1697) <= not a or b;
    layer0_outputs(1698) <= a and not b;
    layer0_outputs(1699) <= b and not a;
    layer0_outputs(1700) <= 1'b1;
    layer0_outputs(1701) <= 1'b0;
    layer0_outputs(1702) <= not a;
    layer0_outputs(1703) <= not b or a;
    layer0_outputs(1704) <= a xor b;
    layer0_outputs(1705) <= 1'b1;
    layer0_outputs(1706) <= not a or b;
    layer0_outputs(1707) <= 1'b1;
    layer0_outputs(1708) <= b and not a;
    layer0_outputs(1709) <= not b;
    layer0_outputs(1710) <= 1'b0;
    layer0_outputs(1711) <= b and not a;
    layer0_outputs(1712) <= not b or a;
    layer0_outputs(1713) <= not (a xor b);
    layer0_outputs(1714) <= a or b;
    layer0_outputs(1715) <= 1'b0;
    layer0_outputs(1716) <= a and not b;
    layer0_outputs(1717) <= a and not b;
    layer0_outputs(1718) <= not b or a;
    layer0_outputs(1719) <= b and not a;
    layer0_outputs(1720) <= not (a or b);
    layer0_outputs(1721) <= not b;
    layer0_outputs(1722) <= 1'b1;
    layer0_outputs(1723) <= b;
    layer0_outputs(1724) <= not (a and b);
    layer0_outputs(1725) <= 1'b0;
    layer0_outputs(1726) <= not a or b;
    layer0_outputs(1727) <= not a or b;
    layer0_outputs(1728) <= a xor b;
    layer0_outputs(1729) <= a or b;
    layer0_outputs(1730) <= not a;
    layer0_outputs(1731) <= b and not a;
    layer0_outputs(1732) <= a or b;
    layer0_outputs(1733) <= not a or b;
    layer0_outputs(1734) <= 1'b0;
    layer0_outputs(1735) <= not a or b;
    layer0_outputs(1736) <= not b;
    layer0_outputs(1737) <= a and not b;
    layer0_outputs(1738) <= 1'b1;
    layer0_outputs(1739) <= not b or a;
    layer0_outputs(1740) <= not (a or b);
    layer0_outputs(1741) <= 1'b1;
    layer0_outputs(1742) <= not b or a;
    layer0_outputs(1743) <= a;
    layer0_outputs(1744) <= b;
    layer0_outputs(1745) <= not a;
    layer0_outputs(1746) <= not (a or b);
    layer0_outputs(1747) <= a and b;
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= 1'b0;
    layer0_outputs(1750) <= not a or b;
    layer0_outputs(1751) <= not (a or b);
    layer0_outputs(1752) <= 1'b0;
    layer0_outputs(1753) <= 1'b0;
    layer0_outputs(1754) <= b;
    layer0_outputs(1755) <= a;
    layer0_outputs(1756) <= b and not a;
    layer0_outputs(1757) <= a and b;
    layer0_outputs(1758) <= a;
    layer0_outputs(1759) <= a;
    layer0_outputs(1760) <= not (a or b);
    layer0_outputs(1761) <= b;
    layer0_outputs(1762) <= not b;
    layer0_outputs(1763) <= not b;
    layer0_outputs(1764) <= a or b;
    layer0_outputs(1765) <= not (a and b);
    layer0_outputs(1766) <= a xor b;
    layer0_outputs(1767) <= not b;
    layer0_outputs(1768) <= a and b;
    layer0_outputs(1769) <= a and b;
    layer0_outputs(1770) <= 1'b0;
    layer0_outputs(1771) <= not a or b;
    layer0_outputs(1772) <= a and not b;
    layer0_outputs(1773) <= a and b;
    layer0_outputs(1774) <= not (a and b);
    layer0_outputs(1775) <= a xor b;
    layer0_outputs(1776) <= a;
    layer0_outputs(1777) <= b and not a;
    layer0_outputs(1778) <= a;
    layer0_outputs(1779) <= not (a xor b);
    layer0_outputs(1780) <= a;
    layer0_outputs(1781) <= not a or b;
    layer0_outputs(1782) <= a xor b;
    layer0_outputs(1783) <= a;
    layer0_outputs(1784) <= 1'b0;
    layer0_outputs(1785) <= not (a or b);
    layer0_outputs(1786) <= not a;
    layer0_outputs(1787) <= 1'b1;
    layer0_outputs(1788) <= not a;
    layer0_outputs(1789) <= a and b;
    layer0_outputs(1790) <= not (a xor b);
    layer0_outputs(1791) <= a and b;
    layer0_outputs(1792) <= not (a and b);
    layer0_outputs(1793) <= 1'b1;
    layer0_outputs(1794) <= not a or b;
    layer0_outputs(1795) <= a and not b;
    layer0_outputs(1796) <= 1'b0;
    layer0_outputs(1797) <= not (a and b);
    layer0_outputs(1798) <= b;
    layer0_outputs(1799) <= b;
    layer0_outputs(1800) <= 1'b1;
    layer0_outputs(1801) <= not a or b;
    layer0_outputs(1802) <= not (a and b);
    layer0_outputs(1803) <= a and b;
    layer0_outputs(1804) <= a;
    layer0_outputs(1805) <= not (a and b);
    layer0_outputs(1806) <= not (a or b);
    layer0_outputs(1807) <= b;
    layer0_outputs(1808) <= not b;
    layer0_outputs(1809) <= a or b;
    layer0_outputs(1810) <= 1'b1;
    layer0_outputs(1811) <= not (a and b);
    layer0_outputs(1812) <= not (a or b);
    layer0_outputs(1813) <= not (a xor b);
    layer0_outputs(1814) <= not (a and b);
    layer0_outputs(1815) <= a and b;
    layer0_outputs(1816) <= not a or b;
    layer0_outputs(1817) <= a;
    layer0_outputs(1818) <= not a;
    layer0_outputs(1819) <= a xor b;
    layer0_outputs(1820) <= a;
    layer0_outputs(1821) <= not a or b;
    layer0_outputs(1822) <= b and not a;
    layer0_outputs(1823) <= b and not a;
    layer0_outputs(1824) <= not (a or b);
    layer0_outputs(1825) <= b;
    layer0_outputs(1826) <= a;
    layer0_outputs(1827) <= b;
    layer0_outputs(1828) <= 1'b0;
    layer0_outputs(1829) <= not a or b;
    layer0_outputs(1830) <= b and not a;
    layer0_outputs(1831) <= not (a xor b);
    layer0_outputs(1832) <= not a;
    layer0_outputs(1833) <= not (a and b);
    layer0_outputs(1834) <= not b;
    layer0_outputs(1835) <= a or b;
    layer0_outputs(1836) <= not b;
    layer0_outputs(1837) <= b;
    layer0_outputs(1838) <= not (a or b);
    layer0_outputs(1839) <= not (a and b);
    layer0_outputs(1840) <= b;
    layer0_outputs(1841) <= not a;
    layer0_outputs(1842) <= b and not a;
    layer0_outputs(1843) <= b;
    layer0_outputs(1844) <= a or b;
    layer0_outputs(1845) <= 1'b1;
    layer0_outputs(1846) <= a or b;
    layer0_outputs(1847) <= not (a or b);
    layer0_outputs(1848) <= a xor b;
    layer0_outputs(1849) <= b;
    layer0_outputs(1850) <= not (a xor b);
    layer0_outputs(1851) <= 1'b1;
    layer0_outputs(1852) <= a xor b;
    layer0_outputs(1853) <= a;
    layer0_outputs(1854) <= a and b;
    layer0_outputs(1855) <= not a or b;
    layer0_outputs(1856) <= a or b;
    layer0_outputs(1857) <= 1'b1;
    layer0_outputs(1858) <= not (a or b);
    layer0_outputs(1859) <= a xor b;
    layer0_outputs(1860) <= not (a or b);
    layer0_outputs(1861) <= a and not b;
    layer0_outputs(1862) <= not (a xor b);
    layer0_outputs(1863) <= a or b;
    layer0_outputs(1864) <= not (a and b);
    layer0_outputs(1865) <= not (a xor b);
    layer0_outputs(1866) <= not (a xor b);
    layer0_outputs(1867) <= not b;
    layer0_outputs(1868) <= not b or a;
    layer0_outputs(1869) <= not a;
    layer0_outputs(1870) <= a;
    layer0_outputs(1871) <= not b;
    layer0_outputs(1872) <= b;
    layer0_outputs(1873) <= b;
    layer0_outputs(1874) <= not a or b;
    layer0_outputs(1875) <= not (a or b);
    layer0_outputs(1876) <= not a;
    layer0_outputs(1877) <= a and b;
    layer0_outputs(1878) <= not (a and b);
    layer0_outputs(1879) <= b;
    layer0_outputs(1880) <= not a;
    layer0_outputs(1881) <= b and not a;
    layer0_outputs(1882) <= not a;
    layer0_outputs(1883) <= a and not b;
    layer0_outputs(1884) <= a xor b;
    layer0_outputs(1885) <= 1'b0;
    layer0_outputs(1886) <= 1'b1;
    layer0_outputs(1887) <= 1'b1;
    layer0_outputs(1888) <= not b;
    layer0_outputs(1889) <= b and not a;
    layer0_outputs(1890) <= 1'b1;
    layer0_outputs(1891) <= a;
    layer0_outputs(1892) <= not a;
    layer0_outputs(1893) <= 1'b0;
    layer0_outputs(1894) <= 1'b1;
    layer0_outputs(1895) <= a or b;
    layer0_outputs(1896) <= b and not a;
    layer0_outputs(1897) <= b and not a;
    layer0_outputs(1898) <= not a or b;
    layer0_outputs(1899) <= 1'b0;
    layer0_outputs(1900) <= not b or a;
    layer0_outputs(1901) <= a and not b;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= b and not a;
    layer0_outputs(1904) <= not b;
    layer0_outputs(1905) <= b;
    layer0_outputs(1906) <= b and not a;
    layer0_outputs(1907) <= b;
    layer0_outputs(1908) <= a;
    layer0_outputs(1909) <= 1'b0;
    layer0_outputs(1910) <= not b or a;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= a and b;
    layer0_outputs(1913) <= not (a or b);
    layer0_outputs(1914) <= not a or b;
    layer0_outputs(1915) <= a and not b;
    layer0_outputs(1916) <= a xor b;
    layer0_outputs(1917) <= 1'b1;
    layer0_outputs(1918) <= a;
    layer0_outputs(1919) <= a and b;
    layer0_outputs(1920) <= 1'b0;
    layer0_outputs(1921) <= not (a and b);
    layer0_outputs(1922) <= a;
    layer0_outputs(1923) <= not a or b;
    layer0_outputs(1924) <= not b or a;
    layer0_outputs(1925) <= b and not a;
    layer0_outputs(1926) <= a and b;
    layer0_outputs(1927) <= b;
    layer0_outputs(1928) <= 1'b0;
    layer0_outputs(1929) <= a and not b;
    layer0_outputs(1930) <= not a;
    layer0_outputs(1931) <= 1'b0;
    layer0_outputs(1932) <= a;
    layer0_outputs(1933) <= a and b;
    layer0_outputs(1934) <= not a or b;
    layer0_outputs(1935) <= a xor b;
    layer0_outputs(1936) <= a and b;
    layer0_outputs(1937) <= not (a and b);
    layer0_outputs(1938) <= b and not a;
    layer0_outputs(1939) <= not (a and b);
    layer0_outputs(1940) <= not (a or b);
    layer0_outputs(1941) <= not (a or b);
    layer0_outputs(1942) <= 1'b0;
    layer0_outputs(1943) <= not a;
    layer0_outputs(1944) <= 1'b1;
    layer0_outputs(1945) <= b and not a;
    layer0_outputs(1946) <= 1'b1;
    layer0_outputs(1947) <= 1'b1;
    layer0_outputs(1948) <= 1'b0;
    layer0_outputs(1949) <= 1'b1;
    layer0_outputs(1950) <= not (a and b);
    layer0_outputs(1951) <= a xor b;
    layer0_outputs(1952) <= not a;
    layer0_outputs(1953) <= not a;
    layer0_outputs(1954) <= not b;
    layer0_outputs(1955) <= not a or b;
    layer0_outputs(1956) <= not a;
    layer0_outputs(1957) <= not (a or b);
    layer0_outputs(1958) <= 1'b0;
    layer0_outputs(1959) <= not a;
    layer0_outputs(1960) <= a or b;
    layer0_outputs(1961) <= a and not b;
    layer0_outputs(1962) <= a and not b;
    layer0_outputs(1963) <= b;
    layer0_outputs(1964) <= not (a or b);
    layer0_outputs(1965) <= not (a and b);
    layer0_outputs(1966) <= b and not a;
    layer0_outputs(1967) <= a or b;
    layer0_outputs(1968) <= not b;
    layer0_outputs(1969) <= b;
    layer0_outputs(1970) <= not (a xor b);
    layer0_outputs(1971) <= not (a or b);
    layer0_outputs(1972) <= not (a or b);
    layer0_outputs(1973) <= b;
    layer0_outputs(1974) <= 1'b0;
    layer0_outputs(1975) <= a;
    layer0_outputs(1976) <= a and not b;
    layer0_outputs(1977) <= not b;
    layer0_outputs(1978) <= a and not b;
    layer0_outputs(1979) <= b;
    layer0_outputs(1980) <= a and not b;
    layer0_outputs(1981) <= not b;
    layer0_outputs(1982) <= not (a xor b);
    layer0_outputs(1983) <= not b or a;
    layer0_outputs(1984) <= b;
    layer0_outputs(1985) <= not a or b;
    layer0_outputs(1986) <= a and not b;
    layer0_outputs(1987) <= a and b;
    layer0_outputs(1988) <= a or b;
    layer0_outputs(1989) <= not b;
    layer0_outputs(1990) <= a;
    layer0_outputs(1991) <= a or b;
    layer0_outputs(1992) <= 1'b0;
    layer0_outputs(1993) <= not b or a;
    layer0_outputs(1994) <= a;
    layer0_outputs(1995) <= 1'b0;
    layer0_outputs(1996) <= not b or a;
    layer0_outputs(1997) <= a xor b;
    layer0_outputs(1998) <= not (a or b);
    layer0_outputs(1999) <= a and not b;
    layer0_outputs(2000) <= 1'b0;
    layer0_outputs(2001) <= b and not a;
    layer0_outputs(2002) <= a or b;
    layer0_outputs(2003) <= not (a or b);
    layer0_outputs(2004) <= not a;
    layer0_outputs(2005) <= 1'b1;
    layer0_outputs(2006) <= a and b;
    layer0_outputs(2007) <= not a;
    layer0_outputs(2008) <= a and b;
    layer0_outputs(2009) <= not (a or b);
    layer0_outputs(2010) <= a xor b;
    layer0_outputs(2011) <= not (a or b);
    layer0_outputs(2012) <= a and not b;
    layer0_outputs(2013) <= a;
    layer0_outputs(2014) <= a or b;
    layer0_outputs(2015) <= not (a or b);
    layer0_outputs(2016) <= not (a xor b);
    layer0_outputs(2017) <= a and b;
    layer0_outputs(2018) <= a or b;
    layer0_outputs(2019) <= 1'b0;
    layer0_outputs(2020) <= not a;
    layer0_outputs(2021) <= 1'b1;
    layer0_outputs(2022) <= a;
    layer0_outputs(2023) <= b and not a;
    layer0_outputs(2024) <= not (a or b);
    layer0_outputs(2025) <= b and not a;
    layer0_outputs(2026) <= not (a xor b);
    layer0_outputs(2027) <= b and not a;
    layer0_outputs(2028) <= 1'b0;
    layer0_outputs(2029) <= a;
    layer0_outputs(2030) <= not a;
    layer0_outputs(2031) <= a and not b;
    layer0_outputs(2032) <= not a;
    layer0_outputs(2033) <= a and b;
    layer0_outputs(2034) <= a;
    layer0_outputs(2035) <= not (a and b);
    layer0_outputs(2036) <= 1'b0;
    layer0_outputs(2037) <= b;
    layer0_outputs(2038) <= not (a xor b);
    layer0_outputs(2039) <= not b;
    layer0_outputs(2040) <= b;
    layer0_outputs(2041) <= 1'b1;
    layer0_outputs(2042) <= not a;
    layer0_outputs(2043) <= not a;
    layer0_outputs(2044) <= a and not b;
    layer0_outputs(2045) <= 1'b0;
    layer0_outputs(2046) <= not (a and b);
    layer0_outputs(2047) <= a and not b;
    layer0_outputs(2048) <= not a or b;
    layer0_outputs(2049) <= a and not b;
    layer0_outputs(2050) <= a and not b;
    layer0_outputs(2051) <= not a;
    layer0_outputs(2052) <= 1'b1;
    layer0_outputs(2053) <= a and not b;
    layer0_outputs(2054) <= a xor b;
    layer0_outputs(2055) <= not b;
    layer0_outputs(2056) <= b;
    layer0_outputs(2057) <= a and b;
    layer0_outputs(2058) <= 1'b0;
    layer0_outputs(2059) <= b and not a;
    layer0_outputs(2060) <= not a;
    layer0_outputs(2061) <= a and not b;
    layer0_outputs(2062) <= a and b;
    layer0_outputs(2063) <= not (a xor b);
    layer0_outputs(2064) <= not b;
    layer0_outputs(2065) <= a and not b;
    layer0_outputs(2066) <= a and not b;
    layer0_outputs(2067) <= a;
    layer0_outputs(2068) <= a and not b;
    layer0_outputs(2069) <= a;
    layer0_outputs(2070) <= a;
    layer0_outputs(2071) <= 1'b1;
    layer0_outputs(2072) <= a or b;
    layer0_outputs(2073) <= not a;
    layer0_outputs(2074) <= a and b;
    layer0_outputs(2075) <= not (a or b);
    layer0_outputs(2076) <= a;
    layer0_outputs(2077) <= a;
    layer0_outputs(2078) <= b;
    layer0_outputs(2079) <= a and not b;
    layer0_outputs(2080) <= not a or b;
    layer0_outputs(2081) <= not (a or b);
    layer0_outputs(2082) <= a or b;
    layer0_outputs(2083) <= not b;
    layer0_outputs(2084) <= not (a or b);
    layer0_outputs(2085) <= not (a or b);
    layer0_outputs(2086) <= 1'b1;
    layer0_outputs(2087) <= 1'b1;
    layer0_outputs(2088) <= a and not b;
    layer0_outputs(2089) <= not a;
    layer0_outputs(2090) <= 1'b0;
    layer0_outputs(2091) <= a and b;
    layer0_outputs(2092) <= a;
    layer0_outputs(2093) <= not (a or b);
    layer0_outputs(2094) <= a;
    layer0_outputs(2095) <= not a or b;
    layer0_outputs(2096) <= not a;
    layer0_outputs(2097) <= not a or b;
    layer0_outputs(2098) <= 1'b1;
    layer0_outputs(2099) <= a and not b;
    layer0_outputs(2100) <= a and b;
    layer0_outputs(2101) <= not (a and b);
    layer0_outputs(2102) <= a;
    layer0_outputs(2103) <= not (a or b);
    layer0_outputs(2104) <= not b or a;
    layer0_outputs(2105) <= not b;
    layer0_outputs(2106) <= not (a xor b);
    layer0_outputs(2107) <= not b;
    layer0_outputs(2108) <= 1'b0;
    layer0_outputs(2109) <= not a;
    layer0_outputs(2110) <= a or b;
    layer0_outputs(2111) <= not (a or b);
    layer0_outputs(2112) <= 1'b1;
    layer0_outputs(2113) <= not a or b;
    layer0_outputs(2114) <= a and not b;
    layer0_outputs(2115) <= a and b;
    layer0_outputs(2116) <= a and b;
    layer0_outputs(2117) <= b and not a;
    layer0_outputs(2118) <= b and not a;
    layer0_outputs(2119) <= not (a or b);
    layer0_outputs(2120) <= a;
    layer0_outputs(2121) <= not a or b;
    layer0_outputs(2122) <= a and not b;
    layer0_outputs(2123) <= a and b;
    layer0_outputs(2124) <= 1'b1;
    layer0_outputs(2125) <= not a;
    layer0_outputs(2126) <= b and not a;
    layer0_outputs(2127) <= not a or b;
    layer0_outputs(2128) <= not b;
    layer0_outputs(2129) <= not a;
    layer0_outputs(2130) <= b and not a;
    layer0_outputs(2131) <= a or b;
    layer0_outputs(2132) <= b and not a;
    layer0_outputs(2133) <= a;
    layer0_outputs(2134) <= a or b;
    layer0_outputs(2135) <= a;
    layer0_outputs(2136) <= not (a xor b);
    layer0_outputs(2137) <= not a or b;
    layer0_outputs(2138) <= not a;
    layer0_outputs(2139) <= a or b;
    layer0_outputs(2140) <= a and b;
    layer0_outputs(2141) <= 1'b0;
    layer0_outputs(2142) <= not a;
    layer0_outputs(2143) <= a or b;
    layer0_outputs(2144) <= 1'b1;
    layer0_outputs(2145) <= not b;
    layer0_outputs(2146) <= a and b;
    layer0_outputs(2147) <= not a;
    layer0_outputs(2148) <= 1'b1;
    layer0_outputs(2149) <= not (a and b);
    layer0_outputs(2150) <= b;
    layer0_outputs(2151) <= a;
    layer0_outputs(2152) <= not b or a;
    layer0_outputs(2153) <= not (a and b);
    layer0_outputs(2154) <= 1'b0;
    layer0_outputs(2155) <= a and not b;
    layer0_outputs(2156) <= 1'b1;
    layer0_outputs(2157) <= not b;
    layer0_outputs(2158) <= not b;
    layer0_outputs(2159) <= 1'b1;
    layer0_outputs(2160) <= 1'b0;
    layer0_outputs(2161) <= a and b;
    layer0_outputs(2162) <= b and not a;
    layer0_outputs(2163) <= 1'b1;
    layer0_outputs(2164) <= a and not b;
    layer0_outputs(2165) <= b;
    layer0_outputs(2166) <= not (a and b);
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= 1'b0;
    layer0_outputs(2169) <= not a;
    layer0_outputs(2170) <= not b;
    layer0_outputs(2171) <= 1'b0;
    layer0_outputs(2172) <= 1'b0;
    layer0_outputs(2173) <= not b;
    layer0_outputs(2174) <= a and not b;
    layer0_outputs(2175) <= not a;
    layer0_outputs(2176) <= 1'b1;
    layer0_outputs(2177) <= 1'b1;
    layer0_outputs(2178) <= not (a or b);
    layer0_outputs(2179) <= not a;
    layer0_outputs(2180) <= a;
    layer0_outputs(2181) <= a xor b;
    layer0_outputs(2182) <= 1'b0;
    layer0_outputs(2183) <= not b or a;
    layer0_outputs(2184) <= not b or a;
    layer0_outputs(2185) <= a or b;
    layer0_outputs(2186) <= b;
    layer0_outputs(2187) <= 1'b1;
    layer0_outputs(2188) <= a xor b;
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= not a;
    layer0_outputs(2191) <= not (a and b);
    layer0_outputs(2192) <= not (a xor b);
    layer0_outputs(2193) <= not b or a;
    layer0_outputs(2194) <= a and not b;
    layer0_outputs(2195) <= not (a and b);
    layer0_outputs(2196) <= a and not b;
    layer0_outputs(2197) <= a;
    layer0_outputs(2198) <= b and not a;
    layer0_outputs(2199) <= b and not a;
    layer0_outputs(2200) <= a and b;
    layer0_outputs(2201) <= not (a or b);
    layer0_outputs(2202) <= a and not b;
    layer0_outputs(2203) <= not a or b;
    layer0_outputs(2204) <= 1'b1;
    layer0_outputs(2205) <= a and not b;
    layer0_outputs(2206) <= b;
    layer0_outputs(2207) <= 1'b1;
    layer0_outputs(2208) <= not b or a;
    layer0_outputs(2209) <= a and not b;
    layer0_outputs(2210) <= not b or a;
    layer0_outputs(2211) <= a and b;
    layer0_outputs(2212) <= not a or b;
    layer0_outputs(2213) <= a and not b;
    layer0_outputs(2214) <= a and b;
    layer0_outputs(2215) <= a;
    layer0_outputs(2216) <= a xor b;
    layer0_outputs(2217) <= not a;
    layer0_outputs(2218) <= not a or b;
    layer0_outputs(2219) <= not (a or b);
    layer0_outputs(2220) <= a and not b;
    layer0_outputs(2221) <= a;
    layer0_outputs(2222) <= b and not a;
    layer0_outputs(2223) <= a and b;
    layer0_outputs(2224) <= a;
    layer0_outputs(2225) <= a and not b;
    layer0_outputs(2226) <= not b;
    layer0_outputs(2227) <= b and not a;
    layer0_outputs(2228) <= not b or a;
    layer0_outputs(2229) <= not b;
    layer0_outputs(2230) <= 1'b0;
    layer0_outputs(2231) <= b;
    layer0_outputs(2232) <= b;
    layer0_outputs(2233) <= b and not a;
    layer0_outputs(2234) <= a and b;
    layer0_outputs(2235) <= not (a and b);
    layer0_outputs(2236) <= not (a xor b);
    layer0_outputs(2237) <= not b or a;
    layer0_outputs(2238) <= 1'b0;
    layer0_outputs(2239) <= not b;
    layer0_outputs(2240) <= a and b;
    layer0_outputs(2241) <= a;
    layer0_outputs(2242) <= 1'b0;
    layer0_outputs(2243) <= a and b;
    layer0_outputs(2244) <= a or b;
    layer0_outputs(2245) <= a xor b;
    layer0_outputs(2246) <= b and not a;
    layer0_outputs(2247) <= b;
    layer0_outputs(2248) <= a or b;
    layer0_outputs(2249) <= 1'b0;
    layer0_outputs(2250) <= b;
    layer0_outputs(2251) <= a and b;
    layer0_outputs(2252) <= not (a and b);
    layer0_outputs(2253) <= not b or a;
    layer0_outputs(2254) <= not a or b;
    layer0_outputs(2255) <= b;
    layer0_outputs(2256) <= not (a and b);
    layer0_outputs(2257) <= not b;
    layer0_outputs(2258) <= a and not b;
    layer0_outputs(2259) <= 1'b1;
    layer0_outputs(2260) <= not (a and b);
    layer0_outputs(2261) <= 1'b1;
    layer0_outputs(2262) <= a and not b;
    layer0_outputs(2263) <= b;
    layer0_outputs(2264) <= not b;
    layer0_outputs(2265) <= b and not a;
    layer0_outputs(2266) <= not (a or b);
    layer0_outputs(2267) <= 1'b1;
    layer0_outputs(2268) <= b;
    layer0_outputs(2269) <= 1'b1;
    layer0_outputs(2270) <= a or b;
    layer0_outputs(2271) <= a and not b;
    layer0_outputs(2272) <= b;
    layer0_outputs(2273) <= 1'b0;
    layer0_outputs(2274) <= not b or a;
    layer0_outputs(2275) <= not a;
    layer0_outputs(2276) <= not b or a;
    layer0_outputs(2277) <= not (a xor b);
    layer0_outputs(2278) <= not (a xor b);
    layer0_outputs(2279) <= not (a or b);
    layer0_outputs(2280) <= a;
    layer0_outputs(2281) <= b;
    layer0_outputs(2282) <= not a;
    layer0_outputs(2283) <= not a;
    layer0_outputs(2284) <= not (a and b);
    layer0_outputs(2285) <= b and not a;
    layer0_outputs(2286) <= b;
    layer0_outputs(2287) <= b and not a;
    layer0_outputs(2288) <= not (a and b);
    layer0_outputs(2289) <= not (a or b);
    layer0_outputs(2290) <= not a or b;
    layer0_outputs(2291) <= b;
    layer0_outputs(2292) <= a and not b;
    layer0_outputs(2293) <= a or b;
    layer0_outputs(2294) <= not a or b;
    layer0_outputs(2295) <= not (a or b);
    layer0_outputs(2296) <= not b;
    layer0_outputs(2297) <= a and b;
    layer0_outputs(2298) <= a;
    layer0_outputs(2299) <= not a or b;
    layer0_outputs(2300) <= b and not a;
    layer0_outputs(2301) <= a or b;
    layer0_outputs(2302) <= not b;
    layer0_outputs(2303) <= a and not b;
    layer0_outputs(2304) <= 1'b0;
    layer0_outputs(2305) <= not a or b;
    layer0_outputs(2306) <= a and not b;
    layer0_outputs(2307) <= not (a or b);
    layer0_outputs(2308) <= 1'b1;
    layer0_outputs(2309) <= 1'b0;
    layer0_outputs(2310) <= a;
    layer0_outputs(2311) <= a or b;
    layer0_outputs(2312) <= not a or b;
    layer0_outputs(2313) <= not (a and b);
    layer0_outputs(2314) <= not (a or b);
    layer0_outputs(2315) <= 1'b0;
    layer0_outputs(2316) <= not (a and b);
    layer0_outputs(2317) <= not b;
    layer0_outputs(2318) <= a and b;
    layer0_outputs(2319) <= 1'b1;
    layer0_outputs(2320) <= a and b;
    layer0_outputs(2321) <= b and not a;
    layer0_outputs(2322) <= not (a or b);
    layer0_outputs(2323) <= not a or b;
    layer0_outputs(2324) <= 1'b1;
    layer0_outputs(2325) <= a and not b;
    layer0_outputs(2326) <= a and b;
    layer0_outputs(2327) <= not (a xor b);
    layer0_outputs(2328) <= not (a or b);
    layer0_outputs(2329) <= not b or a;
    layer0_outputs(2330) <= not b or a;
    layer0_outputs(2331) <= a and b;
    layer0_outputs(2332) <= b and not a;
    layer0_outputs(2333) <= a and not b;
    layer0_outputs(2334) <= a and b;
    layer0_outputs(2335) <= 1'b1;
    layer0_outputs(2336) <= not a;
    layer0_outputs(2337) <= not (a or b);
    layer0_outputs(2338) <= b;
    layer0_outputs(2339) <= 1'b1;
    layer0_outputs(2340) <= not (a and b);
    layer0_outputs(2341) <= a and not b;
    layer0_outputs(2342) <= not a;
    layer0_outputs(2343) <= 1'b0;
    layer0_outputs(2344) <= not a;
    layer0_outputs(2345) <= a;
    layer0_outputs(2346) <= b and not a;
    layer0_outputs(2347) <= a or b;
    layer0_outputs(2348) <= a and not b;
    layer0_outputs(2349) <= not b;
    layer0_outputs(2350) <= b and not a;
    layer0_outputs(2351) <= a or b;
    layer0_outputs(2352) <= a;
    layer0_outputs(2353) <= 1'b0;
    layer0_outputs(2354) <= not a;
    layer0_outputs(2355) <= not (a xor b);
    layer0_outputs(2356) <= not a or b;
    layer0_outputs(2357) <= not (a or b);
    layer0_outputs(2358) <= a or b;
    layer0_outputs(2359) <= 1'b0;
    layer0_outputs(2360) <= not (a or b);
    layer0_outputs(2361) <= not b or a;
    layer0_outputs(2362) <= a and b;
    layer0_outputs(2363) <= a and b;
    layer0_outputs(2364) <= 1'b1;
    layer0_outputs(2365) <= not b or a;
    layer0_outputs(2366) <= 1'b1;
    layer0_outputs(2367) <= b;
    layer0_outputs(2368) <= a xor b;
    layer0_outputs(2369) <= a xor b;
    layer0_outputs(2370) <= not b;
    layer0_outputs(2371) <= not (a and b);
    layer0_outputs(2372) <= a and b;
    layer0_outputs(2373) <= 1'b0;
    layer0_outputs(2374) <= b;
    layer0_outputs(2375) <= a xor b;
    layer0_outputs(2376) <= a;
    layer0_outputs(2377) <= not b;
    layer0_outputs(2378) <= not b or a;
    layer0_outputs(2379) <= not (a or b);
    layer0_outputs(2380) <= a and not b;
    layer0_outputs(2381) <= 1'b1;
    layer0_outputs(2382) <= not b;
    layer0_outputs(2383) <= b and not a;
    layer0_outputs(2384) <= b and not a;
    layer0_outputs(2385) <= not a or b;
    layer0_outputs(2386) <= a and b;
    layer0_outputs(2387) <= a;
    layer0_outputs(2388) <= a and not b;
    layer0_outputs(2389) <= not (a and b);
    layer0_outputs(2390) <= a and not b;
    layer0_outputs(2391) <= b and not a;
    layer0_outputs(2392) <= b and not a;
    layer0_outputs(2393) <= b and not a;
    layer0_outputs(2394) <= a or b;
    layer0_outputs(2395) <= not a;
    layer0_outputs(2396) <= not (a or b);
    layer0_outputs(2397) <= a;
    layer0_outputs(2398) <= not a or b;
    layer0_outputs(2399) <= not a;
    layer0_outputs(2400) <= a and not b;
    layer0_outputs(2401) <= not (a or b);
    layer0_outputs(2402) <= not (a or b);
    layer0_outputs(2403) <= a or b;
    layer0_outputs(2404) <= a or b;
    layer0_outputs(2405) <= not b or a;
    layer0_outputs(2406) <= b;
    layer0_outputs(2407) <= a;
    layer0_outputs(2408) <= not a;
    layer0_outputs(2409) <= a and b;
    layer0_outputs(2410) <= 1'b0;
    layer0_outputs(2411) <= not a or b;
    layer0_outputs(2412) <= not (a or b);
    layer0_outputs(2413) <= 1'b1;
    layer0_outputs(2414) <= 1'b0;
    layer0_outputs(2415) <= not (a or b);
    layer0_outputs(2416) <= 1'b0;
    layer0_outputs(2417) <= not a or b;
    layer0_outputs(2418) <= not (a and b);
    layer0_outputs(2419) <= not a or b;
    layer0_outputs(2420) <= not a;
    layer0_outputs(2421) <= a;
    layer0_outputs(2422) <= not b or a;
    layer0_outputs(2423) <= not (a or b);
    layer0_outputs(2424) <= not (a or b);
    layer0_outputs(2425) <= not a or b;
    layer0_outputs(2426) <= 1'b0;
    layer0_outputs(2427) <= 1'b1;
    layer0_outputs(2428) <= b and not a;
    layer0_outputs(2429) <= not (a and b);
    layer0_outputs(2430) <= not b or a;
    layer0_outputs(2431) <= a;
    layer0_outputs(2432) <= not a;
    layer0_outputs(2433) <= b;
    layer0_outputs(2434) <= b;
    layer0_outputs(2435) <= not b or a;
    layer0_outputs(2436) <= not (a and b);
    layer0_outputs(2437) <= not a;
    layer0_outputs(2438) <= a or b;
    layer0_outputs(2439) <= b;
    layer0_outputs(2440) <= not b or a;
    layer0_outputs(2441) <= not a;
    layer0_outputs(2442) <= not a;
    layer0_outputs(2443) <= 1'b0;
    layer0_outputs(2444) <= a and b;
    layer0_outputs(2445) <= b and not a;
    layer0_outputs(2446) <= not (a or b);
    layer0_outputs(2447) <= a xor b;
    layer0_outputs(2448) <= a xor b;
    layer0_outputs(2449) <= not b;
    layer0_outputs(2450) <= a and b;
    layer0_outputs(2451) <= not (a or b);
    layer0_outputs(2452) <= a;
    layer0_outputs(2453) <= a;
    layer0_outputs(2454) <= not a;
    layer0_outputs(2455) <= b;
    layer0_outputs(2456) <= a;
    layer0_outputs(2457) <= 1'b1;
    layer0_outputs(2458) <= b;
    layer0_outputs(2459) <= not a;
    layer0_outputs(2460) <= b and not a;
    layer0_outputs(2461) <= a or b;
    layer0_outputs(2462) <= a or b;
    layer0_outputs(2463) <= a or b;
    layer0_outputs(2464) <= not b;
    layer0_outputs(2465) <= not (a and b);
    layer0_outputs(2466) <= not a or b;
    layer0_outputs(2467) <= not a;
    layer0_outputs(2468) <= 1'b1;
    layer0_outputs(2469) <= a and b;
    layer0_outputs(2470) <= not b or a;
    layer0_outputs(2471) <= 1'b1;
    layer0_outputs(2472) <= 1'b1;
    layer0_outputs(2473) <= a;
    layer0_outputs(2474) <= b;
    layer0_outputs(2475) <= not a or b;
    layer0_outputs(2476) <= 1'b1;
    layer0_outputs(2477) <= not a;
    layer0_outputs(2478) <= not a or b;
    layer0_outputs(2479) <= not b;
    layer0_outputs(2480) <= 1'b0;
    layer0_outputs(2481) <= not (a and b);
    layer0_outputs(2482) <= a and not b;
    layer0_outputs(2483) <= not a;
    layer0_outputs(2484) <= b;
    layer0_outputs(2485) <= not b or a;
    layer0_outputs(2486) <= 1'b0;
    layer0_outputs(2487) <= not b;
    layer0_outputs(2488) <= b and not a;
    layer0_outputs(2489) <= not b or a;
    layer0_outputs(2490) <= a and b;
    layer0_outputs(2491) <= not a or b;
    layer0_outputs(2492) <= not b;
    layer0_outputs(2493) <= a and not b;
    layer0_outputs(2494) <= not a;
    layer0_outputs(2495) <= not b or a;
    layer0_outputs(2496) <= 1'b1;
    layer0_outputs(2497) <= not (a or b);
    layer0_outputs(2498) <= 1'b0;
    layer0_outputs(2499) <= b;
    layer0_outputs(2500) <= not b;
    layer0_outputs(2501) <= not a;
    layer0_outputs(2502) <= b;
    layer0_outputs(2503) <= a xor b;
    layer0_outputs(2504) <= not (a and b);
    layer0_outputs(2505) <= not (a and b);
    layer0_outputs(2506) <= a;
    layer0_outputs(2507) <= a;
    layer0_outputs(2508) <= not a or b;
    layer0_outputs(2509) <= not b or a;
    layer0_outputs(2510) <= 1'b0;
    layer0_outputs(2511) <= not (a and b);
    layer0_outputs(2512) <= not (a or b);
    layer0_outputs(2513) <= a and not b;
    layer0_outputs(2514) <= a xor b;
    layer0_outputs(2515) <= a;
    layer0_outputs(2516) <= not b;
    layer0_outputs(2517) <= not a or b;
    layer0_outputs(2518) <= a and b;
    layer0_outputs(2519) <= not a;
    layer0_outputs(2520) <= b;
    layer0_outputs(2521) <= a;
    layer0_outputs(2522) <= a or b;
    layer0_outputs(2523) <= a;
    layer0_outputs(2524) <= a;
    layer0_outputs(2525) <= not b or a;
    layer0_outputs(2526) <= not b or a;
    layer0_outputs(2527) <= 1'b1;
    layer0_outputs(2528) <= not b;
    layer0_outputs(2529) <= not a or b;
    layer0_outputs(2530) <= a and b;
    layer0_outputs(2531) <= not b or a;
    layer0_outputs(2532) <= not b;
    layer0_outputs(2533) <= not (a and b);
    layer0_outputs(2534) <= b;
    layer0_outputs(2535) <= 1'b0;
    layer0_outputs(2536) <= not a or b;
    layer0_outputs(2537) <= not b;
    layer0_outputs(2538) <= a;
    layer0_outputs(2539) <= not b;
    layer0_outputs(2540) <= b;
    layer0_outputs(2541) <= a;
    layer0_outputs(2542) <= a xor b;
    layer0_outputs(2543) <= a;
    layer0_outputs(2544) <= 1'b0;
    layer0_outputs(2545) <= a;
    layer0_outputs(2546) <= 1'b1;
    layer0_outputs(2547) <= 1'b0;
    layer0_outputs(2548) <= a or b;
    layer0_outputs(2549) <= 1'b0;
    layer0_outputs(2550) <= b;
    layer0_outputs(2551) <= not (a xor b);
    layer0_outputs(2552) <= a and b;
    layer0_outputs(2553) <= a and not b;
    layer0_outputs(2554) <= not a or b;
    layer0_outputs(2555) <= not b or a;
    layer0_outputs(2556) <= a and not b;
    layer0_outputs(2557) <= a and not b;
    layer0_outputs(2558) <= not (a xor b);
    layer0_outputs(2559) <= a or b;
    layer1_outputs(0) <= not b or a;
    layer1_outputs(1) <= not (a and b);
    layer1_outputs(2) <= not (a and b);
    layer1_outputs(3) <= 1'b1;
    layer1_outputs(4) <= a;
    layer1_outputs(5) <= not a or b;
    layer1_outputs(6) <= b and not a;
    layer1_outputs(7) <= b;
    layer1_outputs(8) <= a or b;
    layer1_outputs(9) <= not b;
    layer1_outputs(10) <= not b;
    layer1_outputs(11) <= not (a or b);
    layer1_outputs(12) <= 1'b0;
    layer1_outputs(13) <= not b or a;
    layer1_outputs(14) <= not a or b;
    layer1_outputs(15) <= not a or b;
    layer1_outputs(16) <= 1'b1;
    layer1_outputs(17) <= b and not a;
    layer1_outputs(18) <= 1'b0;
    layer1_outputs(19) <= 1'b0;
    layer1_outputs(20) <= a and b;
    layer1_outputs(21) <= b;
    layer1_outputs(22) <= a and b;
    layer1_outputs(23) <= not (a or b);
    layer1_outputs(24) <= not (a and b);
    layer1_outputs(25) <= a and not b;
    layer1_outputs(26) <= a or b;
    layer1_outputs(27) <= not (a or b);
    layer1_outputs(28) <= 1'b1;
    layer1_outputs(29) <= a;
    layer1_outputs(30) <= 1'b0;
    layer1_outputs(31) <= not b;
    layer1_outputs(32) <= a and not b;
    layer1_outputs(33) <= not a;
    layer1_outputs(34) <= not (a xor b);
    layer1_outputs(35) <= not (a xor b);
    layer1_outputs(36) <= a;
    layer1_outputs(37) <= a and not b;
    layer1_outputs(38) <= not a or b;
    layer1_outputs(39) <= not (a or b);
    layer1_outputs(40) <= not (a or b);
    layer1_outputs(41) <= a or b;
    layer1_outputs(42) <= b and not a;
    layer1_outputs(43) <= b;
    layer1_outputs(44) <= not b;
    layer1_outputs(45) <= a;
    layer1_outputs(46) <= b;
    layer1_outputs(47) <= 1'b1;
    layer1_outputs(48) <= a or b;
    layer1_outputs(49) <= not (a or b);
    layer1_outputs(50) <= a;
    layer1_outputs(51) <= not b or a;
    layer1_outputs(52) <= 1'b1;
    layer1_outputs(53) <= not a;
    layer1_outputs(54) <= 1'b0;
    layer1_outputs(55) <= a and not b;
    layer1_outputs(56) <= a and not b;
    layer1_outputs(57) <= not (a or b);
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= a;
    layer1_outputs(60) <= 1'b0;
    layer1_outputs(61) <= 1'b1;
    layer1_outputs(62) <= not b or a;
    layer1_outputs(63) <= 1'b1;
    layer1_outputs(64) <= 1'b0;
    layer1_outputs(65) <= a and b;
    layer1_outputs(66) <= a or b;
    layer1_outputs(67) <= not a;
    layer1_outputs(68) <= 1'b0;
    layer1_outputs(69) <= 1'b0;
    layer1_outputs(70) <= a and b;
    layer1_outputs(71) <= a or b;
    layer1_outputs(72) <= a;
    layer1_outputs(73) <= 1'b0;
    layer1_outputs(74) <= b and not a;
    layer1_outputs(75) <= b;
    layer1_outputs(76) <= a;
    layer1_outputs(77) <= not a;
    layer1_outputs(78) <= a and not b;
    layer1_outputs(79) <= b and not a;
    layer1_outputs(80) <= not (a or b);
    layer1_outputs(81) <= not b;
    layer1_outputs(82) <= 1'b0;
    layer1_outputs(83) <= 1'b0;
    layer1_outputs(84) <= b and not a;
    layer1_outputs(85) <= not (a or b);
    layer1_outputs(86) <= not b;
    layer1_outputs(87) <= not b;
    layer1_outputs(88) <= not b;
    layer1_outputs(89) <= not a or b;
    layer1_outputs(90) <= not b;
    layer1_outputs(91) <= a and not b;
    layer1_outputs(92) <= b;
    layer1_outputs(93) <= a and b;
    layer1_outputs(94) <= a or b;
    layer1_outputs(95) <= a and not b;
    layer1_outputs(96) <= a;
    layer1_outputs(97) <= not b or a;
    layer1_outputs(98) <= 1'b0;
    layer1_outputs(99) <= 1'b0;
    layer1_outputs(100) <= a and not b;
    layer1_outputs(101) <= not b;
    layer1_outputs(102) <= not a or b;
    layer1_outputs(103) <= a xor b;
    layer1_outputs(104) <= not b or a;
    layer1_outputs(105) <= a or b;
    layer1_outputs(106) <= not (a and b);
    layer1_outputs(107) <= 1'b1;
    layer1_outputs(108) <= not a;
    layer1_outputs(109) <= a or b;
    layer1_outputs(110) <= 1'b1;
    layer1_outputs(111) <= not (a or b);
    layer1_outputs(112) <= not b or a;
    layer1_outputs(113) <= 1'b1;
    layer1_outputs(114) <= a;
    layer1_outputs(115) <= not b or a;
    layer1_outputs(116) <= 1'b1;
    layer1_outputs(117) <= a or b;
    layer1_outputs(118) <= not (a or b);
    layer1_outputs(119) <= 1'b1;
    layer1_outputs(120) <= not (a or b);
    layer1_outputs(121) <= b and not a;
    layer1_outputs(122) <= a;
    layer1_outputs(123) <= 1'b0;
    layer1_outputs(124) <= not b or a;
    layer1_outputs(125) <= b and not a;
    layer1_outputs(126) <= 1'b1;
    layer1_outputs(127) <= not a;
    layer1_outputs(128) <= a or b;
    layer1_outputs(129) <= not a or b;
    layer1_outputs(130) <= a xor b;
    layer1_outputs(131) <= not (a and b);
    layer1_outputs(132) <= b;
    layer1_outputs(133) <= not a or b;
    layer1_outputs(134) <= not b or a;
    layer1_outputs(135) <= a and not b;
    layer1_outputs(136) <= 1'b0;
    layer1_outputs(137) <= 1'b1;
    layer1_outputs(138) <= b;
    layer1_outputs(139) <= 1'b1;
    layer1_outputs(140) <= not (a or b);
    layer1_outputs(141) <= b;
    layer1_outputs(142) <= a and b;
    layer1_outputs(143) <= not b;
    layer1_outputs(144) <= a and not b;
    layer1_outputs(145) <= 1'b1;
    layer1_outputs(146) <= 1'b0;
    layer1_outputs(147) <= not (a and b);
    layer1_outputs(148) <= not a or b;
    layer1_outputs(149) <= a and not b;
    layer1_outputs(150) <= not b or a;
    layer1_outputs(151) <= b and not a;
    layer1_outputs(152) <= a and b;
    layer1_outputs(153) <= b;
    layer1_outputs(154) <= b and not a;
    layer1_outputs(155) <= not b;
    layer1_outputs(156) <= not a;
    layer1_outputs(157) <= not b;
    layer1_outputs(158) <= 1'b1;
    layer1_outputs(159) <= 1'b0;
    layer1_outputs(160) <= a and b;
    layer1_outputs(161) <= not (a or b);
    layer1_outputs(162) <= 1'b1;
    layer1_outputs(163) <= b and not a;
    layer1_outputs(164) <= not (a xor b);
    layer1_outputs(165) <= 1'b1;
    layer1_outputs(166) <= a;
    layer1_outputs(167) <= 1'b0;
    layer1_outputs(168) <= not b or a;
    layer1_outputs(169) <= not a;
    layer1_outputs(170) <= not a or b;
    layer1_outputs(171) <= not (a or b);
    layer1_outputs(172) <= not b;
    layer1_outputs(173) <= a and not b;
    layer1_outputs(174) <= b and not a;
    layer1_outputs(175) <= not a or b;
    layer1_outputs(176) <= a or b;
    layer1_outputs(177) <= a;
    layer1_outputs(178) <= b;
    layer1_outputs(179) <= 1'b0;
    layer1_outputs(180) <= a and b;
    layer1_outputs(181) <= a or b;
    layer1_outputs(182) <= b;
    layer1_outputs(183) <= b;
    layer1_outputs(184) <= a or b;
    layer1_outputs(185) <= a and not b;
    layer1_outputs(186) <= 1'b0;
    layer1_outputs(187) <= a and not b;
    layer1_outputs(188) <= 1'b0;
    layer1_outputs(189) <= not a or b;
    layer1_outputs(190) <= not a;
    layer1_outputs(191) <= 1'b0;
    layer1_outputs(192) <= a and b;
    layer1_outputs(193) <= b;
    layer1_outputs(194) <= 1'b1;
    layer1_outputs(195) <= not a or b;
    layer1_outputs(196) <= a;
    layer1_outputs(197) <= 1'b0;
    layer1_outputs(198) <= a xor b;
    layer1_outputs(199) <= b and not a;
    layer1_outputs(200) <= a;
    layer1_outputs(201) <= a and b;
    layer1_outputs(202) <= not (a or b);
    layer1_outputs(203) <= 1'b1;
    layer1_outputs(204) <= a and not b;
    layer1_outputs(205) <= 1'b0;
    layer1_outputs(206) <= not (a and b);
    layer1_outputs(207) <= a or b;
    layer1_outputs(208) <= 1'b1;
    layer1_outputs(209) <= 1'b0;
    layer1_outputs(210) <= not (a and b);
    layer1_outputs(211) <= b;
    layer1_outputs(212) <= not (a or b);
    layer1_outputs(213) <= a or b;
    layer1_outputs(214) <= not (a or b);
    layer1_outputs(215) <= a;
    layer1_outputs(216) <= not b;
    layer1_outputs(217) <= b and not a;
    layer1_outputs(218) <= a;
    layer1_outputs(219) <= not (a and b);
    layer1_outputs(220) <= not (a or b);
    layer1_outputs(221) <= a and b;
    layer1_outputs(222) <= not b or a;
    layer1_outputs(223) <= a or b;
    layer1_outputs(224) <= not b or a;
    layer1_outputs(225) <= a and not b;
    layer1_outputs(226) <= not (a or b);
    layer1_outputs(227) <= b and not a;
    layer1_outputs(228) <= not a;
    layer1_outputs(229) <= 1'b0;
    layer1_outputs(230) <= not (a or b);
    layer1_outputs(231) <= not (a and b);
    layer1_outputs(232) <= a;
    layer1_outputs(233) <= 1'b0;
    layer1_outputs(234) <= a and not b;
    layer1_outputs(235) <= not (a and b);
    layer1_outputs(236) <= a and b;
    layer1_outputs(237) <= 1'b1;
    layer1_outputs(238) <= a;
    layer1_outputs(239) <= a and b;
    layer1_outputs(240) <= b;
    layer1_outputs(241) <= not b or a;
    layer1_outputs(242) <= b and not a;
    layer1_outputs(243) <= not a or b;
    layer1_outputs(244) <= not b or a;
    layer1_outputs(245) <= 1'b0;
    layer1_outputs(246) <= not (a or b);
    layer1_outputs(247) <= a and b;
    layer1_outputs(248) <= not a or b;
    layer1_outputs(249) <= not a;
    layer1_outputs(250) <= a and not b;
    layer1_outputs(251) <= not a;
    layer1_outputs(252) <= a and b;
    layer1_outputs(253) <= not (a and b);
    layer1_outputs(254) <= a;
    layer1_outputs(255) <= b;
    layer1_outputs(256) <= 1'b1;
    layer1_outputs(257) <= not a;
    layer1_outputs(258) <= 1'b1;
    layer1_outputs(259) <= 1'b0;
    layer1_outputs(260) <= not b or a;
    layer1_outputs(261) <= not (a and b);
    layer1_outputs(262) <= not (a or b);
    layer1_outputs(263) <= a;
    layer1_outputs(264) <= a;
    layer1_outputs(265) <= a or b;
    layer1_outputs(266) <= not a or b;
    layer1_outputs(267) <= b and not a;
    layer1_outputs(268) <= b;
    layer1_outputs(269) <= b and not a;
    layer1_outputs(270) <= 1'b1;
    layer1_outputs(271) <= not a or b;
    layer1_outputs(272) <= not b or a;
    layer1_outputs(273) <= a or b;
    layer1_outputs(274) <= a and not b;
    layer1_outputs(275) <= a and not b;
    layer1_outputs(276) <= not a;
    layer1_outputs(277) <= 1'b0;
    layer1_outputs(278) <= a and not b;
    layer1_outputs(279) <= b;
    layer1_outputs(280) <= not b;
    layer1_outputs(281) <= a and b;
    layer1_outputs(282) <= a and not b;
    layer1_outputs(283) <= not a or b;
    layer1_outputs(284) <= b and not a;
    layer1_outputs(285) <= a;
    layer1_outputs(286) <= not a or b;
    layer1_outputs(287) <= a and b;
    layer1_outputs(288) <= b;
    layer1_outputs(289) <= b;
    layer1_outputs(290) <= not a or b;
    layer1_outputs(291) <= a and not b;
    layer1_outputs(292) <= not (a or b);
    layer1_outputs(293) <= a and not b;
    layer1_outputs(294) <= not (a and b);
    layer1_outputs(295) <= a and b;
    layer1_outputs(296) <= b and not a;
    layer1_outputs(297) <= not (a and b);
    layer1_outputs(298) <= a and not b;
    layer1_outputs(299) <= b and not a;
    layer1_outputs(300) <= a and b;
    layer1_outputs(301) <= a and b;
    layer1_outputs(302) <= 1'b0;
    layer1_outputs(303) <= a or b;
    layer1_outputs(304) <= a and not b;
    layer1_outputs(305) <= a xor b;
    layer1_outputs(306) <= a or b;
    layer1_outputs(307) <= b and not a;
    layer1_outputs(308) <= b;
    layer1_outputs(309) <= a and not b;
    layer1_outputs(310) <= a or b;
    layer1_outputs(311) <= a and b;
    layer1_outputs(312) <= a and not b;
    layer1_outputs(313) <= 1'b1;
    layer1_outputs(314) <= not b;
    layer1_outputs(315) <= b;
    layer1_outputs(316) <= a and not b;
    layer1_outputs(317) <= not b;
    layer1_outputs(318) <= a and b;
    layer1_outputs(319) <= not (a or b);
    layer1_outputs(320) <= not a;
    layer1_outputs(321) <= not (a or b);
    layer1_outputs(322) <= not a;
    layer1_outputs(323) <= a;
    layer1_outputs(324) <= not a;
    layer1_outputs(325) <= 1'b1;
    layer1_outputs(326) <= a and b;
    layer1_outputs(327) <= 1'b1;
    layer1_outputs(328) <= a and b;
    layer1_outputs(329) <= b and not a;
    layer1_outputs(330) <= a and b;
    layer1_outputs(331) <= a or b;
    layer1_outputs(332) <= a or b;
    layer1_outputs(333) <= a and not b;
    layer1_outputs(334) <= a and b;
    layer1_outputs(335) <= a or b;
    layer1_outputs(336) <= 1'b1;
    layer1_outputs(337) <= b and not a;
    layer1_outputs(338) <= a or b;
    layer1_outputs(339) <= b and not a;
    layer1_outputs(340) <= 1'b1;
    layer1_outputs(341) <= b;
    layer1_outputs(342) <= not (a and b);
    layer1_outputs(343) <= a or b;
    layer1_outputs(344) <= 1'b1;
    layer1_outputs(345) <= not (a xor b);
    layer1_outputs(346) <= b and not a;
    layer1_outputs(347) <= 1'b0;
    layer1_outputs(348) <= b and not a;
    layer1_outputs(349) <= not (a or b);
    layer1_outputs(350) <= a and not b;
    layer1_outputs(351) <= 1'b0;
    layer1_outputs(352) <= not (a xor b);
    layer1_outputs(353) <= not (a and b);
    layer1_outputs(354) <= a;
    layer1_outputs(355) <= not b;
    layer1_outputs(356) <= b;
    layer1_outputs(357) <= not a or b;
    layer1_outputs(358) <= 1'b1;
    layer1_outputs(359) <= a;
    layer1_outputs(360) <= 1'b1;
    layer1_outputs(361) <= a or b;
    layer1_outputs(362) <= not b or a;
    layer1_outputs(363) <= a;
    layer1_outputs(364) <= not b;
    layer1_outputs(365) <= b;
    layer1_outputs(366) <= a or b;
    layer1_outputs(367) <= b and not a;
    layer1_outputs(368) <= not a;
    layer1_outputs(369) <= a or b;
    layer1_outputs(370) <= a and not b;
    layer1_outputs(371) <= not a or b;
    layer1_outputs(372) <= not a;
    layer1_outputs(373) <= b;
    layer1_outputs(374) <= 1'b0;
    layer1_outputs(375) <= not b;
    layer1_outputs(376) <= a;
    layer1_outputs(377) <= a or b;
    layer1_outputs(378) <= 1'b0;
    layer1_outputs(379) <= a or b;
    layer1_outputs(380) <= b;
    layer1_outputs(381) <= not b;
    layer1_outputs(382) <= not b or a;
    layer1_outputs(383) <= not (a or b);
    layer1_outputs(384) <= b;
    layer1_outputs(385) <= not a;
    layer1_outputs(386) <= not b or a;
    layer1_outputs(387) <= b and not a;
    layer1_outputs(388) <= b;
    layer1_outputs(389) <= a or b;
    layer1_outputs(390) <= not b or a;
    layer1_outputs(391) <= a and not b;
    layer1_outputs(392) <= 1'b0;
    layer1_outputs(393) <= not (a and b);
    layer1_outputs(394) <= not b or a;
    layer1_outputs(395) <= not (a or b);
    layer1_outputs(396) <= a and b;
    layer1_outputs(397) <= b and not a;
    layer1_outputs(398) <= 1'b0;
    layer1_outputs(399) <= not b;
    layer1_outputs(400) <= a and not b;
    layer1_outputs(401) <= not (a or b);
    layer1_outputs(402) <= 1'b1;
    layer1_outputs(403) <= 1'b0;
    layer1_outputs(404) <= a;
    layer1_outputs(405) <= 1'b1;
    layer1_outputs(406) <= 1'b0;
    layer1_outputs(407) <= b and not a;
    layer1_outputs(408) <= 1'b0;
    layer1_outputs(409) <= b;
    layer1_outputs(410) <= 1'b1;
    layer1_outputs(411) <= not (a or b);
    layer1_outputs(412) <= a and not b;
    layer1_outputs(413) <= a and b;
    layer1_outputs(414) <= not a;
    layer1_outputs(415) <= not b;
    layer1_outputs(416) <= not (a xor b);
    layer1_outputs(417) <= a;
    layer1_outputs(418) <= not b or a;
    layer1_outputs(419) <= a and not b;
    layer1_outputs(420) <= not b or a;
    layer1_outputs(421) <= not b;
    layer1_outputs(422) <= not a;
    layer1_outputs(423) <= not a;
    layer1_outputs(424) <= not a or b;
    layer1_outputs(425) <= 1'b1;
    layer1_outputs(426) <= not b;
    layer1_outputs(427) <= 1'b1;
    layer1_outputs(428) <= not b or a;
    layer1_outputs(429) <= not b;
    layer1_outputs(430) <= not (a xor b);
    layer1_outputs(431) <= not (a or b);
    layer1_outputs(432) <= 1'b0;
    layer1_outputs(433) <= b and not a;
    layer1_outputs(434) <= not a;
    layer1_outputs(435) <= 1'b1;
    layer1_outputs(436) <= b and not a;
    layer1_outputs(437) <= 1'b1;
    layer1_outputs(438) <= a and b;
    layer1_outputs(439) <= not (a and b);
    layer1_outputs(440) <= not (a and b);
    layer1_outputs(441) <= not (a and b);
    layer1_outputs(442) <= a;
    layer1_outputs(443) <= a xor b;
    layer1_outputs(444) <= not (a or b);
    layer1_outputs(445) <= 1'b1;
    layer1_outputs(446) <= a;
    layer1_outputs(447) <= a;
    layer1_outputs(448) <= not a or b;
    layer1_outputs(449) <= not (a or b);
    layer1_outputs(450) <= 1'b1;
    layer1_outputs(451) <= a and b;
    layer1_outputs(452) <= 1'b0;
    layer1_outputs(453) <= not a;
    layer1_outputs(454) <= not (a or b);
    layer1_outputs(455) <= b and not a;
    layer1_outputs(456) <= a and not b;
    layer1_outputs(457) <= not b;
    layer1_outputs(458) <= not a;
    layer1_outputs(459) <= not b;
    layer1_outputs(460) <= a and not b;
    layer1_outputs(461) <= not (a or b);
    layer1_outputs(462) <= not b or a;
    layer1_outputs(463) <= 1'b0;
    layer1_outputs(464) <= not b;
    layer1_outputs(465) <= a and not b;
    layer1_outputs(466) <= not b;
    layer1_outputs(467) <= 1'b0;
    layer1_outputs(468) <= not b or a;
    layer1_outputs(469) <= not b;
    layer1_outputs(470) <= a;
    layer1_outputs(471) <= a and not b;
    layer1_outputs(472) <= not (a or b);
    layer1_outputs(473) <= 1'b1;
    layer1_outputs(474) <= not (a and b);
    layer1_outputs(475) <= a or b;
    layer1_outputs(476) <= not b;
    layer1_outputs(477) <= a and b;
    layer1_outputs(478) <= 1'b0;
    layer1_outputs(479) <= a and b;
    layer1_outputs(480) <= b and not a;
    layer1_outputs(481) <= a and b;
    layer1_outputs(482) <= not (a and b);
    layer1_outputs(483) <= not a or b;
    layer1_outputs(484) <= not a;
    layer1_outputs(485) <= not b;
    layer1_outputs(486) <= not b or a;
    layer1_outputs(487) <= a;
    layer1_outputs(488) <= a xor b;
    layer1_outputs(489) <= not (a xor b);
    layer1_outputs(490) <= b;
    layer1_outputs(491) <= not a or b;
    layer1_outputs(492) <= not b;
    layer1_outputs(493) <= a and not b;
    layer1_outputs(494) <= a and not b;
    layer1_outputs(495) <= not a or b;
    layer1_outputs(496) <= not a;
    layer1_outputs(497) <= a;
    layer1_outputs(498) <= a;
    layer1_outputs(499) <= a or b;
    layer1_outputs(500) <= 1'b0;
    layer1_outputs(501) <= a and not b;
    layer1_outputs(502) <= not a;
    layer1_outputs(503) <= not b or a;
    layer1_outputs(504) <= b and not a;
    layer1_outputs(505) <= a and not b;
    layer1_outputs(506) <= not (a xor b);
    layer1_outputs(507) <= not b or a;
    layer1_outputs(508) <= a and not b;
    layer1_outputs(509) <= not (a xor b);
    layer1_outputs(510) <= not b;
    layer1_outputs(511) <= not b or a;
    layer1_outputs(512) <= 1'b0;
    layer1_outputs(513) <= not a or b;
    layer1_outputs(514) <= not b or a;
    layer1_outputs(515) <= not a;
    layer1_outputs(516) <= 1'b0;
    layer1_outputs(517) <= a;
    layer1_outputs(518) <= b and not a;
    layer1_outputs(519) <= a;
    layer1_outputs(520) <= not b or a;
    layer1_outputs(521) <= not a or b;
    layer1_outputs(522) <= not a or b;
    layer1_outputs(523) <= not b or a;
    layer1_outputs(524) <= not (a or b);
    layer1_outputs(525) <= not (a and b);
    layer1_outputs(526) <= not b or a;
    layer1_outputs(527) <= not (a and b);
    layer1_outputs(528) <= not b;
    layer1_outputs(529) <= not b;
    layer1_outputs(530) <= not b;
    layer1_outputs(531) <= not (a or b);
    layer1_outputs(532) <= not (a or b);
    layer1_outputs(533) <= 1'b0;
    layer1_outputs(534) <= 1'b1;
    layer1_outputs(535) <= not (a and b);
    layer1_outputs(536) <= not b or a;
    layer1_outputs(537) <= not (a or b);
    layer1_outputs(538) <= not (a and b);
    layer1_outputs(539) <= 1'b0;
    layer1_outputs(540) <= not a or b;
    layer1_outputs(541) <= not (a and b);
    layer1_outputs(542) <= 1'b1;
    layer1_outputs(543) <= 1'b1;
    layer1_outputs(544) <= 1'b0;
    layer1_outputs(545) <= a xor b;
    layer1_outputs(546) <= b and not a;
    layer1_outputs(547) <= a and b;
    layer1_outputs(548) <= b;
    layer1_outputs(549) <= not a or b;
    layer1_outputs(550) <= 1'b0;
    layer1_outputs(551) <= a or b;
    layer1_outputs(552) <= a and b;
    layer1_outputs(553) <= not a or b;
    layer1_outputs(554) <= not (a xor b);
    layer1_outputs(555) <= a or b;
    layer1_outputs(556) <= not (a and b);
    layer1_outputs(557) <= 1'b1;
    layer1_outputs(558) <= 1'b1;
    layer1_outputs(559) <= b and not a;
    layer1_outputs(560) <= a and not b;
    layer1_outputs(561) <= a;
    layer1_outputs(562) <= not (a and b);
    layer1_outputs(563) <= not b;
    layer1_outputs(564) <= not (a and b);
    layer1_outputs(565) <= not a;
    layer1_outputs(566) <= a and not b;
    layer1_outputs(567) <= 1'b0;
    layer1_outputs(568) <= 1'b1;
    layer1_outputs(569) <= a;
    layer1_outputs(570) <= b and not a;
    layer1_outputs(571) <= not b;
    layer1_outputs(572) <= a xor b;
    layer1_outputs(573) <= not a or b;
    layer1_outputs(574) <= 1'b1;
    layer1_outputs(575) <= a;
    layer1_outputs(576) <= not (a or b);
    layer1_outputs(577) <= 1'b0;
    layer1_outputs(578) <= not b or a;
    layer1_outputs(579) <= 1'b1;
    layer1_outputs(580) <= 1'b1;
    layer1_outputs(581) <= not (a or b);
    layer1_outputs(582) <= a and b;
    layer1_outputs(583) <= a and not b;
    layer1_outputs(584) <= not b;
    layer1_outputs(585) <= not (a or b);
    layer1_outputs(586) <= not (a and b);
    layer1_outputs(587) <= not b or a;
    layer1_outputs(588) <= b;
    layer1_outputs(589) <= a and not b;
    layer1_outputs(590) <= not (a and b);
    layer1_outputs(591) <= not b or a;
    layer1_outputs(592) <= a or b;
    layer1_outputs(593) <= not a or b;
    layer1_outputs(594) <= a and not b;
    layer1_outputs(595) <= b and not a;
    layer1_outputs(596) <= b;
    layer1_outputs(597) <= not b or a;
    layer1_outputs(598) <= b and not a;
    layer1_outputs(599) <= not a;
    layer1_outputs(600) <= not (a and b);
    layer1_outputs(601) <= not (a and b);
    layer1_outputs(602) <= a xor b;
    layer1_outputs(603) <= b;
    layer1_outputs(604) <= not a;
    layer1_outputs(605) <= 1'b1;
    layer1_outputs(606) <= a and not b;
    layer1_outputs(607) <= b;
    layer1_outputs(608) <= b and not a;
    layer1_outputs(609) <= a and b;
    layer1_outputs(610) <= a or b;
    layer1_outputs(611) <= not a or b;
    layer1_outputs(612) <= not a or b;
    layer1_outputs(613) <= b;
    layer1_outputs(614) <= 1'b0;
    layer1_outputs(615) <= a and b;
    layer1_outputs(616) <= not (a and b);
    layer1_outputs(617) <= not b;
    layer1_outputs(618) <= not b;
    layer1_outputs(619) <= 1'b1;
    layer1_outputs(620) <= b;
    layer1_outputs(621) <= b and not a;
    layer1_outputs(622) <= b;
    layer1_outputs(623) <= a and not b;
    layer1_outputs(624) <= b and not a;
    layer1_outputs(625) <= not (a xor b);
    layer1_outputs(626) <= 1'b1;
    layer1_outputs(627) <= 1'b0;
    layer1_outputs(628) <= not b or a;
    layer1_outputs(629) <= a and not b;
    layer1_outputs(630) <= 1'b1;
    layer1_outputs(631) <= a or b;
    layer1_outputs(632) <= 1'b0;
    layer1_outputs(633) <= 1'b1;
    layer1_outputs(634) <= a and b;
    layer1_outputs(635) <= a and b;
    layer1_outputs(636) <= not (a and b);
    layer1_outputs(637) <= a;
    layer1_outputs(638) <= a or b;
    layer1_outputs(639) <= not a;
    layer1_outputs(640) <= a and b;
    layer1_outputs(641) <= not (a or b);
    layer1_outputs(642) <= 1'b0;
    layer1_outputs(643) <= not a or b;
    layer1_outputs(644) <= 1'b0;
    layer1_outputs(645) <= a or b;
    layer1_outputs(646) <= not a;
    layer1_outputs(647) <= not (a and b);
    layer1_outputs(648) <= a and not b;
    layer1_outputs(649) <= 1'b0;
    layer1_outputs(650) <= b and not a;
    layer1_outputs(651) <= a and b;
    layer1_outputs(652) <= 1'b0;
    layer1_outputs(653) <= not b or a;
    layer1_outputs(654) <= b;
    layer1_outputs(655) <= a xor b;
    layer1_outputs(656) <= b and not a;
    layer1_outputs(657) <= a and not b;
    layer1_outputs(658) <= not (a and b);
    layer1_outputs(659) <= a or b;
    layer1_outputs(660) <= not b;
    layer1_outputs(661) <= a and b;
    layer1_outputs(662) <= b;
    layer1_outputs(663) <= 1'b1;
    layer1_outputs(664) <= a and b;
    layer1_outputs(665) <= b and not a;
    layer1_outputs(666) <= b;
    layer1_outputs(667) <= not b or a;
    layer1_outputs(668) <= a;
    layer1_outputs(669) <= not b;
    layer1_outputs(670) <= not a or b;
    layer1_outputs(671) <= 1'b0;
    layer1_outputs(672) <= b;
    layer1_outputs(673) <= b;
    layer1_outputs(674) <= 1'b0;
    layer1_outputs(675) <= a or b;
    layer1_outputs(676) <= b and not a;
    layer1_outputs(677) <= 1'b1;
    layer1_outputs(678) <= a or b;
    layer1_outputs(679) <= 1'b1;
    layer1_outputs(680) <= not (a and b);
    layer1_outputs(681) <= a and b;
    layer1_outputs(682) <= not b;
    layer1_outputs(683) <= not a;
    layer1_outputs(684) <= a and not b;
    layer1_outputs(685) <= not (a or b);
    layer1_outputs(686) <= not a or b;
    layer1_outputs(687) <= not b;
    layer1_outputs(688) <= not a;
    layer1_outputs(689) <= not (a and b);
    layer1_outputs(690) <= 1'b1;
    layer1_outputs(691) <= not b;
    layer1_outputs(692) <= not b or a;
    layer1_outputs(693) <= a and b;
    layer1_outputs(694) <= 1'b1;
    layer1_outputs(695) <= b;
    layer1_outputs(696) <= not (a xor b);
    layer1_outputs(697) <= not (a and b);
    layer1_outputs(698) <= 1'b0;
    layer1_outputs(699) <= not a;
    layer1_outputs(700) <= a and b;
    layer1_outputs(701) <= 1'b0;
    layer1_outputs(702) <= not a;
    layer1_outputs(703) <= b and not a;
    layer1_outputs(704) <= not (a and b);
    layer1_outputs(705) <= not (a xor b);
    layer1_outputs(706) <= not (a or b);
    layer1_outputs(707) <= not a or b;
    layer1_outputs(708) <= a or b;
    layer1_outputs(709) <= 1'b0;
    layer1_outputs(710) <= not b or a;
    layer1_outputs(711) <= b;
    layer1_outputs(712) <= b and not a;
    layer1_outputs(713) <= 1'b0;
    layer1_outputs(714) <= a;
    layer1_outputs(715) <= 1'b0;
    layer1_outputs(716) <= a or b;
    layer1_outputs(717) <= 1'b0;
    layer1_outputs(718) <= not a;
    layer1_outputs(719) <= a or b;
    layer1_outputs(720) <= 1'b0;
    layer1_outputs(721) <= 1'b0;
    layer1_outputs(722) <= 1'b0;
    layer1_outputs(723) <= not (a or b);
    layer1_outputs(724) <= not b or a;
    layer1_outputs(725) <= not b or a;
    layer1_outputs(726) <= not a or b;
    layer1_outputs(727) <= 1'b1;
    layer1_outputs(728) <= not b or a;
    layer1_outputs(729) <= b;
    layer1_outputs(730) <= not b;
    layer1_outputs(731) <= a;
    layer1_outputs(732) <= not b or a;
    layer1_outputs(733) <= not (a or b);
    layer1_outputs(734) <= not (a and b);
    layer1_outputs(735) <= not a;
    layer1_outputs(736) <= a and b;
    layer1_outputs(737) <= b and not a;
    layer1_outputs(738) <= not a or b;
    layer1_outputs(739) <= not a or b;
    layer1_outputs(740) <= a and b;
    layer1_outputs(741) <= not a or b;
    layer1_outputs(742) <= not a or b;
    layer1_outputs(743) <= not a or b;
    layer1_outputs(744) <= 1'b0;
    layer1_outputs(745) <= 1'b0;
    layer1_outputs(746) <= 1'b1;
    layer1_outputs(747) <= not (a xor b);
    layer1_outputs(748) <= b and not a;
    layer1_outputs(749) <= a or b;
    layer1_outputs(750) <= not (a or b);
    layer1_outputs(751) <= 1'b1;
    layer1_outputs(752) <= b;
    layer1_outputs(753) <= 1'b0;
    layer1_outputs(754) <= 1'b0;
    layer1_outputs(755) <= not a;
    layer1_outputs(756) <= not a or b;
    layer1_outputs(757) <= not b or a;
    layer1_outputs(758) <= a and b;
    layer1_outputs(759) <= a and not b;
    layer1_outputs(760) <= b and not a;
    layer1_outputs(761) <= 1'b1;
    layer1_outputs(762) <= not b or a;
    layer1_outputs(763) <= a and b;
    layer1_outputs(764) <= a;
    layer1_outputs(765) <= not a or b;
    layer1_outputs(766) <= not (a or b);
    layer1_outputs(767) <= 1'b0;
    layer1_outputs(768) <= a and b;
    layer1_outputs(769) <= not b or a;
    layer1_outputs(770) <= not (a and b);
    layer1_outputs(771) <= not (a and b);
    layer1_outputs(772) <= 1'b1;
    layer1_outputs(773) <= not (a or b);
    layer1_outputs(774) <= b;
    layer1_outputs(775) <= not a;
    layer1_outputs(776) <= not b;
    layer1_outputs(777) <= not b or a;
    layer1_outputs(778) <= a and not b;
    layer1_outputs(779) <= not (a and b);
    layer1_outputs(780) <= 1'b0;
    layer1_outputs(781) <= 1'b0;
    layer1_outputs(782) <= a;
    layer1_outputs(783) <= a xor b;
    layer1_outputs(784) <= a xor b;
    layer1_outputs(785) <= b;
    layer1_outputs(786) <= 1'b0;
    layer1_outputs(787) <= not (a or b);
    layer1_outputs(788) <= b and not a;
    layer1_outputs(789) <= a or b;
    layer1_outputs(790) <= b and not a;
    layer1_outputs(791) <= b;
    layer1_outputs(792) <= not b or a;
    layer1_outputs(793) <= not a or b;
    layer1_outputs(794) <= a and not b;
    layer1_outputs(795) <= 1'b0;
    layer1_outputs(796) <= a and not b;
    layer1_outputs(797) <= not b;
    layer1_outputs(798) <= not (a xor b);
    layer1_outputs(799) <= not b or a;
    layer1_outputs(800) <= 1'b0;
    layer1_outputs(801) <= 1'b1;
    layer1_outputs(802) <= 1'b0;
    layer1_outputs(803) <= not a;
    layer1_outputs(804) <= a and not b;
    layer1_outputs(805) <= not (a and b);
    layer1_outputs(806) <= not b or a;
    layer1_outputs(807) <= not (a and b);
    layer1_outputs(808) <= b;
    layer1_outputs(809) <= not (a and b);
    layer1_outputs(810) <= not (a or b);
    layer1_outputs(811) <= a xor b;
    layer1_outputs(812) <= not a or b;
    layer1_outputs(813) <= a;
    layer1_outputs(814) <= a and not b;
    layer1_outputs(815) <= not (a xor b);
    layer1_outputs(816) <= a;
    layer1_outputs(817) <= not (a and b);
    layer1_outputs(818) <= 1'b1;
    layer1_outputs(819) <= not a or b;
    layer1_outputs(820) <= 1'b1;
    layer1_outputs(821) <= a or b;
    layer1_outputs(822) <= not (a and b);
    layer1_outputs(823) <= not (a and b);
    layer1_outputs(824) <= a xor b;
    layer1_outputs(825) <= not b;
    layer1_outputs(826) <= a and not b;
    layer1_outputs(827) <= not b or a;
    layer1_outputs(828) <= not a;
    layer1_outputs(829) <= not a;
    layer1_outputs(830) <= b and not a;
    layer1_outputs(831) <= not b;
    layer1_outputs(832) <= a or b;
    layer1_outputs(833) <= not (a and b);
    layer1_outputs(834) <= a and not b;
    layer1_outputs(835) <= not (a and b);
    layer1_outputs(836) <= a and b;
    layer1_outputs(837) <= not b or a;
    layer1_outputs(838) <= not (a or b);
    layer1_outputs(839) <= a and not b;
    layer1_outputs(840) <= 1'b0;
    layer1_outputs(841) <= a and b;
    layer1_outputs(842) <= 1'b0;
    layer1_outputs(843) <= a or b;
    layer1_outputs(844) <= not b;
    layer1_outputs(845) <= not a or b;
    layer1_outputs(846) <= 1'b1;
    layer1_outputs(847) <= b;
    layer1_outputs(848) <= not (a and b);
    layer1_outputs(849) <= b;
    layer1_outputs(850) <= a;
    layer1_outputs(851) <= not (a or b);
    layer1_outputs(852) <= b;
    layer1_outputs(853) <= not b;
    layer1_outputs(854) <= a and not b;
    layer1_outputs(855) <= a and b;
    layer1_outputs(856) <= a and not b;
    layer1_outputs(857) <= a and not b;
    layer1_outputs(858) <= not a or b;
    layer1_outputs(859) <= a or b;
    layer1_outputs(860) <= 1'b1;
    layer1_outputs(861) <= a;
    layer1_outputs(862) <= b and not a;
    layer1_outputs(863) <= a;
    layer1_outputs(864) <= a and not b;
    layer1_outputs(865) <= a and not b;
    layer1_outputs(866) <= 1'b0;
    layer1_outputs(867) <= b;
    layer1_outputs(868) <= b;
    layer1_outputs(869) <= 1'b0;
    layer1_outputs(870) <= 1'b0;
    layer1_outputs(871) <= a and b;
    layer1_outputs(872) <= a and not b;
    layer1_outputs(873) <= a;
    layer1_outputs(874) <= a;
    layer1_outputs(875) <= b and not a;
    layer1_outputs(876) <= a and not b;
    layer1_outputs(877) <= a or b;
    layer1_outputs(878) <= not (a and b);
    layer1_outputs(879) <= not (a xor b);
    layer1_outputs(880) <= a and b;
    layer1_outputs(881) <= a or b;
    layer1_outputs(882) <= a;
    layer1_outputs(883) <= not a or b;
    layer1_outputs(884) <= not a or b;
    layer1_outputs(885) <= 1'b1;
    layer1_outputs(886) <= not b;
    layer1_outputs(887) <= not b;
    layer1_outputs(888) <= not b or a;
    layer1_outputs(889) <= not (a or b);
    layer1_outputs(890) <= not b or a;
    layer1_outputs(891) <= b and not a;
    layer1_outputs(892) <= not a or b;
    layer1_outputs(893) <= b and not a;
    layer1_outputs(894) <= b and not a;
    layer1_outputs(895) <= not (a and b);
    layer1_outputs(896) <= not a;
    layer1_outputs(897) <= not (a and b);
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= a;
    layer1_outputs(900) <= 1'b1;
    layer1_outputs(901) <= 1'b1;
    layer1_outputs(902) <= not a;
    layer1_outputs(903) <= 1'b1;
    layer1_outputs(904) <= not (a or b);
    layer1_outputs(905) <= not a or b;
    layer1_outputs(906) <= not (a and b);
    layer1_outputs(907) <= 1'b0;
    layer1_outputs(908) <= b;
    layer1_outputs(909) <= a and not b;
    layer1_outputs(910) <= a;
    layer1_outputs(911) <= not (a and b);
    layer1_outputs(912) <= 1'b1;
    layer1_outputs(913) <= not b;
    layer1_outputs(914) <= not (a xor b);
    layer1_outputs(915) <= not a;
    layer1_outputs(916) <= 1'b0;
    layer1_outputs(917) <= a xor b;
    layer1_outputs(918) <= not b or a;
    layer1_outputs(919) <= not (a or b);
    layer1_outputs(920) <= not b or a;
    layer1_outputs(921) <= not a or b;
    layer1_outputs(922) <= not (a or b);
    layer1_outputs(923) <= b and not a;
    layer1_outputs(924) <= not a;
    layer1_outputs(925) <= b;
    layer1_outputs(926) <= a;
    layer1_outputs(927) <= 1'b0;
    layer1_outputs(928) <= 1'b1;
    layer1_outputs(929) <= not (a or b);
    layer1_outputs(930) <= 1'b0;
    layer1_outputs(931) <= 1'b0;
    layer1_outputs(932) <= a or b;
    layer1_outputs(933) <= 1'b0;
    layer1_outputs(934) <= a and not b;
    layer1_outputs(935) <= a and not b;
    layer1_outputs(936) <= not (a and b);
    layer1_outputs(937) <= a;
    layer1_outputs(938) <= not a or b;
    layer1_outputs(939) <= not (a and b);
    layer1_outputs(940) <= a and b;
    layer1_outputs(941) <= b and not a;
    layer1_outputs(942) <= not a;
    layer1_outputs(943) <= a or b;
    layer1_outputs(944) <= not b or a;
    layer1_outputs(945) <= a and not b;
    layer1_outputs(946) <= 1'b0;
    layer1_outputs(947) <= 1'b1;
    layer1_outputs(948) <= a and b;
    layer1_outputs(949) <= 1'b1;
    layer1_outputs(950) <= not b;
    layer1_outputs(951) <= 1'b0;
    layer1_outputs(952) <= not b;
    layer1_outputs(953) <= not a;
    layer1_outputs(954) <= not b or a;
    layer1_outputs(955) <= 1'b0;
    layer1_outputs(956) <= a or b;
    layer1_outputs(957) <= a and b;
    layer1_outputs(958) <= 1'b0;
    layer1_outputs(959) <= a and not b;
    layer1_outputs(960) <= not (a or b);
    layer1_outputs(961) <= a and b;
    layer1_outputs(962) <= not b or a;
    layer1_outputs(963) <= a and b;
    layer1_outputs(964) <= not a or b;
    layer1_outputs(965) <= a or b;
    layer1_outputs(966) <= not b;
    layer1_outputs(967) <= b and not a;
    layer1_outputs(968) <= not b;
    layer1_outputs(969) <= b;
    layer1_outputs(970) <= a and not b;
    layer1_outputs(971) <= b;
    layer1_outputs(972) <= not (a and b);
    layer1_outputs(973) <= not a;
    layer1_outputs(974) <= a or b;
    layer1_outputs(975) <= a and b;
    layer1_outputs(976) <= a or b;
    layer1_outputs(977) <= b;
    layer1_outputs(978) <= not a;
    layer1_outputs(979) <= a or b;
    layer1_outputs(980) <= not b or a;
    layer1_outputs(981) <= not b;
    layer1_outputs(982) <= not a;
    layer1_outputs(983) <= not a;
    layer1_outputs(984) <= 1'b0;
    layer1_outputs(985) <= a or b;
    layer1_outputs(986) <= a and not b;
    layer1_outputs(987) <= not a or b;
    layer1_outputs(988) <= 1'b0;
    layer1_outputs(989) <= a or b;
    layer1_outputs(990) <= a;
    layer1_outputs(991) <= not a or b;
    layer1_outputs(992) <= not (a and b);
    layer1_outputs(993) <= b;
    layer1_outputs(994) <= a;
    layer1_outputs(995) <= a or b;
    layer1_outputs(996) <= b and not a;
    layer1_outputs(997) <= a or b;
    layer1_outputs(998) <= not a;
    layer1_outputs(999) <= not (a or b);
    layer1_outputs(1000) <= a and not b;
    layer1_outputs(1001) <= a or b;
    layer1_outputs(1002) <= not (a and b);
    layer1_outputs(1003) <= not (a or b);
    layer1_outputs(1004) <= a or b;
    layer1_outputs(1005) <= 1'b1;
    layer1_outputs(1006) <= not (a xor b);
    layer1_outputs(1007) <= not a or b;
    layer1_outputs(1008) <= 1'b1;
    layer1_outputs(1009) <= not (a and b);
    layer1_outputs(1010) <= 1'b0;
    layer1_outputs(1011) <= a or b;
    layer1_outputs(1012) <= a xor b;
    layer1_outputs(1013) <= 1'b0;
    layer1_outputs(1014) <= not a;
    layer1_outputs(1015) <= b and not a;
    layer1_outputs(1016) <= not (a and b);
    layer1_outputs(1017) <= not (a and b);
    layer1_outputs(1018) <= 1'b1;
    layer1_outputs(1019) <= not b or a;
    layer1_outputs(1020) <= not a;
    layer1_outputs(1021) <= a or b;
    layer1_outputs(1022) <= b and not a;
    layer1_outputs(1023) <= not a;
    layer1_outputs(1024) <= a or b;
    layer1_outputs(1025) <= b and not a;
    layer1_outputs(1026) <= not b or a;
    layer1_outputs(1027) <= not (a and b);
    layer1_outputs(1028) <= not (a or b);
    layer1_outputs(1029) <= a and b;
    layer1_outputs(1030) <= not a;
    layer1_outputs(1031) <= 1'b0;
    layer1_outputs(1032) <= not b;
    layer1_outputs(1033) <= not a;
    layer1_outputs(1034) <= 1'b0;
    layer1_outputs(1035) <= not a;
    layer1_outputs(1036) <= a and not b;
    layer1_outputs(1037) <= a or b;
    layer1_outputs(1038) <= not (a or b);
    layer1_outputs(1039) <= 1'b0;
    layer1_outputs(1040) <= 1'b1;
    layer1_outputs(1041) <= 1'b1;
    layer1_outputs(1042) <= not b or a;
    layer1_outputs(1043) <= not (a or b);
    layer1_outputs(1044) <= not b;
    layer1_outputs(1045) <= a and b;
    layer1_outputs(1046) <= b;
    layer1_outputs(1047) <= b and not a;
    layer1_outputs(1048) <= a or b;
    layer1_outputs(1049) <= not a or b;
    layer1_outputs(1050) <= b;
    layer1_outputs(1051) <= a;
    layer1_outputs(1052) <= 1'b1;
    layer1_outputs(1053) <= 1'b1;
    layer1_outputs(1054) <= 1'b1;
    layer1_outputs(1055) <= not (a and b);
    layer1_outputs(1056) <= a;
    layer1_outputs(1057) <= not (a or b);
    layer1_outputs(1058) <= a or b;
    layer1_outputs(1059) <= a xor b;
    layer1_outputs(1060) <= a and not b;
    layer1_outputs(1061) <= not b;
    layer1_outputs(1062) <= not (a or b);
    layer1_outputs(1063) <= b and not a;
    layer1_outputs(1064) <= 1'b1;
    layer1_outputs(1065) <= a;
    layer1_outputs(1066) <= 1'b1;
    layer1_outputs(1067) <= not b or a;
    layer1_outputs(1068) <= a or b;
    layer1_outputs(1069) <= not (a or b);
    layer1_outputs(1070) <= not a or b;
    layer1_outputs(1071) <= 1'b0;
    layer1_outputs(1072) <= 1'b1;
    layer1_outputs(1073) <= not (a or b);
    layer1_outputs(1074) <= not (a or b);
    layer1_outputs(1075) <= a;
    layer1_outputs(1076) <= not a;
    layer1_outputs(1077) <= a;
    layer1_outputs(1078) <= not b;
    layer1_outputs(1079) <= not (a or b);
    layer1_outputs(1080) <= a and not b;
    layer1_outputs(1081) <= not a or b;
    layer1_outputs(1082) <= not a or b;
    layer1_outputs(1083) <= a;
    layer1_outputs(1084) <= 1'b0;
    layer1_outputs(1085) <= not (a and b);
    layer1_outputs(1086) <= a and not b;
    layer1_outputs(1087) <= not b;
    layer1_outputs(1088) <= 1'b0;
    layer1_outputs(1089) <= a and not b;
    layer1_outputs(1090) <= 1'b0;
    layer1_outputs(1091) <= 1'b0;
    layer1_outputs(1092) <= a or b;
    layer1_outputs(1093) <= b;
    layer1_outputs(1094) <= 1'b0;
    layer1_outputs(1095) <= a;
    layer1_outputs(1096) <= 1'b1;
    layer1_outputs(1097) <= a xor b;
    layer1_outputs(1098) <= not a;
    layer1_outputs(1099) <= b;
    layer1_outputs(1100) <= a and not b;
    layer1_outputs(1101) <= not a or b;
    layer1_outputs(1102) <= not a or b;
    layer1_outputs(1103) <= not (a xor b);
    layer1_outputs(1104) <= 1'b0;
    layer1_outputs(1105) <= not a;
    layer1_outputs(1106) <= a and b;
    layer1_outputs(1107) <= a;
    layer1_outputs(1108) <= 1'b1;
    layer1_outputs(1109) <= not a;
    layer1_outputs(1110) <= not b or a;
    layer1_outputs(1111) <= not (a or b);
    layer1_outputs(1112) <= not a or b;
    layer1_outputs(1113) <= a;
    layer1_outputs(1114) <= not (a or b);
    layer1_outputs(1115) <= not a;
    layer1_outputs(1116) <= a and not b;
    layer1_outputs(1117) <= 1'b0;
    layer1_outputs(1118) <= a or b;
    layer1_outputs(1119) <= a xor b;
    layer1_outputs(1120) <= b and not a;
    layer1_outputs(1121) <= not b or a;
    layer1_outputs(1122) <= not b;
    layer1_outputs(1123) <= 1'b0;
    layer1_outputs(1124) <= not b or a;
    layer1_outputs(1125) <= 1'b1;
    layer1_outputs(1126) <= 1'b1;
    layer1_outputs(1127) <= not (a or b);
    layer1_outputs(1128) <= 1'b0;
    layer1_outputs(1129) <= 1'b0;
    layer1_outputs(1130) <= a and b;
    layer1_outputs(1131) <= 1'b1;
    layer1_outputs(1132) <= a and b;
    layer1_outputs(1133) <= not (a xor b);
    layer1_outputs(1134) <= 1'b1;
    layer1_outputs(1135) <= not a or b;
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= not (a or b);
    layer1_outputs(1138) <= a;
    layer1_outputs(1139) <= not b or a;
    layer1_outputs(1140) <= 1'b0;
    layer1_outputs(1141) <= 1'b0;
    layer1_outputs(1142) <= not a or b;
    layer1_outputs(1143) <= a xor b;
    layer1_outputs(1144) <= 1'b1;
    layer1_outputs(1145) <= a and b;
    layer1_outputs(1146) <= 1'b1;
    layer1_outputs(1147) <= a;
    layer1_outputs(1148) <= not a;
    layer1_outputs(1149) <= a or b;
    layer1_outputs(1150) <= a or b;
    layer1_outputs(1151) <= b;
    layer1_outputs(1152) <= b and not a;
    layer1_outputs(1153) <= 1'b0;
    layer1_outputs(1154) <= b;
    layer1_outputs(1155) <= a and b;
    layer1_outputs(1156) <= b;
    layer1_outputs(1157) <= a or b;
    layer1_outputs(1158) <= not a;
    layer1_outputs(1159) <= a or b;
    layer1_outputs(1160) <= b and not a;
    layer1_outputs(1161) <= b;
    layer1_outputs(1162) <= 1'b1;
    layer1_outputs(1163) <= b;
    layer1_outputs(1164) <= b and not a;
    layer1_outputs(1165) <= 1'b1;
    layer1_outputs(1166) <= not a;
    layer1_outputs(1167) <= a or b;
    layer1_outputs(1168) <= b and not a;
    layer1_outputs(1169) <= a and b;
    layer1_outputs(1170) <= a and b;
    layer1_outputs(1171) <= not a or b;
    layer1_outputs(1172) <= not (a and b);
    layer1_outputs(1173) <= not a or b;
    layer1_outputs(1174) <= not (a and b);
    layer1_outputs(1175) <= not (a or b);
    layer1_outputs(1176) <= not b or a;
    layer1_outputs(1177) <= 1'b1;
    layer1_outputs(1178) <= 1'b1;
    layer1_outputs(1179) <= a;
    layer1_outputs(1180) <= a xor b;
    layer1_outputs(1181) <= b;
    layer1_outputs(1182) <= b;
    layer1_outputs(1183) <= not a;
    layer1_outputs(1184) <= not a or b;
    layer1_outputs(1185) <= a xor b;
    layer1_outputs(1186) <= 1'b1;
    layer1_outputs(1187) <= a;
    layer1_outputs(1188) <= 1'b0;
    layer1_outputs(1189) <= not a or b;
    layer1_outputs(1190) <= 1'b1;
    layer1_outputs(1191) <= not (a and b);
    layer1_outputs(1192) <= a or b;
    layer1_outputs(1193) <= b;
    layer1_outputs(1194) <= not (a and b);
    layer1_outputs(1195) <= a;
    layer1_outputs(1196) <= not (a and b);
    layer1_outputs(1197) <= a and b;
    layer1_outputs(1198) <= not b or a;
    layer1_outputs(1199) <= 1'b1;
    layer1_outputs(1200) <= not (a or b);
    layer1_outputs(1201) <= a;
    layer1_outputs(1202) <= a xor b;
    layer1_outputs(1203) <= 1'b1;
    layer1_outputs(1204) <= a xor b;
    layer1_outputs(1205) <= b and not a;
    layer1_outputs(1206) <= a and b;
    layer1_outputs(1207) <= not (a and b);
    layer1_outputs(1208) <= not a;
    layer1_outputs(1209) <= not b or a;
    layer1_outputs(1210) <= b;
    layer1_outputs(1211) <= b and not a;
    layer1_outputs(1212) <= 1'b0;
    layer1_outputs(1213) <= a or b;
    layer1_outputs(1214) <= not a;
    layer1_outputs(1215) <= 1'b0;
    layer1_outputs(1216) <= 1'b0;
    layer1_outputs(1217) <= not (a or b);
    layer1_outputs(1218) <= a and b;
    layer1_outputs(1219) <= not b;
    layer1_outputs(1220) <= a;
    layer1_outputs(1221) <= a xor b;
    layer1_outputs(1222) <= not a;
    layer1_outputs(1223) <= 1'b1;
    layer1_outputs(1224) <= 1'b1;
    layer1_outputs(1225) <= not b;
    layer1_outputs(1226) <= a and b;
    layer1_outputs(1227) <= 1'b1;
    layer1_outputs(1228) <= not a;
    layer1_outputs(1229) <= not b;
    layer1_outputs(1230) <= b and not a;
    layer1_outputs(1231) <= not b;
    layer1_outputs(1232) <= not (a and b);
    layer1_outputs(1233) <= not (a or b);
    layer1_outputs(1234) <= a and not b;
    layer1_outputs(1235) <= b and not a;
    layer1_outputs(1236) <= b;
    layer1_outputs(1237) <= not b;
    layer1_outputs(1238) <= not (a or b);
    layer1_outputs(1239) <= not b;
    layer1_outputs(1240) <= not a;
    layer1_outputs(1241) <= not (a and b);
    layer1_outputs(1242) <= a or b;
    layer1_outputs(1243) <= not (a and b);
    layer1_outputs(1244) <= a and not b;
    layer1_outputs(1245) <= 1'b0;
    layer1_outputs(1246) <= a and b;
    layer1_outputs(1247) <= not a or b;
    layer1_outputs(1248) <= b and not a;
    layer1_outputs(1249) <= not b;
    layer1_outputs(1250) <= not b or a;
    layer1_outputs(1251) <= 1'b1;
    layer1_outputs(1252) <= 1'b1;
    layer1_outputs(1253) <= not a or b;
    layer1_outputs(1254) <= b and not a;
    layer1_outputs(1255) <= a;
    layer1_outputs(1256) <= not b;
    layer1_outputs(1257) <= a and b;
    layer1_outputs(1258) <= not (a and b);
    layer1_outputs(1259) <= a and not b;
    layer1_outputs(1260) <= 1'b0;
    layer1_outputs(1261) <= not (a or b);
    layer1_outputs(1262) <= a and b;
    layer1_outputs(1263) <= a;
    layer1_outputs(1264) <= 1'b0;
    layer1_outputs(1265) <= not b or a;
    layer1_outputs(1266) <= 1'b1;
    layer1_outputs(1267) <= 1'b1;
    layer1_outputs(1268) <= b and not a;
    layer1_outputs(1269) <= b and not a;
    layer1_outputs(1270) <= not (a xor b);
    layer1_outputs(1271) <= not a;
    layer1_outputs(1272) <= 1'b0;
    layer1_outputs(1273) <= 1'b0;
    layer1_outputs(1274) <= 1'b0;
    layer1_outputs(1275) <= a and b;
    layer1_outputs(1276) <= a or b;
    layer1_outputs(1277) <= a and b;
    layer1_outputs(1278) <= not b;
    layer1_outputs(1279) <= a;
    layer1_outputs(1280) <= a and b;
    layer1_outputs(1281) <= a and not b;
    layer1_outputs(1282) <= a and b;
    layer1_outputs(1283) <= 1'b0;
    layer1_outputs(1284) <= not (a and b);
    layer1_outputs(1285) <= a;
    layer1_outputs(1286) <= not a;
    layer1_outputs(1287) <= not (a or b);
    layer1_outputs(1288) <= 1'b1;
    layer1_outputs(1289) <= not a;
    layer1_outputs(1290) <= 1'b0;
    layer1_outputs(1291) <= not a;
    layer1_outputs(1292) <= not (a or b);
    layer1_outputs(1293) <= a;
    layer1_outputs(1294) <= a or b;
    layer1_outputs(1295) <= 1'b1;
    layer1_outputs(1296) <= 1'b0;
    layer1_outputs(1297) <= 1'b1;
    layer1_outputs(1298) <= 1'b0;
    layer1_outputs(1299) <= not a or b;
    layer1_outputs(1300) <= a or b;
    layer1_outputs(1301) <= not (a and b);
    layer1_outputs(1302) <= a and not b;
    layer1_outputs(1303) <= a and b;
    layer1_outputs(1304) <= 1'b0;
    layer1_outputs(1305) <= a;
    layer1_outputs(1306) <= not b or a;
    layer1_outputs(1307) <= not (a xor b);
    layer1_outputs(1308) <= not (a or b);
    layer1_outputs(1309) <= not (a or b);
    layer1_outputs(1310) <= b and not a;
    layer1_outputs(1311) <= b and not a;
    layer1_outputs(1312) <= a;
    layer1_outputs(1313) <= not (a or b);
    layer1_outputs(1314) <= a;
    layer1_outputs(1315) <= not b;
    layer1_outputs(1316) <= a;
    layer1_outputs(1317) <= 1'b1;
    layer1_outputs(1318) <= b;
    layer1_outputs(1319) <= not b or a;
    layer1_outputs(1320) <= 1'b0;
    layer1_outputs(1321) <= not a;
    layer1_outputs(1322) <= 1'b1;
    layer1_outputs(1323) <= a and b;
    layer1_outputs(1324) <= a;
    layer1_outputs(1325) <= a;
    layer1_outputs(1326) <= not b;
    layer1_outputs(1327) <= not (a or b);
    layer1_outputs(1328) <= not a;
    layer1_outputs(1329) <= b and not a;
    layer1_outputs(1330) <= not a or b;
    layer1_outputs(1331) <= 1'b1;
    layer1_outputs(1332) <= b;
    layer1_outputs(1333) <= not b;
    layer1_outputs(1334) <= 1'b1;
    layer1_outputs(1335) <= b;
    layer1_outputs(1336) <= not b;
    layer1_outputs(1337) <= 1'b1;
    layer1_outputs(1338) <= a xor b;
    layer1_outputs(1339) <= a or b;
    layer1_outputs(1340) <= not (a and b);
    layer1_outputs(1341) <= a xor b;
    layer1_outputs(1342) <= b and not a;
    layer1_outputs(1343) <= 1'b1;
    layer1_outputs(1344) <= not (a and b);
    layer1_outputs(1345) <= not (a and b);
    layer1_outputs(1346) <= a and not b;
    layer1_outputs(1347) <= a and b;
    layer1_outputs(1348) <= 1'b1;
    layer1_outputs(1349) <= a and not b;
    layer1_outputs(1350) <= 1'b1;
    layer1_outputs(1351) <= not (a and b);
    layer1_outputs(1352) <= 1'b1;
    layer1_outputs(1353) <= 1'b0;
    layer1_outputs(1354) <= 1'b0;
    layer1_outputs(1355) <= a;
    layer1_outputs(1356) <= a and not b;
    layer1_outputs(1357) <= a or b;
    layer1_outputs(1358) <= a and not b;
    layer1_outputs(1359) <= not b;
    layer1_outputs(1360) <= not b;
    layer1_outputs(1361) <= a and b;
    layer1_outputs(1362) <= a or b;
    layer1_outputs(1363) <= a and not b;
    layer1_outputs(1364) <= not (a and b);
    layer1_outputs(1365) <= not (a xor b);
    layer1_outputs(1366) <= b and not a;
    layer1_outputs(1367) <= 1'b0;
    layer1_outputs(1368) <= a and b;
    layer1_outputs(1369) <= not a;
    layer1_outputs(1370) <= not a or b;
    layer1_outputs(1371) <= 1'b1;
    layer1_outputs(1372) <= b and not a;
    layer1_outputs(1373) <= not b;
    layer1_outputs(1374) <= not (a and b);
    layer1_outputs(1375) <= not (a or b);
    layer1_outputs(1376) <= not b or a;
    layer1_outputs(1377) <= a and not b;
    layer1_outputs(1378) <= not b or a;
    layer1_outputs(1379) <= not a;
    layer1_outputs(1380) <= not a or b;
    layer1_outputs(1381) <= not b or a;
    layer1_outputs(1382) <= 1'b0;
    layer1_outputs(1383) <= not b or a;
    layer1_outputs(1384) <= a and b;
    layer1_outputs(1385) <= a;
    layer1_outputs(1386) <= not a or b;
    layer1_outputs(1387) <= a or b;
    layer1_outputs(1388) <= a and b;
    layer1_outputs(1389) <= not (a and b);
    layer1_outputs(1390) <= a and b;
    layer1_outputs(1391) <= not b;
    layer1_outputs(1392) <= not b;
    layer1_outputs(1393) <= not a;
    layer1_outputs(1394) <= a and b;
    layer1_outputs(1395) <= not a or b;
    layer1_outputs(1396) <= b and not a;
    layer1_outputs(1397) <= not (a and b);
    layer1_outputs(1398) <= not a or b;
    layer1_outputs(1399) <= a and b;
    layer1_outputs(1400) <= a or b;
    layer1_outputs(1401) <= not b;
    layer1_outputs(1402) <= not (a and b);
    layer1_outputs(1403) <= not (a and b);
    layer1_outputs(1404) <= not (a and b);
    layer1_outputs(1405) <= a xor b;
    layer1_outputs(1406) <= not a;
    layer1_outputs(1407) <= b and not a;
    layer1_outputs(1408) <= not b or a;
    layer1_outputs(1409) <= a and b;
    layer1_outputs(1410) <= b;
    layer1_outputs(1411) <= b and not a;
    layer1_outputs(1412) <= not a;
    layer1_outputs(1413) <= a or b;
    layer1_outputs(1414) <= b and not a;
    layer1_outputs(1415) <= a and not b;
    layer1_outputs(1416) <= not b;
    layer1_outputs(1417) <= 1'b1;
    layer1_outputs(1418) <= not b;
    layer1_outputs(1419) <= b;
    layer1_outputs(1420) <= not b or a;
    layer1_outputs(1421) <= not b or a;
    layer1_outputs(1422) <= a and b;
    layer1_outputs(1423) <= 1'b0;
    layer1_outputs(1424) <= not b;
    layer1_outputs(1425) <= 1'b1;
    layer1_outputs(1426) <= not b or a;
    layer1_outputs(1427) <= b and not a;
    layer1_outputs(1428) <= not (a or b);
    layer1_outputs(1429) <= not a;
    layer1_outputs(1430) <= b;
    layer1_outputs(1431) <= a and b;
    layer1_outputs(1432) <= not (a and b);
    layer1_outputs(1433) <= 1'b1;
    layer1_outputs(1434) <= a and not b;
    layer1_outputs(1435) <= a;
    layer1_outputs(1436) <= a or b;
    layer1_outputs(1437) <= not a or b;
    layer1_outputs(1438) <= not b or a;
    layer1_outputs(1439) <= not (a and b);
    layer1_outputs(1440) <= not b;
    layer1_outputs(1441) <= b and not a;
    layer1_outputs(1442) <= a;
    layer1_outputs(1443) <= 1'b1;
    layer1_outputs(1444) <= a or b;
    layer1_outputs(1445) <= 1'b0;
    layer1_outputs(1446) <= not (a xor b);
    layer1_outputs(1447) <= a and b;
    layer1_outputs(1448) <= b;
    layer1_outputs(1449) <= b and not a;
    layer1_outputs(1450) <= 1'b1;
    layer1_outputs(1451) <= not b;
    layer1_outputs(1452) <= not b;
    layer1_outputs(1453) <= a xor b;
    layer1_outputs(1454) <= not b or a;
    layer1_outputs(1455) <= a and not b;
    layer1_outputs(1456) <= b and not a;
    layer1_outputs(1457) <= a;
    layer1_outputs(1458) <= 1'b1;
    layer1_outputs(1459) <= b;
    layer1_outputs(1460) <= a and b;
    layer1_outputs(1461) <= b;
    layer1_outputs(1462) <= not (a or b);
    layer1_outputs(1463) <= 1'b0;
    layer1_outputs(1464) <= not b;
    layer1_outputs(1465) <= not b;
    layer1_outputs(1466) <= not b or a;
    layer1_outputs(1467) <= not (a and b);
    layer1_outputs(1468) <= not (a and b);
    layer1_outputs(1469) <= 1'b1;
    layer1_outputs(1470) <= b and not a;
    layer1_outputs(1471) <= 1'b1;
    layer1_outputs(1472) <= not (a or b);
    layer1_outputs(1473) <= not a;
    layer1_outputs(1474) <= a and not b;
    layer1_outputs(1475) <= not a;
    layer1_outputs(1476) <= not (a and b);
    layer1_outputs(1477) <= not b or a;
    layer1_outputs(1478) <= not (a and b);
    layer1_outputs(1479) <= 1'b1;
    layer1_outputs(1480) <= 1'b0;
    layer1_outputs(1481) <= a and b;
    layer1_outputs(1482) <= a or b;
    layer1_outputs(1483) <= not a or b;
    layer1_outputs(1484) <= a and b;
    layer1_outputs(1485) <= not b;
    layer1_outputs(1486) <= 1'b1;
    layer1_outputs(1487) <= not (a xor b);
    layer1_outputs(1488) <= a and not b;
    layer1_outputs(1489) <= not (a or b);
    layer1_outputs(1490) <= not a;
    layer1_outputs(1491) <= not b or a;
    layer1_outputs(1492) <= not (a and b);
    layer1_outputs(1493) <= not (a and b);
    layer1_outputs(1494) <= not (a or b);
    layer1_outputs(1495) <= a and b;
    layer1_outputs(1496) <= 1'b1;
    layer1_outputs(1497) <= not (a xor b);
    layer1_outputs(1498) <= not (a or b);
    layer1_outputs(1499) <= not b;
    layer1_outputs(1500) <= not b or a;
    layer1_outputs(1501) <= 1'b1;
    layer1_outputs(1502) <= not (a or b);
    layer1_outputs(1503) <= b and not a;
    layer1_outputs(1504) <= not (a or b);
    layer1_outputs(1505) <= b;
    layer1_outputs(1506) <= b;
    layer1_outputs(1507) <= a and b;
    layer1_outputs(1508) <= 1'b1;
    layer1_outputs(1509) <= not b;
    layer1_outputs(1510) <= not a;
    layer1_outputs(1511) <= a and b;
    layer1_outputs(1512) <= a;
    layer1_outputs(1513) <= not a or b;
    layer1_outputs(1514) <= 1'b1;
    layer1_outputs(1515) <= not (a and b);
    layer1_outputs(1516) <= not a;
    layer1_outputs(1517) <= not a;
    layer1_outputs(1518) <= a or b;
    layer1_outputs(1519) <= not (a xor b);
    layer1_outputs(1520) <= b;
    layer1_outputs(1521) <= not a or b;
    layer1_outputs(1522) <= not a;
    layer1_outputs(1523) <= not (a xor b);
    layer1_outputs(1524) <= a and b;
    layer1_outputs(1525) <= not a or b;
    layer1_outputs(1526) <= 1'b0;
    layer1_outputs(1527) <= a and not b;
    layer1_outputs(1528) <= not a or b;
    layer1_outputs(1529) <= not (a xor b);
    layer1_outputs(1530) <= 1'b1;
    layer1_outputs(1531) <= not (a and b);
    layer1_outputs(1532) <= 1'b0;
    layer1_outputs(1533) <= 1'b1;
    layer1_outputs(1534) <= not (a and b);
    layer1_outputs(1535) <= 1'b1;
    layer1_outputs(1536) <= a;
    layer1_outputs(1537) <= 1'b0;
    layer1_outputs(1538) <= not (a or b);
    layer1_outputs(1539) <= b;
    layer1_outputs(1540) <= a or b;
    layer1_outputs(1541) <= not (a or b);
    layer1_outputs(1542) <= not (a and b);
    layer1_outputs(1543) <= 1'b1;
    layer1_outputs(1544) <= not (a and b);
    layer1_outputs(1545) <= a and b;
    layer1_outputs(1546) <= not b or a;
    layer1_outputs(1547) <= not a or b;
    layer1_outputs(1548) <= not a or b;
    layer1_outputs(1549) <= not a or b;
    layer1_outputs(1550) <= not (a xor b);
    layer1_outputs(1551) <= 1'b1;
    layer1_outputs(1552) <= a;
    layer1_outputs(1553) <= not a or b;
    layer1_outputs(1554) <= a and b;
    layer1_outputs(1555) <= not a;
    layer1_outputs(1556) <= a or b;
    layer1_outputs(1557) <= a and b;
    layer1_outputs(1558) <= not (a or b);
    layer1_outputs(1559) <= b and not a;
    layer1_outputs(1560) <= 1'b0;
    layer1_outputs(1561) <= not a or b;
    layer1_outputs(1562) <= 1'b1;
    layer1_outputs(1563) <= a or b;
    layer1_outputs(1564) <= 1'b1;
    layer1_outputs(1565) <= not a or b;
    layer1_outputs(1566) <= not (a or b);
    layer1_outputs(1567) <= 1'b1;
    layer1_outputs(1568) <= not (a or b);
    layer1_outputs(1569) <= 1'b0;
    layer1_outputs(1570) <= not (a or b);
    layer1_outputs(1571) <= not b or a;
    layer1_outputs(1572) <= not b or a;
    layer1_outputs(1573) <= 1'b1;
    layer1_outputs(1574) <= not a;
    layer1_outputs(1575) <= not b or a;
    layer1_outputs(1576) <= a and not b;
    layer1_outputs(1577) <= 1'b0;
    layer1_outputs(1578) <= not a or b;
    layer1_outputs(1579) <= b;
    layer1_outputs(1580) <= a xor b;
    layer1_outputs(1581) <= not (a or b);
    layer1_outputs(1582) <= not (a and b);
    layer1_outputs(1583) <= not b;
    layer1_outputs(1584) <= not (a or b);
    layer1_outputs(1585) <= 1'b0;
    layer1_outputs(1586) <= b and not a;
    layer1_outputs(1587) <= a;
    layer1_outputs(1588) <= 1'b1;
    layer1_outputs(1589) <= not b;
    layer1_outputs(1590) <= not (a xor b);
    layer1_outputs(1591) <= 1'b0;
    layer1_outputs(1592) <= not (a and b);
    layer1_outputs(1593) <= not (a or b);
    layer1_outputs(1594) <= 1'b1;
    layer1_outputs(1595) <= a;
    layer1_outputs(1596) <= a or b;
    layer1_outputs(1597) <= not (a or b);
    layer1_outputs(1598) <= a;
    layer1_outputs(1599) <= not a or b;
    layer1_outputs(1600) <= a xor b;
    layer1_outputs(1601) <= not (a or b);
    layer1_outputs(1602) <= a and not b;
    layer1_outputs(1603) <= a or b;
    layer1_outputs(1604) <= not (a and b);
    layer1_outputs(1605) <= 1'b1;
    layer1_outputs(1606) <= a or b;
    layer1_outputs(1607) <= 1'b1;
    layer1_outputs(1608) <= 1'b1;
    layer1_outputs(1609) <= 1'b0;
    layer1_outputs(1610) <= b and not a;
    layer1_outputs(1611) <= not (a xor b);
    layer1_outputs(1612) <= not a;
    layer1_outputs(1613) <= not a;
    layer1_outputs(1614) <= a;
    layer1_outputs(1615) <= a or b;
    layer1_outputs(1616) <= not a;
    layer1_outputs(1617) <= not b or a;
    layer1_outputs(1618) <= 1'b1;
    layer1_outputs(1619) <= not (a or b);
    layer1_outputs(1620) <= a;
    layer1_outputs(1621) <= not (a and b);
    layer1_outputs(1622) <= not b or a;
    layer1_outputs(1623) <= not (a and b);
    layer1_outputs(1624) <= 1'b0;
    layer1_outputs(1625) <= 1'b0;
    layer1_outputs(1626) <= not (a and b);
    layer1_outputs(1627) <= not a;
    layer1_outputs(1628) <= a and not b;
    layer1_outputs(1629) <= not b or a;
    layer1_outputs(1630) <= not (a and b);
    layer1_outputs(1631) <= not b or a;
    layer1_outputs(1632) <= a and not b;
    layer1_outputs(1633) <= not b or a;
    layer1_outputs(1634) <= 1'b1;
    layer1_outputs(1635) <= 1'b1;
    layer1_outputs(1636) <= 1'b0;
    layer1_outputs(1637) <= a or b;
    layer1_outputs(1638) <= a or b;
    layer1_outputs(1639) <= not (a or b);
    layer1_outputs(1640) <= 1'b1;
    layer1_outputs(1641) <= b;
    layer1_outputs(1642) <= not a;
    layer1_outputs(1643) <= b;
    layer1_outputs(1644) <= 1'b0;
    layer1_outputs(1645) <= not (a and b);
    layer1_outputs(1646) <= a or b;
    layer1_outputs(1647) <= 1'b0;
    layer1_outputs(1648) <= not a or b;
    layer1_outputs(1649) <= a and b;
    layer1_outputs(1650) <= not (a or b);
    layer1_outputs(1651) <= not (a or b);
    layer1_outputs(1652) <= not b;
    layer1_outputs(1653) <= 1'b0;
    layer1_outputs(1654) <= 1'b1;
    layer1_outputs(1655) <= 1'b1;
    layer1_outputs(1656) <= a xor b;
    layer1_outputs(1657) <= a;
    layer1_outputs(1658) <= not b or a;
    layer1_outputs(1659) <= a and b;
    layer1_outputs(1660) <= not a;
    layer1_outputs(1661) <= a or b;
    layer1_outputs(1662) <= not a;
    layer1_outputs(1663) <= not (a or b);
    layer1_outputs(1664) <= a or b;
    layer1_outputs(1665) <= a;
    layer1_outputs(1666) <= a or b;
    layer1_outputs(1667) <= a and b;
    layer1_outputs(1668) <= a and b;
    layer1_outputs(1669) <= b;
    layer1_outputs(1670) <= not (a and b);
    layer1_outputs(1671) <= b;
    layer1_outputs(1672) <= b and not a;
    layer1_outputs(1673) <= b and not a;
    layer1_outputs(1674) <= not a;
    layer1_outputs(1675) <= 1'b0;
    layer1_outputs(1676) <= not (a and b);
    layer1_outputs(1677) <= not a or b;
    layer1_outputs(1678) <= 1'b0;
    layer1_outputs(1679) <= a and b;
    layer1_outputs(1680) <= a or b;
    layer1_outputs(1681) <= not b;
    layer1_outputs(1682) <= a and not b;
    layer1_outputs(1683) <= not b;
    layer1_outputs(1684) <= 1'b1;
    layer1_outputs(1685) <= a;
    layer1_outputs(1686) <= a xor b;
    layer1_outputs(1687) <= 1'b1;
    layer1_outputs(1688) <= a and not b;
    layer1_outputs(1689) <= not a;
    layer1_outputs(1690) <= b and not a;
    layer1_outputs(1691) <= 1'b1;
    layer1_outputs(1692) <= not a or b;
    layer1_outputs(1693) <= 1'b1;
    layer1_outputs(1694) <= 1'b1;
    layer1_outputs(1695) <= 1'b0;
    layer1_outputs(1696) <= 1'b1;
    layer1_outputs(1697) <= not (a or b);
    layer1_outputs(1698) <= not (a and b);
    layer1_outputs(1699) <= a and b;
    layer1_outputs(1700) <= a and not b;
    layer1_outputs(1701) <= 1'b1;
    layer1_outputs(1702) <= a and b;
    layer1_outputs(1703) <= a and not b;
    layer1_outputs(1704) <= a or b;
    layer1_outputs(1705) <= 1'b1;
    layer1_outputs(1706) <= not b or a;
    layer1_outputs(1707) <= a and not b;
    layer1_outputs(1708) <= not a or b;
    layer1_outputs(1709) <= not a or b;
    layer1_outputs(1710) <= b;
    layer1_outputs(1711) <= a and not b;
    layer1_outputs(1712) <= not (a xor b);
    layer1_outputs(1713) <= not a;
    layer1_outputs(1714) <= not (a and b);
    layer1_outputs(1715) <= not (a or b);
    layer1_outputs(1716) <= 1'b0;
    layer1_outputs(1717) <= not a or b;
    layer1_outputs(1718) <= not b;
    layer1_outputs(1719) <= a and not b;
    layer1_outputs(1720) <= a and not b;
    layer1_outputs(1721) <= a and b;
    layer1_outputs(1722) <= not b or a;
    layer1_outputs(1723) <= a and not b;
    layer1_outputs(1724) <= a and b;
    layer1_outputs(1725) <= a and not b;
    layer1_outputs(1726) <= a;
    layer1_outputs(1727) <= not (a or b);
    layer1_outputs(1728) <= a or b;
    layer1_outputs(1729) <= not b;
    layer1_outputs(1730) <= a;
    layer1_outputs(1731) <= a;
    layer1_outputs(1732) <= not (a or b);
    layer1_outputs(1733) <= 1'b0;
    layer1_outputs(1734) <= 1'b0;
    layer1_outputs(1735) <= a and not b;
    layer1_outputs(1736) <= a and b;
    layer1_outputs(1737) <= 1'b0;
    layer1_outputs(1738) <= b;
    layer1_outputs(1739) <= not b or a;
    layer1_outputs(1740) <= not b or a;
    layer1_outputs(1741) <= a and not b;
    layer1_outputs(1742) <= a;
    layer1_outputs(1743) <= 1'b1;
    layer1_outputs(1744) <= not b;
    layer1_outputs(1745) <= 1'b1;
    layer1_outputs(1746) <= 1'b0;
    layer1_outputs(1747) <= a or b;
    layer1_outputs(1748) <= not b or a;
    layer1_outputs(1749) <= not a;
    layer1_outputs(1750) <= b and not a;
    layer1_outputs(1751) <= not a;
    layer1_outputs(1752) <= a and b;
    layer1_outputs(1753) <= not (a and b);
    layer1_outputs(1754) <= a and b;
    layer1_outputs(1755) <= not (a or b);
    layer1_outputs(1756) <= 1'b0;
    layer1_outputs(1757) <= not a;
    layer1_outputs(1758) <= 1'b1;
    layer1_outputs(1759) <= b and not a;
    layer1_outputs(1760) <= 1'b1;
    layer1_outputs(1761) <= not (a and b);
    layer1_outputs(1762) <= not (a or b);
    layer1_outputs(1763) <= not (a or b);
    layer1_outputs(1764) <= a and not b;
    layer1_outputs(1765) <= a and not b;
    layer1_outputs(1766) <= a;
    layer1_outputs(1767) <= not a;
    layer1_outputs(1768) <= not a or b;
    layer1_outputs(1769) <= not b;
    layer1_outputs(1770) <= not (a or b);
    layer1_outputs(1771) <= not a;
    layer1_outputs(1772) <= not a or b;
    layer1_outputs(1773) <= a and b;
    layer1_outputs(1774) <= 1'b1;
    layer1_outputs(1775) <= a;
    layer1_outputs(1776) <= 1'b1;
    layer1_outputs(1777) <= a and not b;
    layer1_outputs(1778) <= not (a or b);
    layer1_outputs(1779) <= b;
    layer1_outputs(1780) <= 1'b0;
    layer1_outputs(1781) <= a and b;
    layer1_outputs(1782) <= 1'b0;
    layer1_outputs(1783) <= a and not b;
    layer1_outputs(1784) <= not b or a;
    layer1_outputs(1785) <= not (a and b);
    layer1_outputs(1786) <= b;
    layer1_outputs(1787) <= b and not a;
    layer1_outputs(1788) <= b and not a;
    layer1_outputs(1789) <= not a or b;
    layer1_outputs(1790) <= not b or a;
    layer1_outputs(1791) <= not a or b;
    layer1_outputs(1792) <= a and not b;
    layer1_outputs(1793) <= 1'b0;
    layer1_outputs(1794) <= not b;
    layer1_outputs(1795) <= 1'b1;
    layer1_outputs(1796) <= 1'b1;
    layer1_outputs(1797) <= a;
    layer1_outputs(1798) <= a and not b;
    layer1_outputs(1799) <= not a or b;
    layer1_outputs(1800) <= 1'b1;
    layer1_outputs(1801) <= b;
    layer1_outputs(1802) <= 1'b1;
    layer1_outputs(1803) <= 1'b1;
    layer1_outputs(1804) <= 1'b1;
    layer1_outputs(1805) <= b and not a;
    layer1_outputs(1806) <= not b or a;
    layer1_outputs(1807) <= a;
    layer1_outputs(1808) <= not (a or b);
    layer1_outputs(1809) <= not a;
    layer1_outputs(1810) <= not (a or b);
    layer1_outputs(1811) <= a and not b;
    layer1_outputs(1812) <= not b;
    layer1_outputs(1813) <= not (a or b);
    layer1_outputs(1814) <= not a;
    layer1_outputs(1815) <= a and not b;
    layer1_outputs(1816) <= b and not a;
    layer1_outputs(1817) <= a and b;
    layer1_outputs(1818) <= not b or a;
    layer1_outputs(1819) <= not b or a;
    layer1_outputs(1820) <= 1'b0;
    layer1_outputs(1821) <= not (a or b);
    layer1_outputs(1822) <= 1'b0;
    layer1_outputs(1823) <= a and b;
    layer1_outputs(1824) <= a and b;
    layer1_outputs(1825) <= b;
    layer1_outputs(1826) <= 1'b1;
    layer1_outputs(1827) <= not (a xor b);
    layer1_outputs(1828) <= 1'b1;
    layer1_outputs(1829) <= not b or a;
    layer1_outputs(1830) <= not (a and b);
    layer1_outputs(1831) <= not b or a;
    layer1_outputs(1832) <= not a or b;
    layer1_outputs(1833) <= 1'b1;
    layer1_outputs(1834) <= not (a and b);
    layer1_outputs(1835) <= b and not a;
    layer1_outputs(1836) <= not a or b;
    layer1_outputs(1837) <= a xor b;
    layer1_outputs(1838) <= 1'b0;
    layer1_outputs(1839) <= a;
    layer1_outputs(1840) <= b and not a;
    layer1_outputs(1841) <= a;
    layer1_outputs(1842) <= a and not b;
    layer1_outputs(1843) <= a or b;
    layer1_outputs(1844) <= not (a or b);
    layer1_outputs(1845) <= 1'b1;
    layer1_outputs(1846) <= not a;
    layer1_outputs(1847) <= not b;
    layer1_outputs(1848) <= b;
    layer1_outputs(1849) <= not (a and b);
    layer1_outputs(1850) <= a;
    layer1_outputs(1851) <= not b;
    layer1_outputs(1852) <= not (a or b);
    layer1_outputs(1853) <= not a;
    layer1_outputs(1854) <= b and not a;
    layer1_outputs(1855) <= not (a or b);
    layer1_outputs(1856) <= a and b;
    layer1_outputs(1857) <= a or b;
    layer1_outputs(1858) <= a;
    layer1_outputs(1859) <= b and not a;
    layer1_outputs(1860) <= b and not a;
    layer1_outputs(1861) <= b and not a;
    layer1_outputs(1862) <= a;
    layer1_outputs(1863) <= a and not b;
    layer1_outputs(1864) <= a and b;
    layer1_outputs(1865) <= 1'b0;
    layer1_outputs(1866) <= not a or b;
    layer1_outputs(1867) <= not b or a;
    layer1_outputs(1868) <= 1'b1;
    layer1_outputs(1869) <= not (a xor b);
    layer1_outputs(1870) <= 1'b1;
    layer1_outputs(1871) <= 1'b0;
    layer1_outputs(1872) <= 1'b0;
    layer1_outputs(1873) <= not a or b;
    layer1_outputs(1874) <= a;
    layer1_outputs(1875) <= not a or b;
    layer1_outputs(1876) <= 1'b1;
    layer1_outputs(1877) <= b and not a;
    layer1_outputs(1878) <= a;
    layer1_outputs(1879) <= 1'b0;
    layer1_outputs(1880) <= a and not b;
    layer1_outputs(1881) <= a and not b;
    layer1_outputs(1882) <= 1'b1;
    layer1_outputs(1883) <= 1'b0;
    layer1_outputs(1884) <= b;
    layer1_outputs(1885) <= 1'b1;
    layer1_outputs(1886) <= 1'b0;
    layer1_outputs(1887) <= not b or a;
    layer1_outputs(1888) <= a xor b;
    layer1_outputs(1889) <= a or b;
    layer1_outputs(1890) <= a;
    layer1_outputs(1891) <= 1'b0;
    layer1_outputs(1892) <= not (a and b);
    layer1_outputs(1893) <= not (a and b);
    layer1_outputs(1894) <= not a or b;
    layer1_outputs(1895) <= a;
    layer1_outputs(1896) <= not (a xor b);
    layer1_outputs(1897) <= 1'b0;
    layer1_outputs(1898) <= a;
    layer1_outputs(1899) <= not a or b;
    layer1_outputs(1900) <= not a or b;
    layer1_outputs(1901) <= not (a or b);
    layer1_outputs(1902) <= 1'b1;
    layer1_outputs(1903) <= a and b;
    layer1_outputs(1904) <= not b or a;
    layer1_outputs(1905) <= b and not a;
    layer1_outputs(1906) <= not b or a;
    layer1_outputs(1907) <= not (a xor b);
    layer1_outputs(1908) <= not a or b;
    layer1_outputs(1909) <= a xor b;
    layer1_outputs(1910) <= 1'b1;
    layer1_outputs(1911) <= a and not b;
    layer1_outputs(1912) <= a and b;
    layer1_outputs(1913) <= a and b;
    layer1_outputs(1914) <= a or b;
    layer1_outputs(1915) <= 1'b1;
    layer1_outputs(1916) <= 1'b0;
    layer1_outputs(1917) <= not a;
    layer1_outputs(1918) <= a or b;
    layer1_outputs(1919) <= a;
    layer1_outputs(1920) <= not (a xor b);
    layer1_outputs(1921) <= a;
    layer1_outputs(1922) <= not b or a;
    layer1_outputs(1923) <= a;
    layer1_outputs(1924) <= a and not b;
    layer1_outputs(1925) <= 1'b0;
    layer1_outputs(1926) <= not b or a;
    layer1_outputs(1927) <= a and b;
    layer1_outputs(1928) <= not a;
    layer1_outputs(1929) <= a xor b;
    layer1_outputs(1930) <= not (a or b);
    layer1_outputs(1931) <= b;
    layer1_outputs(1932) <= a;
    layer1_outputs(1933) <= not (a xor b);
    layer1_outputs(1934) <= a and b;
    layer1_outputs(1935) <= a or b;
    layer1_outputs(1936) <= a;
    layer1_outputs(1937) <= not (a and b);
    layer1_outputs(1938) <= b;
    layer1_outputs(1939) <= not (a and b);
    layer1_outputs(1940) <= b and not a;
    layer1_outputs(1941) <= a and b;
    layer1_outputs(1942) <= a and not b;
    layer1_outputs(1943) <= not b or a;
    layer1_outputs(1944) <= a or b;
    layer1_outputs(1945) <= not (a and b);
    layer1_outputs(1946) <= a and b;
    layer1_outputs(1947) <= a or b;
    layer1_outputs(1948) <= 1'b0;
    layer1_outputs(1949) <= 1'b0;
    layer1_outputs(1950) <= b;
    layer1_outputs(1951) <= 1'b1;
    layer1_outputs(1952) <= 1'b1;
    layer1_outputs(1953) <= 1'b1;
    layer1_outputs(1954) <= not (a xor b);
    layer1_outputs(1955) <= not (a or b);
    layer1_outputs(1956) <= not (a and b);
    layer1_outputs(1957) <= not b or a;
    layer1_outputs(1958) <= a;
    layer1_outputs(1959) <= a;
    layer1_outputs(1960) <= a;
    layer1_outputs(1961) <= a or b;
    layer1_outputs(1962) <= 1'b1;
    layer1_outputs(1963) <= b and not a;
    layer1_outputs(1964) <= a;
    layer1_outputs(1965) <= not a or b;
    layer1_outputs(1966) <= not a;
    layer1_outputs(1967) <= 1'b0;
    layer1_outputs(1968) <= not b;
    layer1_outputs(1969) <= 1'b1;
    layer1_outputs(1970) <= 1'b0;
    layer1_outputs(1971) <= not b;
    layer1_outputs(1972) <= a;
    layer1_outputs(1973) <= a or b;
    layer1_outputs(1974) <= not a or b;
    layer1_outputs(1975) <= 1'b0;
    layer1_outputs(1976) <= 1'b0;
    layer1_outputs(1977) <= 1'b1;
    layer1_outputs(1978) <= 1'b1;
    layer1_outputs(1979) <= not a or b;
    layer1_outputs(1980) <= b;
    layer1_outputs(1981) <= a;
    layer1_outputs(1982) <= 1'b1;
    layer1_outputs(1983) <= b and not a;
    layer1_outputs(1984) <= b and not a;
    layer1_outputs(1985) <= a and not b;
    layer1_outputs(1986) <= not a or b;
    layer1_outputs(1987) <= a or b;
    layer1_outputs(1988) <= not b or a;
    layer1_outputs(1989) <= 1'b0;
    layer1_outputs(1990) <= 1'b0;
    layer1_outputs(1991) <= not (a and b);
    layer1_outputs(1992) <= not a;
    layer1_outputs(1993) <= not b or a;
    layer1_outputs(1994) <= not a or b;
    layer1_outputs(1995) <= b;
    layer1_outputs(1996) <= not a or b;
    layer1_outputs(1997) <= not (a or b);
    layer1_outputs(1998) <= a and b;
    layer1_outputs(1999) <= not (a and b);
    layer1_outputs(2000) <= not (a or b);
    layer1_outputs(2001) <= 1'b1;
    layer1_outputs(2002) <= not a or b;
    layer1_outputs(2003) <= 1'b1;
    layer1_outputs(2004) <= not (a xor b);
    layer1_outputs(2005) <= not b or a;
    layer1_outputs(2006) <= a and not b;
    layer1_outputs(2007) <= a;
    layer1_outputs(2008) <= 1'b0;
    layer1_outputs(2009) <= not (a or b);
    layer1_outputs(2010) <= not b or a;
    layer1_outputs(2011) <= not b or a;
    layer1_outputs(2012) <= 1'b1;
    layer1_outputs(2013) <= a and not b;
    layer1_outputs(2014) <= 1'b1;
    layer1_outputs(2015) <= 1'b0;
    layer1_outputs(2016) <= b;
    layer1_outputs(2017) <= b and not a;
    layer1_outputs(2018) <= a;
    layer1_outputs(2019) <= a and b;
    layer1_outputs(2020) <= a;
    layer1_outputs(2021) <= not b;
    layer1_outputs(2022) <= not b or a;
    layer1_outputs(2023) <= 1'b0;
    layer1_outputs(2024) <= not b or a;
    layer1_outputs(2025) <= not (a and b);
    layer1_outputs(2026) <= not a or b;
    layer1_outputs(2027) <= not a or b;
    layer1_outputs(2028) <= not (a xor b);
    layer1_outputs(2029) <= 1'b1;
    layer1_outputs(2030) <= a and b;
    layer1_outputs(2031) <= 1'b0;
    layer1_outputs(2032) <= a or b;
    layer1_outputs(2033) <= a xor b;
    layer1_outputs(2034) <= not b or a;
    layer1_outputs(2035) <= not b;
    layer1_outputs(2036) <= 1'b0;
    layer1_outputs(2037) <= not a;
    layer1_outputs(2038) <= a;
    layer1_outputs(2039) <= not a or b;
    layer1_outputs(2040) <= b and not a;
    layer1_outputs(2041) <= a;
    layer1_outputs(2042) <= a and not b;
    layer1_outputs(2043) <= not a or b;
    layer1_outputs(2044) <= 1'b1;
    layer1_outputs(2045) <= 1'b0;
    layer1_outputs(2046) <= 1'b0;
    layer1_outputs(2047) <= a or b;
    layer1_outputs(2048) <= not (a or b);
    layer1_outputs(2049) <= 1'b0;
    layer1_outputs(2050) <= not (a or b);
    layer1_outputs(2051) <= not b;
    layer1_outputs(2052) <= not (a xor b);
    layer1_outputs(2053) <= 1'b1;
    layer1_outputs(2054) <= not b or a;
    layer1_outputs(2055) <= 1'b1;
    layer1_outputs(2056) <= not (a and b);
    layer1_outputs(2057) <= b and not a;
    layer1_outputs(2058) <= a or b;
    layer1_outputs(2059) <= b;
    layer1_outputs(2060) <= not b;
    layer1_outputs(2061) <= not a or b;
    layer1_outputs(2062) <= 1'b1;
    layer1_outputs(2063) <= not a or b;
    layer1_outputs(2064) <= not a or b;
    layer1_outputs(2065) <= b;
    layer1_outputs(2066) <= not a;
    layer1_outputs(2067) <= b and not a;
    layer1_outputs(2068) <= 1'b0;
    layer1_outputs(2069) <= a or b;
    layer1_outputs(2070) <= not (a and b);
    layer1_outputs(2071) <= b;
    layer1_outputs(2072) <= a and b;
    layer1_outputs(2073) <= a xor b;
    layer1_outputs(2074) <= not b;
    layer1_outputs(2075) <= 1'b0;
    layer1_outputs(2076) <= not a;
    layer1_outputs(2077) <= not (a and b);
    layer1_outputs(2078) <= not (a or b);
    layer1_outputs(2079) <= not (a and b);
    layer1_outputs(2080) <= b;
    layer1_outputs(2081) <= not a or b;
    layer1_outputs(2082) <= 1'b0;
    layer1_outputs(2083) <= 1'b1;
    layer1_outputs(2084) <= not (a or b);
    layer1_outputs(2085) <= b and not a;
    layer1_outputs(2086) <= a or b;
    layer1_outputs(2087) <= not a or b;
    layer1_outputs(2088) <= b and not a;
    layer1_outputs(2089) <= a and not b;
    layer1_outputs(2090) <= a;
    layer1_outputs(2091) <= not (a or b);
    layer1_outputs(2092) <= a and b;
    layer1_outputs(2093) <= a and not b;
    layer1_outputs(2094) <= not a or b;
    layer1_outputs(2095) <= not a;
    layer1_outputs(2096) <= not b or a;
    layer1_outputs(2097) <= 1'b0;
    layer1_outputs(2098) <= a xor b;
    layer1_outputs(2099) <= not (a and b);
    layer1_outputs(2100) <= not b or a;
    layer1_outputs(2101) <= not (a and b);
    layer1_outputs(2102) <= not b or a;
    layer1_outputs(2103) <= b;
    layer1_outputs(2104) <= a;
    layer1_outputs(2105) <= not b;
    layer1_outputs(2106) <= not b or a;
    layer1_outputs(2107) <= not b;
    layer1_outputs(2108) <= 1'b1;
    layer1_outputs(2109) <= not a;
    layer1_outputs(2110) <= a and not b;
    layer1_outputs(2111) <= a and b;
    layer1_outputs(2112) <= 1'b0;
    layer1_outputs(2113) <= a or b;
    layer1_outputs(2114) <= not b;
    layer1_outputs(2115) <= 1'b1;
    layer1_outputs(2116) <= 1'b0;
    layer1_outputs(2117) <= not (a xor b);
    layer1_outputs(2118) <= not a;
    layer1_outputs(2119) <= not b or a;
    layer1_outputs(2120) <= a xor b;
    layer1_outputs(2121) <= not a or b;
    layer1_outputs(2122) <= not (a and b);
    layer1_outputs(2123) <= a and not b;
    layer1_outputs(2124) <= not b;
    layer1_outputs(2125) <= a and not b;
    layer1_outputs(2126) <= 1'b0;
    layer1_outputs(2127) <= not b;
    layer1_outputs(2128) <= not (a and b);
    layer1_outputs(2129) <= 1'b1;
    layer1_outputs(2130) <= not a or b;
    layer1_outputs(2131) <= not b or a;
    layer1_outputs(2132) <= b and not a;
    layer1_outputs(2133) <= b;
    layer1_outputs(2134) <= 1'b0;
    layer1_outputs(2135) <= not b;
    layer1_outputs(2136) <= not a;
    layer1_outputs(2137) <= not a or b;
    layer1_outputs(2138) <= 1'b0;
    layer1_outputs(2139) <= b;
    layer1_outputs(2140) <= not (a and b);
    layer1_outputs(2141) <= 1'b1;
    layer1_outputs(2142) <= not (a or b);
    layer1_outputs(2143) <= a;
    layer1_outputs(2144) <= b;
    layer1_outputs(2145) <= 1'b1;
    layer1_outputs(2146) <= not (a or b);
    layer1_outputs(2147) <= a and not b;
    layer1_outputs(2148) <= a or b;
    layer1_outputs(2149) <= 1'b0;
    layer1_outputs(2150) <= not a;
    layer1_outputs(2151) <= not (a or b);
    layer1_outputs(2152) <= not b or a;
    layer1_outputs(2153) <= 1'b1;
    layer1_outputs(2154) <= 1'b0;
    layer1_outputs(2155) <= not a or b;
    layer1_outputs(2156) <= not (a and b);
    layer1_outputs(2157) <= a and b;
    layer1_outputs(2158) <= not b or a;
    layer1_outputs(2159) <= not (a and b);
    layer1_outputs(2160) <= not (a and b);
    layer1_outputs(2161) <= not (a or b);
    layer1_outputs(2162) <= not (a and b);
    layer1_outputs(2163) <= not a or b;
    layer1_outputs(2164) <= a xor b;
    layer1_outputs(2165) <= not b or a;
    layer1_outputs(2166) <= 1'b0;
    layer1_outputs(2167) <= not b;
    layer1_outputs(2168) <= not b or a;
    layer1_outputs(2169) <= a or b;
    layer1_outputs(2170) <= b and not a;
    layer1_outputs(2171) <= a;
    layer1_outputs(2172) <= b;
    layer1_outputs(2173) <= 1'b1;
    layer1_outputs(2174) <= not (a and b);
    layer1_outputs(2175) <= 1'b1;
    layer1_outputs(2176) <= b;
    layer1_outputs(2177) <= not (a and b);
    layer1_outputs(2178) <= 1'b1;
    layer1_outputs(2179) <= not (a and b);
    layer1_outputs(2180) <= a and b;
    layer1_outputs(2181) <= 1'b1;
    layer1_outputs(2182) <= a;
    layer1_outputs(2183) <= not a;
    layer1_outputs(2184) <= b and not a;
    layer1_outputs(2185) <= not a;
    layer1_outputs(2186) <= b and not a;
    layer1_outputs(2187) <= a or b;
    layer1_outputs(2188) <= a and b;
    layer1_outputs(2189) <= not (a or b);
    layer1_outputs(2190) <= a and not b;
    layer1_outputs(2191) <= a and b;
    layer1_outputs(2192) <= not a;
    layer1_outputs(2193) <= not (a or b);
    layer1_outputs(2194) <= a and not b;
    layer1_outputs(2195) <= a;
    layer1_outputs(2196) <= not (a and b);
    layer1_outputs(2197) <= 1'b0;
    layer1_outputs(2198) <= b;
    layer1_outputs(2199) <= b;
    layer1_outputs(2200) <= 1'b1;
    layer1_outputs(2201) <= not a or b;
    layer1_outputs(2202) <= a;
    layer1_outputs(2203) <= a xor b;
    layer1_outputs(2204) <= 1'b1;
    layer1_outputs(2205) <= not (a and b);
    layer1_outputs(2206) <= not (a or b);
    layer1_outputs(2207) <= not b;
    layer1_outputs(2208) <= a and not b;
    layer1_outputs(2209) <= 1'b0;
    layer1_outputs(2210) <= not a;
    layer1_outputs(2211) <= not (a xor b);
    layer1_outputs(2212) <= not a or b;
    layer1_outputs(2213) <= not a or b;
    layer1_outputs(2214) <= a xor b;
    layer1_outputs(2215) <= a and not b;
    layer1_outputs(2216) <= a;
    layer1_outputs(2217) <= not (a or b);
    layer1_outputs(2218) <= not b;
    layer1_outputs(2219) <= a or b;
    layer1_outputs(2220) <= 1'b0;
    layer1_outputs(2221) <= a xor b;
    layer1_outputs(2222) <= a and not b;
    layer1_outputs(2223) <= 1'b1;
    layer1_outputs(2224) <= b;
    layer1_outputs(2225) <= not b or a;
    layer1_outputs(2226) <= a;
    layer1_outputs(2227) <= b;
    layer1_outputs(2228) <= a and b;
    layer1_outputs(2229) <= b;
    layer1_outputs(2230) <= b;
    layer1_outputs(2231) <= not (a or b);
    layer1_outputs(2232) <= 1'b1;
    layer1_outputs(2233) <= not a or b;
    layer1_outputs(2234) <= 1'b1;
    layer1_outputs(2235) <= 1'b0;
    layer1_outputs(2236) <= not b;
    layer1_outputs(2237) <= not a;
    layer1_outputs(2238) <= 1'b1;
    layer1_outputs(2239) <= not (a or b);
    layer1_outputs(2240) <= a and b;
    layer1_outputs(2241) <= a and not b;
    layer1_outputs(2242) <= 1'b0;
    layer1_outputs(2243) <= a and b;
    layer1_outputs(2244) <= a or b;
    layer1_outputs(2245) <= not a;
    layer1_outputs(2246) <= not (a or b);
    layer1_outputs(2247) <= a;
    layer1_outputs(2248) <= a;
    layer1_outputs(2249) <= not b or a;
    layer1_outputs(2250) <= not (a or b);
    layer1_outputs(2251) <= 1'b1;
    layer1_outputs(2252) <= 1'b0;
    layer1_outputs(2253) <= b and not a;
    layer1_outputs(2254) <= a and b;
    layer1_outputs(2255) <= a and b;
    layer1_outputs(2256) <= not a;
    layer1_outputs(2257) <= a and b;
    layer1_outputs(2258) <= 1'b0;
    layer1_outputs(2259) <= not (a xor b);
    layer1_outputs(2260) <= not a or b;
    layer1_outputs(2261) <= a or b;
    layer1_outputs(2262) <= b;
    layer1_outputs(2263) <= not (a or b);
    layer1_outputs(2264) <= not b or a;
    layer1_outputs(2265) <= not (a or b);
    layer1_outputs(2266) <= a and not b;
    layer1_outputs(2267) <= a or b;
    layer1_outputs(2268) <= b and not a;
    layer1_outputs(2269) <= not b or a;
    layer1_outputs(2270) <= 1'b1;
    layer1_outputs(2271) <= 1'b0;
    layer1_outputs(2272) <= 1'b1;
    layer1_outputs(2273) <= not (a or b);
    layer1_outputs(2274) <= 1'b0;
    layer1_outputs(2275) <= 1'b0;
    layer1_outputs(2276) <= b;
    layer1_outputs(2277) <= b;
    layer1_outputs(2278) <= not a;
    layer1_outputs(2279) <= a or b;
    layer1_outputs(2280) <= 1'b1;
    layer1_outputs(2281) <= a and b;
    layer1_outputs(2282) <= not (a and b);
    layer1_outputs(2283) <= not a;
    layer1_outputs(2284) <= not (a or b);
    layer1_outputs(2285) <= a and b;
    layer1_outputs(2286) <= b;
    layer1_outputs(2287) <= a or b;
    layer1_outputs(2288) <= not a or b;
    layer1_outputs(2289) <= not (a or b);
    layer1_outputs(2290) <= 1'b0;
    layer1_outputs(2291) <= not (a and b);
    layer1_outputs(2292) <= not a or b;
    layer1_outputs(2293) <= not b or a;
    layer1_outputs(2294) <= 1'b0;
    layer1_outputs(2295) <= not b;
    layer1_outputs(2296) <= a;
    layer1_outputs(2297) <= not (a and b);
    layer1_outputs(2298) <= 1'b1;
    layer1_outputs(2299) <= b and not a;
    layer1_outputs(2300) <= not (a or b);
    layer1_outputs(2301) <= not a;
    layer1_outputs(2302) <= not a;
    layer1_outputs(2303) <= 1'b1;
    layer1_outputs(2304) <= a or b;
    layer1_outputs(2305) <= 1'b1;
    layer1_outputs(2306) <= a xor b;
    layer1_outputs(2307) <= not b;
    layer1_outputs(2308) <= a or b;
    layer1_outputs(2309) <= 1'b1;
    layer1_outputs(2310) <= not b;
    layer1_outputs(2311) <= not b;
    layer1_outputs(2312) <= not b;
    layer1_outputs(2313) <= a or b;
    layer1_outputs(2314) <= a or b;
    layer1_outputs(2315) <= not a or b;
    layer1_outputs(2316) <= not b;
    layer1_outputs(2317) <= b and not a;
    layer1_outputs(2318) <= 1'b0;
    layer1_outputs(2319) <= not (a and b);
    layer1_outputs(2320) <= not b;
    layer1_outputs(2321) <= b;
    layer1_outputs(2322) <= not (a and b);
    layer1_outputs(2323) <= not (a xor b);
    layer1_outputs(2324) <= not (a and b);
    layer1_outputs(2325) <= a xor b;
    layer1_outputs(2326) <= 1'b1;
    layer1_outputs(2327) <= a or b;
    layer1_outputs(2328) <= a or b;
    layer1_outputs(2329) <= not b or a;
    layer1_outputs(2330) <= a xor b;
    layer1_outputs(2331) <= a and not b;
    layer1_outputs(2332) <= not (a or b);
    layer1_outputs(2333) <= a or b;
    layer1_outputs(2334) <= b and not a;
    layer1_outputs(2335) <= a or b;
    layer1_outputs(2336) <= not a or b;
    layer1_outputs(2337) <= not a or b;
    layer1_outputs(2338) <= not b;
    layer1_outputs(2339) <= not (a and b);
    layer1_outputs(2340) <= 1'b0;
    layer1_outputs(2341) <= a and not b;
    layer1_outputs(2342) <= not b or a;
    layer1_outputs(2343) <= a and not b;
    layer1_outputs(2344) <= 1'b1;
    layer1_outputs(2345) <= 1'b0;
    layer1_outputs(2346) <= not (a or b);
    layer1_outputs(2347) <= not a or b;
    layer1_outputs(2348) <= 1'b0;
    layer1_outputs(2349) <= a and not b;
    layer1_outputs(2350) <= not (a or b);
    layer1_outputs(2351) <= not b or a;
    layer1_outputs(2352) <= b and not a;
    layer1_outputs(2353) <= 1'b0;
    layer1_outputs(2354) <= 1'b0;
    layer1_outputs(2355) <= not b or a;
    layer1_outputs(2356) <= a or b;
    layer1_outputs(2357) <= a;
    layer1_outputs(2358) <= b;
    layer1_outputs(2359) <= not (a xor b);
    layer1_outputs(2360) <= 1'b1;
    layer1_outputs(2361) <= not b;
    layer1_outputs(2362) <= a and b;
    layer1_outputs(2363) <= a and not b;
    layer1_outputs(2364) <= a and not b;
    layer1_outputs(2365) <= 1'b1;
    layer1_outputs(2366) <= a and not b;
    layer1_outputs(2367) <= a xor b;
    layer1_outputs(2368) <= not b or a;
    layer1_outputs(2369) <= 1'b1;
    layer1_outputs(2370) <= not a;
    layer1_outputs(2371) <= not b or a;
    layer1_outputs(2372) <= not a or b;
    layer1_outputs(2373) <= 1'b0;
    layer1_outputs(2374) <= 1'b0;
    layer1_outputs(2375) <= a and not b;
    layer1_outputs(2376) <= 1'b0;
    layer1_outputs(2377) <= not a or b;
    layer1_outputs(2378) <= a or b;
    layer1_outputs(2379) <= a;
    layer1_outputs(2380) <= a or b;
    layer1_outputs(2381) <= a or b;
    layer1_outputs(2382) <= not a;
    layer1_outputs(2383) <= not b or a;
    layer1_outputs(2384) <= not a or b;
    layer1_outputs(2385) <= 1'b0;
    layer1_outputs(2386) <= not (a xor b);
    layer1_outputs(2387) <= a;
    layer1_outputs(2388) <= 1'b0;
    layer1_outputs(2389) <= not (a and b);
    layer1_outputs(2390) <= not a or b;
    layer1_outputs(2391) <= a;
    layer1_outputs(2392) <= 1'b1;
    layer1_outputs(2393) <= b and not a;
    layer1_outputs(2394) <= a or b;
    layer1_outputs(2395) <= a;
    layer1_outputs(2396) <= a or b;
    layer1_outputs(2397) <= a and not b;
    layer1_outputs(2398) <= not b or a;
    layer1_outputs(2399) <= a;
    layer1_outputs(2400) <= not b;
    layer1_outputs(2401) <= a and not b;
    layer1_outputs(2402) <= b and not a;
    layer1_outputs(2403) <= a;
    layer1_outputs(2404) <= not b or a;
    layer1_outputs(2405) <= not (a and b);
    layer1_outputs(2406) <= a xor b;
    layer1_outputs(2407) <= 1'b0;
    layer1_outputs(2408) <= a or b;
    layer1_outputs(2409) <= not b or a;
    layer1_outputs(2410) <= not (a or b);
    layer1_outputs(2411) <= not b;
    layer1_outputs(2412) <= b and not a;
    layer1_outputs(2413) <= not a or b;
    layer1_outputs(2414) <= 1'b1;
    layer1_outputs(2415) <= not b or a;
    layer1_outputs(2416) <= a and not b;
    layer1_outputs(2417) <= not (a or b);
    layer1_outputs(2418) <= a;
    layer1_outputs(2419) <= not (a or b);
    layer1_outputs(2420) <= a and not b;
    layer1_outputs(2421) <= not b;
    layer1_outputs(2422) <= not a;
    layer1_outputs(2423) <= not b or a;
    layer1_outputs(2424) <= b;
    layer1_outputs(2425) <= 1'b0;
    layer1_outputs(2426) <= a and b;
    layer1_outputs(2427) <= not (a and b);
    layer1_outputs(2428) <= not (a xor b);
    layer1_outputs(2429) <= a or b;
    layer1_outputs(2430) <= not a;
    layer1_outputs(2431) <= b and not a;
    layer1_outputs(2432) <= not a or b;
    layer1_outputs(2433) <= b and not a;
    layer1_outputs(2434) <= a xor b;
    layer1_outputs(2435) <= a or b;
    layer1_outputs(2436) <= b;
    layer1_outputs(2437) <= 1'b0;
    layer1_outputs(2438) <= b and not a;
    layer1_outputs(2439) <= a and not b;
    layer1_outputs(2440) <= 1'b0;
    layer1_outputs(2441) <= a and not b;
    layer1_outputs(2442) <= a and not b;
    layer1_outputs(2443) <= 1'b0;
    layer1_outputs(2444) <= 1'b1;
    layer1_outputs(2445) <= 1'b0;
    layer1_outputs(2446) <= not b or a;
    layer1_outputs(2447) <= not (a or b);
    layer1_outputs(2448) <= not (a and b);
    layer1_outputs(2449) <= 1'b1;
    layer1_outputs(2450) <= 1'b1;
    layer1_outputs(2451) <= a or b;
    layer1_outputs(2452) <= not (a and b);
    layer1_outputs(2453) <= not a;
    layer1_outputs(2454) <= 1'b1;
    layer1_outputs(2455) <= a;
    layer1_outputs(2456) <= not (a or b);
    layer1_outputs(2457) <= 1'b0;
    layer1_outputs(2458) <= 1'b0;
    layer1_outputs(2459) <= 1'b1;
    layer1_outputs(2460) <= b and not a;
    layer1_outputs(2461) <= a xor b;
    layer1_outputs(2462) <= not (a or b);
    layer1_outputs(2463) <= a or b;
    layer1_outputs(2464) <= a or b;
    layer1_outputs(2465) <= b;
    layer1_outputs(2466) <= 1'b1;
    layer1_outputs(2467) <= not (a xor b);
    layer1_outputs(2468) <= not a;
    layer1_outputs(2469) <= 1'b0;
    layer1_outputs(2470) <= a and not b;
    layer1_outputs(2471) <= 1'b0;
    layer1_outputs(2472) <= a and not b;
    layer1_outputs(2473) <= a and b;
    layer1_outputs(2474) <= 1'b0;
    layer1_outputs(2475) <= not (a xor b);
    layer1_outputs(2476) <= a and b;
    layer1_outputs(2477) <= not b;
    layer1_outputs(2478) <= not b or a;
    layer1_outputs(2479) <= a or b;
    layer1_outputs(2480) <= not (a or b);
    layer1_outputs(2481) <= not (a or b);
    layer1_outputs(2482) <= not (a or b);
    layer1_outputs(2483) <= not (a xor b);
    layer1_outputs(2484) <= 1'b0;
    layer1_outputs(2485) <= not (a and b);
    layer1_outputs(2486) <= 1'b1;
    layer1_outputs(2487) <= not (a or b);
    layer1_outputs(2488) <= a;
    layer1_outputs(2489) <= not b or a;
    layer1_outputs(2490) <= not a;
    layer1_outputs(2491) <= a and not b;
    layer1_outputs(2492) <= not (a or b);
    layer1_outputs(2493) <= a or b;
    layer1_outputs(2494) <= not (a or b);
    layer1_outputs(2495) <= 1'b1;
    layer1_outputs(2496) <= a;
    layer1_outputs(2497) <= not b;
    layer1_outputs(2498) <= b and not a;
    layer1_outputs(2499) <= 1'b0;
    layer1_outputs(2500) <= not a;
    layer1_outputs(2501) <= a and b;
    layer1_outputs(2502) <= b;
    layer1_outputs(2503) <= not (a or b);
    layer1_outputs(2504) <= not (a or b);
    layer1_outputs(2505) <= a or b;
    layer1_outputs(2506) <= 1'b0;
    layer1_outputs(2507) <= not (a or b);
    layer1_outputs(2508) <= not a;
    layer1_outputs(2509) <= a and not b;
    layer1_outputs(2510) <= not (a or b);
    layer1_outputs(2511) <= 1'b0;
    layer1_outputs(2512) <= not b or a;
    layer1_outputs(2513) <= b;
    layer1_outputs(2514) <= 1'b0;
    layer1_outputs(2515) <= a and not b;
    layer1_outputs(2516) <= not a or b;
    layer1_outputs(2517) <= not a;
    layer1_outputs(2518) <= not b or a;
    layer1_outputs(2519) <= a and not b;
    layer1_outputs(2520) <= a and not b;
    layer1_outputs(2521) <= 1'b1;
    layer1_outputs(2522) <= a and not b;
    layer1_outputs(2523) <= b and not a;
    layer1_outputs(2524) <= b and not a;
    layer1_outputs(2525) <= not (a or b);
    layer1_outputs(2526) <= 1'b0;
    layer1_outputs(2527) <= a;
    layer1_outputs(2528) <= not b;
    layer1_outputs(2529) <= a;
    layer1_outputs(2530) <= 1'b1;
    layer1_outputs(2531) <= not b;
    layer1_outputs(2532) <= 1'b1;
    layer1_outputs(2533) <= 1'b0;
    layer1_outputs(2534) <= 1'b1;
    layer1_outputs(2535) <= 1'b1;
    layer1_outputs(2536) <= a;
    layer1_outputs(2537) <= 1'b0;
    layer1_outputs(2538) <= b and not a;
    layer1_outputs(2539) <= a;
    layer1_outputs(2540) <= not a or b;
    layer1_outputs(2541) <= 1'b1;
    layer1_outputs(2542) <= a;
    layer1_outputs(2543) <= not (a and b);
    layer1_outputs(2544) <= a and b;
    layer1_outputs(2545) <= 1'b1;
    layer1_outputs(2546) <= a or b;
    layer1_outputs(2547) <= a and not b;
    layer1_outputs(2548) <= not (a xor b);
    layer1_outputs(2549) <= a or b;
    layer1_outputs(2550) <= b and not a;
    layer1_outputs(2551) <= not b;
    layer1_outputs(2552) <= 1'b0;
    layer1_outputs(2553) <= not b;
    layer1_outputs(2554) <= not (a or b);
    layer1_outputs(2555) <= a or b;
    layer1_outputs(2556) <= 1'b1;
    layer1_outputs(2557) <= a xor b;
    layer1_outputs(2558) <= not b or a;
    layer1_outputs(2559) <= 1'b0;
    layer2_outputs(0) <= b and not a;
    layer2_outputs(1) <= 1'b1;
    layer2_outputs(2) <= a;
    layer2_outputs(3) <= b and not a;
    layer2_outputs(4) <= b and not a;
    layer2_outputs(5) <= a xor b;
    layer2_outputs(6) <= a and not b;
    layer2_outputs(7) <= 1'b0;
    layer2_outputs(8) <= b and not a;
    layer2_outputs(9) <= 1'b1;
    layer2_outputs(10) <= b;
    layer2_outputs(11) <= not a;
    layer2_outputs(12) <= b and not a;
    layer2_outputs(13) <= a and b;
    layer2_outputs(14) <= a and b;
    layer2_outputs(15) <= not b;
    layer2_outputs(16) <= not b;
    layer2_outputs(17) <= not (a and b);
    layer2_outputs(18) <= a or b;
    layer2_outputs(19) <= 1'b0;
    layer2_outputs(20) <= not a or b;
    layer2_outputs(21) <= b and not a;
    layer2_outputs(22) <= b and not a;
    layer2_outputs(23) <= not (a or b);
    layer2_outputs(24) <= not a or b;
    layer2_outputs(25) <= not (a and b);
    layer2_outputs(26) <= b;
    layer2_outputs(27) <= a or b;
    layer2_outputs(28) <= 1'b0;
    layer2_outputs(29) <= a;
    layer2_outputs(30) <= 1'b0;
    layer2_outputs(31) <= 1'b1;
    layer2_outputs(32) <= 1'b0;
    layer2_outputs(33) <= not a or b;
    layer2_outputs(34) <= not a;
    layer2_outputs(35) <= 1'b0;
    layer2_outputs(36) <= not b;
    layer2_outputs(37) <= a or b;
    layer2_outputs(38) <= a and b;
    layer2_outputs(39) <= not a or b;
    layer2_outputs(40) <= not (a and b);
    layer2_outputs(41) <= 1'b0;
    layer2_outputs(42) <= a and not b;
    layer2_outputs(43) <= 1'b0;
    layer2_outputs(44) <= a and not b;
    layer2_outputs(45) <= not (a xor b);
    layer2_outputs(46) <= 1'b0;
    layer2_outputs(47) <= not (a and b);
    layer2_outputs(48) <= b;
    layer2_outputs(49) <= a and b;
    layer2_outputs(50) <= 1'b0;
    layer2_outputs(51) <= not (a and b);
    layer2_outputs(52) <= 1'b1;
    layer2_outputs(53) <= 1'b1;
    layer2_outputs(54) <= not a;
    layer2_outputs(55) <= b;
    layer2_outputs(56) <= not b;
    layer2_outputs(57) <= a;
    layer2_outputs(58) <= 1'b0;
    layer2_outputs(59) <= not a;
    layer2_outputs(60) <= not (a or b);
    layer2_outputs(61) <= not b or a;
    layer2_outputs(62) <= 1'b0;
    layer2_outputs(63) <= not a;
    layer2_outputs(64) <= not b or a;
    layer2_outputs(65) <= a;
    layer2_outputs(66) <= a and not b;
    layer2_outputs(67) <= not b;
    layer2_outputs(68) <= not a;
    layer2_outputs(69) <= a or b;
    layer2_outputs(70) <= b and not a;
    layer2_outputs(71) <= not (a and b);
    layer2_outputs(72) <= 1'b0;
    layer2_outputs(73) <= not b;
    layer2_outputs(74) <= a or b;
    layer2_outputs(75) <= not a or b;
    layer2_outputs(76) <= not a or b;
    layer2_outputs(77) <= 1'b1;
    layer2_outputs(78) <= 1'b1;
    layer2_outputs(79) <= b and not a;
    layer2_outputs(80) <= a and not b;
    layer2_outputs(81) <= not a or b;
    layer2_outputs(82) <= a xor b;
    layer2_outputs(83) <= a and b;
    layer2_outputs(84) <= a and not b;
    layer2_outputs(85) <= 1'b1;
    layer2_outputs(86) <= not b;
    layer2_outputs(87) <= a;
    layer2_outputs(88) <= 1'b0;
    layer2_outputs(89) <= 1'b1;
    layer2_outputs(90) <= a;
    layer2_outputs(91) <= not b;
    layer2_outputs(92) <= a and b;
    layer2_outputs(93) <= not (a or b);
    layer2_outputs(94) <= not (a or b);
    layer2_outputs(95) <= not (a or b);
    layer2_outputs(96) <= not (a and b);
    layer2_outputs(97) <= 1'b0;
    layer2_outputs(98) <= not b;
    layer2_outputs(99) <= 1'b0;
    layer2_outputs(100) <= 1'b1;
    layer2_outputs(101) <= not a;
    layer2_outputs(102) <= not b or a;
    layer2_outputs(103) <= a or b;
    layer2_outputs(104) <= a and not b;
    layer2_outputs(105) <= 1'b0;
    layer2_outputs(106) <= a and not b;
    layer2_outputs(107) <= a;
    layer2_outputs(108) <= not b;
    layer2_outputs(109) <= a and b;
    layer2_outputs(110) <= a or b;
    layer2_outputs(111) <= 1'b1;
    layer2_outputs(112) <= a or b;
    layer2_outputs(113) <= not a;
    layer2_outputs(114) <= a and not b;
    layer2_outputs(115) <= not a or b;
    layer2_outputs(116) <= 1'b1;
    layer2_outputs(117) <= not b;
    layer2_outputs(118) <= not b;
    layer2_outputs(119) <= a and b;
    layer2_outputs(120) <= not (a xor b);
    layer2_outputs(121) <= not b or a;
    layer2_outputs(122) <= not a or b;
    layer2_outputs(123) <= not (a and b);
    layer2_outputs(124) <= b and not a;
    layer2_outputs(125) <= b and not a;
    layer2_outputs(126) <= 1'b0;
    layer2_outputs(127) <= 1'b0;
    layer2_outputs(128) <= b and not a;
    layer2_outputs(129) <= a and not b;
    layer2_outputs(130) <= not (a or b);
    layer2_outputs(131) <= not (a or b);
    layer2_outputs(132) <= a and b;
    layer2_outputs(133) <= not b;
    layer2_outputs(134) <= not a or b;
    layer2_outputs(135) <= 1'b1;
    layer2_outputs(136) <= not a or b;
    layer2_outputs(137) <= b;
    layer2_outputs(138) <= b;
    layer2_outputs(139) <= b;
    layer2_outputs(140) <= 1'b0;
    layer2_outputs(141) <= a and not b;
    layer2_outputs(142) <= not (a or b);
    layer2_outputs(143) <= not a;
    layer2_outputs(144) <= a or b;
    layer2_outputs(145) <= a or b;
    layer2_outputs(146) <= a;
    layer2_outputs(147) <= not (a xor b);
    layer2_outputs(148) <= not a or b;
    layer2_outputs(149) <= 1'b1;
    layer2_outputs(150) <= a or b;
    layer2_outputs(151) <= not (a and b);
    layer2_outputs(152) <= 1'b0;
    layer2_outputs(153) <= not (a or b);
    layer2_outputs(154) <= a and not b;
    layer2_outputs(155) <= 1'b1;
    layer2_outputs(156) <= not a or b;
    layer2_outputs(157) <= not b or a;
    layer2_outputs(158) <= a xor b;
    layer2_outputs(159) <= a and not b;
    layer2_outputs(160) <= 1'b0;
    layer2_outputs(161) <= a and b;
    layer2_outputs(162) <= not b or a;
    layer2_outputs(163) <= not (a and b);
    layer2_outputs(164) <= a and not b;
    layer2_outputs(165) <= b;
    layer2_outputs(166) <= a or b;
    layer2_outputs(167) <= not a or b;
    layer2_outputs(168) <= not b;
    layer2_outputs(169) <= not a;
    layer2_outputs(170) <= a and not b;
    layer2_outputs(171) <= b;
    layer2_outputs(172) <= 1'b1;
    layer2_outputs(173) <= not b;
    layer2_outputs(174) <= a;
    layer2_outputs(175) <= not (a or b);
    layer2_outputs(176) <= not b or a;
    layer2_outputs(177) <= not a or b;
    layer2_outputs(178) <= 1'b0;
    layer2_outputs(179) <= not b or a;
    layer2_outputs(180) <= a;
    layer2_outputs(181) <= a;
    layer2_outputs(182) <= not b;
    layer2_outputs(183) <= 1'b1;
    layer2_outputs(184) <= not a;
    layer2_outputs(185) <= b;
    layer2_outputs(186) <= b and not a;
    layer2_outputs(187) <= b and not a;
    layer2_outputs(188) <= not (a and b);
    layer2_outputs(189) <= 1'b1;
    layer2_outputs(190) <= not b;
    layer2_outputs(191) <= a and b;
    layer2_outputs(192) <= b and not a;
    layer2_outputs(193) <= 1'b1;
    layer2_outputs(194) <= 1'b0;
    layer2_outputs(195) <= a and b;
    layer2_outputs(196) <= not a or b;
    layer2_outputs(197) <= 1'b0;
    layer2_outputs(198) <= not a;
    layer2_outputs(199) <= not b;
    layer2_outputs(200) <= a or b;
    layer2_outputs(201) <= a or b;
    layer2_outputs(202) <= not (a xor b);
    layer2_outputs(203) <= a;
    layer2_outputs(204) <= b and not a;
    layer2_outputs(205) <= b and not a;
    layer2_outputs(206) <= a;
    layer2_outputs(207) <= 1'b0;
    layer2_outputs(208) <= 1'b1;
    layer2_outputs(209) <= b and not a;
    layer2_outputs(210) <= 1'b0;
    layer2_outputs(211) <= not b;
    layer2_outputs(212) <= not (a or b);
    layer2_outputs(213) <= 1'b1;
    layer2_outputs(214) <= a and b;
    layer2_outputs(215) <= b;
    layer2_outputs(216) <= not (a and b);
    layer2_outputs(217) <= not (a or b);
    layer2_outputs(218) <= a and not b;
    layer2_outputs(219) <= not b;
    layer2_outputs(220) <= a and not b;
    layer2_outputs(221) <= not (a and b);
    layer2_outputs(222) <= not a or b;
    layer2_outputs(223) <= not a;
    layer2_outputs(224) <= b and not a;
    layer2_outputs(225) <= 1'b0;
    layer2_outputs(226) <= b and not a;
    layer2_outputs(227) <= a or b;
    layer2_outputs(228) <= a;
    layer2_outputs(229) <= 1'b1;
    layer2_outputs(230) <= a and not b;
    layer2_outputs(231) <= a and b;
    layer2_outputs(232) <= a;
    layer2_outputs(233) <= not a or b;
    layer2_outputs(234) <= 1'b1;
    layer2_outputs(235) <= b;
    layer2_outputs(236) <= not b;
    layer2_outputs(237) <= not a or b;
    layer2_outputs(238) <= b;
    layer2_outputs(239) <= a;
    layer2_outputs(240) <= not a or b;
    layer2_outputs(241) <= not a or b;
    layer2_outputs(242) <= not (a or b);
    layer2_outputs(243) <= a and b;
    layer2_outputs(244) <= not a;
    layer2_outputs(245) <= 1'b1;
    layer2_outputs(246) <= b and not a;
    layer2_outputs(247) <= a;
    layer2_outputs(248) <= 1'b0;
    layer2_outputs(249) <= not a;
    layer2_outputs(250) <= 1'b1;
    layer2_outputs(251) <= not (a or b);
    layer2_outputs(252) <= 1'b1;
    layer2_outputs(253) <= 1'b0;
    layer2_outputs(254) <= 1'b0;
    layer2_outputs(255) <= b and not a;
    layer2_outputs(256) <= a xor b;
    layer2_outputs(257) <= a and not b;
    layer2_outputs(258) <= a and b;
    layer2_outputs(259) <= b and not a;
    layer2_outputs(260) <= not (a or b);
    layer2_outputs(261) <= not b;
    layer2_outputs(262) <= not a;
    layer2_outputs(263) <= not a;
    layer2_outputs(264) <= 1'b0;
    layer2_outputs(265) <= 1'b1;
    layer2_outputs(266) <= a or b;
    layer2_outputs(267) <= b and not a;
    layer2_outputs(268) <= a;
    layer2_outputs(269) <= 1'b1;
    layer2_outputs(270) <= b;
    layer2_outputs(271) <= 1'b1;
    layer2_outputs(272) <= 1'b1;
    layer2_outputs(273) <= not (a and b);
    layer2_outputs(274) <= a and not b;
    layer2_outputs(275) <= not b;
    layer2_outputs(276) <= b;
    layer2_outputs(277) <= not (a or b);
    layer2_outputs(278) <= not (a or b);
    layer2_outputs(279) <= not (a and b);
    layer2_outputs(280) <= not (a and b);
    layer2_outputs(281) <= a and b;
    layer2_outputs(282) <= a xor b;
    layer2_outputs(283) <= 1'b1;
    layer2_outputs(284) <= not (a or b);
    layer2_outputs(285) <= not b;
    layer2_outputs(286) <= a or b;
    layer2_outputs(287) <= a and not b;
    layer2_outputs(288) <= a and not b;
    layer2_outputs(289) <= 1'b1;
    layer2_outputs(290) <= 1'b0;
    layer2_outputs(291) <= a or b;
    layer2_outputs(292) <= not (a or b);
    layer2_outputs(293) <= 1'b1;
    layer2_outputs(294) <= a and b;
    layer2_outputs(295) <= not a;
    layer2_outputs(296) <= a or b;
    layer2_outputs(297) <= not b or a;
    layer2_outputs(298) <= a;
    layer2_outputs(299) <= b and not a;
    layer2_outputs(300) <= not b;
    layer2_outputs(301) <= not a or b;
    layer2_outputs(302) <= a;
    layer2_outputs(303) <= 1'b1;
    layer2_outputs(304) <= a and b;
    layer2_outputs(305) <= a or b;
    layer2_outputs(306) <= not b or a;
    layer2_outputs(307) <= a or b;
    layer2_outputs(308) <= 1'b0;
    layer2_outputs(309) <= not b;
    layer2_outputs(310) <= 1'b0;
    layer2_outputs(311) <= not (a and b);
    layer2_outputs(312) <= not (a and b);
    layer2_outputs(313) <= not (a or b);
    layer2_outputs(314) <= b;
    layer2_outputs(315) <= a and b;
    layer2_outputs(316) <= a or b;
    layer2_outputs(317) <= not a;
    layer2_outputs(318) <= b and not a;
    layer2_outputs(319) <= 1'b0;
    layer2_outputs(320) <= 1'b0;
    layer2_outputs(321) <= a and not b;
    layer2_outputs(322) <= not (a or b);
    layer2_outputs(323) <= 1'b1;
    layer2_outputs(324) <= 1'b0;
    layer2_outputs(325) <= not (a or b);
    layer2_outputs(326) <= not (a xor b);
    layer2_outputs(327) <= not a;
    layer2_outputs(328) <= a and not b;
    layer2_outputs(329) <= not b or a;
    layer2_outputs(330) <= a;
    layer2_outputs(331) <= a and b;
    layer2_outputs(332) <= b;
    layer2_outputs(333) <= not (a and b);
    layer2_outputs(334) <= a or b;
    layer2_outputs(335) <= a and b;
    layer2_outputs(336) <= b and not a;
    layer2_outputs(337) <= a and not b;
    layer2_outputs(338) <= 1'b0;
    layer2_outputs(339) <= a;
    layer2_outputs(340) <= b and not a;
    layer2_outputs(341) <= b and not a;
    layer2_outputs(342) <= not b or a;
    layer2_outputs(343) <= b and not a;
    layer2_outputs(344) <= not (a and b);
    layer2_outputs(345) <= 1'b0;
    layer2_outputs(346) <= a and not b;
    layer2_outputs(347) <= not b or a;
    layer2_outputs(348) <= not b or a;
    layer2_outputs(349) <= a or b;
    layer2_outputs(350) <= not a;
    layer2_outputs(351) <= 1'b0;
    layer2_outputs(352) <= a and b;
    layer2_outputs(353) <= a and not b;
    layer2_outputs(354) <= not b;
    layer2_outputs(355) <= a and not b;
    layer2_outputs(356) <= a and b;
    layer2_outputs(357) <= a;
    layer2_outputs(358) <= not a or b;
    layer2_outputs(359) <= b;
    layer2_outputs(360) <= not b;
    layer2_outputs(361) <= a and not b;
    layer2_outputs(362) <= not b or a;
    layer2_outputs(363) <= a and b;
    layer2_outputs(364) <= not (a or b);
    layer2_outputs(365) <= not (a or b);
    layer2_outputs(366) <= not b or a;
    layer2_outputs(367) <= b and not a;
    layer2_outputs(368) <= not a;
    layer2_outputs(369) <= not a;
    layer2_outputs(370) <= 1'b0;
    layer2_outputs(371) <= a;
    layer2_outputs(372) <= not b or a;
    layer2_outputs(373) <= a and not b;
    layer2_outputs(374) <= not b;
    layer2_outputs(375) <= a or b;
    layer2_outputs(376) <= 1'b1;
    layer2_outputs(377) <= a xor b;
    layer2_outputs(378) <= a or b;
    layer2_outputs(379) <= a and b;
    layer2_outputs(380) <= not a or b;
    layer2_outputs(381) <= 1'b0;
    layer2_outputs(382) <= not (a or b);
    layer2_outputs(383) <= not (a or b);
    layer2_outputs(384) <= b and not a;
    layer2_outputs(385) <= not b;
    layer2_outputs(386) <= 1'b1;
    layer2_outputs(387) <= not (a and b);
    layer2_outputs(388) <= 1'b1;
    layer2_outputs(389) <= not b;
    layer2_outputs(390) <= not (a or b);
    layer2_outputs(391) <= a and b;
    layer2_outputs(392) <= not b;
    layer2_outputs(393) <= a and not b;
    layer2_outputs(394) <= not a;
    layer2_outputs(395) <= 1'b1;
    layer2_outputs(396) <= not a;
    layer2_outputs(397) <= a and b;
    layer2_outputs(398) <= not (a and b);
    layer2_outputs(399) <= a or b;
    layer2_outputs(400) <= a and b;
    layer2_outputs(401) <= 1'b0;
    layer2_outputs(402) <= not a or b;
    layer2_outputs(403) <= not a or b;
    layer2_outputs(404) <= 1'b0;
    layer2_outputs(405) <= b;
    layer2_outputs(406) <= not b or a;
    layer2_outputs(407) <= a and not b;
    layer2_outputs(408) <= a or b;
    layer2_outputs(409) <= a xor b;
    layer2_outputs(410) <= not a;
    layer2_outputs(411) <= 1'b1;
    layer2_outputs(412) <= not (a and b);
    layer2_outputs(413) <= a and not b;
    layer2_outputs(414) <= not a;
    layer2_outputs(415) <= b;
    layer2_outputs(416) <= 1'b0;
    layer2_outputs(417) <= 1'b0;
    layer2_outputs(418) <= a;
    layer2_outputs(419) <= not a or b;
    layer2_outputs(420) <= a and not b;
    layer2_outputs(421) <= a or b;
    layer2_outputs(422) <= 1'b1;
    layer2_outputs(423) <= a and not b;
    layer2_outputs(424) <= not (a and b);
    layer2_outputs(425) <= b and not a;
    layer2_outputs(426) <= 1'b1;
    layer2_outputs(427) <= not (a and b);
    layer2_outputs(428) <= b;
    layer2_outputs(429) <= not (a and b);
    layer2_outputs(430) <= a;
    layer2_outputs(431) <= 1'b1;
    layer2_outputs(432) <= not a;
    layer2_outputs(433) <= a;
    layer2_outputs(434) <= not a or b;
    layer2_outputs(435) <= b and not a;
    layer2_outputs(436) <= not a or b;
    layer2_outputs(437) <= not a;
    layer2_outputs(438) <= not a or b;
    layer2_outputs(439) <= a or b;
    layer2_outputs(440) <= a and not b;
    layer2_outputs(441) <= b and not a;
    layer2_outputs(442) <= 1'b1;
    layer2_outputs(443) <= b;
    layer2_outputs(444) <= not a;
    layer2_outputs(445) <= not b;
    layer2_outputs(446) <= 1'b0;
    layer2_outputs(447) <= a and not b;
    layer2_outputs(448) <= not a;
    layer2_outputs(449) <= 1'b0;
    layer2_outputs(450) <= not a or b;
    layer2_outputs(451) <= not b or a;
    layer2_outputs(452) <= not b;
    layer2_outputs(453) <= not b or a;
    layer2_outputs(454) <= not a or b;
    layer2_outputs(455) <= not a;
    layer2_outputs(456) <= not a or b;
    layer2_outputs(457) <= not a;
    layer2_outputs(458) <= a xor b;
    layer2_outputs(459) <= not a;
    layer2_outputs(460) <= a;
    layer2_outputs(461) <= 1'b1;
    layer2_outputs(462) <= a;
    layer2_outputs(463) <= not a or b;
    layer2_outputs(464) <= 1'b0;
    layer2_outputs(465) <= a and b;
    layer2_outputs(466) <= not (a and b);
    layer2_outputs(467) <= not (a or b);
    layer2_outputs(468) <= 1'b1;
    layer2_outputs(469) <= not (a and b);
    layer2_outputs(470) <= a and b;
    layer2_outputs(471) <= not b or a;
    layer2_outputs(472) <= b;
    layer2_outputs(473) <= not a or b;
    layer2_outputs(474) <= a;
    layer2_outputs(475) <= not b or a;
    layer2_outputs(476) <= not b or a;
    layer2_outputs(477) <= a and not b;
    layer2_outputs(478) <= not a or b;
    layer2_outputs(479) <= not (a and b);
    layer2_outputs(480) <= not b;
    layer2_outputs(481) <= not b;
    layer2_outputs(482) <= a and b;
    layer2_outputs(483) <= a and not b;
    layer2_outputs(484) <= not a or b;
    layer2_outputs(485) <= a;
    layer2_outputs(486) <= not (a and b);
    layer2_outputs(487) <= a or b;
    layer2_outputs(488) <= 1'b1;
    layer2_outputs(489) <= not a or b;
    layer2_outputs(490) <= not b;
    layer2_outputs(491) <= 1'b1;
    layer2_outputs(492) <= 1'b1;
    layer2_outputs(493) <= b and not a;
    layer2_outputs(494) <= 1'b0;
    layer2_outputs(495) <= not b or a;
    layer2_outputs(496) <= not (a and b);
    layer2_outputs(497) <= a;
    layer2_outputs(498) <= a and not b;
    layer2_outputs(499) <= 1'b1;
    layer2_outputs(500) <= a and b;
    layer2_outputs(501) <= b and not a;
    layer2_outputs(502) <= a or b;
    layer2_outputs(503) <= a or b;
    layer2_outputs(504) <= 1'b0;
    layer2_outputs(505) <= not b;
    layer2_outputs(506) <= a and b;
    layer2_outputs(507) <= 1'b0;
    layer2_outputs(508) <= b and not a;
    layer2_outputs(509) <= a and b;
    layer2_outputs(510) <= not b;
    layer2_outputs(511) <= 1'b0;
    layer2_outputs(512) <= b and not a;
    layer2_outputs(513) <= 1'b0;
    layer2_outputs(514) <= a and b;
    layer2_outputs(515) <= a and not b;
    layer2_outputs(516) <= not (a or b);
    layer2_outputs(517) <= not b;
    layer2_outputs(518) <= not a;
    layer2_outputs(519) <= a;
    layer2_outputs(520) <= a and b;
    layer2_outputs(521) <= 1'b1;
    layer2_outputs(522) <= not (a or b);
    layer2_outputs(523) <= b and not a;
    layer2_outputs(524) <= 1'b0;
    layer2_outputs(525) <= not (a or b);
    layer2_outputs(526) <= a and b;
    layer2_outputs(527) <= not b or a;
    layer2_outputs(528) <= 1'b1;
    layer2_outputs(529) <= a and not b;
    layer2_outputs(530) <= a and b;
    layer2_outputs(531) <= b and not a;
    layer2_outputs(532) <= not b or a;
    layer2_outputs(533) <= a or b;
    layer2_outputs(534) <= b;
    layer2_outputs(535) <= a and not b;
    layer2_outputs(536) <= 1'b1;
    layer2_outputs(537) <= a and not b;
    layer2_outputs(538) <= a;
    layer2_outputs(539) <= 1'b0;
    layer2_outputs(540) <= not b;
    layer2_outputs(541) <= not b or a;
    layer2_outputs(542) <= not b or a;
    layer2_outputs(543) <= not (a and b);
    layer2_outputs(544) <= not (a and b);
    layer2_outputs(545) <= not (a and b);
    layer2_outputs(546) <= not (a and b);
    layer2_outputs(547) <= a or b;
    layer2_outputs(548) <= b and not a;
    layer2_outputs(549) <= b;
    layer2_outputs(550) <= a and not b;
    layer2_outputs(551) <= 1'b1;
    layer2_outputs(552) <= not b or a;
    layer2_outputs(553) <= 1'b0;
    layer2_outputs(554) <= a and not b;
    layer2_outputs(555) <= b and not a;
    layer2_outputs(556) <= not b;
    layer2_outputs(557) <= b and not a;
    layer2_outputs(558) <= not b or a;
    layer2_outputs(559) <= 1'b1;
    layer2_outputs(560) <= not (a xor b);
    layer2_outputs(561) <= b;
    layer2_outputs(562) <= not (a or b);
    layer2_outputs(563) <= not (a or b);
    layer2_outputs(564) <= 1'b0;
    layer2_outputs(565) <= a or b;
    layer2_outputs(566) <= not (a and b);
    layer2_outputs(567) <= a and not b;
    layer2_outputs(568) <= a and b;
    layer2_outputs(569) <= 1'b1;
    layer2_outputs(570) <= 1'b0;
    layer2_outputs(571) <= not (a or b);
    layer2_outputs(572) <= not b or a;
    layer2_outputs(573) <= a and not b;
    layer2_outputs(574) <= 1'b1;
    layer2_outputs(575) <= not (a or b);
    layer2_outputs(576) <= 1'b1;
    layer2_outputs(577) <= 1'b1;
    layer2_outputs(578) <= not (a or b);
    layer2_outputs(579) <= 1'b1;
    layer2_outputs(580) <= not a or b;
    layer2_outputs(581) <= 1'b1;
    layer2_outputs(582) <= 1'b0;
    layer2_outputs(583) <= 1'b1;
    layer2_outputs(584) <= not (a and b);
    layer2_outputs(585) <= not b or a;
    layer2_outputs(586) <= b and not a;
    layer2_outputs(587) <= a or b;
    layer2_outputs(588) <= not b;
    layer2_outputs(589) <= not (a or b);
    layer2_outputs(590) <= a or b;
    layer2_outputs(591) <= a and b;
    layer2_outputs(592) <= not (a or b);
    layer2_outputs(593) <= 1'b0;
    layer2_outputs(594) <= a and not b;
    layer2_outputs(595) <= not (a or b);
    layer2_outputs(596) <= b and not a;
    layer2_outputs(597) <= not b;
    layer2_outputs(598) <= b and not a;
    layer2_outputs(599) <= not (a and b);
    layer2_outputs(600) <= b and not a;
    layer2_outputs(601) <= 1'b0;
    layer2_outputs(602) <= not (a and b);
    layer2_outputs(603) <= a or b;
    layer2_outputs(604) <= not (a or b);
    layer2_outputs(605) <= a and b;
    layer2_outputs(606) <= not b or a;
    layer2_outputs(607) <= b and not a;
    layer2_outputs(608) <= a or b;
    layer2_outputs(609) <= 1'b1;
    layer2_outputs(610) <= a;
    layer2_outputs(611) <= not b;
    layer2_outputs(612) <= not b;
    layer2_outputs(613) <= 1'b1;
    layer2_outputs(614) <= not (a or b);
    layer2_outputs(615) <= 1'b0;
    layer2_outputs(616) <= not b or a;
    layer2_outputs(617) <= b and not a;
    layer2_outputs(618) <= a and b;
    layer2_outputs(619) <= b;
    layer2_outputs(620) <= 1'b1;
    layer2_outputs(621) <= a or b;
    layer2_outputs(622) <= 1'b1;
    layer2_outputs(623) <= a or b;
    layer2_outputs(624) <= not b or a;
    layer2_outputs(625) <= 1'b1;
    layer2_outputs(626) <= not b;
    layer2_outputs(627) <= a;
    layer2_outputs(628) <= not (a xor b);
    layer2_outputs(629) <= 1'b1;
    layer2_outputs(630) <= not b or a;
    layer2_outputs(631) <= 1'b1;
    layer2_outputs(632) <= not a;
    layer2_outputs(633) <= a and not b;
    layer2_outputs(634) <= not a;
    layer2_outputs(635) <= a;
    layer2_outputs(636) <= 1'b0;
    layer2_outputs(637) <= 1'b1;
    layer2_outputs(638) <= a;
    layer2_outputs(639) <= 1'b1;
    layer2_outputs(640) <= not (a or b);
    layer2_outputs(641) <= 1'b0;
    layer2_outputs(642) <= not (a or b);
    layer2_outputs(643) <= not b or a;
    layer2_outputs(644) <= 1'b1;
    layer2_outputs(645) <= not a;
    layer2_outputs(646) <= not (a or b);
    layer2_outputs(647) <= 1'b1;
    layer2_outputs(648) <= not (a or b);
    layer2_outputs(649) <= b;
    layer2_outputs(650) <= b and not a;
    layer2_outputs(651) <= not a or b;
    layer2_outputs(652) <= not a;
    layer2_outputs(653) <= a xor b;
    layer2_outputs(654) <= a and b;
    layer2_outputs(655) <= not (a and b);
    layer2_outputs(656) <= not b or a;
    layer2_outputs(657) <= not a;
    layer2_outputs(658) <= 1'b0;
    layer2_outputs(659) <= 1'b0;
    layer2_outputs(660) <= 1'b0;
    layer2_outputs(661) <= not (a and b);
    layer2_outputs(662) <= not a or b;
    layer2_outputs(663) <= a and not b;
    layer2_outputs(664) <= not b;
    layer2_outputs(665) <= not (a or b);
    layer2_outputs(666) <= b and not a;
    layer2_outputs(667) <= a and b;
    layer2_outputs(668) <= b and not a;
    layer2_outputs(669) <= 1'b1;
    layer2_outputs(670) <= b;
    layer2_outputs(671) <= b;
    layer2_outputs(672) <= not b or a;
    layer2_outputs(673) <= a and b;
    layer2_outputs(674) <= not (a or b);
    layer2_outputs(675) <= a and b;
    layer2_outputs(676) <= a and not b;
    layer2_outputs(677) <= not b or a;
    layer2_outputs(678) <= 1'b0;
    layer2_outputs(679) <= not b;
    layer2_outputs(680) <= not (a and b);
    layer2_outputs(681) <= not (a and b);
    layer2_outputs(682) <= not a;
    layer2_outputs(683) <= 1'b0;
    layer2_outputs(684) <= 1'b0;
    layer2_outputs(685) <= not b;
    layer2_outputs(686) <= not b;
    layer2_outputs(687) <= not (a or b);
    layer2_outputs(688) <= a and not b;
    layer2_outputs(689) <= a and not b;
    layer2_outputs(690) <= a and not b;
    layer2_outputs(691) <= b;
    layer2_outputs(692) <= not (a or b);
    layer2_outputs(693) <= a and not b;
    layer2_outputs(694) <= 1'b1;
    layer2_outputs(695) <= a or b;
    layer2_outputs(696) <= 1'b1;
    layer2_outputs(697) <= not (a xor b);
    layer2_outputs(698) <= a and not b;
    layer2_outputs(699) <= b and not a;
    layer2_outputs(700) <= a or b;
    layer2_outputs(701) <= 1'b1;
    layer2_outputs(702) <= not a;
    layer2_outputs(703) <= not (a xor b);
    layer2_outputs(704) <= b;
    layer2_outputs(705) <= a or b;
    layer2_outputs(706) <= a and b;
    layer2_outputs(707) <= a or b;
    layer2_outputs(708) <= a;
    layer2_outputs(709) <= a and b;
    layer2_outputs(710) <= a or b;
    layer2_outputs(711) <= not a or b;
    layer2_outputs(712) <= a and not b;
    layer2_outputs(713) <= 1'b0;
    layer2_outputs(714) <= 1'b1;
    layer2_outputs(715) <= a and b;
    layer2_outputs(716) <= b;
    layer2_outputs(717) <= 1'b1;
    layer2_outputs(718) <= a and b;
    layer2_outputs(719) <= a;
    layer2_outputs(720) <= not a or b;
    layer2_outputs(721) <= not (a or b);
    layer2_outputs(722) <= not (a and b);
    layer2_outputs(723) <= not (a xor b);
    layer2_outputs(724) <= 1'b0;
    layer2_outputs(725) <= not (a xor b);
    layer2_outputs(726) <= a and not b;
    layer2_outputs(727) <= not (a and b);
    layer2_outputs(728) <= not b;
    layer2_outputs(729) <= not (a or b);
    layer2_outputs(730) <= 1'b0;
    layer2_outputs(731) <= not (a and b);
    layer2_outputs(732) <= not (a or b);
    layer2_outputs(733) <= not a;
    layer2_outputs(734) <= not b;
    layer2_outputs(735) <= not b;
    layer2_outputs(736) <= a;
    layer2_outputs(737) <= b;
    layer2_outputs(738) <= not a or b;
    layer2_outputs(739) <= a and not b;
    layer2_outputs(740) <= not (a or b);
    layer2_outputs(741) <= a and b;
    layer2_outputs(742) <= not b;
    layer2_outputs(743) <= 1'b1;
    layer2_outputs(744) <= not a or b;
    layer2_outputs(745) <= a and not b;
    layer2_outputs(746) <= a or b;
    layer2_outputs(747) <= not (a xor b);
    layer2_outputs(748) <= 1'b0;
    layer2_outputs(749) <= not b or a;
    layer2_outputs(750) <= a;
    layer2_outputs(751) <= a and b;
    layer2_outputs(752) <= b and not a;
    layer2_outputs(753) <= not (a or b);
    layer2_outputs(754) <= not b;
    layer2_outputs(755) <= not b or a;
    layer2_outputs(756) <= 1'b1;
    layer2_outputs(757) <= not b or a;
    layer2_outputs(758) <= b;
    layer2_outputs(759) <= a or b;
    layer2_outputs(760) <= 1'b0;
    layer2_outputs(761) <= a and b;
    layer2_outputs(762) <= 1'b1;
    layer2_outputs(763) <= not b;
    layer2_outputs(764) <= 1'b1;
    layer2_outputs(765) <= b;
    layer2_outputs(766) <= 1'b1;
    layer2_outputs(767) <= not (a and b);
    layer2_outputs(768) <= a and b;
    layer2_outputs(769) <= not a;
    layer2_outputs(770) <= not (a or b);
    layer2_outputs(771) <= 1'b0;
    layer2_outputs(772) <= b and not a;
    layer2_outputs(773) <= not a or b;
    layer2_outputs(774) <= not (a xor b);
    layer2_outputs(775) <= 1'b1;
    layer2_outputs(776) <= a;
    layer2_outputs(777) <= not b;
    layer2_outputs(778) <= not a or b;
    layer2_outputs(779) <= a and b;
    layer2_outputs(780) <= b;
    layer2_outputs(781) <= 1'b0;
    layer2_outputs(782) <= 1'b1;
    layer2_outputs(783) <= 1'b1;
    layer2_outputs(784) <= not b;
    layer2_outputs(785) <= a or b;
    layer2_outputs(786) <= not (a and b);
    layer2_outputs(787) <= b and not a;
    layer2_outputs(788) <= not a;
    layer2_outputs(789) <= a and b;
    layer2_outputs(790) <= not b or a;
    layer2_outputs(791) <= a and b;
    layer2_outputs(792) <= a or b;
    layer2_outputs(793) <= a and b;
    layer2_outputs(794) <= 1'b0;
    layer2_outputs(795) <= 1'b1;
    layer2_outputs(796) <= b and not a;
    layer2_outputs(797) <= not a or b;
    layer2_outputs(798) <= a or b;
    layer2_outputs(799) <= a or b;
    layer2_outputs(800) <= b;
    layer2_outputs(801) <= a and not b;
    layer2_outputs(802) <= 1'b0;
    layer2_outputs(803) <= not (a or b);
    layer2_outputs(804) <= not (a and b);
    layer2_outputs(805) <= not (a or b);
    layer2_outputs(806) <= not b;
    layer2_outputs(807) <= b;
    layer2_outputs(808) <= b and not a;
    layer2_outputs(809) <= 1'b0;
    layer2_outputs(810) <= not (a or b);
    layer2_outputs(811) <= 1'b1;
    layer2_outputs(812) <= a xor b;
    layer2_outputs(813) <= not (a or b);
    layer2_outputs(814) <= not a or b;
    layer2_outputs(815) <= not b;
    layer2_outputs(816) <= not b or a;
    layer2_outputs(817) <= a xor b;
    layer2_outputs(818) <= a and b;
    layer2_outputs(819) <= 1'b1;
    layer2_outputs(820) <= not a or b;
    layer2_outputs(821) <= not a;
    layer2_outputs(822) <= not (a and b);
    layer2_outputs(823) <= 1'b0;
    layer2_outputs(824) <= b;
    layer2_outputs(825) <= a or b;
    layer2_outputs(826) <= b;
    layer2_outputs(827) <= not a or b;
    layer2_outputs(828) <= b and not a;
    layer2_outputs(829) <= a and b;
    layer2_outputs(830) <= not a;
    layer2_outputs(831) <= a or b;
    layer2_outputs(832) <= not (a xor b);
    layer2_outputs(833) <= b;
    layer2_outputs(834) <= not a or b;
    layer2_outputs(835) <= b;
    layer2_outputs(836) <= not b;
    layer2_outputs(837) <= not (a or b);
    layer2_outputs(838) <= not b or a;
    layer2_outputs(839) <= 1'b0;
    layer2_outputs(840) <= 1'b0;
    layer2_outputs(841) <= not (a and b);
    layer2_outputs(842) <= a and b;
    layer2_outputs(843) <= 1'b0;
    layer2_outputs(844) <= not a or b;
    layer2_outputs(845) <= 1'b1;
    layer2_outputs(846) <= a and not b;
    layer2_outputs(847) <= not b or a;
    layer2_outputs(848) <= b and not a;
    layer2_outputs(849) <= a;
    layer2_outputs(850) <= 1'b0;
    layer2_outputs(851) <= not a;
    layer2_outputs(852) <= not (a xor b);
    layer2_outputs(853) <= 1'b0;
    layer2_outputs(854) <= 1'b1;
    layer2_outputs(855) <= 1'b1;
    layer2_outputs(856) <= a and not b;
    layer2_outputs(857) <= a and not b;
    layer2_outputs(858) <= a xor b;
    layer2_outputs(859) <= 1'b1;
    layer2_outputs(860) <= a;
    layer2_outputs(861) <= b and not a;
    layer2_outputs(862) <= not b or a;
    layer2_outputs(863) <= not a;
    layer2_outputs(864) <= a;
    layer2_outputs(865) <= a and b;
    layer2_outputs(866) <= not b or a;
    layer2_outputs(867) <= b and not a;
    layer2_outputs(868) <= a;
    layer2_outputs(869) <= a and b;
    layer2_outputs(870) <= 1'b0;
    layer2_outputs(871) <= not (a and b);
    layer2_outputs(872) <= a and not b;
    layer2_outputs(873) <= 1'b1;
    layer2_outputs(874) <= a and b;
    layer2_outputs(875) <= not (a or b);
    layer2_outputs(876) <= not b;
    layer2_outputs(877) <= not a or b;
    layer2_outputs(878) <= not (a and b);
    layer2_outputs(879) <= a and not b;
    layer2_outputs(880) <= 1'b1;
    layer2_outputs(881) <= a and not b;
    layer2_outputs(882) <= a and b;
    layer2_outputs(883) <= not (a or b);
    layer2_outputs(884) <= 1'b0;
    layer2_outputs(885) <= a;
    layer2_outputs(886) <= not a;
    layer2_outputs(887) <= 1'b0;
    layer2_outputs(888) <= 1'b1;
    layer2_outputs(889) <= not (a and b);
    layer2_outputs(890) <= a or b;
    layer2_outputs(891) <= 1'b1;
    layer2_outputs(892) <= not b or a;
    layer2_outputs(893) <= a and b;
    layer2_outputs(894) <= not (a or b);
    layer2_outputs(895) <= not a or b;
    layer2_outputs(896) <= a or b;
    layer2_outputs(897) <= not a;
    layer2_outputs(898) <= not a or b;
    layer2_outputs(899) <= not (a and b);
    layer2_outputs(900) <= a;
    layer2_outputs(901) <= not (a and b);
    layer2_outputs(902) <= not b or a;
    layer2_outputs(903) <= a or b;
    layer2_outputs(904) <= a;
    layer2_outputs(905) <= 1'b0;
    layer2_outputs(906) <= 1'b1;
    layer2_outputs(907) <= not (a and b);
    layer2_outputs(908) <= b;
    layer2_outputs(909) <= a or b;
    layer2_outputs(910) <= not (a or b);
    layer2_outputs(911) <= not b;
    layer2_outputs(912) <= b;
    layer2_outputs(913) <= a and not b;
    layer2_outputs(914) <= b and not a;
    layer2_outputs(915) <= not (a xor b);
    layer2_outputs(916) <= 1'b1;
    layer2_outputs(917) <= not b or a;
    layer2_outputs(918) <= b;
    layer2_outputs(919) <= not (a and b);
    layer2_outputs(920) <= a or b;
    layer2_outputs(921) <= 1'b0;
    layer2_outputs(922) <= not a;
    layer2_outputs(923) <= b;
    layer2_outputs(924) <= not (a or b);
    layer2_outputs(925) <= not b or a;
    layer2_outputs(926) <= b and not a;
    layer2_outputs(927) <= not (a and b);
    layer2_outputs(928) <= a and not b;
    layer2_outputs(929) <= 1'b0;
    layer2_outputs(930) <= a and not b;
    layer2_outputs(931) <= b and not a;
    layer2_outputs(932) <= not (a and b);
    layer2_outputs(933) <= not b or a;
    layer2_outputs(934) <= 1'b0;
    layer2_outputs(935) <= a and not b;
    layer2_outputs(936) <= a and not b;
    layer2_outputs(937) <= not (a and b);
    layer2_outputs(938) <= a;
    layer2_outputs(939) <= not a;
    layer2_outputs(940) <= not b or a;
    layer2_outputs(941) <= not b;
    layer2_outputs(942) <= b;
    layer2_outputs(943) <= not (a and b);
    layer2_outputs(944) <= not b or a;
    layer2_outputs(945) <= a and not b;
    layer2_outputs(946) <= not (a and b);
    layer2_outputs(947) <= 1'b1;
    layer2_outputs(948) <= not b;
    layer2_outputs(949) <= not a;
    layer2_outputs(950) <= b and not a;
    layer2_outputs(951) <= not b;
    layer2_outputs(952) <= b and not a;
    layer2_outputs(953) <= a;
    layer2_outputs(954) <= a or b;
    layer2_outputs(955) <= a or b;
    layer2_outputs(956) <= a and not b;
    layer2_outputs(957) <= 1'b1;
    layer2_outputs(958) <= a and b;
    layer2_outputs(959) <= not (a or b);
    layer2_outputs(960) <= a and not b;
    layer2_outputs(961) <= not b or a;
    layer2_outputs(962) <= not b or a;
    layer2_outputs(963) <= a or b;
    layer2_outputs(964) <= 1'b0;
    layer2_outputs(965) <= not b;
    layer2_outputs(966) <= not (a and b);
    layer2_outputs(967) <= b and not a;
    layer2_outputs(968) <= not a;
    layer2_outputs(969) <= a xor b;
    layer2_outputs(970) <= not b;
    layer2_outputs(971) <= a and not b;
    layer2_outputs(972) <= not b or a;
    layer2_outputs(973) <= b and not a;
    layer2_outputs(974) <= 1'b0;
    layer2_outputs(975) <= 1'b0;
    layer2_outputs(976) <= a or b;
    layer2_outputs(977) <= a or b;
    layer2_outputs(978) <= b;
    layer2_outputs(979) <= not (a or b);
    layer2_outputs(980) <= a and b;
    layer2_outputs(981) <= not (a and b);
    layer2_outputs(982) <= a or b;
    layer2_outputs(983) <= not (a or b);
    layer2_outputs(984) <= not a or b;
    layer2_outputs(985) <= not (a or b);
    layer2_outputs(986) <= not b;
    layer2_outputs(987) <= a;
    layer2_outputs(988) <= 1'b0;
    layer2_outputs(989) <= 1'b0;
    layer2_outputs(990) <= a and b;
    layer2_outputs(991) <= not (a and b);
    layer2_outputs(992) <= 1'b1;
    layer2_outputs(993) <= not (a xor b);
    layer2_outputs(994) <= not (a or b);
    layer2_outputs(995) <= 1'b0;
    layer2_outputs(996) <= not (a or b);
    layer2_outputs(997) <= a;
    layer2_outputs(998) <= 1'b0;
    layer2_outputs(999) <= 1'b0;
    layer2_outputs(1000) <= b;
    layer2_outputs(1001) <= b;
    layer2_outputs(1002) <= 1'b0;
    layer2_outputs(1003) <= not a;
    layer2_outputs(1004) <= a and not b;
    layer2_outputs(1005) <= not (a and b);
    layer2_outputs(1006) <= not (a or b);
    layer2_outputs(1007) <= b;
    layer2_outputs(1008) <= not a;
    layer2_outputs(1009) <= a and b;
    layer2_outputs(1010) <= not a;
    layer2_outputs(1011) <= a and b;
    layer2_outputs(1012) <= not (a and b);
    layer2_outputs(1013) <= not a or b;
    layer2_outputs(1014) <= not a or b;
    layer2_outputs(1015) <= not a;
    layer2_outputs(1016) <= not (a or b);
    layer2_outputs(1017) <= 1'b1;
    layer2_outputs(1018) <= not b or a;
    layer2_outputs(1019) <= not b or a;
    layer2_outputs(1020) <= a and not b;
    layer2_outputs(1021) <= 1'b1;
    layer2_outputs(1022) <= b and not a;
    layer2_outputs(1023) <= 1'b1;
    layer2_outputs(1024) <= b and not a;
    layer2_outputs(1025) <= a and b;
    layer2_outputs(1026) <= a and not b;
    layer2_outputs(1027) <= a or b;
    layer2_outputs(1028) <= a;
    layer2_outputs(1029) <= a and b;
    layer2_outputs(1030) <= a and b;
    layer2_outputs(1031) <= not (a or b);
    layer2_outputs(1032) <= a;
    layer2_outputs(1033) <= a and b;
    layer2_outputs(1034) <= a or b;
    layer2_outputs(1035) <= not a;
    layer2_outputs(1036) <= b and not a;
    layer2_outputs(1037) <= 1'b0;
    layer2_outputs(1038) <= a and b;
    layer2_outputs(1039) <= not a or b;
    layer2_outputs(1040) <= not (a or b);
    layer2_outputs(1041) <= not (a or b);
    layer2_outputs(1042) <= not b or a;
    layer2_outputs(1043) <= 1'b0;
    layer2_outputs(1044) <= a and b;
    layer2_outputs(1045) <= a;
    layer2_outputs(1046) <= not a or b;
    layer2_outputs(1047) <= 1'b1;
    layer2_outputs(1048) <= a;
    layer2_outputs(1049) <= 1'b0;
    layer2_outputs(1050) <= 1'b1;
    layer2_outputs(1051) <= b;
    layer2_outputs(1052) <= a and b;
    layer2_outputs(1053) <= b and not a;
    layer2_outputs(1054) <= not a or b;
    layer2_outputs(1055) <= not (a xor b);
    layer2_outputs(1056) <= a;
    layer2_outputs(1057) <= not (a and b);
    layer2_outputs(1058) <= not b;
    layer2_outputs(1059) <= b;
    layer2_outputs(1060) <= 1'b0;
    layer2_outputs(1061) <= not (a and b);
    layer2_outputs(1062) <= 1'b1;
    layer2_outputs(1063) <= not b or a;
    layer2_outputs(1064) <= 1'b0;
    layer2_outputs(1065) <= b and not a;
    layer2_outputs(1066) <= a;
    layer2_outputs(1067) <= 1'b0;
    layer2_outputs(1068) <= a and not b;
    layer2_outputs(1069) <= a and b;
    layer2_outputs(1070) <= not (a and b);
    layer2_outputs(1071) <= not b or a;
    layer2_outputs(1072) <= not (a xor b);
    layer2_outputs(1073) <= not a;
    layer2_outputs(1074) <= a or b;
    layer2_outputs(1075) <= 1'b1;
    layer2_outputs(1076) <= not b;
    layer2_outputs(1077) <= a or b;
    layer2_outputs(1078) <= a xor b;
    layer2_outputs(1079) <= a;
    layer2_outputs(1080) <= 1'b0;
    layer2_outputs(1081) <= not (a or b);
    layer2_outputs(1082) <= a and not b;
    layer2_outputs(1083) <= not b or a;
    layer2_outputs(1084) <= not b or a;
    layer2_outputs(1085) <= a;
    layer2_outputs(1086) <= 1'b1;
    layer2_outputs(1087) <= 1'b0;
    layer2_outputs(1088) <= a;
    layer2_outputs(1089) <= not (a xor b);
    layer2_outputs(1090) <= a or b;
    layer2_outputs(1091) <= b;
    layer2_outputs(1092) <= a and not b;
    layer2_outputs(1093) <= 1'b0;
    layer2_outputs(1094) <= a;
    layer2_outputs(1095) <= b;
    layer2_outputs(1096) <= 1'b0;
    layer2_outputs(1097) <= a xor b;
    layer2_outputs(1098) <= a and b;
    layer2_outputs(1099) <= a;
    layer2_outputs(1100) <= a or b;
    layer2_outputs(1101) <= 1'b1;
    layer2_outputs(1102) <= not a;
    layer2_outputs(1103) <= a;
    layer2_outputs(1104) <= b and not a;
    layer2_outputs(1105) <= 1'b0;
    layer2_outputs(1106) <= not a or b;
    layer2_outputs(1107) <= a;
    layer2_outputs(1108) <= not (a and b);
    layer2_outputs(1109) <= a and b;
    layer2_outputs(1110) <= not a;
    layer2_outputs(1111) <= b and not a;
    layer2_outputs(1112) <= not a or b;
    layer2_outputs(1113) <= not (a or b);
    layer2_outputs(1114) <= a xor b;
    layer2_outputs(1115) <= not b or a;
    layer2_outputs(1116) <= a;
    layer2_outputs(1117) <= a or b;
    layer2_outputs(1118) <= a and not b;
    layer2_outputs(1119) <= not b or a;
    layer2_outputs(1120) <= 1'b0;
    layer2_outputs(1121) <= a;
    layer2_outputs(1122) <= 1'b1;
    layer2_outputs(1123) <= a and not b;
    layer2_outputs(1124) <= a or b;
    layer2_outputs(1125) <= not a;
    layer2_outputs(1126) <= 1'b1;
    layer2_outputs(1127) <= b;
    layer2_outputs(1128) <= b;
    layer2_outputs(1129) <= not (a and b);
    layer2_outputs(1130) <= not a or b;
    layer2_outputs(1131) <= not (a or b);
    layer2_outputs(1132) <= not a or b;
    layer2_outputs(1133) <= not a or b;
    layer2_outputs(1134) <= not b or a;
    layer2_outputs(1135) <= a and not b;
    layer2_outputs(1136) <= 1'b1;
    layer2_outputs(1137) <= not b;
    layer2_outputs(1138) <= not (a and b);
    layer2_outputs(1139) <= not b or a;
    layer2_outputs(1140) <= b;
    layer2_outputs(1141) <= a;
    layer2_outputs(1142) <= b and not a;
    layer2_outputs(1143) <= not b;
    layer2_outputs(1144) <= a and not b;
    layer2_outputs(1145) <= not a;
    layer2_outputs(1146) <= 1'b0;
    layer2_outputs(1147) <= 1'b1;
    layer2_outputs(1148) <= not a or b;
    layer2_outputs(1149) <= a and b;
    layer2_outputs(1150) <= a and not b;
    layer2_outputs(1151) <= b and not a;
    layer2_outputs(1152) <= b and not a;
    layer2_outputs(1153) <= b;
    layer2_outputs(1154) <= 1'b1;
    layer2_outputs(1155) <= 1'b0;
    layer2_outputs(1156) <= 1'b0;
    layer2_outputs(1157) <= a;
    layer2_outputs(1158) <= not (a or b);
    layer2_outputs(1159) <= not (a or b);
    layer2_outputs(1160) <= a or b;
    layer2_outputs(1161) <= b;
    layer2_outputs(1162) <= not a or b;
    layer2_outputs(1163) <= 1'b0;
    layer2_outputs(1164) <= not a;
    layer2_outputs(1165) <= a and b;
    layer2_outputs(1166) <= b and not a;
    layer2_outputs(1167) <= not b;
    layer2_outputs(1168) <= 1'b1;
    layer2_outputs(1169) <= not a or b;
    layer2_outputs(1170) <= b;
    layer2_outputs(1171) <= not b;
    layer2_outputs(1172) <= not (a or b);
    layer2_outputs(1173) <= a and b;
    layer2_outputs(1174) <= a and b;
    layer2_outputs(1175) <= 1'b0;
    layer2_outputs(1176) <= not (a and b);
    layer2_outputs(1177) <= a or b;
    layer2_outputs(1178) <= 1'b0;
    layer2_outputs(1179) <= a or b;
    layer2_outputs(1180) <= b;
    layer2_outputs(1181) <= not (a or b);
    layer2_outputs(1182) <= a and b;
    layer2_outputs(1183) <= 1'b0;
    layer2_outputs(1184) <= 1'b1;
    layer2_outputs(1185) <= a;
    layer2_outputs(1186) <= a and b;
    layer2_outputs(1187) <= not b;
    layer2_outputs(1188) <= 1'b0;
    layer2_outputs(1189) <= not b;
    layer2_outputs(1190) <= b and not a;
    layer2_outputs(1191) <= b and not a;
    layer2_outputs(1192) <= 1'b1;
    layer2_outputs(1193) <= a and not b;
    layer2_outputs(1194) <= a or b;
    layer2_outputs(1195) <= 1'b0;
    layer2_outputs(1196) <= b;
    layer2_outputs(1197) <= a and b;
    layer2_outputs(1198) <= a;
    layer2_outputs(1199) <= a;
    layer2_outputs(1200) <= b and not a;
    layer2_outputs(1201) <= not a;
    layer2_outputs(1202) <= not a or b;
    layer2_outputs(1203) <= a and not b;
    layer2_outputs(1204) <= not a;
    layer2_outputs(1205) <= not a;
    layer2_outputs(1206) <= 1'b1;
    layer2_outputs(1207) <= a or b;
    layer2_outputs(1208) <= b and not a;
    layer2_outputs(1209) <= not (a or b);
    layer2_outputs(1210) <= b;
    layer2_outputs(1211) <= a and b;
    layer2_outputs(1212) <= a;
    layer2_outputs(1213) <= b and not a;
    layer2_outputs(1214) <= a or b;
    layer2_outputs(1215) <= not b or a;
    layer2_outputs(1216) <= a and not b;
    layer2_outputs(1217) <= not b;
    layer2_outputs(1218) <= b and not a;
    layer2_outputs(1219) <= b;
    layer2_outputs(1220) <= not b or a;
    layer2_outputs(1221) <= a;
    layer2_outputs(1222) <= b and not a;
    layer2_outputs(1223) <= a xor b;
    layer2_outputs(1224) <= not (a xor b);
    layer2_outputs(1225) <= b and not a;
    layer2_outputs(1226) <= a and b;
    layer2_outputs(1227) <= not b or a;
    layer2_outputs(1228) <= not a or b;
    layer2_outputs(1229) <= not a;
    layer2_outputs(1230) <= not a;
    layer2_outputs(1231) <= not a;
    layer2_outputs(1232) <= b and not a;
    layer2_outputs(1233) <= a or b;
    layer2_outputs(1234) <= not a or b;
    layer2_outputs(1235) <= not a;
    layer2_outputs(1236) <= 1'b0;
    layer2_outputs(1237) <= a;
    layer2_outputs(1238) <= not b or a;
    layer2_outputs(1239) <= 1'b1;
    layer2_outputs(1240) <= not a or b;
    layer2_outputs(1241) <= not b or a;
    layer2_outputs(1242) <= not b;
    layer2_outputs(1243) <= b;
    layer2_outputs(1244) <= not (a or b);
    layer2_outputs(1245) <= 1'b0;
    layer2_outputs(1246) <= 1'b1;
    layer2_outputs(1247) <= not a or b;
    layer2_outputs(1248) <= a and b;
    layer2_outputs(1249) <= 1'b0;
    layer2_outputs(1250) <= a;
    layer2_outputs(1251) <= not (a and b);
    layer2_outputs(1252) <= not a or b;
    layer2_outputs(1253) <= a xor b;
    layer2_outputs(1254) <= not b or a;
    layer2_outputs(1255) <= not a or b;
    layer2_outputs(1256) <= not (a and b);
    layer2_outputs(1257) <= 1'b0;
    layer2_outputs(1258) <= not (a or b);
    layer2_outputs(1259) <= 1'b1;
    layer2_outputs(1260) <= 1'b1;
    layer2_outputs(1261) <= b and not a;
    layer2_outputs(1262) <= not (a or b);
    layer2_outputs(1263) <= 1'b0;
    layer2_outputs(1264) <= 1'b0;
    layer2_outputs(1265) <= not (a xor b);
    layer2_outputs(1266) <= not a or b;
    layer2_outputs(1267) <= 1'b0;
    layer2_outputs(1268) <= a;
    layer2_outputs(1269) <= b and not a;
    layer2_outputs(1270) <= not b or a;
    layer2_outputs(1271) <= not b;
    layer2_outputs(1272) <= a and b;
    layer2_outputs(1273) <= not a;
    layer2_outputs(1274) <= not a;
    layer2_outputs(1275) <= not (a and b);
    layer2_outputs(1276) <= 1'b1;
    layer2_outputs(1277) <= a;
    layer2_outputs(1278) <= not b;
    layer2_outputs(1279) <= not b;
    layer2_outputs(1280) <= b;
    layer2_outputs(1281) <= not b;
    layer2_outputs(1282) <= 1'b1;
    layer2_outputs(1283) <= b;
    layer2_outputs(1284) <= a;
    layer2_outputs(1285) <= a or b;
    layer2_outputs(1286) <= a;
    layer2_outputs(1287) <= b and not a;
    layer2_outputs(1288) <= not a;
    layer2_outputs(1289) <= a or b;
    layer2_outputs(1290) <= not (a or b);
    layer2_outputs(1291) <= a and not b;
    layer2_outputs(1292) <= 1'b0;
    layer2_outputs(1293) <= a and not b;
    layer2_outputs(1294) <= not (a and b);
    layer2_outputs(1295) <= not b or a;
    layer2_outputs(1296) <= 1'b1;
    layer2_outputs(1297) <= 1'b0;
    layer2_outputs(1298) <= not a or b;
    layer2_outputs(1299) <= not b or a;
    layer2_outputs(1300) <= not a;
    layer2_outputs(1301) <= 1'b0;
    layer2_outputs(1302) <= not (a and b);
    layer2_outputs(1303) <= 1'b1;
    layer2_outputs(1304) <= 1'b0;
    layer2_outputs(1305) <= not (a xor b);
    layer2_outputs(1306) <= a;
    layer2_outputs(1307) <= a xor b;
    layer2_outputs(1308) <= a xor b;
    layer2_outputs(1309) <= a;
    layer2_outputs(1310) <= 1'b0;
    layer2_outputs(1311) <= 1'b1;
    layer2_outputs(1312) <= 1'b1;
    layer2_outputs(1313) <= b;
    layer2_outputs(1314) <= b;
    layer2_outputs(1315) <= not a or b;
    layer2_outputs(1316) <= not a;
    layer2_outputs(1317) <= not a;
    layer2_outputs(1318) <= b and not a;
    layer2_outputs(1319) <= a and b;
    layer2_outputs(1320) <= 1'b0;
    layer2_outputs(1321) <= not a;
    layer2_outputs(1322) <= a and not b;
    layer2_outputs(1323) <= b and not a;
    layer2_outputs(1324) <= b and not a;
    layer2_outputs(1325) <= not a;
    layer2_outputs(1326) <= 1'b1;
    layer2_outputs(1327) <= a or b;
    layer2_outputs(1328) <= b and not a;
    layer2_outputs(1329) <= not a or b;
    layer2_outputs(1330) <= a and b;
    layer2_outputs(1331) <= b and not a;
    layer2_outputs(1332) <= 1'b1;
    layer2_outputs(1333) <= b;
    layer2_outputs(1334) <= not b;
    layer2_outputs(1335) <= not a;
    layer2_outputs(1336) <= a and not b;
    layer2_outputs(1337) <= a and not b;
    layer2_outputs(1338) <= a;
    layer2_outputs(1339) <= a or b;
    layer2_outputs(1340) <= not a or b;
    layer2_outputs(1341) <= 1'b1;
    layer2_outputs(1342) <= 1'b0;
    layer2_outputs(1343) <= 1'b0;
    layer2_outputs(1344) <= 1'b0;
    layer2_outputs(1345) <= a xor b;
    layer2_outputs(1346) <= not b or a;
    layer2_outputs(1347) <= a;
    layer2_outputs(1348) <= 1'b1;
    layer2_outputs(1349) <= 1'b0;
    layer2_outputs(1350) <= a and not b;
    layer2_outputs(1351) <= a or b;
    layer2_outputs(1352) <= 1'b1;
    layer2_outputs(1353) <= a and not b;
    layer2_outputs(1354) <= not b;
    layer2_outputs(1355) <= a and b;
    layer2_outputs(1356) <= 1'b0;
    layer2_outputs(1357) <= b and not a;
    layer2_outputs(1358) <= 1'b0;
    layer2_outputs(1359) <= a and b;
    layer2_outputs(1360) <= a;
    layer2_outputs(1361) <= a;
    layer2_outputs(1362) <= 1'b0;
    layer2_outputs(1363) <= a and not b;
    layer2_outputs(1364) <= b;
    layer2_outputs(1365) <= not (a xor b);
    layer2_outputs(1366) <= not b;
    layer2_outputs(1367) <= 1'b0;
    layer2_outputs(1368) <= b;
    layer2_outputs(1369) <= not (a and b);
    layer2_outputs(1370) <= 1'b0;
    layer2_outputs(1371) <= a;
    layer2_outputs(1372) <= a;
    layer2_outputs(1373) <= not (a or b);
    layer2_outputs(1374) <= 1'b1;
    layer2_outputs(1375) <= not (a and b);
    layer2_outputs(1376) <= not b or a;
    layer2_outputs(1377) <= a or b;
    layer2_outputs(1378) <= not (a and b);
    layer2_outputs(1379) <= b;
    layer2_outputs(1380) <= not b or a;
    layer2_outputs(1381) <= not a or b;
    layer2_outputs(1382) <= not (a and b);
    layer2_outputs(1383) <= 1'b1;
    layer2_outputs(1384) <= a or b;
    layer2_outputs(1385) <= not a;
    layer2_outputs(1386) <= a and b;
    layer2_outputs(1387) <= not (a and b);
    layer2_outputs(1388) <= not (a or b);
    layer2_outputs(1389) <= a and b;
    layer2_outputs(1390) <= a;
    layer2_outputs(1391) <= b and not a;
    layer2_outputs(1392) <= b;
    layer2_outputs(1393) <= not b;
    layer2_outputs(1394) <= not b;
    layer2_outputs(1395) <= not a or b;
    layer2_outputs(1396) <= a and not b;
    layer2_outputs(1397) <= not a or b;
    layer2_outputs(1398) <= not (a or b);
    layer2_outputs(1399) <= 1'b0;
    layer2_outputs(1400) <= not (a and b);
    layer2_outputs(1401) <= a and not b;
    layer2_outputs(1402) <= b;
    layer2_outputs(1403) <= 1'b0;
    layer2_outputs(1404) <= not (a and b);
    layer2_outputs(1405) <= a and b;
    layer2_outputs(1406) <= b;
    layer2_outputs(1407) <= b;
    layer2_outputs(1408) <= a;
    layer2_outputs(1409) <= not b;
    layer2_outputs(1410) <= b;
    layer2_outputs(1411) <= not a;
    layer2_outputs(1412) <= a xor b;
    layer2_outputs(1413) <= not b;
    layer2_outputs(1414) <= a;
    layer2_outputs(1415) <= not (a or b);
    layer2_outputs(1416) <= not (a or b);
    layer2_outputs(1417) <= 1'b1;
    layer2_outputs(1418) <= b and not a;
    layer2_outputs(1419) <= not a or b;
    layer2_outputs(1420) <= a and not b;
    layer2_outputs(1421) <= b;
    layer2_outputs(1422) <= not a;
    layer2_outputs(1423) <= a or b;
    layer2_outputs(1424) <= b and not a;
    layer2_outputs(1425) <= a and not b;
    layer2_outputs(1426) <= 1'b1;
    layer2_outputs(1427) <= a and b;
    layer2_outputs(1428) <= not (a and b);
    layer2_outputs(1429) <= 1'b0;
    layer2_outputs(1430) <= not (a and b);
    layer2_outputs(1431) <= not (a or b);
    layer2_outputs(1432) <= a and b;
    layer2_outputs(1433) <= b;
    layer2_outputs(1434) <= not (a and b);
    layer2_outputs(1435) <= not b or a;
    layer2_outputs(1436) <= a or b;
    layer2_outputs(1437) <= 1'b1;
    layer2_outputs(1438) <= a and not b;
    layer2_outputs(1439) <= not a or b;
    layer2_outputs(1440) <= not b or a;
    layer2_outputs(1441) <= a and not b;
    layer2_outputs(1442) <= a or b;
    layer2_outputs(1443) <= not a or b;
    layer2_outputs(1444) <= not a;
    layer2_outputs(1445) <= not (a or b);
    layer2_outputs(1446) <= 1'b0;
    layer2_outputs(1447) <= a or b;
    layer2_outputs(1448) <= not (a or b);
    layer2_outputs(1449) <= not (a and b);
    layer2_outputs(1450) <= 1'b0;
    layer2_outputs(1451) <= b and not a;
    layer2_outputs(1452) <= a and not b;
    layer2_outputs(1453) <= b and not a;
    layer2_outputs(1454) <= not (a and b);
    layer2_outputs(1455) <= a and not b;
    layer2_outputs(1456) <= a and not b;
    layer2_outputs(1457) <= not b or a;
    layer2_outputs(1458) <= a or b;
    layer2_outputs(1459) <= not a or b;
    layer2_outputs(1460) <= not a or b;
    layer2_outputs(1461) <= not (a or b);
    layer2_outputs(1462) <= not (a xor b);
    layer2_outputs(1463) <= not (a and b);
    layer2_outputs(1464) <= not (a or b);
    layer2_outputs(1465) <= b and not a;
    layer2_outputs(1466) <= 1'b1;
    layer2_outputs(1467) <= a and b;
    layer2_outputs(1468) <= not a;
    layer2_outputs(1469) <= not (a or b);
    layer2_outputs(1470) <= 1'b0;
    layer2_outputs(1471) <= 1'b0;
    layer2_outputs(1472) <= a and b;
    layer2_outputs(1473) <= not b;
    layer2_outputs(1474) <= not a;
    layer2_outputs(1475) <= a;
    layer2_outputs(1476) <= 1'b1;
    layer2_outputs(1477) <= b and not a;
    layer2_outputs(1478) <= b;
    layer2_outputs(1479) <= 1'b1;
    layer2_outputs(1480) <= not a;
    layer2_outputs(1481) <= not (a or b);
    layer2_outputs(1482) <= 1'b0;
    layer2_outputs(1483) <= 1'b1;
    layer2_outputs(1484) <= not (a and b);
    layer2_outputs(1485) <= 1'b0;
    layer2_outputs(1486) <= a and not b;
    layer2_outputs(1487) <= not b or a;
    layer2_outputs(1488) <= a;
    layer2_outputs(1489) <= not b or a;
    layer2_outputs(1490) <= b;
    layer2_outputs(1491) <= a and b;
    layer2_outputs(1492) <= not a;
    layer2_outputs(1493) <= b and not a;
    layer2_outputs(1494) <= a;
    layer2_outputs(1495) <= a;
    layer2_outputs(1496) <= a or b;
    layer2_outputs(1497) <= a;
    layer2_outputs(1498) <= a and not b;
    layer2_outputs(1499) <= b and not a;
    layer2_outputs(1500) <= 1'b1;
    layer2_outputs(1501) <= a or b;
    layer2_outputs(1502) <= not a or b;
    layer2_outputs(1503) <= 1'b0;
    layer2_outputs(1504) <= 1'b0;
    layer2_outputs(1505) <= 1'b1;
    layer2_outputs(1506) <= b and not a;
    layer2_outputs(1507) <= a and b;
    layer2_outputs(1508) <= a or b;
    layer2_outputs(1509) <= not (a or b);
    layer2_outputs(1510) <= a and not b;
    layer2_outputs(1511) <= not a or b;
    layer2_outputs(1512) <= a;
    layer2_outputs(1513) <= a and b;
    layer2_outputs(1514) <= 1'b1;
    layer2_outputs(1515) <= a or b;
    layer2_outputs(1516) <= a and not b;
    layer2_outputs(1517) <= not b or a;
    layer2_outputs(1518) <= a and not b;
    layer2_outputs(1519) <= not b;
    layer2_outputs(1520) <= not (a or b);
    layer2_outputs(1521) <= 1'b1;
    layer2_outputs(1522) <= not b or a;
    layer2_outputs(1523) <= b;
    layer2_outputs(1524) <= 1'b1;
    layer2_outputs(1525) <= 1'b1;
    layer2_outputs(1526) <= not a or b;
    layer2_outputs(1527) <= 1'b1;
    layer2_outputs(1528) <= not b or a;
    layer2_outputs(1529) <= b;
    layer2_outputs(1530) <= not a;
    layer2_outputs(1531) <= not (a and b);
    layer2_outputs(1532) <= 1'b1;
    layer2_outputs(1533) <= 1'b0;
    layer2_outputs(1534) <= 1'b0;
    layer2_outputs(1535) <= 1'b0;
    layer2_outputs(1536) <= not a;
    layer2_outputs(1537) <= b;
    layer2_outputs(1538) <= not (a and b);
    layer2_outputs(1539) <= b;
    layer2_outputs(1540) <= a and b;
    layer2_outputs(1541) <= a xor b;
    layer2_outputs(1542) <= not b or a;
    layer2_outputs(1543) <= 1'b0;
    layer2_outputs(1544) <= b and not a;
    layer2_outputs(1545) <= not a or b;
    layer2_outputs(1546) <= a;
    layer2_outputs(1547) <= not (a or b);
    layer2_outputs(1548) <= not b or a;
    layer2_outputs(1549) <= 1'b1;
    layer2_outputs(1550) <= a or b;
    layer2_outputs(1551) <= not (a and b);
    layer2_outputs(1552) <= b;
    layer2_outputs(1553) <= not b;
    layer2_outputs(1554) <= not b;
    layer2_outputs(1555) <= 1'b1;
    layer2_outputs(1556) <= b;
    layer2_outputs(1557) <= not (a and b);
    layer2_outputs(1558) <= not (a and b);
    layer2_outputs(1559) <= b;
    layer2_outputs(1560) <= b and not a;
    layer2_outputs(1561) <= not a or b;
    layer2_outputs(1562) <= not (a and b);
    layer2_outputs(1563) <= a and b;
    layer2_outputs(1564) <= 1'b1;
    layer2_outputs(1565) <= 1'b1;
    layer2_outputs(1566) <= not b;
    layer2_outputs(1567) <= 1'b1;
    layer2_outputs(1568) <= not (a or b);
    layer2_outputs(1569) <= not (a or b);
    layer2_outputs(1570) <= 1'b1;
    layer2_outputs(1571) <= b;
    layer2_outputs(1572) <= 1'b1;
    layer2_outputs(1573) <= a;
    layer2_outputs(1574) <= a and not b;
    layer2_outputs(1575) <= a and not b;
    layer2_outputs(1576) <= b and not a;
    layer2_outputs(1577) <= a and b;
    layer2_outputs(1578) <= not a or b;
    layer2_outputs(1579) <= not (a or b);
    layer2_outputs(1580) <= not (a or b);
    layer2_outputs(1581) <= a or b;
    layer2_outputs(1582) <= not b or a;
    layer2_outputs(1583) <= not (a and b);
    layer2_outputs(1584) <= not a;
    layer2_outputs(1585) <= b and not a;
    layer2_outputs(1586) <= a or b;
    layer2_outputs(1587) <= not b;
    layer2_outputs(1588) <= b and not a;
    layer2_outputs(1589) <= a and b;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= a and not b;
    layer2_outputs(1592) <= b and not a;
    layer2_outputs(1593) <= a and not b;
    layer2_outputs(1594) <= not (a or b);
    layer2_outputs(1595) <= b;
    layer2_outputs(1596) <= b and not a;
    layer2_outputs(1597) <= not a;
    layer2_outputs(1598) <= b and not a;
    layer2_outputs(1599) <= 1'b0;
    layer2_outputs(1600) <= 1'b0;
    layer2_outputs(1601) <= not (a and b);
    layer2_outputs(1602) <= not b;
    layer2_outputs(1603) <= not (a and b);
    layer2_outputs(1604) <= a and not b;
    layer2_outputs(1605) <= 1'b1;
    layer2_outputs(1606) <= not b or a;
    layer2_outputs(1607) <= 1'b1;
    layer2_outputs(1608) <= a;
    layer2_outputs(1609) <= 1'b0;
    layer2_outputs(1610) <= not (a and b);
    layer2_outputs(1611) <= not (a and b);
    layer2_outputs(1612) <= b;
    layer2_outputs(1613) <= a;
    layer2_outputs(1614) <= 1'b0;
    layer2_outputs(1615) <= not a;
    layer2_outputs(1616) <= b;
    layer2_outputs(1617) <= not a or b;
    layer2_outputs(1618) <= not (a or b);
    layer2_outputs(1619) <= b and not a;
    layer2_outputs(1620) <= b;
    layer2_outputs(1621) <= a and b;
    layer2_outputs(1622) <= not a;
    layer2_outputs(1623) <= b and not a;
    layer2_outputs(1624) <= a or b;
    layer2_outputs(1625) <= not (a and b);
    layer2_outputs(1626) <= not (a xor b);
    layer2_outputs(1627) <= not (a or b);
    layer2_outputs(1628) <= a and not b;
    layer2_outputs(1629) <= not b or a;
    layer2_outputs(1630) <= not a;
    layer2_outputs(1631) <= not b or a;
    layer2_outputs(1632) <= not b;
    layer2_outputs(1633) <= a and b;
    layer2_outputs(1634) <= b and not a;
    layer2_outputs(1635) <= b;
    layer2_outputs(1636) <= 1'b1;
    layer2_outputs(1637) <= not b;
    layer2_outputs(1638) <= not (a and b);
    layer2_outputs(1639) <= not b;
    layer2_outputs(1640) <= 1'b0;
    layer2_outputs(1641) <= not (a or b);
    layer2_outputs(1642) <= not b or a;
    layer2_outputs(1643) <= a and not b;
    layer2_outputs(1644) <= a and not b;
    layer2_outputs(1645) <= a and b;
    layer2_outputs(1646) <= b;
    layer2_outputs(1647) <= not b or a;
    layer2_outputs(1648) <= 1'b1;
    layer2_outputs(1649) <= not a or b;
    layer2_outputs(1650) <= not b or a;
    layer2_outputs(1651) <= not a or b;
    layer2_outputs(1652) <= a and b;
    layer2_outputs(1653) <= b and not a;
    layer2_outputs(1654) <= a and b;
    layer2_outputs(1655) <= 1'b0;
    layer2_outputs(1656) <= 1'b1;
    layer2_outputs(1657) <= a or b;
    layer2_outputs(1658) <= a;
    layer2_outputs(1659) <= not a or b;
    layer2_outputs(1660) <= not (a xor b);
    layer2_outputs(1661) <= a or b;
    layer2_outputs(1662) <= b;
    layer2_outputs(1663) <= 1'b0;
    layer2_outputs(1664) <= not b;
    layer2_outputs(1665) <= b;
    layer2_outputs(1666) <= b and not a;
    layer2_outputs(1667) <= a and not b;
    layer2_outputs(1668) <= b;
    layer2_outputs(1669) <= not b or a;
    layer2_outputs(1670) <= a and not b;
    layer2_outputs(1671) <= not a or b;
    layer2_outputs(1672) <= a;
    layer2_outputs(1673) <= a and b;
    layer2_outputs(1674) <= 1'b1;
    layer2_outputs(1675) <= a or b;
    layer2_outputs(1676) <= b and not a;
    layer2_outputs(1677) <= 1'b1;
    layer2_outputs(1678) <= a;
    layer2_outputs(1679) <= a or b;
    layer2_outputs(1680) <= b and not a;
    layer2_outputs(1681) <= a;
    layer2_outputs(1682) <= 1'b0;
    layer2_outputs(1683) <= not (a and b);
    layer2_outputs(1684) <= not (a or b);
    layer2_outputs(1685) <= not b or a;
    layer2_outputs(1686) <= not (a or b);
    layer2_outputs(1687) <= b and not a;
    layer2_outputs(1688) <= b and not a;
    layer2_outputs(1689) <= a and not b;
    layer2_outputs(1690) <= not b;
    layer2_outputs(1691) <= not (a and b);
    layer2_outputs(1692) <= a xor b;
    layer2_outputs(1693) <= not a or b;
    layer2_outputs(1694) <= 1'b1;
    layer2_outputs(1695) <= not (a and b);
    layer2_outputs(1696) <= b and not a;
    layer2_outputs(1697) <= not (a or b);
    layer2_outputs(1698) <= 1'b0;
    layer2_outputs(1699) <= not (a xor b);
    layer2_outputs(1700) <= not b or a;
    layer2_outputs(1701) <= a and not b;
    layer2_outputs(1702) <= a xor b;
    layer2_outputs(1703) <= 1'b0;
    layer2_outputs(1704) <= not b;
    layer2_outputs(1705) <= 1'b0;
    layer2_outputs(1706) <= a;
    layer2_outputs(1707) <= not b;
    layer2_outputs(1708) <= not (a and b);
    layer2_outputs(1709) <= b and not a;
    layer2_outputs(1710) <= 1'b0;
    layer2_outputs(1711) <= not (a or b);
    layer2_outputs(1712) <= 1'b1;
    layer2_outputs(1713) <= not (a or b);
    layer2_outputs(1714) <= not b;
    layer2_outputs(1715) <= not b or a;
    layer2_outputs(1716) <= not a;
    layer2_outputs(1717) <= not (a or b);
    layer2_outputs(1718) <= a xor b;
    layer2_outputs(1719) <= a;
    layer2_outputs(1720) <= a and b;
    layer2_outputs(1721) <= not b;
    layer2_outputs(1722) <= 1'b1;
    layer2_outputs(1723) <= 1'b1;
    layer2_outputs(1724) <= b and not a;
    layer2_outputs(1725) <= b and not a;
    layer2_outputs(1726) <= b;
    layer2_outputs(1727) <= not a or b;
    layer2_outputs(1728) <= 1'b0;
    layer2_outputs(1729) <= b and not a;
    layer2_outputs(1730) <= not (a or b);
    layer2_outputs(1731) <= a and b;
    layer2_outputs(1732) <= not b or a;
    layer2_outputs(1733) <= not a;
    layer2_outputs(1734) <= a and not b;
    layer2_outputs(1735) <= a and b;
    layer2_outputs(1736) <= 1'b1;
    layer2_outputs(1737) <= not (a or b);
    layer2_outputs(1738) <= not a or b;
    layer2_outputs(1739) <= a or b;
    layer2_outputs(1740) <= 1'b0;
    layer2_outputs(1741) <= 1'b0;
    layer2_outputs(1742) <= not a;
    layer2_outputs(1743) <= 1'b0;
    layer2_outputs(1744) <= b;
    layer2_outputs(1745) <= a xor b;
    layer2_outputs(1746) <= not a or b;
    layer2_outputs(1747) <= not (a xor b);
    layer2_outputs(1748) <= a or b;
    layer2_outputs(1749) <= not (a and b);
    layer2_outputs(1750) <= 1'b0;
    layer2_outputs(1751) <= a and not b;
    layer2_outputs(1752) <= b and not a;
    layer2_outputs(1753) <= 1'b1;
    layer2_outputs(1754) <= a and b;
    layer2_outputs(1755) <= a or b;
    layer2_outputs(1756) <= 1'b1;
    layer2_outputs(1757) <= b and not a;
    layer2_outputs(1758) <= not b or a;
    layer2_outputs(1759) <= not a or b;
    layer2_outputs(1760) <= b and not a;
    layer2_outputs(1761) <= a;
    layer2_outputs(1762) <= not (a and b);
    layer2_outputs(1763) <= a xor b;
    layer2_outputs(1764) <= a xor b;
    layer2_outputs(1765) <= not a or b;
    layer2_outputs(1766) <= not b or a;
    layer2_outputs(1767) <= a or b;
    layer2_outputs(1768) <= a or b;
    layer2_outputs(1769) <= not a;
    layer2_outputs(1770) <= b and not a;
    layer2_outputs(1771) <= b and not a;
    layer2_outputs(1772) <= not a;
    layer2_outputs(1773) <= 1'b0;
    layer2_outputs(1774) <= not b;
    layer2_outputs(1775) <= 1'b0;
    layer2_outputs(1776) <= b and not a;
    layer2_outputs(1777) <= not (a xor b);
    layer2_outputs(1778) <= 1'b0;
    layer2_outputs(1779) <= a and b;
    layer2_outputs(1780) <= not b;
    layer2_outputs(1781) <= a xor b;
    layer2_outputs(1782) <= not (a or b);
    layer2_outputs(1783) <= not a;
    layer2_outputs(1784) <= 1'b0;
    layer2_outputs(1785) <= b and not a;
    layer2_outputs(1786) <= not b;
    layer2_outputs(1787) <= not a or b;
    layer2_outputs(1788) <= not b;
    layer2_outputs(1789) <= 1'b1;
    layer2_outputs(1790) <= b and not a;
    layer2_outputs(1791) <= not b;
    layer2_outputs(1792) <= not b or a;
    layer2_outputs(1793) <= not b;
    layer2_outputs(1794) <= not b or a;
    layer2_outputs(1795) <= not (a or b);
    layer2_outputs(1796) <= not (a and b);
    layer2_outputs(1797) <= b;
    layer2_outputs(1798) <= a and not b;
    layer2_outputs(1799) <= b and not a;
    layer2_outputs(1800) <= a or b;
    layer2_outputs(1801) <= a;
    layer2_outputs(1802) <= a and not b;
    layer2_outputs(1803) <= 1'b1;
    layer2_outputs(1804) <= b;
    layer2_outputs(1805) <= a and b;
    layer2_outputs(1806) <= 1'b0;
    layer2_outputs(1807) <= 1'b1;
    layer2_outputs(1808) <= a and not b;
    layer2_outputs(1809) <= not a or b;
    layer2_outputs(1810) <= 1'b0;
    layer2_outputs(1811) <= not (a or b);
    layer2_outputs(1812) <= a;
    layer2_outputs(1813) <= not (a or b);
    layer2_outputs(1814) <= 1'b1;
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= a and not b;
    layer2_outputs(1817) <= not b;
    layer2_outputs(1818) <= a;
    layer2_outputs(1819) <= not a or b;
    layer2_outputs(1820) <= not (a or b);
    layer2_outputs(1821) <= a;
    layer2_outputs(1822) <= not b or a;
    layer2_outputs(1823) <= not b or a;
    layer2_outputs(1824) <= not (a or b);
    layer2_outputs(1825) <= not b;
    layer2_outputs(1826) <= b;
    layer2_outputs(1827) <= a and b;
    layer2_outputs(1828) <= 1'b1;
    layer2_outputs(1829) <= 1'b0;
    layer2_outputs(1830) <= not a;
    layer2_outputs(1831) <= b;
    layer2_outputs(1832) <= a and b;
    layer2_outputs(1833) <= b;
    layer2_outputs(1834) <= not a;
    layer2_outputs(1835) <= not (a or b);
    layer2_outputs(1836) <= not b;
    layer2_outputs(1837) <= a and b;
    layer2_outputs(1838) <= not a;
    layer2_outputs(1839) <= not a;
    layer2_outputs(1840) <= b;
    layer2_outputs(1841) <= not (a or b);
    layer2_outputs(1842) <= not (a xor b);
    layer2_outputs(1843) <= not (a and b);
    layer2_outputs(1844) <= b and not a;
    layer2_outputs(1845) <= not b or a;
    layer2_outputs(1846) <= b;
    layer2_outputs(1847) <= not (a or b);
    layer2_outputs(1848) <= not b;
    layer2_outputs(1849) <= 1'b0;
    layer2_outputs(1850) <= 1'b1;
    layer2_outputs(1851) <= b;
    layer2_outputs(1852) <= not a;
    layer2_outputs(1853) <= b and not a;
    layer2_outputs(1854) <= not a;
    layer2_outputs(1855) <= 1'b0;
    layer2_outputs(1856) <= b;
    layer2_outputs(1857) <= not (a or b);
    layer2_outputs(1858) <= not a;
    layer2_outputs(1859) <= not a;
    layer2_outputs(1860) <= not b or a;
    layer2_outputs(1861) <= not a or b;
    layer2_outputs(1862) <= not a;
    layer2_outputs(1863) <= not b or a;
    layer2_outputs(1864) <= not (a and b);
    layer2_outputs(1865) <= a and b;
    layer2_outputs(1866) <= not b;
    layer2_outputs(1867) <= a and b;
    layer2_outputs(1868) <= not a;
    layer2_outputs(1869) <= not b;
    layer2_outputs(1870) <= not a;
    layer2_outputs(1871) <= a and not b;
    layer2_outputs(1872) <= a and b;
    layer2_outputs(1873) <= not a or b;
    layer2_outputs(1874) <= b and not a;
    layer2_outputs(1875) <= not a or b;
    layer2_outputs(1876) <= a;
    layer2_outputs(1877) <= not (a or b);
    layer2_outputs(1878) <= 1'b0;
    layer2_outputs(1879) <= not (a or b);
    layer2_outputs(1880) <= not b;
    layer2_outputs(1881) <= not (a and b);
    layer2_outputs(1882) <= not a or b;
    layer2_outputs(1883) <= not (a or b);
    layer2_outputs(1884) <= not a or b;
    layer2_outputs(1885) <= a and b;
    layer2_outputs(1886) <= not (a or b);
    layer2_outputs(1887) <= b and not a;
    layer2_outputs(1888) <= not a or b;
    layer2_outputs(1889) <= not a or b;
    layer2_outputs(1890) <= 1'b1;
    layer2_outputs(1891) <= not a;
    layer2_outputs(1892) <= a and b;
    layer2_outputs(1893) <= a and not b;
    layer2_outputs(1894) <= b and not a;
    layer2_outputs(1895) <= not a;
    layer2_outputs(1896) <= a and b;
    layer2_outputs(1897) <= not a or b;
    layer2_outputs(1898) <= a;
    layer2_outputs(1899) <= not (a or b);
    layer2_outputs(1900) <= a and b;
    layer2_outputs(1901) <= a or b;
    layer2_outputs(1902) <= not b;
    layer2_outputs(1903) <= 1'b1;
    layer2_outputs(1904) <= a or b;
    layer2_outputs(1905) <= not b or a;
    layer2_outputs(1906) <= not a;
    layer2_outputs(1907) <= not a or b;
    layer2_outputs(1908) <= b and not a;
    layer2_outputs(1909) <= 1'b0;
    layer2_outputs(1910) <= 1'b1;
    layer2_outputs(1911) <= b and not a;
    layer2_outputs(1912) <= b;
    layer2_outputs(1913) <= b;
    layer2_outputs(1914) <= a and b;
    layer2_outputs(1915) <= a and not b;
    layer2_outputs(1916) <= not b or a;
    layer2_outputs(1917) <= a or b;
    layer2_outputs(1918) <= not b;
    layer2_outputs(1919) <= 1'b1;
    layer2_outputs(1920) <= a and not b;
    layer2_outputs(1921) <= 1'b1;
    layer2_outputs(1922) <= not a or b;
    layer2_outputs(1923) <= not a or b;
    layer2_outputs(1924) <= a and b;
    layer2_outputs(1925) <= 1'b0;
    layer2_outputs(1926) <= not b or a;
    layer2_outputs(1927) <= 1'b0;
    layer2_outputs(1928) <= 1'b1;
    layer2_outputs(1929) <= 1'b0;
    layer2_outputs(1930) <= not a or b;
    layer2_outputs(1931) <= 1'b0;
    layer2_outputs(1932) <= not (a or b);
    layer2_outputs(1933) <= 1'b0;
    layer2_outputs(1934) <= 1'b1;
    layer2_outputs(1935) <= a;
    layer2_outputs(1936) <= not (a and b);
    layer2_outputs(1937) <= b;
    layer2_outputs(1938) <= not (a and b);
    layer2_outputs(1939) <= not b or a;
    layer2_outputs(1940) <= 1'b0;
    layer2_outputs(1941) <= not (a or b);
    layer2_outputs(1942) <= b and not a;
    layer2_outputs(1943) <= not (a or b);
    layer2_outputs(1944) <= a or b;
    layer2_outputs(1945) <= b and not a;
    layer2_outputs(1946) <= 1'b0;
    layer2_outputs(1947) <= not b or a;
    layer2_outputs(1948) <= not b or a;
    layer2_outputs(1949) <= not (a or b);
    layer2_outputs(1950) <= not a;
    layer2_outputs(1951) <= not a or b;
    layer2_outputs(1952) <= 1'b0;
    layer2_outputs(1953) <= a and b;
    layer2_outputs(1954) <= 1'b1;
    layer2_outputs(1955) <= not b;
    layer2_outputs(1956) <= a;
    layer2_outputs(1957) <= not a or b;
    layer2_outputs(1958) <= 1'b1;
    layer2_outputs(1959) <= b and not a;
    layer2_outputs(1960) <= not (a or b);
    layer2_outputs(1961) <= not (a or b);
    layer2_outputs(1962) <= a;
    layer2_outputs(1963) <= a and not b;
    layer2_outputs(1964) <= not (a and b);
    layer2_outputs(1965) <= 1'b1;
    layer2_outputs(1966) <= b and not a;
    layer2_outputs(1967) <= not a;
    layer2_outputs(1968) <= a or b;
    layer2_outputs(1969) <= a and b;
    layer2_outputs(1970) <= 1'b0;
    layer2_outputs(1971) <= 1'b0;
    layer2_outputs(1972) <= a and not b;
    layer2_outputs(1973) <= 1'b0;
    layer2_outputs(1974) <= b;
    layer2_outputs(1975) <= 1'b0;
    layer2_outputs(1976) <= not a;
    layer2_outputs(1977) <= not b or a;
    layer2_outputs(1978) <= not a or b;
    layer2_outputs(1979) <= not (a or b);
    layer2_outputs(1980) <= a and not b;
    layer2_outputs(1981) <= not a;
    layer2_outputs(1982) <= a and b;
    layer2_outputs(1983) <= b and not a;
    layer2_outputs(1984) <= not (a xor b);
    layer2_outputs(1985) <= not a;
    layer2_outputs(1986) <= not (a and b);
    layer2_outputs(1987) <= not (a xor b);
    layer2_outputs(1988) <= b and not a;
    layer2_outputs(1989) <= a xor b;
    layer2_outputs(1990) <= 1'b0;
    layer2_outputs(1991) <= a or b;
    layer2_outputs(1992) <= not a or b;
    layer2_outputs(1993) <= not (a or b);
    layer2_outputs(1994) <= b;
    layer2_outputs(1995) <= 1'b1;
    layer2_outputs(1996) <= not b;
    layer2_outputs(1997) <= 1'b1;
    layer2_outputs(1998) <= not (a or b);
    layer2_outputs(1999) <= 1'b0;
    layer2_outputs(2000) <= not (a xor b);
    layer2_outputs(2001) <= not (a xor b);
    layer2_outputs(2002) <= a and not b;
    layer2_outputs(2003) <= 1'b1;
    layer2_outputs(2004) <= a and b;
    layer2_outputs(2005) <= not (a or b);
    layer2_outputs(2006) <= a and b;
    layer2_outputs(2007) <= a and not b;
    layer2_outputs(2008) <= not b or a;
    layer2_outputs(2009) <= a or b;
    layer2_outputs(2010) <= 1'b0;
    layer2_outputs(2011) <= not (a or b);
    layer2_outputs(2012) <= not (a xor b);
    layer2_outputs(2013) <= not b or a;
    layer2_outputs(2014) <= not b or a;
    layer2_outputs(2015) <= not a or b;
    layer2_outputs(2016) <= a;
    layer2_outputs(2017) <= not a or b;
    layer2_outputs(2018) <= a;
    layer2_outputs(2019) <= 1'b1;
    layer2_outputs(2020) <= 1'b1;
    layer2_outputs(2021) <= not (a or b);
    layer2_outputs(2022) <= a and b;
    layer2_outputs(2023) <= a and not b;
    layer2_outputs(2024) <= not b or a;
    layer2_outputs(2025) <= a or b;
    layer2_outputs(2026) <= not a or b;
    layer2_outputs(2027) <= a;
    layer2_outputs(2028) <= a and not b;
    layer2_outputs(2029) <= 1'b0;
    layer2_outputs(2030) <= not (a or b);
    layer2_outputs(2031) <= not a;
    layer2_outputs(2032) <= not b or a;
    layer2_outputs(2033) <= 1'b1;
    layer2_outputs(2034) <= a or b;
    layer2_outputs(2035) <= a;
    layer2_outputs(2036) <= not a;
    layer2_outputs(2037) <= 1'b1;
    layer2_outputs(2038) <= 1'b1;
    layer2_outputs(2039) <= b and not a;
    layer2_outputs(2040) <= not b;
    layer2_outputs(2041) <= 1'b1;
    layer2_outputs(2042) <= not b or a;
    layer2_outputs(2043) <= a or b;
    layer2_outputs(2044) <= b and not a;
    layer2_outputs(2045) <= not (a or b);
    layer2_outputs(2046) <= not a or b;
    layer2_outputs(2047) <= a;
    layer2_outputs(2048) <= not (a and b);
    layer2_outputs(2049) <= not (a and b);
    layer2_outputs(2050) <= 1'b0;
    layer2_outputs(2051) <= 1'b0;
    layer2_outputs(2052) <= not a or b;
    layer2_outputs(2053) <= 1'b1;
    layer2_outputs(2054) <= b and not a;
    layer2_outputs(2055) <= b and not a;
    layer2_outputs(2056) <= b;
    layer2_outputs(2057) <= b;
    layer2_outputs(2058) <= not (a or b);
    layer2_outputs(2059) <= not b;
    layer2_outputs(2060) <= a and not b;
    layer2_outputs(2061) <= 1'b0;
    layer2_outputs(2062) <= a or b;
    layer2_outputs(2063) <= 1'b0;
    layer2_outputs(2064) <= 1'b0;
    layer2_outputs(2065) <= not (a or b);
    layer2_outputs(2066) <= 1'b0;
    layer2_outputs(2067) <= not a;
    layer2_outputs(2068) <= 1'b1;
    layer2_outputs(2069) <= b;
    layer2_outputs(2070) <= 1'b0;
    layer2_outputs(2071) <= a and b;
    layer2_outputs(2072) <= b and not a;
    layer2_outputs(2073) <= 1'b0;
    layer2_outputs(2074) <= not (a and b);
    layer2_outputs(2075) <= a or b;
    layer2_outputs(2076) <= a;
    layer2_outputs(2077) <= not (a and b);
    layer2_outputs(2078) <= a and b;
    layer2_outputs(2079) <= a xor b;
    layer2_outputs(2080) <= 1'b0;
    layer2_outputs(2081) <= a and b;
    layer2_outputs(2082) <= not a;
    layer2_outputs(2083) <= 1'b1;
    layer2_outputs(2084) <= not (a and b);
    layer2_outputs(2085) <= not a;
    layer2_outputs(2086) <= not a or b;
    layer2_outputs(2087) <= b and not a;
    layer2_outputs(2088) <= 1'b1;
    layer2_outputs(2089) <= b;
    layer2_outputs(2090) <= 1'b0;
    layer2_outputs(2091) <= not b or a;
    layer2_outputs(2092) <= not a;
    layer2_outputs(2093) <= not (a and b);
    layer2_outputs(2094) <= not b or a;
    layer2_outputs(2095) <= a xor b;
    layer2_outputs(2096) <= b and not a;
    layer2_outputs(2097) <= not b or a;
    layer2_outputs(2098) <= a xor b;
    layer2_outputs(2099) <= b and not a;
    layer2_outputs(2100) <= a or b;
    layer2_outputs(2101) <= a and b;
    layer2_outputs(2102) <= not a;
    layer2_outputs(2103) <= a;
    layer2_outputs(2104) <= not a;
    layer2_outputs(2105) <= 1'b0;
    layer2_outputs(2106) <= a xor b;
    layer2_outputs(2107) <= a and not b;
    layer2_outputs(2108) <= b;
    layer2_outputs(2109) <= not a;
    layer2_outputs(2110) <= not (a and b);
    layer2_outputs(2111) <= a;
    layer2_outputs(2112) <= not (a and b);
    layer2_outputs(2113) <= b and not a;
    layer2_outputs(2114) <= 1'b0;
    layer2_outputs(2115) <= 1'b0;
    layer2_outputs(2116) <= not (a and b);
    layer2_outputs(2117) <= not b;
    layer2_outputs(2118) <= 1'b1;
    layer2_outputs(2119) <= not a;
    layer2_outputs(2120) <= a or b;
    layer2_outputs(2121) <= 1'b0;
    layer2_outputs(2122) <= not (a or b);
    layer2_outputs(2123) <= not b or a;
    layer2_outputs(2124) <= a and b;
    layer2_outputs(2125) <= b and not a;
    layer2_outputs(2126) <= not (a or b);
    layer2_outputs(2127) <= 1'b0;
    layer2_outputs(2128) <= a and b;
    layer2_outputs(2129) <= a and not b;
    layer2_outputs(2130) <= 1'b1;
    layer2_outputs(2131) <= a;
    layer2_outputs(2132) <= a and b;
    layer2_outputs(2133) <= not (a and b);
    layer2_outputs(2134) <= not b;
    layer2_outputs(2135) <= 1'b1;
    layer2_outputs(2136) <= 1'b0;
    layer2_outputs(2137) <= a or b;
    layer2_outputs(2138) <= 1'b0;
    layer2_outputs(2139) <= 1'b1;
    layer2_outputs(2140) <= not b or a;
    layer2_outputs(2141) <= b;
    layer2_outputs(2142) <= not (a and b);
    layer2_outputs(2143) <= a;
    layer2_outputs(2144) <= a or b;
    layer2_outputs(2145) <= a;
    layer2_outputs(2146) <= 1'b0;
    layer2_outputs(2147) <= not (a or b);
    layer2_outputs(2148) <= not a;
    layer2_outputs(2149) <= 1'b0;
    layer2_outputs(2150) <= not (a and b);
    layer2_outputs(2151) <= 1'b1;
    layer2_outputs(2152) <= not (a or b);
    layer2_outputs(2153) <= not (a or b);
    layer2_outputs(2154) <= not (a xor b);
    layer2_outputs(2155) <= a and b;
    layer2_outputs(2156) <= a;
    layer2_outputs(2157) <= a and not b;
    layer2_outputs(2158) <= not b or a;
    layer2_outputs(2159) <= a or b;
    layer2_outputs(2160) <= b;
    layer2_outputs(2161) <= not (a or b);
    layer2_outputs(2162) <= a;
    layer2_outputs(2163) <= a;
    layer2_outputs(2164) <= not b or a;
    layer2_outputs(2165) <= b and not a;
    layer2_outputs(2166) <= not b;
    layer2_outputs(2167) <= b;
    layer2_outputs(2168) <= 1'b0;
    layer2_outputs(2169) <= b and not a;
    layer2_outputs(2170) <= not a or b;
    layer2_outputs(2171) <= not a or b;
    layer2_outputs(2172) <= 1'b0;
    layer2_outputs(2173) <= not b;
    layer2_outputs(2174) <= a and b;
    layer2_outputs(2175) <= 1'b0;
    layer2_outputs(2176) <= not (a or b);
    layer2_outputs(2177) <= not (a or b);
    layer2_outputs(2178) <= 1'b1;
    layer2_outputs(2179) <= 1'b1;
    layer2_outputs(2180) <= 1'b0;
    layer2_outputs(2181) <= not a;
    layer2_outputs(2182) <= 1'b0;
    layer2_outputs(2183) <= 1'b1;
    layer2_outputs(2184) <= a and not b;
    layer2_outputs(2185) <= 1'b1;
    layer2_outputs(2186) <= 1'b1;
    layer2_outputs(2187) <= b and not a;
    layer2_outputs(2188) <= not (a or b);
    layer2_outputs(2189) <= not b;
    layer2_outputs(2190) <= not b or a;
    layer2_outputs(2191) <= 1'b0;
    layer2_outputs(2192) <= not (a and b);
    layer2_outputs(2193) <= a or b;
    layer2_outputs(2194) <= a and b;
    layer2_outputs(2195) <= a or b;
    layer2_outputs(2196) <= not (a and b);
    layer2_outputs(2197) <= 1'b0;
    layer2_outputs(2198) <= 1'b1;
    layer2_outputs(2199) <= not (a and b);
    layer2_outputs(2200) <= 1'b0;
    layer2_outputs(2201) <= a and not b;
    layer2_outputs(2202) <= not a;
    layer2_outputs(2203) <= a xor b;
    layer2_outputs(2204) <= 1'b1;
    layer2_outputs(2205) <= 1'b0;
    layer2_outputs(2206) <= 1'b0;
    layer2_outputs(2207) <= not b or a;
    layer2_outputs(2208) <= 1'b1;
    layer2_outputs(2209) <= a and b;
    layer2_outputs(2210) <= b;
    layer2_outputs(2211) <= not b or a;
    layer2_outputs(2212) <= not (a and b);
    layer2_outputs(2213) <= not a;
    layer2_outputs(2214) <= not a or b;
    layer2_outputs(2215) <= not (a and b);
    layer2_outputs(2216) <= b;
    layer2_outputs(2217) <= 1'b1;
    layer2_outputs(2218) <= 1'b0;
    layer2_outputs(2219) <= 1'b1;
    layer2_outputs(2220) <= b and not a;
    layer2_outputs(2221) <= b and not a;
    layer2_outputs(2222) <= a or b;
    layer2_outputs(2223) <= not (a or b);
    layer2_outputs(2224) <= b and not a;
    layer2_outputs(2225) <= not a or b;
    layer2_outputs(2226) <= 1'b0;
    layer2_outputs(2227) <= a and not b;
    layer2_outputs(2228) <= not (a and b);
    layer2_outputs(2229) <= not b;
    layer2_outputs(2230) <= a;
    layer2_outputs(2231) <= a and b;
    layer2_outputs(2232) <= not a;
    layer2_outputs(2233) <= not a;
    layer2_outputs(2234) <= 1'b0;
    layer2_outputs(2235) <= 1'b1;
    layer2_outputs(2236) <= a and b;
    layer2_outputs(2237) <= not (a or b);
    layer2_outputs(2238) <= not (a and b);
    layer2_outputs(2239) <= not a or b;
    layer2_outputs(2240) <= not b;
    layer2_outputs(2241) <= a and not b;
    layer2_outputs(2242) <= not a;
    layer2_outputs(2243) <= b;
    layer2_outputs(2244) <= b and not a;
    layer2_outputs(2245) <= b and not a;
    layer2_outputs(2246) <= not a or b;
    layer2_outputs(2247) <= not b or a;
    layer2_outputs(2248) <= a;
    layer2_outputs(2249) <= not b;
    layer2_outputs(2250) <= a;
    layer2_outputs(2251) <= a xor b;
    layer2_outputs(2252) <= not (a and b);
    layer2_outputs(2253) <= a and not b;
    layer2_outputs(2254) <= a;
    layer2_outputs(2255) <= b and not a;
    layer2_outputs(2256) <= not a or b;
    layer2_outputs(2257) <= a and not b;
    layer2_outputs(2258) <= 1'b1;
    layer2_outputs(2259) <= not a;
    layer2_outputs(2260) <= 1'b1;
    layer2_outputs(2261) <= 1'b1;
    layer2_outputs(2262) <= not b;
    layer2_outputs(2263) <= 1'b0;
    layer2_outputs(2264) <= not b;
    layer2_outputs(2265) <= a or b;
    layer2_outputs(2266) <= a and not b;
    layer2_outputs(2267) <= b and not a;
    layer2_outputs(2268) <= not (a or b);
    layer2_outputs(2269) <= not b or a;
    layer2_outputs(2270) <= a;
    layer2_outputs(2271) <= 1'b0;
    layer2_outputs(2272) <= not a;
    layer2_outputs(2273) <= b and not a;
    layer2_outputs(2274) <= not (a and b);
    layer2_outputs(2275) <= not b or a;
    layer2_outputs(2276) <= a and not b;
    layer2_outputs(2277) <= 1'b0;
    layer2_outputs(2278) <= a and not b;
    layer2_outputs(2279) <= not a or b;
    layer2_outputs(2280) <= not (a or b);
    layer2_outputs(2281) <= not b or a;
    layer2_outputs(2282) <= a and b;
    layer2_outputs(2283) <= not a or b;
    layer2_outputs(2284) <= a and b;
    layer2_outputs(2285) <= b;
    layer2_outputs(2286) <= 1'b1;
    layer2_outputs(2287) <= b;
    layer2_outputs(2288) <= 1'b0;
    layer2_outputs(2289) <= a and not b;
    layer2_outputs(2290) <= not a;
    layer2_outputs(2291) <= 1'b0;
    layer2_outputs(2292) <= not a or b;
    layer2_outputs(2293) <= not a or b;
    layer2_outputs(2294) <= 1'b0;
    layer2_outputs(2295) <= not b;
    layer2_outputs(2296) <= a and b;
    layer2_outputs(2297) <= 1'b0;
    layer2_outputs(2298) <= not a or b;
    layer2_outputs(2299) <= b and not a;
    layer2_outputs(2300) <= a and b;
    layer2_outputs(2301) <= not b;
    layer2_outputs(2302) <= b;
    layer2_outputs(2303) <= not (a and b);
    layer2_outputs(2304) <= not a;
    layer2_outputs(2305) <= not a;
    layer2_outputs(2306) <= b and not a;
    layer2_outputs(2307) <= a and b;
    layer2_outputs(2308) <= 1'b1;
    layer2_outputs(2309) <= 1'b0;
    layer2_outputs(2310) <= not b;
    layer2_outputs(2311) <= a and b;
    layer2_outputs(2312) <= not a or b;
    layer2_outputs(2313) <= 1'b1;
    layer2_outputs(2314) <= not a;
    layer2_outputs(2315) <= not (a or b);
    layer2_outputs(2316) <= 1'b1;
    layer2_outputs(2317) <= not a or b;
    layer2_outputs(2318) <= not a;
    layer2_outputs(2319) <= not (a xor b);
    layer2_outputs(2320) <= not (a or b);
    layer2_outputs(2321) <= not (a and b);
    layer2_outputs(2322) <= not (a and b);
    layer2_outputs(2323) <= b and not a;
    layer2_outputs(2324) <= 1'b1;
    layer2_outputs(2325) <= b and not a;
    layer2_outputs(2326) <= a or b;
    layer2_outputs(2327) <= a and b;
    layer2_outputs(2328) <= a and not b;
    layer2_outputs(2329) <= not a or b;
    layer2_outputs(2330) <= b and not a;
    layer2_outputs(2331) <= not (a xor b);
    layer2_outputs(2332) <= b;
    layer2_outputs(2333) <= not a;
    layer2_outputs(2334) <= b;
    layer2_outputs(2335) <= not a;
    layer2_outputs(2336) <= a;
    layer2_outputs(2337) <= not (a or b);
    layer2_outputs(2338) <= a and b;
    layer2_outputs(2339) <= a or b;
    layer2_outputs(2340) <= 1'b0;
    layer2_outputs(2341) <= not a;
    layer2_outputs(2342) <= 1'b0;
    layer2_outputs(2343) <= 1'b0;
    layer2_outputs(2344) <= not b or a;
    layer2_outputs(2345) <= 1'b0;
    layer2_outputs(2346) <= b and not a;
    layer2_outputs(2347) <= not a or b;
    layer2_outputs(2348) <= not a;
    layer2_outputs(2349) <= 1'b1;
    layer2_outputs(2350) <= a and b;
    layer2_outputs(2351) <= a or b;
    layer2_outputs(2352) <= not a;
    layer2_outputs(2353) <= a xor b;
    layer2_outputs(2354) <= b;
    layer2_outputs(2355) <= a or b;
    layer2_outputs(2356) <= a and b;
    layer2_outputs(2357) <= not b or a;
    layer2_outputs(2358) <= a xor b;
    layer2_outputs(2359) <= a and b;
    layer2_outputs(2360) <= a and b;
    layer2_outputs(2361) <= not a or b;
    layer2_outputs(2362) <= 1'b1;
    layer2_outputs(2363) <= 1'b1;
    layer2_outputs(2364) <= not (a or b);
    layer2_outputs(2365) <= a;
    layer2_outputs(2366) <= 1'b1;
    layer2_outputs(2367) <= b;
    layer2_outputs(2368) <= not a or b;
    layer2_outputs(2369) <= 1'b1;
    layer2_outputs(2370) <= 1'b1;
    layer2_outputs(2371) <= not a or b;
    layer2_outputs(2372) <= b and not a;
    layer2_outputs(2373) <= not b;
    layer2_outputs(2374) <= 1'b0;
    layer2_outputs(2375) <= not (a xor b);
    layer2_outputs(2376) <= not b;
    layer2_outputs(2377) <= a and b;
    layer2_outputs(2378) <= a and b;
    layer2_outputs(2379) <= b;
    layer2_outputs(2380) <= not a;
    layer2_outputs(2381) <= not (a and b);
    layer2_outputs(2382) <= a;
    layer2_outputs(2383) <= 1'b0;
    layer2_outputs(2384) <= b and not a;
    layer2_outputs(2385) <= not b;
    layer2_outputs(2386) <= a and not b;
    layer2_outputs(2387) <= not (a or b);
    layer2_outputs(2388) <= not b or a;
    layer2_outputs(2389) <= not (a xor b);
    layer2_outputs(2390) <= a or b;
    layer2_outputs(2391) <= not b;
    layer2_outputs(2392) <= not (a or b);
    layer2_outputs(2393) <= a and not b;
    layer2_outputs(2394) <= not b;
    layer2_outputs(2395) <= a and not b;
    layer2_outputs(2396) <= a and not b;
    layer2_outputs(2397) <= not (a xor b);
    layer2_outputs(2398) <= a and b;
    layer2_outputs(2399) <= b and not a;
    layer2_outputs(2400) <= not b;
    layer2_outputs(2401) <= 1'b1;
    layer2_outputs(2402) <= a or b;
    layer2_outputs(2403) <= b and not a;
    layer2_outputs(2404) <= a;
    layer2_outputs(2405) <= b and not a;
    layer2_outputs(2406) <= b;
    layer2_outputs(2407) <= not a;
    layer2_outputs(2408) <= not (a or b);
    layer2_outputs(2409) <= a and b;
    layer2_outputs(2410) <= 1'b1;
    layer2_outputs(2411) <= not (a and b);
    layer2_outputs(2412) <= not b;
    layer2_outputs(2413) <= a xor b;
    layer2_outputs(2414) <= not b;
    layer2_outputs(2415) <= 1'b0;
    layer2_outputs(2416) <= not (a and b);
    layer2_outputs(2417) <= not b;
    layer2_outputs(2418) <= not a;
    layer2_outputs(2419) <= b and not a;
    layer2_outputs(2420) <= b;
    layer2_outputs(2421) <= b and not a;
    layer2_outputs(2422) <= not (a and b);
    layer2_outputs(2423) <= a or b;
    layer2_outputs(2424) <= a;
    layer2_outputs(2425) <= b and not a;
    layer2_outputs(2426) <= 1'b0;
    layer2_outputs(2427) <= 1'b1;
    layer2_outputs(2428) <= a or b;
    layer2_outputs(2429) <= 1'b0;
    layer2_outputs(2430) <= not (a or b);
    layer2_outputs(2431) <= 1'b1;
    layer2_outputs(2432) <= not b or a;
    layer2_outputs(2433) <= a or b;
    layer2_outputs(2434) <= b;
    layer2_outputs(2435) <= not a;
    layer2_outputs(2436) <= b;
    layer2_outputs(2437) <= a and b;
    layer2_outputs(2438) <= a or b;
    layer2_outputs(2439) <= not (a or b);
    layer2_outputs(2440) <= not a or b;
    layer2_outputs(2441) <= a or b;
    layer2_outputs(2442) <= not a or b;
    layer2_outputs(2443) <= not (a or b);
    layer2_outputs(2444) <= 1'b1;
    layer2_outputs(2445) <= not b or a;
    layer2_outputs(2446) <= not a or b;
    layer2_outputs(2447) <= a or b;
    layer2_outputs(2448) <= not (a xor b);
    layer2_outputs(2449) <= 1'b1;
    layer2_outputs(2450) <= 1'b1;
    layer2_outputs(2451) <= a and not b;
    layer2_outputs(2452) <= not (a and b);
    layer2_outputs(2453) <= not b or a;
    layer2_outputs(2454) <= not (a or b);
    layer2_outputs(2455) <= not (a and b);
    layer2_outputs(2456) <= not (a or b);
    layer2_outputs(2457) <= a or b;
    layer2_outputs(2458) <= not b or a;
    layer2_outputs(2459) <= not b or a;
    layer2_outputs(2460) <= not b or a;
    layer2_outputs(2461) <= a and not b;
    layer2_outputs(2462) <= a or b;
    layer2_outputs(2463) <= 1'b0;
    layer2_outputs(2464) <= a and b;
    layer2_outputs(2465) <= not a;
    layer2_outputs(2466) <= b;
    layer2_outputs(2467) <= not a or b;
    layer2_outputs(2468) <= a and not b;
    layer2_outputs(2469) <= not a or b;
    layer2_outputs(2470) <= 1'b0;
    layer2_outputs(2471) <= a;
    layer2_outputs(2472) <= not (a and b);
    layer2_outputs(2473) <= not a;
    layer2_outputs(2474) <= a and not b;
    layer2_outputs(2475) <= b;
    layer2_outputs(2476) <= a;
    layer2_outputs(2477) <= b;
    layer2_outputs(2478) <= b and not a;
    layer2_outputs(2479) <= 1'b1;
    layer2_outputs(2480) <= 1'b0;
    layer2_outputs(2481) <= a;
    layer2_outputs(2482) <= 1'b1;
    layer2_outputs(2483) <= b and not a;
    layer2_outputs(2484) <= not a or b;
    layer2_outputs(2485) <= not (a and b);
    layer2_outputs(2486) <= a;
    layer2_outputs(2487) <= b and not a;
    layer2_outputs(2488) <= b and not a;
    layer2_outputs(2489) <= not a or b;
    layer2_outputs(2490) <= not (a or b);
    layer2_outputs(2491) <= a;
    layer2_outputs(2492) <= b;
    layer2_outputs(2493) <= not (a and b);
    layer2_outputs(2494) <= not b or a;
    layer2_outputs(2495) <= b;
    layer2_outputs(2496) <= a or b;
    layer2_outputs(2497) <= a and b;
    layer2_outputs(2498) <= 1'b1;
    layer2_outputs(2499) <= a;
    layer2_outputs(2500) <= not a or b;
    layer2_outputs(2501) <= not b;
    layer2_outputs(2502) <= a and b;
    layer2_outputs(2503) <= b;
    layer2_outputs(2504) <= not (a or b);
    layer2_outputs(2505) <= not a or b;
    layer2_outputs(2506) <= not (a and b);
    layer2_outputs(2507) <= not b or a;
    layer2_outputs(2508) <= b and not a;
    layer2_outputs(2509) <= a and b;
    layer2_outputs(2510) <= not a or b;
    layer2_outputs(2511) <= a and not b;
    layer2_outputs(2512) <= a and b;
    layer2_outputs(2513) <= not b or a;
    layer2_outputs(2514) <= not a or b;
    layer2_outputs(2515) <= 1'b1;
    layer2_outputs(2516) <= not b;
    layer2_outputs(2517) <= b and not a;
    layer2_outputs(2518) <= a;
    layer2_outputs(2519) <= a and not b;
    layer2_outputs(2520) <= not b;
    layer2_outputs(2521) <= not (a or b);
    layer2_outputs(2522) <= b and not a;
    layer2_outputs(2523) <= a and not b;
    layer2_outputs(2524) <= a and not b;
    layer2_outputs(2525) <= 1'b1;
    layer2_outputs(2526) <= b and not a;
    layer2_outputs(2527) <= 1'b1;
    layer2_outputs(2528) <= a and not b;
    layer2_outputs(2529) <= a or b;
    layer2_outputs(2530) <= a;
    layer2_outputs(2531) <= 1'b1;
    layer2_outputs(2532) <= b and not a;
    layer2_outputs(2533) <= not (a or b);
    layer2_outputs(2534) <= not (a xor b);
    layer2_outputs(2535) <= not (a or b);
    layer2_outputs(2536) <= a and not b;
    layer2_outputs(2537) <= a and b;
    layer2_outputs(2538) <= not b;
    layer2_outputs(2539) <= a and b;
    layer2_outputs(2540) <= 1'b0;
    layer2_outputs(2541) <= a and b;
    layer2_outputs(2542) <= a or b;
    layer2_outputs(2543) <= 1'b1;
    layer2_outputs(2544) <= not b;
    layer2_outputs(2545) <= a and not b;
    layer2_outputs(2546) <= not a or b;
    layer2_outputs(2547) <= 1'b0;
    layer2_outputs(2548) <= 1'b1;
    layer2_outputs(2549) <= not b or a;
    layer2_outputs(2550) <= a and not b;
    layer2_outputs(2551) <= a and not b;
    layer2_outputs(2552) <= 1'b1;
    layer2_outputs(2553) <= not a or b;
    layer2_outputs(2554) <= 1'b1;
    layer2_outputs(2555) <= a and b;
    layer2_outputs(2556) <= not a or b;
    layer2_outputs(2557) <= a and b;
    layer2_outputs(2558) <= not (a or b);
    layer2_outputs(2559) <= a or b;
    layer3_outputs(0) <= not a or b;
    layer3_outputs(1) <= b;
    layer3_outputs(2) <= a and b;
    layer3_outputs(3) <= not b or a;
    layer3_outputs(4) <= b and not a;
    layer3_outputs(5) <= not (a and b);
    layer3_outputs(6) <= a and not b;
    layer3_outputs(7) <= not b;
    layer3_outputs(8) <= b and not a;
    layer3_outputs(9) <= not a or b;
    layer3_outputs(10) <= a;
    layer3_outputs(11) <= a or b;
    layer3_outputs(12) <= not a or b;
    layer3_outputs(13) <= 1'b0;
    layer3_outputs(14) <= not (a or b);
    layer3_outputs(15) <= not a or b;
    layer3_outputs(16) <= 1'b0;
    layer3_outputs(17) <= not a or b;
    layer3_outputs(18) <= not (a or b);
    layer3_outputs(19) <= a;
    layer3_outputs(20) <= a and b;
    layer3_outputs(21) <= a and not b;
    layer3_outputs(22) <= b and not a;
    layer3_outputs(23) <= 1'b1;
    layer3_outputs(24) <= not b;
    layer3_outputs(25) <= not a;
    layer3_outputs(26) <= 1'b0;
    layer3_outputs(27) <= not (a or b);
    layer3_outputs(28) <= b;
    layer3_outputs(29) <= a or b;
    layer3_outputs(30) <= not (a and b);
    layer3_outputs(31) <= a or b;
    layer3_outputs(32) <= a and not b;
    layer3_outputs(33) <= not a;
    layer3_outputs(34) <= not (a and b);
    layer3_outputs(35) <= a and b;
    layer3_outputs(36) <= a and not b;
    layer3_outputs(37) <= a and not b;
    layer3_outputs(38) <= a and b;
    layer3_outputs(39) <= 1'b0;
    layer3_outputs(40) <= a or b;
    layer3_outputs(41) <= not (a and b);
    layer3_outputs(42) <= 1'b0;
    layer3_outputs(43) <= a;
    layer3_outputs(44) <= not a;
    layer3_outputs(45) <= not a or b;
    layer3_outputs(46) <= 1'b0;
    layer3_outputs(47) <= a;
    layer3_outputs(48) <= a and not b;
    layer3_outputs(49) <= b;
    layer3_outputs(50) <= b;
    layer3_outputs(51) <= not a or b;
    layer3_outputs(52) <= 1'b0;
    layer3_outputs(53) <= 1'b0;
    layer3_outputs(54) <= a or b;
    layer3_outputs(55) <= not (a or b);
    layer3_outputs(56) <= a and not b;
    layer3_outputs(57) <= a and not b;
    layer3_outputs(58) <= a and b;
    layer3_outputs(59) <= 1'b0;
    layer3_outputs(60) <= a and not b;
    layer3_outputs(61) <= not (a or b);
    layer3_outputs(62) <= not b;
    layer3_outputs(63) <= not (a and b);
    layer3_outputs(64) <= b and not a;
    layer3_outputs(65) <= not a or b;
    layer3_outputs(66) <= 1'b1;
    layer3_outputs(67) <= a and b;
    layer3_outputs(68) <= a or b;
    layer3_outputs(69) <= not (a or b);
    layer3_outputs(70) <= not b;
    layer3_outputs(71) <= not b or a;
    layer3_outputs(72) <= a and not b;
    layer3_outputs(73) <= not (a or b);
    layer3_outputs(74) <= not (a and b);
    layer3_outputs(75) <= 1'b0;
    layer3_outputs(76) <= not (a or b);
    layer3_outputs(77) <= a;
    layer3_outputs(78) <= a and b;
    layer3_outputs(79) <= a and b;
    layer3_outputs(80) <= not a or b;
    layer3_outputs(81) <= a and not b;
    layer3_outputs(82) <= not a or b;
    layer3_outputs(83) <= not a;
    layer3_outputs(84) <= 1'b0;
    layer3_outputs(85) <= not b or a;
    layer3_outputs(86) <= a;
    layer3_outputs(87) <= a and not b;
    layer3_outputs(88) <= not a;
    layer3_outputs(89) <= not b or a;
    layer3_outputs(90) <= not b or a;
    layer3_outputs(91) <= 1'b0;
    layer3_outputs(92) <= b and not a;
    layer3_outputs(93) <= b and not a;
    layer3_outputs(94) <= a;
    layer3_outputs(95) <= 1'b0;
    layer3_outputs(96) <= not a;
    layer3_outputs(97) <= a and not b;
    layer3_outputs(98) <= 1'b1;
    layer3_outputs(99) <= a and b;
    layer3_outputs(100) <= a or b;
    layer3_outputs(101) <= not (a or b);
    layer3_outputs(102) <= 1'b1;
    layer3_outputs(103) <= 1'b1;
    layer3_outputs(104) <= b;
    layer3_outputs(105) <= not (a or b);
    layer3_outputs(106) <= a and not b;
    layer3_outputs(107) <= 1'b1;
    layer3_outputs(108) <= not a or b;
    layer3_outputs(109) <= not (a and b);
    layer3_outputs(110) <= 1'b1;
    layer3_outputs(111) <= not b;
    layer3_outputs(112) <= not b or a;
    layer3_outputs(113) <= a;
    layer3_outputs(114) <= b and not a;
    layer3_outputs(115) <= b;
    layer3_outputs(116) <= a or b;
    layer3_outputs(117) <= not a or b;
    layer3_outputs(118) <= 1'b1;
    layer3_outputs(119) <= 1'b0;
    layer3_outputs(120) <= 1'b1;
    layer3_outputs(121) <= b;
    layer3_outputs(122) <= 1'b1;
    layer3_outputs(123) <= a and b;
    layer3_outputs(124) <= 1'b0;
    layer3_outputs(125) <= a and not b;
    layer3_outputs(126) <= a and b;
    layer3_outputs(127) <= a and not b;
    layer3_outputs(128) <= 1'b1;
    layer3_outputs(129) <= 1'b0;
    layer3_outputs(130) <= 1'b0;
    layer3_outputs(131) <= b;
    layer3_outputs(132) <= 1'b1;
    layer3_outputs(133) <= 1'b1;
    layer3_outputs(134) <= not b or a;
    layer3_outputs(135) <= a and not b;
    layer3_outputs(136) <= a and b;
    layer3_outputs(137) <= not b;
    layer3_outputs(138) <= 1'b1;
    layer3_outputs(139) <= not (a or b);
    layer3_outputs(140) <= not b or a;
    layer3_outputs(141) <= not (a or b);
    layer3_outputs(142) <= a or b;
    layer3_outputs(143) <= a and b;
    layer3_outputs(144) <= not (a or b);
    layer3_outputs(145) <= a and b;
    layer3_outputs(146) <= not (a or b);
    layer3_outputs(147) <= not (a or b);
    layer3_outputs(148) <= a;
    layer3_outputs(149) <= not b;
    layer3_outputs(150) <= not (a and b);
    layer3_outputs(151) <= not b;
    layer3_outputs(152) <= a or b;
    layer3_outputs(153) <= a and b;
    layer3_outputs(154) <= a;
    layer3_outputs(155) <= 1'b1;
    layer3_outputs(156) <= a or b;
    layer3_outputs(157) <= a xor b;
    layer3_outputs(158) <= not (a or b);
    layer3_outputs(159) <= not b or a;
    layer3_outputs(160) <= 1'b1;
    layer3_outputs(161) <= a and b;
    layer3_outputs(162) <= 1'b1;
    layer3_outputs(163) <= not a or b;
    layer3_outputs(164) <= not (a and b);
    layer3_outputs(165) <= a or b;
    layer3_outputs(166) <= a and not b;
    layer3_outputs(167) <= not b or a;
    layer3_outputs(168) <= not (a or b);
    layer3_outputs(169) <= 1'b1;
    layer3_outputs(170) <= not a;
    layer3_outputs(171) <= not a;
    layer3_outputs(172) <= b;
    layer3_outputs(173) <= not a;
    layer3_outputs(174) <= a and b;
    layer3_outputs(175) <= not a or b;
    layer3_outputs(176) <= a or b;
    layer3_outputs(177) <= a and b;
    layer3_outputs(178) <= not b;
    layer3_outputs(179) <= b;
    layer3_outputs(180) <= not a or b;
    layer3_outputs(181) <= a and not b;
    layer3_outputs(182) <= not (a or b);
    layer3_outputs(183) <= not (a xor b);
    layer3_outputs(184) <= a and not b;
    layer3_outputs(185) <= not b or a;
    layer3_outputs(186) <= not (a and b);
    layer3_outputs(187) <= a and not b;
    layer3_outputs(188) <= not (a and b);
    layer3_outputs(189) <= a or b;
    layer3_outputs(190) <= 1'b0;
    layer3_outputs(191) <= not a or b;
    layer3_outputs(192) <= b and not a;
    layer3_outputs(193) <= not b or a;
    layer3_outputs(194) <= a and b;
    layer3_outputs(195) <= a and not b;
    layer3_outputs(196) <= a xor b;
    layer3_outputs(197) <= 1'b1;
    layer3_outputs(198) <= a or b;
    layer3_outputs(199) <= b and not a;
    layer3_outputs(200) <= a and not b;
    layer3_outputs(201) <= not a or b;
    layer3_outputs(202) <= b and not a;
    layer3_outputs(203) <= not b or a;
    layer3_outputs(204) <= a;
    layer3_outputs(205) <= 1'b0;
    layer3_outputs(206) <= b and not a;
    layer3_outputs(207) <= not b;
    layer3_outputs(208) <= not b;
    layer3_outputs(209) <= a;
    layer3_outputs(210) <= not (a or b);
    layer3_outputs(211) <= not b or a;
    layer3_outputs(212) <= a and not b;
    layer3_outputs(213) <= not b or a;
    layer3_outputs(214) <= not b or a;
    layer3_outputs(215) <= b and not a;
    layer3_outputs(216) <= not b;
    layer3_outputs(217) <= not b or a;
    layer3_outputs(218) <= not b;
    layer3_outputs(219) <= not (a or b);
    layer3_outputs(220) <= 1'b0;
    layer3_outputs(221) <= b;
    layer3_outputs(222) <= not a or b;
    layer3_outputs(223) <= 1'b0;
    layer3_outputs(224) <= not (a or b);
    layer3_outputs(225) <= 1'b0;
    layer3_outputs(226) <= a and not b;
    layer3_outputs(227) <= a;
    layer3_outputs(228) <= a or b;
    layer3_outputs(229) <= a or b;
    layer3_outputs(230) <= not (a or b);
    layer3_outputs(231) <= not (a and b);
    layer3_outputs(232) <= not (a xor b);
    layer3_outputs(233) <= not (a xor b);
    layer3_outputs(234) <= a or b;
    layer3_outputs(235) <= 1'b1;
    layer3_outputs(236) <= 1'b1;
    layer3_outputs(237) <= not a;
    layer3_outputs(238) <= b and not a;
    layer3_outputs(239) <= a;
    layer3_outputs(240) <= a xor b;
    layer3_outputs(241) <= 1'b0;
    layer3_outputs(242) <= a and b;
    layer3_outputs(243) <= not a or b;
    layer3_outputs(244) <= 1'b0;
    layer3_outputs(245) <= not (a and b);
    layer3_outputs(246) <= a or b;
    layer3_outputs(247) <= a or b;
    layer3_outputs(248) <= a and b;
    layer3_outputs(249) <= b and not a;
    layer3_outputs(250) <= not a or b;
    layer3_outputs(251) <= not b or a;
    layer3_outputs(252) <= a or b;
    layer3_outputs(253) <= 1'b1;
    layer3_outputs(254) <= not b;
    layer3_outputs(255) <= 1'b0;
    layer3_outputs(256) <= a or b;
    layer3_outputs(257) <= not (a or b);
    layer3_outputs(258) <= b;
    layer3_outputs(259) <= b;
    layer3_outputs(260) <= a and b;
    layer3_outputs(261) <= 1'b0;
    layer3_outputs(262) <= a or b;
    layer3_outputs(263) <= a xor b;
    layer3_outputs(264) <= not (a or b);
    layer3_outputs(265) <= not a or b;
    layer3_outputs(266) <= not b;
    layer3_outputs(267) <= a and not b;
    layer3_outputs(268) <= 1'b0;
    layer3_outputs(269) <= a;
    layer3_outputs(270) <= not (a and b);
    layer3_outputs(271) <= not (a and b);
    layer3_outputs(272) <= a and b;
    layer3_outputs(273) <= not a or b;
    layer3_outputs(274) <= 1'b0;
    layer3_outputs(275) <= not (a or b);
    layer3_outputs(276) <= b and not a;
    layer3_outputs(277) <= b and not a;
    layer3_outputs(278) <= not (a and b);
    layer3_outputs(279) <= b;
    layer3_outputs(280) <= not (a or b);
    layer3_outputs(281) <= b;
    layer3_outputs(282) <= not (a or b);
    layer3_outputs(283) <= a and not b;
    layer3_outputs(284) <= not b;
    layer3_outputs(285) <= a and not b;
    layer3_outputs(286) <= a and not b;
    layer3_outputs(287) <= not (a or b);
    layer3_outputs(288) <= 1'b0;
    layer3_outputs(289) <= a and not b;
    layer3_outputs(290) <= not b;
    layer3_outputs(291) <= not (a or b);
    layer3_outputs(292) <= b and not a;
    layer3_outputs(293) <= not a or b;
    layer3_outputs(294) <= not b;
    layer3_outputs(295) <= a;
    layer3_outputs(296) <= 1'b1;
    layer3_outputs(297) <= not a or b;
    layer3_outputs(298) <= b;
    layer3_outputs(299) <= a and b;
    layer3_outputs(300) <= not a or b;
    layer3_outputs(301) <= not b;
    layer3_outputs(302) <= 1'b0;
    layer3_outputs(303) <= b and not a;
    layer3_outputs(304) <= not a or b;
    layer3_outputs(305) <= not (a and b);
    layer3_outputs(306) <= a and b;
    layer3_outputs(307) <= not (a and b);
    layer3_outputs(308) <= not (a and b);
    layer3_outputs(309) <= 1'b1;
    layer3_outputs(310) <= a xor b;
    layer3_outputs(311) <= b and not a;
    layer3_outputs(312) <= not (a or b);
    layer3_outputs(313) <= a and b;
    layer3_outputs(314) <= not a or b;
    layer3_outputs(315) <= not a or b;
    layer3_outputs(316) <= 1'b1;
    layer3_outputs(317) <= a or b;
    layer3_outputs(318) <= not a or b;
    layer3_outputs(319) <= a and b;
    layer3_outputs(320) <= a and not b;
    layer3_outputs(321) <= not b;
    layer3_outputs(322) <= not a;
    layer3_outputs(323) <= a and b;
    layer3_outputs(324) <= not (a or b);
    layer3_outputs(325) <= not b;
    layer3_outputs(326) <= 1'b1;
    layer3_outputs(327) <= not (a and b);
    layer3_outputs(328) <= not b or a;
    layer3_outputs(329) <= a;
    layer3_outputs(330) <= not (a xor b);
    layer3_outputs(331) <= a and not b;
    layer3_outputs(332) <= a and b;
    layer3_outputs(333) <= not a or b;
    layer3_outputs(334) <= a and not b;
    layer3_outputs(335) <= 1'b0;
    layer3_outputs(336) <= 1'b0;
    layer3_outputs(337) <= a;
    layer3_outputs(338) <= 1'b0;
    layer3_outputs(339) <= not a or b;
    layer3_outputs(340) <= a;
    layer3_outputs(341) <= 1'b0;
    layer3_outputs(342) <= not b;
    layer3_outputs(343) <= b;
    layer3_outputs(344) <= not a;
    layer3_outputs(345) <= a or b;
    layer3_outputs(346) <= a or b;
    layer3_outputs(347) <= not a or b;
    layer3_outputs(348) <= a and b;
    layer3_outputs(349) <= a and not b;
    layer3_outputs(350) <= not a;
    layer3_outputs(351) <= a and not b;
    layer3_outputs(352) <= a or b;
    layer3_outputs(353) <= 1'b1;
    layer3_outputs(354) <= 1'b1;
    layer3_outputs(355) <= a;
    layer3_outputs(356) <= b and not a;
    layer3_outputs(357) <= not (a and b);
    layer3_outputs(358) <= not b or a;
    layer3_outputs(359) <= b and not a;
    layer3_outputs(360) <= a xor b;
    layer3_outputs(361) <= not b;
    layer3_outputs(362) <= not a;
    layer3_outputs(363) <= not (a and b);
    layer3_outputs(364) <= a and b;
    layer3_outputs(365) <= a and b;
    layer3_outputs(366) <= a or b;
    layer3_outputs(367) <= not (a and b);
    layer3_outputs(368) <= not (a or b);
    layer3_outputs(369) <= a xor b;
    layer3_outputs(370) <= a;
    layer3_outputs(371) <= a and not b;
    layer3_outputs(372) <= a and not b;
    layer3_outputs(373) <= not b or a;
    layer3_outputs(374) <= not b;
    layer3_outputs(375) <= not b;
    layer3_outputs(376) <= not (a xor b);
    layer3_outputs(377) <= not a or b;
    layer3_outputs(378) <= not b;
    layer3_outputs(379) <= not a or b;
    layer3_outputs(380) <= not a or b;
    layer3_outputs(381) <= a and not b;
    layer3_outputs(382) <= not (a or b);
    layer3_outputs(383) <= not (a or b);
    layer3_outputs(384) <= not (a xor b);
    layer3_outputs(385) <= a and not b;
    layer3_outputs(386) <= not (a xor b);
    layer3_outputs(387) <= not (a and b);
    layer3_outputs(388) <= not (a and b);
    layer3_outputs(389) <= not b;
    layer3_outputs(390) <= a;
    layer3_outputs(391) <= 1'b0;
    layer3_outputs(392) <= not (a and b);
    layer3_outputs(393) <= a and b;
    layer3_outputs(394) <= not (a and b);
    layer3_outputs(395) <= not b or a;
    layer3_outputs(396) <= a;
    layer3_outputs(397) <= b and not a;
    layer3_outputs(398) <= 1'b1;
    layer3_outputs(399) <= not (a and b);
    layer3_outputs(400) <= a;
    layer3_outputs(401) <= 1'b1;
    layer3_outputs(402) <= a and not b;
    layer3_outputs(403) <= a and not b;
    layer3_outputs(404) <= b and not a;
    layer3_outputs(405) <= not a or b;
    layer3_outputs(406) <= not (a xor b);
    layer3_outputs(407) <= not b;
    layer3_outputs(408) <= not b;
    layer3_outputs(409) <= not (a or b);
    layer3_outputs(410) <= 1'b1;
    layer3_outputs(411) <= not b;
    layer3_outputs(412) <= not a or b;
    layer3_outputs(413) <= not (a and b);
    layer3_outputs(414) <= a and b;
    layer3_outputs(415) <= not a or b;
    layer3_outputs(416) <= a and b;
    layer3_outputs(417) <= not a or b;
    layer3_outputs(418) <= not (a and b);
    layer3_outputs(419) <= 1'b1;
    layer3_outputs(420) <= b;
    layer3_outputs(421) <= a;
    layer3_outputs(422) <= b;
    layer3_outputs(423) <= a or b;
    layer3_outputs(424) <= a or b;
    layer3_outputs(425) <= b;
    layer3_outputs(426) <= b and not a;
    layer3_outputs(427) <= not a or b;
    layer3_outputs(428) <= 1'b1;
    layer3_outputs(429) <= not a;
    layer3_outputs(430) <= a and not b;
    layer3_outputs(431) <= 1'b0;
    layer3_outputs(432) <= not (a and b);
    layer3_outputs(433) <= a and b;
    layer3_outputs(434) <= not a or b;
    layer3_outputs(435) <= b;
    layer3_outputs(436) <= not a;
    layer3_outputs(437) <= not b;
    layer3_outputs(438) <= b and not a;
    layer3_outputs(439) <= not a;
    layer3_outputs(440) <= a xor b;
    layer3_outputs(441) <= b and not a;
    layer3_outputs(442) <= not (a and b);
    layer3_outputs(443) <= a;
    layer3_outputs(444) <= not a or b;
    layer3_outputs(445) <= b;
    layer3_outputs(446) <= not (a and b);
    layer3_outputs(447) <= 1'b1;
    layer3_outputs(448) <= not (a or b);
    layer3_outputs(449) <= 1'b1;
    layer3_outputs(450) <= a xor b;
    layer3_outputs(451) <= b and not a;
    layer3_outputs(452) <= b and not a;
    layer3_outputs(453) <= not (a or b);
    layer3_outputs(454) <= a and b;
    layer3_outputs(455) <= a and not b;
    layer3_outputs(456) <= not a;
    layer3_outputs(457) <= b;
    layer3_outputs(458) <= not a or b;
    layer3_outputs(459) <= b and not a;
    layer3_outputs(460) <= not (a and b);
    layer3_outputs(461) <= a or b;
    layer3_outputs(462) <= 1'b1;
    layer3_outputs(463) <= b;
    layer3_outputs(464) <= 1'b1;
    layer3_outputs(465) <= a or b;
    layer3_outputs(466) <= not b;
    layer3_outputs(467) <= 1'b1;
    layer3_outputs(468) <= 1'b1;
    layer3_outputs(469) <= a and b;
    layer3_outputs(470) <= not (a and b);
    layer3_outputs(471) <= a or b;
    layer3_outputs(472) <= not (a xor b);
    layer3_outputs(473) <= not a or b;
    layer3_outputs(474) <= 1'b1;
    layer3_outputs(475) <= b and not a;
    layer3_outputs(476) <= not (a or b);
    layer3_outputs(477) <= a and b;
    layer3_outputs(478) <= a;
    layer3_outputs(479) <= a and not b;
    layer3_outputs(480) <= not a;
    layer3_outputs(481) <= 1'b0;
    layer3_outputs(482) <= b;
    layer3_outputs(483) <= not (a and b);
    layer3_outputs(484) <= not (a xor b);
    layer3_outputs(485) <= a and b;
    layer3_outputs(486) <= b;
    layer3_outputs(487) <= 1'b0;
    layer3_outputs(488) <= not b or a;
    layer3_outputs(489) <= b;
    layer3_outputs(490) <= not a or b;
    layer3_outputs(491) <= a and b;
    layer3_outputs(492) <= not b or a;
    layer3_outputs(493) <= b;
    layer3_outputs(494) <= 1'b1;
    layer3_outputs(495) <= not a or b;
    layer3_outputs(496) <= a and not b;
    layer3_outputs(497) <= not b or a;
    layer3_outputs(498) <= not a;
    layer3_outputs(499) <= not (a and b);
    layer3_outputs(500) <= a;
    layer3_outputs(501) <= not a;
    layer3_outputs(502) <= not b or a;
    layer3_outputs(503) <= a;
    layer3_outputs(504) <= a and b;
    layer3_outputs(505) <= not a or b;
    layer3_outputs(506) <= b;
    layer3_outputs(507) <= a or b;
    layer3_outputs(508) <= a or b;
    layer3_outputs(509) <= b and not a;
    layer3_outputs(510) <= not a or b;
    layer3_outputs(511) <= not (a and b);
    layer3_outputs(512) <= a and not b;
    layer3_outputs(513) <= 1'b0;
    layer3_outputs(514) <= a and b;
    layer3_outputs(515) <= not b or a;
    layer3_outputs(516) <= 1'b1;
    layer3_outputs(517) <= a or b;
    layer3_outputs(518) <= not (a and b);
    layer3_outputs(519) <= a and not b;
    layer3_outputs(520) <= not a or b;
    layer3_outputs(521) <= not b;
    layer3_outputs(522) <= a;
    layer3_outputs(523) <= b;
    layer3_outputs(524) <= not b;
    layer3_outputs(525) <= b;
    layer3_outputs(526) <= 1'b1;
    layer3_outputs(527) <= b and not a;
    layer3_outputs(528) <= not a or b;
    layer3_outputs(529) <= 1'b1;
    layer3_outputs(530) <= not a or b;
    layer3_outputs(531) <= b;
    layer3_outputs(532) <= 1'b0;
    layer3_outputs(533) <= not (a or b);
    layer3_outputs(534) <= b;
    layer3_outputs(535) <= not (a or b);
    layer3_outputs(536) <= a or b;
    layer3_outputs(537) <= a xor b;
    layer3_outputs(538) <= a and not b;
    layer3_outputs(539) <= a;
    layer3_outputs(540) <= 1'b1;
    layer3_outputs(541) <= a and not b;
    layer3_outputs(542) <= not b or a;
    layer3_outputs(543) <= 1'b0;
    layer3_outputs(544) <= a;
    layer3_outputs(545) <= a and not b;
    layer3_outputs(546) <= 1'b1;
    layer3_outputs(547) <= not b;
    layer3_outputs(548) <= not (a or b);
    layer3_outputs(549) <= a;
    layer3_outputs(550) <= not b or a;
    layer3_outputs(551) <= not a or b;
    layer3_outputs(552) <= not b or a;
    layer3_outputs(553) <= 1'b1;
    layer3_outputs(554) <= not b;
    layer3_outputs(555) <= not a;
    layer3_outputs(556) <= not b;
    layer3_outputs(557) <= b;
    layer3_outputs(558) <= not a or b;
    layer3_outputs(559) <= b and not a;
    layer3_outputs(560) <= 1'b1;
    layer3_outputs(561) <= 1'b1;
    layer3_outputs(562) <= not (a xor b);
    layer3_outputs(563) <= 1'b0;
    layer3_outputs(564) <= b and not a;
    layer3_outputs(565) <= a and b;
    layer3_outputs(566) <= not (a or b);
    layer3_outputs(567) <= a;
    layer3_outputs(568) <= not a;
    layer3_outputs(569) <= a or b;
    layer3_outputs(570) <= 1'b1;
    layer3_outputs(571) <= a and not b;
    layer3_outputs(572) <= 1'b1;
    layer3_outputs(573) <= a or b;
    layer3_outputs(574) <= not a or b;
    layer3_outputs(575) <= a and b;
    layer3_outputs(576) <= b and not a;
    layer3_outputs(577) <= not b or a;
    layer3_outputs(578) <= b and not a;
    layer3_outputs(579) <= b;
    layer3_outputs(580) <= b and not a;
    layer3_outputs(581) <= b and not a;
    layer3_outputs(582) <= not (a or b);
    layer3_outputs(583) <= a or b;
    layer3_outputs(584) <= not b;
    layer3_outputs(585) <= a or b;
    layer3_outputs(586) <= b and not a;
    layer3_outputs(587) <= not a or b;
    layer3_outputs(588) <= 1'b0;
    layer3_outputs(589) <= a or b;
    layer3_outputs(590) <= not b or a;
    layer3_outputs(591) <= not a;
    layer3_outputs(592) <= not (a and b);
    layer3_outputs(593) <= 1'b1;
    layer3_outputs(594) <= not b or a;
    layer3_outputs(595) <= a and b;
    layer3_outputs(596) <= b;
    layer3_outputs(597) <= not a;
    layer3_outputs(598) <= not a or b;
    layer3_outputs(599) <= a and b;
    layer3_outputs(600) <= 1'b1;
    layer3_outputs(601) <= a and b;
    layer3_outputs(602) <= not a;
    layer3_outputs(603) <= not a or b;
    layer3_outputs(604) <= a and not b;
    layer3_outputs(605) <= not b;
    layer3_outputs(606) <= not (a and b);
    layer3_outputs(607) <= b and not a;
    layer3_outputs(608) <= not (a and b);
    layer3_outputs(609) <= not a or b;
    layer3_outputs(610) <= not a or b;
    layer3_outputs(611) <= b and not a;
    layer3_outputs(612) <= b and not a;
    layer3_outputs(613) <= 1'b1;
    layer3_outputs(614) <= 1'b0;
    layer3_outputs(615) <= not a;
    layer3_outputs(616) <= a or b;
    layer3_outputs(617) <= not a or b;
    layer3_outputs(618) <= a and not b;
    layer3_outputs(619) <= not (a or b);
    layer3_outputs(620) <= a;
    layer3_outputs(621) <= a and not b;
    layer3_outputs(622) <= b;
    layer3_outputs(623) <= not a;
    layer3_outputs(624) <= not (a and b);
    layer3_outputs(625) <= b;
    layer3_outputs(626) <= 1'b0;
    layer3_outputs(627) <= a or b;
    layer3_outputs(628) <= not (a and b);
    layer3_outputs(629) <= not (a or b);
    layer3_outputs(630) <= 1'b0;
    layer3_outputs(631) <= a and not b;
    layer3_outputs(632) <= 1'b1;
    layer3_outputs(633) <= not (a xor b);
    layer3_outputs(634) <= 1'b0;
    layer3_outputs(635) <= b;
    layer3_outputs(636) <= 1'b0;
    layer3_outputs(637) <= not a;
    layer3_outputs(638) <= b and not a;
    layer3_outputs(639) <= b;
    layer3_outputs(640) <= a and b;
    layer3_outputs(641) <= b and not a;
    layer3_outputs(642) <= not a or b;
    layer3_outputs(643) <= a or b;
    layer3_outputs(644) <= a;
    layer3_outputs(645) <= a and b;
    layer3_outputs(646) <= b and not a;
    layer3_outputs(647) <= 1'b0;
    layer3_outputs(648) <= not b;
    layer3_outputs(649) <= 1'b1;
    layer3_outputs(650) <= a and not b;
    layer3_outputs(651) <= b and not a;
    layer3_outputs(652) <= 1'b0;
    layer3_outputs(653) <= not a;
    layer3_outputs(654) <= 1'b1;
    layer3_outputs(655) <= not (a or b);
    layer3_outputs(656) <= a or b;
    layer3_outputs(657) <= not a;
    layer3_outputs(658) <= 1'b0;
    layer3_outputs(659) <= a;
    layer3_outputs(660) <= 1'b0;
    layer3_outputs(661) <= a or b;
    layer3_outputs(662) <= 1'b1;
    layer3_outputs(663) <= not a;
    layer3_outputs(664) <= not (a and b);
    layer3_outputs(665) <= a or b;
    layer3_outputs(666) <= b;
    layer3_outputs(667) <= a and b;
    layer3_outputs(668) <= not b or a;
    layer3_outputs(669) <= a and not b;
    layer3_outputs(670) <= b;
    layer3_outputs(671) <= 1'b1;
    layer3_outputs(672) <= not (a and b);
    layer3_outputs(673) <= a and not b;
    layer3_outputs(674) <= not (a and b);
    layer3_outputs(675) <= 1'b0;
    layer3_outputs(676) <= b and not a;
    layer3_outputs(677) <= a xor b;
    layer3_outputs(678) <= not b;
    layer3_outputs(679) <= not b or a;
    layer3_outputs(680) <= not b or a;
    layer3_outputs(681) <= not (a and b);
    layer3_outputs(682) <= not (a xor b);
    layer3_outputs(683) <= 1'b0;
    layer3_outputs(684) <= a and not b;
    layer3_outputs(685) <= not (a and b);
    layer3_outputs(686) <= a and not b;
    layer3_outputs(687) <= not a;
    layer3_outputs(688) <= not b or a;
    layer3_outputs(689) <= 1'b1;
    layer3_outputs(690) <= not b or a;
    layer3_outputs(691) <= a;
    layer3_outputs(692) <= a and b;
    layer3_outputs(693) <= a;
    layer3_outputs(694) <= not (a and b);
    layer3_outputs(695) <= a;
    layer3_outputs(696) <= 1'b1;
    layer3_outputs(697) <= not a or b;
    layer3_outputs(698) <= not (a or b);
    layer3_outputs(699) <= not (a or b);
    layer3_outputs(700) <= not b or a;
    layer3_outputs(701) <= a and not b;
    layer3_outputs(702) <= a and not b;
    layer3_outputs(703) <= 1'b1;
    layer3_outputs(704) <= b and not a;
    layer3_outputs(705) <= b and not a;
    layer3_outputs(706) <= not (a and b);
    layer3_outputs(707) <= not (a and b);
    layer3_outputs(708) <= a and b;
    layer3_outputs(709) <= not a or b;
    layer3_outputs(710) <= 1'b1;
    layer3_outputs(711) <= a and b;
    layer3_outputs(712) <= not (a and b);
    layer3_outputs(713) <= a or b;
    layer3_outputs(714) <= b and not a;
    layer3_outputs(715) <= a and not b;
    layer3_outputs(716) <= not (a and b);
    layer3_outputs(717) <= not a;
    layer3_outputs(718) <= not a;
    layer3_outputs(719) <= a and b;
    layer3_outputs(720) <= b and not a;
    layer3_outputs(721) <= b;
    layer3_outputs(722) <= 1'b0;
    layer3_outputs(723) <= not a;
    layer3_outputs(724) <= a and b;
    layer3_outputs(725) <= not b or a;
    layer3_outputs(726) <= not (a or b);
    layer3_outputs(727) <= not b;
    layer3_outputs(728) <= a and b;
    layer3_outputs(729) <= not (a and b);
    layer3_outputs(730) <= not (a and b);
    layer3_outputs(731) <= b;
    layer3_outputs(732) <= b;
    layer3_outputs(733) <= a;
    layer3_outputs(734) <= 1'b1;
    layer3_outputs(735) <= a or b;
    layer3_outputs(736) <= b and not a;
    layer3_outputs(737) <= not (a and b);
    layer3_outputs(738) <= b;
    layer3_outputs(739) <= not b or a;
    layer3_outputs(740) <= not (a or b);
    layer3_outputs(741) <= a;
    layer3_outputs(742) <= not b or a;
    layer3_outputs(743) <= a;
    layer3_outputs(744) <= not (a xor b);
    layer3_outputs(745) <= not (a or b);
    layer3_outputs(746) <= not a;
    layer3_outputs(747) <= not b or a;
    layer3_outputs(748) <= not a;
    layer3_outputs(749) <= a;
    layer3_outputs(750) <= a;
    layer3_outputs(751) <= a;
    layer3_outputs(752) <= not (a or b);
    layer3_outputs(753) <= not a or b;
    layer3_outputs(754) <= 1'b1;
    layer3_outputs(755) <= a or b;
    layer3_outputs(756) <= not (a and b);
    layer3_outputs(757) <= not (a and b);
    layer3_outputs(758) <= 1'b0;
    layer3_outputs(759) <= not (a and b);
    layer3_outputs(760) <= b;
    layer3_outputs(761) <= 1'b1;
    layer3_outputs(762) <= a;
    layer3_outputs(763) <= b;
    layer3_outputs(764) <= 1'b1;
    layer3_outputs(765) <= a and not b;
    layer3_outputs(766) <= not b or a;
    layer3_outputs(767) <= a and not b;
    layer3_outputs(768) <= not a or b;
    layer3_outputs(769) <= 1'b0;
    layer3_outputs(770) <= not a or b;
    layer3_outputs(771) <= b;
    layer3_outputs(772) <= a;
    layer3_outputs(773) <= b;
    layer3_outputs(774) <= b;
    layer3_outputs(775) <= 1'b0;
    layer3_outputs(776) <= not b or a;
    layer3_outputs(777) <= not b or a;
    layer3_outputs(778) <= 1'b0;
    layer3_outputs(779) <= b and not a;
    layer3_outputs(780) <= a;
    layer3_outputs(781) <= not (a and b);
    layer3_outputs(782) <= not b;
    layer3_outputs(783) <= a;
    layer3_outputs(784) <= not (a or b);
    layer3_outputs(785) <= 1'b0;
    layer3_outputs(786) <= a and b;
    layer3_outputs(787) <= not (a or b);
    layer3_outputs(788) <= not b;
    layer3_outputs(789) <= a and not b;
    layer3_outputs(790) <= b and not a;
    layer3_outputs(791) <= 1'b1;
    layer3_outputs(792) <= a;
    layer3_outputs(793) <= not b;
    layer3_outputs(794) <= not (a and b);
    layer3_outputs(795) <= a;
    layer3_outputs(796) <= not (a and b);
    layer3_outputs(797) <= a or b;
    layer3_outputs(798) <= 1'b1;
    layer3_outputs(799) <= a or b;
    layer3_outputs(800) <= b and not a;
    layer3_outputs(801) <= not b;
    layer3_outputs(802) <= a and not b;
    layer3_outputs(803) <= b and not a;
    layer3_outputs(804) <= a xor b;
    layer3_outputs(805) <= a;
    layer3_outputs(806) <= 1'b0;
    layer3_outputs(807) <= b and not a;
    layer3_outputs(808) <= a or b;
    layer3_outputs(809) <= a and not b;
    layer3_outputs(810) <= a;
    layer3_outputs(811) <= a;
    layer3_outputs(812) <= not (a or b);
    layer3_outputs(813) <= a;
    layer3_outputs(814) <= a;
    layer3_outputs(815) <= not a or b;
    layer3_outputs(816) <= a xor b;
    layer3_outputs(817) <= not b or a;
    layer3_outputs(818) <= a;
    layer3_outputs(819) <= a and not b;
    layer3_outputs(820) <= not (a and b);
    layer3_outputs(821) <= not a or b;
    layer3_outputs(822) <= b and not a;
    layer3_outputs(823) <= a and not b;
    layer3_outputs(824) <= not a;
    layer3_outputs(825) <= a or b;
    layer3_outputs(826) <= a and b;
    layer3_outputs(827) <= not b or a;
    layer3_outputs(828) <= 1'b0;
    layer3_outputs(829) <= a and b;
    layer3_outputs(830) <= not (a or b);
    layer3_outputs(831) <= b and not a;
    layer3_outputs(832) <= a and not b;
    layer3_outputs(833) <= a or b;
    layer3_outputs(834) <= not a or b;
    layer3_outputs(835) <= 1'b1;
    layer3_outputs(836) <= a;
    layer3_outputs(837) <= a and not b;
    layer3_outputs(838) <= not (a or b);
    layer3_outputs(839) <= a and b;
    layer3_outputs(840) <= b and not a;
    layer3_outputs(841) <= b and not a;
    layer3_outputs(842) <= a and not b;
    layer3_outputs(843) <= not a or b;
    layer3_outputs(844) <= b;
    layer3_outputs(845) <= b and not a;
    layer3_outputs(846) <= not (a or b);
    layer3_outputs(847) <= not (a or b);
    layer3_outputs(848) <= not a;
    layer3_outputs(849) <= a and not b;
    layer3_outputs(850) <= b;
    layer3_outputs(851) <= a and not b;
    layer3_outputs(852) <= b and not a;
    layer3_outputs(853) <= not b or a;
    layer3_outputs(854) <= not (a and b);
    layer3_outputs(855) <= a and b;
    layer3_outputs(856) <= a xor b;
    layer3_outputs(857) <= 1'b0;
    layer3_outputs(858) <= b and not a;
    layer3_outputs(859) <= not (a or b);
    layer3_outputs(860) <= not a;
    layer3_outputs(861) <= not (a or b);
    layer3_outputs(862) <= 1'b1;
    layer3_outputs(863) <= not a;
    layer3_outputs(864) <= a or b;
    layer3_outputs(865) <= not a;
    layer3_outputs(866) <= not (a and b);
    layer3_outputs(867) <= 1'b0;
    layer3_outputs(868) <= 1'b1;
    layer3_outputs(869) <= a and not b;
    layer3_outputs(870) <= a or b;
    layer3_outputs(871) <= not (a and b);
    layer3_outputs(872) <= not (a or b);
    layer3_outputs(873) <= b and not a;
    layer3_outputs(874) <= not a;
    layer3_outputs(875) <= a and not b;
    layer3_outputs(876) <= 1'b0;
    layer3_outputs(877) <= 1'b1;
    layer3_outputs(878) <= not a;
    layer3_outputs(879) <= a;
    layer3_outputs(880) <= not b or a;
    layer3_outputs(881) <= not a;
    layer3_outputs(882) <= a and b;
    layer3_outputs(883) <= a;
    layer3_outputs(884) <= a and b;
    layer3_outputs(885) <= a xor b;
    layer3_outputs(886) <= 1'b1;
    layer3_outputs(887) <= a and b;
    layer3_outputs(888) <= not a or b;
    layer3_outputs(889) <= b and not a;
    layer3_outputs(890) <= a;
    layer3_outputs(891) <= not a;
    layer3_outputs(892) <= not (a and b);
    layer3_outputs(893) <= a and not b;
    layer3_outputs(894) <= not (a or b);
    layer3_outputs(895) <= 1'b0;
    layer3_outputs(896) <= not b or a;
    layer3_outputs(897) <= a or b;
    layer3_outputs(898) <= not b;
    layer3_outputs(899) <= not (a and b);
    layer3_outputs(900) <= a;
    layer3_outputs(901) <= not a or b;
    layer3_outputs(902) <= a and b;
    layer3_outputs(903) <= 1'b1;
    layer3_outputs(904) <= a;
    layer3_outputs(905) <= not (a and b);
    layer3_outputs(906) <= not a or b;
    layer3_outputs(907) <= 1'b1;
    layer3_outputs(908) <= a or b;
    layer3_outputs(909) <= not a or b;
    layer3_outputs(910) <= a;
    layer3_outputs(911) <= 1'b1;
    layer3_outputs(912) <= not b;
    layer3_outputs(913) <= not (a and b);
    layer3_outputs(914) <= a and b;
    layer3_outputs(915) <= not b or a;
    layer3_outputs(916) <= a and b;
    layer3_outputs(917) <= b;
    layer3_outputs(918) <= a;
    layer3_outputs(919) <= b and not a;
    layer3_outputs(920) <= 1'b0;
    layer3_outputs(921) <= b;
    layer3_outputs(922) <= b and not a;
    layer3_outputs(923) <= not b or a;
    layer3_outputs(924) <= not (a and b);
    layer3_outputs(925) <= a or b;
    layer3_outputs(926) <= 1'b1;
    layer3_outputs(927) <= a or b;
    layer3_outputs(928) <= a and b;
    layer3_outputs(929) <= b and not a;
    layer3_outputs(930) <= not b or a;
    layer3_outputs(931) <= a and b;
    layer3_outputs(932) <= not (a or b);
    layer3_outputs(933) <= 1'b1;
    layer3_outputs(934) <= 1'b1;
    layer3_outputs(935) <= a and not b;
    layer3_outputs(936) <= a;
    layer3_outputs(937) <= a or b;
    layer3_outputs(938) <= b;
    layer3_outputs(939) <= not a;
    layer3_outputs(940) <= b and not a;
    layer3_outputs(941) <= a and not b;
    layer3_outputs(942) <= not a;
    layer3_outputs(943) <= not b or a;
    layer3_outputs(944) <= b and not a;
    layer3_outputs(945) <= not (a or b);
    layer3_outputs(946) <= not (a and b);
    layer3_outputs(947) <= 1'b0;
    layer3_outputs(948) <= b and not a;
    layer3_outputs(949) <= a or b;
    layer3_outputs(950) <= 1'b1;
    layer3_outputs(951) <= not (a xor b);
    layer3_outputs(952) <= not (a or b);
    layer3_outputs(953) <= a and not b;
    layer3_outputs(954) <= not b or a;
    layer3_outputs(955) <= a or b;
    layer3_outputs(956) <= b and not a;
    layer3_outputs(957) <= b and not a;
    layer3_outputs(958) <= 1'b1;
    layer3_outputs(959) <= 1'b1;
    layer3_outputs(960) <= not a or b;
    layer3_outputs(961) <= not a;
    layer3_outputs(962) <= a or b;
    layer3_outputs(963) <= a or b;
    layer3_outputs(964) <= a and b;
    layer3_outputs(965) <= a or b;
    layer3_outputs(966) <= 1'b0;
    layer3_outputs(967) <= not (a and b);
    layer3_outputs(968) <= 1'b0;
    layer3_outputs(969) <= a;
    layer3_outputs(970) <= not b;
    layer3_outputs(971) <= not (a or b);
    layer3_outputs(972) <= b;
    layer3_outputs(973) <= a and b;
    layer3_outputs(974) <= 1'b1;
    layer3_outputs(975) <= not b or a;
    layer3_outputs(976) <= not (a or b);
    layer3_outputs(977) <= 1'b1;
    layer3_outputs(978) <= not (a and b);
    layer3_outputs(979) <= not a or b;
    layer3_outputs(980) <= not b or a;
    layer3_outputs(981) <= 1'b0;
    layer3_outputs(982) <= b;
    layer3_outputs(983) <= a and b;
    layer3_outputs(984) <= not (a or b);
    layer3_outputs(985) <= not b or a;
    layer3_outputs(986) <= a and b;
    layer3_outputs(987) <= a;
    layer3_outputs(988) <= not (a and b);
    layer3_outputs(989) <= a or b;
    layer3_outputs(990) <= a and b;
    layer3_outputs(991) <= a or b;
    layer3_outputs(992) <= b;
    layer3_outputs(993) <= not (a or b);
    layer3_outputs(994) <= 1'b0;
    layer3_outputs(995) <= 1'b0;
    layer3_outputs(996) <= not a or b;
    layer3_outputs(997) <= not a or b;
    layer3_outputs(998) <= not b or a;
    layer3_outputs(999) <= not (a and b);
    layer3_outputs(1000) <= not a;
    layer3_outputs(1001) <= not (a or b);
    layer3_outputs(1002) <= not (a xor b);
    layer3_outputs(1003) <= not (a or b);
    layer3_outputs(1004) <= a xor b;
    layer3_outputs(1005) <= b and not a;
    layer3_outputs(1006) <= a and b;
    layer3_outputs(1007) <= not b or a;
    layer3_outputs(1008) <= not (a or b);
    layer3_outputs(1009) <= not b or a;
    layer3_outputs(1010) <= a;
    layer3_outputs(1011) <= not (a or b);
    layer3_outputs(1012) <= 1'b1;
    layer3_outputs(1013) <= 1'b0;
    layer3_outputs(1014) <= not (a and b);
    layer3_outputs(1015) <= not a or b;
    layer3_outputs(1016) <= b;
    layer3_outputs(1017) <= not (a or b);
    layer3_outputs(1018) <= b and not a;
    layer3_outputs(1019) <= b and not a;
    layer3_outputs(1020) <= not a or b;
    layer3_outputs(1021) <= not b or a;
    layer3_outputs(1022) <= not b or a;
    layer3_outputs(1023) <= not a;
    layer3_outputs(1024) <= b;
    layer3_outputs(1025) <= a;
    layer3_outputs(1026) <= 1'b1;
    layer3_outputs(1027) <= not a;
    layer3_outputs(1028) <= 1'b0;
    layer3_outputs(1029) <= not b;
    layer3_outputs(1030) <= a or b;
    layer3_outputs(1031) <= b and not a;
    layer3_outputs(1032) <= a;
    layer3_outputs(1033) <= a xor b;
    layer3_outputs(1034) <= not b;
    layer3_outputs(1035) <= not a;
    layer3_outputs(1036) <= a and b;
    layer3_outputs(1037) <= not a;
    layer3_outputs(1038) <= 1'b1;
    layer3_outputs(1039) <= not a;
    layer3_outputs(1040) <= not a;
    layer3_outputs(1041) <= not a or b;
    layer3_outputs(1042) <= a and b;
    layer3_outputs(1043) <= not (a or b);
    layer3_outputs(1044) <= a;
    layer3_outputs(1045) <= a or b;
    layer3_outputs(1046) <= a and not b;
    layer3_outputs(1047) <= a and not b;
    layer3_outputs(1048) <= not a or b;
    layer3_outputs(1049) <= a and not b;
    layer3_outputs(1050) <= a;
    layer3_outputs(1051) <= not b or a;
    layer3_outputs(1052) <= not (a and b);
    layer3_outputs(1053) <= not a or b;
    layer3_outputs(1054) <= not b;
    layer3_outputs(1055) <= not a;
    layer3_outputs(1056) <= not (a and b);
    layer3_outputs(1057) <= not a or b;
    layer3_outputs(1058) <= b and not a;
    layer3_outputs(1059) <= 1'b0;
    layer3_outputs(1060) <= b and not a;
    layer3_outputs(1061) <= a xor b;
    layer3_outputs(1062) <= a and not b;
    layer3_outputs(1063) <= a;
    layer3_outputs(1064) <= not b;
    layer3_outputs(1065) <= not (a or b);
    layer3_outputs(1066) <= b and not a;
    layer3_outputs(1067) <= a;
    layer3_outputs(1068) <= a and b;
    layer3_outputs(1069) <= a;
    layer3_outputs(1070) <= not (a or b);
    layer3_outputs(1071) <= a xor b;
    layer3_outputs(1072) <= b and not a;
    layer3_outputs(1073) <= b and not a;
    layer3_outputs(1074) <= a;
    layer3_outputs(1075) <= a and b;
    layer3_outputs(1076) <= not a;
    layer3_outputs(1077) <= a and not b;
    layer3_outputs(1078) <= a;
    layer3_outputs(1079) <= b;
    layer3_outputs(1080) <= 1'b0;
    layer3_outputs(1081) <= a;
    layer3_outputs(1082) <= not b or a;
    layer3_outputs(1083) <= 1'b1;
    layer3_outputs(1084) <= b and not a;
    layer3_outputs(1085) <= 1'b1;
    layer3_outputs(1086) <= not (a and b);
    layer3_outputs(1087) <= a and b;
    layer3_outputs(1088) <= not (a or b);
    layer3_outputs(1089) <= a;
    layer3_outputs(1090) <= not a;
    layer3_outputs(1091) <= a or b;
    layer3_outputs(1092) <= not (a and b);
    layer3_outputs(1093) <= not b or a;
    layer3_outputs(1094) <= a and not b;
    layer3_outputs(1095) <= not (a and b);
    layer3_outputs(1096) <= not b;
    layer3_outputs(1097) <= not b;
    layer3_outputs(1098) <= 1'b1;
    layer3_outputs(1099) <= not b or a;
    layer3_outputs(1100) <= b;
    layer3_outputs(1101) <= 1'b1;
    layer3_outputs(1102) <= not (a and b);
    layer3_outputs(1103) <= not (a or b);
    layer3_outputs(1104) <= a and not b;
    layer3_outputs(1105) <= 1'b0;
    layer3_outputs(1106) <= b;
    layer3_outputs(1107) <= 1'b0;
    layer3_outputs(1108) <= not (a and b);
    layer3_outputs(1109) <= 1'b0;
    layer3_outputs(1110) <= not b;
    layer3_outputs(1111) <= 1'b1;
    layer3_outputs(1112) <= not b;
    layer3_outputs(1113) <= 1'b1;
    layer3_outputs(1114) <= not (a and b);
    layer3_outputs(1115) <= not a or b;
    layer3_outputs(1116) <= 1'b0;
    layer3_outputs(1117) <= not (a or b);
    layer3_outputs(1118) <= a and b;
    layer3_outputs(1119) <= b and not a;
    layer3_outputs(1120) <= a and not b;
    layer3_outputs(1121) <= a and b;
    layer3_outputs(1122) <= not a or b;
    layer3_outputs(1123) <= b and not a;
    layer3_outputs(1124) <= not a or b;
    layer3_outputs(1125) <= not a;
    layer3_outputs(1126) <= a;
    layer3_outputs(1127) <= not a or b;
    layer3_outputs(1128) <= 1'b0;
    layer3_outputs(1129) <= a and not b;
    layer3_outputs(1130) <= not a;
    layer3_outputs(1131) <= a or b;
    layer3_outputs(1132) <= not b or a;
    layer3_outputs(1133) <= not (a or b);
    layer3_outputs(1134) <= not a;
    layer3_outputs(1135) <= not b or a;
    layer3_outputs(1136) <= b;
    layer3_outputs(1137) <= a and b;
    layer3_outputs(1138) <= not (a and b);
    layer3_outputs(1139) <= a and not b;
    layer3_outputs(1140) <= a or b;
    layer3_outputs(1141) <= not b or a;
    layer3_outputs(1142) <= a;
    layer3_outputs(1143) <= a and b;
    layer3_outputs(1144) <= not b;
    layer3_outputs(1145) <= 1'b1;
    layer3_outputs(1146) <= not (a and b);
    layer3_outputs(1147) <= a or b;
    layer3_outputs(1148) <= not b or a;
    layer3_outputs(1149) <= b and not a;
    layer3_outputs(1150) <= a and not b;
    layer3_outputs(1151) <= a and b;
    layer3_outputs(1152) <= 1'b1;
    layer3_outputs(1153) <= b and not a;
    layer3_outputs(1154) <= not (a and b);
    layer3_outputs(1155) <= a and b;
    layer3_outputs(1156) <= a;
    layer3_outputs(1157) <= a and not b;
    layer3_outputs(1158) <= a and not b;
    layer3_outputs(1159) <= 1'b0;
    layer3_outputs(1160) <= a and not b;
    layer3_outputs(1161) <= a;
    layer3_outputs(1162) <= b;
    layer3_outputs(1163) <= not (a xor b);
    layer3_outputs(1164) <= not a;
    layer3_outputs(1165) <= not b or a;
    layer3_outputs(1166) <= 1'b0;
    layer3_outputs(1167) <= a or b;
    layer3_outputs(1168) <= not (a or b);
    layer3_outputs(1169) <= not b or a;
    layer3_outputs(1170) <= a;
    layer3_outputs(1171) <= not b;
    layer3_outputs(1172) <= not a or b;
    layer3_outputs(1173) <= a;
    layer3_outputs(1174) <= a;
    layer3_outputs(1175) <= 1'b1;
    layer3_outputs(1176) <= not b or a;
    layer3_outputs(1177) <= not b or a;
    layer3_outputs(1178) <= 1'b0;
    layer3_outputs(1179) <= 1'b0;
    layer3_outputs(1180) <= a and b;
    layer3_outputs(1181) <= not b;
    layer3_outputs(1182) <= a;
    layer3_outputs(1183) <= not a or b;
    layer3_outputs(1184) <= not b or a;
    layer3_outputs(1185) <= a and b;
    layer3_outputs(1186) <= not a;
    layer3_outputs(1187) <= 1'b0;
    layer3_outputs(1188) <= not b or a;
    layer3_outputs(1189) <= not b or a;
    layer3_outputs(1190) <= not (a or b);
    layer3_outputs(1191) <= a;
    layer3_outputs(1192) <= a;
    layer3_outputs(1193) <= 1'b0;
    layer3_outputs(1194) <= not a or b;
    layer3_outputs(1195) <= b and not a;
    layer3_outputs(1196) <= 1'b0;
    layer3_outputs(1197) <= a and not b;
    layer3_outputs(1198) <= 1'b1;
    layer3_outputs(1199) <= 1'b0;
    layer3_outputs(1200) <= a;
    layer3_outputs(1201) <= 1'b0;
    layer3_outputs(1202) <= b and not a;
    layer3_outputs(1203) <= b and not a;
    layer3_outputs(1204) <= 1'b1;
    layer3_outputs(1205) <= b;
    layer3_outputs(1206) <= a and b;
    layer3_outputs(1207) <= not b;
    layer3_outputs(1208) <= not (a or b);
    layer3_outputs(1209) <= b and not a;
    layer3_outputs(1210) <= a and not b;
    layer3_outputs(1211) <= not (a and b);
    layer3_outputs(1212) <= not a;
    layer3_outputs(1213) <= a or b;
    layer3_outputs(1214) <= not (a and b);
    layer3_outputs(1215) <= a and not b;
    layer3_outputs(1216) <= a and b;
    layer3_outputs(1217) <= not (a and b);
    layer3_outputs(1218) <= 1'b0;
    layer3_outputs(1219) <= not b or a;
    layer3_outputs(1220) <= 1'b1;
    layer3_outputs(1221) <= 1'b0;
    layer3_outputs(1222) <= a xor b;
    layer3_outputs(1223) <= not b;
    layer3_outputs(1224) <= a;
    layer3_outputs(1225) <= not (a and b);
    layer3_outputs(1226) <= b and not a;
    layer3_outputs(1227) <= a or b;
    layer3_outputs(1228) <= b;
    layer3_outputs(1229) <= a or b;
    layer3_outputs(1230) <= not (a xor b);
    layer3_outputs(1231) <= a and not b;
    layer3_outputs(1232) <= not b;
    layer3_outputs(1233) <= a and not b;
    layer3_outputs(1234) <= not b or a;
    layer3_outputs(1235) <= not b;
    layer3_outputs(1236) <= b and not a;
    layer3_outputs(1237) <= not b;
    layer3_outputs(1238) <= not (a and b);
    layer3_outputs(1239) <= 1'b1;
    layer3_outputs(1240) <= 1'b0;
    layer3_outputs(1241) <= not a;
    layer3_outputs(1242) <= a and not b;
    layer3_outputs(1243) <= not b;
    layer3_outputs(1244) <= a xor b;
    layer3_outputs(1245) <= not a or b;
    layer3_outputs(1246) <= a or b;
    layer3_outputs(1247) <= 1'b0;
    layer3_outputs(1248) <= not b;
    layer3_outputs(1249) <= not b or a;
    layer3_outputs(1250) <= a and b;
    layer3_outputs(1251) <= not a or b;
    layer3_outputs(1252) <= a;
    layer3_outputs(1253) <= not a;
    layer3_outputs(1254) <= not b;
    layer3_outputs(1255) <= not (a or b);
    layer3_outputs(1256) <= 1'b0;
    layer3_outputs(1257) <= b;
    layer3_outputs(1258) <= a and b;
    layer3_outputs(1259) <= not (a or b);
    layer3_outputs(1260) <= not b or a;
    layer3_outputs(1261) <= a and not b;
    layer3_outputs(1262) <= b;
    layer3_outputs(1263) <= a;
    layer3_outputs(1264) <= a;
    layer3_outputs(1265) <= not a or b;
    layer3_outputs(1266) <= b and not a;
    layer3_outputs(1267) <= b;
    layer3_outputs(1268) <= 1'b0;
    layer3_outputs(1269) <= not a;
    layer3_outputs(1270) <= not (a or b);
    layer3_outputs(1271) <= not b or a;
    layer3_outputs(1272) <= not (a or b);
    layer3_outputs(1273) <= a and b;
    layer3_outputs(1274) <= b and not a;
    layer3_outputs(1275) <= 1'b1;
    layer3_outputs(1276) <= not b;
    layer3_outputs(1277) <= not b or a;
    layer3_outputs(1278) <= b and not a;
    layer3_outputs(1279) <= not (a or b);
    layer3_outputs(1280) <= 1'b1;
    layer3_outputs(1281) <= b;
    layer3_outputs(1282) <= b and not a;
    layer3_outputs(1283) <= not (a or b);
    layer3_outputs(1284) <= not a;
    layer3_outputs(1285) <= b and not a;
    layer3_outputs(1286) <= not (a xor b);
    layer3_outputs(1287) <= not (a or b);
    layer3_outputs(1288) <= 1'b0;
    layer3_outputs(1289) <= a and b;
    layer3_outputs(1290) <= 1'b0;
    layer3_outputs(1291) <= a and not b;
    layer3_outputs(1292) <= b and not a;
    layer3_outputs(1293) <= b;
    layer3_outputs(1294) <= b and not a;
    layer3_outputs(1295) <= not b;
    layer3_outputs(1296) <= a or b;
    layer3_outputs(1297) <= not (a and b);
    layer3_outputs(1298) <= not (a or b);
    layer3_outputs(1299) <= not a;
    layer3_outputs(1300) <= 1'b0;
    layer3_outputs(1301) <= not a;
    layer3_outputs(1302) <= not a;
    layer3_outputs(1303) <= b and not a;
    layer3_outputs(1304) <= not a or b;
    layer3_outputs(1305) <= b;
    layer3_outputs(1306) <= not b or a;
    layer3_outputs(1307) <= not a;
    layer3_outputs(1308) <= not b;
    layer3_outputs(1309) <= 1'b0;
    layer3_outputs(1310) <= b and not a;
    layer3_outputs(1311) <= 1'b1;
    layer3_outputs(1312) <= 1'b1;
    layer3_outputs(1313) <= not b or a;
    layer3_outputs(1314) <= not b or a;
    layer3_outputs(1315) <= a xor b;
    layer3_outputs(1316) <= a and b;
    layer3_outputs(1317) <= not b or a;
    layer3_outputs(1318) <= a and b;
    layer3_outputs(1319) <= not b;
    layer3_outputs(1320) <= 1'b1;
    layer3_outputs(1321) <= b and not a;
    layer3_outputs(1322) <= a or b;
    layer3_outputs(1323) <= not b;
    layer3_outputs(1324) <= not b or a;
    layer3_outputs(1325) <= a xor b;
    layer3_outputs(1326) <= not (a or b);
    layer3_outputs(1327) <= b;
    layer3_outputs(1328) <= not b or a;
    layer3_outputs(1329) <= a and b;
    layer3_outputs(1330) <= a;
    layer3_outputs(1331) <= a and b;
    layer3_outputs(1332) <= not (a or b);
    layer3_outputs(1333) <= a and not b;
    layer3_outputs(1334) <= a and b;
    layer3_outputs(1335) <= not (a or b);
    layer3_outputs(1336) <= not (a or b);
    layer3_outputs(1337) <= not (a and b);
    layer3_outputs(1338) <= not a;
    layer3_outputs(1339) <= b and not a;
    layer3_outputs(1340) <= not b or a;
    layer3_outputs(1341) <= a and not b;
    layer3_outputs(1342) <= a and b;
    layer3_outputs(1343) <= a xor b;
    layer3_outputs(1344) <= not b or a;
    layer3_outputs(1345) <= a and b;
    layer3_outputs(1346) <= 1'b1;
    layer3_outputs(1347) <= not (a or b);
    layer3_outputs(1348) <= a and not b;
    layer3_outputs(1349) <= b;
    layer3_outputs(1350) <= a and b;
    layer3_outputs(1351) <= not a;
    layer3_outputs(1352) <= not b;
    layer3_outputs(1353) <= not b;
    layer3_outputs(1354) <= not a;
    layer3_outputs(1355) <= not a or b;
    layer3_outputs(1356) <= 1'b0;
    layer3_outputs(1357) <= not (a and b);
    layer3_outputs(1358) <= 1'b0;
    layer3_outputs(1359) <= 1'b0;
    layer3_outputs(1360) <= 1'b1;
    layer3_outputs(1361) <= b;
    layer3_outputs(1362) <= a or b;
    layer3_outputs(1363) <= 1'b1;
    layer3_outputs(1364) <= 1'b0;
    layer3_outputs(1365) <= b and not a;
    layer3_outputs(1366) <= not (a and b);
    layer3_outputs(1367) <= a or b;
    layer3_outputs(1368) <= a;
    layer3_outputs(1369) <= a and not b;
    layer3_outputs(1370) <= not (a and b);
    layer3_outputs(1371) <= a;
    layer3_outputs(1372) <= 1'b0;
    layer3_outputs(1373) <= 1'b1;
    layer3_outputs(1374) <= not a;
    layer3_outputs(1375) <= a and b;
    layer3_outputs(1376) <= not a;
    layer3_outputs(1377) <= not (a or b);
    layer3_outputs(1378) <= not (a and b);
    layer3_outputs(1379) <= 1'b0;
    layer3_outputs(1380) <= not (a and b);
    layer3_outputs(1381) <= 1'b0;
    layer3_outputs(1382) <= b;
    layer3_outputs(1383) <= a and b;
    layer3_outputs(1384) <= a and not b;
    layer3_outputs(1385) <= not a or b;
    layer3_outputs(1386) <= not b or a;
    layer3_outputs(1387) <= not b or a;
    layer3_outputs(1388) <= not b;
    layer3_outputs(1389) <= not (a and b);
    layer3_outputs(1390) <= b;
    layer3_outputs(1391) <= 1'b0;
    layer3_outputs(1392) <= not a;
    layer3_outputs(1393) <= b and not a;
    layer3_outputs(1394) <= a;
    layer3_outputs(1395) <= not (a and b);
    layer3_outputs(1396) <= not a;
    layer3_outputs(1397) <= not (a or b);
    layer3_outputs(1398) <= b;
    layer3_outputs(1399) <= not (a and b);
    layer3_outputs(1400) <= 1'b0;
    layer3_outputs(1401) <= not b or a;
    layer3_outputs(1402) <= b;
    layer3_outputs(1403) <= not (a and b);
    layer3_outputs(1404) <= 1'b0;
    layer3_outputs(1405) <= not a or b;
    layer3_outputs(1406) <= a and b;
    layer3_outputs(1407) <= not a;
    layer3_outputs(1408) <= not a;
    layer3_outputs(1409) <= 1'b0;
    layer3_outputs(1410) <= not b;
    layer3_outputs(1411) <= not a or b;
    layer3_outputs(1412) <= not b or a;
    layer3_outputs(1413) <= not (a and b);
    layer3_outputs(1414) <= not (a and b);
    layer3_outputs(1415) <= 1'b0;
    layer3_outputs(1416) <= a and not b;
    layer3_outputs(1417) <= a and not b;
    layer3_outputs(1418) <= not b or a;
    layer3_outputs(1419) <= not (a and b);
    layer3_outputs(1420) <= a or b;
    layer3_outputs(1421) <= b and not a;
    layer3_outputs(1422) <= not b or a;
    layer3_outputs(1423) <= a;
    layer3_outputs(1424) <= b;
    layer3_outputs(1425) <= not (a or b);
    layer3_outputs(1426) <= b and not a;
    layer3_outputs(1427) <= not (a and b);
    layer3_outputs(1428) <= not a;
    layer3_outputs(1429) <= a;
    layer3_outputs(1430) <= a and b;
    layer3_outputs(1431) <= 1'b1;
    layer3_outputs(1432) <= not (a or b);
    layer3_outputs(1433) <= not a;
    layer3_outputs(1434) <= a or b;
    layer3_outputs(1435) <= not a or b;
    layer3_outputs(1436) <= b;
    layer3_outputs(1437) <= not b;
    layer3_outputs(1438) <= 1'b1;
    layer3_outputs(1439) <= 1'b0;
    layer3_outputs(1440) <= not b;
    layer3_outputs(1441) <= 1'b0;
    layer3_outputs(1442) <= not (a and b);
    layer3_outputs(1443) <= not a or b;
    layer3_outputs(1444) <= not a or b;
    layer3_outputs(1445) <= not b;
    layer3_outputs(1446) <= a and b;
    layer3_outputs(1447) <= b and not a;
    layer3_outputs(1448) <= a and b;
    layer3_outputs(1449) <= a and not b;
    layer3_outputs(1450) <= not b;
    layer3_outputs(1451) <= b and not a;
    layer3_outputs(1452) <= b and not a;
    layer3_outputs(1453) <= not (a and b);
    layer3_outputs(1454) <= b;
    layer3_outputs(1455) <= b;
    layer3_outputs(1456) <= a and b;
    layer3_outputs(1457) <= not a;
    layer3_outputs(1458) <= b;
    layer3_outputs(1459) <= b;
    layer3_outputs(1460) <= not (a and b);
    layer3_outputs(1461) <= b and not a;
    layer3_outputs(1462) <= not b;
    layer3_outputs(1463) <= a or b;
    layer3_outputs(1464) <= not a or b;
    layer3_outputs(1465) <= not (a and b);
    layer3_outputs(1466) <= a;
    layer3_outputs(1467) <= a and b;
    layer3_outputs(1468) <= b;
    layer3_outputs(1469) <= a and not b;
    layer3_outputs(1470) <= not a or b;
    layer3_outputs(1471) <= 1'b0;
    layer3_outputs(1472) <= not (a or b);
    layer3_outputs(1473) <= b;
    layer3_outputs(1474) <= b;
    layer3_outputs(1475) <= 1'b0;
    layer3_outputs(1476) <= not b or a;
    layer3_outputs(1477) <= a;
    layer3_outputs(1478) <= not b;
    layer3_outputs(1479) <= a or b;
    layer3_outputs(1480) <= 1'b1;
    layer3_outputs(1481) <= a;
    layer3_outputs(1482) <= a and b;
    layer3_outputs(1483) <= 1'b0;
    layer3_outputs(1484) <= not b;
    layer3_outputs(1485) <= not b or a;
    layer3_outputs(1486) <= a;
    layer3_outputs(1487) <= not b;
    layer3_outputs(1488) <= a and not b;
    layer3_outputs(1489) <= 1'b1;
    layer3_outputs(1490) <= not a;
    layer3_outputs(1491) <= not (a and b);
    layer3_outputs(1492) <= not a or b;
    layer3_outputs(1493) <= a;
    layer3_outputs(1494) <= not a or b;
    layer3_outputs(1495) <= b and not a;
    layer3_outputs(1496) <= not b;
    layer3_outputs(1497) <= b;
    layer3_outputs(1498) <= not a;
    layer3_outputs(1499) <= not b or a;
    layer3_outputs(1500) <= not (a and b);
    layer3_outputs(1501) <= b and not a;
    layer3_outputs(1502) <= not b;
    layer3_outputs(1503) <= a and b;
    layer3_outputs(1504) <= not b or a;
    layer3_outputs(1505) <= 1'b1;
    layer3_outputs(1506) <= 1'b0;
    layer3_outputs(1507) <= not (a or b);
    layer3_outputs(1508) <= a;
    layer3_outputs(1509) <= 1'b1;
    layer3_outputs(1510) <= b;
    layer3_outputs(1511) <= not (a and b);
    layer3_outputs(1512) <= b and not a;
    layer3_outputs(1513) <= not (a or b);
    layer3_outputs(1514) <= b;
    layer3_outputs(1515) <= not a or b;
    layer3_outputs(1516) <= 1'b0;
    layer3_outputs(1517) <= b;
    layer3_outputs(1518) <= not b or a;
    layer3_outputs(1519) <= not a or b;
    layer3_outputs(1520) <= a xor b;
    layer3_outputs(1521) <= not b or a;
    layer3_outputs(1522) <= b and not a;
    layer3_outputs(1523) <= not (a xor b);
    layer3_outputs(1524) <= not a;
    layer3_outputs(1525) <= not (a or b);
    layer3_outputs(1526) <= not a or b;
    layer3_outputs(1527) <= 1'b0;
    layer3_outputs(1528) <= not b or a;
    layer3_outputs(1529) <= 1'b1;
    layer3_outputs(1530) <= a and b;
    layer3_outputs(1531) <= not b or a;
    layer3_outputs(1532) <= not (a and b);
    layer3_outputs(1533) <= a;
    layer3_outputs(1534) <= a and not b;
    layer3_outputs(1535) <= not (a or b);
    layer3_outputs(1536) <= not a or b;
    layer3_outputs(1537) <= a xor b;
    layer3_outputs(1538) <= not a or b;
    layer3_outputs(1539) <= not b;
    layer3_outputs(1540) <= not (a or b);
    layer3_outputs(1541) <= a and b;
    layer3_outputs(1542) <= not b or a;
    layer3_outputs(1543) <= 1'b0;
    layer3_outputs(1544) <= b and not a;
    layer3_outputs(1545) <= a and b;
    layer3_outputs(1546) <= a xor b;
    layer3_outputs(1547) <= a or b;
    layer3_outputs(1548) <= 1'b0;
    layer3_outputs(1549) <= not (a and b);
    layer3_outputs(1550) <= a and b;
    layer3_outputs(1551) <= not a or b;
    layer3_outputs(1552) <= b and not a;
    layer3_outputs(1553) <= not (a or b);
    layer3_outputs(1554) <= not b;
    layer3_outputs(1555) <= not (a or b);
    layer3_outputs(1556) <= a and b;
    layer3_outputs(1557) <= a or b;
    layer3_outputs(1558) <= 1'b0;
    layer3_outputs(1559) <= a or b;
    layer3_outputs(1560) <= b and not a;
    layer3_outputs(1561) <= a and not b;
    layer3_outputs(1562) <= not b;
    layer3_outputs(1563) <= not (a and b);
    layer3_outputs(1564) <= a and b;
    layer3_outputs(1565) <= not b or a;
    layer3_outputs(1566) <= a and b;
    layer3_outputs(1567) <= a and not b;
    layer3_outputs(1568) <= not a;
    layer3_outputs(1569) <= b and not a;
    layer3_outputs(1570) <= a and not b;
    layer3_outputs(1571) <= 1'b0;
    layer3_outputs(1572) <= b;
    layer3_outputs(1573) <= a or b;
    layer3_outputs(1574) <= not (a and b);
    layer3_outputs(1575) <= a xor b;
    layer3_outputs(1576) <= not b or a;
    layer3_outputs(1577) <= b;
    layer3_outputs(1578) <= 1'b1;
    layer3_outputs(1579) <= 1'b1;
    layer3_outputs(1580) <= not a;
    layer3_outputs(1581) <= not b or a;
    layer3_outputs(1582) <= not (a or b);
    layer3_outputs(1583) <= b;
    layer3_outputs(1584) <= 1'b1;
    layer3_outputs(1585) <= 1'b1;
    layer3_outputs(1586) <= 1'b0;
    layer3_outputs(1587) <= b;
    layer3_outputs(1588) <= a and not b;
    layer3_outputs(1589) <= 1'b0;
    layer3_outputs(1590) <= a and b;
    layer3_outputs(1591) <= a or b;
    layer3_outputs(1592) <= a or b;
    layer3_outputs(1593) <= 1'b1;
    layer3_outputs(1594) <= 1'b0;
    layer3_outputs(1595) <= a;
    layer3_outputs(1596) <= not (a and b);
    layer3_outputs(1597) <= a;
    layer3_outputs(1598) <= 1'b0;
    layer3_outputs(1599) <= not a or b;
    layer3_outputs(1600) <= 1'b1;
    layer3_outputs(1601) <= b;
    layer3_outputs(1602) <= 1'b0;
    layer3_outputs(1603) <= 1'b0;
    layer3_outputs(1604) <= b and not a;
    layer3_outputs(1605) <= not (a or b);
    layer3_outputs(1606) <= 1'b0;
    layer3_outputs(1607) <= 1'b0;
    layer3_outputs(1608) <= b and not a;
    layer3_outputs(1609) <= 1'b0;
    layer3_outputs(1610) <= not (a or b);
    layer3_outputs(1611) <= not (a or b);
    layer3_outputs(1612) <= not (a and b);
    layer3_outputs(1613) <= 1'b1;
    layer3_outputs(1614) <= not (a and b);
    layer3_outputs(1615) <= a and not b;
    layer3_outputs(1616) <= 1'b0;
    layer3_outputs(1617) <= 1'b1;
    layer3_outputs(1618) <= not b or a;
    layer3_outputs(1619) <= a or b;
    layer3_outputs(1620) <= b;
    layer3_outputs(1621) <= a and b;
    layer3_outputs(1622) <= not b or a;
    layer3_outputs(1623) <= 1'b0;
    layer3_outputs(1624) <= 1'b1;
    layer3_outputs(1625) <= b and not a;
    layer3_outputs(1626) <= a and not b;
    layer3_outputs(1627) <= a or b;
    layer3_outputs(1628) <= not b or a;
    layer3_outputs(1629) <= not a;
    layer3_outputs(1630) <= a and b;
    layer3_outputs(1631) <= not a;
    layer3_outputs(1632) <= a;
    layer3_outputs(1633) <= a or b;
    layer3_outputs(1634) <= 1'b0;
    layer3_outputs(1635) <= not (a or b);
    layer3_outputs(1636) <= not b or a;
    layer3_outputs(1637) <= not a or b;
    layer3_outputs(1638) <= 1'b0;
    layer3_outputs(1639) <= not a;
    layer3_outputs(1640) <= b;
    layer3_outputs(1641) <= not a or b;
    layer3_outputs(1642) <= not a or b;
    layer3_outputs(1643) <= 1'b1;
    layer3_outputs(1644) <= a or b;
    layer3_outputs(1645) <= a and b;
    layer3_outputs(1646) <= 1'b0;
    layer3_outputs(1647) <= b and not a;
    layer3_outputs(1648) <= b;
    layer3_outputs(1649) <= b and not a;
    layer3_outputs(1650) <= 1'b0;
    layer3_outputs(1651) <= not b or a;
    layer3_outputs(1652) <= not a;
    layer3_outputs(1653) <= not (a xor b);
    layer3_outputs(1654) <= b and not a;
    layer3_outputs(1655) <= a;
    layer3_outputs(1656) <= not b or a;
    layer3_outputs(1657) <= not b;
    layer3_outputs(1658) <= a and b;
    layer3_outputs(1659) <= not (a and b);
    layer3_outputs(1660) <= 1'b1;
    layer3_outputs(1661) <= b and not a;
    layer3_outputs(1662) <= a and not b;
    layer3_outputs(1663) <= 1'b0;
    layer3_outputs(1664) <= not a;
    layer3_outputs(1665) <= not a or b;
    layer3_outputs(1666) <= not (a and b);
    layer3_outputs(1667) <= 1'b0;
    layer3_outputs(1668) <= a and b;
    layer3_outputs(1669) <= not a or b;
    layer3_outputs(1670) <= 1'b1;
    layer3_outputs(1671) <= not b or a;
    layer3_outputs(1672) <= a and not b;
    layer3_outputs(1673) <= a and b;
    layer3_outputs(1674) <= not (a and b);
    layer3_outputs(1675) <= a or b;
    layer3_outputs(1676) <= not a;
    layer3_outputs(1677) <= not b or a;
    layer3_outputs(1678) <= not b;
    layer3_outputs(1679) <= b;
    layer3_outputs(1680) <= not a or b;
    layer3_outputs(1681) <= a and not b;
    layer3_outputs(1682) <= a and not b;
    layer3_outputs(1683) <= 1'b1;
    layer3_outputs(1684) <= 1'b1;
    layer3_outputs(1685) <= not (a and b);
    layer3_outputs(1686) <= not a or b;
    layer3_outputs(1687) <= not b or a;
    layer3_outputs(1688) <= not a or b;
    layer3_outputs(1689) <= a or b;
    layer3_outputs(1690) <= not (a and b);
    layer3_outputs(1691) <= b;
    layer3_outputs(1692) <= a;
    layer3_outputs(1693) <= not (a xor b);
    layer3_outputs(1694) <= 1'b0;
    layer3_outputs(1695) <= not (a and b);
    layer3_outputs(1696) <= not b;
    layer3_outputs(1697) <= not a or b;
    layer3_outputs(1698) <= not b or a;
    layer3_outputs(1699) <= 1'b0;
    layer3_outputs(1700) <= b and not a;
    layer3_outputs(1701) <= not a or b;
    layer3_outputs(1702) <= a xor b;
    layer3_outputs(1703) <= a or b;
    layer3_outputs(1704) <= a;
    layer3_outputs(1705) <= not b or a;
    layer3_outputs(1706) <= not (a xor b);
    layer3_outputs(1707) <= b;
    layer3_outputs(1708) <= not a;
    layer3_outputs(1709) <= not a;
    layer3_outputs(1710) <= not (a and b);
    layer3_outputs(1711) <= a and not b;
    layer3_outputs(1712) <= a and not b;
    layer3_outputs(1713) <= not a or b;
    layer3_outputs(1714) <= a and b;
    layer3_outputs(1715) <= a and b;
    layer3_outputs(1716) <= not b;
    layer3_outputs(1717) <= not a or b;
    layer3_outputs(1718) <= b;
    layer3_outputs(1719) <= a and b;
    layer3_outputs(1720) <= b;
    layer3_outputs(1721) <= a and b;
    layer3_outputs(1722) <= a and not b;
    layer3_outputs(1723) <= not (a or b);
    layer3_outputs(1724) <= 1'b1;
    layer3_outputs(1725) <= not (a and b);
    layer3_outputs(1726) <= a or b;
    layer3_outputs(1727) <= a and b;
    layer3_outputs(1728) <= not (a or b);
    layer3_outputs(1729) <= not a;
    layer3_outputs(1730) <= a and b;
    layer3_outputs(1731) <= not (a and b);
    layer3_outputs(1732) <= a and not b;
    layer3_outputs(1733) <= not b or a;
    layer3_outputs(1734) <= 1'b0;
    layer3_outputs(1735) <= a;
    layer3_outputs(1736) <= a and b;
    layer3_outputs(1737) <= a and b;
    layer3_outputs(1738) <= a and not b;
    layer3_outputs(1739) <= not a;
    layer3_outputs(1740) <= a;
    layer3_outputs(1741) <= not a or b;
    layer3_outputs(1742) <= a and not b;
    layer3_outputs(1743) <= not a or b;
    layer3_outputs(1744) <= 1'b0;
    layer3_outputs(1745) <= b;
    layer3_outputs(1746) <= a xor b;
    layer3_outputs(1747) <= b and not a;
    layer3_outputs(1748) <= not b;
    layer3_outputs(1749) <= not a or b;
    layer3_outputs(1750) <= a and b;
    layer3_outputs(1751) <= a and b;
    layer3_outputs(1752) <= 1'b1;
    layer3_outputs(1753) <= not (a or b);
    layer3_outputs(1754) <= not b or a;
    layer3_outputs(1755) <= a and b;
    layer3_outputs(1756) <= not a;
    layer3_outputs(1757) <= 1'b0;
    layer3_outputs(1758) <= a;
    layer3_outputs(1759) <= not (a or b);
    layer3_outputs(1760) <= not b or a;
    layer3_outputs(1761) <= not a or b;
    layer3_outputs(1762) <= not a or b;
    layer3_outputs(1763) <= not b or a;
    layer3_outputs(1764) <= not b;
    layer3_outputs(1765) <= 1'b0;
    layer3_outputs(1766) <= a and b;
    layer3_outputs(1767) <= a and b;
    layer3_outputs(1768) <= not a or b;
    layer3_outputs(1769) <= b and not a;
    layer3_outputs(1770) <= not a;
    layer3_outputs(1771) <= not b;
    layer3_outputs(1772) <= not b or a;
    layer3_outputs(1773) <= a;
    layer3_outputs(1774) <= not a;
    layer3_outputs(1775) <= b;
    layer3_outputs(1776) <= not (a or b);
    layer3_outputs(1777) <= b and not a;
    layer3_outputs(1778) <= a;
    layer3_outputs(1779) <= 1'b0;
    layer3_outputs(1780) <= 1'b1;
    layer3_outputs(1781) <= not (a and b);
    layer3_outputs(1782) <= 1'b0;
    layer3_outputs(1783) <= a;
    layer3_outputs(1784) <= a or b;
    layer3_outputs(1785) <= b;
    layer3_outputs(1786) <= not a or b;
    layer3_outputs(1787) <= 1'b1;
    layer3_outputs(1788) <= b;
    layer3_outputs(1789) <= not b or a;
    layer3_outputs(1790) <= b;
    layer3_outputs(1791) <= b;
    layer3_outputs(1792) <= a or b;
    layer3_outputs(1793) <= b;
    layer3_outputs(1794) <= not b;
    layer3_outputs(1795) <= not (a and b);
    layer3_outputs(1796) <= not (a or b);
    layer3_outputs(1797) <= a and b;
    layer3_outputs(1798) <= not a or b;
    layer3_outputs(1799) <= not a or b;
    layer3_outputs(1800) <= a and b;
    layer3_outputs(1801) <= a;
    layer3_outputs(1802) <= not a or b;
    layer3_outputs(1803) <= not (a and b);
    layer3_outputs(1804) <= b;
    layer3_outputs(1805) <= b;
    layer3_outputs(1806) <= not a or b;
    layer3_outputs(1807) <= a;
    layer3_outputs(1808) <= a and b;
    layer3_outputs(1809) <= a and not b;
    layer3_outputs(1810) <= not b;
    layer3_outputs(1811) <= not a;
    layer3_outputs(1812) <= a and b;
    layer3_outputs(1813) <= 1'b0;
    layer3_outputs(1814) <= 1'b0;
    layer3_outputs(1815) <= not (a and b);
    layer3_outputs(1816) <= 1'b1;
    layer3_outputs(1817) <= b;
    layer3_outputs(1818) <= b;
    layer3_outputs(1819) <= 1'b1;
    layer3_outputs(1820) <= not a;
    layer3_outputs(1821) <= 1'b0;
    layer3_outputs(1822) <= not (a or b);
    layer3_outputs(1823) <= a or b;
    layer3_outputs(1824) <= not a or b;
    layer3_outputs(1825) <= not (a or b);
    layer3_outputs(1826) <= a and b;
    layer3_outputs(1827) <= not b or a;
    layer3_outputs(1828) <= not b or a;
    layer3_outputs(1829) <= 1'b0;
    layer3_outputs(1830) <= 1'b1;
    layer3_outputs(1831) <= a and b;
    layer3_outputs(1832) <= 1'b0;
    layer3_outputs(1833) <= not (a and b);
    layer3_outputs(1834) <= 1'b0;
    layer3_outputs(1835) <= a and b;
    layer3_outputs(1836) <= 1'b0;
    layer3_outputs(1837) <= a;
    layer3_outputs(1838) <= not a or b;
    layer3_outputs(1839) <= not (a or b);
    layer3_outputs(1840) <= not a or b;
    layer3_outputs(1841) <= not b;
    layer3_outputs(1842) <= not a or b;
    layer3_outputs(1843) <= 1'b0;
    layer3_outputs(1844) <= a or b;
    layer3_outputs(1845) <= b and not a;
    layer3_outputs(1846) <= not b or a;
    layer3_outputs(1847) <= a and not b;
    layer3_outputs(1848) <= b;
    layer3_outputs(1849) <= 1'b0;
    layer3_outputs(1850) <= b and not a;
    layer3_outputs(1851) <= a and b;
    layer3_outputs(1852) <= b and not a;
    layer3_outputs(1853) <= a and not b;
    layer3_outputs(1854) <= not a;
    layer3_outputs(1855) <= not a or b;
    layer3_outputs(1856) <= a;
    layer3_outputs(1857) <= not a;
    layer3_outputs(1858) <= b and not a;
    layer3_outputs(1859) <= not (a and b);
    layer3_outputs(1860) <= b and not a;
    layer3_outputs(1861) <= a;
    layer3_outputs(1862) <= a or b;
    layer3_outputs(1863) <= b and not a;
    layer3_outputs(1864) <= not b;
    layer3_outputs(1865) <= b and not a;
    layer3_outputs(1866) <= b and not a;
    layer3_outputs(1867) <= a;
    layer3_outputs(1868) <= not b or a;
    layer3_outputs(1869) <= b and not a;
    layer3_outputs(1870) <= not a;
    layer3_outputs(1871) <= a and not b;
    layer3_outputs(1872) <= not (a and b);
    layer3_outputs(1873) <= not a;
    layer3_outputs(1874) <= not b;
    layer3_outputs(1875) <= not b or a;
    layer3_outputs(1876) <= not a;
    layer3_outputs(1877) <= not (a or b);
    layer3_outputs(1878) <= a;
    layer3_outputs(1879) <= not b;
    layer3_outputs(1880) <= a and not b;
    layer3_outputs(1881) <= b and not a;
    layer3_outputs(1882) <= 1'b0;
    layer3_outputs(1883) <= b and not a;
    layer3_outputs(1884) <= a;
    layer3_outputs(1885) <= not b;
    layer3_outputs(1886) <= a or b;
    layer3_outputs(1887) <= not (a and b);
    layer3_outputs(1888) <= not (a and b);
    layer3_outputs(1889) <= not (a or b);
    layer3_outputs(1890) <= b and not a;
    layer3_outputs(1891) <= not b or a;
    layer3_outputs(1892) <= not a;
    layer3_outputs(1893) <= not (a and b);
    layer3_outputs(1894) <= a;
    layer3_outputs(1895) <= a;
    layer3_outputs(1896) <= a and not b;
    layer3_outputs(1897) <= 1'b0;
    layer3_outputs(1898) <= a and b;
    layer3_outputs(1899) <= a;
    layer3_outputs(1900) <= 1'b1;
    layer3_outputs(1901) <= b;
    layer3_outputs(1902) <= not (a and b);
    layer3_outputs(1903) <= 1'b1;
    layer3_outputs(1904) <= not (a and b);
    layer3_outputs(1905) <= 1'b0;
    layer3_outputs(1906) <= b;
    layer3_outputs(1907) <= not (a and b);
    layer3_outputs(1908) <= b;
    layer3_outputs(1909) <= 1'b1;
    layer3_outputs(1910) <= not (a and b);
    layer3_outputs(1911) <= a and b;
    layer3_outputs(1912) <= a or b;
    layer3_outputs(1913) <= a;
    layer3_outputs(1914) <= not b;
    layer3_outputs(1915) <= b;
    layer3_outputs(1916) <= 1'b1;
    layer3_outputs(1917) <= 1'b0;
    layer3_outputs(1918) <= a or b;
    layer3_outputs(1919) <= 1'b0;
    layer3_outputs(1920) <= not (a or b);
    layer3_outputs(1921) <= 1'b1;
    layer3_outputs(1922) <= a or b;
    layer3_outputs(1923) <= not b or a;
    layer3_outputs(1924) <= 1'b0;
    layer3_outputs(1925) <= 1'b0;
    layer3_outputs(1926) <= 1'b1;
    layer3_outputs(1927) <= not (a and b);
    layer3_outputs(1928) <= b and not a;
    layer3_outputs(1929) <= b;
    layer3_outputs(1930) <= not b or a;
    layer3_outputs(1931) <= a;
    layer3_outputs(1932) <= a or b;
    layer3_outputs(1933) <= a or b;
    layer3_outputs(1934) <= b and not a;
    layer3_outputs(1935) <= not b or a;
    layer3_outputs(1936) <= not (a and b);
    layer3_outputs(1937) <= a or b;
    layer3_outputs(1938) <= a and b;
    layer3_outputs(1939) <= b and not a;
    layer3_outputs(1940) <= a or b;
    layer3_outputs(1941) <= not (a and b);
    layer3_outputs(1942) <= a and not b;
    layer3_outputs(1943) <= 1'b0;
    layer3_outputs(1944) <= not b;
    layer3_outputs(1945) <= 1'b1;
    layer3_outputs(1946) <= not a or b;
    layer3_outputs(1947) <= not (a or b);
    layer3_outputs(1948) <= b and not a;
    layer3_outputs(1949) <= a and not b;
    layer3_outputs(1950) <= a or b;
    layer3_outputs(1951) <= not (a or b);
    layer3_outputs(1952) <= a and not b;
    layer3_outputs(1953) <= a;
    layer3_outputs(1954) <= b and not a;
    layer3_outputs(1955) <= not (a xor b);
    layer3_outputs(1956) <= not a or b;
    layer3_outputs(1957) <= 1'b0;
    layer3_outputs(1958) <= a and b;
    layer3_outputs(1959) <= not a or b;
    layer3_outputs(1960) <= a or b;
    layer3_outputs(1961) <= not b or a;
    layer3_outputs(1962) <= a or b;
    layer3_outputs(1963) <= not a;
    layer3_outputs(1964) <= 1'b1;
    layer3_outputs(1965) <= b;
    layer3_outputs(1966) <= 1'b0;
    layer3_outputs(1967) <= 1'b0;
    layer3_outputs(1968) <= not b;
    layer3_outputs(1969) <= a and b;
    layer3_outputs(1970) <= not (a xor b);
    layer3_outputs(1971) <= not b;
    layer3_outputs(1972) <= not b or a;
    layer3_outputs(1973) <= not (a and b);
    layer3_outputs(1974) <= 1'b0;
    layer3_outputs(1975) <= not (a and b);
    layer3_outputs(1976) <= not b or a;
    layer3_outputs(1977) <= not a;
    layer3_outputs(1978) <= not b;
    layer3_outputs(1979) <= not b or a;
    layer3_outputs(1980) <= a;
    layer3_outputs(1981) <= not b or a;
    layer3_outputs(1982) <= 1'b0;
    layer3_outputs(1983) <= a or b;
    layer3_outputs(1984) <= not b;
    layer3_outputs(1985) <= not a;
    layer3_outputs(1986) <= not b or a;
    layer3_outputs(1987) <= not b;
    layer3_outputs(1988) <= a and not b;
    layer3_outputs(1989) <= 1'b1;
    layer3_outputs(1990) <= 1'b1;
    layer3_outputs(1991) <= a;
    layer3_outputs(1992) <= 1'b0;
    layer3_outputs(1993) <= b;
    layer3_outputs(1994) <= b and not a;
    layer3_outputs(1995) <= not a;
    layer3_outputs(1996) <= b;
    layer3_outputs(1997) <= not b or a;
    layer3_outputs(1998) <= not a;
    layer3_outputs(1999) <= not b;
    layer3_outputs(2000) <= not b or a;
    layer3_outputs(2001) <= not a or b;
    layer3_outputs(2002) <= not a or b;
    layer3_outputs(2003) <= 1'b0;
    layer3_outputs(2004) <= b and not a;
    layer3_outputs(2005) <= not a or b;
    layer3_outputs(2006) <= a and not b;
    layer3_outputs(2007) <= 1'b1;
    layer3_outputs(2008) <= 1'b1;
    layer3_outputs(2009) <= not (a or b);
    layer3_outputs(2010) <= a;
    layer3_outputs(2011) <= 1'b0;
    layer3_outputs(2012) <= b and not a;
    layer3_outputs(2013) <= b and not a;
    layer3_outputs(2014) <= not (a or b);
    layer3_outputs(2015) <= not a;
    layer3_outputs(2016) <= not (a and b);
    layer3_outputs(2017) <= not (a and b);
    layer3_outputs(2018) <= not (a and b);
    layer3_outputs(2019) <= not b;
    layer3_outputs(2020) <= a and b;
    layer3_outputs(2021) <= not (a or b);
    layer3_outputs(2022) <= a;
    layer3_outputs(2023) <= not (a or b);
    layer3_outputs(2024) <= a;
    layer3_outputs(2025) <= a;
    layer3_outputs(2026) <= a and b;
    layer3_outputs(2027) <= not b or a;
    layer3_outputs(2028) <= not b or a;
    layer3_outputs(2029) <= not a or b;
    layer3_outputs(2030) <= 1'b0;
    layer3_outputs(2031) <= not (a or b);
    layer3_outputs(2032) <= a;
    layer3_outputs(2033) <= a and not b;
    layer3_outputs(2034) <= b and not a;
    layer3_outputs(2035) <= not a;
    layer3_outputs(2036) <= not a;
    layer3_outputs(2037) <= not (a and b);
    layer3_outputs(2038) <= 1'b0;
    layer3_outputs(2039) <= 1'b1;
    layer3_outputs(2040) <= a or b;
    layer3_outputs(2041) <= not a or b;
    layer3_outputs(2042) <= a and b;
    layer3_outputs(2043) <= not b or a;
    layer3_outputs(2044) <= a or b;
    layer3_outputs(2045) <= b;
    layer3_outputs(2046) <= not a;
    layer3_outputs(2047) <= 1'b0;
    layer3_outputs(2048) <= a and b;
    layer3_outputs(2049) <= b and not a;
    layer3_outputs(2050) <= not (a and b);
    layer3_outputs(2051) <= a and b;
    layer3_outputs(2052) <= not (a xor b);
    layer3_outputs(2053) <= not (a and b);
    layer3_outputs(2054) <= b;
    layer3_outputs(2055) <= not a or b;
    layer3_outputs(2056) <= not (a and b);
    layer3_outputs(2057) <= b;
    layer3_outputs(2058) <= not a;
    layer3_outputs(2059) <= 1'b1;
    layer3_outputs(2060) <= a xor b;
    layer3_outputs(2061) <= not b or a;
    layer3_outputs(2062) <= not (a or b);
    layer3_outputs(2063) <= not b;
    layer3_outputs(2064) <= 1'b0;
    layer3_outputs(2065) <= a and not b;
    layer3_outputs(2066) <= not (a or b);
    layer3_outputs(2067) <= not a;
    layer3_outputs(2068) <= 1'b1;
    layer3_outputs(2069) <= 1'b0;
    layer3_outputs(2070) <= not b or a;
    layer3_outputs(2071) <= not b;
    layer3_outputs(2072) <= a and b;
    layer3_outputs(2073) <= a;
    layer3_outputs(2074) <= b and not a;
    layer3_outputs(2075) <= not (a or b);
    layer3_outputs(2076) <= not b;
    layer3_outputs(2077) <= a or b;
    layer3_outputs(2078) <= not (a or b);
    layer3_outputs(2079) <= not (a and b);
    layer3_outputs(2080) <= b;
    layer3_outputs(2081) <= a and not b;
    layer3_outputs(2082) <= not (a or b);
    layer3_outputs(2083) <= not a;
    layer3_outputs(2084) <= a and b;
    layer3_outputs(2085) <= not (a and b);
    layer3_outputs(2086) <= a and not b;
    layer3_outputs(2087) <= 1'b0;
    layer3_outputs(2088) <= a;
    layer3_outputs(2089) <= a and b;
    layer3_outputs(2090) <= 1'b0;
    layer3_outputs(2091) <= not b;
    layer3_outputs(2092) <= 1'b0;
    layer3_outputs(2093) <= a and b;
    layer3_outputs(2094) <= a;
    layer3_outputs(2095) <= 1'b0;
    layer3_outputs(2096) <= 1'b1;
    layer3_outputs(2097) <= a and not b;
    layer3_outputs(2098) <= a and b;
    layer3_outputs(2099) <= a or b;
    layer3_outputs(2100) <= not (a or b);
    layer3_outputs(2101) <= 1'b1;
    layer3_outputs(2102) <= 1'b1;
    layer3_outputs(2103) <= not (a and b);
    layer3_outputs(2104) <= not a or b;
    layer3_outputs(2105) <= not a;
    layer3_outputs(2106) <= 1'b0;
    layer3_outputs(2107) <= 1'b0;
    layer3_outputs(2108) <= not b or a;
    layer3_outputs(2109) <= not a;
    layer3_outputs(2110) <= not b;
    layer3_outputs(2111) <= not (a and b);
    layer3_outputs(2112) <= not (a or b);
    layer3_outputs(2113) <= not a;
    layer3_outputs(2114) <= 1'b0;
    layer3_outputs(2115) <= not b or a;
    layer3_outputs(2116) <= a;
    layer3_outputs(2117) <= not a or b;
    layer3_outputs(2118) <= not a or b;
    layer3_outputs(2119) <= b;
    layer3_outputs(2120) <= b and not a;
    layer3_outputs(2121) <= not (a or b);
    layer3_outputs(2122) <= 1'b0;
    layer3_outputs(2123) <= a and b;
    layer3_outputs(2124) <= a;
    layer3_outputs(2125) <= not b;
    layer3_outputs(2126) <= not b;
    layer3_outputs(2127) <= 1'b1;
    layer3_outputs(2128) <= a and not b;
    layer3_outputs(2129) <= not (a or b);
    layer3_outputs(2130) <= not b or a;
    layer3_outputs(2131) <= 1'b1;
    layer3_outputs(2132) <= not b;
    layer3_outputs(2133) <= not a or b;
    layer3_outputs(2134) <= a;
    layer3_outputs(2135) <= 1'b1;
    layer3_outputs(2136) <= b and not a;
    layer3_outputs(2137) <= 1'b0;
    layer3_outputs(2138) <= a or b;
    layer3_outputs(2139) <= b;
    layer3_outputs(2140) <= not b or a;
    layer3_outputs(2141) <= a and b;
    layer3_outputs(2142) <= b and not a;
    layer3_outputs(2143) <= 1'b1;
    layer3_outputs(2144) <= 1'b0;
    layer3_outputs(2145) <= a or b;
    layer3_outputs(2146) <= not b or a;
    layer3_outputs(2147) <= b and not a;
    layer3_outputs(2148) <= 1'b1;
    layer3_outputs(2149) <= not b or a;
    layer3_outputs(2150) <= not (a or b);
    layer3_outputs(2151) <= not (a or b);
    layer3_outputs(2152) <= a and not b;
    layer3_outputs(2153) <= not b or a;
    layer3_outputs(2154) <= 1'b1;
    layer3_outputs(2155) <= a and b;
    layer3_outputs(2156) <= a;
    layer3_outputs(2157) <= not (a xor b);
    layer3_outputs(2158) <= not a;
    layer3_outputs(2159) <= not a;
    layer3_outputs(2160) <= not b;
    layer3_outputs(2161) <= not (a or b);
    layer3_outputs(2162) <= a and b;
    layer3_outputs(2163) <= not a;
    layer3_outputs(2164) <= not (a or b);
    layer3_outputs(2165) <= 1'b1;
    layer3_outputs(2166) <= b and not a;
    layer3_outputs(2167) <= b;
    layer3_outputs(2168) <= a and not b;
    layer3_outputs(2169) <= not b or a;
    layer3_outputs(2170) <= 1'b0;
    layer3_outputs(2171) <= 1'b1;
    layer3_outputs(2172) <= a and b;
    layer3_outputs(2173) <= a and not b;
    layer3_outputs(2174) <= b;
    layer3_outputs(2175) <= 1'b1;
    layer3_outputs(2176) <= a;
    layer3_outputs(2177) <= not b or a;
    layer3_outputs(2178) <= a and b;
    layer3_outputs(2179) <= a and b;
    layer3_outputs(2180) <= a and not b;
    layer3_outputs(2181) <= 1'b0;
    layer3_outputs(2182) <= not a;
    layer3_outputs(2183) <= a and not b;
    layer3_outputs(2184) <= 1'b1;
    layer3_outputs(2185) <= 1'b0;
    layer3_outputs(2186) <= not b;
    layer3_outputs(2187) <= not a or b;
    layer3_outputs(2188) <= 1'b1;
    layer3_outputs(2189) <= not a or b;
    layer3_outputs(2190) <= not b;
    layer3_outputs(2191) <= a and not b;
    layer3_outputs(2192) <= not b;
    layer3_outputs(2193) <= not a;
    layer3_outputs(2194) <= not b;
    layer3_outputs(2195) <= not b or a;
    layer3_outputs(2196) <= not a or b;
    layer3_outputs(2197) <= not b or a;
    layer3_outputs(2198) <= 1'b1;
    layer3_outputs(2199) <= not a or b;
    layer3_outputs(2200) <= not a or b;
    layer3_outputs(2201) <= 1'b1;
    layer3_outputs(2202) <= a or b;
    layer3_outputs(2203) <= b;
    layer3_outputs(2204) <= 1'b1;
    layer3_outputs(2205) <= 1'b1;
    layer3_outputs(2206) <= not b;
    layer3_outputs(2207) <= a and not b;
    layer3_outputs(2208) <= b and not a;
    layer3_outputs(2209) <= a;
    layer3_outputs(2210) <= not (a and b);
    layer3_outputs(2211) <= a or b;
    layer3_outputs(2212) <= not a;
    layer3_outputs(2213) <= 1'b0;
    layer3_outputs(2214) <= not (a or b);
    layer3_outputs(2215) <= not a or b;
    layer3_outputs(2216) <= not b;
    layer3_outputs(2217) <= 1'b1;
    layer3_outputs(2218) <= a or b;
    layer3_outputs(2219) <= a or b;
    layer3_outputs(2220) <= not (a or b);
    layer3_outputs(2221) <= 1'b1;
    layer3_outputs(2222) <= not a or b;
    layer3_outputs(2223) <= a and not b;
    layer3_outputs(2224) <= not (a or b);
    layer3_outputs(2225) <= b;
    layer3_outputs(2226) <= not b;
    layer3_outputs(2227) <= not a or b;
    layer3_outputs(2228) <= not b;
    layer3_outputs(2229) <= 1'b1;
    layer3_outputs(2230) <= a or b;
    layer3_outputs(2231) <= not a or b;
    layer3_outputs(2232) <= not (a or b);
    layer3_outputs(2233) <= 1'b1;
    layer3_outputs(2234) <= not b;
    layer3_outputs(2235) <= a and not b;
    layer3_outputs(2236) <= not b;
    layer3_outputs(2237) <= b;
    layer3_outputs(2238) <= not b;
    layer3_outputs(2239) <= a and not b;
    layer3_outputs(2240) <= 1'b1;
    layer3_outputs(2241) <= b and not a;
    layer3_outputs(2242) <= not b or a;
    layer3_outputs(2243) <= a;
    layer3_outputs(2244) <= a;
    layer3_outputs(2245) <= not b;
    layer3_outputs(2246) <= not b or a;
    layer3_outputs(2247) <= a and b;
    layer3_outputs(2248) <= not b;
    layer3_outputs(2249) <= not b;
    layer3_outputs(2250) <= a and b;
    layer3_outputs(2251) <= not a;
    layer3_outputs(2252) <= not b or a;
    layer3_outputs(2253) <= a and not b;
    layer3_outputs(2254) <= 1'b0;
    layer3_outputs(2255) <= a or b;
    layer3_outputs(2256) <= b;
    layer3_outputs(2257) <= 1'b0;
    layer3_outputs(2258) <= not b;
    layer3_outputs(2259) <= not b;
    layer3_outputs(2260) <= a or b;
    layer3_outputs(2261) <= not a;
    layer3_outputs(2262) <= 1'b0;
    layer3_outputs(2263) <= a or b;
    layer3_outputs(2264) <= not a;
    layer3_outputs(2265) <= not b;
    layer3_outputs(2266) <= not b or a;
    layer3_outputs(2267) <= a;
    layer3_outputs(2268) <= not a or b;
    layer3_outputs(2269) <= b;
    layer3_outputs(2270) <= a or b;
    layer3_outputs(2271) <= not a;
    layer3_outputs(2272) <= b and not a;
    layer3_outputs(2273) <= not (a xor b);
    layer3_outputs(2274) <= not a or b;
    layer3_outputs(2275) <= 1'b1;
    layer3_outputs(2276) <= not a or b;
    layer3_outputs(2277) <= not (a and b);
    layer3_outputs(2278) <= a and not b;
    layer3_outputs(2279) <= not b or a;
    layer3_outputs(2280) <= a xor b;
    layer3_outputs(2281) <= not (a and b);
    layer3_outputs(2282) <= b;
    layer3_outputs(2283) <= not a or b;
    layer3_outputs(2284) <= a and not b;
    layer3_outputs(2285) <= 1'b1;
    layer3_outputs(2286) <= not b or a;
    layer3_outputs(2287) <= not (a or b);
    layer3_outputs(2288) <= a or b;
    layer3_outputs(2289) <= b and not a;
    layer3_outputs(2290) <= not a;
    layer3_outputs(2291) <= 1'b1;
    layer3_outputs(2292) <= 1'b1;
    layer3_outputs(2293) <= b and not a;
    layer3_outputs(2294) <= b;
    layer3_outputs(2295) <= 1'b0;
    layer3_outputs(2296) <= 1'b0;
    layer3_outputs(2297) <= a and not b;
    layer3_outputs(2298) <= not b or a;
    layer3_outputs(2299) <= not (a and b);
    layer3_outputs(2300) <= not (a or b);
    layer3_outputs(2301) <= not (a or b);
    layer3_outputs(2302) <= not a;
    layer3_outputs(2303) <= a and b;
    layer3_outputs(2304) <= a;
    layer3_outputs(2305) <= a xor b;
    layer3_outputs(2306) <= a or b;
    layer3_outputs(2307) <= a and b;
    layer3_outputs(2308) <= not (a or b);
    layer3_outputs(2309) <= b;
    layer3_outputs(2310) <= not b or a;
    layer3_outputs(2311) <= not b or a;
    layer3_outputs(2312) <= not (a or b);
    layer3_outputs(2313) <= a and b;
    layer3_outputs(2314) <= not b;
    layer3_outputs(2315) <= not a;
    layer3_outputs(2316) <= a or b;
    layer3_outputs(2317) <= a xor b;
    layer3_outputs(2318) <= 1'b1;
    layer3_outputs(2319) <= b and not a;
    layer3_outputs(2320) <= a or b;
    layer3_outputs(2321) <= 1'b0;
    layer3_outputs(2322) <= a or b;
    layer3_outputs(2323) <= not a or b;
    layer3_outputs(2324) <= not b;
    layer3_outputs(2325) <= b and not a;
    layer3_outputs(2326) <= a;
    layer3_outputs(2327) <= b;
    layer3_outputs(2328) <= not b;
    layer3_outputs(2329) <= a and not b;
    layer3_outputs(2330) <= 1'b0;
    layer3_outputs(2331) <= 1'b0;
    layer3_outputs(2332) <= not (a xor b);
    layer3_outputs(2333) <= not a or b;
    layer3_outputs(2334) <= a and not b;
    layer3_outputs(2335) <= a and not b;
    layer3_outputs(2336) <= a and not b;
    layer3_outputs(2337) <= not b or a;
    layer3_outputs(2338) <= a and not b;
    layer3_outputs(2339) <= a and b;
    layer3_outputs(2340) <= b;
    layer3_outputs(2341) <= not (a or b);
    layer3_outputs(2342) <= a and b;
    layer3_outputs(2343) <= not a or b;
    layer3_outputs(2344) <= not b or a;
    layer3_outputs(2345) <= b;
    layer3_outputs(2346) <= 1'b1;
    layer3_outputs(2347) <= 1'b1;
    layer3_outputs(2348) <= not (a or b);
    layer3_outputs(2349) <= a and not b;
    layer3_outputs(2350) <= a;
    layer3_outputs(2351) <= a and b;
    layer3_outputs(2352) <= not b or a;
    layer3_outputs(2353) <= 1'b1;
    layer3_outputs(2354) <= not (a or b);
    layer3_outputs(2355) <= not (a and b);
    layer3_outputs(2356) <= a or b;
    layer3_outputs(2357) <= not b or a;
    layer3_outputs(2358) <= a and not b;
    layer3_outputs(2359) <= a;
    layer3_outputs(2360) <= a or b;
    layer3_outputs(2361) <= 1'b0;
    layer3_outputs(2362) <= a or b;
    layer3_outputs(2363) <= a or b;
    layer3_outputs(2364) <= a and not b;
    layer3_outputs(2365) <= a and not b;
    layer3_outputs(2366) <= a and not b;
    layer3_outputs(2367) <= a;
    layer3_outputs(2368) <= 1'b1;
    layer3_outputs(2369) <= a and not b;
    layer3_outputs(2370) <= b;
    layer3_outputs(2371) <= b and not a;
    layer3_outputs(2372) <= a and not b;
    layer3_outputs(2373) <= a;
    layer3_outputs(2374) <= a or b;
    layer3_outputs(2375) <= not a or b;
    layer3_outputs(2376) <= 1'b0;
    layer3_outputs(2377) <= a;
    layer3_outputs(2378) <= 1'b0;
    layer3_outputs(2379) <= not (a or b);
    layer3_outputs(2380) <= not b;
    layer3_outputs(2381) <= a and b;
    layer3_outputs(2382) <= a and b;
    layer3_outputs(2383) <= b and not a;
    layer3_outputs(2384) <= b and not a;
    layer3_outputs(2385) <= a and b;
    layer3_outputs(2386) <= not (a and b);
    layer3_outputs(2387) <= b and not a;
    layer3_outputs(2388) <= not b;
    layer3_outputs(2389) <= a or b;
    layer3_outputs(2390) <= 1'b1;
    layer3_outputs(2391) <= not b or a;
    layer3_outputs(2392) <= not a or b;
    layer3_outputs(2393) <= b;
    layer3_outputs(2394) <= 1'b1;
    layer3_outputs(2395) <= 1'b1;
    layer3_outputs(2396) <= a or b;
    layer3_outputs(2397) <= not (a xor b);
    layer3_outputs(2398) <= a and b;
    layer3_outputs(2399) <= b;
    layer3_outputs(2400) <= 1'b0;
    layer3_outputs(2401) <= not b;
    layer3_outputs(2402) <= a or b;
    layer3_outputs(2403) <= not (a or b);
    layer3_outputs(2404) <= not a or b;
    layer3_outputs(2405) <= 1'b1;
    layer3_outputs(2406) <= 1'b0;
    layer3_outputs(2407) <= not a or b;
    layer3_outputs(2408) <= not (a and b);
    layer3_outputs(2409) <= 1'b1;
    layer3_outputs(2410) <= a xor b;
    layer3_outputs(2411) <= a and not b;
    layer3_outputs(2412) <= a;
    layer3_outputs(2413) <= not a;
    layer3_outputs(2414) <= not b or a;
    layer3_outputs(2415) <= not a or b;
    layer3_outputs(2416) <= not (a xor b);
    layer3_outputs(2417) <= 1'b0;
    layer3_outputs(2418) <= 1'b1;
    layer3_outputs(2419) <= a;
    layer3_outputs(2420) <= b and not a;
    layer3_outputs(2421) <= 1'b0;
    layer3_outputs(2422) <= not (a and b);
    layer3_outputs(2423) <= not (a and b);
    layer3_outputs(2424) <= not b or a;
    layer3_outputs(2425) <= a and b;
    layer3_outputs(2426) <= a or b;
    layer3_outputs(2427) <= not a;
    layer3_outputs(2428) <= not a or b;
    layer3_outputs(2429) <= b;
    layer3_outputs(2430) <= not (a or b);
    layer3_outputs(2431) <= a;
    layer3_outputs(2432) <= a;
    layer3_outputs(2433) <= not b;
    layer3_outputs(2434) <= a;
    layer3_outputs(2435) <= a and b;
    layer3_outputs(2436) <= not (a or b);
    layer3_outputs(2437) <= b;
    layer3_outputs(2438) <= 1'b0;
    layer3_outputs(2439) <= not (a or b);
    layer3_outputs(2440) <= not (a xor b);
    layer3_outputs(2441) <= a and b;
    layer3_outputs(2442) <= b and not a;
    layer3_outputs(2443) <= b;
    layer3_outputs(2444) <= a;
    layer3_outputs(2445) <= not (a and b);
    layer3_outputs(2446) <= not (a xor b);
    layer3_outputs(2447) <= not (a or b);
    layer3_outputs(2448) <= 1'b1;
    layer3_outputs(2449) <= not a;
    layer3_outputs(2450) <= 1'b1;
    layer3_outputs(2451) <= b;
    layer3_outputs(2452) <= a;
    layer3_outputs(2453) <= b;
    layer3_outputs(2454) <= a;
    layer3_outputs(2455) <= not b;
    layer3_outputs(2456) <= not (a or b);
    layer3_outputs(2457) <= a and b;
    layer3_outputs(2458) <= not (a or b);
    layer3_outputs(2459) <= b;
    layer3_outputs(2460) <= not (a or b);
    layer3_outputs(2461) <= not a or b;
    layer3_outputs(2462) <= b and not a;
    layer3_outputs(2463) <= a or b;
    layer3_outputs(2464) <= a;
    layer3_outputs(2465) <= b and not a;
    layer3_outputs(2466) <= not b or a;
    layer3_outputs(2467) <= not a or b;
    layer3_outputs(2468) <= b;
    layer3_outputs(2469) <= a and not b;
    layer3_outputs(2470) <= a xor b;
    layer3_outputs(2471) <= not b;
    layer3_outputs(2472) <= a;
    layer3_outputs(2473) <= not a or b;
    layer3_outputs(2474) <= b;
    layer3_outputs(2475) <= not a;
    layer3_outputs(2476) <= not a or b;
    layer3_outputs(2477) <= not b;
    layer3_outputs(2478) <= 1'b0;
    layer3_outputs(2479) <= b;
    layer3_outputs(2480) <= b and not a;
    layer3_outputs(2481) <= b;
    layer3_outputs(2482) <= not (a or b);
    layer3_outputs(2483) <= 1'b1;
    layer3_outputs(2484) <= not b;
    layer3_outputs(2485) <= not b or a;
    layer3_outputs(2486) <= a;
    layer3_outputs(2487) <= not b or a;
    layer3_outputs(2488) <= b and not a;
    layer3_outputs(2489) <= a and b;
    layer3_outputs(2490) <= a;
    layer3_outputs(2491) <= b and not a;
    layer3_outputs(2492) <= a and not b;
    layer3_outputs(2493) <= a xor b;
    layer3_outputs(2494) <= not (a xor b);
    layer3_outputs(2495) <= not b or a;
    layer3_outputs(2496) <= b and not a;
    layer3_outputs(2497) <= not b or a;
    layer3_outputs(2498) <= not b;
    layer3_outputs(2499) <= b;
    layer3_outputs(2500) <= not a or b;
    layer3_outputs(2501) <= not b;
    layer3_outputs(2502) <= not (a or b);
    layer3_outputs(2503) <= not b;
    layer3_outputs(2504) <= a or b;
    layer3_outputs(2505) <= 1'b0;
    layer3_outputs(2506) <= a xor b;
    layer3_outputs(2507) <= not b or a;
    layer3_outputs(2508) <= a xor b;
    layer3_outputs(2509) <= a and not b;
    layer3_outputs(2510) <= not b or a;
    layer3_outputs(2511) <= 1'b0;
    layer3_outputs(2512) <= not a;
    layer3_outputs(2513) <= not a or b;
    layer3_outputs(2514) <= 1'b1;
    layer3_outputs(2515) <= 1'b1;
    layer3_outputs(2516) <= a;
    layer3_outputs(2517) <= a;
    layer3_outputs(2518) <= 1'b0;
    layer3_outputs(2519) <= a and b;
    layer3_outputs(2520) <= not a or b;
    layer3_outputs(2521) <= a and not b;
    layer3_outputs(2522) <= 1'b1;
    layer3_outputs(2523) <= a or b;
    layer3_outputs(2524) <= not (a or b);
    layer3_outputs(2525) <= 1'b1;
    layer3_outputs(2526) <= a and b;
    layer3_outputs(2527) <= 1'b0;
    layer3_outputs(2528) <= 1'b1;
    layer3_outputs(2529) <= a;
    layer3_outputs(2530) <= not b or a;
    layer3_outputs(2531) <= not b or a;
    layer3_outputs(2532) <= not a or b;
    layer3_outputs(2533) <= a and b;
    layer3_outputs(2534) <= a and b;
    layer3_outputs(2535) <= a xor b;
    layer3_outputs(2536) <= not b;
    layer3_outputs(2537) <= not (a and b);
    layer3_outputs(2538) <= a and not b;
    layer3_outputs(2539) <= b and not a;
    layer3_outputs(2540) <= not a;
    layer3_outputs(2541) <= not b;
    layer3_outputs(2542) <= not (a or b);
    layer3_outputs(2543) <= a and b;
    layer3_outputs(2544) <= not b or a;
    layer3_outputs(2545) <= 1'b0;
    layer3_outputs(2546) <= a xor b;
    layer3_outputs(2547) <= not a or b;
    layer3_outputs(2548) <= a;
    layer3_outputs(2549) <= 1'b0;
    layer3_outputs(2550) <= a and not b;
    layer3_outputs(2551) <= not (a or b);
    layer3_outputs(2552) <= a xor b;
    layer3_outputs(2553) <= a;
    layer3_outputs(2554) <= not b or a;
    layer3_outputs(2555) <= b;
    layer3_outputs(2556) <= not a;
    layer3_outputs(2557) <= not (a and b);
    layer3_outputs(2558) <= a and b;
    layer3_outputs(2559) <= a or b;
    layer4_outputs(0) <= not a or b;
    layer4_outputs(1) <= not b or a;
    layer4_outputs(2) <= a and b;
    layer4_outputs(3) <= not a or b;
    layer4_outputs(4) <= b;
    layer4_outputs(5) <= b;
    layer4_outputs(6) <= not (a and b);
    layer4_outputs(7) <= 1'b1;
    layer4_outputs(8) <= a or b;
    layer4_outputs(9) <= a xor b;
    layer4_outputs(10) <= a and b;
    layer4_outputs(11) <= b;
    layer4_outputs(12) <= not b or a;
    layer4_outputs(13) <= not a;
    layer4_outputs(14) <= b and not a;
    layer4_outputs(15) <= a and not b;
    layer4_outputs(16) <= a;
    layer4_outputs(17) <= not a or b;
    layer4_outputs(18) <= 1'b0;
    layer4_outputs(19) <= not (a and b);
    layer4_outputs(20) <= not a or b;
    layer4_outputs(21) <= not a or b;
    layer4_outputs(22) <= a and not b;
    layer4_outputs(23) <= a or b;
    layer4_outputs(24) <= a and not b;
    layer4_outputs(25) <= 1'b1;
    layer4_outputs(26) <= 1'b0;
    layer4_outputs(27) <= b;
    layer4_outputs(28) <= a;
    layer4_outputs(29) <= 1'b0;
    layer4_outputs(30) <= not (a or b);
    layer4_outputs(31) <= not a or b;
    layer4_outputs(32) <= a;
    layer4_outputs(33) <= not (a or b);
    layer4_outputs(34) <= not (a and b);
    layer4_outputs(35) <= a and b;
    layer4_outputs(36) <= a or b;
    layer4_outputs(37) <= not b or a;
    layer4_outputs(38) <= not (a and b);
    layer4_outputs(39) <= a;
    layer4_outputs(40) <= b and not a;
    layer4_outputs(41) <= not (a or b);
    layer4_outputs(42) <= a;
    layer4_outputs(43) <= b;
    layer4_outputs(44) <= not b;
    layer4_outputs(45) <= not (a and b);
    layer4_outputs(46) <= b;
    layer4_outputs(47) <= b and not a;
    layer4_outputs(48) <= not a or b;
    layer4_outputs(49) <= not a or b;
    layer4_outputs(50) <= a and not b;
    layer4_outputs(51) <= a and b;
    layer4_outputs(52) <= a and b;
    layer4_outputs(53) <= b;
    layer4_outputs(54) <= b;
    layer4_outputs(55) <= not b;
    layer4_outputs(56) <= a xor b;
    layer4_outputs(57) <= a or b;
    layer4_outputs(58) <= not a;
    layer4_outputs(59) <= not a;
    layer4_outputs(60) <= not b;
    layer4_outputs(61) <= b;
    layer4_outputs(62) <= not (a xor b);
    layer4_outputs(63) <= not (a and b);
    layer4_outputs(64) <= a and b;
    layer4_outputs(65) <= a or b;
    layer4_outputs(66) <= a and b;
    layer4_outputs(67) <= not a or b;
    layer4_outputs(68) <= not (a and b);
    layer4_outputs(69) <= not b;
    layer4_outputs(70) <= a;
    layer4_outputs(71) <= b;
    layer4_outputs(72) <= a and not b;
    layer4_outputs(73) <= not b or a;
    layer4_outputs(74) <= not a or b;
    layer4_outputs(75) <= not b;
    layer4_outputs(76) <= a;
    layer4_outputs(77) <= a xor b;
    layer4_outputs(78) <= not (a and b);
    layer4_outputs(79) <= not a or b;
    layer4_outputs(80) <= 1'b0;
    layer4_outputs(81) <= 1'b1;
    layer4_outputs(82) <= not a or b;
    layer4_outputs(83) <= a and not b;
    layer4_outputs(84) <= not a;
    layer4_outputs(85) <= not b;
    layer4_outputs(86) <= 1'b1;
    layer4_outputs(87) <= 1'b1;
    layer4_outputs(88) <= not (a or b);
    layer4_outputs(89) <= not a;
    layer4_outputs(90) <= not (a or b);
    layer4_outputs(91) <= b and not a;
    layer4_outputs(92) <= a and not b;
    layer4_outputs(93) <= b;
    layer4_outputs(94) <= 1'b1;
    layer4_outputs(95) <= not a or b;
    layer4_outputs(96) <= b and not a;
    layer4_outputs(97) <= 1'b1;
    layer4_outputs(98) <= 1'b0;
    layer4_outputs(99) <= not b;
    layer4_outputs(100) <= not (a or b);
    layer4_outputs(101) <= not (a and b);
    layer4_outputs(102) <= not (a and b);
    layer4_outputs(103) <= not a;
    layer4_outputs(104) <= not a or b;
    layer4_outputs(105) <= b;
    layer4_outputs(106) <= not (a or b);
    layer4_outputs(107) <= b and not a;
    layer4_outputs(108) <= not b or a;
    layer4_outputs(109) <= a;
    layer4_outputs(110) <= 1'b1;
    layer4_outputs(111) <= a or b;
    layer4_outputs(112) <= not (a and b);
    layer4_outputs(113) <= a and b;
    layer4_outputs(114) <= not (a or b);
    layer4_outputs(115) <= not b;
    layer4_outputs(116) <= a and b;
    layer4_outputs(117) <= not (a xor b);
    layer4_outputs(118) <= 1'b0;
    layer4_outputs(119) <= a;
    layer4_outputs(120) <= b;
    layer4_outputs(121) <= a and b;
    layer4_outputs(122) <= not a or b;
    layer4_outputs(123) <= a or b;
    layer4_outputs(124) <= not a or b;
    layer4_outputs(125) <= a;
    layer4_outputs(126) <= not a;
    layer4_outputs(127) <= not (a xor b);
    layer4_outputs(128) <= a;
    layer4_outputs(129) <= b and not a;
    layer4_outputs(130) <= not a;
    layer4_outputs(131) <= 1'b0;
    layer4_outputs(132) <= b;
    layer4_outputs(133) <= b;
    layer4_outputs(134) <= not (a or b);
    layer4_outputs(135) <= a;
    layer4_outputs(136) <= not b or a;
    layer4_outputs(137) <= a and b;
    layer4_outputs(138) <= 1'b0;
    layer4_outputs(139) <= not a;
    layer4_outputs(140) <= a or b;
    layer4_outputs(141) <= 1'b1;
    layer4_outputs(142) <= a or b;
    layer4_outputs(143) <= a and b;
    layer4_outputs(144) <= a or b;
    layer4_outputs(145) <= not b or a;
    layer4_outputs(146) <= a and not b;
    layer4_outputs(147) <= a or b;
    layer4_outputs(148) <= a xor b;
    layer4_outputs(149) <= a;
    layer4_outputs(150) <= not b;
    layer4_outputs(151) <= not b;
    layer4_outputs(152) <= a and b;
    layer4_outputs(153) <= a or b;
    layer4_outputs(154) <= 1'b1;
    layer4_outputs(155) <= a and b;
    layer4_outputs(156) <= not a;
    layer4_outputs(157) <= not b;
    layer4_outputs(158) <= not b;
    layer4_outputs(159) <= not a;
    layer4_outputs(160) <= not b or a;
    layer4_outputs(161) <= a and not b;
    layer4_outputs(162) <= not b or a;
    layer4_outputs(163) <= a or b;
    layer4_outputs(164) <= a and not b;
    layer4_outputs(165) <= not b or a;
    layer4_outputs(166) <= 1'b1;
    layer4_outputs(167) <= b and not a;
    layer4_outputs(168) <= a and not b;
    layer4_outputs(169) <= a xor b;
    layer4_outputs(170) <= not a;
    layer4_outputs(171) <= not b;
    layer4_outputs(172) <= not b or a;
    layer4_outputs(173) <= a;
    layer4_outputs(174) <= 1'b0;
    layer4_outputs(175) <= not b;
    layer4_outputs(176) <= not a or b;
    layer4_outputs(177) <= 1'b1;
    layer4_outputs(178) <= 1'b1;
    layer4_outputs(179) <= 1'b0;
    layer4_outputs(180) <= not b or a;
    layer4_outputs(181) <= b;
    layer4_outputs(182) <= b;
    layer4_outputs(183) <= not (a and b);
    layer4_outputs(184) <= b;
    layer4_outputs(185) <= not a or b;
    layer4_outputs(186) <= 1'b0;
    layer4_outputs(187) <= a;
    layer4_outputs(188) <= not a or b;
    layer4_outputs(189) <= not b;
    layer4_outputs(190) <= b and not a;
    layer4_outputs(191) <= 1'b1;
    layer4_outputs(192) <= b and not a;
    layer4_outputs(193) <= not (a or b);
    layer4_outputs(194) <= not b;
    layer4_outputs(195) <= 1'b0;
    layer4_outputs(196) <= 1'b0;
    layer4_outputs(197) <= not b or a;
    layer4_outputs(198) <= not b or a;
    layer4_outputs(199) <= not a or b;
    layer4_outputs(200) <= b and not a;
    layer4_outputs(201) <= a and not b;
    layer4_outputs(202) <= a and not b;
    layer4_outputs(203) <= a and b;
    layer4_outputs(204) <= b and not a;
    layer4_outputs(205) <= not b or a;
    layer4_outputs(206) <= not a;
    layer4_outputs(207) <= b and not a;
    layer4_outputs(208) <= b and not a;
    layer4_outputs(209) <= 1'b0;
    layer4_outputs(210) <= a and b;
    layer4_outputs(211) <= a and not b;
    layer4_outputs(212) <= 1'b0;
    layer4_outputs(213) <= 1'b1;
    layer4_outputs(214) <= not b or a;
    layer4_outputs(215) <= not a;
    layer4_outputs(216) <= 1'b1;
    layer4_outputs(217) <= not (a or b);
    layer4_outputs(218) <= a and not b;
    layer4_outputs(219) <= a;
    layer4_outputs(220) <= a and not b;
    layer4_outputs(221) <= not (a or b);
    layer4_outputs(222) <= b and not a;
    layer4_outputs(223) <= not b;
    layer4_outputs(224) <= not (a and b);
    layer4_outputs(225) <= b;
    layer4_outputs(226) <= a and not b;
    layer4_outputs(227) <= b;
    layer4_outputs(228) <= a and b;
    layer4_outputs(229) <= not a or b;
    layer4_outputs(230) <= not (a xor b);
    layer4_outputs(231) <= a;
    layer4_outputs(232) <= 1'b1;
    layer4_outputs(233) <= b and not a;
    layer4_outputs(234) <= not a;
    layer4_outputs(235) <= not a or b;
    layer4_outputs(236) <= a and not b;
    layer4_outputs(237) <= not b or a;
    layer4_outputs(238) <= a and b;
    layer4_outputs(239) <= not (a xor b);
    layer4_outputs(240) <= a or b;
    layer4_outputs(241) <= b and not a;
    layer4_outputs(242) <= a;
    layer4_outputs(243) <= a or b;
    layer4_outputs(244) <= b and not a;
    layer4_outputs(245) <= not a;
    layer4_outputs(246) <= a;
    layer4_outputs(247) <= not b;
    layer4_outputs(248) <= a;
    layer4_outputs(249) <= a and b;
    layer4_outputs(250) <= a;
    layer4_outputs(251) <= not b or a;
    layer4_outputs(252) <= a;
    layer4_outputs(253) <= b;
    layer4_outputs(254) <= not (a or b);
    layer4_outputs(255) <= not b or a;
    layer4_outputs(256) <= not a or b;
    layer4_outputs(257) <= a;
    layer4_outputs(258) <= b and not a;
    layer4_outputs(259) <= not (a and b);
    layer4_outputs(260) <= not (a and b);
    layer4_outputs(261) <= not a;
    layer4_outputs(262) <= a;
    layer4_outputs(263) <= not b;
    layer4_outputs(264) <= not b;
    layer4_outputs(265) <= not (a and b);
    layer4_outputs(266) <= not (a and b);
    layer4_outputs(267) <= a;
    layer4_outputs(268) <= not (a or b);
    layer4_outputs(269) <= b and not a;
    layer4_outputs(270) <= not a or b;
    layer4_outputs(271) <= b and not a;
    layer4_outputs(272) <= not (a and b);
    layer4_outputs(273) <= a and not b;
    layer4_outputs(274) <= a;
    layer4_outputs(275) <= not b or a;
    layer4_outputs(276) <= not (a xor b);
    layer4_outputs(277) <= a and not b;
    layer4_outputs(278) <= not (a or b);
    layer4_outputs(279) <= 1'b1;
    layer4_outputs(280) <= a xor b;
    layer4_outputs(281) <= 1'b0;
    layer4_outputs(282) <= not (a xor b);
    layer4_outputs(283) <= b;
    layer4_outputs(284) <= not a or b;
    layer4_outputs(285) <= not b or a;
    layer4_outputs(286) <= not a or b;
    layer4_outputs(287) <= not a or b;
    layer4_outputs(288) <= not (a or b);
    layer4_outputs(289) <= a;
    layer4_outputs(290) <= not (a and b);
    layer4_outputs(291) <= not b or a;
    layer4_outputs(292) <= not a;
    layer4_outputs(293) <= a and not b;
    layer4_outputs(294) <= a or b;
    layer4_outputs(295) <= 1'b0;
    layer4_outputs(296) <= not (a or b);
    layer4_outputs(297) <= not a or b;
    layer4_outputs(298) <= not a;
    layer4_outputs(299) <= not a or b;
    layer4_outputs(300) <= a and b;
    layer4_outputs(301) <= not b;
    layer4_outputs(302) <= a and not b;
    layer4_outputs(303) <= a;
    layer4_outputs(304) <= not a;
    layer4_outputs(305) <= 1'b0;
    layer4_outputs(306) <= not a;
    layer4_outputs(307) <= a or b;
    layer4_outputs(308) <= a;
    layer4_outputs(309) <= a or b;
    layer4_outputs(310) <= not a;
    layer4_outputs(311) <= not a or b;
    layer4_outputs(312) <= not b;
    layer4_outputs(313) <= not (a and b);
    layer4_outputs(314) <= not (a and b);
    layer4_outputs(315) <= not (a or b);
    layer4_outputs(316) <= not b or a;
    layer4_outputs(317) <= a or b;
    layer4_outputs(318) <= not a;
    layer4_outputs(319) <= not (a or b);
    layer4_outputs(320) <= b and not a;
    layer4_outputs(321) <= not (a and b);
    layer4_outputs(322) <= not b or a;
    layer4_outputs(323) <= not b;
    layer4_outputs(324) <= 1'b0;
    layer4_outputs(325) <= not a;
    layer4_outputs(326) <= not a;
    layer4_outputs(327) <= a;
    layer4_outputs(328) <= a;
    layer4_outputs(329) <= a;
    layer4_outputs(330) <= b;
    layer4_outputs(331) <= a or b;
    layer4_outputs(332) <= a and not b;
    layer4_outputs(333) <= a and not b;
    layer4_outputs(334) <= a;
    layer4_outputs(335) <= a and not b;
    layer4_outputs(336) <= not a or b;
    layer4_outputs(337) <= not a;
    layer4_outputs(338) <= not (a or b);
    layer4_outputs(339) <= not a;
    layer4_outputs(340) <= not (a or b);
    layer4_outputs(341) <= not a;
    layer4_outputs(342) <= a and not b;
    layer4_outputs(343) <= not a;
    layer4_outputs(344) <= not (a and b);
    layer4_outputs(345) <= not (a and b);
    layer4_outputs(346) <= a and b;
    layer4_outputs(347) <= b;
    layer4_outputs(348) <= not a or b;
    layer4_outputs(349) <= not a or b;
    layer4_outputs(350) <= not a or b;
    layer4_outputs(351) <= a and b;
    layer4_outputs(352) <= 1'b0;
    layer4_outputs(353) <= not a;
    layer4_outputs(354) <= b;
    layer4_outputs(355) <= not a or b;
    layer4_outputs(356) <= b;
    layer4_outputs(357) <= a and b;
    layer4_outputs(358) <= not a;
    layer4_outputs(359) <= a or b;
    layer4_outputs(360) <= b and not a;
    layer4_outputs(361) <= not (a or b);
    layer4_outputs(362) <= not (a and b);
    layer4_outputs(363) <= a and b;
    layer4_outputs(364) <= not a or b;
    layer4_outputs(365) <= not a;
    layer4_outputs(366) <= 1'b1;
    layer4_outputs(367) <= a and b;
    layer4_outputs(368) <= not (a or b);
    layer4_outputs(369) <= a and not b;
    layer4_outputs(370) <= not b;
    layer4_outputs(371) <= a;
    layer4_outputs(372) <= b and not a;
    layer4_outputs(373) <= a or b;
    layer4_outputs(374) <= not a;
    layer4_outputs(375) <= not b or a;
    layer4_outputs(376) <= a and b;
    layer4_outputs(377) <= a or b;
    layer4_outputs(378) <= a and b;
    layer4_outputs(379) <= a;
    layer4_outputs(380) <= not b;
    layer4_outputs(381) <= not (a and b);
    layer4_outputs(382) <= 1'b1;
    layer4_outputs(383) <= 1'b1;
    layer4_outputs(384) <= 1'b1;
    layer4_outputs(385) <= b and not a;
    layer4_outputs(386) <= not b;
    layer4_outputs(387) <= 1'b0;
    layer4_outputs(388) <= not (a or b);
    layer4_outputs(389) <= not a;
    layer4_outputs(390) <= a and b;
    layer4_outputs(391) <= 1'b1;
    layer4_outputs(392) <= not b;
    layer4_outputs(393) <= a;
    layer4_outputs(394) <= not b or a;
    layer4_outputs(395) <= not (a and b);
    layer4_outputs(396) <= a and not b;
    layer4_outputs(397) <= not b;
    layer4_outputs(398) <= not (a and b);
    layer4_outputs(399) <= not (a and b);
    layer4_outputs(400) <= a and b;
    layer4_outputs(401) <= not (a or b);
    layer4_outputs(402) <= b and not a;
    layer4_outputs(403) <= not (a and b);
    layer4_outputs(404) <= 1'b1;
    layer4_outputs(405) <= not a or b;
    layer4_outputs(406) <= a xor b;
    layer4_outputs(407) <= not (a and b);
    layer4_outputs(408) <= 1'b0;
    layer4_outputs(409) <= 1'b0;
    layer4_outputs(410) <= b and not a;
    layer4_outputs(411) <= not b;
    layer4_outputs(412) <= a or b;
    layer4_outputs(413) <= not b or a;
    layer4_outputs(414) <= b and not a;
    layer4_outputs(415) <= not b;
    layer4_outputs(416) <= not (a and b);
    layer4_outputs(417) <= a;
    layer4_outputs(418) <= 1'b1;
    layer4_outputs(419) <= not a or b;
    layer4_outputs(420) <= not b or a;
    layer4_outputs(421) <= not (a or b);
    layer4_outputs(422) <= a xor b;
    layer4_outputs(423) <= 1'b1;
    layer4_outputs(424) <= b;
    layer4_outputs(425) <= not (a and b);
    layer4_outputs(426) <= not a;
    layer4_outputs(427) <= not b or a;
    layer4_outputs(428) <= not b;
    layer4_outputs(429) <= not b or a;
    layer4_outputs(430) <= not b or a;
    layer4_outputs(431) <= not (a or b);
    layer4_outputs(432) <= a and b;
    layer4_outputs(433) <= a;
    layer4_outputs(434) <= 1'b0;
    layer4_outputs(435) <= b and not a;
    layer4_outputs(436) <= not b or a;
    layer4_outputs(437) <= not b;
    layer4_outputs(438) <= not b;
    layer4_outputs(439) <= a and not b;
    layer4_outputs(440) <= a and not b;
    layer4_outputs(441) <= 1'b0;
    layer4_outputs(442) <= b;
    layer4_outputs(443) <= 1'b0;
    layer4_outputs(444) <= not (a xor b);
    layer4_outputs(445) <= not (a or b);
    layer4_outputs(446) <= not a or b;
    layer4_outputs(447) <= a or b;
    layer4_outputs(448) <= 1'b1;
    layer4_outputs(449) <= not b;
    layer4_outputs(450) <= b and not a;
    layer4_outputs(451) <= not (a or b);
    layer4_outputs(452) <= a and b;
    layer4_outputs(453) <= not (a or b);
    layer4_outputs(454) <= not b;
    layer4_outputs(455) <= a and b;
    layer4_outputs(456) <= a and b;
    layer4_outputs(457) <= not (a and b);
    layer4_outputs(458) <= not (a or b);
    layer4_outputs(459) <= a and not b;
    layer4_outputs(460) <= not a;
    layer4_outputs(461) <= not (a or b);
    layer4_outputs(462) <= a or b;
    layer4_outputs(463) <= a and not b;
    layer4_outputs(464) <= 1'b1;
    layer4_outputs(465) <= 1'b1;
    layer4_outputs(466) <= not b;
    layer4_outputs(467) <= a and not b;
    layer4_outputs(468) <= not (a or b);
    layer4_outputs(469) <= a and b;
    layer4_outputs(470) <= 1'b1;
    layer4_outputs(471) <= b and not a;
    layer4_outputs(472) <= a and not b;
    layer4_outputs(473) <= not b;
    layer4_outputs(474) <= not a or b;
    layer4_outputs(475) <= b;
    layer4_outputs(476) <= 1'b0;
    layer4_outputs(477) <= not a;
    layer4_outputs(478) <= a and not b;
    layer4_outputs(479) <= not b or a;
    layer4_outputs(480) <= a and b;
    layer4_outputs(481) <= b;
    layer4_outputs(482) <= a and not b;
    layer4_outputs(483) <= a and b;
    layer4_outputs(484) <= a and b;
    layer4_outputs(485) <= a or b;
    layer4_outputs(486) <= a and not b;
    layer4_outputs(487) <= 1'b1;
    layer4_outputs(488) <= b and not a;
    layer4_outputs(489) <= 1'b1;
    layer4_outputs(490) <= not a or b;
    layer4_outputs(491) <= a and b;
    layer4_outputs(492) <= not (a or b);
    layer4_outputs(493) <= b;
    layer4_outputs(494) <= not (a or b);
    layer4_outputs(495) <= a;
    layer4_outputs(496) <= not (a or b);
    layer4_outputs(497) <= b;
    layer4_outputs(498) <= not a;
    layer4_outputs(499) <= not b or a;
    layer4_outputs(500) <= 1'b1;
    layer4_outputs(501) <= not a;
    layer4_outputs(502) <= b and not a;
    layer4_outputs(503) <= not b;
    layer4_outputs(504) <= not (a or b);
    layer4_outputs(505) <= a or b;
    layer4_outputs(506) <= b;
    layer4_outputs(507) <= not b;
    layer4_outputs(508) <= a;
    layer4_outputs(509) <= not b;
    layer4_outputs(510) <= 1'b1;
    layer4_outputs(511) <= b;
    layer4_outputs(512) <= b and not a;
    layer4_outputs(513) <= not b or a;
    layer4_outputs(514) <= 1'b1;
    layer4_outputs(515) <= 1'b1;
    layer4_outputs(516) <= 1'b1;
    layer4_outputs(517) <= not (a or b);
    layer4_outputs(518) <= b;
    layer4_outputs(519) <= not b or a;
    layer4_outputs(520) <= a;
    layer4_outputs(521) <= 1'b1;
    layer4_outputs(522) <= not (a or b);
    layer4_outputs(523) <= not (a and b);
    layer4_outputs(524) <= b and not a;
    layer4_outputs(525) <= 1'b0;
    layer4_outputs(526) <= a or b;
    layer4_outputs(527) <= not b or a;
    layer4_outputs(528) <= b;
    layer4_outputs(529) <= a and not b;
    layer4_outputs(530) <= not b or a;
    layer4_outputs(531) <= not (a and b);
    layer4_outputs(532) <= a and not b;
    layer4_outputs(533) <= a or b;
    layer4_outputs(534) <= not b;
    layer4_outputs(535) <= b and not a;
    layer4_outputs(536) <= not b;
    layer4_outputs(537) <= 1'b0;
    layer4_outputs(538) <= not b or a;
    layer4_outputs(539) <= not b;
    layer4_outputs(540) <= 1'b1;
    layer4_outputs(541) <= 1'b0;
    layer4_outputs(542) <= not b;
    layer4_outputs(543) <= b;
    layer4_outputs(544) <= not (a and b);
    layer4_outputs(545) <= a and b;
    layer4_outputs(546) <= a and b;
    layer4_outputs(547) <= a;
    layer4_outputs(548) <= not a;
    layer4_outputs(549) <= not (a xor b);
    layer4_outputs(550) <= not b;
    layer4_outputs(551) <= b;
    layer4_outputs(552) <= a and b;
    layer4_outputs(553) <= 1'b1;
    layer4_outputs(554) <= a;
    layer4_outputs(555) <= not b or a;
    layer4_outputs(556) <= a or b;
    layer4_outputs(557) <= a and not b;
    layer4_outputs(558) <= a xor b;
    layer4_outputs(559) <= a xor b;
    layer4_outputs(560) <= a and not b;
    layer4_outputs(561) <= a;
    layer4_outputs(562) <= not b;
    layer4_outputs(563) <= not a;
    layer4_outputs(564) <= 1'b0;
    layer4_outputs(565) <= a and not b;
    layer4_outputs(566) <= a and not b;
    layer4_outputs(567) <= a or b;
    layer4_outputs(568) <= not (a and b);
    layer4_outputs(569) <= not b or a;
    layer4_outputs(570) <= b and not a;
    layer4_outputs(571) <= a and not b;
    layer4_outputs(572) <= not a;
    layer4_outputs(573) <= b;
    layer4_outputs(574) <= not a;
    layer4_outputs(575) <= not b or a;
    layer4_outputs(576) <= not b or a;
    layer4_outputs(577) <= not b or a;
    layer4_outputs(578) <= not a or b;
    layer4_outputs(579) <= a and not b;
    layer4_outputs(580) <= not (a xor b);
    layer4_outputs(581) <= a and b;
    layer4_outputs(582) <= not a;
    layer4_outputs(583) <= not b or a;
    layer4_outputs(584) <= not b or a;
    layer4_outputs(585) <= not b or a;
    layer4_outputs(586) <= b;
    layer4_outputs(587) <= a and b;
    layer4_outputs(588) <= a and not b;
    layer4_outputs(589) <= not b or a;
    layer4_outputs(590) <= a and b;
    layer4_outputs(591) <= a or b;
    layer4_outputs(592) <= not a or b;
    layer4_outputs(593) <= a and b;
    layer4_outputs(594) <= a xor b;
    layer4_outputs(595) <= a or b;
    layer4_outputs(596) <= a;
    layer4_outputs(597) <= not b or a;
    layer4_outputs(598) <= not a or b;
    layer4_outputs(599) <= not a or b;
    layer4_outputs(600) <= not a or b;
    layer4_outputs(601) <= not (a and b);
    layer4_outputs(602) <= not (a and b);
    layer4_outputs(603) <= 1'b1;
    layer4_outputs(604) <= b;
    layer4_outputs(605) <= not b or a;
    layer4_outputs(606) <= a and b;
    layer4_outputs(607) <= a and not b;
    layer4_outputs(608) <= not a;
    layer4_outputs(609) <= not a;
    layer4_outputs(610) <= 1'b1;
    layer4_outputs(611) <= not b;
    layer4_outputs(612) <= not (a and b);
    layer4_outputs(613) <= not b or a;
    layer4_outputs(614) <= b and not a;
    layer4_outputs(615) <= a and not b;
    layer4_outputs(616) <= not a or b;
    layer4_outputs(617) <= 1'b1;
    layer4_outputs(618) <= not b or a;
    layer4_outputs(619) <= a and not b;
    layer4_outputs(620) <= b and not a;
    layer4_outputs(621) <= 1'b0;
    layer4_outputs(622) <= a and b;
    layer4_outputs(623) <= b;
    layer4_outputs(624) <= not b or a;
    layer4_outputs(625) <= 1'b0;
    layer4_outputs(626) <= a and not b;
    layer4_outputs(627) <= a and b;
    layer4_outputs(628) <= not a or b;
    layer4_outputs(629) <= a or b;
    layer4_outputs(630) <= 1'b1;
    layer4_outputs(631) <= not a or b;
    layer4_outputs(632) <= not a;
    layer4_outputs(633) <= not a or b;
    layer4_outputs(634) <= a and not b;
    layer4_outputs(635) <= a;
    layer4_outputs(636) <= b;
    layer4_outputs(637) <= b;
    layer4_outputs(638) <= not a or b;
    layer4_outputs(639) <= not a;
    layer4_outputs(640) <= not b;
    layer4_outputs(641) <= a or b;
    layer4_outputs(642) <= not b or a;
    layer4_outputs(643) <= not b or a;
    layer4_outputs(644) <= not (a or b);
    layer4_outputs(645) <= not (a and b);
    layer4_outputs(646) <= a;
    layer4_outputs(647) <= a;
    layer4_outputs(648) <= a or b;
    layer4_outputs(649) <= 1'b0;
    layer4_outputs(650) <= 1'b1;
    layer4_outputs(651) <= a and not b;
    layer4_outputs(652) <= a and not b;
    layer4_outputs(653) <= a and not b;
    layer4_outputs(654) <= a;
    layer4_outputs(655) <= 1'b1;
    layer4_outputs(656) <= not a;
    layer4_outputs(657) <= not (a xor b);
    layer4_outputs(658) <= not b;
    layer4_outputs(659) <= not (a and b);
    layer4_outputs(660) <= b and not a;
    layer4_outputs(661) <= not (a or b);
    layer4_outputs(662) <= 1'b0;
    layer4_outputs(663) <= a;
    layer4_outputs(664) <= not b or a;
    layer4_outputs(665) <= a or b;
    layer4_outputs(666) <= a;
    layer4_outputs(667) <= 1'b0;
    layer4_outputs(668) <= a and b;
    layer4_outputs(669) <= a and not b;
    layer4_outputs(670) <= not (a and b);
    layer4_outputs(671) <= not b or a;
    layer4_outputs(672) <= b;
    layer4_outputs(673) <= not b;
    layer4_outputs(674) <= not b;
    layer4_outputs(675) <= not (a or b);
    layer4_outputs(676) <= b;
    layer4_outputs(677) <= not b or a;
    layer4_outputs(678) <= a and not b;
    layer4_outputs(679) <= 1'b1;
    layer4_outputs(680) <= not b or a;
    layer4_outputs(681) <= not (a and b);
    layer4_outputs(682) <= b;
    layer4_outputs(683) <= 1'b1;
    layer4_outputs(684) <= not (a or b);
    layer4_outputs(685) <= 1'b0;
    layer4_outputs(686) <= a;
    layer4_outputs(687) <= not a or b;
    layer4_outputs(688) <= a and b;
    layer4_outputs(689) <= a and not b;
    layer4_outputs(690) <= not (a or b);
    layer4_outputs(691) <= not a;
    layer4_outputs(692) <= not a;
    layer4_outputs(693) <= b and not a;
    layer4_outputs(694) <= not (a xor b);
    layer4_outputs(695) <= not (a or b);
    layer4_outputs(696) <= 1'b0;
    layer4_outputs(697) <= 1'b1;
    layer4_outputs(698) <= not (a or b);
    layer4_outputs(699) <= 1'b1;
    layer4_outputs(700) <= 1'b1;
    layer4_outputs(701) <= a or b;
    layer4_outputs(702) <= a;
    layer4_outputs(703) <= not b or a;
    layer4_outputs(704) <= a;
    layer4_outputs(705) <= a;
    layer4_outputs(706) <= b;
    layer4_outputs(707) <= not a;
    layer4_outputs(708) <= not b or a;
    layer4_outputs(709) <= b and not a;
    layer4_outputs(710) <= not b or a;
    layer4_outputs(711) <= 1'b0;
    layer4_outputs(712) <= a;
    layer4_outputs(713) <= b;
    layer4_outputs(714) <= not a;
    layer4_outputs(715) <= 1'b0;
    layer4_outputs(716) <= not a or b;
    layer4_outputs(717) <= a and not b;
    layer4_outputs(718) <= 1'b0;
    layer4_outputs(719) <= b and not a;
    layer4_outputs(720) <= not a;
    layer4_outputs(721) <= a and b;
    layer4_outputs(722) <= 1'b1;
    layer4_outputs(723) <= not a;
    layer4_outputs(724) <= b and not a;
    layer4_outputs(725) <= b and not a;
    layer4_outputs(726) <= a or b;
    layer4_outputs(727) <= a and not b;
    layer4_outputs(728) <= 1'b1;
    layer4_outputs(729) <= not a or b;
    layer4_outputs(730) <= a and b;
    layer4_outputs(731) <= not b or a;
    layer4_outputs(732) <= a or b;
    layer4_outputs(733) <= a and not b;
    layer4_outputs(734) <= a;
    layer4_outputs(735) <= not a or b;
    layer4_outputs(736) <= 1'b1;
    layer4_outputs(737) <= not b;
    layer4_outputs(738) <= b;
    layer4_outputs(739) <= 1'b1;
    layer4_outputs(740) <= not a or b;
    layer4_outputs(741) <= not a;
    layer4_outputs(742) <= a and not b;
    layer4_outputs(743) <= a;
    layer4_outputs(744) <= not a;
    layer4_outputs(745) <= not a;
    layer4_outputs(746) <= not b;
    layer4_outputs(747) <= b and not a;
    layer4_outputs(748) <= not (a and b);
    layer4_outputs(749) <= not (a and b);
    layer4_outputs(750) <= not b or a;
    layer4_outputs(751) <= not b or a;
    layer4_outputs(752) <= a and not b;
    layer4_outputs(753) <= b and not a;
    layer4_outputs(754) <= b;
    layer4_outputs(755) <= not (a xor b);
    layer4_outputs(756) <= b;
    layer4_outputs(757) <= not (a or b);
    layer4_outputs(758) <= a;
    layer4_outputs(759) <= a or b;
    layer4_outputs(760) <= a;
    layer4_outputs(761) <= a and not b;
    layer4_outputs(762) <= a and not b;
    layer4_outputs(763) <= b;
    layer4_outputs(764) <= a or b;
    layer4_outputs(765) <= not (a xor b);
    layer4_outputs(766) <= not a;
    layer4_outputs(767) <= not (a and b);
    layer4_outputs(768) <= 1'b1;
    layer4_outputs(769) <= a xor b;
    layer4_outputs(770) <= b;
    layer4_outputs(771) <= b;
    layer4_outputs(772) <= a or b;
    layer4_outputs(773) <= not a or b;
    layer4_outputs(774) <= a and not b;
    layer4_outputs(775) <= a xor b;
    layer4_outputs(776) <= a;
    layer4_outputs(777) <= b;
    layer4_outputs(778) <= a and not b;
    layer4_outputs(779) <= not (a and b);
    layer4_outputs(780) <= not a or b;
    layer4_outputs(781) <= a and not b;
    layer4_outputs(782) <= not b or a;
    layer4_outputs(783) <= not b;
    layer4_outputs(784) <= a or b;
    layer4_outputs(785) <= not b;
    layer4_outputs(786) <= not b;
    layer4_outputs(787) <= a xor b;
    layer4_outputs(788) <= a and b;
    layer4_outputs(789) <= a;
    layer4_outputs(790) <= 1'b1;
    layer4_outputs(791) <= b;
    layer4_outputs(792) <= not (a or b);
    layer4_outputs(793) <= a and not b;
    layer4_outputs(794) <= b and not a;
    layer4_outputs(795) <= not (a xor b);
    layer4_outputs(796) <= a;
    layer4_outputs(797) <= not b;
    layer4_outputs(798) <= not b;
    layer4_outputs(799) <= 1'b1;
    layer4_outputs(800) <= a or b;
    layer4_outputs(801) <= not (a or b);
    layer4_outputs(802) <= not (a or b);
    layer4_outputs(803) <= a xor b;
    layer4_outputs(804) <= a;
    layer4_outputs(805) <= a and not b;
    layer4_outputs(806) <= b;
    layer4_outputs(807) <= b;
    layer4_outputs(808) <= a and b;
    layer4_outputs(809) <= not (a and b);
    layer4_outputs(810) <= a or b;
    layer4_outputs(811) <= 1'b0;
    layer4_outputs(812) <= not b or a;
    layer4_outputs(813) <= 1'b1;
    layer4_outputs(814) <= 1'b0;
    layer4_outputs(815) <= a;
    layer4_outputs(816) <= not b;
    layer4_outputs(817) <= not b or a;
    layer4_outputs(818) <= not b or a;
    layer4_outputs(819) <= 1'b0;
    layer4_outputs(820) <= a and not b;
    layer4_outputs(821) <= not (a or b);
    layer4_outputs(822) <= not a or b;
    layer4_outputs(823) <= b;
    layer4_outputs(824) <= b and not a;
    layer4_outputs(825) <= 1'b1;
    layer4_outputs(826) <= a or b;
    layer4_outputs(827) <= b;
    layer4_outputs(828) <= not b;
    layer4_outputs(829) <= 1'b0;
    layer4_outputs(830) <= not (a and b);
    layer4_outputs(831) <= not (a and b);
    layer4_outputs(832) <= a;
    layer4_outputs(833) <= a or b;
    layer4_outputs(834) <= not b;
    layer4_outputs(835) <= not a;
    layer4_outputs(836) <= not b;
    layer4_outputs(837) <= not (a and b);
    layer4_outputs(838) <= a or b;
    layer4_outputs(839) <= not a or b;
    layer4_outputs(840) <= not a;
    layer4_outputs(841) <= not a or b;
    layer4_outputs(842) <= not (a and b);
    layer4_outputs(843) <= not b or a;
    layer4_outputs(844) <= b and not a;
    layer4_outputs(845) <= b;
    layer4_outputs(846) <= b and not a;
    layer4_outputs(847) <= not (a and b);
    layer4_outputs(848) <= not b or a;
    layer4_outputs(849) <= a and not b;
    layer4_outputs(850) <= 1'b0;
    layer4_outputs(851) <= not a;
    layer4_outputs(852) <= b;
    layer4_outputs(853) <= 1'b1;
    layer4_outputs(854) <= b and not a;
    layer4_outputs(855) <= b and not a;
    layer4_outputs(856) <= a and not b;
    layer4_outputs(857) <= not b or a;
    layer4_outputs(858) <= not (a or b);
    layer4_outputs(859) <= b;
    layer4_outputs(860) <= a and b;
    layer4_outputs(861) <= a xor b;
    layer4_outputs(862) <= a or b;
    layer4_outputs(863) <= not (a or b);
    layer4_outputs(864) <= not b or a;
    layer4_outputs(865) <= a and b;
    layer4_outputs(866) <= a;
    layer4_outputs(867) <= a and b;
    layer4_outputs(868) <= b;
    layer4_outputs(869) <= 1'b0;
    layer4_outputs(870) <= not b or a;
    layer4_outputs(871) <= not a;
    layer4_outputs(872) <= a and b;
    layer4_outputs(873) <= not a;
    layer4_outputs(874) <= b and not a;
    layer4_outputs(875) <= b and not a;
    layer4_outputs(876) <= not a or b;
    layer4_outputs(877) <= a;
    layer4_outputs(878) <= not (a and b);
    layer4_outputs(879) <= 1'b1;
    layer4_outputs(880) <= a and not b;
    layer4_outputs(881) <= not b;
    layer4_outputs(882) <= b and not a;
    layer4_outputs(883) <= 1'b0;
    layer4_outputs(884) <= not (a and b);
    layer4_outputs(885) <= b;
    layer4_outputs(886) <= b;
    layer4_outputs(887) <= 1'b0;
    layer4_outputs(888) <= not a;
    layer4_outputs(889) <= b and not a;
    layer4_outputs(890) <= a and not b;
    layer4_outputs(891) <= not a or b;
    layer4_outputs(892) <= a and not b;
    layer4_outputs(893) <= a;
    layer4_outputs(894) <= not b;
    layer4_outputs(895) <= b;
    layer4_outputs(896) <= not b;
    layer4_outputs(897) <= b and not a;
    layer4_outputs(898) <= 1'b0;
    layer4_outputs(899) <= not a or b;
    layer4_outputs(900) <= not b or a;
    layer4_outputs(901) <= a;
    layer4_outputs(902) <= not b or a;
    layer4_outputs(903) <= 1'b0;
    layer4_outputs(904) <= not b or a;
    layer4_outputs(905) <= a xor b;
    layer4_outputs(906) <= not b or a;
    layer4_outputs(907) <= not (a and b);
    layer4_outputs(908) <= a and not b;
    layer4_outputs(909) <= a;
    layer4_outputs(910) <= a or b;
    layer4_outputs(911) <= a and b;
    layer4_outputs(912) <= 1'b0;
    layer4_outputs(913) <= 1'b0;
    layer4_outputs(914) <= not (a and b);
    layer4_outputs(915) <= a;
    layer4_outputs(916) <= a or b;
    layer4_outputs(917) <= 1'b1;
    layer4_outputs(918) <= a xor b;
    layer4_outputs(919) <= a or b;
    layer4_outputs(920) <= a;
    layer4_outputs(921) <= not b or a;
    layer4_outputs(922) <= not b or a;
    layer4_outputs(923) <= not a;
    layer4_outputs(924) <= not b;
    layer4_outputs(925) <= a and not b;
    layer4_outputs(926) <= b and not a;
    layer4_outputs(927) <= not (a and b);
    layer4_outputs(928) <= a and b;
    layer4_outputs(929) <= a;
    layer4_outputs(930) <= a or b;
    layer4_outputs(931) <= not (a and b);
    layer4_outputs(932) <= not (a or b);
    layer4_outputs(933) <= a;
    layer4_outputs(934) <= not (a and b);
    layer4_outputs(935) <= not (a and b);
    layer4_outputs(936) <= b and not a;
    layer4_outputs(937) <= a or b;
    layer4_outputs(938) <= a;
    layer4_outputs(939) <= 1'b0;
    layer4_outputs(940) <= b;
    layer4_outputs(941) <= 1'b0;
    layer4_outputs(942) <= 1'b0;
    layer4_outputs(943) <= a or b;
    layer4_outputs(944) <= b;
    layer4_outputs(945) <= a and not b;
    layer4_outputs(946) <= a;
    layer4_outputs(947) <= a or b;
    layer4_outputs(948) <= a and not b;
    layer4_outputs(949) <= not b or a;
    layer4_outputs(950) <= a or b;
    layer4_outputs(951) <= not (a or b);
    layer4_outputs(952) <= a and not b;
    layer4_outputs(953) <= not a or b;
    layer4_outputs(954) <= not a;
    layer4_outputs(955) <= a and b;
    layer4_outputs(956) <= not a;
    layer4_outputs(957) <= a and not b;
    layer4_outputs(958) <= a and b;
    layer4_outputs(959) <= not b or a;
    layer4_outputs(960) <= 1'b1;
    layer4_outputs(961) <= not a;
    layer4_outputs(962) <= not (a and b);
    layer4_outputs(963) <= 1'b1;
    layer4_outputs(964) <= not (a or b);
    layer4_outputs(965) <= a and not b;
    layer4_outputs(966) <= not (a or b);
    layer4_outputs(967) <= a and b;
    layer4_outputs(968) <= a;
    layer4_outputs(969) <= not a;
    layer4_outputs(970) <= not (a xor b);
    layer4_outputs(971) <= a;
    layer4_outputs(972) <= a and b;
    layer4_outputs(973) <= a and b;
    layer4_outputs(974) <= not (a or b);
    layer4_outputs(975) <= a;
    layer4_outputs(976) <= not (a and b);
    layer4_outputs(977) <= not a or b;
    layer4_outputs(978) <= not b;
    layer4_outputs(979) <= a;
    layer4_outputs(980) <= 1'b1;
    layer4_outputs(981) <= a xor b;
    layer4_outputs(982) <= b and not a;
    layer4_outputs(983) <= b;
    layer4_outputs(984) <= b and not a;
    layer4_outputs(985) <= 1'b1;
    layer4_outputs(986) <= b;
    layer4_outputs(987) <= 1'b0;
    layer4_outputs(988) <= not a;
    layer4_outputs(989) <= 1'b1;
    layer4_outputs(990) <= a or b;
    layer4_outputs(991) <= b and not a;
    layer4_outputs(992) <= not a;
    layer4_outputs(993) <= not (a or b);
    layer4_outputs(994) <= 1'b1;
    layer4_outputs(995) <= not (a xor b);
    layer4_outputs(996) <= a and not b;
    layer4_outputs(997) <= a xor b;
    layer4_outputs(998) <= 1'b1;
    layer4_outputs(999) <= not (a or b);
    layer4_outputs(1000) <= a or b;
    layer4_outputs(1001) <= not (a and b);
    layer4_outputs(1002) <= a and not b;
    layer4_outputs(1003) <= a xor b;
    layer4_outputs(1004) <= not b or a;
    layer4_outputs(1005) <= not (a and b);
    layer4_outputs(1006) <= not b;
    layer4_outputs(1007) <= not a or b;
    layer4_outputs(1008) <= a;
    layer4_outputs(1009) <= a xor b;
    layer4_outputs(1010) <= not b;
    layer4_outputs(1011) <= a;
    layer4_outputs(1012) <= a and not b;
    layer4_outputs(1013) <= not a or b;
    layer4_outputs(1014) <= a and b;
    layer4_outputs(1015) <= 1'b1;
    layer4_outputs(1016) <= not a;
    layer4_outputs(1017) <= b and not a;
    layer4_outputs(1018) <= a and not b;
    layer4_outputs(1019) <= 1'b0;
    layer4_outputs(1020) <= a and not b;
    layer4_outputs(1021) <= a or b;
    layer4_outputs(1022) <= not b or a;
    layer4_outputs(1023) <= b and not a;
    layer4_outputs(1024) <= a or b;
    layer4_outputs(1025) <= b;
    layer4_outputs(1026) <= not b or a;
    layer4_outputs(1027) <= a;
    layer4_outputs(1028) <= not (a or b);
    layer4_outputs(1029) <= not b;
    layer4_outputs(1030) <= a;
    layer4_outputs(1031) <= a and not b;
    layer4_outputs(1032) <= a and not b;
    layer4_outputs(1033) <= not b or a;
    layer4_outputs(1034) <= not a;
    layer4_outputs(1035) <= 1'b1;
    layer4_outputs(1036) <= 1'b0;
    layer4_outputs(1037) <= a and not b;
    layer4_outputs(1038) <= b and not a;
    layer4_outputs(1039) <= not a;
    layer4_outputs(1040) <= not (a or b);
    layer4_outputs(1041) <= a and not b;
    layer4_outputs(1042) <= not a or b;
    layer4_outputs(1043) <= not b;
    layer4_outputs(1044) <= not (a and b);
    layer4_outputs(1045) <= a and not b;
    layer4_outputs(1046) <= not a or b;
    layer4_outputs(1047) <= 1'b1;
    layer4_outputs(1048) <= b and not a;
    layer4_outputs(1049) <= a and not b;
    layer4_outputs(1050) <= b;
    layer4_outputs(1051) <= not a or b;
    layer4_outputs(1052) <= b;
    layer4_outputs(1053) <= a and not b;
    layer4_outputs(1054) <= not b;
    layer4_outputs(1055) <= 1'b0;
    layer4_outputs(1056) <= a and b;
    layer4_outputs(1057) <= not (a xor b);
    layer4_outputs(1058) <= 1'b1;
    layer4_outputs(1059) <= b and not a;
    layer4_outputs(1060) <= 1'b0;
    layer4_outputs(1061) <= not b;
    layer4_outputs(1062) <= not b or a;
    layer4_outputs(1063) <= not (a or b);
    layer4_outputs(1064) <= not a or b;
    layer4_outputs(1065) <= not (a or b);
    layer4_outputs(1066) <= not b or a;
    layer4_outputs(1067) <= 1'b0;
    layer4_outputs(1068) <= a and b;
    layer4_outputs(1069) <= not b or a;
    layer4_outputs(1070) <= 1'b0;
    layer4_outputs(1071) <= a and not b;
    layer4_outputs(1072) <= 1'b0;
    layer4_outputs(1073) <= not (a or b);
    layer4_outputs(1074) <= not b or a;
    layer4_outputs(1075) <= a or b;
    layer4_outputs(1076) <= not a or b;
    layer4_outputs(1077) <= 1'b1;
    layer4_outputs(1078) <= b and not a;
    layer4_outputs(1079) <= not a;
    layer4_outputs(1080) <= not b or a;
    layer4_outputs(1081) <= a;
    layer4_outputs(1082) <= not (a xor b);
    layer4_outputs(1083) <= not (a and b);
    layer4_outputs(1084) <= not (a and b);
    layer4_outputs(1085) <= a;
    layer4_outputs(1086) <= a and not b;
    layer4_outputs(1087) <= not b;
    layer4_outputs(1088) <= a and not b;
    layer4_outputs(1089) <= b;
    layer4_outputs(1090) <= b and not a;
    layer4_outputs(1091) <= b;
    layer4_outputs(1092) <= a and b;
    layer4_outputs(1093) <= 1'b0;
    layer4_outputs(1094) <= not b;
    layer4_outputs(1095) <= not (a and b);
    layer4_outputs(1096) <= b and not a;
    layer4_outputs(1097) <= b and not a;
    layer4_outputs(1098) <= 1'b1;
    layer4_outputs(1099) <= not a;
    layer4_outputs(1100) <= a or b;
    layer4_outputs(1101) <= 1'b0;
    layer4_outputs(1102) <= not b;
    layer4_outputs(1103) <= b;
    layer4_outputs(1104) <= not a;
    layer4_outputs(1105) <= a;
    layer4_outputs(1106) <= not a or b;
    layer4_outputs(1107) <= a;
    layer4_outputs(1108) <= 1'b1;
    layer4_outputs(1109) <= not b or a;
    layer4_outputs(1110) <= a;
    layer4_outputs(1111) <= a or b;
    layer4_outputs(1112) <= not (a and b);
    layer4_outputs(1113) <= a and b;
    layer4_outputs(1114) <= not b;
    layer4_outputs(1115) <= a or b;
    layer4_outputs(1116) <= 1'b0;
    layer4_outputs(1117) <= not (a or b);
    layer4_outputs(1118) <= not a or b;
    layer4_outputs(1119) <= not a or b;
    layer4_outputs(1120) <= not (a and b);
    layer4_outputs(1121) <= b;
    layer4_outputs(1122) <= not b or a;
    layer4_outputs(1123) <= 1'b1;
    layer4_outputs(1124) <= a and b;
    layer4_outputs(1125) <= not a or b;
    layer4_outputs(1126) <= not b;
    layer4_outputs(1127) <= not b;
    layer4_outputs(1128) <= 1'b1;
    layer4_outputs(1129) <= a;
    layer4_outputs(1130) <= 1'b0;
    layer4_outputs(1131) <= 1'b0;
    layer4_outputs(1132) <= not a or b;
    layer4_outputs(1133) <= b;
    layer4_outputs(1134) <= b;
    layer4_outputs(1135) <= a or b;
    layer4_outputs(1136) <= not (a or b);
    layer4_outputs(1137) <= not (a or b);
    layer4_outputs(1138) <= a or b;
    layer4_outputs(1139) <= not (a xor b);
    layer4_outputs(1140) <= not a or b;
    layer4_outputs(1141) <= not b or a;
    layer4_outputs(1142) <= 1'b0;
    layer4_outputs(1143) <= b;
    layer4_outputs(1144) <= a;
    layer4_outputs(1145) <= not a;
    layer4_outputs(1146) <= not (a and b);
    layer4_outputs(1147) <= 1'b1;
    layer4_outputs(1148) <= not (a or b);
    layer4_outputs(1149) <= not (a and b);
    layer4_outputs(1150) <= not (a or b);
    layer4_outputs(1151) <= a or b;
    layer4_outputs(1152) <= a or b;
    layer4_outputs(1153) <= a;
    layer4_outputs(1154) <= a and not b;
    layer4_outputs(1155) <= not a or b;
    layer4_outputs(1156) <= 1'b0;
    layer4_outputs(1157) <= a or b;
    layer4_outputs(1158) <= a and not b;
    layer4_outputs(1159) <= a;
    layer4_outputs(1160) <= not (a and b);
    layer4_outputs(1161) <= not (a and b);
    layer4_outputs(1162) <= a;
    layer4_outputs(1163) <= not a;
    layer4_outputs(1164) <= 1'b1;
    layer4_outputs(1165) <= 1'b1;
    layer4_outputs(1166) <= not b or a;
    layer4_outputs(1167) <= not (a or b);
    layer4_outputs(1168) <= b;
    layer4_outputs(1169) <= not (a or b);
    layer4_outputs(1170) <= not (a or b);
    layer4_outputs(1171) <= not (a or b);
    layer4_outputs(1172) <= not a or b;
    layer4_outputs(1173) <= 1'b0;
    layer4_outputs(1174) <= 1'b0;
    layer4_outputs(1175) <= not a or b;
    layer4_outputs(1176) <= 1'b1;
    layer4_outputs(1177) <= b;
    layer4_outputs(1178) <= a;
    layer4_outputs(1179) <= not b;
    layer4_outputs(1180) <= b;
    layer4_outputs(1181) <= not b or a;
    layer4_outputs(1182) <= a or b;
    layer4_outputs(1183) <= not b or a;
    layer4_outputs(1184) <= not (a and b);
    layer4_outputs(1185) <= a and not b;
    layer4_outputs(1186) <= not a;
    layer4_outputs(1187) <= not b or a;
    layer4_outputs(1188) <= a and not b;
    layer4_outputs(1189) <= not a;
    layer4_outputs(1190) <= a and not b;
    layer4_outputs(1191) <= not b;
    layer4_outputs(1192) <= a or b;
    layer4_outputs(1193) <= b and not a;
    layer4_outputs(1194) <= not (a or b);
    layer4_outputs(1195) <= not (a or b);
    layer4_outputs(1196) <= b and not a;
    layer4_outputs(1197) <= not a;
    layer4_outputs(1198) <= b;
    layer4_outputs(1199) <= a and b;
    layer4_outputs(1200) <= a;
    layer4_outputs(1201) <= b;
    layer4_outputs(1202) <= a or b;
    layer4_outputs(1203) <= not a or b;
    layer4_outputs(1204) <= not (a xor b);
    layer4_outputs(1205) <= 1'b0;
    layer4_outputs(1206) <= not a or b;
    layer4_outputs(1207) <= not b;
    layer4_outputs(1208) <= 1'b0;
    layer4_outputs(1209) <= not a;
    layer4_outputs(1210) <= a and b;
    layer4_outputs(1211) <= a and b;
    layer4_outputs(1212) <= not a or b;
    layer4_outputs(1213) <= not a or b;
    layer4_outputs(1214) <= not b or a;
    layer4_outputs(1215) <= not a or b;
    layer4_outputs(1216) <= not (a or b);
    layer4_outputs(1217) <= not (a and b);
    layer4_outputs(1218) <= a;
    layer4_outputs(1219) <= b and not a;
    layer4_outputs(1220) <= not (a and b);
    layer4_outputs(1221) <= b;
    layer4_outputs(1222) <= not (a or b);
    layer4_outputs(1223) <= b;
    layer4_outputs(1224) <= 1'b0;
    layer4_outputs(1225) <= not a;
    layer4_outputs(1226) <= a or b;
    layer4_outputs(1227) <= not (a and b);
    layer4_outputs(1228) <= a or b;
    layer4_outputs(1229) <= b;
    layer4_outputs(1230) <= a or b;
    layer4_outputs(1231) <= not a;
    layer4_outputs(1232) <= not b or a;
    layer4_outputs(1233) <= not (a or b);
    layer4_outputs(1234) <= a or b;
    layer4_outputs(1235) <= not b;
    layer4_outputs(1236) <= b and not a;
    layer4_outputs(1237) <= not b;
    layer4_outputs(1238) <= not a;
    layer4_outputs(1239) <= a or b;
    layer4_outputs(1240) <= 1'b0;
    layer4_outputs(1241) <= a;
    layer4_outputs(1242) <= a and b;
    layer4_outputs(1243) <= not b or a;
    layer4_outputs(1244) <= 1'b0;
    layer4_outputs(1245) <= a and not b;
    layer4_outputs(1246) <= not (a and b);
    layer4_outputs(1247) <= not a;
    layer4_outputs(1248) <= b and not a;
    layer4_outputs(1249) <= not b;
    layer4_outputs(1250) <= b and not a;
    layer4_outputs(1251) <= not a;
    layer4_outputs(1252) <= 1'b0;
    layer4_outputs(1253) <= a and not b;
    layer4_outputs(1254) <= not b or a;
    layer4_outputs(1255) <= a;
    layer4_outputs(1256) <= 1'b0;
    layer4_outputs(1257) <= a;
    layer4_outputs(1258) <= not b or a;
    layer4_outputs(1259) <= b;
    layer4_outputs(1260) <= b;
    layer4_outputs(1261) <= not (a and b);
    layer4_outputs(1262) <= not (a or b);
    layer4_outputs(1263) <= b;
    layer4_outputs(1264) <= not b or a;
    layer4_outputs(1265) <= not (a and b);
    layer4_outputs(1266) <= not (a and b);
    layer4_outputs(1267) <= not b;
    layer4_outputs(1268) <= not b;
    layer4_outputs(1269) <= a;
    layer4_outputs(1270) <= 1'b0;
    layer4_outputs(1271) <= a and not b;
    layer4_outputs(1272) <= not (a or b);
    layer4_outputs(1273) <= a and not b;
    layer4_outputs(1274) <= 1'b1;
    layer4_outputs(1275) <= not a or b;
    layer4_outputs(1276) <= a and not b;
    layer4_outputs(1277) <= not a;
    layer4_outputs(1278) <= not a or b;
    layer4_outputs(1279) <= not a or b;
    layer4_outputs(1280) <= 1'b1;
    layer4_outputs(1281) <= a or b;
    layer4_outputs(1282) <= not a or b;
    layer4_outputs(1283) <= not (a or b);
    layer4_outputs(1284) <= 1'b1;
    layer4_outputs(1285) <= a and b;
    layer4_outputs(1286) <= not b or a;
    layer4_outputs(1287) <= a and not b;
    layer4_outputs(1288) <= 1'b0;
    layer4_outputs(1289) <= b;
    layer4_outputs(1290) <= not (a or b);
    layer4_outputs(1291) <= a xor b;
    layer4_outputs(1292) <= a and not b;
    layer4_outputs(1293) <= 1'b1;
    layer4_outputs(1294) <= not (a or b);
    layer4_outputs(1295) <= b and not a;
    layer4_outputs(1296) <= b and not a;
    layer4_outputs(1297) <= a or b;
    layer4_outputs(1298) <= b and not a;
    layer4_outputs(1299) <= a and not b;
    layer4_outputs(1300) <= not a or b;
    layer4_outputs(1301) <= 1'b1;
    layer4_outputs(1302) <= not a;
    layer4_outputs(1303) <= not (a or b);
    layer4_outputs(1304) <= a;
    layer4_outputs(1305) <= b and not a;
    layer4_outputs(1306) <= 1'b0;
    layer4_outputs(1307) <= a or b;
    layer4_outputs(1308) <= not a or b;
    layer4_outputs(1309) <= not (a or b);
    layer4_outputs(1310) <= a;
    layer4_outputs(1311) <= not (a or b);
    layer4_outputs(1312) <= a or b;
    layer4_outputs(1313) <= a and b;
    layer4_outputs(1314) <= not a or b;
    layer4_outputs(1315) <= a;
    layer4_outputs(1316) <= not a or b;
    layer4_outputs(1317) <= b;
    layer4_outputs(1318) <= not (a or b);
    layer4_outputs(1319) <= not a or b;
    layer4_outputs(1320) <= not (a and b);
    layer4_outputs(1321) <= a and not b;
    layer4_outputs(1322) <= not b;
    layer4_outputs(1323) <= not b;
    layer4_outputs(1324) <= 1'b0;
    layer4_outputs(1325) <= a or b;
    layer4_outputs(1326) <= a;
    layer4_outputs(1327) <= a;
    layer4_outputs(1328) <= not a or b;
    layer4_outputs(1329) <= a and b;
    layer4_outputs(1330) <= not b or a;
    layer4_outputs(1331) <= 1'b0;
    layer4_outputs(1332) <= not b;
    layer4_outputs(1333) <= not (a and b);
    layer4_outputs(1334) <= not b;
    layer4_outputs(1335) <= 1'b0;
    layer4_outputs(1336) <= b and not a;
    layer4_outputs(1337) <= a and b;
    layer4_outputs(1338) <= a and b;
    layer4_outputs(1339) <= not (a and b);
    layer4_outputs(1340) <= 1'b1;
    layer4_outputs(1341) <= not b;
    layer4_outputs(1342) <= b and not a;
    layer4_outputs(1343) <= a or b;
    layer4_outputs(1344) <= not a or b;
    layer4_outputs(1345) <= a or b;
    layer4_outputs(1346) <= not (a and b);
    layer4_outputs(1347) <= not (a and b);
    layer4_outputs(1348) <= a and not b;
    layer4_outputs(1349) <= a;
    layer4_outputs(1350) <= not (a or b);
    layer4_outputs(1351) <= not (a or b);
    layer4_outputs(1352) <= not b;
    layer4_outputs(1353) <= 1'b1;
    layer4_outputs(1354) <= not (a or b);
    layer4_outputs(1355) <= 1'b0;
    layer4_outputs(1356) <= not b or a;
    layer4_outputs(1357) <= b;
    layer4_outputs(1358) <= a and b;
    layer4_outputs(1359) <= not a or b;
    layer4_outputs(1360) <= b and not a;
    layer4_outputs(1361) <= not (a or b);
    layer4_outputs(1362) <= b;
    layer4_outputs(1363) <= not (a xor b);
    layer4_outputs(1364) <= not a;
    layer4_outputs(1365) <= not a;
    layer4_outputs(1366) <= not (a and b);
    layer4_outputs(1367) <= a xor b;
    layer4_outputs(1368) <= a;
    layer4_outputs(1369) <= not a;
    layer4_outputs(1370) <= not a or b;
    layer4_outputs(1371) <= b;
    layer4_outputs(1372) <= not b;
    layer4_outputs(1373) <= 1'b0;
    layer4_outputs(1374) <= not a;
    layer4_outputs(1375) <= not b or a;
    layer4_outputs(1376) <= a and b;
    layer4_outputs(1377) <= b and not a;
    layer4_outputs(1378) <= not b;
    layer4_outputs(1379) <= a and b;
    layer4_outputs(1380) <= a and b;
    layer4_outputs(1381) <= not b or a;
    layer4_outputs(1382) <= not b;
    layer4_outputs(1383) <= not b or a;
    layer4_outputs(1384) <= not a or b;
    layer4_outputs(1385) <= not a;
    layer4_outputs(1386) <= b and not a;
    layer4_outputs(1387) <= 1'b0;
    layer4_outputs(1388) <= a;
    layer4_outputs(1389) <= 1'b0;
    layer4_outputs(1390) <= a and b;
    layer4_outputs(1391) <= not a or b;
    layer4_outputs(1392) <= not b or a;
    layer4_outputs(1393) <= b;
    layer4_outputs(1394) <= not a;
    layer4_outputs(1395) <= not (a and b);
    layer4_outputs(1396) <= b;
    layer4_outputs(1397) <= a;
    layer4_outputs(1398) <= b;
    layer4_outputs(1399) <= not b;
    layer4_outputs(1400) <= not b;
    layer4_outputs(1401) <= not (a and b);
    layer4_outputs(1402) <= a and b;
    layer4_outputs(1403) <= not (a and b);
    layer4_outputs(1404) <= not a;
    layer4_outputs(1405) <= not (a or b);
    layer4_outputs(1406) <= not a or b;
    layer4_outputs(1407) <= not a;
    layer4_outputs(1408) <= 1'b1;
    layer4_outputs(1409) <= not a;
    layer4_outputs(1410) <= 1'b0;
    layer4_outputs(1411) <= 1'b1;
    layer4_outputs(1412) <= a and not b;
    layer4_outputs(1413) <= a or b;
    layer4_outputs(1414) <= not (a and b);
    layer4_outputs(1415) <= a and b;
    layer4_outputs(1416) <= not a or b;
    layer4_outputs(1417) <= b;
    layer4_outputs(1418) <= not a;
    layer4_outputs(1419) <= b;
    layer4_outputs(1420) <= b;
    layer4_outputs(1421) <= a and b;
    layer4_outputs(1422) <= 1'b0;
    layer4_outputs(1423) <= a or b;
    layer4_outputs(1424) <= b and not a;
    layer4_outputs(1425) <= not a or b;
    layer4_outputs(1426) <= a or b;
    layer4_outputs(1427) <= a;
    layer4_outputs(1428) <= 1'b1;
    layer4_outputs(1429) <= 1'b0;
    layer4_outputs(1430) <= a;
    layer4_outputs(1431) <= 1'b0;
    layer4_outputs(1432) <= not b or a;
    layer4_outputs(1433) <= not (a and b);
    layer4_outputs(1434) <= not a or b;
    layer4_outputs(1435) <= b and not a;
    layer4_outputs(1436) <= not a;
    layer4_outputs(1437) <= a and b;
    layer4_outputs(1438) <= not b;
    layer4_outputs(1439) <= a and b;
    layer4_outputs(1440) <= not (a or b);
    layer4_outputs(1441) <= 1'b0;
    layer4_outputs(1442) <= a;
    layer4_outputs(1443) <= a;
    layer4_outputs(1444) <= not a;
    layer4_outputs(1445) <= 1'b0;
    layer4_outputs(1446) <= a;
    layer4_outputs(1447) <= not b;
    layer4_outputs(1448) <= not b or a;
    layer4_outputs(1449) <= a and b;
    layer4_outputs(1450) <= 1'b0;
    layer4_outputs(1451) <= 1'b0;
    layer4_outputs(1452) <= not b or a;
    layer4_outputs(1453) <= not (a and b);
    layer4_outputs(1454) <= not (a and b);
    layer4_outputs(1455) <= 1'b0;
    layer4_outputs(1456) <= a xor b;
    layer4_outputs(1457) <= 1'b0;
    layer4_outputs(1458) <= b;
    layer4_outputs(1459) <= a;
    layer4_outputs(1460) <= not a or b;
    layer4_outputs(1461) <= 1'b1;
    layer4_outputs(1462) <= 1'b1;
    layer4_outputs(1463) <= not (a or b);
    layer4_outputs(1464) <= b and not a;
    layer4_outputs(1465) <= not a;
    layer4_outputs(1466) <= b;
    layer4_outputs(1467) <= a and b;
    layer4_outputs(1468) <= a or b;
    layer4_outputs(1469) <= not b or a;
    layer4_outputs(1470) <= a or b;
    layer4_outputs(1471) <= b and not a;
    layer4_outputs(1472) <= a;
    layer4_outputs(1473) <= not (a or b);
    layer4_outputs(1474) <= a;
    layer4_outputs(1475) <= b;
    layer4_outputs(1476) <= a and not b;
    layer4_outputs(1477) <= 1'b1;
    layer4_outputs(1478) <= 1'b1;
    layer4_outputs(1479) <= a xor b;
    layer4_outputs(1480) <= b and not a;
    layer4_outputs(1481) <= a;
    layer4_outputs(1482) <= 1'b1;
    layer4_outputs(1483) <= 1'b1;
    layer4_outputs(1484) <= 1'b0;
    layer4_outputs(1485) <= not b or a;
    layer4_outputs(1486) <= not (a or b);
    layer4_outputs(1487) <= not (a and b);
    layer4_outputs(1488) <= not b or a;
    layer4_outputs(1489) <= 1'b0;
    layer4_outputs(1490) <= not b;
    layer4_outputs(1491) <= b;
    layer4_outputs(1492) <= b;
    layer4_outputs(1493) <= a and b;
    layer4_outputs(1494) <= a or b;
    layer4_outputs(1495) <= 1'b1;
    layer4_outputs(1496) <= a and b;
    layer4_outputs(1497) <= not b or a;
    layer4_outputs(1498) <= 1'b1;
    layer4_outputs(1499) <= b and not a;
    layer4_outputs(1500) <= not (a and b);
    layer4_outputs(1501) <= a;
    layer4_outputs(1502) <= 1'b0;
    layer4_outputs(1503) <= a xor b;
    layer4_outputs(1504) <= not (a or b);
    layer4_outputs(1505) <= a and b;
    layer4_outputs(1506) <= 1'b0;
    layer4_outputs(1507) <= not (a and b);
    layer4_outputs(1508) <= a or b;
    layer4_outputs(1509) <= not b;
    layer4_outputs(1510) <= 1'b0;
    layer4_outputs(1511) <= a and b;
    layer4_outputs(1512) <= not b;
    layer4_outputs(1513) <= not a;
    layer4_outputs(1514) <= 1'b0;
    layer4_outputs(1515) <= a;
    layer4_outputs(1516) <= b and not a;
    layer4_outputs(1517) <= 1'b0;
    layer4_outputs(1518) <= not a;
    layer4_outputs(1519) <= not b;
    layer4_outputs(1520) <= not b;
    layer4_outputs(1521) <= 1'b0;
    layer4_outputs(1522) <= not a;
    layer4_outputs(1523) <= 1'b0;
    layer4_outputs(1524) <= not a or b;
    layer4_outputs(1525) <= a;
    layer4_outputs(1526) <= a and not b;
    layer4_outputs(1527) <= not a or b;
    layer4_outputs(1528) <= not a or b;
    layer4_outputs(1529) <= not (a and b);
    layer4_outputs(1530) <= b;
    layer4_outputs(1531) <= b and not a;
    layer4_outputs(1532) <= a xor b;
    layer4_outputs(1533) <= not b;
    layer4_outputs(1534) <= a;
    layer4_outputs(1535) <= b and not a;
    layer4_outputs(1536) <= a and not b;
    layer4_outputs(1537) <= 1'b0;
    layer4_outputs(1538) <= a and not b;
    layer4_outputs(1539) <= not (a xor b);
    layer4_outputs(1540) <= not a;
    layer4_outputs(1541) <= not a;
    layer4_outputs(1542) <= 1'b0;
    layer4_outputs(1543) <= not b or a;
    layer4_outputs(1544) <= a and not b;
    layer4_outputs(1545) <= not b or a;
    layer4_outputs(1546) <= not a;
    layer4_outputs(1547) <= not b;
    layer4_outputs(1548) <= 1'b0;
    layer4_outputs(1549) <= a and b;
    layer4_outputs(1550) <= a and not b;
    layer4_outputs(1551) <= not b;
    layer4_outputs(1552) <= a;
    layer4_outputs(1553) <= not a or b;
    layer4_outputs(1554) <= b;
    layer4_outputs(1555) <= b;
    layer4_outputs(1556) <= not a or b;
    layer4_outputs(1557) <= 1'b0;
    layer4_outputs(1558) <= not a or b;
    layer4_outputs(1559) <= a or b;
    layer4_outputs(1560) <= a and not b;
    layer4_outputs(1561) <= not (a and b);
    layer4_outputs(1562) <= not b;
    layer4_outputs(1563) <= b;
    layer4_outputs(1564) <= a and not b;
    layer4_outputs(1565) <= b;
    layer4_outputs(1566) <= not (a or b);
    layer4_outputs(1567) <= 1'b1;
    layer4_outputs(1568) <= a and not b;
    layer4_outputs(1569) <= not b;
    layer4_outputs(1570) <= 1'b1;
    layer4_outputs(1571) <= not a or b;
    layer4_outputs(1572) <= a or b;
    layer4_outputs(1573) <= a and b;
    layer4_outputs(1574) <= b and not a;
    layer4_outputs(1575) <= 1'b0;
    layer4_outputs(1576) <= not a or b;
    layer4_outputs(1577) <= 1'b0;
    layer4_outputs(1578) <= not b or a;
    layer4_outputs(1579) <= not a;
    layer4_outputs(1580) <= not (a xor b);
    layer4_outputs(1581) <= not b or a;
    layer4_outputs(1582) <= not (a and b);
    layer4_outputs(1583) <= a;
    layer4_outputs(1584) <= b;
    layer4_outputs(1585) <= not (a and b);
    layer4_outputs(1586) <= not (a or b);
    layer4_outputs(1587) <= 1'b0;
    layer4_outputs(1588) <= not (a or b);
    layer4_outputs(1589) <= a;
    layer4_outputs(1590) <= a or b;
    layer4_outputs(1591) <= 1'b0;
    layer4_outputs(1592) <= b;
    layer4_outputs(1593) <= 1'b0;
    layer4_outputs(1594) <= not b or a;
    layer4_outputs(1595) <= not b;
    layer4_outputs(1596) <= not a;
    layer4_outputs(1597) <= not (a or b);
    layer4_outputs(1598) <= 1'b1;
    layer4_outputs(1599) <= not (a or b);
    layer4_outputs(1600) <= a or b;
    layer4_outputs(1601) <= b and not a;
    layer4_outputs(1602) <= b;
    layer4_outputs(1603) <= a or b;
    layer4_outputs(1604) <= not b or a;
    layer4_outputs(1605) <= not a or b;
    layer4_outputs(1606) <= 1'b0;
    layer4_outputs(1607) <= not a or b;
    layer4_outputs(1608) <= not a or b;
    layer4_outputs(1609) <= not (a or b);
    layer4_outputs(1610) <= not (a or b);
    layer4_outputs(1611) <= b and not a;
    layer4_outputs(1612) <= b;
    layer4_outputs(1613) <= a xor b;
    layer4_outputs(1614) <= a xor b;
    layer4_outputs(1615) <= b and not a;
    layer4_outputs(1616) <= not (a and b);
    layer4_outputs(1617) <= a and b;
    layer4_outputs(1618) <= not (a and b);
    layer4_outputs(1619) <= not (a or b);
    layer4_outputs(1620) <= 1'b0;
    layer4_outputs(1621) <= b;
    layer4_outputs(1622) <= 1'b1;
    layer4_outputs(1623) <= a and b;
    layer4_outputs(1624) <= not (a or b);
    layer4_outputs(1625) <= not b or a;
    layer4_outputs(1626) <= not (a or b);
    layer4_outputs(1627) <= a or b;
    layer4_outputs(1628) <= a or b;
    layer4_outputs(1629) <= not a;
    layer4_outputs(1630) <= a;
    layer4_outputs(1631) <= a or b;
    layer4_outputs(1632) <= a and b;
    layer4_outputs(1633) <= 1'b1;
    layer4_outputs(1634) <= not (a and b);
    layer4_outputs(1635) <= not (a and b);
    layer4_outputs(1636) <= not a or b;
    layer4_outputs(1637) <= not b or a;
    layer4_outputs(1638) <= a and not b;
    layer4_outputs(1639) <= b and not a;
    layer4_outputs(1640) <= 1'b0;
    layer4_outputs(1641) <= not (a xor b);
    layer4_outputs(1642) <= 1'b0;
    layer4_outputs(1643) <= b and not a;
    layer4_outputs(1644) <= not b or a;
    layer4_outputs(1645) <= 1'b1;
    layer4_outputs(1646) <= a;
    layer4_outputs(1647) <= not a;
    layer4_outputs(1648) <= a and not b;
    layer4_outputs(1649) <= b and not a;
    layer4_outputs(1650) <= not (a or b);
    layer4_outputs(1651) <= not (a and b);
    layer4_outputs(1652) <= not b or a;
    layer4_outputs(1653) <= not b or a;
    layer4_outputs(1654) <= a;
    layer4_outputs(1655) <= not a;
    layer4_outputs(1656) <= a;
    layer4_outputs(1657) <= not a or b;
    layer4_outputs(1658) <= a or b;
    layer4_outputs(1659) <= not (a and b);
    layer4_outputs(1660) <= not a;
    layer4_outputs(1661) <= a;
    layer4_outputs(1662) <= a or b;
    layer4_outputs(1663) <= b and not a;
    layer4_outputs(1664) <= a;
    layer4_outputs(1665) <= not b;
    layer4_outputs(1666) <= a and not b;
    layer4_outputs(1667) <= not (a and b);
    layer4_outputs(1668) <= a and b;
    layer4_outputs(1669) <= a;
    layer4_outputs(1670) <= not (a xor b);
    layer4_outputs(1671) <= not (a or b);
    layer4_outputs(1672) <= not b or a;
    layer4_outputs(1673) <= b;
    layer4_outputs(1674) <= a or b;
    layer4_outputs(1675) <= a and b;
    layer4_outputs(1676) <= b;
    layer4_outputs(1677) <= b;
    layer4_outputs(1678) <= not (a and b);
    layer4_outputs(1679) <= a or b;
    layer4_outputs(1680) <= not (a or b);
    layer4_outputs(1681) <= not (a or b);
    layer4_outputs(1682) <= not b;
    layer4_outputs(1683) <= 1'b0;
    layer4_outputs(1684) <= not (a and b);
    layer4_outputs(1685) <= 1'b0;
    layer4_outputs(1686) <= not a;
    layer4_outputs(1687) <= not b or a;
    layer4_outputs(1688) <= 1'b0;
    layer4_outputs(1689) <= a;
    layer4_outputs(1690) <= a;
    layer4_outputs(1691) <= not (a and b);
    layer4_outputs(1692) <= not b;
    layer4_outputs(1693) <= b and not a;
    layer4_outputs(1694) <= not b;
    layer4_outputs(1695) <= not a;
    layer4_outputs(1696) <= not a or b;
    layer4_outputs(1697) <= not a or b;
    layer4_outputs(1698) <= not b or a;
    layer4_outputs(1699) <= 1'b1;
    layer4_outputs(1700) <= not b;
    layer4_outputs(1701) <= a and not b;
    layer4_outputs(1702) <= a and b;
    layer4_outputs(1703) <= a and b;
    layer4_outputs(1704) <= not (a and b);
    layer4_outputs(1705) <= a or b;
    layer4_outputs(1706) <= not (a and b);
    layer4_outputs(1707) <= 1'b1;
    layer4_outputs(1708) <= a and b;
    layer4_outputs(1709) <= not a or b;
    layer4_outputs(1710) <= not b;
    layer4_outputs(1711) <= not a or b;
    layer4_outputs(1712) <= b;
    layer4_outputs(1713) <= a;
    layer4_outputs(1714) <= not (a and b);
    layer4_outputs(1715) <= 1'b1;
    layer4_outputs(1716) <= a or b;
    layer4_outputs(1717) <= 1'b0;
    layer4_outputs(1718) <= a and not b;
    layer4_outputs(1719) <= 1'b1;
    layer4_outputs(1720) <= not a;
    layer4_outputs(1721) <= not (a and b);
    layer4_outputs(1722) <= a or b;
    layer4_outputs(1723) <= b and not a;
    layer4_outputs(1724) <= not (a or b);
    layer4_outputs(1725) <= not a or b;
    layer4_outputs(1726) <= a and b;
    layer4_outputs(1727) <= a and b;
    layer4_outputs(1728) <= not a;
    layer4_outputs(1729) <= b;
    layer4_outputs(1730) <= not b or a;
    layer4_outputs(1731) <= not a;
    layer4_outputs(1732) <= 1'b1;
    layer4_outputs(1733) <= b;
    layer4_outputs(1734) <= a and not b;
    layer4_outputs(1735) <= a;
    layer4_outputs(1736) <= a and b;
    layer4_outputs(1737) <= not a;
    layer4_outputs(1738) <= a and not b;
    layer4_outputs(1739) <= not (a or b);
    layer4_outputs(1740) <= not (a xor b);
    layer4_outputs(1741) <= b;
    layer4_outputs(1742) <= 1'b0;
    layer4_outputs(1743) <= not b or a;
    layer4_outputs(1744) <= 1'b1;
    layer4_outputs(1745) <= 1'b0;
    layer4_outputs(1746) <= a or b;
    layer4_outputs(1747) <= a;
    layer4_outputs(1748) <= not (a xor b);
    layer4_outputs(1749) <= not (a and b);
    layer4_outputs(1750) <= not b or a;
    layer4_outputs(1751) <= 1'b1;
    layer4_outputs(1752) <= 1'b0;
    layer4_outputs(1753) <= not (a or b);
    layer4_outputs(1754) <= not (a and b);
    layer4_outputs(1755) <= not (a or b);
    layer4_outputs(1756) <= a and b;
    layer4_outputs(1757) <= not a or b;
    layer4_outputs(1758) <= not b;
    layer4_outputs(1759) <= a or b;
    layer4_outputs(1760) <= a;
    layer4_outputs(1761) <= b;
    layer4_outputs(1762) <= not a;
    layer4_outputs(1763) <= 1'b0;
    layer4_outputs(1764) <= 1'b0;
    layer4_outputs(1765) <= not b or a;
    layer4_outputs(1766) <= a or b;
    layer4_outputs(1767) <= not a or b;
    layer4_outputs(1768) <= not b or a;
    layer4_outputs(1769) <= not b;
    layer4_outputs(1770) <= not (a and b);
    layer4_outputs(1771) <= not (a and b);
    layer4_outputs(1772) <= b;
    layer4_outputs(1773) <= a or b;
    layer4_outputs(1774) <= not (a and b);
    layer4_outputs(1775) <= a;
    layer4_outputs(1776) <= a xor b;
    layer4_outputs(1777) <= b;
    layer4_outputs(1778) <= a and b;
    layer4_outputs(1779) <= a and not b;
    layer4_outputs(1780) <= a xor b;
    layer4_outputs(1781) <= a and not b;
    layer4_outputs(1782) <= a and b;
    layer4_outputs(1783) <= b and not a;
    layer4_outputs(1784) <= a and not b;
    layer4_outputs(1785) <= 1'b0;
    layer4_outputs(1786) <= a and not b;
    layer4_outputs(1787) <= not b or a;
    layer4_outputs(1788) <= a;
    layer4_outputs(1789) <= 1'b1;
    layer4_outputs(1790) <= not a or b;
    layer4_outputs(1791) <= b and not a;
    layer4_outputs(1792) <= a and not b;
    layer4_outputs(1793) <= 1'b0;
    layer4_outputs(1794) <= not a or b;
    layer4_outputs(1795) <= 1'b0;
    layer4_outputs(1796) <= not b;
    layer4_outputs(1797) <= 1'b0;
    layer4_outputs(1798) <= a;
    layer4_outputs(1799) <= not b or a;
    layer4_outputs(1800) <= not b;
    layer4_outputs(1801) <= not b;
    layer4_outputs(1802) <= a and b;
    layer4_outputs(1803) <= not (a xor b);
    layer4_outputs(1804) <= not (a or b);
    layer4_outputs(1805) <= 1'b0;
    layer4_outputs(1806) <= a and not b;
    layer4_outputs(1807) <= not a or b;
    layer4_outputs(1808) <= 1'b0;
    layer4_outputs(1809) <= 1'b1;
    layer4_outputs(1810) <= not (a and b);
    layer4_outputs(1811) <= not (a or b);
    layer4_outputs(1812) <= a and not b;
    layer4_outputs(1813) <= not (a or b);
    layer4_outputs(1814) <= not (a or b);
    layer4_outputs(1815) <= not (a and b);
    layer4_outputs(1816) <= not b;
    layer4_outputs(1817) <= a and not b;
    layer4_outputs(1818) <= a or b;
    layer4_outputs(1819) <= a and not b;
    layer4_outputs(1820) <= not (a and b);
    layer4_outputs(1821) <= not b;
    layer4_outputs(1822) <= not (a and b);
    layer4_outputs(1823) <= a;
    layer4_outputs(1824) <= not b or a;
    layer4_outputs(1825) <= not (a or b);
    layer4_outputs(1826) <= 1'b1;
    layer4_outputs(1827) <= 1'b0;
    layer4_outputs(1828) <= b and not a;
    layer4_outputs(1829) <= b and not a;
    layer4_outputs(1830) <= not (a or b);
    layer4_outputs(1831) <= a;
    layer4_outputs(1832) <= a or b;
    layer4_outputs(1833) <= b and not a;
    layer4_outputs(1834) <= not (a or b);
    layer4_outputs(1835) <= not b;
    layer4_outputs(1836) <= not b;
    layer4_outputs(1837) <= b and not a;
    layer4_outputs(1838) <= a or b;
    layer4_outputs(1839) <= not a or b;
    layer4_outputs(1840) <= a and b;
    layer4_outputs(1841) <= 1'b1;
    layer4_outputs(1842) <= not (a and b);
    layer4_outputs(1843) <= b;
    layer4_outputs(1844) <= a or b;
    layer4_outputs(1845) <= not b or a;
    layer4_outputs(1846) <= a or b;
    layer4_outputs(1847) <= a or b;
    layer4_outputs(1848) <= a or b;
    layer4_outputs(1849) <= not (a and b);
    layer4_outputs(1850) <= not b;
    layer4_outputs(1851) <= a and not b;
    layer4_outputs(1852) <= b and not a;
    layer4_outputs(1853) <= not b or a;
    layer4_outputs(1854) <= a and not b;
    layer4_outputs(1855) <= b;
    layer4_outputs(1856) <= a and b;
    layer4_outputs(1857) <= not (a and b);
    layer4_outputs(1858) <= 1'b1;
    layer4_outputs(1859) <= a or b;
    layer4_outputs(1860) <= b;
    layer4_outputs(1861) <= not b or a;
    layer4_outputs(1862) <= 1'b0;
    layer4_outputs(1863) <= not (a and b);
    layer4_outputs(1864) <= not a;
    layer4_outputs(1865) <= b;
    layer4_outputs(1866) <= not b;
    layer4_outputs(1867) <= not a;
    layer4_outputs(1868) <= a;
    layer4_outputs(1869) <= b and not a;
    layer4_outputs(1870) <= not a or b;
    layer4_outputs(1871) <= a and b;
    layer4_outputs(1872) <= not b;
    layer4_outputs(1873) <= not b or a;
    layer4_outputs(1874) <= 1'b0;
    layer4_outputs(1875) <= a or b;
    layer4_outputs(1876) <= not a;
    layer4_outputs(1877) <= not b;
    layer4_outputs(1878) <= not (a or b);
    layer4_outputs(1879) <= a and b;
    layer4_outputs(1880) <= not (a or b);
    layer4_outputs(1881) <= a and b;
    layer4_outputs(1882) <= a or b;
    layer4_outputs(1883) <= not (a or b);
    layer4_outputs(1884) <= a;
    layer4_outputs(1885) <= a;
    layer4_outputs(1886) <= not (a and b);
    layer4_outputs(1887) <= not a or b;
    layer4_outputs(1888) <= not b;
    layer4_outputs(1889) <= not b or a;
    layer4_outputs(1890) <= 1'b1;
    layer4_outputs(1891) <= b;
    layer4_outputs(1892) <= b;
    layer4_outputs(1893) <= a;
    layer4_outputs(1894) <= a or b;
    layer4_outputs(1895) <= not (a and b);
    layer4_outputs(1896) <= a and b;
    layer4_outputs(1897) <= not (a and b);
    layer4_outputs(1898) <= a and not b;
    layer4_outputs(1899) <= a and b;
    layer4_outputs(1900) <= a and not b;
    layer4_outputs(1901) <= not (a and b);
    layer4_outputs(1902) <= b and not a;
    layer4_outputs(1903) <= b;
    layer4_outputs(1904) <= b;
    layer4_outputs(1905) <= not b or a;
    layer4_outputs(1906) <= 1'b1;
    layer4_outputs(1907) <= a and not b;
    layer4_outputs(1908) <= not b or a;
    layer4_outputs(1909) <= 1'b1;
    layer4_outputs(1910) <= 1'b1;
    layer4_outputs(1911) <= not a;
    layer4_outputs(1912) <= a;
    layer4_outputs(1913) <= not b;
    layer4_outputs(1914) <= not b;
    layer4_outputs(1915) <= not b;
    layer4_outputs(1916) <= not b or a;
    layer4_outputs(1917) <= not (a and b);
    layer4_outputs(1918) <= not (a and b);
    layer4_outputs(1919) <= not (a or b);
    layer4_outputs(1920) <= a and not b;
    layer4_outputs(1921) <= not (a xor b);
    layer4_outputs(1922) <= not (a or b);
    layer4_outputs(1923) <= not (a or b);
    layer4_outputs(1924) <= not a;
    layer4_outputs(1925) <= not a;
    layer4_outputs(1926) <= not (a or b);
    layer4_outputs(1927) <= a and not b;
    layer4_outputs(1928) <= a xor b;
    layer4_outputs(1929) <= b and not a;
    layer4_outputs(1930) <= not a or b;
    layer4_outputs(1931) <= a and not b;
    layer4_outputs(1932) <= b and not a;
    layer4_outputs(1933) <= not (a xor b);
    layer4_outputs(1934) <= not a;
    layer4_outputs(1935) <= not a;
    layer4_outputs(1936) <= not b or a;
    layer4_outputs(1937) <= not a or b;
    layer4_outputs(1938) <= a and b;
    layer4_outputs(1939) <= 1'b0;
    layer4_outputs(1940) <= b and not a;
    layer4_outputs(1941) <= b;
    layer4_outputs(1942) <= not (a and b);
    layer4_outputs(1943) <= a and b;
    layer4_outputs(1944) <= a or b;
    layer4_outputs(1945) <= not b;
    layer4_outputs(1946) <= not b;
    layer4_outputs(1947) <= not b;
    layer4_outputs(1948) <= not (a and b);
    layer4_outputs(1949) <= not a or b;
    layer4_outputs(1950) <= a;
    layer4_outputs(1951) <= a or b;
    layer4_outputs(1952) <= 1'b0;
    layer4_outputs(1953) <= not (a and b);
    layer4_outputs(1954) <= b and not a;
    layer4_outputs(1955) <= 1'b0;
    layer4_outputs(1956) <= not a;
    layer4_outputs(1957) <= 1'b0;
    layer4_outputs(1958) <= not (a or b);
    layer4_outputs(1959) <= a or b;
    layer4_outputs(1960) <= not b;
    layer4_outputs(1961) <= 1'b1;
    layer4_outputs(1962) <= a;
    layer4_outputs(1963) <= a and not b;
    layer4_outputs(1964) <= 1'b1;
    layer4_outputs(1965) <= 1'b1;
    layer4_outputs(1966) <= a;
    layer4_outputs(1967) <= not (a or b);
    layer4_outputs(1968) <= a xor b;
    layer4_outputs(1969) <= b and not a;
    layer4_outputs(1970) <= not a or b;
    layer4_outputs(1971) <= 1'b0;
    layer4_outputs(1972) <= not (a and b);
    layer4_outputs(1973) <= a;
    layer4_outputs(1974) <= a;
    layer4_outputs(1975) <= a and b;
    layer4_outputs(1976) <= 1'b1;
    layer4_outputs(1977) <= b and not a;
    layer4_outputs(1978) <= b and not a;
    layer4_outputs(1979) <= b and not a;
    layer4_outputs(1980) <= b;
    layer4_outputs(1981) <= b;
    layer4_outputs(1982) <= a or b;
    layer4_outputs(1983) <= not b or a;
    layer4_outputs(1984) <= a xor b;
    layer4_outputs(1985) <= 1'b0;
    layer4_outputs(1986) <= b and not a;
    layer4_outputs(1987) <= not (a and b);
    layer4_outputs(1988) <= a and not b;
    layer4_outputs(1989) <= not a or b;
    layer4_outputs(1990) <= a and b;
    layer4_outputs(1991) <= not a;
    layer4_outputs(1992) <= not (a or b);
    layer4_outputs(1993) <= a xor b;
    layer4_outputs(1994) <= 1'b1;
    layer4_outputs(1995) <= b;
    layer4_outputs(1996) <= not a;
    layer4_outputs(1997) <= not a or b;
    layer4_outputs(1998) <= b;
    layer4_outputs(1999) <= not b or a;
    layer4_outputs(2000) <= 1'b0;
    layer4_outputs(2001) <= b;
    layer4_outputs(2002) <= not b or a;
    layer4_outputs(2003) <= 1'b1;
    layer4_outputs(2004) <= not b or a;
    layer4_outputs(2005) <= not (a xor b);
    layer4_outputs(2006) <= not b;
    layer4_outputs(2007) <= not a;
    layer4_outputs(2008) <= a and not b;
    layer4_outputs(2009) <= 1'b0;
    layer4_outputs(2010) <= a;
    layer4_outputs(2011) <= a or b;
    layer4_outputs(2012) <= b;
    layer4_outputs(2013) <= a and not b;
    layer4_outputs(2014) <= not a or b;
    layer4_outputs(2015) <= not (a or b);
    layer4_outputs(2016) <= not (a and b);
    layer4_outputs(2017) <= a xor b;
    layer4_outputs(2018) <= not (a or b);
    layer4_outputs(2019) <= not b or a;
    layer4_outputs(2020) <= 1'b1;
    layer4_outputs(2021) <= a and not b;
    layer4_outputs(2022) <= not a;
    layer4_outputs(2023) <= not a or b;
    layer4_outputs(2024) <= a;
    layer4_outputs(2025) <= not (a and b);
    layer4_outputs(2026) <= not (a xor b);
    layer4_outputs(2027) <= a;
    layer4_outputs(2028) <= b;
    layer4_outputs(2029) <= not (a and b);
    layer4_outputs(2030) <= not b or a;
    layer4_outputs(2031) <= not a;
    layer4_outputs(2032) <= a and b;
    layer4_outputs(2033) <= not b or a;
    layer4_outputs(2034) <= a or b;
    layer4_outputs(2035) <= b and not a;
    layer4_outputs(2036) <= not a;
    layer4_outputs(2037) <= not a;
    layer4_outputs(2038) <= a and not b;
    layer4_outputs(2039) <= not (a and b);
    layer4_outputs(2040) <= a and not b;
    layer4_outputs(2041) <= b and not a;
    layer4_outputs(2042) <= not b or a;
    layer4_outputs(2043) <= a or b;
    layer4_outputs(2044) <= b and not a;
    layer4_outputs(2045) <= not a or b;
    layer4_outputs(2046) <= a xor b;
    layer4_outputs(2047) <= 1'b1;
    layer4_outputs(2048) <= not (a and b);
    layer4_outputs(2049) <= not (a or b);
    layer4_outputs(2050) <= not (a and b);
    layer4_outputs(2051) <= a and not b;
    layer4_outputs(2052) <= not (a and b);
    layer4_outputs(2053) <= not b;
    layer4_outputs(2054) <= not b or a;
    layer4_outputs(2055) <= 1'b1;
    layer4_outputs(2056) <= 1'b1;
    layer4_outputs(2057) <= b;
    layer4_outputs(2058) <= not b or a;
    layer4_outputs(2059) <= a or b;
    layer4_outputs(2060) <= not (a and b);
    layer4_outputs(2061) <= a or b;
    layer4_outputs(2062) <= not a or b;
    layer4_outputs(2063) <= 1'b0;
    layer4_outputs(2064) <= 1'b1;
    layer4_outputs(2065) <= a and b;
    layer4_outputs(2066) <= not a or b;
    layer4_outputs(2067) <= b;
    layer4_outputs(2068) <= a xor b;
    layer4_outputs(2069) <= not (a or b);
    layer4_outputs(2070) <= a and b;
    layer4_outputs(2071) <= a;
    layer4_outputs(2072) <= not a;
    layer4_outputs(2073) <= not a or b;
    layer4_outputs(2074) <= not b;
    layer4_outputs(2075) <= not b;
    layer4_outputs(2076) <= 1'b1;
    layer4_outputs(2077) <= 1'b1;
    layer4_outputs(2078) <= a;
    layer4_outputs(2079) <= 1'b1;
    layer4_outputs(2080) <= a or b;
    layer4_outputs(2081) <= a and b;
    layer4_outputs(2082) <= a xor b;
    layer4_outputs(2083) <= a;
    layer4_outputs(2084) <= not (a and b);
    layer4_outputs(2085) <= a or b;
    layer4_outputs(2086) <= 1'b0;
    layer4_outputs(2087) <= a or b;
    layer4_outputs(2088) <= 1'b0;
    layer4_outputs(2089) <= a and b;
    layer4_outputs(2090) <= 1'b1;
    layer4_outputs(2091) <= not a;
    layer4_outputs(2092) <= not (a and b);
    layer4_outputs(2093) <= a;
    layer4_outputs(2094) <= not (a and b);
    layer4_outputs(2095) <= 1'b1;
    layer4_outputs(2096) <= 1'b0;
    layer4_outputs(2097) <= b and not a;
    layer4_outputs(2098) <= not b;
    layer4_outputs(2099) <= not a or b;
    layer4_outputs(2100) <= not (a and b);
    layer4_outputs(2101) <= b and not a;
    layer4_outputs(2102) <= 1'b0;
    layer4_outputs(2103) <= not (a or b);
    layer4_outputs(2104) <= a and not b;
    layer4_outputs(2105) <= not a;
    layer4_outputs(2106) <= not (a or b);
    layer4_outputs(2107) <= not b or a;
    layer4_outputs(2108) <= not (a xor b);
    layer4_outputs(2109) <= not a;
    layer4_outputs(2110) <= 1'b1;
    layer4_outputs(2111) <= not b or a;
    layer4_outputs(2112) <= not a or b;
    layer4_outputs(2113) <= 1'b0;
    layer4_outputs(2114) <= not b or a;
    layer4_outputs(2115) <= not a or b;
    layer4_outputs(2116) <= 1'b0;
    layer4_outputs(2117) <= a or b;
    layer4_outputs(2118) <= a and b;
    layer4_outputs(2119) <= not b or a;
    layer4_outputs(2120) <= not (a or b);
    layer4_outputs(2121) <= not b;
    layer4_outputs(2122) <= not (a and b);
    layer4_outputs(2123) <= a or b;
    layer4_outputs(2124) <= 1'b0;
    layer4_outputs(2125) <= a and b;
    layer4_outputs(2126) <= not a;
    layer4_outputs(2127) <= a and b;
    layer4_outputs(2128) <= a and b;
    layer4_outputs(2129) <= b and not a;
    layer4_outputs(2130) <= a or b;
    layer4_outputs(2131) <= not (a xor b);
    layer4_outputs(2132) <= not a or b;
    layer4_outputs(2133) <= not b;
    layer4_outputs(2134) <= not (a or b);
    layer4_outputs(2135) <= 1'b0;
    layer4_outputs(2136) <= not (a or b);
    layer4_outputs(2137) <= not (a and b);
    layer4_outputs(2138) <= a and b;
    layer4_outputs(2139) <= a;
    layer4_outputs(2140) <= not b;
    layer4_outputs(2141) <= not b or a;
    layer4_outputs(2142) <= a and b;
    layer4_outputs(2143) <= not b or a;
    layer4_outputs(2144) <= 1'b1;
    layer4_outputs(2145) <= b and not a;
    layer4_outputs(2146) <= a;
    layer4_outputs(2147) <= not b or a;
    layer4_outputs(2148) <= a and b;
    layer4_outputs(2149) <= not (a and b);
    layer4_outputs(2150) <= not a;
    layer4_outputs(2151) <= a and not b;
    layer4_outputs(2152) <= a xor b;
    layer4_outputs(2153) <= not a or b;
    layer4_outputs(2154) <= not (a or b);
    layer4_outputs(2155) <= a;
    layer4_outputs(2156) <= a and not b;
    layer4_outputs(2157) <= not b;
    layer4_outputs(2158) <= not b;
    layer4_outputs(2159) <= a and b;
    layer4_outputs(2160) <= not b;
    layer4_outputs(2161) <= a and not b;
    layer4_outputs(2162) <= a or b;
    layer4_outputs(2163) <= a and b;
    layer4_outputs(2164) <= b;
    layer4_outputs(2165) <= a;
    layer4_outputs(2166) <= 1'b0;
    layer4_outputs(2167) <= a and not b;
    layer4_outputs(2168) <= a or b;
    layer4_outputs(2169) <= 1'b1;
    layer4_outputs(2170) <= a and b;
    layer4_outputs(2171) <= a or b;
    layer4_outputs(2172) <= b;
    layer4_outputs(2173) <= b and not a;
    layer4_outputs(2174) <= not a;
    layer4_outputs(2175) <= not b;
    layer4_outputs(2176) <= not b;
    layer4_outputs(2177) <= a;
    layer4_outputs(2178) <= not a;
    layer4_outputs(2179) <= a or b;
    layer4_outputs(2180) <= a and b;
    layer4_outputs(2181) <= not (a or b);
    layer4_outputs(2182) <= not b;
    layer4_outputs(2183) <= not a;
    layer4_outputs(2184) <= a or b;
    layer4_outputs(2185) <= a and not b;
    layer4_outputs(2186) <= a and not b;
    layer4_outputs(2187) <= 1'b0;
    layer4_outputs(2188) <= not b;
    layer4_outputs(2189) <= a;
    layer4_outputs(2190) <= b and not a;
    layer4_outputs(2191) <= a or b;
    layer4_outputs(2192) <= 1'b1;
    layer4_outputs(2193) <= a;
    layer4_outputs(2194) <= 1'b0;
    layer4_outputs(2195) <= 1'b0;
    layer4_outputs(2196) <= not (a or b);
    layer4_outputs(2197) <= b;
    layer4_outputs(2198) <= not (a or b);
    layer4_outputs(2199) <= b;
    layer4_outputs(2200) <= a;
    layer4_outputs(2201) <= not b;
    layer4_outputs(2202) <= not b;
    layer4_outputs(2203) <= not a;
    layer4_outputs(2204) <= b;
    layer4_outputs(2205) <= not a;
    layer4_outputs(2206) <= not b;
    layer4_outputs(2207) <= not a;
    layer4_outputs(2208) <= a and not b;
    layer4_outputs(2209) <= 1'b1;
    layer4_outputs(2210) <= b and not a;
    layer4_outputs(2211) <= a and b;
    layer4_outputs(2212) <= not a;
    layer4_outputs(2213) <= b;
    layer4_outputs(2214) <= b;
    layer4_outputs(2215) <= a;
    layer4_outputs(2216) <= not a or b;
    layer4_outputs(2217) <= a and b;
    layer4_outputs(2218) <= not a;
    layer4_outputs(2219) <= a or b;
    layer4_outputs(2220) <= not (a or b);
    layer4_outputs(2221) <= not (a or b);
    layer4_outputs(2222) <= not (a and b);
    layer4_outputs(2223) <= not a;
    layer4_outputs(2224) <= not (a and b);
    layer4_outputs(2225) <= not b;
    layer4_outputs(2226) <= not a;
    layer4_outputs(2227) <= a and b;
    layer4_outputs(2228) <= a;
    layer4_outputs(2229) <= not a or b;
    layer4_outputs(2230) <= a and not b;
    layer4_outputs(2231) <= b;
    layer4_outputs(2232) <= b;
    layer4_outputs(2233) <= not a;
    layer4_outputs(2234) <= not b or a;
    layer4_outputs(2235) <= not (a xor b);
    layer4_outputs(2236) <= not a;
    layer4_outputs(2237) <= a and b;
    layer4_outputs(2238) <= b;
    layer4_outputs(2239) <= b;
    layer4_outputs(2240) <= b;
    layer4_outputs(2241) <= not a;
    layer4_outputs(2242) <= a or b;
    layer4_outputs(2243) <= a and b;
    layer4_outputs(2244) <= not a;
    layer4_outputs(2245) <= not a;
    layer4_outputs(2246) <= not b;
    layer4_outputs(2247) <= b;
    layer4_outputs(2248) <= b;
    layer4_outputs(2249) <= a and not b;
    layer4_outputs(2250) <= 1'b0;
    layer4_outputs(2251) <= not b or a;
    layer4_outputs(2252) <= 1'b0;
    layer4_outputs(2253) <= a or b;
    layer4_outputs(2254) <= a and not b;
    layer4_outputs(2255) <= a;
    layer4_outputs(2256) <= not (a or b);
    layer4_outputs(2257) <= 1'b1;
    layer4_outputs(2258) <= not (a or b);
    layer4_outputs(2259) <= not (a or b);
    layer4_outputs(2260) <= not a or b;
    layer4_outputs(2261) <= 1'b0;
    layer4_outputs(2262) <= b;
    layer4_outputs(2263) <= not (a and b);
    layer4_outputs(2264) <= a and not b;
    layer4_outputs(2265) <= not a or b;
    layer4_outputs(2266) <= not (a or b);
    layer4_outputs(2267) <= a and b;
    layer4_outputs(2268) <= not b;
    layer4_outputs(2269) <= not b or a;
    layer4_outputs(2270) <= not a;
    layer4_outputs(2271) <= a or b;
    layer4_outputs(2272) <= a or b;
    layer4_outputs(2273) <= 1'b1;
    layer4_outputs(2274) <= b and not a;
    layer4_outputs(2275) <= 1'b1;
    layer4_outputs(2276) <= 1'b1;
    layer4_outputs(2277) <= 1'b1;
    layer4_outputs(2278) <= b and not a;
    layer4_outputs(2279) <= not b;
    layer4_outputs(2280) <= a;
    layer4_outputs(2281) <= not (a and b);
    layer4_outputs(2282) <= not a or b;
    layer4_outputs(2283) <= b and not a;
    layer4_outputs(2284) <= a and b;
    layer4_outputs(2285) <= not (a xor b);
    layer4_outputs(2286) <= not (a or b);
    layer4_outputs(2287) <= not a;
    layer4_outputs(2288) <= 1'b1;
    layer4_outputs(2289) <= a or b;
    layer4_outputs(2290) <= a and not b;
    layer4_outputs(2291) <= a and b;
    layer4_outputs(2292) <= not b or a;
    layer4_outputs(2293) <= not b;
    layer4_outputs(2294) <= a and b;
    layer4_outputs(2295) <= not (a and b);
    layer4_outputs(2296) <= a or b;
    layer4_outputs(2297) <= a;
    layer4_outputs(2298) <= 1'b1;
    layer4_outputs(2299) <= a and b;
    layer4_outputs(2300) <= not a;
    layer4_outputs(2301) <= b and not a;
    layer4_outputs(2302) <= not (a and b);
    layer4_outputs(2303) <= not a;
    layer4_outputs(2304) <= a or b;
    layer4_outputs(2305) <= not a or b;
    layer4_outputs(2306) <= not b;
    layer4_outputs(2307) <= not a;
    layer4_outputs(2308) <= b;
    layer4_outputs(2309) <= b and not a;
    layer4_outputs(2310) <= b;
    layer4_outputs(2311) <= b;
    layer4_outputs(2312) <= 1'b0;
    layer4_outputs(2313) <= 1'b0;
    layer4_outputs(2314) <= b and not a;
    layer4_outputs(2315) <= a;
    layer4_outputs(2316) <= a;
    layer4_outputs(2317) <= a and not b;
    layer4_outputs(2318) <= a and b;
    layer4_outputs(2319) <= 1'b1;
    layer4_outputs(2320) <= b and not a;
    layer4_outputs(2321) <= a;
    layer4_outputs(2322) <= b and not a;
    layer4_outputs(2323) <= 1'b0;
    layer4_outputs(2324) <= a;
    layer4_outputs(2325) <= not (a and b);
    layer4_outputs(2326) <= not (a and b);
    layer4_outputs(2327) <= b and not a;
    layer4_outputs(2328) <= b;
    layer4_outputs(2329) <= b;
    layer4_outputs(2330) <= a xor b;
    layer4_outputs(2331) <= not b;
    layer4_outputs(2332) <= not b;
    layer4_outputs(2333) <= not b;
    layer4_outputs(2334) <= a and not b;
    layer4_outputs(2335) <= a and b;
    layer4_outputs(2336) <= not (a or b);
    layer4_outputs(2337) <= 1'b0;
    layer4_outputs(2338) <= a or b;
    layer4_outputs(2339) <= b and not a;
    layer4_outputs(2340) <= not b;
    layer4_outputs(2341) <= a and not b;
    layer4_outputs(2342) <= a and b;
    layer4_outputs(2343) <= 1'b1;
    layer4_outputs(2344) <= 1'b1;
    layer4_outputs(2345) <= a;
    layer4_outputs(2346) <= 1'b1;
    layer4_outputs(2347) <= b;
    layer4_outputs(2348) <= a and not b;
    layer4_outputs(2349) <= b;
    layer4_outputs(2350) <= a or b;
    layer4_outputs(2351) <= not b;
    layer4_outputs(2352) <= a and not b;
    layer4_outputs(2353) <= not a or b;
    layer4_outputs(2354) <= not (a and b);
    layer4_outputs(2355) <= a and not b;
    layer4_outputs(2356) <= not b;
    layer4_outputs(2357) <= not a;
    layer4_outputs(2358) <= 1'b0;
    layer4_outputs(2359) <= not b;
    layer4_outputs(2360) <= a and not b;
    layer4_outputs(2361) <= not a;
    layer4_outputs(2362) <= not b;
    layer4_outputs(2363) <= not (a and b);
    layer4_outputs(2364) <= 1'b0;
    layer4_outputs(2365) <= a and not b;
    layer4_outputs(2366) <= not a or b;
    layer4_outputs(2367) <= not (a or b);
    layer4_outputs(2368) <= b and not a;
    layer4_outputs(2369) <= not a or b;
    layer4_outputs(2370) <= 1'b1;
    layer4_outputs(2371) <= a and b;
    layer4_outputs(2372) <= not (a or b);
    layer4_outputs(2373) <= not (a xor b);
    layer4_outputs(2374) <= not b or a;
    layer4_outputs(2375) <= b and not a;
    layer4_outputs(2376) <= not a;
    layer4_outputs(2377) <= not a or b;
    layer4_outputs(2378) <= a and not b;
    layer4_outputs(2379) <= not b;
    layer4_outputs(2380) <= not (a or b);
    layer4_outputs(2381) <= not b or a;
    layer4_outputs(2382) <= a and not b;
    layer4_outputs(2383) <= 1'b0;
    layer4_outputs(2384) <= b;
    layer4_outputs(2385) <= not b;
    layer4_outputs(2386) <= not a or b;
    layer4_outputs(2387) <= not b or a;
    layer4_outputs(2388) <= not a or b;
    layer4_outputs(2389) <= not (a and b);
    layer4_outputs(2390) <= not (a or b);
    layer4_outputs(2391) <= not b;
    layer4_outputs(2392) <= not b;
    layer4_outputs(2393) <= 1'b1;
    layer4_outputs(2394) <= not a;
    layer4_outputs(2395) <= not b;
    layer4_outputs(2396) <= not (a and b);
    layer4_outputs(2397) <= not a;
    layer4_outputs(2398) <= a and not b;
    layer4_outputs(2399) <= not a;
    layer4_outputs(2400) <= b and not a;
    layer4_outputs(2401) <= 1'b1;
    layer4_outputs(2402) <= not a or b;
    layer4_outputs(2403) <= 1'b0;
    layer4_outputs(2404) <= not a;
    layer4_outputs(2405) <= a xor b;
    layer4_outputs(2406) <= not b or a;
    layer4_outputs(2407) <= a and b;
    layer4_outputs(2408) <= not a or b;
    layer4_outputs(2409) <= not a or b;
    layer4_outputs(2410) <= a or b;
    layer4_outputs(2411) <= a and not b;
    layer4_outputs(2412) <= a;
    layer4_outputs(2413) <= a and b;
    layer4_outputs(2414) <= not (a and b);
    layer4_outputs(2415) <= not a;
    layer4_outputs(2416) <= b and not a;
    layer4_outputs(2417) <= b;
    layer4_outputs(2418) <= not (a or b);
    layer4_outputs(2419) <= 1'b1;
    layer4_outputs(2420) <= not (a and b);
    layer4_outputs(2421) <= not b;
    layer4_outputs(2422) <= a and not b;
    layer4_outputs(2423) <= not a;
    layer4_outputs(2424) <= not a;
    layer4_outputs(2425) <= not (a or b);
    layer4_outputs(2426) <= a and b;
    layer4_outputs(2427) <= not a;
    layer4_outputs(2428) <= 1'b1;
    layer4_outputs(2429) <= not b;
    layer4_outputs(2430) <= a;
    layer4_outputs(2431) <= 1'b0;
    layer4_outputs(2432) <= not (a or b);
    layer4_outputs(2433) <= not b;
    layer4_outputs(2434) <= not (a and b);
    layer4_outputs(2435) <= not b;
    layer4_outputs(2436) <= not a or b;
    layer4_outputs(2437) <= a or b;
    layer4_outputs(2438) <= 1'b0;
    layer4_outputs(2439) <= not a;
    layer4_outputs(2440) <= not a or b;
    layer4_outputs(2441) <= a and b;
    layer4_outputs(2442) <= a and not b;
    layer4_outputs(2443) <= not b;
    layer4_outputs(2444) <= not a;
    layer4_outputs(2445) <= not a or b;
    layer4_outputs(2446) <= not b;
    layer4_outputs(2447) <= a and not b;
    layer4_outputs(2448) <= not b;
    layer4_outputs(2449) <= a or b;
    layer4_outputs(2450) <= 1'b1;
    layer4_outputs(2451) <= a or b;
    layer4_outputs(2452) <= 1'b0;
    layer4_outputs(2453) <= not (a and b);
    layer4_outputs(2454) <= not b or a;
    layer4_outputs(2455) <= not (a and b);
    layer4_outputs(2456) <= not a or b;
    layer4_outputs(2457) <= a or b;
    layer4_outputs(2458) <= not b or a;
    layer4_outputs(2459) <= 1'b0;
    layer4_outputs(2460) <= not a;
    layer4_outputs(2461) <= not b;
    layer4_outputs(2462) <= a or b;
    layer4_outputs(2463) <= not b or a;
    layer4_outputs(2464) <= b;
    layer4_outputs(2465) <= not a;
    layer4_outputs(2466) <= a and not b;
    layer4_outputs(2467) <= 1'b0;
    layer4_outputs(2468) <= b;
    layer4_outputs(2469) <= a and b;
    layer4_outputs(2470) <= not (a and b);
    layer4_outputs(2471) <= not b or a;
    layer4_outputs(2472) <= a and b;
    layer4_outputs(2473) <= not (a xor b);
    layer4_outputs(2474) <= not b;
    layer4_outputs(2475) <= not a;
    layer4_outputs(2476) <= not (a and b);
    layer4_outputs(2477) <= a and b;
    layer4_outputs(2478) <= a;
    layer4_outputs(2479) <= 1'b0;
    layer4_outputs(2480) <= 1'b1;
    layer4_outputs(2481) <= not (a and b);
    layer4_outputs(2482) <= not a or b;
    layer4_outputs(2483) <= b and not a;
    layer4_outputs(2484) <= not b or a;
    layer4_outputs(2485) <= not a;
    layer4_outputs(2486) <= not b;
    layer4_outputs(2487) <= not a or b;
    layer4_outputs(2488) <= not b or a;
    layer4_outputs(2489) <= not b or a;
    layer4_outputs(2490) <= a or b;
    layer4_outputs(2491) <= a and not b;
    layer4_outputs(2492) <= not b;
    layer4_outputs(2493) <= not b or a;
    layer4_outputs(2494) <= a;
    layer4_outputs(2495) <= not b;
    layer4_outputs(2496) <= not (a or b);
    layer4_outputs(2497) <= a and b;
    layer4_outputs(2498) <= not (a or b);
    layer4_outputs(2499) <= not (a or b);
    layer4_outputs(2500) <= not a;
    layer4_outputs(2501) <= not a;
    layer4_outputs(2502) <= not b;
    layer4_outputs(2503) <= not b or a;
    layer4_outputs(2504) <= not (a and b);
    layer4_outputs(2505) <= b and not a;
    layer4_outputs(2506) <= a and not b;
    layer4_outputs(2507) <= not a;
    layer4_outputs(2508) <= b and not a;
    layer4_outputs(2509) <= a and b;
    layer4_outputs(2510) <= a;
    layer4_outputs(2511) <= not a;
    layer4_outputs(2512) <= b and not a;
    layer4_outputs(2513) <= a and not b;
    layer4_outputs(2514) <= not b;
    layer4_outputs(2515) <= 1'b0;
    layer4_outputs(2516) <= b and not a;
    layer4_outputs(2517) <= 1'b1;
    layer4_outputs(2518) <= not a;
    layer4_outputs(2519) <= not (a and b);
    layer4_outputs(2520) <= b;
    layer4_outputs(2521) <= not b;
    layer4_outputs(2522) <= a and not b;
    layer4_outputs(2523) <= not (a or b);
    layer4_outputs(2524) <= not (a xor b);
    layer4_outputs(2525) <= not a;
    layer4_outputs(2526) <= a;
    layer4_outputs(2527) <= not a or b;
    layer4_outputs(2528) <= not (a or b);
    layer4_outputs(2529) <= not (a or b);
    layer4_outputs(2530) <= a;
    layer4_outputs(2531) <= not a;
    layer4_outputs(2532) <= not b or a;
    layer4_outputs(2533) <= not a;
    layer4_outputs(2534) <= b;
    layer4_outputs(2535) <= b;
    layer4_outputs(2536) <= not b;
    layer4_outputs(2537) <= not a or b;
    layer4_outputs(2538) <= not a or b;
    layer4_outputs(2539) <= a and not b;
    layer4_outputs(2540) <= a and b;
    layer4_outputs(2541) <= not a;
    layer4_outputs(2542) <= a or b;
    layer4_outputs(2543) <= not (a or b);
    layer4_outputs(2544) <= 1'b0;
    layer4_outputs(2545) <= not (a or b);
    layer4_outputs(2546) <= not a;
    layer4_outputs(2547) <= 1'b1;
    layer4_outputs(2548) <= a and b;
    layer4_outputs(2549) <= a and b;
    layer4_outputs(2550) <= not a;
    layer4_outputs(2551) <= a and not b;
    layer4_outputs(2552) <= b;
    layer4_outputs(2553) <= a;
    layer4_outputs(2554) <= not b or a;
    layer4_outputs(2555) <= 1'b1;
    layer4_outputs(2556) <= a and b;
    layer4_outputs(2557) <= not (a xor b);
    layer4_outputs(2558) <= a;
    layer4_outputs(2559) <= b;
    layer5_outputs(0) <= a;
    layer5_outputs(1) <= not (a and b);
    layer5_outputs(2) <= not a;
    layer5_outputs(3) <= not a or b;
    layer5_outputs(4) <= not (a and b);
    layer5_outputs(5) <= a;
    layer5_outputs(6) <= b and not a;
    layer5_outputs(7) <= b and not a;
    layer5_outputs(8) <= 1'b1;
    layer5_outputs(9) <= a and b;
    layer5_outputs(10) <= a or b;
    layer5_outputs(11) <= a or b;
    layer5_outputs(12) <= b and not a;
    layer5_outputs(13) <= 1'b1;
    layer5_outputs(14) <= not b or a;
    layer5_outputs(15) <= a and not b;
    layer5_outputs(16) <= not b;
    layer5_outputs(17) <= b and not a;
    layer5_outputs(18) <= not a;
    layer5_outputs(19) <= 1'b0;
    layer5_outputs(20) <= not (a and b);
    layer5_outputs(21) <= not a;
    layer5_outputs(22) <= not b;
    layer5_outputs(23) <= not a;
    layer5_outputs(24) <= a;
    layer5_outputs(25) <= a xor b;
    layer5_outputs(26) <= 1'b0;
    layer5_outputs(27) <= not a or b;
    layer5_outputs(28) <= not b;
    layer5_outputs(29) <= a and b;
    layer5_outputs(30) <= not a;
    layer5_outputs(31) <= not (a xor b);
    layer5_outputs(32) <= b and not a;
    layer5_outputs(33) <= not b;
    layer5_outputs(34) <= a and not b;
    layer5_outputs(35) <= not a;
    layer5_outputs(36) <= not b;
    layer5_outputs(37) <= not a;
    layer5_outputs(38) <= 1'b0;
    layer5_outputs(39) <= not (a or b);
    layer5_outputs(40) <= a and b;
    layer5_outputs(41) <= not b or a;
    layer5_outputs(42) <= not b or a;
    layer5_outputs(43) <= b;
    layer5_outputs(44) <= a and not b;
    layer5_outputs(45) <= a xor b;
    layer5_outputs(46) <= 1'b1;
    layer5_outputs(47) <= not a;
    layer5_outputs(48) <= 1'b0;
    layer5_outputs(49) <= 1'b1;
    layer5_outputs(50) <= not a;
    layer5_outputs(51) <= not b;
    layer5_outputs(52) <= b;
    layer5_outputs(53) <= not a;
    layer5_outputs(54) <= a and not b;
    layer5_outputs(55) <= not a or b;
    layer5_outputs(56) <= a and b;
    layer5_outputs(57) <= b;
    layer5_outputs(58) <= a and b;
    layer5_outputs(59) <= b;
    layer5_outputs(60) <= 1'b1;
    layer5_outputs(61) <= not a;
    layer5_outputs(62) <= a;
    layer5_outputs(63) <= b and not a;
    layer5_outputs(64) <= a or b;
    layer5_outputs(65) <= not b or a;
    layer5_outputs(66) <= a and b;
    layer5_outputs(67) <= a and not b;
    layer5_outputs(68) <= a and b;
    layer5_outputs(69) <= not (a or b);
    layer5_outputs(70) <= not b or a;
    layer5_outputs(71) <= a and not b;
    layer5_outputs(72) <= not a;
    layer5_outputs(73) <= not (a and b);
    layer5_outputs(74) <= not (a or b);
    layer5_outputs(75) <= a and not b;
    layer5_outputs(76) <= a or b;
    layer5_outputs(77) <= not a or b;
    layer5_outputs(78) <= not (a or b);
    layer5_outputs(79) <= not (a and b);
    layer5_outputs(80) <= 1'b0;
    layer5_outputs(81) <= not a;
    layer5_outputs(82) <= b and not a;
    layer5_outputs(83) <= not (a or b);
    layer5_outputs(84) <= not a;
    layer5_outputs(85) <= not b or a;
    layer5_outputs(86) <= 1'b1;
    layer5_outputs(87) <= a or b;
    layer5_outputs(88) <= 1'b1;
    layer5_outputs(89) <= a;
    layer5_outputs(90) <= a and b;
    layer5_outputs(91) <= not a or b;
    layer5_outputs(92) <= not (a or b);
    layer5_outputs(93) <= not a or b;
    layer5_outputs(94) <= a and b;
    layer5_outputs(95) <= a or b;
    layer5_outputs(96) <= not a or b;
    layer5_outputs(97) <= not a;
    layer5_outputs(98) <= b and not a;
    layer5_outputs(99) <= a;
    layer5_outputs(100) <= a;
    layer5_outputs(101) <= not a or b;
    layer5_outputs(102) <= not a;
    layer5_outputs(103) <= not b;
    layer5_outputs(104) <= not a;
    layer5_outputs(105) <= not a;
    layer5_outputs(106) <= b and not a;
    layer5_outputs(107) <= 1'b1;
    layer5_outputs(108) <= not b;
    layer5_outputs(109) <= not b;
    layer5_outputs(110) <= not a or b;
    layer5_outputs(111) <= not b or a;
    layer5_outputs(112) <= a and b;
    layer5_outputs(113) <= 1'b1;
    layer5_outputs(114) <= not (a and b);
    layer5_outputs(115) <= a and not b;
    layer5_outputs(116) <= 1'b0;
    layer5_outputs(117) <= a or b;
    layer5_outputs(118) <= a;
    layer5_outputs(119) <= not (a and b);
    layer5_outputs(120) <= 1'b1;
    layer5_outputs(121) <= 1'b0;
    layer5_outputs(122) <= not b;
    layer5_outputs(123) <= not b;
    layer5_outputs(124) <= b;
    layer5_outputs(125) <= a and b;
    layer5_outputs(126) <= b;
    layer5_outputs(127) <= not (a and b);
    layer5_outputs(128) <= not a or b;
    layer5_outputs(129) <= not (a and b);
    layer5_outputs(130) <= a or b;
    layer5_outputs(131) <= not a or b;
    layer5_outputs(132) <= 1'b0;
    layer5_outputs(133) <= a and not b;
    layer5_outputs(134) <= not (a and b);
    layer5_outputs(135) <= 1'b0;
    layer5_outputs(136) <= a xor b;
    layer5_outputs(137) <= not b;
    layer5_outputs(138) <= not (a or b);
    layer5_outputs(139) <= 1'b1;
    layer5_outputs(140) <= not (a and b);
    layer5_outputs(141) <= 1'b0;
    layer5_outputs(142) <= not (a or b);
    layer5_outputs(143) <= a xor b;
    layer5_outputs(144) <= not a;
    layer5_outputs(145) <= 1'b1;
    layer5_outputs(146) <= a and b;
    layer5_outputs(147) <= not a or b;
    layer5_outputs(148) <= not a or b;
    layer5_outputs(149) <= not (a or b);
    layer5_outputs(150) <= a and not b;
    layer5_outputs(151) <= not b;
    layer5_outputs(152) <= a and not b;
    layer5_outputs(153) <= not a or b;
    layer5_outputs(154) <= not b or a;
    layer5_outputs(155) <= b;
    layer5_outputs(156) <= not (a or b);
    layer5_outputs(157) <= not a;
    layer5_outputs(158) <= not a or b;
    layer5_outputs(159) <= not (a or b);
    layer5_outputs(160) <= not (a and b);
    layer5_outputs(161) <= not a or b;
    layer5_outputs(162) <= a and b;
    layer5_outputs(163) <= b and not a;
    layer5_outputs(164) <= a;
    layer5_outputs(165) <= not a or b;
    layer5_outputs(166) <= b and not a;
    layer5_outputs(167) <= not b;
    layer5_outputs(168) <= a or b;
    layer5_outputs(169) <= not b;
    layer5_outputs(170) <= b;
    layer5_outputs(171) <= not b;
    layer5_outputs(172) <= a;
    layer5_outputs(173) <= a;
    layer5_outputs(174) <= not b;
    layer5_outputs(175) <= not a or b;
    layer5_outputs(176) <= 1'b1;
    layer5_outputs(177) <= 1'b0;
    layer5_outputs(178) <= 1'b1;
    layer5_outputs(179) <= a and not b;
    layer5_outputs(180) <= a;
    layer5_outputs(181) <= not b or a;
    layer5_outputs(182) <= not b;
    layer5_outputs(183) <= not a or b;
    layer5_outputs(184) <= a;
    layer5_outputs(185) <= a;
    layer5_outputs(186) <= b;
    layer5_outputs(187) <= not (a or b);
    layer5_outputs(188) <= not b or a;
    layer5_outputs(189) <= 1'b0;
    layer5_outputs(190) <= 1'b1;
    layer5_outputs(191) <= a;
    layer5_outputs(192) <= b;
    layer5_outputs(193) <= b;
    layer5_outputs(194) <= a and not b;
    layer5_outputs(195) <= not a or b;
    layer5_outputs(196) <= not b;
    layer5_outputs(197) <= a and b;
    layer5_outputs(198) <= not a;
    layer5_outputs(199) <= not (a or b);
    layer5_outputs(200) <= a;
    layer5_outputs(201) <= a and b;
    layer5_outputs(202) <= b;
    layer5_outputs(203) <= not b;
    layer5_outputs(204) <= not (a and b);
    layer5_outputs(205) <= not b;
    layer5_outputs(206) <= not b or a;
    layer5_outputs(207) <= a or b;
    layer5_outputs(208) <= b;
    layer5_outputs(209) <= not (a and b);
    layer5_outputs(210) <= a and b;
    layer5_outputs(211) <= not (a and b);
    layer5_outputs(212) <= 1'b0;
    layer5_outputs(213) <= 1'b1;
    layer5_outputs(214) <= a and b;
    layer5_outputs(215) <= not a;
    layer5_outputs(216) <= not (a and b);
    layer5_outputs(217) <= not b;
    layer5_outputs(218) <= a;
    layer5_outputs(219) <= a or b;
    layer5_outputs(220) <= not a;
    layer5_outputs(221) <= b;
    layer5_outputs(222) <= not a;
    layer5_outputs(223) <= a or b;
    layer5_outputs(224) <= a and not b;
    layer5_outputs(225) <= a and not b;
    layer5_outputs(226) <= b;
    layer5_outputs(227) <= not (a or b);
    layer5_outputs(228) <= b;
    layer5_outputs(229) <= not (a or b);
    layer5_outputs(230) <= 1'b1;
    layer5_outputs(231) <= b;
    layer5_outputs(232) <= a and not b;
    layer5_outputs(233) <= a and b;
    layer5_outputs(234) <= a and b;
    layer5_outputs(235) <= not a;
    layer5_outputs(236) <= a xor b;
    layer5_outputs(237) <= b;
    layer5_outputs(238) <= not b or a;
    layer5_outputs(239) <= not b;
    layer5_outputs(240) <= not a;
    layer5_outputs(241) <= a;
    layer5_outputs(242) <= b;
    layer5_outputs(243) <= not b or a;
    layer5_outputs(244) <= not a or b;
    layer5_outputs(245) <= a or b;
    layer5_outputs(246) <= not a or b;
    layer5_outputs(247) <= b;
    layer5_outputs(248) <= a or b;
    layer5_outputs(249) <= not (a and b);
    layer5_outputs(250) <= a and not b;
    layer5_outputs(251) <= not b;
    layer5_outputs(252) <= not a;
    layer5_outputs(253) <= not (a or b);
    layer5_outputs(254) <= a or b;
    layer5_outputs(255) <= b and not a;
    layer5_outputs(256) <= a and not b;
    layer5_outputs(257) <= b;
    layer5_outputs(258) <= a and not b;
    layer5_outputs(259) <= 1'b1;
    layer5_outputs(260) <= a;
    layer5_outputs(261) <= not b;
    layer5_outputs(262) <= not b or a;
    layer5_outputs(263) <= 1'b0;
    layer5_outputs(264) <= a and b;
    layer5_outputs(265) <= a;
    layer5_outputs(266) <= a or b;
    layer5_outputs(267) <= a and not b;
    layer5_outputs(268) <= not b or a;
    layer5_outputs(269) <= b and not a;
    layer5_outputs(270) <= a;
    layer5_outputs(271) <= a and not b;
    layer5_outputs(272) <= b;
    layer5_outputs(273) <= a;
    layer5_outputs(274) <= a;
    layer5_outputs(275) <= b;
    layer5_outputs(276) <= not a or b;
    layer5_outputs(277) <= not (a and b);
    layer5_outputs(278) <= not (a xor b);
    layer5_outputs(279) <= 1'b1;
    layer5_outputs(280) <= not a or b;
    layer5_outputs(281) <= not a or b;
    layer5_outputs(282) <= not (a and b);
    layer5_outputs(283) <= not a or b;
    layer5_outputs(284) <= not b or a;
    layer5_outputs(285) <= 1'b1;
    layer5_outputs(286) <= not a or b;
    layer5_outputs(287) <= b;
    layer5_outputs(288) <= a or b;
    layer5_outputs(289) <= not a;
    layer5_outputs(290) <= a and not b;
    layer5_outputs(291) <= not (a or b);
    layer5_outputs(292) <= not a;
    layer5_outputs(293) <= not (a or b);
    layer5_outputs(294) <= b and not a;
    layer5_outputs(295) <= b and not a;
    layer5_outputs(296) <= not a;
    layer5_outputs(297) <= 1'b1;
    layer5_outputs(298) <= not b;
    layer5_outputs(299) <= a and not b;
    layer5_outputs(300) <= not (a and b);
    layer5_outputs(301) <= not a;
    layer5_outputs(302) <= not a;
    layer5_outputs(303) <= not a;
    layer5_outputs(304) <= not (a xor b);
    layer5_outputs(305) <= not b or a;
    layer5_outputs(306) <= not b;
    layer5_outputs(307) <= not (a or b);
    layer5_outputs(308) <= a;
    layer5_outputs(309) <= not a or b;
    layer5_outputs(310) <= 1'b0;
    layer5_outputs(311) <= a xor b;
    layer5_outputs(312) <= a and b;
    layer5_outputs(313) <= a;
    layer5_outputs(314) <= a;
    layer5_outputs(315) <= not (a and b);
    layer5_outputs(316) <= a or b;
    layer5_outputs(317) <= not (a or b);
    layer5_outputs(318) <= not a;
    layer5_outputs(319) <= a xor b;
    layer5_outputs(320) <= a or b;
    layer5_outputs(321) <= not a;
    layer5_outputs(322) <= not a or b;
    layer5_outputs(323) <= not (a xor b);
    layer5_outputs(324) <= b;
    layer5_outputs(325) <= a or b;
    layer5_outputs(326) <= b and not a;
    layer5_outputs(327) <= not b;
    layer5_outputs(328) <= b;
    layer5_outputs(329) <= not b or a;
    layer5_outputs(330) <= not a;
    layer5_outputs(331) <= not a or b;
    layer5_outputs(332) <= b and not a;
    layer5_outputs(333) <= not b or a;
    layer5_outputs(334) <= 1'b0;
    layer5_outputs(335) <= not (a or b);
    layer5_outputs(336) <= a;
    layer5_outputs(337) <= not a or b;
    layer5_outputs(338) <= a or b;
    layer5_outputs(339) <= a and b;
    layer5_outputs(340) <= not b;
    layer5_outputs(341) <= a and b;
    layer5_outputs(342) <= not (a xor b);
    layer5_outputs(343) <= not (a xor b);
    layer5_outputs(344) <= b;
    layer5_outputs(345) <= b and not a;
    layer5_outputs(346) <= not b;
    layer5_outputs(347) <= a;
    layer5_outputs(348) <= 1'b0;
    layer5_outputs(349) <= not a or b;
    layer5_outputs(350) <= not b;
    layer5_outputs(351) <= b;
    layer5_outputs(352) <= b;
    layer5_outputs(353) <= b;
    layer5_outputs(354) <= b;
    layer5_outputs(355) <= b and not a;
    layer5_outputs(356) <= not b;
    layer5_outputs(357) <= 1'b1;
    layer5_outputs(358) <= b;
    layer5_outputs(359) <= b;
    layer5_outputs(360) <= not a;
    layer5_outputs(361) <= 1'b1;
    layer5_outputs(362) <= a or b;
    layer5_outputs(363) <= b;
    layer5_outputs(364) <= not a;
    layer5_outputs(365) <= not b;
    layer5_outputs(366) <= not (a or b);
    layer5_outputs(367) <= not a;
    layer5_outputs(368) <= not b;
    layer5_outputs(369) <= b;
    layer5_outputs(370) <= 1'b1;
    layer5_outputs(371) <= not a or b;
    layer5_outputs(372) <= a and not b;
    layer5_outputs(373) <= not (a and b);
    layer5_outputs(374) <= not a;
    layer5_outputs(375) <= not a;
    layer5_outputs(376) <= not b or a;
    layer5_outputs(377) <= not b or a;
    layer5_outputs(378) <= not (a or b);
    layer5_outputs(379) <= not b;
    layer5_outputs(380) <= not b or a;
    layer5_outputs(381) <= not a;
    layer5_outputs(382) <= not (a or b);
    layer5_outputs(383) <= 1'b1;
    layer5_outputs(384) <= not a;
    layer5_outputs(385) <= not (a and b);
    layer5_outputs(386) <= not a;
    layer5_outputs(387) <= b;
    layer5_outputs(388) <= not b or a;
    layer5_outputs(389) <= a;
    layer5_outputs(390) <= not (a or b);
    layer5_outputs(391) <= a;
    layer5_outputs(392) <= a or b;
    layer5_outputs(393) <= not b;
    layer5_outputs(394) <= b;
    layer5_outputs(395) <= a xor b;
    layer5_outputs(396) <= b and not a;
    layer5_outputs(397) <= not b;
    layer5_outputs(398) <= not (a or b);
    layer5_outputs(399) <= not b;
    layer5_outputs(400) <= a xor b;
    layer5_outputs(401) <= b;
    layer5_outputs(402) <= not b;
    layer5_outputs(403) <= not a;
    layer5_outputs(404) <= 1'b0;
    layer5_outputs(405) <= a;
    layer5_outputs(406) <= not (a or b);
    layer5_outputs(407) <= b and not a;
    layer5_outputs(408) <= not a;
    layer5_outputs(409) <= not b;
    layer5_outputs(410) <= not b or a;
    layer5_outputs(411) <= not b or a;
    layer5_outputs(412) <= 1'b0;
    layer5_outputs(413) <= not (a or b);
    layer5_outputs(414) <= not (a or b);
    layer5_outputs(415) <= 1'b0;
    layer5_outputs(416) <= not a;
    layer5_outputs(417) <= not a or b;
    layer5_outputs(418) <= not a;
    layer5_outputs(419) <= a;
    layer5_outputs(420) <= not (a xor b);
    layer5_outputs(421) <= not b or a;
    layer5_outputs(422) <= not (a or b);
    layer5_outputs(423) <= not b or a;
    layer5_outputs(424) <= a;
    layer5_outputs(425) <= 1'b0;
    layer5_outputs(426) <= a or b;
    layer5_outputs(427) <= 1'b1;
    layer5_outputs(428) <= not a or b;
    layer5_outputs(429) <= a and b;
    layer5_outputs(430) <= a and not b;
    layer5_outputs(431) <= b;
    layer5_outputs(432) <= not a;
    layer5_outputs(433) <= a and not b;
    layer5_outputs(434) <= a and not b;
    layer5_outputs(435) <= not b or a;
    layer5_outputs(436) <= not a;
    layer5_outputs(437) <= not (a or b);
    layer5_outputs(438) <= not a;
    layer5_outputs(439) <= not a;
    layer5_outputs(440) <= not (a xor b);
    layer5_outputs(441) <= not b;
    layer5_outputs(442) <= a and not b;
    layer5_outputs(443) <= a or b;
    layer5_outputs(444) <= not b;
    layer5_outputs(445) <= not a;
    layer5_outputs(446) <= not b or a;
    layer5_outputs(447) <= a or b;
    layer5_outputs(448) <= a and not b;
    layer5_outputs(449) <= not b;
    layer5_outputs(450) <= not b;
    layer5_outputs(451) <= not a;
    layer5_outputs(452) <= not a;
    layer5_outputs(453) <= a and not b;
    layer5_outputs(454) <= not b or a;
    layer5_outputs(455) <= b;
    layer5_outputs(456) <= not (a or b);
    layer5_outputs(457) <= b and not a;
    layer5_outputs(458) <= b;
    layer5_outputs(459) <= not a or b;
    layer5_outputs(460) <= not b;
    layer5_outputs(461) <= a;
    layer5_outputs(462) <= not a;
    layer5_outputs(463) <= not b or a;
    layer5_outputs(464) <= not a;
    layer5_outputs(465) <= not b;
    layer5_outputs(466) <= not a;
    layer5_outputs(467) <= not b;
    layer5_outputs(468) <= a and b;
    layer5_outputs(469) <= 1'b1;
    layer5_outputs(470) <= a or b;
    layer5_outputs(471) <= b and not a;
    layer5_outputs(472) <= not b;
    layer5_outputs(473) <= 1'b0;
    layer5_outputs(474) <= not (a or b);
    layer5_outputs(475) <= not b or a;
    layer5_outputs(476) <= a or b;
    layer5_outputs(477) <= b;
    layer5_outputs(478) <= a or b;
    layer5_outputs(479) <= 1'b1;
    layer5_outputs(480) <= not a;
    layer5_outputs(481) <= b;
    layer5_outputs(482) <= b and not a;
    layer5_outputs(483) <= not a;
    layer5_outputs(484) <= a and b;
    layer5_outputs(485) <= 1'b0;
    layer5_outputs(486) <= a;
    layer5_outputs(487) <= a;
    layer5_outputs(488) <= not a;
    layer5_outputs(489) <= not b;
    layer5_outputs(490) <= not a or b;
    layer5_outputs(491) <= a and b;
    layer5_outputs(492) <= b and not a;
    layer5_outputs(493) <= not b;
    layer5_outputs(494) <= b and not a;
    layer5_outputs(495) <= a;
    layer5_outputs(496) <= b and not a;
    layer5_outputs(497) <= b;
    layer5_outputs(498) <= 1'b0;
    layer5_outputs(499) <= not b;
    layer5_outputs(500) <= not b or a;
    layer5_outputs(501) <= b;
    layer5_outputs(502) <= not b;
    layer5_outputs(503) <= a;
    layer5_outputs(504) <= not (a or b);
    layer5_outputs(505) <= not (a or b);
    layer5_outputs(506) <= not b;
    layer5_outputs(507) <= not (a and b);
    layer5_outputs(508) <= a;
    layer5_outputs(509) <= not a;
    layer5_outputs(510) <= a;
    layer5_outputs(511) <= a and b;
    layer5_outputs(512) <= not (a or b);
    layer5_outputs(513) <= a and not b;
    layer5_outputs(514) <= 1'b0;
    layer5_outputs(515) <= a and b;
    layer5_outputs(516) <= not a;
    layer5_outputs(517) <= a or b;
    layer5_outputs(518) <= not (a xor b);
    layer5_outputs(519) <= not b;
    layer5_outputs(520) <= not a or b;
    layer5_outputs(521) <= b;
    layer5_outputs(522) <= not (a and b);
    layer5_outputs(523) <= b;
    layer5_outputs(524) <= not a;
    layer5_outputs(525) <= a xor b;
    layer5_outputs(526) <= not b;
    layer5_outputs(527) <= not b or a;
    layer5_outputs(528) <= a or b;
    layer5_outputs(529) <= a and b;
    layer5_outputs(530) <= b;
    layer5_outputs(531) <= a;
    layer5_outputs(532) <= 1'b1;
    layer5_outputs(533) <= b;
    layer5_outputs(534) <= 1'b1;
    layer5_outputs(535) <= 1'b0;
    layer5_outputs(536) <= not b or a;
    layer5_outputs(537) <= not a or b;
    layer5_outputs(538) <= b and not a;
    layer5_outputs(539) <= b and not a;
    layer5_outputs(540) <= not b or a;
    layer5_outputs(541) <= a or b;
    layer5_outputs(542) <= not b or a;
    layer5_outputs(543) <= a or b;
    layer5_outputs(544) <= not b;
    layer5_outputs(545) <= not b or a;
    layer5_outputs(546) <= a and not b;
    layer5_outputs(547) <= a and not b;
    layer5_outputs(548) <= not a or b;
    layer5_outputs(549) <= not (a and b);
    layer5_outputs(550) <= a;
    layer5_outputs(551) <= not a or b;
    layer5_outputs(552) <= b;
    layer5_outputs(553) <= a;
    layer5_outputs(554) <= b and not a;
    layer5_outputs(555) <= b;
    layer5_outputs(556) <= a and b;
    layer5_outputs(557) <= not (a or b);
    layer5_outputs(558) <= not a;
    layer5_outputs(559) <= not (a and b);
    layer5_outputs(560) <= a and b;
    layer5_outputs(561) <= not b or a;
    layer5_outputs(562) <= not a or b;
    layer5_outputs(563) <= a and b;
    layer5_outputs(564) <= 1'b0;
    layer5_outputs(565) <= not a;
    layer5_outputs(566) <= a;
    layer5_outputs(567) <= a or b;
    layer5_outputs(568) <= not a;
    layer5_outputs(569) <= a or b;
    layer5_outputs(570) <= not a;
    layer5_outputs(571) <= not (a and b);
    layer5_outputs(572) <= a and b;
    layer5_outputs(573) <= not b;
    layer5_outputs(574) <= not a;
    layer5_outputs(575) <= a;
    layer5_outputs(576) <= 1'b0;
    layer5_outputs(577) <= a;
    layer5_outputs(578) <= not (a xor b);
    layer5_outputs(579) <= b;
    layer5_outputs(580) <= not a;
    layer5_outputs(581) <= a and b;
    layer5_outputs(582) <= not b;
    layer5_outputs(583) <= b and not a;
    layer5_outputs(584) <= b;
    layer5_outputs(585) <= not a or b;
    layer5_outputs(586) <= 1'b0;
    layer5_outputs(587) <= 1'b0;
    layer5_outputs(588) <= not a or b;
    layer5_outputs(589) <= not b or a;
    layer5_outputs(590) <= not (a or b);
    layer5_outputs(591) <= 1'b1;
    layer5_outputs(592) <= a;
    layer5_outputs(593) <= not (a and b);
    layer5_outputs(594) <= not (a xor b);
    layer5_outputs(595) <= b;
    layer5_outputs(596) <= not a;
    layer5_outputs(597) <= 1'b1;
    layer5_outputs(598) <= not b;
    layer5_outputs(599) <= not b;
    layer5_outputs(600) <= a and b;
    layer5_outputs(601) <= a and not b;
    layer5_outputs(602) <= a;
    layer5_outputs(603) <= a and b;
    layer5_outputs(604) <= a and not b;
    layer5_outputs(605) <= a and b;
    layer5_outputs(606) <= a;
    layer5_outputs(607) <= not a;
    layer5_outputs(608) <= b and not a;
    layer5_outputs(609) <= not b;
    layer5_outputs(610) <= a and b;
    layer5_outputs(611) <= not b or a;
    layer5_outputs(612) <= not (a and b);
    layer5_outputs(613) <= not b or a;
    layer5_outputs(614) <= not a or b;
    layer5_outputs(615) <= not (a or b);
    layer5_outputs(616) <= not (a xor b);
    layer5_outputs(617) <= a;
    layer5_outputs(618) <= 1'b0;
    layer5_outputs(619) <= a or b;
    layer5_outputs(620) <= not b;
    layer5_outputs(621) <= a;
    layer5_outputs(622) <= 1'b1;
    layer5_outputs(623) <= a and not b;
    layer5_outputs(624) <= not b;
    layer5_outputs(625) <= not a or b;
    layer5_outputs(626) <= not b;
    layer5_outputs(627) <= not (a or b);
    layer5_outputs(628) <= b;
    layer5_outputs(629) <= not a;
    layer5_outputs(630) <= not b;
    layer5_outputs(631) <= 1'b0;
    layer5_outputs(632) <= a xor b;
    layer5_outputs(633) <= b;
    layer5_outputs(634) <= a or b;
    layer5_outputs(635) <= 1'b0;
    layer5_outputs(636) <= not (a and b);
    layer5_outputs(637) <= not b;
    layer5_outputs(638) <= b and not a;
    layer5_outputs(639) <= a and b;
    layer5_outputs(640) <= 1'b1;
    layer5_outputs(641) <= b;
    layer5_outputs(642) <= b;
    layer5_outputs(643) <= a;
    layer5_outputs(644) <= not b;
    layer5_outputs(645) <= a and b;
    layer5_outputs(646) <= not (a and b);
    layer5_outputs(647) <= a;
    layer5_outputs(648) <= not a;
    layer5_outputs(649) <= a;
    layer5_outputs(650) <= not a or b;
    layer5_outputs(651) <= a;
    layer5_outputs(652) <= not a or b;
    layer5_outputs(653) <= not a or b;
    layer5_outputs(654) <= 1'b0;
    layer5_outputs(655) <= 1'b0;
    layer5_outputs(656) <= not b;
    layer5_outputs(657) <= not (a and b);
    layer5_outputs(658) <= a and b;
    layer5_outputs(659) <= not a or b;
    layer5_outputs(660) <= not a or b;
    layer5_outputs(661) <= b;
    layer5_outputs(662) <= not a;
    layer5_outputs(663) <= not (a xor b);
    layer5_outputs(664) <= not b;
    layer5_outputs(665) <= not a;
    layer5_outputs(666) <= 1'b0;
    layer5_outputs(667) <= not a;
    layer5_outputs(668) <= a or b;
    layer5_outputs(669) <= a and b;
    layer5_outputs(670) <= a and not b;
    layer5_outputs(671) <= 1'b0;
    layer5_outputs(672) <= not (a and b);
    layer5_outputs(673) <= not a;
    layer5_outputs(674) <= b and not a;
    layer5_outputs(675) <= a;
    layer5_outputs(676) <= b;
    layer5_outputs(677) <= b and not a;
    layer5_outputs(678) <= not (a or b);
    layer5_outputs(679) <= 1'b1;
    layer5_outputs(680) <= b;
    layer5_outputs(681) <= b and not a;
    layer5_outputs(682) <= not a;
    layer5_outputs(683) <= not b or a;
    layer5_outputs(684) <= not (a or b);
    layer5_outputs(685) <= not (a and b);
    layer5_outputs(686) <= not (a and b);
    layer5_outputs(687) <= not a;
    layer5_outputs(688) <= b and not a;
    layer5_outputs(689) <= not b;
    layer5_outputs(690) <= a;
    layer5_outputs(691) <= b;
    layer5_outputs(692) <= b and not a;
    layer5_outputs(693) <= not b;
    layer5_outputs(694) <= not (a xor b);
    layer5_outputs(695) <= a and not b;
    layer5_outputs(696) <= a;
    layer5_outputs(697) <= not b;
    layer5_outputs(698) <= a xor b;
    layer5_outputs(699) <= not a or b;
    layer5_outputs(700) <= b;
    layer5_outputs(701) <= a;
    layer5_outputs(702) <= not a or b;
    layer5_outputs(703) <= a and not b;
    layer5_outputs(704) <= not b;
    layer5_outputs(705) <= not (a or b);
    layer5_outputs(706) <= not b or a;
    layer5_outputs(707) <= b;
    layer5_outputs(708) <= 1'b0;
    layer5_outputs(709) <= a and b;
    layer5_outputs(710) <= b;
    layer5_outputs(711) <= not b or a;
    layer5_outputs(712) <= b and not a;
    layer5_outputs(713) <= not (a and b);
    layer5_outputs(714) <= 1'b1;
    layer5_outputs(715) <= not (a or b);
    layer5_outputs(716) <= b;
    layer5_outputs(717) <= a and not b;
    layer5_outputs(718) <= not (a and b);
    layer5_outputs(719) <= b and not a;
    layer5_outputs(720) <= not (a xor b);
    layer5_outputs(721) <= not a or b;
    layer5_outputs(722) <= 1'b1;
    layer5_outputs(723) <= b;
    layer5_outputs(724) <= a xor b;
    layer5_outputs(725) <= a;
    layer5_outputs(726) <= not a;
    layer5_outputs(727) <= b;
    layer5_outputs(728) <= b;
    layer5_outputs(729) <= not a or b;
    layer5_outputs(730) <= not a;
    layer5_outputs(731) <= a;
    layer5_outputs(732) <= not a or b;
    layer5_outputs(733) <= not a or b;
    layer5_outputs(734) <= not a or b;
    layer5_outputs(735) <= not a;
    layer5_outputs(736) <= b;
    layer5_outputs(737) <= a and not b;
    layer5_outputs(738) <= 1'b1;
    layer5_outputs(739) <= not b;
    layer5_outputs(740) <= 1'b1;
    layer5_outputs(741) <= not a or b;
    layer5_outputs(742) <= not (a and b);
    layer5_outputs(743) <= 1'b0;
    layer5_outputs(744) <= not (a or b);
    layer5_outputs(745) <= a and b;
    layer5_outputs(746) <= not (a and b);
    layer5_outputs(747) <= not (a xor b);
    layer5_outputs(748) <= b and not a;
    layer5_outputs(749) <= a or b;
    layer5_outputs(750) <= a and not b;
    layer5_outputs(751) <= not a or b;
    layer5_outputs(752) <= a and not b;
    layer5_outputs(753) <= a;
    layer5_outputs(754) <= not a;
    layer5_outputs(755) <= 1'b1;
    layer5_outputs(756) <= not b or a;
    layer5_outputs(757) <= a and b;
    layer5_outputs(758) <= b and not a;
    layer5_outputs(759) <= not a or b;
    layer5_outputs(760) <= 1'b1;
    layer5_outputs(761) <= not (a and b);
    layer5_outputs(762) <= a;
    layer5_outputs(763) <= a and not b;
    layer5_outputs(764) <= not a or b;
    layer5_outputs(765) <= not (a or b);
    layer5_outputs(766) <= b;
    layer5_outputs(767) <= b;
    layer5_outputs(768) <= not b;
    layer5_outputs(769) <= not b or a;
    layer5_outputs(770) <= 1'b1;
    layer5_outputs(771) <= not (a or b);
    layer5_outputs(772) <= not a;
    layer5_outputs(773) <= a;
    layer5_outputs(774) <= not a or b;
    layer5_outputs(775) <= a;
    layer5_outputs(776) <= b and not a;
    layer5_outputs(777) <= b;
    layer5_outputs(778) <= not b;
    layer5_outputs(779) <= not b or a;
    layer5_outputs(780) <= b;
    layer5_outputs(781) <= not a or b;
    layer5_outputs(782) <= b and not a;
    layer5_outputs(783) <= not a;
    layer5_outputs(784) <= 1'b1;
    layer5_outputs(785) <= a and not b;
    layer5_outputs(786) <= a or b;
    layer5_outputs(787) <= not b or a;
    layer5_outputs(788) <= not (a or b);
    layer5_outputs(789) <= a and b;
    layer5_outputs(790) <= not (a and b);
    layer5_outputs(791) <= a and b;
    layer5_outputs(792) <= not (a and b);
    layer5_outputs(793) <= 1'b1;
    layer5_outputs(794) <= a xor b;
    layer5_outputs(795) <= a and not b;
    layer5_outputs(796) <= a and not b;
    layer5_outputs(797) <= a;
    layer5_outputs(798) <= 1'b1;
    layer5_outputs(799) <= not (a and b);
    layer5_outputs(800) <= a and b;
    layer5_outputs(801) <= a and not b;
    layer5_outputs(802) <= a;
    layer5_outputs(803) <= not b;
    layer5_outputs(804) <= not (a or b);
    layer5_outputs(805) <= not b or a;
    layer5_outputs(806) <= not b;
    layer5_outputs(807) <= b and not a;
    layer5_outputs(808) <= not b;
    layer5_outputs(809) <= b;
    layer5_outputs(810) <= not (a or b);
    layer5_outputs(811) <= not a;
    layer5_outputs(812) <= not b or a;
    layer5_outputs(813) <= not a;
    layer5_outputs(814) <= not (a and b);
    layer5_outputs(815) <= 1'b0;
    layer5_outputs(816) <= 1'b0;
    layer5_outputs(817) <= b and not a;
    layer5_outputs(818) <= 1'b0;
    layer5_outputs(819) <= a;
    layer5_outputs(820) <= a;
    layer5_outputs(821) <= not (a and b);
    layer5_outputs(822) <= b and not a;
    layer5_outputs(823) <= not a;
    layer5_outputs(824) <= a;
    layer5_outputs(825) <= b;
    layer5_outputs(826) <= not b;
    layer5_outputs(827) <= b;
    layer5_outputs(828) <= not (a xor b);
    layer5_outputs(829) <= not a;
    layer5_outputs(830) <= not a or b;
    layer5_outputs(831) <= a or b;
    layer5_outputs(832) <= not b or a;
    layer5_outputs(833) <= a;
    layer5_outputs(834) <= b;
    layer5_outputs(835) <= not b;
    layer5_outputs(836) <= not a;
    layer5_outputs(837) <= not (a or b);
    layer5_outputs(838) <= b;
    layer5_outputs(839) <= a or b;
    layer5_outputs(840) <= not b;
    layer5_outputs(841) <= b;
    layer5_outputs(842) <= a;
    layer5_outputs(843) <= not b;
    layer5_outputs(844) <= not a or b;
    layer5_outputs(845) <= not b or a;
    layer5_outputs(846) <= not b;
    layer5_outputs(847) <= a xor b;
    layer5_outputs(848) <= not b;
    layer5_outputs(849) <= a and not b;
    layer5_outputs(850) <= a and not b;
    layer5_outputs(851) <= not b;
    layer5_outputs(852) <= a;
    layer5_outputs(853) <= a;
    layer5_outputs(854) <= not b or a;
    layer5_outputs(855) <= a xor b;
    layer5_outputs(856) <= not b;
    layer5_outputs(857) <= not b;
    layer5_outputs(858) <= not a;
    layer5_outputs(859) <= not (a or b);
    layer5_outputs(860) <= a and b;
    layer5_outputs(861) <= a or b;
    layer5_outputs(862) <= a;
    layer5_outputs(863) <= b;
    layer5_outputs(864) <= b and not a;
    layer5_outputs(865) <= a;
    layer5_outputs(866) <= not a;
    layer5_outputs(867) <= 1'b0;
    layer5_outputs(868) <= a and b;
    layer5_outputs(869) <= a and b;
    layer5_outputs(870) <= a;
    layer5_outputs(871) <= not a or b;
    layer5_outputs(872) <= a and b;
    layer5_outputs(873) <= b;
    layer5_outputs(874) <= 1'b0;
    layer5_outputs(875) <= not (a xor b);
    layer5_outputs(876) <= not (a and b);
    layer5_outputs(877) <= 1'b0;
    layer5_outputs(878) <= not (a xor b);
    layer5_outputs(879) <= not b;
    layer5_outputs(880) <= b;
    layer5_outputs(881) <= not a or b;
    layer5_outputs(882) <= not (a xor b);
    layer5_outputs(883) <= a and not b;
    layer5_outputs(884) <= not b or a;
    layer5_outputs(885) <= not b or a;
    layer5_outputs(886) <= not (a or b);
    layer5_outputs(887) <= not a or b;
    layer5_outputs(888) <= b;
    layer5_outputs(889) <= not (a or b);
    layer5_outputs(890) <= not (a xor b);
    layer5_outputs(891) <= b;
    layer5_outputs(892) <= 1'b0;
    layer5_outputs(893) <= not (a xor b);
    layer5_outputs(894) <= a or b;
    layer5_outputs(895) <= b and not a;
    layer5_outputs(896) <= 1'b0;
    layer5_outputs(897) <= a and not b;
    layer5_outputs(898) <= a xor b;
    layer5_outputs(899) <= a;
    layer5_outputs(900) <= not a;
    layer5_outputs(901) <= not b;
    layer5_outputs(902) <= 1'b1;
    layer5_outputs(903) <= not b;
    layer5_outputs(904) <= a;
    layer5_outputs(905) <= not a or b;
    layer5_outputs(906) <= not b or a;
    layer5_outputs(907) <= a and not b;
    layer5_outputs(908) <= not (a and b);
    layer5_outputs(909) <= not (a or b);
    layer5_outputs(910) <= not a;
    layer5_outputs(911) <= not b;
    layer5_outputs(912) <= a xor b;
    layer5_outputs(913) <= a;
    layer5_outputs(914) <= not (a and b);
    layer5_outputs(915) <= not a or b;
    layer5_outputs(916) <= not a or b;
    layer5_outputs(917) <= a or b;
    layer5_outputs(918) <= a and not b;
    layer5_outputs(919) <= a xor b;
    layer5_outputs(920) <= 1'b0;
    layer5_outputs(921) <= not (a and b);
    layer5_outputs(922) <= a and b;
    layer5_outputs(923) <= not a;
    layer5_outputs(924) <= not a;
    layer5_outputs(925) <= b;
    layer5_outputs(926) <= b;
    layer5_outputs(927) <= not a;
    layer5_outputs(928) <= 1'b1;
    layer5_outputs(929) <= 1'b1;
    layer5_outputs(930) <= a and b;
    layer5_outputs(931) <= a and not b;
    layer5_outputs(932) <= not (a xor b);
    layer5_outputs(933) <= a xor b;
    layer5_outputs(934) <= not b or a;
    layer5_outputs(935) <= b;
    layer5_outputs(936) <= a;
    layer5_outputs(937) <= a;
    layer5_outputs(938) <= not (a xor b);
    layer5_outputs(939) <= a;
    layer5_outputs(940) <= a;
    layer5_outputs(941) <= not a or b;
    layer5_outputs(942) <= a and b;
    layer5_outputs(943) <= not a or b;
    layer5_outputs(944) <= not (a or b);
    layer5_outputs(945) <= a and b;
    layer5_outputs(946) <= not b or a;
    layer5_outputs(947) <= not (a or b);
    layer5_outputs(948) <= b;
    layer5_outputs(949) <= not a;
    layer5_outputs(950) <= a;
    layer5_outputs(951) <= a and b;
    layer5_outputs(952) <= a or b;
    layer5_outputs(953) <= a or b;
    layer5_outputs(954) <= not (a or b);
    layer5_outputs(955) <= a and not b;
    layer5_outputs(956) <= b and not a;
    layer5_outputs(957) <= not a;
    layer5_outputs(958) <= not (a xor b);
    layer5_outputs(959) <= not a or b;
    layer5_outputs(960) <= 1'b0;
    layer5_outputs(961) <= not b or a;
    layer5_outputs(962) <= not b;
    layer5_outputs(963) <= 1'b0;
    layer5_outputs(964) <= not b;
    layer5_outputs(965) <= 1'b1;
    layer5_outputs(966) <= not a or b;
    layer5_outputs(967) <= b and not a;
    layer5_outputs(968) <= a and b;
    layer5_outputs(969) <= not b;
    layer5_outputs(970) <= b;
    layer5_outputs(971) <= not a;
    layer5_outputs(972) <= not a;
    layer5_outputs(973) <= a;
    layer5_outputs(974) <= not (a and b);
    layer5_outputs(975) <= not a;
    layer5_outputs(976) <= a or b;
    layer5_outputs(977) <= a;
    layer5_outputs(978) <= 1'b0;
    layer5_outputs(979) <= b and not a;
    layer5_outputs(980) <= not a or b;
    layer5_outputs(981) <= a and b;
    layer5_outputs(982) <= not a;
    layer5_outputs(983) <= not (a and b);
    layer5_outputs(984) <= not b or a;
    layer5_outputs(985) <= a;
    layer5_outputs(986) <= b and not a;
    layer5_outputs(987) <= not (a and b);
    layer5_outputs(988) <= not b;
    layer5_outputs(989) <= a and b;
    layer5_outputs(990) <= a;
    layer5_outputs(991) <= not a or b;
    layer5_outputs(992) <= not (a and b);
    layer5_outputs(993) <= not a or b;
    layer5_outputs(994) <= 1'b1;
    layer5_outputs(995) <= a and not b;
    layer5_outputs(996) <= a and b;
    layer5_outputs(997) <= a and not b;
    layer5_outputs(998) <= a;
    layer5_outputs(999) <= not a or b;
    layer5_outputs(1000) <= b and not a;
    layer5_outputs(1001) <= not b;
    layer5_outputs(1002) <= a and b;
    layer5_outputs(1003) <= not (a xor b);
    layer5_outputs(1004) <= not (a and b);
    layer5_outputs(1005) <= not b;
    layer5_outputs(1006) <= b;
    layer5_outputs(1007) <= a;
    layer5_outputs(1008) <= b and not a;
    layer5_outputs(1009) <= a and b;
    layer5_outputs(1010) <= a;
    layer5_outputs(1011) <= b and not a;
    layer5_outputs(1012) <= not (a and b);
    layer5_outputs(1013) <= b and not a;
    layer5_outputs(1014) <= not (a and b);
    layer5_outputs(1015) <= a or b;
    layer5_outputs(1016) <= not (a and b);
    layer5_outputs(1017) <= not a;
    layer5_outputs(1018) <= b and not a;
    layer5_outputs(1019) <= not a or b;
    layer5_outputs(1020) <= not a;
    layer5_outputs(1021) <= not (a and b);
    layer5_outputs(1022) <= a or b;
    layer5_outputs(1023) <= a and not b;
    layer5_outputs(1024) <= b;
    layer5_outputs(1025) <= b and not a;
    layer5_outputs(1026) <= not (a xor b);
    layer5_outputs(1027) <= not (a and b);
    layer5_outputs(1028) <= not b or a;
    layer5_outputs(1029) <= b and not a;
    layer5_outputs(1030) <= a;
    layer5_outputs(1031) <= not a or b;
    layer5_outputs(1032) <= a;
    layer5_outputs(1033) <= not (a or b);
    layer5_outputs(1034) <= a xor b;
    layer5_outputs(1035) <= 1'b1;
    layer5_outputs(1036) <= not a;
    layer5_outputs(1037) <= 1'b1;
    layer5_outputs(1038) <= a and b;
    layer5_outputs(1039) <= a;
    layer5_outputs(1040) <= a;
    layer5_outputs(1041) <= not a;
    layer5_outputs(1042) <= a and b;
    layer5_outputs(1043) <= not a or b;
    layer5_outputs(1044) <= not a;
    layer5_outputs(1045) <= not a;
    layer5_outputs(1046) <= not a;
    layer5_outputs(1047) <= a or b;
    layer5_outputs(1048) <= not (a and b);
    layer5_outputs(1049) <= a and not b;
    layer5_outputs(1050) <= 1'b1;
    layer5_outputs(1051) <= not (a or b);
    layer5_outputs(1052) <= not (a or b);
    layer5_outputs(1053) <= not b or a;
    layer5_outputs(1054) <= not (a and b);
    layer5_outputs(1055) <= b and not a;
    layer5_outputs(1056) <= a;
    layer5_outputs(1057) <= 1'b1;
    layer5_outputs(1058) <= a xor b;
    layer5_outputs(1059) <= not b;
    layer5_outputs(1060) <= not (a xor b);
    layer5_outputs(1061) <= not b;
    layer5_outputs(1062) <= not (a or b);
    layer5_outputs(1063) <= not b or a;
    layer5_outputs(1064) <= not b or a;
    layer5_outputs(1065) <= a;
    layer5_outputs(1066) <= a or b;
    layer5_outputs(1067) <= a;
    layer5_outputs(1068) <= 1'b0;
    layer5_outputs(1069) <= a and not b;
    layer5_outputs(1070) <= b;
    layer5_outputs(1071) <= not b;
    layer5_outputs(1072) <= 1'b0;
    layer5_outputs(1073) <= not a or b;
    layer5_outputs(1074) <= not b or a;
    layer5_outputs(1075) <= not a or b;
    layer5_outputs(1076) <= not a;
    layer5_outputs(1077) <= a and not b;
    layer5_outputs(1078) <= b and not a;
    layer5_outputs(1079) <= b and not a;
    layer5_outputs(1080) <= not a;
    layer5_outputs(1081) <= 1'b0;
    layer5_outputs(1082) <= not (a and b);
    layer5_outputs(1083) <= a and b;
    layer5_outputs(1084) <= b and not a;
    layer5_outputs(1085) <= not a or b;
    layer5_outputs(1086) <= not a;
    layer5_outputs(1087) <= not (a xor b);
    layer5_outputs(1088) <= 1'b1;
    layer5_outputs(1089) <= a;
    layer5_outputs(1090) <= b;
    layer5_outputs(1091) <= not b;
    layer5_outputs(1092) <= a or b;
    layer5_outputs(1093) <= not b;
    layer5_outputs(1094) <= 1'b1;
    layer5_outputs(1095) <= not (a and b);
    layer5_outputs(1096) <= not a or b;
    layer5_outputs(1097) <= a or b;
    layer5_outputs(1098) <= a or b;
    layer5_outputs(1099) <= a and not b;
    layer5_outputs(1100) <= b;
    layer5_outputs(1101) <= not (a or b);
    layer5_outputs(1102) <= not a;
    layer5_outputs(1103) <= not (a or b);
    layer5_outputs(1104) <= b;
    layer5_outputs(1105) <= a;
    layer5_outputs(1106) <= not b;
    layer5_outputs(1107) <= not (a or b);
    layer5_outputs(1108) <= a and b;
    layer5_outputs(1109) <= b and not a;
    layer5_outputs(1110) <= not b or a;
    layer5_outputs(1111) <= not (a or b);
    layer5_outputs(1112) <= not b or a;
    layer5_outputs(1113) <= b;
    layer5_outputs(1114) <= a and b;
    layer5_outputs(1115) <= not b;
    layer5_outputs(1116) <= not b or a;
    layer5_outputs(1117) <= not b or a;
    layer5_outputs(1118) <= b and not a;
    layer5_outputs(1119) <= not a;
    layer5_outputs(1120) <= not a;
    layer5_outputs(1121) <= b;
    layer5_outputs(1122) <= a or b;
    layer5_outputs(1123) <= not b;
    layer5_outputs(1124) <= b;
    layer5_outputs(1125) <= b and not a;
    layer5_outputs(1126) <= a;
    layer5_outputs(1127) <= a;
    layer5_outputs(1128) <= b;
    layer5_outputs(1129) <= not a;
    layer5_outputs(1130) <= not a;
    layer5_outputs(1131) <= not (a and b);
    layer5_outputs(1132) <= a and b;
    layer5_outputs(1133) <= not b or a;
    layer5_outputs(1134) <= a;
    layer5_outputs(1135) <= not (a and b);
    layer5_outputs(1136) <= not b or a;
    layer5_outputs(1137) <= not b or a;
    layer5_outputs(1138) <= not a;
    layer5_outputs(1139) <= not a;
    layer5_outputs(1140) <= a or b;
    layer5_outputs(1141) <= a and b;
    layer5_outputs(1142) <= not b;
    layer5_outputs(1143) <= 1'b0;
    layer5_outputs(1144) <= not b;
    layer5_outputs(1145) <= not (a xor b);
    layer5_outputs(1146) <= not a;
    layer5_outputs(1147) <= not (a or b);
    layer5_outputs(1148) <= not b;
    layer5_outputs(1149) <= not b;
    layer5_outputs(1150) <= not a;
    layer5_outputs(1151) <= b;
    layer5_outputs(1152) <= a and b;
    layer5_outputs(1153) <= not (a or b);
    layer5_outputs(1154) <= a;
    layer5_outputs(1155) <= a or b;
    layer5_outputs(1156) <= not (a or b);
    layer5_outputs(1157) <= 1'b1;
    layer5_outputs(1158) <= a;
    layer5_outputs(1159) <= b and not a;
    layer5_outputs(1160) <= not (a and b);
    layer5_outputs(1161) <= 1'b1;
    layer5_outputs(1162) <= a and not b;
    layer5_outputs(1163) <= not a or b;
    layer5_outputs(1164) <= a;
    layer5_outputs(1165) <= not a or b;
    layer5_outputs(1166) <= 1'b1;
    layer5_outputs(1167) <= a or b;
    layer5_outputs(1168) <= not (a xor b);
    layer5_outputs(1169) <= a;
    layer5_outputs(1170) <= a and not b;
    layer5_outputs(1171) <= b;
    layer5_outputs(1172) <= not (a and b);
    layer5_outputs(1173) <= not (a or b);
    layer5_outputs(1174) <= b and not a;
    layer5_outputs(1175) <= 1'b0;
    layer5_outputs(1176) <= not b;
    layer5_outputs(1177) <= b;
    layer5_outputs(1178) <= not b;
    layer5_outputs(1179) <= not (a or b);
    layer5_outputs(1180) <= a;
    layer5_outputs(1181) <= not a;
    layer5_outputs(1182) <= a and not b;
    layer5_outputs(1183) <= a and not b;
    layer5_outputs(1184) <= not a;
    layer5_outputs(1185) <= a;
    layer5_outputs(1186) <= a and not b;
    layer5_outputs(1187) <= a or b;
    layer5_outputs(1188) <= a;
    layer5_outputs(1189) <= a or b;
    layer5_outputs(1190) <= not b;
    layer5_outputs(1191) <= not b;
    layer5_outputs(1192) <= a or b;
    layer5_outputs(1193) <= 1'b0;
    layer5_outputs(1194) <= b;
    layer5_outputs(1195) <= b;
    layer5_outputs(1196) <= 1'b1;
    layer5_outputs(1197) <= 1'b0;
    layer5_outputs(1198) <= not (a and b);
    layer5_outputs(1199) <= not b;
    layer5_outputs(1200) <= b;
    layer5_outputs(1201) <= a;
    layer5_outputs(1202) <= a;
    layer5_outputs(1203) <= a;
    layer5_outputs(1204) <= not b;
    layer5_outputs(1205) <= not a;
    layer5_outputs(1206) <= a and b;
    layer5_outputs(1207) <= not (a and b);
    layer5_outputs(1208) <= a;
    layer5_outputs(1209) <= not b or a;
    layer5_outputs(1210) <= a or b;
    layer5_outputs(1211) <= a xor b;
    layer5_outputs(1212) <= a;
    layer5_outputs(1213) <= not (a and b);
    layer5_outputs(1214) <= b;
    layer5_outputs(1215) <= not b;
    layer5_outputs(1216) <= not a or b;
    layer5_outputs(1217) <= not b;
    layer5_outputs(1218) <= b;
    layer5_outputs(1219) <= not a;
    layer5_outputs(1220) <= a;
    layer5_outputs(1221) <= a;
    layer5_outputs(1222) <= not b;
    layer5_outputs(1223) <= a and b;
    layer5_outputs(1224) <= not a;
    layer5_outputs(1225) <= not b;
    layer5_outputs(1226) <= not (a or b);
    layer5_outputs(1227) <= a and not b;
    layer5_outputs(1228) <= not (a or b);
    layer5_outputs(1229) <= not a;
    layer5_outputs(1230) <= not a or b;
    layer5_outputs(1231) <= not (a and b);
    layer5_outputs(1232) <= a xor b;
    layer5_outputs(1233) <= not a;
    layer5_outputs(1234) <= not (a and b);
    layer5_outputs(1235) <= not a;
    layer5_outputs(1236) <= not b or a;
    layer5_outputs(1237) <= a and not b;
    layer5_outputs(1238) <= 1'b1;
    layer5_outputs(1239) <= a and not b;
    layer5_outputs(1240) <= not b;
    layer5_outputs(1241) <= not a or b;
    layer5_outputs(1242) <= not (a and b);
    layer5_outputs(1243) <= a and b;
    layer5_outputs(1244) <= not a;
    layer5_outputs(1245) <= b;
    layer5_outputs(1246) <= not b;
    layer5_outputs(1247) <= a and b;
    layer5_outputs(1248) <= 1'b0;
    layer5_outputs(1249) <= b;
    layer5_outputs(1250) <= b;
    layer5_outputs(1251) <= 1'b0;
    layer5_outputs(1252) <= b;
    layer5_outputs(1253) <= a;
    layer5_outputs(1254) <= not (a or b);
    layer5_outputs(1255) <= not (a or b);
    layer5_outputs(1256) <= not (a and b);
    layer5_outputs(1257) <= 1'b1;
    layer5_outputs(1258) <= a;
    layer5_outputs(1259) <= not (a or b);
    layer5_outputs(1260) <= a xor b;
    layer5_outputs(1261) <= b;
    layer5_outputs(1262) <= b;
    layer5_outputs(1263) <= a;
    layer5_outputs(1264) <= 1'b1;
    layer5_outputs(1265) <= not a or b;
    layer5_outputs(1266) <= a or b;
    layer5_outputs(1267) <= not a;
    layer5_outputs(1268) <= not (a and b);
    layer5_outputs(1269) <= not b;
    layer5_outputs(1270) <= not a;
    layer5_outputs(1271) <= a and not b;
    layer5_outputs(1272) <= not (a or b);
    layer5_outputs(1273) <= not a or b;
    layer5_outputs(1274) <= not a or b;
    layer5_outputs(1275) <= b;
    layer5_outputs(1276) <= not a;
    layer5_outputs(1277) <= a or b;
    layer5_outputs(1278) <= b and not a;
    layer5_outputs(1279) <= a and b;
    layer5_outputs(1280) <= not b;
    layer5_outputs(1281) <= b;
    layer5_outputs(1282) <= not (a xor b);
    layer5_outputs(1283) <= 1'b1;
    layer5_outputs(1284) <= not a;
    layer5_outputs(1285) <= b and not a;
    layer5_outputs(1286) <= a and b;
    layer5_outputs(1287) <= not a;
    layer5_outputs(1288) <= not a or b;
    layer5_outputs(1289) <= a and not b;
    layer5_outputs(1290) <= not (a xor b);
    layer5_outputs(1291) <= 1'b0;
    layer5_outputs(1292) <= not b or a;
    layer5_outputs(1293) <= a;
    layer5_outputs(1294) <= a or b;
    layer5_outputs(1295) <= a xor b;
    layer5_outputs(1296) <= not b or a;
    layer5_outputs(1297) <= not b;
    layer5_outputs(1298) <= not b or a;
    layer5_outputs(1299) <= b;
    layer5_outputs(1300) <= b and not a;
    layer5_outputs(1301) <= a and b;
    layer5_outputs(1302) <= a;
    layer5_outputs(1303) <= a or b;
    layer5_outputs(1304) <= not a;
    layer5_outputs(1305) <= b;
    layer5_outputs(1306) <= a and b;
    layer5_outputs(1307) <= not (a or b);
    layer5_outputs(1308) <= b and not a;
    layer5_outputs(1309) <= a and b;
    layer5_outputs(1310) <= not a or b;
    layer5_outputs(1311) <= not a or b;
    layer5_outputs(1312) <= a or b;
    layer5_outputs(1313) <= a;
    layer5_outputs(1314) <= a and not b;
    layer5_outputs(1315) <= not a or b;
    layer5_outputs(1316) <= a or b;
    layer5_outputs(1317) <= not (a and b);
    layer5_outputs(1318) <= not b or a;
    layer5_outputs(1319) <= a;
    layer5_outputs(1320) <= b;
    layer5_outputs(1321) <= not (a and b);
    layer5_outputs(1322) <= not a or b;
    layer5_outputs(1323) <= not b;
    layer5_outputs(1324) <= a or b;
    layer5_outputs(1325) <= b;
    layer5_outputs(1326) <= not b or a;
    layer5_outputs(1327) <= not (a xor b);
    layer5_outputs(1328) <= b and not a;
    layer5_outputs(1329) <= not b;
    layer5_outputs(1330) <= not b;
    layer5_outputs(1331) <= b and not a;
    layer5_outputs(1332) <= not b;
    layer5_outputs(1333) <= a;
    layer5_outputs(1334) <= not a;
    layer5_outputs(1335) <= b and not a;
    layer5_outputs(1336) <= not a or b;
    layer5_outputs(1337) <= not a;
    layer5_outputs(1338) <= not b or a;
    layer5_outputs(1339) <= a or b;
    layer5_outputs(1340) <= not a or b;
    layer5_outputs(1341) <= b;
    layer5_outputs(1342) <= a;
    layer5_outputs(1343) <= not a;
    layer5_outputs(1344) <= b;
    layer5_outputs(1345) <= not (a and b);
    layer5_outputs(1346) <= not b or a;
    layer5_outputs(1347) <= a;
    layer5_outputs(1348) <= not (a or b);
    layer5_outputs(1349) <= 1'b0;
    layer5_outputs(1350) <= b;
    layer5_outputs(1351) <= 1'b0;
    layer5_outputs(1352) <= a or b;
    layer5_outputs(1353) <= not a;
    layer5_outputs(1354) <= a and not b;
    layer5_outputs(1355) <= not b or a;
    layer5_outputs(1356) <= not b;
    layer5_outputs(1357) <= a;
    layer5_outputs(1358) <= not (a and b);
    layer5_outputs(1359) <= b;
    layer5_outputs(1360) <= 1'b0;
    layer5_outputs(1361) <= a;
    layer5_outputs(1362) <= 1'b1;
    layer5_outputs(1363) <= b and not a;
    layer5_outputs(1364) <= a and b;
    layer5_outputs(1365) <= a and not b;
    layer5_outputs(1366) <= not (a or b);
    layer5_outputs(1367) <= not (a xor b);
    layer5_outputs(1368) <= a and b;
    layer5_outputs(1369) <= not b;
    layer5_outputs(1370) <= not a;
    layer5_outputs(1371) <= not b;
    layer5_outputs(1372) <= a xor b;
    layer5_outputs(1373) <= not b;
    layer5_outputs(1374) <= a and not b;
    layer5_outputs(1375) <= a and not b;
    layer5_outputs(1376) <= b and not a;
    layer5_outputs(1377) <= not b or a;
    layer5_outputs(1378) <= a and not b;
    layer5_outputs(1379) <= b;
    layer5_outputs(1380) <= not (a or b);
    layer5_outputs(1381) <= not a or b;
    layer5_outputs(1382) <= b;
    layer5_outputs(1383) <= 1'b1;
    layer5_outputs(1384) <= b;
    layer5_outputs(1385) <= a and b;
    layer5_outputs(1386) <= a or b;
    layer5_outputs(1387) <= 1'b0;
    layer5_outputs(1388) <= b;
    layer5_outputs(1389) <= 1'b1;
    layer5_outputs(1390) <= a and not b;
    layer5_outputs(1391) <= not b or a;
    layer5_outputs(1392) <= not a;
    layer5_outputs(1393) <= b;
    layer5_outputs(1394) <= not b;
    layer5_outputs(1395) <= b and not a;
    layer5_outputs(1396) <= not b;
    layer5_outputs(1397) <= b and not a;
    layer5_outputs(1398) <= a;
    layer5_outputs(1399) <= a or b;
    layer5_outputs(1400) <= b;
    layer5_outputs(1401) <= a and b;
    layer5_outputs(1402) <= not (a or b);
    layer5_outputs(1403) <= a or b;
    layer5_outputs(1404) <= not (a xor b);
    layer5_outputs(1405) <= 1'b0;
    layer5_outputs(1406) <= not a;
    layer5_outputs(1407) <= not (a and b);
    layer5_outputs(1408) <= not b;
    layer5_outputs(1409) <= b;
    layer5_outputs(1410) <= a and b;
    layer5_outputs(1411) <= not (a or b);
    layer5_outputs(1412) <= 1'b0;
    layer5_outputs(1413) <= not b;
    layer5_outputs(1414) <= not (a or b);
    layer5_outputs(1415) <= b and not a;
    layer5_outputs(1416) <= not b or a;
    layer5_outputs(1417) <= a and b;
    layer5_outputs(1418) <= not a;
    layer5_outputs(1419) <= not (a or b);
    layer5_outputs(1420) <= a;
    layer5_outputs(1421) <= not b;
    layer5_outputs(1422) <= not b;
    layer5_outputs(1423) <= a and b;
    layer5_outputs(1424) <= a and b;
    layer5_outputs(1425) <= b;
    layer5_outputs(1426) <= not b or a;
    layer5_outputs(1427) <= not b or a;
    layer5_outputs(1428) <= b and not a;
    layer5_outputs(1429) <= not (a and b);
    layer5_outputs(1430) <= not b;
    layer5_outputs(1431) <= b and not a;
    layer5_outputs(1432) <= a;
    layer5_outputs(1433) <= b and not a;
    layer5_outputs(1434) <= not (a or b);
    layer5_outputs(1435) <= not b;
    layer5_outputs(1436) <= a and not b;
    layer5_outputs(1437) <= not b or a;
    layer5_outputs(1438) <= not b or a;
    layer5_outputs(1439) <= a and b;
    layer5_outputs(1440) <= a;
    layer5_outputs(1441) <= not (a and b);
    layer5_outputs(1442) <= a or b;
    layer5_outputs(1443) <= not (a or b);
    layer5_outputs(1444) <= a;
    layer5_outputs(1445) <= not a or b;
    layer5_outputs(1446) <= a or b;
    layer5_outputs(1447) <= 1'b0;
    layer5_outputs(1448) <= not a or b;
    layer5_outputs(1449) <= 1'b0;
    layer5_outputs(1450) <= not (a and b);
    layer5_outputs(1451) <= a and b;
    layer5_outputs(1452) <= a;
    layer5_outputs(1453) <= b;
    layer5_outputs(1454) <= a and not b;
    layer5_outputs(1455) <= not (a or b);
    layer5_outputs(1456) <= not b or a;
    layer5_outputs(1457) <= b;
    layer5_outputs(1458) <= a;
    layer5_outputs(1459) <= not b;
    layer5_outputs(1460) <= a;
    layer5_outputs(1461) <= not b or a;
    layer5_outputs(1462) <= a and not b;
    layer5_outputs(1463) <= not a;
    layer5_outputs(1464) <= 1'b1;
    layer5_outputs(1465) <= a or b;
    layer5_outputs(1466) <= b;
    layer5_outputs(1467) <= a and not b;
    layer5_outputs(1468) <= not (a and b);
    layer5_outputs(1469) <= a and not b;
    layer5_outputs(1470) <= not a;
    layer5_outputs(1471) <= b;
    layer5_outputs(1472) <= not a;
    layer5_outputs(1473) <= 1'b1;
    layer5_outputs(1474) <= a;
    layer5_outputs(1475) <= b and not a;
    layer5_outputs(1476) <= b and not a;
    layer5_outputs(1477) <= a xor b;
    layer5_outputs(1478) <= a xor b;
    layer5_outputs(1479) <= not b;
    layer5_outputs(1480) <= not (a or b);
    layer5_outputs(1481) <= 1'b1;
    layer5_outputs(1482) <= a xor b;
    layer5_outputs(1483) <= b and not a;
    layer5_outputs(1484) <= b and not a;
    layer5_outputs(1485) <= b;
    layer5_outputs(1486) <= b and not a;
    layer5_outputs(1487) <= a;
    layer5_outputs(1488) <= not (a and b);
    layer5_outputs(1489) <= b;
    layer5_outputs(1490) <= not a or b;
    layer5_outputs(1491) <= not a;
    layer5_outputs(1492) <= a and b;
    layer5_outputs(1493) <= not b or a;
    layer5_outputs(1494) <= a xor b;
    layer5_outputs(1495) <= 1'b1;
    layer5_outputs(1496) <= a or b;
    layer5_outputs(1497) <= a and not b;
    layer5_outputs(1498) <= not a or b;
    layer5_outputs(1499) <= a;
    layer5_outputs(1500) <= not b or a;
    layer5_outputs(1501) <= a;
    layer5_outputs(1502) <= not a;
    layer5_outputs(1503) <= a or b;
    layer5_outputs(1504) <= not b;
    layer5_outputs(1505) <= b and not a;
    layer5_outputs(1506) <= not a;
    layer5_outputs(1507) <= 1'b1;
    layer5_outputs(1508) <= b;
    layer5_outputs(1509) <= a and not b;
    layer5_outputs(1510) <= not a;
    layer5_outputs(1511) <= 1'b0;
    layer5_outputs(1512) <= not a;
    layer5_outputs(1513) <= b and not a;
    layer5_outputs(1514) <= a and b;
    layer5_outputs(1515) <= a;
    layer5_outputs(1516) <= a;
    layer5_outputs(1517) <= 1'b1;
    layer5_outputs(1518) <= a;
    layer5_outputs(1519) <= not a or b;
    layer5_outputs(1520) <= b and not a;
    layer5_outputs(1521) <= not a;
    layer5_outputs(1522) <= 1'b0;
    layer5_outputs(1523) <= not a or b;
    layer5_outputs(1524) <= not a or b;
    layer5_outputs(1525) <= not (a xor b);
    layer5_outputs(1526) <= not a;
    layer5_outputs(1527) <= a and b;
    layer5_outputs(1528) <= not b or a;
    layer5_outputs(1529) <= not (a and b);
    layer5_outputs(1530) <= not b or a;
    layer5_outputs(1531) <= b;
    layer5_outputs(1532) <= b and not a;
    layer5_outputs(1533) <= not (a xor b);
    layer5_outputs(1534) <= a or b;
    layer5_outputs(1535) <= not a;
    layer5_outputs(1536) <= not (a and b);
    layer5_outputs(1537) <= a;
    layer5_outputs(1538) <= a and b;
    layer5_outputs(1539) <= a and b;
    layer5_outputs(1540) <= a and b;
    layer5_outputs(1541) <= not (a and b);
    layer5_outputs(1542) <= b;
    layer5_outputs(1543) <= a and b;
    layer5_outputs(1544) <= not b;
    layer5_outputs(1545) <= not b;
    layer5_outputs(1546) <= a;
    layer5_outputs(1547) <= not b or a;
    layer5_outputs(1548) <= a and b;
    layer5_outputs(1549) <= a and b;
    layer5_outputs(1550) <= not b or a;
    layer5_outputs(1551) <= not (a or b);
    layer5_outputs(1552) <= not (a or b);
    layer5_outputs(1553) <= not (a and b);
    layer5_outputs(1554) <= b;
    layer5_outputs(1555) <= not (a or b);
    layer5_outputs(1556) <= not a or b;
    layer5_outputs(1557) <= b and not a;
    layer5_outputs(1558) <= not b;
    layer5_outputs(1559) <= not a or b;
    layer5_outputs(1560) <= a or b;
    layer5_outputs(1561) <= a and not b;
    layer5_outputs(1562) <= not b or a;
    layer5_outputs(1563) <= a and not b;
    layer5_outputs(1564) <= not a;
    layer5_outputs(1565) <= b and not a;
    layer5_outputs(1566) <= not a or b;
    layer5_outputs(1567) <= a and not b;
    layer5_outputs(1568) <= not a or b;
    layer5_outputs(1569) <= not (a or b);
    layer5_outputs(1570) <= not a;
    layer5_outputs(1571) <= b;
    layer5_outputs(1572) <= not b or a;
    layer5_outputs(1573) <= not b;
    layer5_outputs(1574) <= a or b;
    layer5_outputs(1575) <= not (a or b);
    layer5_outputs(1576) <= not (a or b);
    layer5_outputs(1577) <= not b or a;
    layer5_outputs(1578) <= a and not b;
    layer5_outputs(1579) <= not (a and b);
    layer5_outputs(1580) <= not (a and b);
    layer5_outputs(1581) <= a and b;
    layer5_outputs(1582) <= a xor b;
    layer5_outputs(1583) <= a and b;
    layer5_outputs(1584) <= a;
    layer5_outputs(1585) <= b;
    layer5_outputs(1586) <= not b;
    layer5_outputs(1587) <= not (a or b);
    layer5_outputs(1588) <= b and not a;
    layer5_outputs(1589) <= not b or a;
    layer5_outputs(1590) <= 1'b1;
    layer5_outputs(1591) <= a and b;
    layer5_outputs(1592) <= not b or a;
    layer5_outputs(1593) <= not a;
    layer5_outputs(1594) <= a;
    layer5_outputs(1595) <= b and not a;
    layer5_outputs(1596) <= 1'b0;
    layer5_outputs(1597) <= 1'b1;
    layer5_outputs(1598) <= b;
    layer5_outputs(1599) <= not a or b;
    layer5_outputs(1600) <= not (a and b);
    layer5_outputs(1601) <= not (a and b);
    layer5_outputs(1602) <= a;
    layer5_outputs(1603) <= not (a xor b);
    layer5_outputs(1604) <= 1'b0;
    layer5_outputs(1605) <= not a;
    layer5_outputs(1606) <= b;
    layer5_outputs(1607) <= not (a or b);
    layer5_outputs(1608) <= a and b;
    layer5_outputs(1609) <= not a;
    layer5_outputs(1610) <= not (a and b);
    layer5_outputs(1611) <= not (a xor b);
    layer5_outputs(1612) <= a and not b;
    layer5_outputs(1613) <= not a;
    layer5_outputs(1614) <= a and b;
    layer5_outputs(1615) <= not (a or b);
    layer5_outputs(1616) <= not a;
    layer5_outputs(1617) <= a;
    layer5_outputs(1618) <= not a or b;
    layer5_outputs(1619) <= b;
    layer5_outputs(1620) <= not a;
    layer5_outputs(1621) <= 1'b0;
    layer5_outputs(1622) <= 1'b0;
    layer5_outputs(1623) <= b and not a;
    layer5_outputs(1624) <= a and not b;
    layer5_outputs(1625) <= a xor b;
    layer5_outputs(1626) <= a or b;
    layer5_outputs(1627) <= not b;
    layer5_outputs(1628) <= a;
    layer5_outputs(1629) <= 1'b1;
    layer5_outputs(1630) <= b;
    layer5_outputs(1631) <= not a or b;
    layer5_outputs(1632) <= a and not b;
    layer5_outputs(1633) <= not b;
    layer5_outputs(1634) <= b;
    layer5_outputs(1635) <= b;
    layer5_outputs(1636) <= b and not a;
    layer5_outputs(1637) <= a and not b;
    layer5_outputs(1638) <= b;
    layer5_outputs(1639) <= not a;
    layer5_outputs(1640) <= b and not a;
    layer5_outputs(1641) <= not a;
    layer5_outputs(1642) <= not (a or b);
    layer5_outputs(1643) <= not a;
    layer5_outputs(1644) <= not (a or b);
    layer5_outputs(1645) <= a;
    layer5_outputs(1646) <= a;
    layer5_outputs(1647) <= not (a and b);
    layer5_outputs(1648) <= not a;
    layer5_outputs(1649) <= not (a and b);
    layer5_outputs(1650) <= a and not b;
    layer5_outputs(1651) <= not (a or b);
    layer5_outputs(1652) <= b and not a;
    layer5_outputs(1653) <= b;
    layer5_outputs(1654) <= b and not a;
    layer5_outputs(1655) <= a and not b;
    layer5_outputs(1656) <= 1'b0;
    layer5_outputs(1657) <= a and not b;
    layer5_outputs(1658) <= not a;
    layer5_outputs(1659) <= a and b;
    layer5_outputs(1660) <= not b or a;
    layer5_outputs(1661) <= a or b;
    layer5_outputs(1662) <= a;
    layer5_outputs(1663) <= not a;
    layer5_outputs(1664) <= not a;
    layer5_outputs(1665) <= not (a or b);
    layer5_outputs(1666) <= a;
    layer5_outputs(1667) <= not a;
    layer5_outputs(1668) <= not b or a;
    layer5_outputs(1669) <= not a or b;
    layer5_outputs(1670) <= a;
    layer5_outputs(1671) <= not (a or b);
    layer5_outputs(1672) <= 1'b1;
    layer5_outputs(1673) <= b;
    layer5_outputs(1674) <= 1'b0;
    layer5_outputs(1675) <= b;
    layer5_outputs(1676) <= b and not a;
    layer5_outputs(1677) <= not a or b;
    layer5_outputs(1678) <= not a;
    layer5_outputs(1679) <= a or b;
    layer5_outputs(1680) <= 1'b0;
    layer5_outputs(1681) <= 1'b1;
    layer5_outputs(1682) <= a;
    layer5_outputs(1683) <= a;
    layer5_outputs(1684) <= a and b;
    layer5_outputs(1685) <= b;
    layer5_outputs(1686) <= 1'b1;
    layer5_outputs(1687) <= not a or b;
    layer5_outputs(1688) <= not b;
    layer5_outputs(1689) <= not a;
    layer5_outputs(1690) <= a or b;
    layer5_outputs(1691) <= not (a or b);
    layer5_outputs(1692) <= a and b;
    layer5_outputs(1693) <= 1'b1;
    layer5_outputs(1694) <= not b;
    layer5_outputs(1695) <= not a;
    layer5_outputs(1696) <= b;
    layer5_outputs(1697) <= not a;
    layer5_outputs(1698) <= a or b;
    layer5_outputs(1699) <= not a or b;
    layer5_outputs(1700) <= not (a xor b);
    layer5_outputs(1701) <= not a or b;
    layer5_outputs(1702) <= a or b;
    layer5_outputs(1703) <= a and b;
    layer5_outputs(1704) <= a;
    layer5_outputs(1705) <= not b or a;
    layer5_outputs(1706) <= a and not b;
    layer5_outputs(1707) <= b;
    layer5_outputs(1708) <= a and b;
    layer5_outputs(1709) <= not b;
    layer5_outputs(1710) <= not a or b;
    layer5_outputs(1711) <= a xor b;
    layer5_outputs(1712) <= not b or a;
    layer5_outputs(1713) <= a;
    layer5_outputs(1714) <= not b or a;
    layer5_outputs(1715) <= not a;
    layer5_outputs(1716) <= not a;
    layer5_outputs(1717) <= not a;
    layer5_outputs(1718) <= not (a or b);
    layer5_outputs(1719) <= not (a and b);
    layer5_outputs(1720) <= a and not b;
    layer5_outputs(1721) <= not a;
    layer5_outputs(1722) <= a or b;
    layer5_outputs(1723) <= not a;
    layer5_outputs(1724) <= a or b;
    layer5_outputs(1725) <= b and not a;
    layer5_outputs(1726) <= a;
    layer5_outputs(1727) <= not (a or b);
    layer5_outputs(1728) <= a and b;
    layer5_outputs(1729) <= not b;
    layer5_outputs(1730) <= a xor b;
    layer5_outputs(1731) <= b;
    layer5_outputs(1732) <= not b;
    layer5_outputs(1733) <= not a;
    layer5_outputs(1734) <= not a;
    layer5_outputs(1735) <= a;
    layer5_outputs(1736) <= 1'b1;
    layer5_outputs(1737) <= not (a or b);
    layer5_outputs(1738) <= not b;
    layer5_outputs(1739) <= a and not b;
    layer5_outputs(1740) <= not a or b;
    layer5_outputs(1741) <= a;
    layer5_outputs(1742) <= 1'b0;
    layer5_outputs(1743) <= not b;
    layer5_outputs(1744) <= not a;
    layer5_outputs(1745) <= a and not b;
    layer5_outputs(1746) <= a;
    layer5_outputs(1747) <= not a or b;
    layer5_outputs(1748) <= not a;
    layer5_outputs(1749) <= not b;
    layer5_outputs(1750) <= 1'b1;
    layer5_outputs(1751) <= not (a xor b);
    layer5_outputs(1752) <= a and not b;
    layer5_outputs(1753) <= not (a or b);
    layer5_outputs(1754) <= not (a and b);
    layer5_outputs(1755) <= not b or a;
    layer5_outputs(1756) <= not b or a;
    layer5_outputs(1757) <= not b;
    layer5_outputs(1758) <= a;
    layer5_outputs(1759) <= a and not b;
    layer5_outputs(1760) <= 1'b1;
    layer5_outputs(1761) <= b and not a;
    layer5_outputs(1762) <= a or b;
    layer5_outputs(1763) <= not (a and b);
    layer5_outputs(1764) <= not (a and b);
    layer5_outputs(1765) <= not b;
    layer5_outputs(1766) <= 1'b1;
    layer5_outputs(1767) <= not a;
    layer5_outputs(1768) <= not a;
    layer5_outputs(1769) <= not a or b;
    layer5_outputs(1770) <= not a;
    layer5_outputs(1771) <= not (a or b);
    layer5_outputs(1772) <= not a;
    layer5_outputs(1773) <= not a or b;
    layer5_outputs(1774) <= a xor b;
    layer5_outputs(1775) <= a and b;
    layer5_outputs(1776) <= a and b;
    layer5_outputs(1777) <= b;
    layer5_outputs(1778) <= not (a or b);
    layer5_outputs(1779) <= b and not a;
    layer5_outputs(1780) <= not a or b;
    layer5_outputs(1781) <= not (a or b);
    layer5_outputs(1782) <= not a or b;
    layer5_outputs(1783) <= not (a and b);
    layer5_outputs(1784) <= not a or b;
    layer5_outputs(1785) <= 1'b1;
    layer5_outputs(1786) <= not (a or b);
    layer5_outputs(1787) <= not b;
    layer5_outputs(1788) <= not (a or b);
    layer5_outputs(1789) <= b;
    layer5_outputs(1790) <= b;
    layer5_outputs(1791) <= b;
    layer5_outputs(1792) <= not (a and b);
    layer5_outputs(1793) <= not b or a;
    layer5_outputs(1794) <= not (a and b);
    layer5_outputs(1795) <= not a or b;
    layer5_outputs(1796) <= not (a and b);
    layer5_outputs(1797) <= 1'b0;
    layer5_outputs(1798) <= not (a and b);
    layer5_outputs(1799) <= not a;
    layer5_outputs(1800) <= a and b;
    layer5_outputs(1801) <= 1'b0;
    layer5_outputs(1802) <= not (a and b);
    layer5_outputs(1803) <= not b or a;
    layer5_outputs(1804) <= a xor b;
    layer5_outputs(1805) <= b and not a;
    layer5_outputs(1806) <= a;
    layer5_outputs(1807) <= not (a and b);
    layer5_outputs(1808) <= a xor b;
    layer5_outputs(1809) <= not (a and b);
    layer5_outputs(1810) <= not a;
    layer5_outputs(1811) <= not a;
    layer5_outputs(1812) <= not b;
    layer5_outputs(1813) <= not a;
    layer5_outputs(1814) <= not a;
    layer5_outputs(1815) <= not b or a;
    layer5_outputs(1816) <= not b;
    layer5_outputs(1817) <= b;
    layer5_outputs(1818) <= not b;
    layer5_outputs(1819) <= not b or a;
    layer5_outputs(1820) <= b and not a;
    layer5_outputs(1821) <= a;
    layer5_outputs(1822) <= not (a xor b);
    layer5_outputs(1823) <= not (a and b);
    layer5_outputs(1824) <= a;
    layer5_outputs(1825) <= a or b;
    layer5_outputs(1826) <= a and not b;
    layer5_outputs(1827) <= a and b;
    layer5_outputs(1828) <= 1'b0;
    layer5_outputs(1829) <= not b;
    layer5_outputs(1830) <= b;
    layer5_outputs(1831) <= not a or b;
    layer5_outputs(1832) <= not (a or b);
    layer5_outputs(1833) <= not (a or b);
    layer5_outputs(1834) <= a and b;
    layer5_outputs(1835) <= not (a and b);
    layer5_outputs(1836) <= a and b;
    layer5_outputs(1837) <= not a;
    layer5_outputs(1838) <= b;
    layer5_outputs(1839) <= not a;
    layer5_outputs(1840) <= not b;
    layer5_outputs(1841) <= not (a and b);
    layer5_outputs(1842) <= a or b;
    layer5_outputs(1843) <= a;
    layer5_outputs(1844) <= not b;
    layer5_outputs(1845) <= not (a or b);
    layer5_outputs(1846) <= b;
    layer5_outputs(1847) <= not b;
    layer5_outputs(1848) <= not a or b;
    layer5_outputs(1849) <= not a;
    layer5_outputs(1850) <= a xor b;
    layer5_outputs(1851) <= a xor b;
    layer5_outputs(1852) <= a;
    layer5_outputs(1853) <= b;
    layer5_outputs(1854) <= not b;
    layer5_outputs(1855) <= a or b;
    layer5_outputs(1856) <= not (a xor b);
    layer5_outputs(1857) <= not b or a;
    layer5_outputs(1858) <= a and b;
    layer5_outputs(1859) <= a xor b;
    layer5_outputs(1860) <= a and not b;
    layer5_outputs(1861) <= not a or b;
    layer5_outputs(1862) <= a and not b;
    layer5_outputs(1863) <= a;
    layer5_outputs(1864) <= b;
    layer5_outputs(1865) <= a or b;
    layer5_outputs(1866) <= a and not b;
    layer5_outputs(1867) <= b;
    layer5_outputs(1868) <= not (a or b);
    layer5_outputs(1869) <= a and b;
    layer5_outputs(1870) <= a or b;
    layer5_outputs(1871) <= not b or a;
    layer5_outputs(1872) <= a;
    layer5_outputs(1873) <= not a;
    layer5_outputs(1874) <= a and not b;
    layer5_outputs(1875) <= not b;
    layer5_outputs(1876) <= b and not a;
    layer5_outputs(1877) <= not b;
    layer5_outputs(1878) <= not a or b;
    layer5_outputs(1879) <= a and b;
    layer5_outputs(1880) <= a and not b;
    layer5_outputs(1881) <= a and not b;
    layer5_outputs(1882) <= not a or b;
    layer5_outputs(1883) <= not b;
    layer5_outputs(1884) <= b;
    layer5_outputs(1885) <= not b or a;
    layer5_outputs(1886) <= not b;
    layer5_outputs(1887) <= not a;
    layer5_outputs(1888) <= b;
    layer5_outputs(1889) <= b and not a;
    layer5_outputs(1890) <= not b;
    layer5_outputs(1891) <= not (a or b);
    layer5_outputs(1892) <= not a;
    layer5_outputs(1893) <= 1'b0;
    layer5_outputs(1894) <= b and not a;
    layer5_outputs(1895) <= a xor b;
    layer5_outputs(1896) <= a and not b;
    layer5_outputs(1897) <= 1'b1;
    layer5_outputs(1898) <= not a or b;
    layer5_outputs(1899) <= not (a xor b);
    layer5_outputs(1900) <= b and not a;
    layer5_outputs(1901) <= a and b;
    layer5_outputs(1902) <= b;
    layer5_outputs(1903) <= a or b;
    layer5_outputs(1904) <= not (a and b);
    layer5_outputs(1905) <= not b or a;
    layer5_outputs(1906) <= a and not b;
    layer5_outputs(1907) <= a or b;
    layer5_outputs(1908) <= not a;
    layer5_outputs(1909) <= not a or b;
    layer5_outputs(1910) <= not (a or b);
    layer5_outputs(1911) <= a and not b;
    layer5_outputs(1912) <= 1'b0;
    layer5_outputs(1913) <= 1'b0;
    layer5_outputs(1914) <= b;
    layer5_outputs(1915) <= a and not b;
    layer5_outputs(1916) <= a;
    layer5_outputs(1917) <= a;
    layer5_outputs(1918) <= a and b;
    layer5_outputs(1919) <= a and not b;
    layer5_outputs(1920) <= a and b;
    layer5_outputs(1921) <= a;
    layer5_outputs(1922) <= b;
    layer5_outputs(1923) <= not (a or b);
    layer5_outputs(1924) <= b and not a;
    layer5_outputs(1925) <= 1'b1;
    layer5_outputs(1926) <= a and not b;
    layer5_outputs(1927) <= a;
    layer5_outputs(1928) <= 1'b0;
    layer5_outputs(1929) <= b and not a;
    layer5_outputs(1930) <= b and not a;
    layer5_outputs(1931) <= a or b;
    layer5_outputs(1932) <= 1'b1;
    layer5_outputs(1933) <= not (a and b);
    layer5_outputs(1934) <= not (a and b);
    layer5_outputs(1935) <= a and not b;
    layer5_outputs(1936) <= not a;
    layer5_outputs(1937) <= not b;
    layer5_outputs(1938) <= not b or a;
    layer5_outputs(1939) <= not a;
    layer5_outputs(1940) <= a;
    layer5_outputs(1941) <= not (a and b);
    layer5_outputs(1942) <= a or b;
    layer5_outputs(1943) <= not a;
    layer5_outputs(1944) <= 1'b0;
    layer5_outputs(1945) <= not b or a;
    layer5_outputs(1946) <= b;
    layer5_outputs(1947) <= a;
    layer5_outputs(1948) <= a;
    layer5_outputs(1949) <= not b;
    layer5_outputs(1950) <= b and not a;
    layer5_outputs(1951) <= a and not b;
    layer5_outputs(1952) <= not (a and b);
    layer5_outputs(1953) <= a or b;
    layer5_outputs(1954) <= not (a xor b);
    layer5_outputs(1955) <= not (a and b);
    layer5_outputs(1956) <= not (a or b);
    layer5_outputs(1957) <= not a or b;
    layer5_outputs(1958) <= a or b;
    layer5_outputs(1959) <= not b or a;
    layer5_outputs(1960) <= b;
    layer5_outputs(1961) <= b and not a;
    layer5_outputs(1962) <= not a;
    layer5_outputs(1963) <= b;
    layer5_outputs(1964) <= b;
    layer5_outputs(1965) <= b;
    layer5_outputs(1966) <= not (a or b);
    layer5_outputs(1967) <= 1'b1;
    layer5_outputs(1968) <= a;
    layer5_outputs(1969) <= a or b;
    layer5_outputs(1970) <= a or b;
    layer5_outputs(1971) <= a and b;
    layer5_outputs(1972) <= not b;
    layer5_outputs(1973) <= a or b;
    layer5_outputs(1974) <= a and not b;
    layer5_outputs(1975) <= not (a and b);
    layer5_outputs(1976) <= a and not b;
    layer5_outputs(1977) <= a and b;
    layer5_outputs(1978) <= not a;
    layer5_outputs(1979) <= not (a or b);
    layer5_outputs(1980) <= not (a xor b);
    layer5_outputs(1981) <= not a;
    layer5_outputs(1982) <= a and not b;
    layer5_outputs(1983) <= b;
    layer5_outputs(1984) <= not b;
    layer5_outputs(1985) <= b and not a;
    layer5_outputs(1986) <= a and b;
    layer5_outputs(1987) <= a and not b;
    layer5_outputs(1988) <= not (a xor b);
    layer5_outputs(1989) <= a;
    layer5_outputs(1990) <= 1'b1;
    layer5_outputs(1991) <= not a;
    layer5_outputs(1992) <= a;
    layer5_outputs(1993) <= a or b;
    layer5_outputs(1994) <= b and not a;
    layer5_outputs(1995) <= not (a and b);
    layer5_outputs(1996) <= not a or b;
    layer5_outputs(1997) <= 1'b0;
    layer5_outputs(1998) <= not a or b;
    layer5_outputs(1999) <= b and not a;
    layer5_outputs(2000) <= not a;
    layer5_outputs(2001) <= b;
    layer5_outputs(2002) <= a and b;
    layer5_outputs(2003) <= not (a or b);
    layer5_outputs(2004) <= not b or a;
    layer5_outputs(2005) <= not (a or b);
    layer5_outputs(2006) <= not b or a;
    layer5_outputs(2007) <= b and not a;
    layer5_outputs(2008) <= a;
    layer5_outputs(2009) <= a and not b;
    layer5_outputs(2010) <= a and b;
    layer5_outputs(2011) <= not b or a;
    layer5_outputs(2012) <= not a;
    layer5_outputs(2013) <= 1'b1;
    layer5_outputs(2014) <= not (a and b);
    layer5_outputs(2015) <= b;
    layer5_outputs(2016) <= b;
    layer5_outputs(2017) <= not a;
    layer5_outputs(2018) <= b;
    layer5_outputs(2019) <= a or b;
    layer5_outputs(2020) <= not a;
    layer5_outputs(2021) <= not a or b;
    layer5_outputs(2022) <= 1'b0;
    layer5_outputs(2023) <= a and b;
    layer5_outputs(2024) <= not b;
    layer5_outputs(2025) <= a or b;
    layer5_outputs(2026) <= b;
    layer5_outputs(2027) <= a xor b;
    layer5_outputs(2028) <= a;
    layer5_outputs(2029) <= a and not b;
    layer5_outputs(2030) <= not a;
    layer5_outputs(2031) <= b;
    layer5_outputs(2032) <= a and b;
    layer5_outputs(2033) <= b;
    layer5_outputs(2034) <= a and not b;
    layer5_outputs(2035) <= a and b;
    layer5_outputs(2036) <= a or b;
    layer5_outputs(2037) <= b and not a;
    layer5_outputs(2038) <= 1'b0;
    layer5_outputs(2039) <= a and not b;
    layer5_outputs(2040) <= not a;
    layer5_outputs(2041) <= not a;
    layer5_outputs(2042) <= a and b;
    layer5_outputs(2043) <= not (a and b);
    layer5_outputs(2044) <= 1'b1;
    layer5_outputs(2045) <= not (a and b);
    layer5_outputs(2046) <= b and not a;
    layer5_outputs(2047) <= not (a and b);
    layer5_outputs(2048) <= not b or a;
    layer5_outputs(2049) <= not b;
    layer5_outputs(2050) <= not (a and b);
    layer5_outputs(2051) <= 1'b0;
    layer5_outputs(2052) <= not a;
    layer5_outputs(2053) <= not (a and b);
    layer5_outputs(2054) <= not b or a;
    layer5_outputs(2055) <= b;
    layer5_outputs(2056) <= a and b;
    layer5_outputs(2057) <= not b;
    layer5_outputs(2058) <= not a;
    layer5_outputs(2059) <= a and not b;
    layer5_outputs(2060) <= not (a and b);
    layer5_outputs(2061) <= not a;
    layer5_outputs(2062) <= 1'b1;
    layer5_outputs(2063) <= b and not a;
    layer5_outputs(2064) <= not (a xor b);
    layer5_outputs(2065) <= not (a or b);
    layer5_outputs(2066) <= b;
    layer5_outputs(2067) <= b;
    layer5_outputs(2068) <= b and not a;
    layer5_outputs(2069) <= a or b;
    layer5_outputs(2070) <= not (a or b);
    layer5_outputs(2071) <= b;
    layer5_outputs(2072) <= not b or a;
    layer5_outputs(2073) <= a and b;
    layer5_outputs(2074) <= b and not a;
    layer5_outputs(2075) <= 1'b0;
    layer5_outputs(2076) <= not (a and b);
    layer5_outputs(2077) <= b and not a;
    layer5_outputs(2078) <= not a;
    layer5_outputs(2079) <= not b or a;
    layer5_outputs(2080) <= not b;
    layer5_outputs(2081) <= not b;
    layer5_outputs(2082) <= not b;
    layer5_outputs(2083) <= a;
    layer5_outputs(2084) <= not b;
    layer5_outputs(2085) <= not a;
    layer5_outputs(2086) <= a;
    layer5_outputs(2087) <= not a or b;
    layer5_outputs(2088) <= a and not b;
    layer5_outputs(2089) <= not a;
    layer5_outputs(2090) <= 1'b0;
    layer5_outputs(2091) <= not b;
    layer5_outputs(2092) <= not b;
    layer5_outputs(2093) <= not b;
    layer5_outputs(2094) <= not (a and b);
    layer5_outputs(2095) <= not a or b;
    layer5_outputs(2096) <= 1'b1;
    layer5_outputs(2097) <= a and b;
    layer5_outputs(2098) <= a and not b;
    layer5_outputs(2099) <= not b or a;
    layer5_outputs(2100) <= a and not b;
    layer5_outputs(2101) <= not a;
    layer5_outputs(2102) <= not (a and b);
    layer5_outputs(2103) <= not a;
    layer5_outputs(2104) <= 1'b1;
    layer5_outputs(2105) <= a and not b;
    layer5_outputs(2106) <= a and not b;
    layer5_outputs(2107) <= not b or a;
    layer5_outputs(2108) <= not (a xor b);
    layer5_outputs(2109) <= a;
    layer5_outputs(2110) <= not b or a;
    layer5_outputs(2111) <= not (a or b);
    layer5_outputs(2112) <= not b or a;
    layer5_outputs(2113) <= b and not a;
    layer5_outputs(2114) <= a and b;
    layer5_outputs(2115) <= not (a or b);
    layer5_outputs(2116) <= not b;
    layer5_outputs(2117) <= 1'b0;
    layer5_outputs(2118) <= a;
    layer5_outputs(2119) <= b;
    layer5_outputs(2120) <= not b or a;
    layer5_outputs(2121) <= a and b;
    layer5_outputs(2122) <= b and not a;
    layer5_outputs(2123) <= not (a or b);
    layer5_outputs(2124) <= not (a and b);
    layer5_outputs(2125) <= not b;
    layer5_outputs(2126) <= b;
    layer5_outputs(2127) <= not (a xor b);
    layer5_outputs(2128) <= b and not a;
    layer5_outputs(2129) <= not (a and b);
    layer5_outputs(2130) <= not a;
    layer5_outputs(2131) <= a and b;
    layer5_outputs(2132) <= not a or b;
    layer5_outputs(2133) <= a;
    layer5_outputs(2134) <= not (a and b);
    layer5_outputs(2135) <= a;
    layer5_outputs(2136) <= a;
    layer5_outputs(2137) <= not b;
    layer5_outputs(2138) <= 1'b1;
    layer5_outputs(2139) <= not a or b;
    layer5_outputs(2140) <= a and b;
    layer5_outputs(2141) <= not a;
    layer5_outputs(2142) <= b;
    layer5_outputs(2143) <= not (a and b);
    layer5_outputs(2144) <= a and not b;
    layer5_outputs(2145) <= 1'b1;
    layer5_outputs(2146) <= not (a xor b);
    layer5_outputs(2147) <= 1'b1;
    layer5_outputs(2148) <= 1'b0;
    layer5_outputs(2149) <= a xor b;
    layer5_outputs(2150) <= a or b;
    layer5_outputs(2151) <= b;
    layer5_outputs(2152) <= a xor b;
    layer5_outputs(2153) <= not b;
    layer5_outputs(2154) <= b;
    layer5_outputs(2155) <= not a or b;
    layer5_outputs(2156) <= not a or b;
    layer5_outputs(2157) <= not a;
    layer5_outputs(2158) <= not b or a;
    layer5_outputs(2159) <= a xor b;
    layer5_outputs(2160) <= not (a or b);
    layer5_outputs(2161) <= b;
    layer5_outputs(2162) <= not a;
    layer5_outputs(2163) <= not a or b;
    layer5_outputs(2164) <= a;
    layer5_outputs(2165) <= b;
    layer5_outputs(2166) <= not b;
    layer5_outputs(2167) <= a;
    layer5_outputs(2168) <= a;
    layer5_outputs(2169) <= 1'b1;
    layer5_outputs(2170) <= a or b;
    layer5_outputs(2171) <= not (a xor b);
    layer5_outputs(2172) <= b;
    layer5_outputs(2173) <= a and not b;
    layer5_outputs(2174) <= not b or a;
    layer5_outputs(2175) <= b;
    layer5_outputs(2176) <= not b or a;
    layer5_outputs(2177) <= not b;
    layer5_outputs(2178) <= not a;
    layer5_outputs(2179) <= b;
    layer5_outputs(2180) <= b;
    layer5_outputs(2181) <= 1'b0;
    layer5_outputs(2182) <= not (a and b);
    layer5_outputs(2183) <= not b or a;
    layer5_outputs(2184) <= not a;
    layer5_outputs(2185) <= not b or a;
    layer5_outputs(2186) <= a xor b;
    layer5_outputs(2187) <= not a;
    layer5_outputs(2188) <= not a;
    layer5_outputs(2189) <= b and not a;
    layer5_outputs(2190) <= a and not b;
    layer5_outputs(2191) <= b;
    layer5_outputs(2192) <= not (a and b);
    layer5_outputs(2193) <= a;
    layer5_outputs(2194) <= not b;
    layer5_outputs(2195) <= b and not a;
    layer5_outputs(2196) <= not b;
    layer5_outputs(2197) <= b;
    layer5_outputs(2198) <= not a;
    layer5_outputs(2199) <= b and not a;
    layer5_outputs(2200) <= not (a and b);
    layer5_outputs(2201) <= 1'b1;
    layer5_outputs(2202) <= 1'b1;
    layer5_outputs(2203) <= not a;
    layer5_outputs(2204) <= not a or b;
    layer5_outputs(2205) <= not (a or b);
    layer5_outputs(2206) <= a and b;
    layer5_outputs(2207) <= not (a or b);
    layer5_outputs(2208) <= a;
    layer5_outputs(2209) <= 1'b0;
    layer5_outputs(2210) <= not (a or b);
    layer5_outputs(2211) <= a xor b;
    layer5_outputs(2212) <= not b;
    layer5_outputs(2213) <= a or b;
    layer5_outputs(2214) <= a and b;
    layer5_outputs(2215) <= 1'b0;
    layer5_outputs(2216) <= not b or a;
    layer5_outputs(2217) <= not (a and b);
    layer5_outputs(2218) <= not (a and b);
    layer5_outputs(2219) <= b and not a;
    layer5_outputs(2220) <= b;
    layer5_outputs(2221) <= a and not b;
    layer5_outputs(2222) <= not a or b;
    layer5_outputs(2223) <= 1'b0;
    layer5_outputs(2224) <= a or b;
    layer5_outputs(2225) <= 1'b1;
    layer5_outputs(2226) <= a and b;
    layer5_outputs(2227) <= not a or b;
    layer5_outputs(2228) <= 1'b0;
    layer5_outputs(2229) <= not b;
    layer5_outputs(2230) <= a or b;
    layer5_outputs(2231) <= not a;
    layer5_outputs(2232) <= not b;
    layer5_outputs(2233) <= not (a and b);
    layer5_outputs(2234) <= a xor b;
    layer5_outputs(2235) <= not a or b;
    layer5_outputs(2236) <= 1'b1;
    layer5_outputs(2237) <= b;
    layer5_outputs(2238) <= not (a or b);
    layer5_outputs(2239) <= b;
    layer5_outputs(2240) <= not (a or b);
    layer5_outputs(2241) <= not a or b;
    layer5_outputs(2242) <= b and not a;
    layer5_outputs(2243) <= b;
    layer5_outputs(2244) <= b;
    layer5_outputs(2245) <= not b;
    layer5_outputs(2246) <= 1'b1;
    layer5_outputs(2247) <= not b or a;
    layer5_outputs(2248) <= a and not b;
    layer5_outputs(2249) <= a and b;
    layer5_outputs(2250) <= a;
    layer5_outputs(2251) <= a;
    layer5_outputs(2252) <= a and b;
    layer5_outputs(2253) <= b and not a;
    layer5_outputs(2254) <= a and not b;
    layer5_outputs(2255) <= a and not b;
    layer5_outputs(2256) <= a;
    layer5_outputs(2257) <= a or b;
    layer5_outputs(2258) <= not a or b;
    layer5_outputs(2259) <= not a;
    layer5_outputs(2260) <= b and not a;
    layer5_outputs(2261) <= not (a and b);
    layer5_outputs(2262) <= not b;
    layer5_outputs(2263) <= a and not b;
    layer5_outputs(2264) <= not a;
    layer5_outputs(2265) <= not (a xor b);
    layer5_outputs(2266) <= a and b;
    layer5_outputs(2267) <= a;
    layer5_outputs(2268) <= a and not b;
    layer5_outputs(2269) <= a xor b;
    layer5_outputs(2270) <= b;
    layer5_outputs(2271) <= b and not a;
    layer5_outputs(2272) <= a;
    layer5_outputs(2273) <= 1'b1;
    layer5_outputs(2274) <= a xor b;
    layer5_outputs(2275) <= a and not b;
    layer5_outputs(2276) <= not (a or b);
    layer5_outputs(2277) <= a and not b;
    layer5_outputs(2278) <= not b;
    layer5_outputs(2279) <= a;
    layer5_outputs(2280) <= a or b;
    layer5_outputs(2281) <= b and not a;
    layer5_outputs(2282) <= a and not b;
    layer5_outputs(2283) <= a and not b;
    layer5_outputs(2284) <= b;
    layer5_outputs(2285) <= b and not a;
    layer5_outputs(2286) <= not b;
    layer5_outputs(2287) <= not (a and b);
    layer5_outputs(2288) <= not (a and b);
    layer5_outputs(2289) <= not b or a;
    layer5_outputs(2290) <= a and b;
    layer5_outputs(2291) <= not (a or b);
    layer5_outputs(2292) <= b and not a;
    layer5_outputs(2293) <= b;
    layer5_outputs(2294) <= b and not a;
    layer5_outputs(2295) <= not a or b;
    layer5_outputs(2296) <= a or b;
    layer5_outputs(2297) <= b;
    layer5_outputs(2298) <= 1'b0;
    layer5_outputs(2299) <= not a;
    layer5_outputs(2300) <= b;
    layer5_outputs(2301) <= b and not a;
    layer5_outputs(2302) <= not a;
    layer5_outputs(2303) <= b;
    layer5_outputs(2304) <= a and not b;
    layer5_outputs(2305) <= a or b;
    layer5_outputs(2306) <= b and not a;
    layer5_outputs(2307) <= not a or b;
    layer5_outputs(2308) <= not a;
    layer5_outputs(2309) <= b and not a;
    layer5_outputs(2310) <= not a;
    layer5_outputs(2311) <= a or b;
    layer5_outputs(2312) <= a;
    layer5_outputs(2313) <= not a or b;
    layer5_outputs(2314) <= not a or b;
    layer5_outputs(2315) <= not b;
    layer5_outputs(2316) <= not a or b;
    layer5_outputs(2317) <= not (a or b);
    layer5_outputs(2318) <= 1'b0;
    layer5_outputs(2319) <= not (a and b);
    layer5_outputs(2320) <= not a;
    layer5_outputs(2321) <= a and b;
    layer5_outputs(2322) <= not (a and b);
    layer5_outputs(2323) <= not (a or b);
    layer5_outputs(2324) <= a and b;
    layer5_outputs(2325) <= b;
    layer5_outputs(2326) <= not (a or b);
    layer5_outputs(2327) <= a;
    layer5_outputs(2328) <= not (a and b);
    layer5_outputs(2329) <= not (a or b);
    layer5_outputs(2330) <= a and b;
    layer5_outputs(2331) <= a;
    layer5_outputs(2332) <= a and not b;
    layer5_outputs(2333) <= a and not b;
    layer5_outputs(2334) <= not a;
    layer5_outputs(2335) <= b and not a;
    layer5_outputs(2336) <= a;
    layer5_outputs(2337) <= a xor b;
    layer5_outputs(2338) <= not b;
    layer5_outputs(2339) <= not (a or b);
    layer5_outputs(2340) <= a and not b;
    layer5_outputs(2341) <= not a or b;
    layer5_outputs(2342) <= a;
    layer5_outputs(2343) <= b and not a;
    layer5_outputs(2344) <= a;
    layer5_outputs(2345) <= not a;
    layer5_outputs(2346) <= b and not a;
    layer5_outputs(2347) <= not b;
    layer5_outputs(2348) <= not a or b;
    layer5_outputs(2349) <= a and not b;
    layer5_outputs(2350) <= a and not b;
    layer5_outputs(2351) <= 1'b0;
    layer5_outputs(2352) <= 1'b0;
    layer5_outputs(2353) <= a xor b;
    layer5_outputs(2354) <= not (a or b);
    layer5_outputs(2355) <= not (a and b);
    layer5_outputs(2356) <= b and not a;
    layer5_outputs(2357) <= a;
    layer5_outputs(2358) <= b and not a;
    layer5_outputs(2359) <= not (a and b);
    layer5_outputs(2360) <= not b;
    layer5_outputs(2361) <= not (a or b);
    layer5_outputs(2362) <= b;
    layer5_outputs(2363) <= not a;
    layer5_outputs(2364) <= b and not a;
    layer5_outputs(2365) <= not b or a;
    layer5_outputs(2366) <= a;
    layer5_outputs(2367) <= a;
    layer5_outputs(2368) <= b;
    layer5_outputs(2369) <= not (a or b);
    layer5_outputs(2370) <= not a or b;
    layer5_outputs(2371) <= b and not a;
    layer5_outputs(2372) <= not b;
    layer5_outputs(2373) <= not (a and b);
    layer5_outputs(2374) <= a and not b;
    layer5_outputs(2375) <= not a or b;
    layer5_outputs(2376) <= a;
    layer5_outputs(2377) <= a and not b;
    layer5_outputs(2378) <= not a;
    layer5_outputs(2379) <= not b;
    layer5_outputs(2380) <= not b or a;
    layer5_outputs(2381) <= a and b;
    layer5_outputs(2382) <= a or b;
    layer5_outputs(2383) <= a;
    layer5_outputs(2384) <= 1'b0;
    layer5_outputs(2385) <= a or b;
    layer5_outputs(2386) <= not b;
    layer5_outputs(2387) <= not a or b;
    layer5_outputs(2388) <= not a;
    layer5_outputs(2389) <= a and b;
    layer5_outputs(2390) <= b;
    layer5_outputs(2391) <= b;
    layer5_outputs(2392) <= not (a and b);
    layer5_outputs(2393) <= not a or b;
    layer5_outputs(2394) <= not (a and b);
    layer5_outputs(2395) <= not b or a;
    layer5_outputs(2396) <= a or b;
    layer5_outputs(2397) <= b;
    layer5_outputs(2398) <= a;
    layer5_outputs(2399) <= b and not a;
    layer5_outputs(2400) <= not (a or b);
    layer5_outputs(2401) <= not a or b;
    layer5_outputs(2402) <= not a or b;
    layer5_outputs(2403) <= b and not a;
    layer5_outputs(2404) <= not (a and b);
    layer5_outputs(2405) <= not (a and b);
    layer5_outputs(2406) <= not (a and b);
    layer5_outputs(2407) <= a and not b;
    layer5_outputs(2408) <= not a;
    layer5_outputs(2409) <= a and b;
    layer5_outputs(2410) <= a and b;
    layer5_outputs(2411) <= 1'b1;
    layer5_outputs(2412) <= not (a and b);
    layer5_outputs(2413) <= not b or a;
    layer5_outputs(2414) <= 1'b1;
    layer5_outputs(2415) <= a and b;
    layer5_outputs(2416) <= b;
    layer5_outputs(2417) <= 1'b1;
    layer5_outputs(2418) <= not b;
    layer5_outputs(2419) <= a and not b;
    layer5_outputs(2420) <= not (a or b);
    layer5_outputs(2421) <= not (a and b);
    layer5_outputs(2422) <= not b or a;
    layer5_outputs(2423) <= 1'b0;
    layer5_outputs(2424) <= a and not b;
    layer5_outputs(2425) <= 1'b1;
    layer5_outputs(2426) <= b and not a;
    layer5_outputs(2427) <= b and not a;
    layer5_outputs(2428) <= a;
    layer5_outputs(2429) <= a and not b;
    layer5_outputs(2430) <= not b;
    layer5_outputs(2431) <= not a or b;
    layer5_outputs(2432) <= a;
    layer5_outputs(2433) <= not a;
    layer5_outputs(2434) <= a and b;
    layer5_outputs(2435) <= not a or b;
    layer5_outputs(2436) <= b;
    layer5_outputs(2437) <= not b;
    layer5_outputs(2438) <= a or b;
    layer5_outputs(2439) <= a;
    layer5_outputs(2440) <= not b or a;
    layer5_outputs(2441) <= not b;
    layer5_outputs(2442) <= b;
    layer5_outputs(2443) <= not (a or b);
    layer5_outputs(2444) <= 1'b1;
    layer5_outputs(2445) <= not b;
    layer5_outputs(2446) <= not b or a;
    layer5_outputs(2447) <= not (a xor b);
    layer5_outputs(2448) <= not b or a;
    layer5_outputs(2449) <= b and not a;
    layer5_outputs(2450) <= not (a and b);
    layer5_outputs(2451) <= b;
    layer5_outputs(2452) <= b and not a;
    layer5_outputs(2453) <= not a;
    layer5_outputs(2454) <= not b or a;
    layer5_outputs(2455) <= a and b;
    layer5_outputs(2456) <= a;
    layer5_outputs(2457) <= not b;
    layer5_outputs(2458) <= b;
    layer5_outputs(2459) <= not a;
    layer5_outputs(2460) <= a and b;
    layer5_outputs(2461) <= not (a or b);
    layer5_outputs(2462) <= a and b;
    layer5_outputs(2463) <= not b or a;
    layer5_outputs(2464) <= not a;
    layer5_outputs(2465) <= not a;
    layer5_outputs(2466) <= not b or a;
    layer5_outputs(2467) <= not b or a;
    layer5_outputs(2468) <= b;
    layer5_outputs(2469) <= b and not a;
    layer5_outputs(2470) <= a;
    layer5_outputs(2471) <= not (a or b);
    layer5_outputs(2472) <= 1'b0;
    layer5_outputs(2473) <= not (a or b);
    layer5_outputs(2474) <= not a or b;
    layer5_outputs(2475) <= not b or a;
    layer5_outputs(2476) <= not b or a;
    layer5_outputs(2477) <= not (a and b);
    layer5_outputs(2478) <= 1'b0;
    layer5_outputs(2479) <= 1'b1;
    layer5_outputs(2480) <= 1'b0;
    layer5_outputs(2481) <= not a or b;
    layer5_outputs(2482) <= a or b;
    layer5_outputs(2483) <= b;
    layer5_outputs(2484) <= a and b;
    layer5_outputs(2485) <= not a or b;
    layer5_outputs(2486) <= a and b;
    layer5_outputs(2487) <= b and not a;
    layer5_outputs(2488) <= a;
    layer5_outputs(2489) <= not a;
    layer5_outputs(2490) <= a xor b;
    layer5_outputs(2491) <= a;
    layer5_outputs(2492) <= a and b;
    layer5_outputs(2493) <= not b;
    layer5_outputs(2494) <= a and not b;
    layer5_outputs(2495) <= 1'b1;
    layer5_outputs(2496) <= a and b;
    layer5_outputs(2497) <= a and b;
    layer5_outputs(2498) <= b;
    layer5_outputs(2499) <= 1'b0;
    layer5_outputs(2500) <= not b or a;
    layer5_outputs(2501) <= not (a or b);
    layer5_outputs(2502) <= not b;
    layer5_outputs(2503) <= not a;
    layer5_outputs(2504) <= a;
    layer5_outputs(2505) <= b;
    layer5_outputs(2506) <= a and not b;
    layer5_outputs(2507) <= not (a and b);
    layer5_outputs(2508) <= a and b;
    layer5_outputs(2509) <= a;
    layer5_outputs(2510) <= 1'b1;
    layer5_outputs(2511) <= b and not a;
    layer5_outputs(2512) <= not b;
    layer5_outputs(2513) <= a or b;
    layer5_outputs(2514) <= not b;
    layer5_outputs(2515) <= b and not a;
    layer5_outputs(2516) <= not b;
    layer5_outputs(2517) <= not a or b;
    layer5_outputs(2518) <= b;
    layer5_outputs(2519) <= a;
    layer5_outputs(2520) <= a or b;
    layer5_outputs(2521) <= a or b;
    layer5_outputs(2522) <= not (a and b);
    layer5_outputs(2523) <= 1'b0;
    layer5_outputs(2524) <= b and not a;
    layer5_outputs(2525) <= not a;
    layer5_outputs(2526) <= b and not a;
    layer5_outputs(2527) <= a;
    layer5_outputs(2528) <= not b;
    layer5_outputs(2529) <= not b;
    layer5_outputs(2530) <= a and b;
    layer5_outputs(2531) <= not (a and b);
    layer5_outputs(2532) <= b and not a;
    layer5_outputs(2533) <= a and not b;
    layer5_outputs(2534) <= not b;
    layer5_outputs(2535) <= b;
    layer5_outputs(2536) <= not (a and b);
    layer5_outputs(2537) <= b and not a;
    layer5_outputs(2538) <= a or b;
    layer5_outputs(2539) <= not b;
    layer5_outputs(2540) <= not a;
    layer5_outputs(2541) <= a or b;
    layer5_outputs(2542) <= 1'b0;
    layer5_outputs(2543) <= not b;
    layer5_outputs(2544) <= not b or a;
    layer5_outputs(2545) <= not b;
    layer5_outputs(2546) <= not (a and b);
    layer5_outputs(2547) <= not b;
    layer5_outputs(2548) <= b and not a;
    layer5_outputs(2549) <= a;
    layer5_outputs(2550) <= not (a xor b);
    layer5_outputs(2551) <= a or b;
    layer5_outputs(2552) <= not (a and b);
    layer5_outputs(2553) <= not b;
    layer5_outputs(2554) <= a and b;
    layer5_outputs(2555) <= not a;
    layer5_outputs(2556) <= a and b;
    layer5_outputs(2557) <= b;
    layer5_outputs(2558) <= not (a or b);
    layer5_outputs(2559) <= not a or b;
    layer6_outputs(0) <= a and b;
    layer6_outputs(1) <= not (a or b);
    layer6_outputs(2) <= not (a and b);
    layer6_outputs(3) <= 1'b1;
    layer6_outputs(4) <= b;
    layer6_outputs(5) <= a and b;
    layer6_outputs(6) <= not a or b;
    layer6_outputs(7) <= not (a or b);
    layer6_outputs(8) <= not a;
    layer6_outputs(9) <= a and b;
    layer6_outputs(10) <= not a or b;
    layer6_outputs(11) <= a and b;
    layer6_outputs(12) <= a xor b;
    layer6_outputs(13) <= a and b;
    layer6_outputs(14) <= a;
    layer6_outputs(15) <= b and not a;
    layer6_outputs(16) <= not (a xor b);
    layer6_outputs(17) <= b;
    layer6_outputs(18) <= not (a and b);
    layer6_outputs(19) <= not b;
    layer6_outputs(20) <= a or b;
    layer6_outputs(21) <= a and not b;
    layer6_outputs(22) <= a and not b;
    layer6_outputs(23) <= a xor b;
    layer6_outputs(24) <= not (a and b);
    layer6_outputs(25) <= not a;
    layer6_outputs(26) <= not a;
    layer6_outputs(27) <= not a;
    layer6_outputs(28) <= not a;
    layer6_outputs(29) <= not b or a;
    layer6_outputs(30) <= a;
    layer6_outputs(31) <= a;
    layer6_outputs(32) <= b;
    layer6_outputs(33) <= a and b;
    layer6_outputs(34) <= not b;
    layer6_outputs(35) <= not (a and b);
    layer6_outputs(36) <= a and b;
    layer6_outputs(37) <= a and b;
    layer6_outputs(38) <= a;
    layer6_outputs(39) <= a or b;
    layer6_outputs(40) <= a and not b;
    layer6_outputs(41) <= not a or b;
    layer6_outputs(42) <= not (a and b);
    layer6_outputs(43) <= not (a or b);
    layer6_outputs(44) <= a or b;
    layer6_outputs(45) <= a;
    layer6_outputs(46) <= a;
    layer6_outputs(47) <= not (a xor b);
    layer6_outputs(48) <= a or b;
    layer6_outputs(49) <= b;
    layer6_outputs(50) <= b and not a;
    layer6_outputs(51) <= not (a xor b);
    layer6_outputs(52) <= b;
    layer6_outputs(53) <= 1'b1;
    layer6_outputs(54) <= a;
    layer6_outputs(55) <= b;
    layer6_outputs(56) <= a;
    layer6_outputs(57) <= b;
    layer6_outputs(58) <= a;
    layer6_outputs(59) <= not b;
    layer6_outputs(60) <= a or b;
    layer6_outputs(61) <= b and not a;
    layer6_outputs(62) <= not b or a;
    layer6_outputs(63) <= not (a and b);
    layer6_outputs(64) <= a and not b;
    layer6_outputs(65) <= not a or b;
    layer6_outputs(66) <= not a;
    layer6_outputs(67) <= a and b;
    layer6_outputs(68) <= a;
    layer6_outputs(69) <= not a;
    layer6_outputs(70) <= not (a or b);
    layer6_outputs(71) <= not a;
    layer6_outputs(72) <= a or b;
    layer6_outputs(73) <= not b;
    layer6_outputs(74) <= a and not b;
    layer6_outputs(75) <= a;
    layer6_outputs(76) <= not a or b;
    layer6_outputs(77) <= a or b;
    layer6_outputs(78) <= a or b;
    layer6_outputs(79) <= a and not b;
    layer6_outputs(80) <= not b or a;
    layer6_outputs(81) <= b;
    layer6_outputs(82) <= b;
    layer6_outputs(83) <= b;
    layer6_outputs(84) <= not b;
    layer6_outputs(85) <= b and not a;
    layer6_outputs(86) <= 1'b1;
    layer6_outputs(87) <= a;
    layer6_outputs(88) <= not b or a;
    layer6_outputs(89) <= not a or b;
    layer6_outputs(90) <= a xor b;
    layer6_outputs(91) <= b;
    layer6_outputs(92) <= a and b;
    layer6_outputs(93) <= b;
    layer6_outputs(94) <= not (a and b);
    layer6_outputs(95) <= not b or a;
    layer6_outputs(96) <= not a;
    layer6_outputs(97) <= not (a or b);
    layer6_outputs(98) <= not b or a;
    layer6_outputs(99) <= a and b;
    layer6_outputs(100) <= not (a xor b);
    layer6_outputs(101) <= a;
    layer6_outputs(102) <= not b;
    layer6_outputs(103) <= b and not a;
    layer6_outputs(104) <= not (a and b);
    layer6_outputs(105) <= b;
    layer6_outputs(106) <= not a;
    layer6_outputs(107) <= a and not b;
    layer6_outputs(108) <= b and not a;
    layer6_outputs(109) <= not a or b;
    layer6_outputs(110) <= a;
    layer6_outputs(111) <= not a;
    layer6_outputs(112) <= not a;
    layer6_outputs(113) <= b;
    layer6_outputs(114) <= not b;
    layer6_outputs(115) <= not a or b;
    layer6_outputs(116) <= not (a or b);
    layer6_outputs(117) <= a and b;
    layer6_outputs(118) <= a;
    layer6_outputs(119) <= not a;
    layer6_outputs(120) <= not (a xor b);
    layer6_outputs(121) <= b and not a;
    layer6_outputs(122) <= not (a xor b);
    layer6_outputs(123) <= not a or b;
    layer6_outputs(124) <= not a or b;
    layer6_outputs(125) <= a or b;
    layer6_outputs(126) <= not (a and b);
    layer6_outputs(127) <= a;
    layer6_outputs(128) <= not a;
    layer6_outputs(129) <= a;
    layer6_outputs(130) <= not a;
    layer6_outputs(131) <= not a;
    layer6_outputs(132) <= not (a or b);
    layer6_outputs(133) <= not b or a;
    layer6_outputs(134) <= not b;
    layer6_outputs(135) <= b and not a;
    layer6_outputs(136) <= not (a or b);
    layer6_outputs(137) <= b and not a;
    layer6_outputs(138) <= not (a and b);
    layer6_outputs(139) <= not b;
    layer6_outputs(140) <= 1'b0;
    layer6_outputs(141) <= not a or b;
    layer6_outputs(142) <= not (a and b);
    layer6_outputs(143) <= a and not b;
    layer6_outputs(144) <= not (a and b);
    layer6_outputs(145) <= b and not a;
    layer6_outputs(146) <= not a;
    layer6_outputs(147) <= a and b;
    layer6_outputs(148) <= b;
    layer6_outputs(149) <= not (a or b);
    layer6_outputs(150) <= a and b;
    layer6_outputs(151) <= not b;
    layer6_outputs(152) <= not (a or b);
    layer6_outputs(153) <= a;
    layer6_outputs(154) <= not a;
    layer6_outputs(155) <= a and b;
    layer6_outputs(156) <= a and not b;
    layer6_outputs(157) <= not b;
    layer6_outputs(158) <= b;
    layer6_outputs(159) <= b and not a;
    layer6_outputs(160) <= a;
    layer6_outputs(161) <= a;
    layer6_outputs(162) <= 1'b1;
    layer6_outputs(163) <= a and b;
    layer6_outputs(164) <= a;
    layer6_outputs(165) <= a xor b;
    layer6_outputs(166) <= not (a or b);
    layer6_outputs(167) <= a and not b;
    layer6_outputs(168) <= b;
    layer6_outputs(169) <= a and b;
    layer6_outputs(170) <= not b;
    layer6_outputs(171) <= not b or a;
    layer6_outputs(172) <= not a;
    layer6_outputs(173) <= a and b;
    layer6_outputs(174) <= b;
    layer6_outputs(175) <= not a;
    layer6_outputs(176) <= 1'b1;
    layer6_outputs(177) <= b;
    layer6_outputs(178) <= 1'b0;
    layer6_outputs(179) <= not b or a;
    layer6_outputs(180) <= a;
    layer6_outputs(181) <= not a or b;
    layer6_outputs(182) <= not a;
    layer6_outputs(183) <= b and not a;
    layer6_outputs(184) <= not (a or b);
    layer6_outputs(185) <= a;
    layer6_outputs(186) <= a and b;
    layer6_outputs(187) <= a xor b;
    layer6_outputs(188) <= b and not a;
    layer6_outputs(189) <= b;
    layer6_outputs(190) <= not (a or b);
    layer6_outputs(191) <= not (a or b);
    layer6_outputs(192) <= not (a and b);
    layer6_outputs(193) <= b;
    layer6_outputs(194) <= not (a xor b);
    layer6_outputs(195) <= not (a and b);
    layer6_outputs(196) <= a and not b;
    layer6_outputs(197) <= a;
    layer6_outputs(198) <= not b or a;
    layer6_outputs(199) <= a and b;
    layer6_outputs(200) <= not (a and b);
    layer6_outputs(201) <= not b;
    layer6_outputs(202) <= b and not a;
    layer6_outputs(203) <= b;
    layer6_outputs(204) <= a and not b;
    layer6_outputs(205) <= not b;
    layer6_outputs(206) <= not (a xor b);
    layer6_outputs(207) <= a xor b;
    layer6_outputs(208) <= a or b;
    layer6_outputs(209) <= a;
    layer6_outputs(210) <= not (a xor b);
    layer6_outputs(211) <= b;
    layer6_outputs(212) <= not a;
    layer6_outputs(213) <= a;
    layer6_outputs(214) <= not (a xor b);
    layer6_outputs(215) <= a and not b;
    layer6_outputs(216) <= a and b;
    layer6_outputs(217) <= a;
    layer6_outputs(218) <= a;
    layer6_outputs(219) <= a;
    layer6_outputs(220) <= b;
    layer6_outputs(221) <= b;
    layer6_outputs(222) <= not b;
    layer6_outputs(223) <= b;
    layer6_outputs(224) <= a and not b;
    layer6_outputs(225) <= b and not a;
    layer6_outputs(226) <= not (a and b);
    layer6_outputs(227) <= a and b;
    layer6_outputs(228) <= not b;
    layer6_outputs(229) <= a or b;
    layer6_outputs(230) <= a or b;
    layer6_outputs(231) <= a and b;
    layer6_outputs(232) <= a or b;
    layer6_outputs(233) <= a and not b;
    layer6_outputs(234) <= not (a and b);
    layer6_outputs(235) <= not (a or b);
    layer6_outputs(236) <= not b or a;
    layer6_outputs(237) <= not (a or b);
    layer6_outputs(238) <= not (a xor b);
    layer6_outputs(239) <= b and not a;
    layer6_outputs(240) <= b and not a;
    layer6_outputs(241) <= not a or b;
    layer6_outputs(242) <= not (a or b);
    layer6_outputs(243) <= not a;
    layer6_outputs(244) <= not a or b;
    layer6_outputs(245) <= not (a and b);
    layer6_outputs(246) <= a;
    layer6_outputs(247) <= a and b;
    layer6_outputs(248) <= a and b;
    layer6_outputs(249) <= b and not a;
    layer6_outputs(250) <= b and not a;
    layer6_outputs(251) <= a and not b;
    layer6_outputs(252) <= b;
    layer6_outputs(253) <= not b or a;
    layer6_outputs(254) <= 1'b0;
    layer6_outputs(255) <= a or b;
    layer6_outputs(256) <= not b or a;
    layer6_outputs(257) <= 1'b1;
    layer6_outputs(258) <= a;
    layer6_outputs(259) <= 1'b1;
    layer6_outputs(260) <= not a;
    layer6_outputs(261) <= not b;
    layer6_outputs(262) <= not b;
    layer6_outputs(263) <= not a;
    layer6_outputs(264) <= not (a xor b);
    layer6_outputs(265) <= not (a and b);
    layer6_outputs(266) <= not a;
    layer6_outputs(267) <= not a;
    layer6_outputs(268) <= a;
    layer6_outputs(269) <= not b or a;
    layer6_outputs(270) <= 1'b0;
    layer6_outputs(271) <= b and not a;
    layer6_outputs(272) <= not (a and b);
    layer6_outputs(273) <= not b;
    layer6_outputs(274) <= not (a or b);
    layer6_outputs(275) <= not a or b;
    layer6_outputs(276) <= b and not a;
    layer6_outputs(277) <= not a or b;
    layer6_outputs(278) <= a and b;
    layer6_outputs(279) <= b;
    layer6_outputs(280) <= not a or b;
    layer6_outputs(281) <= a and not b;
    layer6_outputs(282) <= 1'b1;
    layer6_outputs(283) <= a and not b;
    layer6_outputs(284) <= not (a or b);
    layer6_outputs(285) <= a;
    layer6_outputs(286) <= not a or b;
    layer6_outputs(287) <= not b;
    layer6_outputs(288) <= 1'b0;
    layer6_outputs(289) <= a and not b;
    layer6_outputs(290) <= b;
    layer6_outputs(291) <= a and not b;
    layer6_outputs(292) <= not (a or b);
    layer6_outputs(293) <= a;
    layer6_outputs(294) <= a and b;
    layer6_outputs(295) <= not (a or b);
    layer6_outputs(296) <= not (a and b);
    layer6_outputs(297) <= a xor b;
    layer6_outputs(298) <= b;
    layer6_outputs(299) <= not (a xor b);
    layer6_outputs(300) <= not a or b;
    layer6_outputs(301) <= not b;
    layer6_outputs(302) <= a;
    layer6_outputs(303) <= not a or b;
    layer6_outputs(304) <= not (a or b);
    layer6_outputs(305) <= not (a or b);
    layer6_outputs(306) <= b;
    layer6_outputs(307) <= not a;
    layer6_outputs(308) <= not b or a;
    layer6_outputs(309) <= b;
    layer6_outputs(310) <= a and b;
    layer6_outputs(311) <= not (a or b);
    layer6_outputs(312) <= not b;
    layer6_outputs(313) <= not b or a;
    layer6_outputs(314) <= not b or a;
    layer6_outputs(315) <= a or b;
    layer6_outputs(316) <= b;
    layer6_outputs(317) <= not b;
    layer6_outputs(318) <= a and not b;
    layer6_outputs(319) <= a and b;
    layer6_outputs(320) <= a;
    layer6_outputs(321) <= a and not b;
    layer6_outputs(322) <= a and not b;
    layer6_outputs(323) <= not b or a;
    layer6_outputs(324) <= b and not a;
    layer6_outputs(325) <= a;
    layer6_outputs(326) <= b;
    layer6_outputs(327) <= not b;
    layer6_outputs(328) <= not a;
    layer6_outputs(329) <= not b or a;
    layer6_outputs(330) <= not b;
    layer6_outputs(331) <= b;
    layer6_outputs(332) <= 1'b1;
    layer6_outputs(333) <= a;
    layer6_outputs(334) <= a xor b;
    layer6_outputs(335) <= b and not a;
    layer6_outputs(336) <= a;
    layer6_outputs(337) <= a xor b;
    layer6_outputs(338) <= a or b;
    layer6_outputs(339) <= a and b;
    layer6_outputs(340) <= not b;
    layer6_outputs(341) <= a and b;
    layer6_outputs(342) <= not b;
    layer6_outputs(343) <= a or b;
    layer6_outputs(344) <= not b or a;
    layer6_outputs(345) <= b and not a;
    layer6_outputs(346) <= not (a or b);
    layer6_outputs(347) <= a;
    layer6_outputs(348) <= a xor b;
    layer6_outputs(349) <= a;
    layer6_outputs(350) <= a and not b;
    layer6_outputs(351) <= b;
    layer6_outputs(352) <= a and b;
    layer6_outputs(353) <= not a;
    layer6_outputs(354) <= a;
    layer6_outputs(355) <= a;
    layer6_outputs(356) <= a;
    layer6_outputs(357) <= not b;
    layer6_outputs(358) <= a or b;
    layer6_outputs(359) <= not (a or b);
    layer6_outputs(360) <= a or b;
    layer6_outputs(361) <= not a;
    layer6_outputs(362) <= not a;
    layer6_outputs(363) <= b;
    layer6_outputs(364) <= not b or a;
    layer6_outputs(365) <= not (a or b);
    layer6_outputs(366) <= a or b;
    layer6_outputs(367) <= not b;
    layer6_outputs(368) <= not (a xor b);
    layer6_outputs(369) <= not (a or b);
    layer6_outputs(370) <= a;
    layer6_outputs(371) <= not a or b;
    layer6_outputs(372) <= not b or a;
    layer6_outputs(373) <= a;
    layer6_outputs(374) <= not a;
    layer6_outputs(375) <= not b;
    layer6_outputs(376) <= b and not a;
    layer6_outputs(377) <= b and not a;
    layer6_outputs(378) <= b;
    layer6_outputs(379) <= 1'b0;
    layer6_outputs(380) <= b and not a;
    layer6_outputs(381) <= a;
    layer6_outputs(382) <= not (a xor b);
    layer6_outputs(383) <= a and not b;
    layer6_outputs(384) <= a;
    layer6_outputs(385) <= not (a or b);
    layer6_outputs(386) <= not a;
    layer6_outputs(387) <= not b;
    layer6_outputs(388) <= a;
    layer6_outputs(389) <= not (a and b);
    layer6_outputs(390) <= b and not a;
    layer6_outputs(391) <= a or b;
    layer6_outputs(392) <= a xor b;
    layer6_outputs(393) <= a or b;
    layer6_outputs(394) <= not b;
    layer6_outputs(395) <= not a;
    layer6_outputs(396) <= not (a and b);
    layer6_outputs(397) <= b;
    layer6_outputs(398) <= 1'b1;
    layer6_outputs(399) <= b;
    layer6_outputs(400) <= a;
    layer6_outputs(401) <= a and not b;
    layer6_outputs(402) <= not a;
    layer6_outputs(403) <= b;
    layer6_outputs(404) <= 1'b0;
    layer6_outputs(405) <= b and not a;
    layer6_outputs(406) <= 1'b0;
    layer6_outputs(407) <= b;
    layer6_outputs(408) <= not (a xor b);
    layer6_outputs(409) <= not a;
    layer6_outputs(410) <= 1'b0;
    layer6_outputs(411) <= 1'b0;
    layer6_outputs(412) <= not a;
    layer6_outputs(413) <= b and not a;
    layer6_outputs(414) <= not a or b;
    layer6_outputs(415) <= a;
    layer6_outputs(416) <= not a or b;
    layer6_outputs(417) <= 1'b1;
    layer6_outputs(418) <= not (a and b);
    layer6_outputs(419) <= not (a and b);
    layer6_outputs(420) <= not b or a;
    layer6_outputs(421) <= a and not b;
    layer6_outputs(422) <= a and not b;
    layer6_outputs(423) <= not (a xor b);
    layer6_outputs(424) <= a or b;
    layer6_outputs(425) <= not a;
    layer6_outputs(426) <= a or b;
    layer6_outputs(427) <= not b;
    layer6_outputs(428) <= not (a and b);
    layer6_outputs(429) <= b;
    layer6_outputs(430) <= a;
    layer6_outputs(431) <= not b or a;
    layer6_outputs(432) <= b;
    layer6_outputs(433) <= not a;
    layer6_outputs(434) <= b and not a;
    layer6_outputs(435) <= a;
    layer6_outputs(436) <= a xor b;
    layer6_outputs(437) <= not a;
    layer6_outputs(438) <= not b or a;
    layer6_outputs(439) <= not a;
    layer6_outputs(440) <= a and b;
    layer6_outputs(441) <= b and not a;
    layer6_outputs(442) <= b;
    layer6_outputs(443) <= not b;
    layer6_outputs(444) <= not a or b;
    layer6_outputs(445) <= not a or b;
    layer6_outputs(446) <= not a;
    layer6_outputs(447) <= not a;
    layer6_outputs(448) <= a;
    layer6_outputs(449) <= a and b;
    layer6_outputs(450) <= a and not b;
    layer6_outputs(451) <= not (a xor b);
    layer6_outputs(452) <= a xor b;
    layer6_outputs(453) <= not a or b;
    layer6_outputs(454) <= a and b;
    layer6_outputs(455) <= not a;
    layer6_outputs(456) <= not (a and b);
    layer6_outputs(457) <= not b;
    layer6_outputs(458) <= not (a or b);
    layer6_outputs(459) <= b;
    layer6_outputs(460) <= a and b;
    layer6_outputs(461) <= a;
    layer6_outputs(462) <= not b or a;
    layer6_outputs(463) <= not b;
    layer6_outputs(464) <= b and not a;
    layer6_outputs(465) <= b;
    layer6_outputs(466) <= 1'b1;
    layer6_outputs(467) <= not (a and b);
    layer6_outputs(468) <= not a;
    layer6_outputs(469) <= not a or b;
    layer6_outputs(470) <= a;
    layer6_outputs(471) <= a and b;
    layer6_outputs(472) <= not (a xor b);
    layer6_outputs(473) <= not (a xor b);
    layer6_outputs(474) <= b;
    layer6_outputs(475) <= not b;
    layer6_outputs(476) <= a;
    layer6_outputs(477) <= not (a or b);
    layer6_outputs(478) <= not a or b;
    layer6_outputs(479) <= not (a or b);
    layer6_outputs(480) <= not (a or b);
    layer6_outputs(481) <= a or b;
    layer6_outputs(482) <= a xor b;
    layer6_outputs(483) <= b and not a;
    layer6_outputs(484) <= a;
    layer6_outputs(485) <= b and not a;
    layer6_outputs(486) <= a;
    layer6_outputs(487) <= not (a xor b);
    layer6_outputs(488) <= not a;
    layer6_outputs(489) <= not (a and b);
    layer6_outputs(490) <= not b;
    layer6_outputs(491) <= not b;
    layer6_outputs(492) <= a;
    layer6_outputs(493) <= a and not b;
    layer6_outputs(494) <= b;
    layer6_outputs(495) <= b and not a;
    layer6_outputs(496) <= b;
    layer6_outputs(497) <= not (a or b);
    layer6_outputs(498) <= b and not a;
    layer6_outputs(499) <= not a;
    layer6_outputs(500) <= not a or b;
    layer6_outputs(501) <= not (a or b);
    layer6_outputs(502) <= not (a or b);
    layer6_outputs(503) <= a or b;
    layer6_outputs(504) <= b;
    layer6_outputs(505) <= not (a and b);
    layer6_outputs(506) <= a and b;
    layer6_outputs(507) <= a;
    layer6_outputs(508) <= not a;
    layer6_outputs(509) <= not (a xor b);
    layer6_outputs(510) <= a;
    layer6_outputs(511) <= not a or b;
    layer6_outputs(512) <= not a or b;
    layer6_outputs(513) <= b and not a;
    layer6_outputs(514) <= a;
    layer6_outputs(515) <= not a or b;
    layer6_outputs(516) <= not b;
    layer6_outputs(517) <= a;
    layer6_outputs(518) <= not (a and b);
    layer6_outputs(519) <= 1'b1;
    layer6_outputs(520) <= not a or b;
    layer6_outputs(521) <= not a;
    layer6_outputs(522) <= a or b;
    layer6_outputs(523) <= b and not a;
    layer6_outputs(524) <= not (a or b);
    layer6_outputs(525) <= a xor b;
    layer6_outputs(526) <= a and not b;
    layer6_outputs(527) <= a and not b;
    layer6_outputs(528) <= not (a or b);
    layer6_outputs(529) <= b;
    layer6_outputs(530) <= not b;
    layer6_outputs(531) <= a xor b;
    layer6_outputs(532) <= not a or b;
    layer6_outputs(533) <= not a;
    layer6_outputs(534) <= b;
    layer6_outputs(535) <= b;
    layer6_outputs(536) <= b;
    layer6_outputs(537) <= a or b;
    layer6_outputs(538) <= a xor b;
    layer6_outputs(539) <= not b;
    layer6_outputs(540) <= b;
    layer6_outputs(541) <= not a or b;
    layer6_outputs(542) <= not (a or b);
    layer6_outputs(543) <= a and not b;
    layer6_outputs(544) <= a and b;
    layer6_outputs(545) <= not (a and b);
    layer6_outputs(546) <= not b;
    layer6_outputs(547) <= not a;
    layer6_outputs(548) <= a and not b;
    layer6_outputs(549) <= not (a or b);
    layer6_outputs(550) <= not (a and b);
    layer6_outputs(551) <= a;
    layer6_outputs(552) <= a;
    layer6_outputs(553) <= a and not b;
    layer6_outputs(554) <= not a;
    layer6_outputs(555) <= not (a xor b);
    layer6_outputs(556) <= not b;
    layer6_outputs(557) <= not (a and b);
    layer6_outputs(558) <= b and not a;
    layer6_outputs(559) <= not b or a;
    layer6_outputs(560) <= not (a or b);
    layer6_outputs(561) <= b;
    layer6_outputs(562) <= not (a xor b);
    layer6_outputs(563) <= not b or a;
    layer6_outputs(564) <= not (a and b);
    layer6_outputs(565) <= a and not b;
    layer6_outputs(566) <= a and not b;
    layer6_outputs(567) <= a and not b;
    layer6_outputs(568) <= not (a and b);
    layer6_outputs(569) <= b and not a;
    layer6_outputs(570) <= a and b;
    layer6_outputs(571) <= b;
    layer6_outputs(572) <= not b or a;
    layer6_outputs(573) <= not a or b;
    layer6_outputs(574) <= not (a and b);
    layer6_outputs(575) <= not b;
    layer6_outputs(576) <= a;
    layer6_outputs(577) <= b;
    layer6_outputs(578) <= not a or b;
    layer6_outputs(579) <= not b;
    layer6_outputs(580) <= a or b;
    layer6_outputs(581) <= b and not a;
    layer6_outputs(582) <= not a or b;
    layer6_outputs(583) <= not b;
    layer6_outputs(584) <= not (a and b);
    layer6_outputs(585) <= not a or b;
    layer6_outputs(586) <= not a or b;
    layer6_outputs(587) <= not b or a;
    layer6_outputs(588) <= b and not a;
    layer6_outputs(589) <= not b;
    layer6_outputs(590) <= not (a or b);
    layer6_outputs(591) <= not (a and b);
    layer6_outputs(592) <= 1'b0;
    layer6_outputs(593) <= a and not b;
    layer6_outputs(594) <= b;
    layer6_outputs(595) <= not a or b;
    layer6_outputs(596) <= not a;
    layer6_outputs(597) <= 1'b1;
    layer6_outputs(598) <= not a;
    layer6_outputs(599) <= b;
    layer6_outputs(600) <= not a or b;
    layer6_outputs(601) <= not a;
    layer6_outputs(602) <= a and b;
    layer6_outputs(603) <= not (a and b);
    layer6_outputs(604) <= 1'b1;
    layer6_outputs(605) <= not (a or b);
    layer6_outputs(606) <= not b;
    layer6_outputs(607) <= 1'b1;
    layer6_outputs(608) <= a and not b;
    layer6_outputs(609) <= not a;
    layer6_outputs(610) <= not b;
    layer6_outputs(611) <= b and not a;
    layer6_outputs(612) <= a and b;
    layer6_outputs(613) <= not (a and b);
    layer6_outputs(614) <= not a;
    layer6_outputs(615) <= not a;
    layer6_outputs(616) <= b;
    layer6_outputs(617) <= b;
    layer6_outputs(618) <= not (a or b);
    layer6_outputs(619) <= not b;
    layer6_outputs(620) <= a;
    layer6_outputs(621) <= a and b;
    layer6_outputs(622) <= a;
    layer6_outputs(623) <= not b;
    layer6_outputs(624) <= not b;
    layer6_outputs(625) <= not (a or b);
    layer6_outputs(626) <= a and b;
    layer6_outputs(627) <= a xor b;
    layer6_outputs(628) <= b;
    layer6_outputs(629) <= not a;
    layer6_outputs(630) <= not b;
    layer6_outputs(631) <= a and not b;
    layer6_outputs(632) <= b;
    layer6_outputs(633) <= 1'b0;
    layer6_outputs(634) <= not a;
    layer6_outputs(635) <= a;
    layer6_outputs(636) <= a and b;
    layer6_outputs(637) <= b;
    layer6_outputs(638) <= a;
    layer6_outputs(639) <= a xor b;
    layer6_outputs(640) <= a and b;
    layer6_outputs(641) <= not b;
    layer6_outputs(642) <= a or b;
    layer6_outputs(643) <= a and not b;
    layer6_outputs(644) <= a and b;
    layer6_outputs(645) <= not (a or b);
    layer6_outputs(646) <= not (a xor b);
    layer6_outputs(647) <= not b;
    layer6_outputs(648) <= not b;
    layer6_outputs(649) <= b;
    layer6_outputs(650) <= b;
    layer6_outputs(651) <= b;
    layer6_outputs(652) <= b;
    layer6_outputs(653) <= a and b;
    layer6_outputs(654) <= b;
    layer6_outputs(655) <= a;
    layer6_outputs(656) <= not a or b;
    layer6_outputs(657) <= not (a or b);
    layer6_outputs(658) <= not a;
    layer6_outputs(659) <= not b;
    layer6_outputs(660) <= not a or b;
    layer6_outputs(661) <= a;
    layer6_outputs(662) <= not (a or b);
    layer6_outputs(663) <= b;
    layer6_outputs(664) <= b;
    layer6_outputs(665) <= not a;
    layer6_outputs(666) <= a xor b;
    layer6_outputs(667) <= not a;
    layer6_outputs(668) <= 1'b1;
    layer6_outputs(669) <= a;
    layer6_outputs(670) <= a;
    layer6_outputs(671) <= not (a or b);
    layer6_outputs(672) <= a;
    layer6_outputs(673) <= a;
    layer6_outputs(674) <= not a;
    layer6_outputs(675) <= b;
    layer6_outputs(676) <= a and b;
    layer6_outputs(677) <= 1'b0;
    layer6_outputs(678) <= not (a and b);
    layer6_outputs(679) <= not a;
    layer6_outputs(680) <= b;
    layer6_outputs(681) <= a and b;
    layer6_outputs(682) <= a;
    layer6_outputs(683) <= not a or b;
    layer6_outputs(684) <= not a or b;
    layer6_outputs(685) <= a or b;
    layer6_outputs(686) <= not b;
    layer6_outputs(687) <= b;
    layer6_outputs(688) <= b and not a;
    layer6_outputs(689) <= b and not a;
    layer6_outputs(690) <= not b or a;
    layer6_outputs(691) <= b;
    layer6_outputs(692) <= a and b;
    layer6_outputs(693) <= not b;
    layer6_outputs(694) <= a;
    layer6_outputs(695) <= not a;
    layer6_outputs(696) <= not b;
    layer6_outputs(697) <= not (a and b);
    layer6_outputs(698) <= b;
    layer6_outputs(699) <= b;
    layer6_outputs(700) <= not (a or b);
    layer6_outputs(701) <= b;
    layer6_outputs(702) <= b;
    layer6_outputs(703) <= a and not b;
    layer6_outputs(704) <= a xor b;
    layer6_outputs(705) <= a and not b;
    layer6_outputs(706) <= a;
    layer6_outputs(707) <= not a or b;
    layer6_outputs(708) <= a and b;
    layer6_outputs(709) <= not a;
    layer6_outputs(710) <= not (a or b);
    layer6_outputs(711) <= not (a or b);
    layer6_outputs(712) <= not (a or b);
    layer6_outputs(713) <= not a;
    layer6_outputs(714) <= not (a and b);
    layer6_outputs(715) <= not a or b;
    layer6_outputs(716) <= 1'b1;
    layer6_outputs(717) <= a or b;
    layer6_outputs(718) <= a or b;
    layer6_outputs(719) <= b;
    layer6_outputs(720) <= not (a or b);
    layer6_outputs(721) <= a;
    layer6_outputs(722) <= not (a and b);
    layer6_outputs(723) <= a or b;
    layer6_outputs(724) <= a and b;
    layer6_outputs(725) <= a and b;
    layer6_outputs(726) <= not (a and b);
    layer6_outputs(727) <= 1'b0;
    layer6_outputs(728) <= not (a or b);
    layer6_outputs(729) <= not a;
    layer6_outputs(730) <= a;
    layer6_outputs(731) <= 1'b1;
    layer6_outputs(732) <= not (a and b);
    layer6_outputs(733) <= a and not b;
    layer6_outputs(734) <= a;
    layer6_outputs(735) <= a and not b;
    layer6_outputs(736) <= a and not b;
    layer6_outputs(737) <= not a;
    layer6_outputs(738) <= a and not b;
    layer6_outputs(739) <= b;
    layer6_outputs(740) <= a or b;
    layer6_outputs(741) <= a;
    layer6_outputs(742) <= b;
    layer6_outputs(743) <= not b or a;
    layer6_outputs(744) <= not b;
    layer6_outputs(745) <= not (a xor b);
    layer6_outputs(746) <= a or b;
    layer6_outputs(747) <= b and not a;
    layer6_outputs(748) <= not a;
    layer6_outputs(749) <= b and not a;
    layer6_outputs(750) <= not (a xor b);
    layer6_outputs(751) <= a and b;
    layer6_outputs(752) <= not a or b;
    layer6_outputs(753) <= not a;
    layer6_outputs(754) <= a xor b;
    layer6_outputs(755) <= b and not a;
    layer6_outputs(756) <= not b;
    layer6_outputs(757) <= b;
    layer6_outputs(758) <= not a or b;
    layer6_outputs(759) <= not a;
    layer6_outputs(760) <= b;
    layer6_outputs(761) <= not a;
    layer6_outputs(762) <= not (a xor b);
    layer6_outputs(763) <= b and not a;
    layer6_outputs(764) <= not b or a;
    layer6_outputs(765) <= not b;
    layer6_outputs(766) <= not b;
    layer6_outputs(767) <= a xor b;
    layer6_outputs(768) <= not a;
    layer6_outputs(769) <= not a or b;
    layer6_outputs(770) <= not b;
    layer6_outputs(771) <= a;
    layer6_outputs(772) <= not (a or b);
    layer6_outputs(773) <= b and not a;
    layer6_outputs(774) <= not (a and b);
    layer6_outputs(775) <= not a;
    layer6_outputs(776) <= not a;
    layer6_outputs(777) <= not (a and b);
    layer6_outputs(778) <= a or b;
    layer6_outputs(779) <= b;
    layer6_outputs(780) <= 1'b0;
    layer6_outputs(781) <= b;
    layer6_outputs(782) <= not b;
    layer6_outputs(783) <= a;
    layer6_outputs(784) <= not b;
    layer6_outputs(785) <= a;
    layer6_outputs(786) <= not (a and b);
    layer6_outputs(787) <= a or b;
    layer6_outputs(788) <= not a or b;
    layer6_outputs(789) <= not b;
    layer6_outputs(790) <= not (a xor b);
    layer6_outputs(791) <= not b;
    layer6_outputs(792) <= b;
    layer6_outputs(793) <= not a or b;
    layer6_outputs(794) <= not a or b;
    layer6_outputs(795) <= b and not a;
    layer6_outputs(796) <= not (a or b);
    layer6_outputs(797) <= not (a or b);
    layer6_outputs(798) <= a and not b;
    layer6_outputs(799) <= not b or a;
    layer6_outputs(800) <= a;
    layer6_outputs(801) <= not a or b;
    layer6_outputs(802) <= b;
    layer6_outputs(803) <= not a or b;
    layer6_outputs(804) <= not b or a;
    layer6_outputs(805) <= not b;
    layer6_outputs(806) <= not b;
    layer6_outputs(807) <= b;
    layer6_outputs(808) <= a and not b;
    layer6_outputs(809) <= a xor b;
    layer6_outputs(810) <= b;
    layer6_outputs(811) <= not (a or b);
    layer6_outputs(812) <= not (a or b);
    layer6_outputs(813) <= not (a or b);
    layer6_outputs(814) <= a;
    layer6_outputs(815) <= a or b;
    layer6_outputs(816) <= 1'b0;
    layer6_outputs(817) <= not a or b;
    layer6_outputs(818) <= not a;
    layer6_outputs(819) <= b;
    layer6_outputs(820) <= not (a xor b);
    layer6_outputs(821) <= 1'b1;
    layer6_outputs(822) <= not a or b;
    layer6_outputs(823) <= b and not a;
    layer6_outputs(824) <= b;
    layer6_outputs(825) <= not a;
    layer6_outputs(826) <= not (a xor b);
    layer6_outputs(827) <= a;
    layer6_outputs(828) <= not a;
    layer6_outputs(829) <= a;
    layer6_outputs(830) <= not (a and b);
    layer6_outputs(831) <= a xor b;
    layer6_outputs(832) <= not a;
    layer6_outputs(833) <= 1'b0;
    layer6_outputs(834) <= 1'b0;
    layer6_outputs(835) <= not (a or b);
    layer6_outputs(836) <= a and b;
    layer6_outputs(837) <= a and not b;
    layer6_outputs(838) <= a and not b;
    layer6_outputs(839) <= a and b;
    layer6_outputs(840) <= not b;
    layer6_outputs(841) <= a;
    layer6_outputs(842) <= not (a and b);
    layer6_outputs(843) <= not a;
    layer6_outputs(844) <= a or b;
    layer6_outputs(845) <= not (a and b);
    layer6_outputs(846) <= a xor b;
    layer6_outputs(847) <= not (a and b);
    layer6_outputs(848) <= a and b;
    layer6_outputs(849) <= a;
    layer6_outputs(850) <= not (a and b);
    layer6_outputs(851) <= a and b;
    layer6_outputs(852) <= a and not b;
    layer6_outputs(853) <= a and b;
    layer6_outputs(854) <= not b;
    layer6_outputs(855) <= not b;
    layer6_outputs(856) <= not a;
    layer6_outputs(857) <= a and not b;
    layer6_outputs(858) <= a or b;
    layer6_outputs(859) <= a and not b;
    layer6_outputs(860) <= 1'b1;
    layer6_outputs(861) <= not (a or b);
    layer6_outputs(862) <= a;
    layer6_outputs(863) <= a;
    layer6_outputs(864) <= b;
    layer6_outputs(865) <= a or b;
    layer6_outputs(866) <= b;
    layer6_outputs(867) <= 1'b1;
    layer6_outputs(868) <= not (a and b);
    layer6_outputs(869) <= not b or a;
    layer6_outputs(870) <= a and b;
    layer6_outputs(871) <= b;
    layer6_outputs(872) <= not (a xor b);
    layer6_outputs(873) <= not b;
    layer6_outputs(874) <= b;
    layer6_outputs(875) <= a and not b;
    layer6_outputs(876) <= not (a and b);
    layer6_outputs(877) <= not a;
    layer6_outputs(878) <= a xor b;
    layer6_outputs(879) <= not a;
    layer6_outputs(880) <= not (a and b);
    layer6_outputs(881) <= a and not b;
    layer6_outputs(882) <= a and not b;
    layer6_outputs(883) <= not b;
    layer6_outputs(884) <= not b;
    layer6_outputs(885) <= b and not a;
    layer6_outputs(886) <= not a;
    layer6_outputs(887) <= 1'b1;
    layer6_outputs(888) <= b;
    layer6_outputs(889) <= a xor b;
    layer6_outputs(890) <= a;
    layer6_outputs(891) <= not a or b;
    layer6_outputs(892) <= not (a xor b);
    layer6_outputs(893) <= not b;
    layer6_outputs(894) <= a and not b;
    layer6_outputs(895) <= a and b;
    layer6_outputs(896) <= not (a and b);
    layer6_outputs(897) <= b;
    layer6_outputs(898) <= not a or b;
    layer6_outputs(899) <= not b or a;
    layer6_outputs(900) <= a or b;
    layer6_outputs(901) <= not (a and b);
    layer6_outputs(902) <= not b;
    layer6_outputs(903) <= not b or a;
    layer6_outputs(904) <= b;
    layer6_outputs(905) <= a or b;
    layer6_outputs(906) <= not (a or b);
    layer6_outputs(907) <= not b;
    layer6_outputs(908) <= b and not a;
    layer6_outputs(909) <= not b;
    layer6_outputs(910) <= b and not a;
    layer6_outputs(911) <= a and not b;
    layer6_outputs(912) <= not (a and b);
    layer6_outputs(913) <= not b;
    layer6_outputs(914) <= a and b;
    layer6_outputs(915) <= a;
    layer6_outputs(916) <= a;
    layer6_outputs(917) <= a or b;
    layer6_outputs(918) <= b and not a;
    layer6_outputs(919) <= b;
    layer6_outputs(920) <= b and not a;
    layer6_outputs(921) <= b and not a;
    layer6_outputs(922) <= b;
    layer6_outputs(923) <= b and not a;
    layer6_outputs(924) <= not (a or b);
    layer6_outputs(925) <= not b or a;
    layer6_outputs(926) <= not b or a;
    layer6_outputs(927) <= a or b;
    layer6_outputs(928) <= b;
    layer6_outputs(929) <= not a or b;
    layer6_outputs(930) <= a and b;
    layer6_outputs(931) <= a and b;
    layer6_outputs(932) <= a or b;
    layer6_outputs(933) <= not b;
    layer6_outputs(934) <= not a or b;
    layer6_outputs(935) <= not b or a;
    layer6_outputs(936) <= not (a xor b);
    layer6_outputs(937) <= not a;
    layer6_outputs(938) <= not b or a;
    layer6_outputs(939) <= a xor b;
    layer6_outputs(940) <= a or b;
    layer6_outputs(941) <= 1'b1;
    layer6_outputs(942) <= not b;
    layer6_outputs(943) <= b;
    layer6_outputs(944) <= not b or a;
    layer6_outputs(945) <= b;
    layer6_outputs(946) <= not (a or b);
    layer6_outputs(947) <= a;
    layer6_outputs(948) <= not a or b;
    layer6_outputs(949) <= not a;
    layer6_outputs(950) <= a;
    layer6_outputs(951) <= a;
    layer6_outputs(952) <= a and b;
    layer6_outputs(953) <= not a;
    layer6_outputs(954) <= a and b;
    layer6_outputs(955) <= not (a and b);
    layer6_outputs(956) <= not (a or b);
    layer6_outputs(957) <= not (a and b);
    layer6_outputs(958) <= a or b;
    layer6_outputs(959) <= not a;
    layer6_outputs(960) <= not b or a;
    layer6_outputs(961) <= a xor b;
    layer6_outputs(962) <= not (a or b);
    layer6_outputs(963) <= a and not b;
    layer6_outputs(964) <= not b;
    layer6_outputs(965) <= a or b;
    layer6_outputs(966) <= not (a or b);
    layer6_outputs(967) <= not a or b;
    layer6_outputs(968) <= a;
    layer6_outputs(969) <= b and not a;
    layer6_outputs(970) <= 1'b1;
    layer6_outputs(971) <= b and not a;
    layer6_outputs(972) <= a;
    layer6_outputs(973) <= a and b;
    layer6_outputs(974) <= a;
    layer6_outputs(975) <= not a or b;
    layer6_outputs(976) <= not b;
    layer6_outputs(977) <= 1'b0;
    layer6_outputs(978) <= a and b;
    layer6_outputs(979) <= b;
    layer6_outputs(980) <= not (a or b);
    layer6_outputs(981) <= not (a xor b);
    layer6_outputs(982) <= not b or a;
    layer6_outputs(983) <= not a;
    layer6_outputs(984) <= not b;
    layer6_outputs(985) <= not (a and b);
    layer6_outputs(986) <= a;
    layer6_outputs(987) <= a and b;
    layer6_outputs(988) <= a xor b;
    layer6_outputs(989) <= not (a and b);
    layer6_outputs(990) <= a or b;
    layer6_outputs(991) <= not b;
    layer6_outputs(992) <= not (a or b);
    layer6_outputs(993) <= not a or b;
    layer6_outputs(994) <= b;
    layer6_outputs(995) <= not a;
    layer6_outputs(996) <= b and not a;
    layer6_outputs(997) <= 1'b1;
    layer6_outputs(998) <= not (a and b);
    layer6_outputs(999) <= b and not a;
    layer6_outputs(1000) <= not b;
    layer6_outputs(1001) <= not (a xor b);
    layer6_outputs(1002) <= b;
    layer6_outputs(1003) <= b;
    layer6_outputs(1004) <= 1'b0;
    layer6_outputs(1005) <= b;
    layer6_outputs(1006) <= b;
    layer6_outputs(1007) <= not b or a;
    layer6_outputs(1008) <= a or b;
    layer6_outputs(1009) <= a or b;
    layer6_outputs(1010) <= b;
    layer6_outputs(1011) <= not (a or b);
    layer6_outputs(1012) <= not b;
    layer6_outputs(1013) <= not b or a;
    layer6_outputs(1014) <= not a or b;
    layer6_outputs(1015) <= not b;
    layer6_outputs(1016) <= a and b;
    layer6_outputs(1017) <= not (a and b);
    layer6_outputs(1018) <= a or b;
    layer6_outputs(1019) <= not a;
    layer6_outputs(1020) <= a and b;
    layer6_outputs(1021) <= not (a and b);
    layer6_outputs(1022) <= not b;
    layer6_outputs(1023) <= not (a xor b);
    layer6_outputs(1024) <= a and not b;
    layer6_outputs(1025) <= a;
    layer6_outputs(1026) <= not a;
    layer6_outputs(1027) <= not (a or b);
    layer6_outputs(1028) <= b;
    layer6_outputs(1029) <= not a;
    layer6_outputs(1030) <= a;
    layer6_outputs(1031) <= b;
    layer6_outputs(1032) <= not (a xor b);
    layer6_outputs(1033) <= not a;
    layer6_outputs(1034) <= a and b;
    layer6_outputs(1035) <= b;
    layer6_outputs(1036) <= a;
    layer6_outputs(1037) <= not (a and b);
    layer6_outputs(1038) <= not a or b;
    layer6_outputs(1039) <= not (a and b);
    layer6_outputs(1040) <= 1'b1;
    layer6_outputs(1041) <= not a or b;
    layer6_outputs(1042) <= not (a or b);
    layer6_outputs(1043) <= not a;
    layer6_outputs(1044) <= a and not b;
    layer6_outputs(1045) <= not a or b;
    layer6_outputs(1046) <= not a or b;
    layer6_outputs(1047) <= not b;
    layer6_outputs(1048) <= not (a and b);
    layer6_outputs(1049) <= not a or b;
    layer6_outputs(1050) <= b;
    layer6_outputs(1051) <= not (a or b);
    layer6_outputs(1052) <= not b or a;
    layer6_outputs(1053) <= not b;
    layer6_outputs(1054) <= a;
    layer6_outputs(1055) <= not b;
    layer6_outputs(1056) <= b;
    layer6_outputs(1057) <= 1'b0;
    layer6_outputs(1058) <= a xor b;
    layer6_outputs(1059) <= a or b;
    layer6_outputs(1060) <= not b or a;
    layer6_outputs(1061) <= a or b;
    layer6_outputs(1062) <= not b;
    layer6_outputs(1063) <= not (a and b);
    layer6_outputs(1064) <= not (a or b);
    layer6_outputs(1065) <= not b or a;
    layer6_outputs(1066) <= not (a and b);
    layer6_outputs(1067) <= not a;
    layer6_outputs(1068) <= not (a and b);
    layer6_outputs(1069) <= not (a or b);
    layer6_outputs(1070) <= a;
    layer6_outputs(1071) <= not a;
    layer6_outputs(1072) <= not (a or b);
    layer6_outputs(1073) <= not a or b;
    layer6_outputs(1074) <= not a or b;
    layer6_outputs(1075) <= not a;
    layer6_outputs(1076) <= b and not a;
    layer6_outputs(1077) <= not b or a;
    layer6_outputs(1078) <= not (a xor b);
    layer6_outputs(1079) <= not (a and b);
    layer6_outputs(1080) <= a or b;
    layer6_outputs(1081) <= not b;
    layer6_outputs(1082) <= not b;
    layer6_outputs(1083) <= a;
    layer6_outputs(1084) <= a;
    layer6_outputs(1085) <= not a;
    layer6_outputs(1086) <= not (a and b);
    layer6_outputs(1087) <= not (a or b);
    layer6_outputs(1088) <= a xor b;
    layer6_outputs(1089) <= not (a or b);
    layer6_outputs(1090) <= b;
    layer6_outputs(1091) <= not (a xor b);
    layer6_outputs(1092) <= b;
    layer6_outputs(1093) <= not (a xor b);
    layer6_outputs(1094) <= not a or b;
    layer6_outputs(1095) <= not (a and b);
    layer6_outputs(1096) <= not b;
    layer6_outputs(1097) <= not (a or b);
    layer6_outputs(1098) <= a and b;
    layer6_outputs(1099) <= a and not b;
    layer6_outputs(1100) <= b;
    layer6_outputs(1101) <= not (a and b);
    layer6_outputs(1102) <= not a;
    layer6_outputs(1103) <= not b or a;
    layer6_outputs(1104) <= b;
    layer6_outputs(1105) <= a and b;
    layer6_outputs(1106) <= not (a xor b);
    layer6_outputs(1107) <= not (a xor b);
    layer6_outputs(1108) <= not (a and b);
    layer6_outputs(1109) <= not a;
    layer6_outputs(1110) <= b;
    layer6_outputs(1111) <= not b or a;
    layer6_outputs(1112) <= a;
    layer6_outputs(1113) <= b and not a;
    layer6_outputs(1114) <= not a;
    layer6_outputs(1115) <= not (a and b);
    layer6_outputs(1116) <= a and b;
    layer6_outputs(1117) <= b;
    layer6_outputs(1118) <= a or b;
    layer6_outputs(1119) <= not b or a;
    layer6_outputs(1120) <= not b;
    layer6_outputs(1121) <= not (a xor b);
    layer6_outputs(1122) <= not (a and b);
    layer6_outputs(1123) <= a;
    layer6_outputs(1124) <= a xor b;
    layer6_outputs(1125) <= a;
    layer6_outputs(1126) <= not (a and b);
    layer6_outputs(1127) <= not b;
    layer6_outputs(1128) <= not (a xor b);
    layer6_outputs(1129) <= not b;
    layer6_outputs(1130) <= not b or a;
    layer6_outputs(1131) <= not a or b;
    layer6_outputs(1132) <= not (a or b);
    layer6_outputs(1133) <= b and not a;
    layer6_outputs(1134) <= b and not a;
    layer6_outputs(1135) <= not b;
    layer6_outputs(1136) <= b;
    layer6_outputs(1137) <= b and not a;
    layer6_outputs(1138) <= not b;
    layer6_outputs(1139) <= not (a or b);
    layer6_outputs(1140) <= a and not b;
    layer6_outputs(1141) <= b and not a;
    layer6_outputs(1142) <= 1'b0;
    layer6_outputs(1143) <= not b;
    layer6_outputs(1144) <= not b;
    layer6_outputs(1145) <= not b;
    layer6_outputs(1146) <= not a;
    layer6_outputs(1147) <= not b;
    layer6_outputs(1148) <= not b;
    layer6_outputs(1149) <= b and not a;
    layer6_outputs(1150) <= not (a xor b);
    layer6_outputs(1151) <= a;
    layer6_outputs(1152) <= b and not a;
    layer6_outputs(1153) <= not (a and b);
    layer6_outputs(1154) <= not a;
    layer6_outputs(1155) <= not b;
    layer6_outputs(1156) <= b;
    layer6_outputs(1157) <= a or b;
    layer6_outputs(1158) <= not b or a;
    layer6_outputs(1159) <= a;
    layer6_outputs(1160) <= a and b;
    layer6_outputs(1161) <= a and not b;
    layer6_outputs(1162) <= 1'b1;
    layer6_outputs(1163) <= 1'b0;
    layer6_outputs(1164) <= a or b;
    layer6_outputs(1165) <= a;
    layer6_outputs(1166) <= not a;
    layer6_outputs(1167) <= a;
    layer6_outputs(1168) <= not (a xor b);
    layer6_outputs(1169) <= not b;
    layer6_outputs(1170) <= b and not a;
    layer6_outputs(1171) <= b and not a;
    layer6_outputs(1172) <= b;
    layer6_outputs(1173) <= a;
    layer6_outputs(1174) <= b and not a;
    layer6_outputs(1175) <= not b;
    layer6_outputs(1176) <= not a;
    layer6_outputs(1177) <= not b or a;
    layer6_outputs(1178) <= not b or a;
    layer6_outputs(1179) <= not (a or b);
    layer6_outputs(1180) <= b;
    layer6_outputs(1181) <= not b;
    layer6_outputs(1182) <= not (a xor b);
    layer6_outputs(1183) <= not a or b;
    layer6_outputs(1184) <= not (a xor b);
    layer6_outputs(1185) <= not a or b;
    layer6_outputs(1186) <= not (a and b);
    layer6_outputs(1187) <= not a;
    layer6_outputs(1188) <= not a;
    layer6_outputs(1189) <= not a or b;
    layer6_outputs(1190) <= a and b;
    layer6_outputs(1191) <= not b;
    layer6_outputs(1192) <= not a or b;
    layer6_outputs(1193) <= a;
    layer6_outputs(1194) <= not (a and b);
    layer6_outputs(1195) <= a and b;
    layer6_outputs(1196) <= a xor b;
    layer6_outputs(1197) <= a and not b;
    layer6_outputs(1198) <= a xor b;
    layer6_outputs(1199) <= a and b;
    layer6_outputs(1200) <= b;
    layer6_outputs(1201) <= not (a or b);
    layer6_outputs(1202) <= a;
    layer6_outputs(1203) <= not a;
    layer6_outputs(1204) <= not (a and b);
    layer6_outputs(1205) <= not b;
    layer6_outputs(1206) <= not a or b;
    layer6_outputs(1207) <= not a;
    layer6_outputs(1208) <= not (a and b);
    layer6_outputs(1209) <= not (a and b);
    layer6_outputs(1210) <= 1'b1;
    layer6_outputs(1211) <= not b;
    layer6_outputs(1212) <= 1'b0;
    layer6_outputs(1213) <= a;
    layer6_outputs(1214) <= 1'b1;
    layer6_outputs(1215) <= not b;
    layer6_outputs(1216) <= not (a or b);
    layer6_outputs(1217) <= not (a xor b);
    layer6_outputs(1218) <= a;
    layer6_outputs(1219) <= not a or b;
    layer6_outputs(1220) <= b;
    layer6_outputs(1221) <= not a;
    layer6_outputs(1222) <= not a;
    layer6_outputs(1223) <= not a;
    layer6_outputs(1224) <= a or b;
    layer6_outputs(1225) <= a or b;
    layer6_outputs(1226) <= b and not a;
    layer6_outputs(1227) <= a and not b;
    layer6_outputs(1228) <= not a;
    layer6_outputs(1229) <= a;
    layer6_outputs(1230) <= a and not b;
    layer6_outputs(1231) <= a xor b;
    layer6_outputs(1232) <= not (a xor b);
    layer6_outputs(1233) <= not b;
    layer6_outputs(1234) <= b and not a;
    layer6_outputs(1235) <= a and b;
    layer6_outputs(1236) <= not (a xor b);
    layer6_outputs(1237) <= a;
    layer6_outputs(1238) <= a or b;
    layer6_outputs(1239) <= 1'b0;
    layer6_outputs(1240) <= a;
    layer6_outputs(1241) <= not b;
    layer6_outputs(1242) <= a and not b;
    layer6_outputs(1243) <= 1'b1;
    layer6_outputs(1244) <= a;
    layer6_outputs(1245) <= not (a or b);
    layer6_outputs(1246) <= a and not b;
    layer6_outputs(1247) <= not b;
    layer6_outputs(1248) <= b and not a;
    layer6_outputs(1249) <= a and b;
    layer6_outputs(1250) <= not a;
    layer6_outputs(1251) <= a;
    layer6_outputs(1252) <= a;
    layer6_outputs(1253) <= not a or b;
    layer6_outputs(1254) <= a or b;
    layer6_outputs(1255) <= b;
    layer6_outputs(1256) <= a or b;
    layer6_outputs(1257) <= a xor b;
    layer6_outputs(1258) <= a or b;
    layer6_outputs(1259) <= 1'b0;
    layer6_outputs(1260) <= a and b;
    layer6_outputs(1261) <= b;
    layer6_outputs(1262) <= b and not a;
    layer6_outputs(1263) <= not (a or b);
    layer6_outputs(1264) <= not (a and b);
    layer6_outputs(1265) <= b and not a;
    layer6_outputs(1266) <= a and not b;
    layer6_outputs(1267) <= b;
    layer6_outputs(1268) <= a and b;
    layer6_outputs(1269) <= not a;
    layer6_outputs(1270) <= a xor b;
    layer6_outputs(1271) <= not b or a;
    layer6_outputs(1272) <= not (a or b);
    layer6_outputs(1273) <= a and b;
    layer6_outputs(1274) <= not a;
    layer6_outputs(1275) <= not (a and b);
    layer6_outputs(1276) <= a and not b;
    layer6_outputs(1277) <= not a;
    layer6_outputs(1278) <= a xor b;
    layer6_outputs(1279) <= b and not a;
    layer6_outputs(1280) <= not b;
    layer6_outputs(1281) <= not (a or b);
    layer6_outputs(1282) <= not b;
    layer6_outputs(1283) <= not (a or b);
    layer6_outputs(1284) <= not a or b;
    layer6_outputs(1285) <= not a;
    layer6_outputs(1286) <= b and not a;
    layer6_outputs(1287) <= a xor b;
    layer6_outputs(1288) <= a or b;
    layer6_outputs(1289) <= a or b;
    layer6_outputs(1290) <= a and not b;
    layer6_outputs(1291) <= a;
    layer6_outputs(1292) <= a;
    layer6_outputs(1293) <= not (a xor b);
    layer6_outputs(1294) <= not (a and b);
    layer6_outputs(1295) <= b and not a;
    layer6_outputs(1296) <= not b or a;
    layer6_outputs(1297) <= not (a or b);
    layer6_outputs(1298) <= not b or a;
    layer6_outputs(1299) <= not (a xor b);
    layer6_outputs(1300) <= 1'b1;
    layer6_outputs(1301) <= a and b;
    layer6_outputs(1302) <= not (a or b);
    layer6_outputs(1303) <= not (a xor b);
    layer6_outputs(1304) <= a and b;
    layer6_outputs(1305) <= a;
    layer6_outputs(1306) <= a or b;
    layer6_outputs(1307) <= not (a and b);
    layer6_outputs(1308) <= not a or b;
    layer6_outputs(1309) <= not (a or b);
    layer6_outputs(1310) <= not b;
    layer6_outputs(1311) <= b;
    layer6_outputs(1312) <= not b or a;
    layer6_outputs(1313) <= not b;
    layer6_outputs(1314) <= not b;
    layer6_outputs(1315) <= a;
    layer6_outputs(1316) <= a;
    layer6_outputs(1317) <= not a;
    layer6_outputs(1318) <= a;
    layer6_outputs(1319) <= not a;
    layer6_outputs(1320) <= b;
    layer6_outputs(1321) <= a;
    layer6_outputs(1322) <= a;
    layer6_outputs(1323) <= b;
    layer6_outputs(1324) <= not (a xor b);
    layer6_outputs(1325) <= a and not b;
    layer6_outputs(1326) <= a;
    layer6_outputs(1327) <= a and not b;
    layer6_outputs(1328) <= a xor b;
    layer6_outputs(1329) <= b and not a;
    layer6_outputs(1330) <= a and not b;
    layer6_outputs(1331) <= b;
    layer6_outputs(1332) <= not (a or b);
    layer6_outputs(1333) <= a and b;
    layer6_outputs(1334) <= 1'b1;
    layer6_outputs(1335) <= b and not a;
    layer6_outputs(1336) <= not b;
    layer6_outputs(1337) <= not b or a;
    layer6_outputs(1338) <= 1'b0;
    layer6_outputs(1339) <= b;
    layer6_outputs(1340) <= a and not b;
    layer6_outputs(1341) <= a;
    layer6_outputs(1342) <= a or b;
    layer6_outputs(1343) <= not b;
    layer6_outputs(1344) <= not (a or b);
    layer6_outputs(1345) <= not a;
    layer6_outputs(1346) <= not (a or b);
    layer6_outputs(1347) <= not a;
    layer6_outputs(1348) <= b;
    layer6_outputs(1349) <= b and not a;
    layer6_outputs(1350) <= not a;
    layer6_outputs(1351) <= a xor b;
    layer6_outputs(1352) <= b and not a;
    layer6_outputs(1353) <= not a;
    layer6_outputs(1354) <= not b;
    layer6_outputs(1355) <= a;
    layer6_outputs(1356) <= b and not a;
    layer6_outputs(1357) <= a;
    layer6_outputs(1358) <= not (a and b);
    layer6_outputs(1359) <= not b or a;
    layer6_outputs(1360) <= b;
    layer6_outputs(1361) <= not a or b;
    layer6_outputs(1362) <= b and not a;
    layer6_outputs(1363) <= b and not a;
    layer6_outputs(1364) <= b;
    layer6_outputs(1365) <= a or b;
    layer6_outputs(1366) <= a xor b;
    layer6_outputs(1367) <= not (a or b);
    layer6_outputs(1368) <= not a or b;
    layer6_outputs(1369) <= a and not b;
    layer6_outputs(1370) <= 1'b1;
    layer6_outputs(1371) <= not (a or b);
    layer6_outputs(1372) <= 1'b0;
    layer6_outputs(1373) <= a and b;
    layer6_outputs(1374) <= a and not b;
    layer6_outputs(1375) <= a;
    layer6_outputs(1376) <= not a;
    layer6_outputs(1377) <= b;
    layer6_outputs(1378) <= a;
    layer6_outputs(1379) <= not b or a;
    layer6_outputs(1380) <= not (a xor b);
    layer6_outputs(1381) <= not a;
    layer6_outputs(1382) <= not (a and b);
    layer6_outputs(1383) <= not b or a;
    layer6_outputs(1384) <= not (a and b);
    layer6_outputs(1385) <= b and not a;
    layer6_outputs(1386) <= b and not a;
    layer6_outputs(1387) <= a and not b;
    layer6_outputs(1388) <= not a;
    layer6_outputs(1389) <= a;
    layer6_outputs(1390) <= 1'b1;
    layer6_outputs(1391) <= not b;
    layer6_outputs(1392) <= a;
    layer6_outputs(1393) <= not (a and b);
    layer6_outputs(1394) <= b;
    layer6_outputs(1395) <= not (a or b);
    layer6_outputs(1396) <= b;
    layer6_outputs(1397) <= b;
    layer6_outputs(1398) <= a;
    layer6_outputs(1399) <= a and b;
    layer6_outputs(1400) <= not a;
    layer6_outputs(1401) <= not a or b;
    layer6_outputs(1402) <= not b or a;
    layer6_outputs(1403) <= not a;
    layer6_outputs(1404) <= a and not b;
    layer6_outputs(1405) <= not b;
    layer6_outputs(1406) <= not (a and b);
    layer6_outputs(1407) <= not (a xor b);
    layer6_outputs(1408) <= not (a xor b);
    layer6_outputs(1409) <= not (a and b);
    layer6_outputs(1410) <= a;
    layer6_outputs(1411) <= not (a xor b);
    layer6_outputs(1412) <= not a;
    layer6_outputs(1413) <= not a;
    layer6_outputs(1414) <= not (a or b);
    layer6_outputs(1415) <= a and not b;
    layer6_outputs(1416) <= a or b;
    layer6_outputs(1417) <= not a;
    layer6_outputs(1418) <= a and b;
    layer6_outputs(1419) <= not a;
    layer6_outputs(1420) <= not (a and b);
    layer6_outputs(1421) <= not (a or b);
    layer6_outputs(1422) <= a and not b;
    layer6_outputs(1423) <= not b or a;
    layer6_outputs(1424) <= not b;
    layer6_outputs(1425) <= not b or a;
    layer6_outputs(1426) <= a or b;
    layer6_outputs(1427) <= not a;
    layer6_outputs(1428) <= 1'b0;
    layer6_outputs(1429) <= a;
    layer6_outputs(1430) <= not a or b;
    layer6_outputs(1431) <= a;
    layer6_outputs(1432) <= not (a and b);
    layer6_outputs(1433) <= a or b;
    layer6_outputs(1434) <= not (a xor b);
    layer6_outputs(1435) <= not b or a;
    layer6_outputs(1436) <= b and not a;
    layer6_outputs(1437) <= a;
    layer6_outputs(1438) <= not (a or b);
    layer6_outputs(1439) <= a or b;
    layer6_outputs(1440) <= not (a and b);
    layer6_outputs(1441) <= a;
    layer6_outputs(1442) <= not (a and b);
    layer6_outputs(1443) <= b;
    layer6_outputs(1444) <= a or b;
    layer6_outputs(1445) <= b;
    layer6_outputs(1446) <= not b;
    layer6_outputs(1447) <= a;
    layer6_outputs(1448) <= 1'b0;
    layer6_outputs(1449) <= a and b;
    layer6_outputs(1450) <= not a;
    layer6_outputs(1451) <= a or b;
    layer6_outputs(1452) <= not a;
    layer6_outputs(1453) <= not (a and b);
    layer6_outputs(1454) <= not b or a;
    layer6_outputs(1455) <= a;
    layer6_outputs(1456) <= not a;
    layer6_outputs(1457) <= a and b;
    layer6_outputs(1458) <= not (a or b);
    layer6_outputs(1459) <= not b;
    layer6_outputs(1460) <= not (a xor b);
    layer6_outputs(1461) <= b and not a;
    layer6_outputs(1462) <= not a or b;
    layer6_outputs(1463) <= a;
    layer6_outputs(1464) <= 1'b0;
    layer6_outputs(1465) <= b and not a;
    layer6_outputs(1466) <= b;
    layer6_outputs(1467) <= a;
    layer6_outputs(1468) <= a;
    layer6_outputs(1469) <= a or b;
    layer6_outputs(1470) <= not a or b;
    layer6_outputs(1471) <= not a or b;
    layer6_outputs(1472) <= not a or b;
    layer6_outputs(1473) <= a;
    layer6_outputs(1474) <= b and not a;
    layer6_outputs(1475) <= b;
    layer6_outputs(1476) <= not (a and b);
    layer6_outputs(1477) <= b;
    layer6_outputs(1478) <= 1'b1;
    layer6_outputs(1479) <= 1'b1;
    layer6_outputs(1480) <= not a;
    layer6_outputs(1481) <= not (a or b);
    layer6_outputs(1482) <= a xor b;
    layer6_outputs(1483) <= a xor b;
    layer6_outputs(1484) <= a;
    layer6_outputs(1485) <= 1'b0;
    layer6_outputs(1486) <= 1'b1;
    layer6_outputs(1487) <= not a;
    layer6_outputs(1488) <= not b;
    layer6_outputs(1489) <= not (a and b);
    layer6_outputs(1490) <= a or b;
    layer6_outputs(1491) <= a or b;
    layer6_outputs(1492) <= a;
    layer6_outputs(1493) <= a or b;
    layer6_outputs(1494) <= b;
    layer6_outputs(1495) <= not a;
    layer6_outputs(1496) <= b;
    layer6_outputs(1497) <= not a or b;
    layer6_outputs(1498) <= b;
    layer6_outputs(1499) <= not (a or b);
    layer6_outputs(1500) <= a xor b;
    layer6_outputs(1501) <= a or b;
    layer6_outputs(1502) <= a;
    layer6_outputs(1503) <= not (a and b);
    layer6_outputs(1504) <= not b;
    layer6_outputs(1505) <= not (a and b);
    layer6_outputs(1506) <= a;
    layer6_outputs(1507) <= not (a or b);
    layer6_outputs(1508) <= not a;
    layer6_outputs(1509) <= a;
    layer6_outputs(1510) <= a or b;
    layer6_outputs(1511) <= b and not a;
    layer6_outputs(1512) <= a;
    layer6_outputs(1513) <= not (a or b);
    layer6_outputs(1514) <= a or b;
    layer6_outputs(1515) <= not (a or b);
    layer6_outputs(1516) <= b;
    layer6_outputs(1517) <= not (a and b);
    layer6_outputs(1518) <= not (a or b);
    layer6_outputs(1519) <= b;
    layer6_outputs(1520) <= b;
    layer6_outputs(1521) <= a xor b;
    layer6_outputs(1522) <= not (a or b);
    layer6_outputs(1523) <= a;
    layer6_outputs(1524) <= b and not a;
    layer6_outputs(1525) <= not (a xor b);
    layer6_outputs(1526) <= a;
    layer6_outputs(1527) <= not (a or b);
    layer6_outputs(1528) <= a and b;
    layer6_outputs(1529) <= not b;
    layer6_outputs(1530) <= not a;
    layer6_outputs(1531) <= not a;
    layer6_outputs(1532) <= b;
    layer6_outputs(1533) <= a and not b;
    layer6_outputs(1534) <= not (a and b);
    layer6_outputs(1535) <= b;
    layer6_outputs(1536) <= not (a or b);
    layer6_outputs(1537) <= a and not b;
    layer6_outputs(1538) <= a and not b;
    layer6_outputs(1539) <= not b or a;
    layer6_outputs(1540) <= a;
    layer6_outputs(1541) <= not a;
    layer6_outputs(1542) <= a and not b;
    layer6_outputs(1543) <= b;
    layer6_outputs(1544) <= not (a or b);
    layer6_outputs(1545) <= a and b;
    layer6_outputs(1546) <= not (a xor b);
    layer6_outputs(1547) <= a;
    layer6_outputs(1548) <= a or b;
    layer6_outputs(1549) <= b;
    layer6_outputs(1550) <= a or b;
    layer6_outputs(1551) <= a or b;
    layer6_outputs(1552) <= 1'b0;
    layer6_outputs(1553) <= not a;
    layer6_outputs(1554) <= not a or b;
    layer6_outputs(1555) <= a and b;
    layer6_outputs(1556) <= not (a xor b);
    layer6_outputs(1557) <= a and b;
    layer6_outputs(1558) <= not (a or b);
    layer6_outputs(1559) <= a or b;
    layer6_outputs(1560) <= not (a and b);
    layer6_outputs(1561) <= not (a and b);
    layer6_outputs(1562) <= b and not a;
    layer6_outputs(1563) <= not b or a;
    layer6_outputs(1564) <= b and not a;
    layer6_outputs(1565) <= not a;
    layer6_outputs(1566) <= a and not b;
    layer6_outputs(1567) <= not (a xor b);
    layer6_outputs(1568) <= b;
    layer6_outputs(1569) <= b;
    layer6_outputs(1570) <= not a;
    layer6_outputs(1571) <= not b or a;
    layer6_outputs(1572) <= not (a and b);
    layer6_outputs(1573) <= not b or a;
    layer6_outputs(1574) <= b;
    layer6_outputs(1575) <= not (a or b);
    layer6_outputs(1576) <= not (a or b);
    layer6_outputs(1577) <= b;
    layer6_outputs(1578) <= not (a or b);
    layer6_outputs(1579) <= a or b;
    layer6_outputs(1580) <= 1'b1;
    layer6_outputs(1581) <= a and not b;
    layer6_outputs(1582) <= b;
    layer6_outputs(1583) <= not (a xor b);
    layer6_outputs(1584) <= a;
    layer6_outputs(1585) <= 1'b0;
    layer6_outputs(1586) <= b and not a;
    layer6_outputs(1587) <= not b or a;
    layer6_outputs(1588) <= a and not b;
    layer6_outputs(1589) <= not (a or b);
    layer6_outputs(1590) <= not b or a;
    layer6_outputs(1591) <= 1'b0;
    layer6_outputs(1592) <= a or b;
    layer6_outputs(1593) <= not b;
    layer6_outputs(1594) <= a and not b;
    layer6_outputs(1595) <= a xor b;
    layer6_outputs(1596) <= a and not b;
    layer6_outputs(1597) <= not b;
    layer6_outputs(1598) <= a and not b;
    layer6_outputs(1599) <= a;
    layer6_outputs(1600) <= a;
    layer6_outputs(1601) <= a;
    layer6_outputs(1602) <= 1'b0;
    layer6_outputs(1603) <= a and b;
    layer6_outputs(1604) <= b and not a;
    layer6_outputs(1605) <= a and b;
    layer6_outputs(1606) <= a xor b;
    layer6_outputs(1607) <= a;
    layer6_outputs(1608) <= not (a and b);
    layer6_outputs(1609) <= not (a xor b);
    layer6_outputs(1610) <= not b;
    layer6_outputs(1611) <= not a;
    layer6_outputs(1612) <= a xor b;
    layer6_outputs(1613) <= 1'b0;
    layer6_outputs(1614) <= a and not b;
    layer6_outputs(1615) <= 1'b0;
    layer6_outputs(1616) <= b;
    layer6_outputs(1617) <= not b;
    layer6_outputs(1618) <= not b or a;
    layer6_outputs(1619) <= a xor b;
    layer6_outputs(1620) <= b;
    layer6_outputs(1621) <= b and not a;
    layer6_outputs(1622) <= a and b;
    layer6_outputs(1623) <= not a;
    layer6_outputs(1624) <= a and b;
    layer6_outputs(1625) <= not b or a;
    layer6_outputs(1626) <= a and b;
    layer6_outputs(1627) <= a and not b;
    layer6_outputs(1628) <= not (a and b);
    layer6_outputs(1629) <= not (a and b);
    layer6_outputs(1630) <= not (a xor b);
    layer6_outputs(1631) <= not a;
    layer6_outputs(1632) <= a;
    layer6_outputs(1633) <= not (a xor b);
    layer6_outputs(1634) <= b;
    layer6_outputs(1635) <= not a;
    layer6_outputs(1636) <= a xor b;
    layer6_outputs(1637) <= 1'b1;
    layer6_outputs(1638) <= b and not a;
    layer6_outputs(1639) <= a;
    layer6_outputs(1640) <= not a;
    layer6_outputs(1641) <= a or b;
    layer6_outputs(1642) <= a and not b;
    layer6_outputs(1643) <= not (a or b);
    layer6_outputs(1644) <= not b;
    layer6_outputs(1645) <= not (a or b);
    layer6_outputs(1646) <= not a or b;
    layer6_outputs(1647) <= not b;
    layer6_outputs(1648) <= not b;
    layer6_outputs(1649) <= not b;
    layer6_outputs(1650) <= a and not b;
    layer6_outputs(1651) <= not b or a;
    layer6_outputs(1652) <= not a;
    layer6_outputs(1653) <= not b or a;
    layer6_outputs(1654) <= a or b;
    layer6_outputs(1655) <= a;
    layer6_outputs(1656) <= a;
    layer6_outputs(1657) <= a or b;
    layer6_outputs(1658) <= a or b;
    layer6_outputs(1659) <= a and not b;
    layer6_outputs(1660) <= a xor b;
    layer6_outputs(1661) <= not (a or b);
    layer6_outputs(1662) <= a or b;
    layer6_outputs(1663) <= not (a and b);
    layer6_outputs(1664) <= not b or a;
    layer6_outputs(1665) <= a;
    layer6_outputs(1666) <= b;
    layer6_outputs(1667) <= b;
    layer6_outputs(1668) <= b;
    layer6_outputs(1669) <= a or b;
    layer6_outputs(1670) <= not (a and b);
    layer6_outputs(1671) <= a;
    layer6_outputs(1672) <= a and b;
    layer6_outputs(1673) <= a;
    layer6_outputs(1674) <= not b;
    layer6_outputs(1675) <= a and not b;
    layer6_outputs(1676) <= not a;
    layer6_outputs(1677) <= a;
    layer6_outputs(1678) <= a or b;
    layer6_outputs(1679) <= not a;
    layer6_outputs(1680) <= not a or b;
    layer6_outputs(1681) <= not b;
    layer6_outputs(1682) <= a and not b;
    layer6_outputs(1683) <= not a or b;
    layer6_outputs(1684) <= not a;
    layer6_outputs(1685) <= not b or a;
    layer6_outputs(1686) <= b;
    layer6_outputs(1687) <= not a;
    layer6_outputs(1688) <= not b;
    layer6_outputs(1689) <= not (a or b);
    layer6_outputs(1690) <= not (a and b);
    layer6_outputs(1691) <= not b;
    layer6_outputs(1692) <= not b or a;
    layer6_outputs(1693) <= b;
    layer6_outputs(1694) <= not a;
    layer6_outputs(1695) <= b;
    layer6_outputs(1696) <= not (a or b);
    layer6_outputs(1697) <= not a;
    layer6_outputs(1698) <= a xor b;
    layer6_outputs(1699) <= a or b;
    layer6_outputs(1700) <= not a;
    layer6_outputs(1701) <= a;
    layer6_outputs(1702) <= a or b;
    layer6_outputs(1703) <= not b;
    layer6_outputs(1704) <= b;
    layer6_outputs(1705) <= not b;
    layer6_outputs(1706) <= not b;
    layer6_outputs(1707) <= a xor b;
    layer6_outputs(1708) <= not (a or b);
    layer6_outputs(1709) <= not b;
    layer6_outputs(1710) <= not b;
    layer6_outputs(1711) <= not (a and b);
    layer6_outputs(1712) <= a and b;
    layer6_outputs(1713) <= not (a or b);
    layer6_outputs(1714) <= not a;
    layer6_outputs(1715) <= not a;
    layer6_outputs(1716) <= 1'b1;
    layer6_outputs(1717) <= not b or a;
    layer6_outputs(1718) <= not a;
    layer6_outputs(1719) <= b;
    layer6_outputs(1720) <= not a;
    layer6_outputs(1721) <= a and not b;
    layer6_outputs(1722) <= not b;
    layer6_outputs(1723) <= not (a or b);
    layer6_outputs(1724) <= a;
    layer6_outputs(1725) <= a or b;
    layer6_outputs(1726) <= b;
    layer6_outputs(1727) <= a and not b;
    layer6_outputs(1728) <= not (a and b);
    layer6_outputs(1729) <= not a;
    layer6_outputs(1730) <= b;
    layer6_outputs(1731) <= b and not a;
    layer6_outputs(1732) <= not a;
    layer6_outputs(1733) <= 1'b1;
    layer6_outputs(1734) <= b;
    layer6_outputs(1735) <= not a;
    layer6_outputs(1736) <= not b or a;
    layer6_outputs(1737) <= not a;
    layer6_outputs(1738) <= b;
    layer6_outputs(1739) <= not a;
    layer6_outputs(1740) <= not a or b;
    layer6_outputs(1741) <= not (a or b);
    layer6_outputs(1742) <= a xor b;
    layer6_outputs(1743) <= a xor b;
    layer6_outputs(1744) <= b and not a;
    layer6_outputs(1745) <= not a or b;
    layer6_outputs(1746) <= not b or a;
    layer6_outputs(1747) <= 1'b0;
    layer6_outputs(1748) <= b and not a;
    layer6_outputs(1749) <= b and not a;
    layer6_outputs(1750) <= not a;
    layer6_outputs(1751) <= a;
    layer6_outputs(1752) <= a;
    layer6_outputs(1753) <= not a or b;
    layer6_outputs(1754) <= not (a or b);
    layer6_outputs(1755) <= b;
    layer6_outputs(1756) <= a or b;
    layer6_outputs(1757) <= not (a and b);
    layer6_outputs(1758) <= b;
    layer6_outputs(1759) <= not (a or b);
    layer6_outputs(1760) <= a and not b;
    layer6_outputs(1761) <= a;
    layer6_outputs(1762) <= b and not a;
    layer6_outputs(1763) <= not b or a;
    layer6_outputs(1764) <= not (a xor b);
    layer6_outputs(1765) <= b;
    layer6_outputs(1766) <= a;
    layer6_outputs(1767) <= not (a xor b);
    layer6_outputs(1768) <= a or b;
    layer6_outputs(1769) <= b;
    layer6_outputs(1770) <= a and b;
    layer6_outputs(1771) <= a;
    layer6_outputs(1772) <= not a;
    layer6_outputs(1773) <= not a or b;
    layer6_outputs(1774) <= a xor b;
    layer6_outputs(1775) <= not b;
    layer6_outputs(1776) <= b;
    layer6_outputs(1777) <= b;
    layer6_outputs(1778) <= a and b;
    layer6_outputs(1779) <= not (a and b);
    layer6_outputs(1780) <= a and b;
    layer6_outputs(1781) <= a and b;
    layer6_outputs(1782) <= not (a and b);
    layer6_outputs(1783) <= a and b;
    layer6_outputs(1784) <= not a;
    layer6_outputs(1785) <= not b;
    layer6_outputs(1786) <= a;
    layer6_outputs(1787) <= b;
    layer6_outputs(1788) <= not b;
    layer6_outputs(1789) <= a;
    layer6_outputs(1790) <= not a;
    layer6_outputs(1791) <= not b;
    layer6_outputs(1792) <= not b or a;
    layer6_outputs(1793) <= b;
    layer6_outputs(1794) <= b and not a;
    layer6_outputs(1795) <= b;
    layer6_outputs(1796) <= not b;
    layer6_outputs(1797) <= a and not b;
    layer6_outputs(1798) <= b;
    layer6_outputs(1799) <= a or b;
    layer6_outputs(1800) <= b;
    layer6_outputs(1801) <= b and not a;
    layer6_outputs(1802) <= not a;
    layer6_outputs(1803) <= a and not b;
    layer6_outputs(1804) <= a and b;
    layer6_outputs(1805) <= a or b;
    layer6_outputs(1806) <= not a or b;
    layer6_outputs(1807) <= b;
    layer6_outputs(1808) <= a and b;
    layer6_outputs(1809) <= not a or b;
    layer6_outputs(1810) <= not b;
    layer6_outputs(1811) <= 1'b1;
    layer6_outputs(1812) <= a;
    layer6_outputs(1813) <= not a or b;
    layer6_outputs(1814) <= a;
    layer6_outputs(1815) <= not (a or b);
    layer6_outputs(1816) <= a and not b;
    layer6_outputs(1817) <= not a;
    layer6_outputs(1818) <= b;
    layer6_outputs(1819) <= a;
    layer6_outputs(1820) <= not (a xor b);
    layer6_outputs(1821) <= not b;
    layer6_outputs(1822) <= b and not a;
    layer6_outputs(1823) <= a and b;
    layer6_outputs(1824) <= a;
    layer6_outputs(1825) <= not (a xor b);
    layer6_outputs(1826) <= b and not a;
    layer6_outputs(1827) <= b;
    layer6_outputs(1828) <= a xor b;
    layer6_outputs(1829) <= not (a xor b);
    layer6_outputs(1830) <= not a;
    layer6_outputs(1831) <= not a or b;
    layer6_outputs(1832) <= 1'b1;
    layer6_outputs(1833) <= not b;
    layer6_outputs(1834) <= a and not b;
    layer6_outputs(1835) <= not (a and b);
    layer6_outputs(1836) <= a and b;
    layer6_outputs(1837) <= a xor b;
    layer6_outputs(1838) <= a;
    layer6_outputs(1839) <= not a;
    layer6_outputs(1840) <= not a or b;
    layer6_outputs(1841) <= not b;
    layer6_outputs(1842) <= a and b;
    layer6_outputs(1843) <= a and not b;
    layer6_outputs(1844) <= not b;
    layer6_outputs(1845) <= b and not a;
    layer6_outputs(1846) <= a and b;
    layer6_outputs(1847) <= not b or a;
    layer6_outputs(1848) <= a or b;
    layer6_outputs(1849) <= b;
    layer6_outputs(1850) <= not (a and b);
    layer6_outputs(1851) <= a or b;
    layer6_outputs(1852) <= a or b;
    layer6_outputs(1853) <= not a;
    layer6_outputs(1854) <= a and b;
    layer6_outputs(1855) <= a and not b;
    layer6_outputs(1856) <= not (a or b);
    layer6_outputs(1857) <= a or b;
    layer6_outputs(1858) <= a and not b;
    layer6_outputs(1859) <= not b;
    layer6_outputs(1860) <= not (a or b);
    layer6_outputs(1861) <= not (a and b);
    layer6_outputs(1862) <= a or b;
    layer6_outputs(1863) <= not b;
    layer6_outputs(1864) <= not b;
    layer6_outputs(1865) <= b;
    layer6_outputs(1866) <= not (a or b);
    layer6_outputs(1867) <= not (a or b);
    layer6_outputs(1868) <= not a or b;
    layer6_outputs(1869) <= not a;
    layer6_outputs(1870) <= b and not a;
    layer6_outputs(1871) <= 1'b0;
    layer6_outputs(1872) <= not a;
    layer6_outputs(1873) <= a and not b;
    layer6_outputs(1874) <= b;
    layer6_outputs(1875) <= not b;
    layer6_outputs(1876) <= not b or a;
    layer6_outputs(1877) <= a;
    layer6_outputs(1878) <= b;
    layer6_outputs(1879) <= not b;
    layer6_outputs(1880) <= b;
    layer6_outputs(1881) <= not (a or b);
    layer6_outputs(1882) <= b;
    layer6_outputs(1883) <= b;
    layer6_outputs(1884) <= 1'b1;
    layer6_outputs(1885) <= not b;
    layer6_outputs(1886) <= not b or a;
    layer6_outputs(1887) <= not (a or b);
    layer6_outputs(1888) <= b;
    layer6_outputs(1889) <= b;
    layer6_outputs(1890) <= a;
    layer6_outputs(1891) <= not b or a;
    layer6_outputs(1892) <= a and not b;
    layer6_outputs(1893) <= not b or a;
    layer6_outputs(1894) <= not a or b;
    layer6_outputs(1895) <= not a or b;
    layer6_outputs(1896) <= not (a and b);
    layer6_outputs(1897) <= a or b;
    layer6_outputs(1898) <= b and not a;
    layer6_outputs(1899) <= b;
    layer6_outputs(1900) <= b;
    layer6_outputs(1901) <= b;
    layer6_outputs(1902) <= b and not a;
    layer6_outputs(1903) <= a and not b;
    layer6_outputs(1904) <= b;
    layer6_outputs(1905) <= a;
    layer6_outputs(1906) <= a or b;
    layer6_outputs(1907) <= not (a xor b);
    layer6_outputs(1908) <= not (a xor b);
    layer6_outputs(1909) <= b and not a;
    layer6_outputs(1910) <= not (a or b);
    layer6_outputs(1911) <= 1'b0;
    layer6_outputs(1912) <= b and not a;
    layer6_outputs(1913) <= not (a or b);
    layer6_outputs(1914) <= not a or b;
    layer6_outputs(1915) <= a and b;
    layer6_outputs(1916) <= not b;
    layer6_outputs(1917) <= not (a and b);
    layer6_outputs(1918) <= b and not a;
    layer6_outputs(1919) <= a and b;
    layer6_outputs(1920) <= b;
    layer6_outputs(1921) <= not a;
    layer6_outputs(1922) <= not b;
    layer6_outputs(1923) <= a and not b;
    layer6_outputs(1924) <= not b;
    layer6_outputs(1925) <= b;
    layer6_outputs(1926) <= a;
    layer6_outputs(1927) <= not b;
    layer6_outputs(1928) <= a;
    layer6_outputs(1929) <= a and not b;
    layer6_outputs(1930) <= not a or b;
    layer6_outputs(1931) <= b and not a;
    layer6_outputs(1932) <= not (a or b);
    layer6_outputs(1933) <= a and not b;
    layer6_outputs(1934) <= a;
    layer6_outputs(1935) <= a and b;
    layer6_outputs(1936) <= 1'b1;
    layer6_outputs(1937) <= a xor b;
    layer6_outputs(1938) <= not a or b;
    layer6_outputs(1939) <= not b or a;
    layer6_outputs(1940) <= not a;
    layer6_outputs(1941) <= b;
    layer6_outputs(1942) <= not b or a;
    layer6_outputs(1943) <= b;
    layer6_outputs(1944) <= not a or b;
    layer6_outputs(1945) <= not b;
    layer6_outputs(1946) <= a;
    layer6_outputs(1947) <= a;
    layer6_outputs(1948) <= not a;
    layer6_outputs(1949) <= not (a and b);
    layer6_outputs(1950) <= a and not b;
    layer6_outputs(1951) <= a and not b;
    layer6_outputs(1952) <= not (a or b);
    layer6_outputs(1953) <= b;
    layer6_outputs(1954) <= a;
    layer6_outputs(1955) <= a;
    layer6_outputs(1956) <= b;
    layer6_outputs(1957) <= a and b;
    layer6_outputs(1958) <= not a;
    layer6_outputs(1959) <= not (a and b);
    layer6_outputs(1960) <= not a or b;
    layer6_outputs(1961) <= a and not b;
    layer6_outputs(1962) <= a xor b;
    layer6_outputs(1963) <= not a or b;
    layer6_outputs(1964) <= a or b;
    layer6_outputs(1965) <= not (a or b);
    layer6_outputs(1966) <= a;
    layer6_outputs(1967) <= not b;
    layer6_outputs(1968) <= not (a or b);
    layer6_outputs(1969) <= a;
    layer6_outputs(1970) <= not b;
    layer6_outputs(1971) <= a and not b;
    layer6_outputs(1972) <= a xor b;
    layer6_outputs(1973) <= a and not b;
    layer6_outputs(1974) <= b;
    layer6_outputs(1975) <= not a;
    layer6_outputs(1976) <= not b;
    layer6_outputs(1977) <= a xor b;
    layer6_outputs(1978) <= not (a or b);
    layer6_outputs(1979) <= not b or a;
    layer6_outputs(1980) <= not (a and b);
    layer6_outputs(1981) <= a or b;
    layer6_outputs(1982) <= not b;
    layer6_outputs(1983) <= a and not b;
    layer6_outputs(1984) <= a and not b;
    layer6_outputs(1985) <= 1'b1;
    layer6_outputs(1986) <= b;
    layer6_outputs(1987) <= a or b;
    layer6_outputs(1988) <= not (a xor b);
    layer6_outputs(1989) <= a and not b;
    layer6_outputs(1990) <= not a;
    layer6_outputs(1991) <= a or b;
    layer6_outputs(1992) <= a or b;
    layer6_outputs(1993) <= not b;
    layer6_outputs(1994) <= not (a and b);
    layer6_outputs(1995) <= a or b;
    layer6_outputs(1996) <= not (a or b);
    layer6_outputs(1997) <= b and not a;
    layer6_outputs(1998) <= not b;
    layer6_outputs(1999) <= a and not b;
    layer6_outputs(2000) <= a and not b;
    layer6_outputs(2001) <= a and b;
    layer6_outputs(2002) <= a or b;
    layer6_outputs(2003) <= a or b;
    layer6_outputs(2004) <= not a;
    layer6_outputs(2005) <= b and not a;
    layer6_outputs(2006) <= b;
    layer6_outputs(2007) <= a or b;
    layer6_outputs(2008) <= not (a xor b);
    layer6_outputs(2009) <= 1'b0;
    layer6_outputs(2010) <= not (a and b);
    layer6_outputs(2011) <= not (a or b);
    layer6_outputs(2012) <= a and not b;
    layer6_outputs(2013) <= not b;
    layer6_outputs(2014) <= a xor b;
    layer6_outputs(2015) <= not (a xor b);
    layer6_outputs(2016) <= a xor b;
    layer6_outputs(2017) <= a;
    layer6_outputs(2018) <= a and b;
    layer6_outputs(2019) <= a;
    layer6_outputs(2020) <= a;
    layer6_outputs(2021) <= a;
    layer6_outputs(2022) <= not a;
    layer6_outputs(2023) <= a;
    layer6_outputs(2024) <= not b;
    layer6_outputs(2025) <= not a;
    layer6_outputs(2026) <= not (a or b);
    layer6_outputs(2027) <= not b;
    layer6_outputs(2028) <= a and b;
    layer6_outputs(2029) <= not a or b;
    layer6_outputs(2030) <= a and not b;
    layer6_outputs(2031) <= a or b;
    layer6_outputs(2032) <= b;
    layer6_outputs(2033) <= b;
    layer6_outputs(2034) <= a;
    layer6_outputs(2035) <= not a;
    layer6_outputs(2036) <= not (a xor b);
    layer6_outputs(2037) <= not a;
    layer6_outputs(2038) <= not a;
    layer6_outputs(2039) <= not b or a;
    layer6_outputs(2040) <= not b;
    layer6_outputs(2041) <= a;
    layer6_outputs(2042) <= a and b;
    layer6_outputs(2043) <= not b or a;
    layer6_outputs(2044) <= not b;
    layer6_outputs(2045) <= a;
    layer6_outputs(2046) <= a;
    layer6_outputs(2047) <= not (a xor b);
    layer6_outputs(2048) <= b;
    layer6_outputs(2049) <= not a;
    layer6_outputs(2050) <= not a or b;
    layer6_outputs(2051) <= 1'b1;
    layer6_outputs(2052) <= b;
    layer6_outputs(2053) <= a;
    layer6_outputs(2054) <= a or b;
    layer6_outputs(2055) <= not b;
    layer6_outputs(2056) <= a;
    layer6_outputs(2057) <= b and not a;
    layer6_outputs(2058) <= not a;
    layer6_outputs(2059) <= b;
    layer6_outputs(2060) <= a;
    layer6_outputs(2061) <= b;
    layer6_outputs(2062) <= not (a or b);
    layer6_outputs(2063) <= not a;
    layer6_outputs(2064) <= not a or b;
    layer6_outputs(2065) <= 1'b0;
    layer6_outputs(2066) <= not (a xor b);
    layer6_outputs(2067) <= not b or a;
    layer6_outputs(2068) <= not b;
    layer6_outputs(2069) <= b and not a;
    layer6_outputs(2070) <= not (a and b);
    layer6_outputs(2071) <= not b;
    layer6_outputs(2072) <= 1'b0;
    layer6_outputs(2073) <= not a;
    layer6_outputs(2074) <= a;
    layer6_outputs(2075) <= not a or b;
    layer6_outputs(2076) <= not a;
    layer6_outputs(2077) <= b;
    layer6_outputs(2078) <= b;
    layer6_outputs(2079) <= b;
    layer6_outputs(2080) <= not b or a;
    layer6_outputs(2081) <= not b;
    layer6_outputs(2082) <= b;
    layer6_outputs(2083) <= not a;
    layer6_outputs(2084) <= not (a or b);
    layer6_outputs(2085) <= a or b;
    layer6_outputs(2086) <= not (a and b);
    layer6_outputs(2087) <= not a or b;
    layer6_outputs(2088) <= a xor b;
    layer6_outputs(2089) <= not b or a;
    layer6_outputs(2090) <= a;
    layer6_outputs(2091) <= not a;
    layer6_outputs(2092) <= a;
    layer6_outputs(2093) <= a or b;
    layer6_outputs(2094) <= a xor b;
    layer6_outputs(2095) <= not (a and b);
    layer6_outputs(2096) <= b;
    layer6_outputs(2097) <= not a or b;
    layer6_outputs(2098) <= not a;
    layer6_outputs(2099) <= a and b;
    layer6_outputs(2100) <= a or b;
    layer6_outputs(2101) <= not (a xor b);
    layer6_outputs(2102) <= not b or a;
    layer6_outputs(2103) <= a;
    layer6_outputs(2104) <= a and b;
    layer6_outputs(2105) <= b and not a;
    layer6_outputs(2106) <= b;
    layer6_outputs(2107) <= not a;
    layer6_outputs(2108) <= b;
    layer6_outputs(2109) <= a and b;
    layer6_outputs(2110) <= a;
    layer6_outputs(2111) <= 1'b0;
    layer6_outputs(2112) <= not b;
    layer6_outputs(2113) <= not (a or b);
    layer6_outputs(2114) <= not b;
    layer6_outputs(2115) <= b;
    layer6_outputs(2116) <= a or b;
    layer6_outputs(2117) <= not (a and b);
    layer6_outputs(2118) <= a;
    layer6_outputs(2119) <= b;
    layer6_outputs(2120) <= not (a xor b);
    layer6_outputs(2121) <= not (a and b);
    layer6_outputs(2122) <= b;
    layer6_outputs(2123) <= not b;
    layer6_outputs(2124) <= a and b;
    layer6_outputs(2125) <= b and not a;
    layer6_outputs(2126) <= b;
    layer6_outputs(2127) <= a;
    layer6_outputs(2128) <= b;
    layer6_outputs(2129) <= a and not b;
    layer6_outputs(2130) <= not a;
    layer6_outputs(2131) <= b;
    layer6_outputs(2132) <= a;
    layer6_outputs(2133) <= not b;
    layer6_outputs(2134) <= not a or b;
    layer6_outputs(2135) <= not (a xor b);
    layer6_outputs(2136) <= not b;
    layer6_outputs(2137) <= a or b;
    layer6_outputs(2138) <= not (a or b);
    layer6_outputs(2139) <= b and not a;
    layer6_outputs(2140) <= not a;
    layer6_outputs(2141) <= 1'b1;
    layer6_outputs(2142) <= not b or a;
    layer6_outputs(2143) <= a and not b;
    layer6_outputs(2144) <= b and not a;
    layer6_outputs(2145) <= b;
    layer6_outputs(2146) <= b and not a;
    layer6_outputs(2147) <= a or b;
    layer6_outputs(2148) <= a or b;
    layer6_outputs(2149) <= not a;
    layer6_outputs(2150) <= not (a or b);
    layer6_outputs(2151) <= b;
    layer6_outputs(2152) <= not a;
    layer6_outputs(2153) <= not a;
    layer6_outputs(2154) <= not a;
    layer6_outputs(2155) <= not (a and b);
    layer6_outputs(2156) <= a;
    layer6_outputs(2157) <= not a;
    layer6_outputs(2158) <= not (a or b);
    layer6_outputs(2159) <= b and not a;
    layer6_outputs(2160) <= not a;
    layer6_outputs(2161) <= not b or a;
    layer6_outputs(2162) <= a;
    layer6_outputs(2163) <= 1'b0;
    layer6_outputs(2164) <= b;
    layer6_outputs(2165) <= a;
    layer6_outputs(2166) <= not a;
    layer6_outputs(2167) <= b;
    layer6_outputs(2168) <= not (a or b);
    layer6_outputs(2169) <= not a;
    layer6_outputs(2170) <= a and not b;
    layer6_outputs(2171) <= b;
    layer6_outputs(2172) <= 1'b1;
    layer6_outputs(2173) <= not (a and b);
    layer6_outputs(2174) <= a;
    layer6_outputs(2175) <= a;
    layer6_outputs(2176) <= not b;
    layer6_outputs(2177) <= not (a and b);
    layer6_outputs(2178) <= not b or a;
    layer6_outputs(2179) <= 1'b1;
    layer6_outputs(2180) <= not b;
    layer6_outputs(2181) <= a and b;
    layer6_outputs(2182) <= not (a or b);
    layer6_outputs(2183) <= not (a or b);
    layer6_outputs(2184) <= not a;
    layer6_outputs(2185) <= a;
    layer6_outputs(2186) <= b;
    layer6_outputs(2187) <= a and not b;
    layer6_outputs(2188) <= b;
    layer6_outputs(2189) <= not b;
    layer6_outputs(2190) <= a;
    layer6_outputs(2191) <= not b or a;
    layer6_outputs(2192) <= a;
    layer6_outputs(2193) <= not b;
    layer6_outputs(2194) <= a or b;
    layer6_outputs(2195) <= b and not a;
    layer6_outputs(2196) <= not (a xor b);
    layer6_outputs(2197) <= not (a xor b);
    layer6_outputs(2198) <= a or b;
    layer6_outputs(2199) <= not a;
    layer6_outputs(2200) <= a and b;
    layer6_outputs(2201) <= not a;
    layer6_outputs(2202) <= not a;
    layer6_outputs(2203) <= a xor b;
    layer6_outputs(2204) <= not (a and b);
    layer6_outputs(2205) <= b;
    layer6_outputs(2206) <= not a;
    layer6_outputs(2207) <= a;
    layer6_outputs(2208) <= not (a and b);
    layer6_outputs(2209) <= b and not a;
    layer6_outputs(2210) <= a and b;
    layer6_outputs(2211) <= not (a or b);
    layer6_outputs(2212) <= not (a or b);
    layer6_outputs(2213) <= 1'b1;
    layer6_outputs(2214) <= 1'b0;
    layer6_outputs(2215) <= a and not b;
    layer6_outputs(2216) <= not b or a;
    layer6_outputs(2217) <= a xor b;
    layer6_outputs(2218) <= b;
    layer6_outputs(2219) <= b and not a;
    layer6_outputs(2220) <= 1'b0;
    layer6_outputs(2221) <= b;
    layer6_outputs(2222) <= not a or b;
    layer6_outputs(2223) <= not b or a;
    layer6_outputs(2224) <= not a or b;
    layer6_outputs(2225) <= b;
    layer6_outputs(2226) <= not a;
    layer6_outputs(2227) <= not a or b;
    layer6_outputs(2228) <= not b;
    layer6_outputs(2229) <= not (a and b);
    layer6_outputs(2230) <= a xor b;
    layer6_outputs(2231) <= a and b;
    layer6_outputs(2232) <= not (a or b);
    layer6_outputs(2233) <= not (a and b);
    layer6_outputs(2234) <= not b or a;
    layer6_outputs(2235) <= not (a and b);
    layer6_outputs(2236) <= not b or a;
    layer6_outputs(2237) <= a xor b;
    layer6_outputs(2238) <= b;
    layer6_outputs(2239) <= b and not a;
    layer6_outputs(2240) <= not a;
    layer6_outputs(2241) <= b and not a;
    layer6_outputs(2242) <= a;
    layer6_outputs(2243) <= a and not b;
    layer6_outputs(2244) <= not b or a;
    layer6_outputs(2245) <= not b;
    layer6_outputs(2246) <= b;
    layer6_outputs(2247) <= not b or a;
    layer6_outputs(2248) <= a xor b;
    layer6_outputs(2249) <= not b;
    layer6_outputs(2250) <= b and not a;
    layer6_outputs(2251) <= not b;
    layer6_outputs(2252) <= not a or b;
    layer6_outputs(2253) <= not (a or b);
    layer6_outputs(2254) <= a and b;
    layer6_outputs(2255) <= 1'b0;
    layer6_outputs(2256) <= not b;
    layer6_outputs(2257) <= not (a or b);
    layer6_outputs(2258) <= b;
    layer6_outputs(2259) <= not a;
    layer6_outputs(2260) <= b;
    layer6_outputs(2261) <= not b;
    layer6_outputs(2262) <= a and not b;
    layer6_outputs(2263) <= a and not b;
    layer6_outputs(2264) <= not b;
    layer6_outputs(2265) <= a and b;
    layer6_outputs(2266) <= a or b;
    layer6_outputs(2267) <= not b or a;
    layer6_outputs(2268) <= b;
    layer6_outputs(2269) <= a and not b;
    layer6_outputs(2270) <= not a or b;
    layer6_outputs(2271) <= not b;
    layer6_outputs(2272) <= not b;
    layer6_outputs(2273) <= not (a or b);
    layer6_outputs(2274) <= not b;
    layer6_outputs(2275) <= not b;
    layer6_outputs(2276) <= not a;
    layer6_outputs(2277) <= a and not b;
    layer6_outputs(2278) <= b;
    layer6_outputs(2279) <= a and b;
    layer6_outputs(2280) <= not a or b;
    layer6_outputs(2281) <= not (a or b);
    layer6_outputs(2282) <= not (a and b);
    layer6_outputs(2283) <= a or b;
    layer6_outputs(2284) <= not a;
    layer6_outputs(2285) <= not (a xor b);
    layer6_outputs(2286) <= not (a or b);
    layer6_outputs(2287) <= not a;
    layer6_outputs(2288) <= a and b;
    layer6_outputs(2289) <= a and not b;
    layer6_outputs(2290) <= b;
    layer6_outputs(2291) <= a;
    layer6_outputs(2292) <= 1'b0;
    layer6_outputs(2293) <= not a;
    layer6_outputs(2294) <= a and b;
    layer6_outputs(2295) <= not a or b;
    layer6_outputs(2296) <= a and not b;
    layer6_outputs(2297) <= not (a and b);
    layer6_outputs(2298) <= not a;
    layer6_outputs(2299) <= not b or a;
    layer6_outputs(2300) <= a xor b;
    layer6_outputs(2301) <= not a;
    layer6_outputs(2302) <= a;
    layer6_outputs(2303) <= not (a xor b);
    layer6_outputs(2304) <= b;
    layer6_outputs(2305) <= a;
    layer6_outputs(2306) <= a and b;
    layer6_outputs(2307) <= not a or b;
    layer6_outputs(2308) <= b;
    layer6_outputs(2309) <= not a;
    layer6_outputs(2310) <= b and not a;
    layer6_outputs(2311) <= a xor b;
    layer6_outputs(2312) <= not a;
    layer6_outputs(2313) <= not (a xor b);
    layer6_outputs(2314) <= not b or a;
    layer6_outputs(2315) <= not b;
    layer6_outputs(2316) <= not a;
    layer6_outputs(2317) <= not b or a;
    layer6_outputs(2318) <= 1'b0;
    layer6_outputs(2319) <= not (a or b);
    layer6_outputs(2320) <= not b;
    layer6_outputs(2321) <= b;
    layer6_outputs(2322) <= 1'b1;
    layer6_outputs(2323) <= not b;
    layer6_outputs(2324) <= a xor b;
    layer6_outputs(2325) <= not b;
    layer6_outputs(2326) <= not b;
    layer6_outputs(2327) <= b;
    layer6_outputs(2328) <= b and not a;
    layer6_outputs(2329) <= 1'b1;
    layer6_outputs(2330) <= a and not b;
    layer6_outputs(2331) <= a;
    layer6_outputs(2332) <= 1'b1;
    layer6_outputs(2333) <= b;
    layer6_outputs(2334) <= 1'b0;
    layer6_outputs(2335) <= b;
    layer6_outputs(2336) <= b;
    layer6_outputs(2337) <= b and not a;
    layer6_outputs(2338) <= not (a xor b);
    layer6_outputs(2339) <= a;
    layer6_outputs(2340) <= not a or b;
    layer6_outputs(2341) <= a;
    layer6_outputs(2342) <= not b;
    layer6_outputs(2343) <= not a;
    layer6_outputs(2344) <= a;
    layer6_outputs(2345) <= a and not b;
    layer6_outputs(2346) <= not b or a;
    layer6_outputs(2347) <= a;
    layer6_outputs(2348) <= not (a or b);
    layer6_outputs(2349) <= not a;
    layer6_outputs(2350) <= not a;
    layer6_outputs(2351) <= b;
    layer6_outputs(2352) <= a and b;
    layer6_outputs(2353) <= a and b;
    layer6_outputs(2354) <= not b or a;
    layer6_outputs(2355) <= not (a or b);
    layer6_outputs(2356) <= not (a xor b);
    layer6_outputs(2357) <= not b;
    layer6_outputs(2358) <= a xor b;
    layer6_outputs(2359) <= b;
    layer6_outputs(2360) <= a or b;
    layer6_outputs(2361) <= not a or b;
    layer6_outputs(2362) <= b;
    layer6_outputs(2363) <= not b or a;
    layer6_outputs(2364) <= a and not b;
    layer6_outputs(2365) <= b;
    layer6_outputs(2366) <= a and b;
    layer6_outputs(2367) <= 1'b0;
    layer6_outputs(2368) <= not (a or b);
    layer6_outputs(2369) <= b and not a;
    layer6_outputs(2370) <= b;
    layer6_outputs(2371) <= a or b;
    layer6_outputs(2372) <= not a;
    layer6_outputs(2373) <= not a;
    layer6_outputs(2374) <= a and not b;
    layer6_outputs(2375) <= a or b;
    layer6_outputs(2376) <= not a or b;
    layer6_outputs(2377) <= a;
    layer6_outputs(2378) <= not b or a;
    layer6_outputs(2379) <= not b;
    layer6_outputs(2380) <= not (a xor b);
    layer6_outputs(2381) <= not a or b;
    layer6_outputs(2382) <= not a;
    layer6_outputs(2383) <= a;
    layer6_outputs(2384) <= not a;
    layer6_outputs(2385) <= 1'b0;
    layer6_outputs(2386) <= a or b;
    layer6_outputs(2387) <= b;
    layer6_outputs(2388) <= b and not a;
    layer6_outputs(2389) <= b and not a;
    layer6_outputs(2390) <= b;
    layer6_outputs(2391) <= a and not b;
    layer6_outputs(2392) <= a and not b;
    layer6_outputs(2393) <= not b;
    layer6_outputs(2394) <= a and b;
    layer6_outputs(2395) <= a;
    layer6_outputs(2396) <= a and not b;
    layer6_outputs(2397) <= b and not a;
    layer6_outputs(2398) <= not a or b;
    layer6_outputs(2399) <= not b;
    layer6_outputs(2400) <= a;
    layer6_outputs(2401) <= a xor b;
    layer6_outputs(2402) <= a;
    layer6_outputs(2403) <= not (a or b);
    layer6_outputs(2404) <= b;
    layer6_outputs(2405) <= b;
    layer6_outputs(2406) <= a;
    layer6_outputs(2407) <= b;
    layer6_outputs(2408) <= 1'b0;
    layer6_outputs(2409) <= not b;
    layer6_outputs(2410) <= not (a or b);
    layer6_outputs(2411) <= b and not a;
    layer6_outputs(2412) <= not a;
    layer6_outputs(2413) <= a;
    layer6_outputs(2414) <= 1'b1;
    layer6_outputs(2415) <= b;
    layer6_outputs(2416) <= 1'b0;
    layer6_outputs(2417) <= a xor b;
    layer6_outputs(2418) <= not a;
    layer6_outputs(2419) <= not (a and b);
    layer6_outputs(2420) <= b;
    layer6_outputs(2421) <= b and not a;
    layer6_outputs(2422) <= not (a and b);
    layer6_outputs(2423) <= a and not b;
    layer6_outputs(2424) <= not (a xor b);
    layer6_outputs(2425) <= a and not b;
    layer6_outputs(2426) <= a;
    layer6_outputs(2427) <= b and not a;
    layer6_outputs(2428) <= 1'b0;
    layer6_outputs(2429) <= b;
    layer6_outputs(2430) <= a and b;
    layer6_outputs(2431) <= a or b;
    layer6_outputs(2432) <= a xor b;
    layer6_outputs(2433) <= not b;
    layer6_outputs(2434) <= a;
    layer6_outputs(2435) <= a;
    layer6_outputs(2436) <= a and b;
    layer6_outputs(2437) <= not (a or b);
    layer6_outputs(2438) <= not b;
    layer6_outputs(2439) <= not (a xor b);
    layer6_outputs(2440) <= not (a and b);
    layer6_outputs(2441) <= not (a or b);
    layer6_outputs(2442) <= a;
    layer6_outputs(2443) <= not a;
    layer6_outputs(2444) <= b;
    layer6_outputs(2445) <= b;
    layer6_outputs(2446) <= a;
    layer6_outputs(2447) <= b and not a;
    layer6_outputs(2448) <= a or b;
    layer6_outputs(2449) <= b;
    layer6_outputs(2450) <= not a;
    layer6_outputs(2451) <= a xor b;
    layer6_outputs(2452) <= 1'b0;
    layer6_outputs(2453) <= a and not b;
    layer6_outputs(2454) <= b and not a;
    layer6_outputs(2455) <= not b;
    layer6_outputs(2456) <= not b;
    layer6_outputs(2457) <= b;
    layer6_outputs(2458) <= not a;
    layer6_outputs(2459) <= not (a or b);
    layer6_outputs(2460) <= not a;
    layer6_outputs(2461) <= a;
    layer6_outputs(2462) <= a;
    layer6_outputs(2463) <= a xor b;
    layer6_outputs(2464) <= a and b;
    layer6_outputs(2465) <= a;
    layer6_outputs(2466) <= not a;
    layer6_outputs(2467) <= not (a and b);
    layer6_outputs(2468) <= a;
    layer6_outputs(2469) <= b;
    layer6_outputs(2470) <= 1'b0;
    layer6_outputs(2471) <= b and not a;
    layer6_outputs(2472) <= not (a and b);
    layer6_outputs(2473) <= not b or a;
    layer6_outputs(2474) <= 1'b1;
    layer6_outputs(2475) <= not (a or b);
    layer6_outputs(2476) <= not (a or b);
    layer6_outputs(2477) <= not (a xor b);
    layer6_outputs(2478) <= not a;
    layer6_outputs(2479) <= b and not a;
    layer6_outputs(2480) <= b;
    layer6_outputs(2481) <= not (a and b);
    layer6_outputs(2482) <= not a;
    layer6_outputs(2483) <= not (a or b);
    layer6_outputs(2484) <= not (a or b);
    layer6_outputs(2485) <= not b;
    layer6_outputs(2486) <= not b;
    layer6_outputs(2487) <= a or b;
    layer6_outputs(2488) <= a;
    layer6_outputs(2489) <= not a or b;
    layer6_outputs(2490) <= a and b;
    layer6_outputs(2491) <= a;
    layer6_outputs(2492) <= b;
    layer6_outputs(2493) <= not b or a;
    layer6_outputs(2494) <= not (a xor b);
    layer6_outputs(2495) <= not b;
    layer6_outputs(2496) <= a;
    layer6_outputs(2497) <= a and b;
    layer6_outputs(2498) <= a;
    layer6_outputs(2499) <= a;
    layer6_outputs(2500) <= a xor b;
    layer6_outputs(2501) <= a xor b;
    layer6_outputs(2502) <= a and b;
    layer6_outputs(2503) <= a and not b;
    layer6_outputs(2504) <= not (a and b);
    layer6_outputs(2505) <= a;
    layer6_outputs(2506) <= not a;
    layer6_outputs(2507) <= b;
    layer6_outputs(2508) <= a or b;
    layer6_outputs(2509) <= not (a or b);
    layer6_outputs(2510) <= b and not a;
    layer6_outputs(2511) <= not a;
    layer6_outputs(2512) <= b;
    layer6_outputs(2513) <= a or b;
    layer6_outputs(2514) <= not b;
    layer6_outputs(2515) <= not a or b;
    layer6_outputs(2516) <= not a or b;
    layer6_outputs(2517) <= not b;
    layer6_outputs(2518) <= b;
    layer6_outputs(2519) <= not b;
    layer6_outputs(2520) <= b;
    layer6_outputs(2521) <= not (a xor b);
    layer6_outputs(2522) <= not a;
    layer6_outputs(2523) <= a or b;
    layer6_outputs(2524) <= not a;
    layer6_outputs(2525) <= a xor b;
    layer6_outputs(2526) <= b;
    layer6_outputs(2527) <= not b;
    layer6_outputs(2528) <= not b or a;
    layer6_outputs(2529) <= not b;
    layer6_outputs(2530) <= not (a xor b);
    layer6_outputs(2531) <= not a;
    layer6_outputs(2532) <= not (a or b);
    layer6_outputs(2533) <= 1'b1;
    layer6_outputs(2534) <= not a;
    layer6_outputs(2535) <= not a;
    layer6_outputs(2536) <= a;
    layer6_outputs(2537) <= b;
    layer6_outputs(2538) <= not (a and b);
    layer6_outputs(2539) <= a xor b;
    layer6_outputs(2540) <= not (a or b);
    layer6_outputs(2541) <= b;
    layer6_outputs(2542) <= not (a and b);
    layer6_outputs(2543) <= 1'b1;
    layer6_outputs(2544) <= not a or b;
    layer6_outputs(2545) <= not b or a;
    layer6_outputs(2546) <= b;
    layer6_outputs(2547) <= b and not a;
    layer6_outputs(2548) <= b;
    layer6_outputs(2549) <= a or b;
    layer6_outputs(2550) <= not a or b;
    layer6_outputs(2551) <= a or b;
    layer6_outputs(2552) <= a and not b;
    layer6_outputs(2553) <= b;
    layer6_outputs(2554) <= not b or a;
    layer6_outputs(2555) <= b;
    layer6_outputs(2556) <= b;
    layer6_outputs(2557) <= a and not b;
    layer6_outputs(2558) <= not (a and b);
    layer6_outputs(2559) <= not b or a;
    layer7_outputs(0) <= not a;
    layer7_outputs(1) <= not a;
    layer7_outputs(2) <= a;
    layer7_outputs(3) <= a;
    layer7_outputs(4) <= a and b;
    layer7_outputs(5) <= not (a or b);
    layer7_outputs(6) <= a or b;
    layer7_outputs(7) <= not (a and b);
    layer7_outputs(8) <= a;
    layer7_outputs(9) <= not (a xor b);
    layer7_outputs(10) <= not b;
    layer7_outputs(11) <= not (a xor b);
    layer7_outputs(12) <= not a;
    layer7_outputs(13) <= b;
    layer7_outputs(14) <= a;
    layer7_outputs(15) <= not (a and b);
    layer7_outputs(16) <= a or b;
    layer7_outputs(17) <= a;
    layer7_outputs(18) <= b;
    layer7_outputs(19) <= not b;
    layer7_outputs(20) <= not b;
    layer7_outputs(21) <= a xor b;
    layer7_outputs(22) <= not (a and b);
    layer7_outputs(23) <= b;
    layer7_outputs(24) <= not a or b;
    layer7_outputs(25) <= a;
    layer7_outputs(26) <= not b;
    layer7_outputs(27) <= not (a xor b);
    layer7_outputs(28) <= not (a or b);
    layer7_outputs(29) <= b;
    layer7_outputs(30) <= not a;
    layer7_outputs(31) <= a or b;
    layer7_outputs(32) <= not a;
    layer7_outputs(33) <= a and not b;
    layer7_outputs(34) <= a and b;
    layer7_outputs(35) <= a;
    layer7_outputs(36) <= a or b;
    layer7_outputs(37) <= not (a or b);
    layer7_outputs(38) <= not (a xor b);
    layer7_outputs(39) <= a xor b;
    layer7_outputs(40) <= b and not a;
    layer7_outputs(41) <= not b;
    layer7_outputs(42) <= not b or a;
    layer7_outputs(43) <= b and not a;
    layer7_outputs(44) <= not a;
    layer7_outputs(45) <= a;
    layer7_outputs(46) <= not a;
    layer7_outputs(47) <= not a;
    layer7_outputs(48) <= not a;
    layer7_outputs(49) <= a xor b;
    layer7_outputs(50) <= not a;
    layer7_outputs(51) <= not (a and b);
    layer7_outputs(52) <= b;
    layer7_outputs(53) <= not (a and b);
    layer7_outputs(54) <= a and b;
    layer7_outputs(55) <= a and b;
    layer7_outputs(56) <= not (a and b);
    layer7_outputs(57) <= a and b;
    layer7_outputs(58) <= a;
    layer7_outputs(59) <= a;
    layer7_outputs(60) <= not (a xor b);
    layer7_outputs(61) <= a or b;
    layer7_outputs(62) <= a xor b;
    layer7_outputs(63) <= not a or b;
    layer7_outputs(64) <= not a or b;
    layer7_outputs(65) <= not a;
    layer7_outputs(66) <= not b or a;
    layer7_outputs(67) <= a and b;
    layer7_outputs(68) <= not a or b;
    layer7_outputs(69) <= not (a or b);
    layer7_outputs(70) <= not a;
    layer7_outputs(71) <= not (a and b);
    layer7_outputs(72) <= a;
    layer7_outputs(73) <= a xor b;
    layer7_outputs(74) <= b and not a;
    layer7_outputs(75) <= not (a xor b);
    layer7_outputs(76) <= a and b;
    layer7_outputs(77) <= not b;
    layer7_outputs(78) <= a;
    layer7_outputs(79) <= a and not b;
    layer7_outputs(80) <= a xor b;
    layer7_outputs(81) <= a;
    layer7_outputs(82) <= not (a or b);
    layer7_outputs(83) <= not a;
    layer7_outputs(84) <= a xor b;
    layer7_outputs(85) <= b;
    layer7_outputs(86) <= not (a or b);
    layer7_outputs(87) <= b and not a;
    layer7_outputs(88) <= a;
    layer7_outputs(89) <= not (a and b);
    layer7_outputs(90) <= not b or a;
    layer7_outputs(91) <= not a;
    layer7_outputs(92) <= 1'b1;
    layer7_outputs(93) <= not (a or b);
    layer7_outputs(94) <= not b;
    layer7_outputs(95) <= not b or a;
    layer7_outputs(96) <= a and not b;
    layer7_outputs(97) <= b;
    layer7_outputs(98) <= not (a or b);
    layer7_outputs(99) <= a;
    layer7_outputs(100) <= not b;
    layer7_outputs(101) <= not a or b;
    layer7_outputs(102) <= not (a and b);
    layer7_outputs(103) <= not (a xor b);
    layer7_outputs(104) <= not b;
    layer7_outputs(105) <= b;
    layer7_outputs(106) <= a or b;
    layer7_outputs(107) <= not b or a;
    layer7_outputs(108) <= b;
    layer7_outputs(109) <= b and not a;
    layer7_outputs(110) <= a;
    layer7_outputs(111) <= not a;
    layer7_outputs(112) <= a and not b;
    layer7_outputs(113) <= not a;
    layer7_outputs(114) <= not (a or b);
    layer7_outputs(115) <= a and b;
    layer7_outputs(116) <= b and not a;
    layer7_outputs(117) <= not b;
    layer7_outputs(118) <= b and not a;
    layer7_outputs(119) <= not a or b;
    layer7_outputs(120) <= b;
    layer7_outputs(121) <= not a;
    layer7_outputs(122) <= not (a xor b);
    layer7_outputs(123) <= not b;
    layer7_outputs(124) <= not (a and b);
    layer7_outputs(125) <= not (a and b);
    layer7_outputs(126) <= a or b;
    layer7_outputs(127) <= a or b;
    layer7_outputs(128) <= a xor b;
    layer7_outputs(129) <= not (a xor b);
    layer7_outputs(130) <= not a;
    layer7_outputs(131) <= b;
    layer7_outputs(132) <= b;
    layer7_outputs(133) <= a or b;
    layer7_outputs(134) <= not b or a;
    layer7_outputs(135) <= a or b;
    layer7_outputs(136) <= b;
    layer7_outputs(137) <= a or b;
    layer7_outputs(138) <= 1'b1;
    layer7_outputs(139) <= not b or a;
    layer7_outputs(140) <= not (a or b);
    layer7_outputs(141) <= not (a or b);
    layer7_outputs(142) <= a or b;
    layer7_outputs(143) <= not (a xor b);
    layer7_outputs(144) <= a;
    layer7_outputs(145) <= b;
    layer7_outputs(146) <= not a;
    layer7_outputs(147) <= not a or b;
    layer7_outputs(148) <= a and b;
    layer7_outputs(149) <= a xor b;
    layer7_outputs(150) <= not (a or b);
    layer7_outputs(151) <= not (a xor b);
    layer7_outputs(152) <= not b;
    layer7_outputs(153) <= 1'b0;
    layer7_outputs(154) <= not b;
    layer7_outputs(155) <= not b;
    layer7_outputs(156) <= not (a or b);
    layer7_outputs(157) <= not (a or b);
    layer7_outputs(158) <= not a or b;
    layer7_outputs(159) <= a;
    layer7_outputs(160) <= not a;
    layer7_outputs(161) <= not b or a;
    layer7_outputs(162) <= a;
    layer7_outputs(163) <= not b;
    layer7_outputs(164) <= a or b;
    layer7_outputs(165) <= not b;
    layer7_outputs(166) <= a or b;
    layer7_outputs(167) <= not b or a;
    layer7_outputs(168) <= not a;
    layer7_outputs(169) <= not b or a;
    layer7_outputs(170) <= a and b;
    layer7_outputs(171) <= not b or a;
    layer7_outputs(172) <= not b;
    layer7_outputs(173) <= a xor b;
    layer7_outputs(174) <= a;
    layer7_outputs(175) <= not (a xor b);
    layer7_outputs(176) <= a;
    layer7_outputs(177) <= not b;
    layer7_outputs(178) <= not a or b;
    layer7_outputs(179) <= not a;
    layer7_outputs(180) <= a xor b;
    layer7_outputs(181) <= a;
    layer7_outputs(182) <= a;
    layer7_outputs(183) <= b;
    layer7_outputs(184) <= not (a xor b);
    layer7_outputs(185) <= b;
    layer7_outputs(186) <= b;
    layer7_outputs(187) <= b;
    layer7_outputs(188) <= b;
    layer7_outputs(189) <= not (a and b);
    layer7_outputs(190) <= not a or b;
    layer7_outputs(191) <= not b or a;
    layer7_outputs(192) <= b;
    layer7_outputs(193) <= not b;
    layer7_outputs(194) <= a and not b;
    layer7_outputs(195) <= not (a and b);
    layer7_outputs(196) <= not b;
    layer7_outputs(197) <= b;
    layer7_outputs(198) <= a and not b;
    layer7_outputs(199) <= not (a xor b);
    layer7_outputs(200) <= not (a or b);
    layer7_outputs(201) <= a;
    layer7_outputs(202) <= not a;
    layer7_outputs(203) <= a and not b;
    layer7_outputs(204) <= a xor b;
    layer7_outputs(205) <= a and b;
    layer7_outputs(206) <= b;
    layer7_outputs(207) <= not b or a;
    layer7_outputs(208) <= not b;
    layer7_outputs(209) <= not a;
    layer7_outputs(210) <= a;
    layer7_outputs(211) <= a;
    layer7_outputs(212) <= not b;
    layer7_outputs(213) <= not a;
    layer7_outputs(214) <= not b or a;
    layer7_outputs(215) <= not (a xor b);
    layer7_outputs(216) <= not a or b;
    layer7_outputs(217) <= a;
    layer7_outputs(218) <= a or b;
    layer7_outputs(219) <= not (a or b);
    layer7_outputs(220) <= b;
    layer7_outputs(221) <= a and b;
    layer7_outputs(222) <= a;
    layer7_outputs(223) <= a xor b;
    layer7_outputs(224) <= 1'b0;
    layer7_outputs(225) <= a;
    layer7_outputs(226) <= b;
    layer7_outputs(227) <= not (a and b);
    layer7_outputs(228) <= not (a xor b);
    layer7_outputs(229) <= a;
    layer7_outputs(230) <= not (a or b);
    layer7_outputs(231) <= not b;
    layer7_outputs(232) <= not (a or b);
    layer7_outputs(233) <= not a;
    layer7_outputs(234) <= a;
    layer7_outputs(235) <= a and b;
    layer7_outputs(236) <= 1'b1;
    layer7_outputs(237) <= b;
    layer7_outputs(238) <= a xor b;
    layer7_outputs(239) <= b and not a;
    layer7_outputs(240) <= a and b;
    layer7_outputs(241) <= not (a and b);
    layer7_outputs(242) <= a;
    layer7_outputs(243) <= not (a or b);
    layer7_outputs(244) <= a;
    layer7_outputs(245) <= a xor b;
    layer7_outputs(246) <= not b or a;
    layer7_outputs(247) <= a;
    layer7_outputs(248) <= not a;
    layer7_outputs(249) <= a;
    layer7_outputs(250) <= b;
    layer7_outputs(251) <= not b;
    layer7_outputs(252) <= not b or a;
    layer7_outputs(253) <= not b;
    layer7_outputs(254) <= a and b;
    layer7_outputs(255) <= not (a or b);
    layer7_outputs(256) <= a xor b;
    layer7_outputs(257) <= b;
    layer7_outputs(258) <= b and not a;
    layer7_outputs(259) <= 1'b1;
    layer7_outputs(260) <= b;
    layer7_outputs(261) <= not b;
    layer7_outputs(262) <= a;
    layer7_outputs(263) <= b;
    layer7_outputs(264) <= not (a xor b);
    layer7_outputs(265) <= not a or b;
    layer7_outputs(266) <= not a;
    layer7_outputs(267) <= b and not a;
    layer7_outputs(268) <= a or b;
    layer7_outputs(269) <= not b;
    layer7_outputs(270) <= not b or a;
    layer7_outputs(271) <= not b or a;
    layer7_outputs(272) <= not a or b;
    layer7_outputs(273) <= not (a xor b);
    layer7_outputs(274) <= not b;
    layer7_outputs(275) <= a;
    layer7_outputs(276) <= not a;
    layer7_outputs(277) <= a xor b;
    layer7_outputs(278) <= a;
    layer7_outputs(279) <= not (a xor b);
    layer7_outputs(280) <= 1'b0;
    layer7_outputs(281) <= not a or b;
    layer7_outputs(282) <= b and not a;
    layer7_outputs(283) <= a and b;
    layer7_outputs(284) <= not (a and b);
    layer7_outputs(285) <= not (a and b);
    layer7_outputs(286) <= not b;
    layer7_outputs(287) <= not b;
    layer7_outputs(288) <= not a;
    layer7_outputs(289) <= b;
    layer7_outputs(290) <= a xor b;
    layer7_outputs(291) <= b;
    layer7_outputs(292) <= not a;
    layer7_outputs(293) <= not b;
    layer7_outputs(294) <= b;
    layer7_outputs(295) <= not b;
    layer7_outputs(296) <= b and not a;
    layer7_outputs(297) <= a and b;
    layer7_outputs(298) <= not a;
    layer7_outputs(299) <= b;
    layer7_outputs(300) <= a;
    layer7_outputs(301) <= b;
    layer7_outputs(302) <= not b or a;
    layer7_outputs(303) <= a;
    layer7_outputs(304) <= b;
    layer7_outputs(305) <= not a or b;
    layer7_outputs(306) <= 1'b0;
    layer7_outputs(307) <= a and b;
    layer7_outputs(308) <= not a;
    layer7_outputs(309) <= not a;
    layer7_outputs(310) <= 1'b0;
    layer7_outputs(311) <= 1'b1;
    layer7_outputs(312) <= not a or b;
    layer7_outputs(313) <= a and b;
    layer7_outputs(314) <= a;
    layer7_outputs(315) <= a;
    layer7_outputs(316) <= b and not a;
    layer7_outputs(317) <= not (a and b);
    layer7_outputs(318) <= a;
    layer7_outputs(319) <= a;
    layer7_outputs(320) <= a or b;
    layer7_outputs(321) <= not a or b;
    layer7_outputs(322) <= a;
    layer7_outputs(323) <= not (a and b);
    layer7_outputs(324) <= b and not a;
    layer7_outputs(325) <= not b or a;
    layer7_outputs(326) <= not a;
    layer7_outputs(327) <= not (a or b);
    layer7_outputs(328) <= a or b;
    layer7_outputs(329) <= not (a and b);
    layer7_outputs(330) <= a and not b;
    layer7_outputs(331) <= not a;
    layer7_outputs(332) <= a and b;
    layer7_outputs(333) <= a xor b;
    layer7_outputs(334) <= b;
    layer7_outputs(335) <= not (a xor b);
    layer7_outputs(336) <= not b;
    layer7_outputs(337) <= b and not a;
    layer7_outputs(338) <= a xor b;
    layer7_outputs(339) <= a and b;
    layer7_outputs(340) <= not b;
    layer7_outputs(341) <= not (a xor b);
    layer7_outputs(342) <= a;
    layer7_outputs(343) <= b;
    layer7_outputs(344) <= b and not a;
    layer7_outputs(345) <= a xor b;
    layer7_outputs(346) <= 1'b0;
    layer7_outputs(347) <= not b;
    layer7_outputs(348) <= b and not a;
    layer7_outputs(349) <= b and not a;
    layer7_outputs(350) <= not b or a;
    layer7_outputs(351) <= b;
    layer7_outputs(352) <= a or b;
    layer7_outputs(353) <= a and not b;
    layer7_outputs(354) <= b and not a;
    layer7_outputs(355) <= not (a xor b);
    layer7_outputs(356) <= 1'b0;
    layer7_outputs(357) <= not b or a;
    layer7_outputs(358) <= not b or a;
    layer7_outputs(359) <= a xor b;
    layer7_outputs(360) <= b;
    layer7_outputs(361) <= not b or a;
    layer7_outputs(362) <= not (a and b);
    layer7_outputs(363) <= a;
    layer7_outputs(364) <= not (a or b);
    layer7_outputs(365) <= not a;
    layer7_outputs(366) <= a xor b;
    layer7_outputs(367) <= not a or b;
    layer7_outputs(368) <= a xor b;
    layer7_outputs(369) <= not (a or b);
    layer7_outputs(370) <= not (a or b);
    layer7_outputs(371) <= not a;
    layer7_outputs(372) <= a or b;
    layer7_outputs(373) <= a xor b;
    layer7_outputs(374) <= a and b;
    layer7_outputs(375) <= b;
    layer7_outputs(376) <= a xor b;
    layer7_outputs(377) <= a and b;
    layer7_outputs(378) <= a and not b;
    layer7_outputs(379) <= not b;
    layer7_outputs(380) <= not b or a;
    layer7_outputs(381) <= not b;
    layer7_outputs(382) <= not a;
    layer7_outputs(383) <= b;
    layer7_outputs(384) <= a or b;
    layer7_outputs(385) <= a and b;
    layer7_outputs(386) <= a and b;
    layer7_outputs(387) <= a and not b;
    layer7_outputs(388) <= a or b;
    layer7_outputs(389) <= a xor b;
    layer7_outputs(390) <= not a;
    layer7_outputs(391) <= not a;
    layer7_outputs(392) <= b;
    layer7_outputs(393) <= b and not a;
    layer7_outputs(394) <= not b;
    layer7_outputs(395) <= a and not b;
    layer7_outputs(396) <= b;
    layer7_outputs(397) <= not (a or b);
    layer7_outputs(398) <= not (a xor b);
    layer7_outputs(399) <= a or b;
    layer7_outputs(400) <= b;
    layer7_outputs(401) <= not a or b;
    layer7_outputs(402) <= b and not a;
    layer7_outputs(403) <= a;
    layer7_outputs(404) <= b;
    layer7_outputs(405) <= not b;
    layer7_outputs(406) <= a xor b;
    layer7_outputs(407) <= b;
    layer7_outputs(408) <= not a or b;
    layer7_outputs(409) <= not b;
    layer7_outputs(410) <= b;
    layer7_outputs(411) <= a xor b;
    layer7_outputs(412) <= not (a or b);
    layer7_outputs(413) <= b;
    layer7_outputs(414) <= a and not b;
    layer7_outputs(415) <= a or b;
    layer7_outputs(416) <= not a;
    layer7_outputs(417) <= not a or b;
    layer7_outputs(418) <= b;
    layer7_outputs(419) <= not (a or b);
    layer7_outputs(420) <= a and not b;
    layer7_outputs(421) <= b;
    layer7_outputs(422) <= a;
    layer7_outputs(423) <= a and not b;
    layer7_outputs(424) <= not (a or b);
    layer7_outputs(425) <= b and not a;
    layer7_outputs(426) <= b;
    layer7_outputs(427) <= a and b;
    layer7_outputs(428) <= b;
    layer7_outputs(429) <= not a or b;
    layer7_outputs(430) <= not b;
    layer7_outputs(431) <= a or b;
    layer7_outputs(432) <= b;
    layer7_outputs(433) <= not a;
    layer7_outputs(434) <= not b;
    layer7_outputs(435) <= a;
    layer7_outputs(436) <= a;
    layer7_outputs(437) <= not (a or b);
    layer7_outputs(438) <= not a or b;
    layer7_outputs(439) <= a xor b;
    layer7_outputs(440) <= not a or b;
    layer7_outputs(441) <= not b or a;
    layer7_outputs(442) <= not b;
    layer7_outputs(443) <= a or b;
    layer7_outputs(444) <= a and b;
    layer7_outputs(445) <= not (a or b);
    layer7_outputs(446) <= a or b;
    layer7_outputs(447) <= not a;
    layer7_outputs(448) <= b and not a;
    layer7_outputs(449) <= not (a or b);
    layer7_outputs(450) <= not b or a;
    layer7_outputs(451) <= a and not b;
    layer7_outputs(452) <= not a or b;
    layer7_outputs(453) <= b;
    layer7_outputs(454) <= not (a or b);
    layer7_outputs(455) <= b;
    layer7_outputs(456) <= a;
    layer7_outputs(457) <= not b;
    layer7_outputs(458) <= not a or b;
    layer7_outputs(459) <= a and b;
    layer7_outputs(460) <= not a;
    layer7_outputs(461) <= not b or a;
    layer7_outputs(462) <= a and b;
    layer7_outputs(463) <= not (a and b);
    layer7_outputs(464) <= a or b;
    layer7_outputs(465) <= a;
    layer7_outputs(466) <= a;
    layer7_outputs(467) <= not b;
    layer7_outputs(468) <= a;
    layer7_outputs(469) <= not (a or b);
    layer7_outputs(470) <= a or b;
    layer7_outputs(471) <= a or b;
    layer7_outputs(472) <= a and not b;
    layer7_outputs(473) <= a and not b;
    layer7_outputs(474) <= b and not a;
    layer7_outputs(475) <= a xor b;
    layer7_outputs(476) <= not (a or b);
    layer7_outputs(477) <= b;
    layer7_outputs(478) <= not (a and b);
    layer7_outputs(479) <= not (a or b);
    layer7_outputs(480) <= a and b;
    layer7_outputs(481) <= not (a xor b);
    layer7_outputs(482) <= b;
    layer7_outputs(483) <= not (a or b);
    layer7_outputs(484) <= a and not b;
    layer7_outputs(485) <= not (a and b);
    layer7_outputs(486) <= a xor b;
    layer7_outputs(487) <= not (a and b);
    layer7_outputs(488) <= a or b;
    layer7_outputs(489) <= not b or a;
    layer7_outputs(490) <= a and not b;
    layer7_outputs(491) <= b;
    layer7_outputs(492) <= b and not a;
    layer7_outputs(493) <= a and b;
    layer7_outputs(494) <= a and not b;
    layer7_outputs(495) <= not (a and b);
    layer7_outputs(496) <= a and b;
    layer7_outputs(497) <= a and not b;
    layer7_outputs(498) <= b;
    layer7_outputs(499) <= not a;
    layer7_outputs(500) <= not (a or b);
    layer7_outputs(501) <= not (a or b);
    layer7_outputs(502) <= not a or b;
    layer7_outputs(503) <= not (a or b);
    layer7_outputs(504) <= b;
    layer7_outputs(505) <= a or b;
    layer7_outputs(506) <= not b or a;
    layer7_outputs(507) <= not b or a;
    layer7_outputs(508) <= a xor b;
    layer7_outputs(509) <= b and not a;
    layer7_outputs(510) <= b and not a;
    layer7_outputs(511) <= not a;
    layer7_outputs(512) <= 1'b1;
    layer7_outputs(513) <= b and not a;
    layer7_outputs(514) <= not (a and b);
    layer7_outputs(515) <= a or b;
    layer7_outputs(516) <= b and not a;
    layer7_outputs(517) <= a;
    layer7_outputs(518) <= not (a and b);
    layer7_outputs(519) <= not b;
    layer7_outputs(520) <= not a;
    layer7_outputs(521) <= a and not b;
    layer7_outputs(522) <= not (a or b);
    layer7_outputs(523) <= b;
    layer7_outputs(524) <= not a;
    layer7_outputs(525) <= b;
    layer7_outputs(526) <= not b or a;
    layer7_outputs(527) <= a;
    layer7_outputs(528) <= not (a and b);
    layer7_outputs(529) <= not (a or b);
    layer7_outputs(530) <= not a;
    layer7_outputs(531) <= a;
    layer7_outputs(532) <= b;
    layer7_outputs(533) <= b and not a;
    layer7_outputs(534) <= a;
    layer7_outputs(535) <= b;
    layer7_outputs(536) <= a or b;
    layer7_outputs(537) <= not (a or b);
    layer7_outputs(538) <= not (a and b);
    layer7_outputs(539) <= a;
    layer7_outputs(540) <= a and not b;
    layer7_outputs(541) <= a;
    layer7_outputs(542) <= a;
    layer7_outputs(543) <= b;
    layer7_outputs(544) <= not b or a;
    layer7_outputs(545) <= not a or b;
    layer7_outputs(546) <= not (a or b);
    layer7_outputs(547) <= b and not a;
    layer7_outputs(548) <= not a;
    layer7_outputs(549) <= not a;
    layer7_outputs(550) <= b;
    layer7_outputs(551) <= a;
    layer7_outputs(552) <= not b or a;
    layer7_outputs(553) <= not a or b;
    layer7_outputs(554) <= not a;
    layer7_outputs(555) <= not a;
    layer7_outputs(556) <= not b;
    layer7_outputs(557) <= b;
    layer7_outputs(558) <= b and not a;
    layer7_outputs(559) <= not a;
    layer7_outputs(560) <= not a;
    layer7_outputs(561) <= b;
    layer7_outputs(562) <= b;
    layer7_outputs(563) <= a and not b;
    layer7_outputs(564) <= not a;
    layer7_outputs(565) <= a;
    layer7_outputs(566) <= not (a xor b);
    layer7_outputs(567) <= not a;
    layer7_outputs(568) <= not b;
    layer7_outputs(569) <= a and b;
    layer7_outputs(570) <= not a or b;
    layer7_outputs(571) <= not (a and b);
    layer7_outputs(572) <= a and not b;
    layer7_outputs(573) <= a;
    layer7_outputs(574) <= b and not a;
    layer7_outputs(575) <= a xor b;
    layer7_outputs(576) <= 1'b0;
    layer7_outputs(577) <= not (a or b);
    layer7_outputs(578) <= not a or b;
    layer7_outputs(579) <= not a;
    layer7_outputs(580) <= not a;
    layer7_outputs(581) <= a and not b;
    layer7_outputs(582) <= a;
    layer7_outputs(583) <= a;
    layer7_outputs(584) <= a or b;
    layer7_outputs(585) <= not b;
    layer7_outputs(586) <= a and not b;
    layer7_outputs(587) <= not (a xor b);
    layer7_outputs(588) <= a or b;
    layer7_outputs(589) <= a;
    layer7_outputs(590) <= a and b;
    layer7_outputs(591) <= b;
    layer7_outputs(592) <= b;
    layer7_outputs(593) <= b;
    layer7_outputs(594) <= b;
    layer7_outputs(595) <= b and not a;
    layer7_outputs(596) <= not a or b;
    layer7_outputs(597) <= not b or a;
    layer7_outputs(598) <= b;
    layer7_outputs(599) <= a;
    layer7_outputs(600) <= not a or b;
    layer7_outputs(601) <= a and not b;
    layer7_outputs(602) <= not b or a;
    layer7_outputs(603) <= not a;
    layer7_outputs(604) <= a xor b;
    layer7_outputs(605) <= not b;
    layer7_outputs(606) <= not (a xor b);
    layer7_outputs(607) <= a and not b;
    layer7_outputs(608) <= a or b;
    layer7_outputs(609) <= not (a xor b);
    layer7_outputs(610) <= a xor b;
    layer7_outputs(611) <= a and b;
    layer7_outputs(612) <= b and not a;
    layer7_outputs(613) <= a xor b;
    layer7_outputs(614) <= not a;
    layer7_outputs(615) <= not (a and b);
    layer7_outputs(616) <= a;
    layer7_outputs(617) <= not a;
    layer7_outputs(618) <= not (a xor b);
    layer7_outputs(619) <= a or b;
    layer7_outputs(620) <= a xor b;
    layer7_outputs(621) <= b;
    layer7_outputs(622) <= not (a and b);
    layer7_outputs(623) <= a xor b;
    layer7_outputs(624) <= not (a or b);
    layer7_outputs(625) <= a and not b;
    layer7_outputs(626) <= b and not a;
    layer7_outputs(627) <= b;
    layer7_outputs(628) <= b and not a;
    layer7_outputs(629) <= a;
    layer7_outputs(630) <= not b;
    layer7_outputs(631) <= not b or a;
    layer7_outputs(632) <= b;
    layer7_outputs(633) <= not b;
    layer7_outputs(634) <= a xor b;
    layer7_outputs(635) <= not a;
    layer7_outputs(636) <= not b;
    layer7_outputs(637) <= not a;
    layer7_outputs(638) <= not (a and b);
    layer7_outputs(639) <= b;
    layer7_outputs(640) <= b and not a;
    layer7_outputs(641) <= b;
    layer7_outputs(642) <= a xor b;
    layer7_outputs(643) <= a or b;
    layer7_outputs(644) <= not b;
    layer7_outputs(645) <= a and b;
    layer7_outputs(646) <= a;
    layer7_outputs(647) <= b;
    layer7_outputs(648) <= b;
    layer7_outputs(649) <= not b;
    layer7_outputs(650) <= a;
    layer7_outputs(651) <= b and not a;
    layer7_outputs(652) <= 1'b1;
    layer7_outputs(653) <= not a or b;
    layer7_outputs(654) <= not b;
    layer7_outputs(655) <= not b or a;
    layer7_outputs(656) <= a xor b;
    layer7_outputs(657) <= not a;
    layer7_outputs(658) <= not a or b;
    layer7_outputs(659) <= a;
    layer7_outputs(660) <= a or b;
    layer7_outputs(661) <= b;
    layer7_outputs(662) <= not (a xor b);
    layer7_outputs(663) <= a;
    layer7_outputs(664) <= not b;
    layer7_outputs(665) <= b;
    layer7_outputs(666) <= a or b;
    layer7_outputs(667) <= not a;
    layer7_outputs(668) <= b and not a;
    layer7_outputs(669) <= not (a or b);
    layer7_outputs(670) <= a xor b;
    layer7_outputs(671) <= a or b;
    layer7_outputs(672) <= a;
    layer7_outputs(673) <= not a or b;
    layer7_outputs(674) <= not (a or b);
    layer7_outputs(675) <= a;
    layer7_outputs(676) <= not a;
    layer7_outputs(677) <= b;
    layer7_outputs(678) <= b;
    layer7_outputs(679) <= a xor b;
    layer7_outputs(680) <= a and b;
    layer7_outputs(681) <= not b;
    layer7_outputs(682) <= not b or a;
    layer7_outputs(683) <= not (a and b);
    layer7_outputs(684) <= not b or a;
    layer7_outputs(685) <= b;
    layer7_outputs(686) <= not (a and b);
    layer7_outputs(687) <= not a;
    layer7_outputs(688) <= a;
    layer7_outputs(689) <= a xor b;
    layer7_outputs(690) <= not (a and b);
    layer7_outputs(691) <= not a;
    layer7_outputs(692) <= not a;
    layer7_outputs(693) <= b and not a;
    layer7_outputs(694) <= b and not a;
    layer7_outputs(695) <= not a or b;
    layer7_outputs(696) <= not a or b;
    layer7_outputs(697) <= not (a or b);
    layer7_outputs(698) <= a or b;
    layer7_outputs(699) <= not (a or b);
    layer7_outputs(700) <= a and b;
    layer7_outputs(701) <= b;
    layer7_outputs(702) <= not (a or b);
    layer7_outputs(703) <= a or b;
    layer7_outputs(704) <= not (a and b);
    layer7_outputs(705) <= b;
    layer7_outputs(706) <= a and not b;
    layer7_outputs(707) <= b;
    layer7_outputs(708) <= a;
    layer7_outputs(709) <= b and not a;
    layer7_outputs(710) <= not b;
    layer7_outputs(711) <= a;
    layer7_outputs(712) <= a;
    layer7_outputs(713) <= a;
    layer7_outputs(714) <= a and not b;
    layer7_outputs(715) <= a and b;
    layer7_outputs(716) <= not a;
    layer7_outputs(717) <= not a;
    layer7_outputs(718) <= not b or a;
    layer7_outputs(719) <= not a;
    layer7_outputs(720) <= not (a xor b);
    layer7_outputs(721) <= a or b;
    layer7_outputs(722) <= a and b;
    layer7_outputs(723) <= not (a or b);
    layer7_outputs(724) <= b;
    layer7_outputs(725) <= not (a or b);
    layer7_outputs(726) <= not a or b;
    layer7_outputs(727) <= b and not a;
    layer7_outputs(728) <= not (a xor b);
    layer7_outputs(729) <= a;
    layer7_outputs(730) <= not (a and b);
    layer7_outputs(731) <= a and b;
    layer7_outputs(732) <= a and b;
    layer7_outputs(733) <= a;
    layer7_outputs(734) <= a;
    layer7_outputs(735) <= a xor b;
    layer7_outputs(736) <= not (a xor b);
    layer7_outputs(737) <= not b;
    layer7_outputs(738) <= a and not b;
    layer7_outputs(739) <= not (a and b);
    layer7_outputs(740) <= a xor b;
    layer7_outputs(741) <= not (a xor b);
    layer7_outputs(742) <= not b;
    layer7_outputs(743) <= not b;
    layer7_outputs(744) <= b;
    layer7_outputs(745) <= a;
    layer7_outputs(746) <= not b;
    layer7_outputs(747) <= a or b;
    layer7_outputs(748) <= not b;
    layer7_outputs(749) <= not (a or b);
    layer7_outputs(750) <= not a;
    layer7_outputs(751) <= not (a xor b);
    layer7_outputs(752) <= not b or a;
    layer7_outputs(753) <= 1'b1;
    layer7_outputs(754) <= not b;
    layer7_outputs(755) <= not (a or b);
    layer7_outputs(756) <= a and not b;
    layer7_outputs(757) <= not a;
    layer7_outputs(758) <= not (a or b);
    layer7_outputs(759) <= a and not b;
    layer7_outputs(760) <= not a;
    layer7_outputs(761) <= a and not b;
    layer7_outputs(762) <= not (a or b);
    layer7_outputs(763) <= a;
    layer7_outputs(764) <= a or b;
    layer7_outputs(765) <= b;
    layer7_outputs(766) <= a and not b;
    layer7_outputs(767) <= not b;
    layer7_outputs(768) <= not (a and b);
    layer7_outputs(769) <= not a;
    layer7_outputs(770) <= not a;
    layer7_outputs(771) <= a or b;
    layer7_outputs(772) <= not (a and b);
    layer7_outputs(773) <= a;
    layer7_outputs(774) <= not b;
    layer7_outputs(775) <= a or b;
    layer7_outputs(776) <= b;
    layer7_outputs(777) <= not a;
    layer7_outputs(778) <= a xor b;
    layer7_outputs(779) <= not b;
    layer7_outputs(780) <= not (a xor b);
    layer7_outputs(781) <= a;
    layer7_outputs(782) <= not b;
    layer7_outputs(783) <= a;
    layer7_outputs(784) <= b and not a;
    layer7_outputs(785) <= b;
    layer7_outputs(786) <= not a;
    layer7_outputs(787) <= not b;
    layer7_outputs(788) <= a or b;
    layer7_outputs(789) <= a;
    layer7_outputs(790) <= b and not a;
    layer7_outputs(791) <= a xor b;
    layer7_outputs(792) <= b;
    layer7_outputs(793) <= not b;
    layer7_outputs(794) <= b;
    layer7_outputs(795) <= not a;
    layer7_outputs(796) <= not (a xor b);
    layer7_outputs(797) <= not a;
    layer7_outputs(798) <= not b;
    layer7_outputs(799) <= b;
    layer7_outputs(800) <= not (a or b);
    layer7_outputs(801) <= not (a or b);
    layer7_outputs(802) <= a and b;
    layer7_outputs(803) <= b;
    layer7_outputs(804) <= not a;
    layer7_outputs(805) <= not a or b;
    layer7_outputs(806) <= a or b;
    layer7_outputs(807) <= b;
    layer7_outputs(808) <= not a;
    layer7_outputs(809) <= not a;
    layer7_outputs(810) <= a;
    layer7_outputs(811) <= b and not a;
    layer7_outputs(812) <= a and not b;
    layer7_outputs(813) <= a and b;
    layer7_outputs(814) <= b and not a;
    layer7_outputs(815) <= a and not b;
    layer7_outputs(816) <= a and not b;
    layer7_outputs(817) <= not a;
    layer7_outputs(818) <= not a;
    layer7_outputs(819) <= b;
    layer7_outputs(820) <= b;
    layer7_outputs(821) <= not b or a;
    layer7_outputs(822) <= b;
    layer7_outputs(823) <= not (a xor b);
    layer7_outputs(824) <= not a;
    layer7_outputs(825) <= not a or b;
    layer7_outputs(826) <= not b;
    layer7_outputs(827) <= 1'b1;
    layer7_outputs(828) <= not a;
    layer7_outputs(829) <= b;
    layer7_outputs(830) <= not a or b;
    layer7_outputs(831) <= b;
    layer7_outputs(832) <= b;
    layer7_outputs(833) <= not (a xor b);
    layer7_outputs(834) <= not (a xor b);
    layer7_outputs(835) <= not (a and b);
    layer7_outputs(836) <= not b;
    layer7_outputs(837) <= a or b;
    layer7_outputs(838) <= not a or b;
    layer7_outputs(839) <= not a;
    layer7_outputs(840) <= a xor b;
    layer7_outputs(841) <= not (a xor b);
    layer7_outputs(842) <= not b;
    layer7_outputs(843) <= a;
    layer7_outputs(844) <= not a or b;
    layer7_outputs(845) <= not a;
    layer7_outputs(846) <= b;
    layer7_outputs(847) <= a or b;
    layer7_outputs(848) <= not b;
    layer7_outputs(849) <= b;
    layer7_outputs(850) <= a and not b;
    layer7_outputs(851) <= not b or a;
    layer7_outputs(852) <= not b;
    layer7_outputs(853) <= not a;
    layer7_outputs(854) <= b;
    layer7_outputs(855) <= not b or a;
    layer7_outputs(856) <= not (a or b);
    layer7_outputs(857) <= not a;
    layer7_outputs(858) <= a and not b;
    layer7_outputs(859) <= not a;
    layer7_outputs(860) <= not b;
    layer7_outputs(861) <= not (a or b);
    layer7_outputs(862) <= not a or b;
    layer7_outputs(863) <= b;
    layer7_outputs(864) <= b;
    layer7_outputs(865) <= not a;
    layer7_outputs(866) <= not a;
    layer7_outputs(867) <= not a or b;
    layer7_outputs(868) <= b;
    layer7_outputs(869) <= a xor b;
    layer7_outputs(870) <= not a or b;
    layer7_outputs(871) <= not (a xor b);
    layer7_outputs(872) <= a or b;
    layer7_outputs(873) <= not b or a;
    layer7_outputs(874) <= a;
    layer7_outputs(875) <= a xor b;
    layer7_outputs(876) <= not a or b;
    layer7_outputs(877) <= not (a xor b);
    layer7_outputs(878) <= a and b;
    layer7_outputs(879) <= b and not a;
    layer7_outputs(880) <= not (a and b);
    layer7_outputs(881) <= b;
    layer7_outputs(882) <= a and not b;
    layer7_outputs(883) <= not b or a;
    layer7_outputs(884) <= not a or b;
    layer7_outputs(885) <= a;
    layer7_outputs(886) <= 1'b1;
    layer7_outputs(887) <= 1'b1;
    layer7_outputs(888) <= not (a xor b);
    layer7_outputs(889) <= not (a xor b);
    layer7_outputs(890) <= not b;
    layer7_outputs(891) <= not (a or b);
    layer7_outputs(892) <= not a;
    layer7_outputs(893) <= a and not b;
    layer7_outputs(894) <= not b;
    layer7_outputs(895) <= b;
    layer7_outputs(896) <= a and b;
    layer7_outputs(897) <= not b;
    layer7_outputs(898) <= a and not b;
    layer7_outputs(899) <= not a or b;
    layer7_outputs(900) <= b and not a;
    layer7_outputs(901) <= a;
    layer7_outputs(902) <= not a;
    layer7_outputs(903) <= not a;
    layer7_outputs(904) <= a;
    layer7_outputs(905) <= not b;
    layer7_outputs(906) <= b;
    layer7_outputs(907) <= not (a xor b);
    layer7_outputs(908) <= a xor b;
    layer7_outputs(909) <= b;
    layer7_outputs(910) <= b;
    layer7_outputs(911) <= not (a or b);
    layer7_outputs(912) <= b;
    layer7_outputs(913) <= a xor b;
    layer7_outputs(914) <= 1'b0;
    layer7_outputs(915) <= not a or b;
    layer7_outputs(916) <= not a;
    layer7_outputs(917) <= b;
    layer7_outputs(918) <= b;
    layer7_outputs(919) <= not (a or b);
    layer7_outputs(920) <= not b;
    layer7_outputs(921) <= a;
    layer7_outputs(922) <= b;
    layer7_outputs(923) <= not b or a;
    layer7_outputs(924) <= not (a or b);
    layer7_outputs(925) <= not (a and b);
    layer7_outputs(926) <= not (a xor b);
    layer7_outputs(927) <= not (a and b);
    layer7_outputs(928) <= b and not a;
    layer7_outputs(929) <= 1'b1;
    layer7_outputs(930) <= b;
    layer7_outputs(931) <= not (a and b);
    layer7_outputs(932) <= not (a xor b);
    layer7_outputs(933) <= not a;
    layer7_outputs(934) <= b;
    layer7_outputs(935) <= not a;
    layer7_outputs(936) <= not b;
    layer7_outputs(937) <= not a;
    layer7_outputs(938) <= b and not a;
    layer7_outputs(939) <= not (a or b);
    layer7_outputs(940) <= not (a and b);
    layer7_outputs(941) <= not b;
    layer7_outputs(942) <= a;
    layer7_outputs(943) <= a;
    layer7_outputs(944) <= not b;
    layer7_outputs(945) <= not b;
    layer7_outputs(946) <= not a or b;
    layer7_outputs(947) <= a and b;
    layer7_outputs(948) <= a;
    layer7_outputs(949) <= not b;
    layer7_outputs(950) <= not a;
    layer7_outputs(951) <= not (a and b);
    layer7_outputs(952) <= not a;
    layer7_outputs(953) <= 1'b0;
    layer7_outputs(954) <= not a;
    layer7_outputs(955) <= a;
    layer7_outputs(956) <= b;
    layer7_outputs(957) <= not b;
    layer7_outputs(958) <= not a or b;
    layer7_outputs(959) <= not (a and b);
    layer7_outputs(960) <= 1'b0;
    layer7_outputs(961) <= not (a and b);
    layer7_outputs(962) <= not (a and b);
    layer7_outputs(963) <= a or b;
    layer7_outputs(964) <= not a or b;
    layer7_outputs(965) <= not (a and b);
    layer7_outputs(966) <= not (a xor b);
    layer7_outputs(967) <= a xor b;
    layer7_outputs(968) <= not (a or b);
    layer7_outputs(969) <= not a;
    layer7_outputs(970) <= not a or b;
    layer7_outputs(971) <= a xor b;
    layer7_outputs(972) <= b;
    layer7_outputs(973) <= a and not b;
    layer7_outputs(974) <= not b;
    layer7_outputs(975) <= b and not a;
    layer7_outputs(976) <= a;
    layer7_outputs(977) <= b;
    layer7_outputs(978) <= not (a xor b);
    layer7_outputs(979) <= not (a xor b);
    layer7_outputs(980) <= not a;
    layer7_outputs(981) <= a xor b;
    layer7_outputs(982) <= not (a xor b);
    layer7_outputs(983) <= not a or b;
    layer7_outputs(984) <= a xor b;
    layer7_outputs(985) <= not a or b;
    layer7_outputs(986) <= not b;
    layer7_outputs(987) <= a;
    layer7_outputs(988) <= a and not b;
    layer7_outputs(989) <= 1'b1;
    layer7_outputs(990) <= a;
    layer7_outputs(991) <= not b;
    layer7_outputs(992) <= not b or a;
    layer7_outputs(993) <= not b or a;
    layer7_outputs(994) <= not (a and b);
    layer7_outputs(995) <= a or b;
    layer7_outputs(996) <= not b;
    layer7_outputs(997) <= not b;
    layer7_outputs(998) <= not a;
    layer7_outputs(999) <= a and b;
    layer7_outputs(1000) <= not (a or b);
    layer7_outputs(1001) <= b;
    layer7_outputs(1002) <= not a or b;
    layer7_outputs(1003) <= not b;
    layer7_outputs(1004) <= not b;
    layer7_outputs(1005) <= not a;
    layer7_outputs(1006) <= a;
    layer7_outputs(1007) <= not a;
    layer7_outputs(1008) <= not b;
    layer7_outputs(1009) <= a;
    layer7_outputs(1010) <= not b or a;
    layer7_outputs(1011) <= not a;
    layer7_outputs(1012) <= not a;
    layer7_outputs(1013) <= a and not b;
    layer7_outputs(1014) <= a;
    layer7_outputs(1015) <= not a;
    layer7_outputs(1016) <= b;
    layer7_outputs(1017) <= a;
    layer7_outputs(1018) <= a;
    layer7_outputs(1019) <= not a;
    layer7_outputs(1020) <= b;
    layer7_outputs(1021) <= not b or a;
    layer7_outputs(1022) <= not (a or b);
    layer7_outputs(1023) <= not (a xor b);
    layer7_outputs(1024) <= a;
    layer7_outputs(1025) <= not (a xor b);
    layer7_outputs(1026) <= not a or b;
    layer7_outputs(1027) <= not a;
    layer7_outputs(1028) <= not a or b;
    layer7_outputs(1029) <= not a;
    layer7_outputs(1030) <= not (a or b);
    layer7_outputs(1031) <= a and not b;
    layer7_outputs(1032) <= not (a and b);
    layer7_outputs(1033) <= a xor b;
    layer7_outputs(1034) <= b;
    layer7_outputs(1035) <= a or b;
    layer7_outputs(1036) <= b;
    layer7_outputs(1037) <= not a or b;
    layer7_outputs(1038) <= not a;
    layer7_outputs(1039) <= not (a xor b);
    layer7_outputs(1040) <= a;
    layer7_outputs(1041) <= not (a xor b);
    layer7_outputs(1042) <= not a;
    layer7_outputs(1043) <= b;
    layer7_outputs(1044) <= not (a and b);
    layer7_outputs(1045) <= not b or a;
    layer7_outputs(1046) <= not (a and b);
    layer7_outputs(1047) <= not a;
    layer7_outputs(1048) <= not (a or b);
    layer7_outputs(1049) <= a or b;
    layer7_outputs(1050) <= not b;
    layer7_outputs(1051) <= 1'b0;
    layer7_outputs(1052) <= b;
    layer7_outputs(1053) <= not b;
    layer7_outputs(1054) <= not a;
    layer7_outputs(1055) <= b and not a;
    layer7_outputs(1056) <= a;
    layer7_outputs(1057) <= b;
    layer7_outputs(1058) <= a and b;
    layer7_outputs(1059) <= b;
    layer7_outputs(1060) <= not a or b;
    layer7_outputs(1061) <= b;
    layer7_outputs(1062) <= b and not a;
    layer7_outputs(1063) <= not a;
    layer7_outputs(1064) <= a;
    layer7_outputs(1065) <= not a or b;
    layer7_outputs(1066) <= not b;
    layer7_outputs(1067) <= not (a xor b);
    layer7_outputs(1068) <= not (a xor b);
    layer7_outputs(1069) <= b and not a;
    layer7_outputs(1070) <= not b;
    layer7_outputs(1071) <= not b;
    layer7_outputs(1072) <= not b;
    layer7_outputs(1073) <= not b;
    layer7_outputs(1074) <= b;
    layer7_outputs(1075) <= not (a xor b);
    layer7_outputs(1076) <= 1'b0;
    layer7_outputs(1077) <= not a;
    layer7_outputs(1078) <= a or b;
    layer7_outputs(1079) <= a and not b;
    layer7_outputs(1080) <= not (a xor b);
    layer7_outputs(1081) <= a and b;
    layer7_outputs(1082) <= not (a or b);
    layer7_outputs(1083) <= b and not a;
    layer7_outputs(1084) <= a;
    layer7_outputs(1085) <= a or b;
    layer7_outputs(1086) <= a;
    layer7_outputs(1087) <= b;
    layer7_outputs(1088) <= a xor b;
    layer7_outputs(1089) <= a;
    layer7_outputs(1090) <= b and not a;
    layer7_outputs(1091) <= a and not b;
    layer7_outputs(1092) <= a xor b;
    layer7_outputs(1093) <= a xor b;
    layer7_outputs(1094) <= b and not a;
    layer7_outputs(1095) <= not b;
    layer7_outputs(1096) <= not b;
    layer7_outputs(1097) <= not b or a;
    layer7_outputs(1098) <= not (a or b);
    layer7_outputs(1099) <= a and not b;
    layer7_outputs(1100) <= a xor b;
    layer7_outputs(1101) <= a;
    layer7_outputs(1102) <= a and b;
    layer7_outputs(1103) <= not b or a;
    layer7_outputs(1104) <= a and not b;
    layer7_outputs(1105) <= a or b;
    layer7_outputs(1106) <= not b or a;
    layer7_outputs(1107) <= not (a xor b);
    layer7_outputs(1108) <= not (a or b);
    layer7_outputs(1109) <= not (a xor b);
    layer7_outputs(1110) <= b and not a;
    layer7_outputs(1111) <= not (a xor b);
    layer7_outputs(1112) <= not b;
    layer7_outputs(1113) <= not a;
    layer7_outputs(1114) <= a;
    layer7_outputs(1115) <= not a;
    layer7_outputs(1116) <= 1'b0;
    layer7_outputs(1117) <= not a;
    layer7_outputs(1118) <= a;
    layer7_outputs(1119) <= b;
    layer7_outputs(1120) <= b;
    layer7_outputs(1121) <= not a;
    layer7_outputs(1122) <= not a;
    layer7_outputs(1123) <= not (a and b);
    layer7_outputs(1124) <= a and not b;
    layer7_outputs(1125) <= a and b;
    layer7_outputs(1126) <= not b;
    layer7_outputs(1127) <= a and not b;
    layer7_outputs(1128) <= a or b;
    layer7_outputs(1129) <= not b or a;
    layer7_outputs(1130) <= a;
    layer7_outputs(1131) <= a or b;
    layer7_outputs(1132) <= a;
    layer7_outputs(1133) <= not a;
    layer7_outputs(1134) <= not b;
    layer7_outputs(1135) <= not a or b;
    layer7_outputs(1136) <= 1'b0;
    layer7_outputs(1137) <= 1'b0;
    layer7_outputs(1138) <= a xor b;
    layer7_outputs(1139) <= not (a and b);
    layer7_outputs(1140) <= not (a and b);
    layer7_outputs(1141) <= not a;
    layer7_outputs(1142) <= not a or b;
    layer7_outputs(1143) <= not a;
    layer7_outputs(1144) <= not (a xor b);
    layer7_outputs(1145) <= 1'b0;
    layer7_outputs(1146) <= not a or b;
    layer7_outputs(1147) <= a xor b;
    layer7_outputs(1148) <= b and not a;
    layer7_outputs(1149) <= a and not b;
    layer7_outputs(1150) <= b;
    layer7_outputs(1151) <= b;
    layer7_outputs(1152) <= b;
    layer7_outputs(1153) <= b and not a;
    layer7_outputs(1154) <= not (a or b);
    layer7_outputs(1155) <= not (a or b);
    layer7_outputs(1156) <= b and not a;
    layer7_outputs(1157) <= not a;
    layer7_outputs(1158) <= b and not a;
    layer7_outputs(1159) <= not a;
    layer7_outputs(1160) <= a and b;
    layer7_outputs(1161) <= not b;
    layer7_outputs(1162) <= not (a and b);
    layer7_outputs(1163) <= not b;
    layer7_outputs(1164) <= b;
    layer7_outputs(1165) <= not a;
    layer7_outputs(1166) <= a;
    layer7_outputs(1167) <= a;
    layer7_outputs(1168) <= not b;
    layer7_outputs(1169) <= not a;
    layer7_outputs(1170) <= a and not b;
    layer7_outputs(1171) <= a and b;
    layer7_outputs(1172) <= not (a xor b);
    layer7_outputs(1173) <= not (a and b);
    layer7_outputs(1174) <= a xor b;
    layer7_outputs(1175) <= not b or a;
    layer7_outputs(1176) <= not (a and b);
    layer7_outputs(1177) <= a and b;
    layer7_outputs(1178) <= not b or a;
    layer7_outputs(1179) <= a and b;
    layer7_outputs(1180) <= not b or a;
    layer7_outputs(1181) <= not b;
    layer7_outputs(1182) <= a and b;
    layer7_outputs(1183) <= a and b;
    layer7_outputs(1184) <= b;
    layer7_outputs(1185) <= a;
    layer7_outputs(1186) <= not b;
    layer7_outputs(1187) <= not (a and b);
    layer7_outputs(1188) <= not b;
    layer7_outputs(1189) <= not (a xor b);
    layer7_outputs(1190) <= not a;
    layer7_outputs(1191) <= not a;
    layer7_outputs(1192) <= b and not a;
    layer7_outputs(1193) <= a xor b;
    layer7_outputs(1194) <= b;
    layer7_outputs(1195) <= b;
    layer7_outputs(1196) <= not a;
    layer7_outputs(1197) <= b and not a;
    layer7_outputs(1198) <= a and b;
    layer7_outputs(1199) <= not (a or b);
    layer7_outputs(1200) <= a and not b;
    layer7_outputs(1201) <= b and not a;
    layer7_outputs(1202) <= a xor b;
    layer7_outputs(1203) <= not (a or b);
    layer7_outputs(1204) <= a and b;
    layer7_outputs(1205) <= not a;
    layer7_outputs(1206) <= not (a or b);
    layer7_outputs(1207) <= not a;
    layer7_outputs(1208) <= a and not b;
    layer7_outputs(1209) <= b and not a;
    layer7_outputs(1210) <= not a;
    layer7_outputs(1211) <= a and not b;
    layer7_outputs(1212) <= a;
    layer7_outputs(1213) <= b;
    layer7_outputs(1214) <= b and not a;
    layer7_outputs(1215) <= not b;
    layer7_outputs(1216) <= a and b;
    layer7_outputs(1217) <= not a;
    layer7_outputs(1218) <= b;
    layer7_outputs(1219) <= b and not a;
    layer7_outputs(1220) <= not b;
    layer7_outputs(1221) <= not b;
    layer7_outputs(1222) <= not (a xor b);
    layer7_outputs(1223) <= not a or b;
    layer7_outputs(1224) <= a or b;
    layer7_outputs(1225) <= not a;
    layer7_outputs(1226) <= not b;
    layer7_outputs(1227) <= not b;
    layer7_outputs(1228) <= a and b;
    layer7_outputs(1229) <= not (a xor b);
    layer7_outputs(1230) <= a and not b;
    layer7_outputs(1231) <= not a or b;
    layer7_outputs(1232) <= not (a or b);
    layer7_outputs(1233) <= not a;
    layer7_outputs(1234) <= b;
    layer7_outputs(1235) <= a and not b;
    layer7_outputs(1236) <= a;
    layer7_outputs(1237) <= not (a or b);
    layer7_outputs(1238) <= a and b;
    layer7_outputs(1239) <= a;
    layer7_outputs(1240) <= a and b;
    layer7_outputs(1241) <= not a;
    layer7_outputs(1242) <= not (a and b);
    layer7_outputs(1243) <= not a;
    layer7_outputs(1244) <= not (a or b);
    layer7_outputs(1245) <= not (a and b);
    layer7_outputs(1246) <= not (a or b);
    layer7_outputs(1247) <= a;
    layer7_outputs(1248) <= not (a xor b);
    layer7_outputs(1249) <= not a;
    layer7_outputs(1250) <= b and not a;
    layer7_outputs(1251) <= a and b;
    layer7_outputs(1252) <= not a;
    layer7_outputs(1253) <= not a;
    layer7_outputs(1254) <= not b;
    layer7_outputs(1255) <= not (a or b);
    layer7_outputs(1256) <= not a;
    layer7_outputs(1257) <= a;
    layer7_outputs(1258) <= not b;
    layer7_outputs(1259) <= b;
    layer7_outputs(1260) <= a xor b;
    layer7_outputs(1261) <= a and b;
    layer7_outputs(1262) <= a and b;
    layer7_outputs(1263) <= a and b;
    layer7_outputs(1264) <= not a;
    layer7_outputs(1265) <= not (a xor b);
    layer7_outputs(1266) <= not a or b;
    layer7_outputs(1267) <= b;
    layer7_outputs(1268) <= a xor b;
    layer7_outputs(1269) <= not b;
    layer7_outputs(1270) <= a xor b;
    layer7_outputs(1271) <= not a;
    layer7_outputs(1272) <= not a;
    layer7_outputs(1273) <= not b or a;
    layer7_outputs(1274) <= a;
    layer7_outputs(1275) <= b;
    layer7_outputs(1276) <= a xor b;
    layer7_outputs(1277) <= not a or b;
    layer7_outputs(1278) <= not a or b;
    layer7_outputs(1279) <= not (a and b);
    layer7_outputs(1280) <= a;
    layer7_outputs(1281) <= not b;
    layer7_outputs(1282) <= a or b;
    layer7_outputs(1283) <= a;
    layer7_outputs(1284) <= b;
    layer7_outputs(1285) <= a;
    layer7_outputs(1286) <= a xor b;
    layer7_outputs(1287) <= not b;
    layer7_outputs(1288) <= not a or b;
    layer7_outputs(1289) <= not b or a;
    layer7_outputs(1290) <= not b;
    layer7_outputs(1291) <= a;
    layer7_outputs(1292) <= a xor b;
    layer7_outputs(1293) <= a and not b;
    layer7_outputs(1294) <= not (a or b);
    layer7_outputs(1295) <= not (a xor b);
    layer7_outputs(1296) <= not (a or b);
    layer7_outputs(1297) <= a and b;
    layer7_outputs(1298) <= a;
    layer7_outputs(1299) <= a or b;
    layer7_outputs(1300) <= not a;
    layer7_outputs(1301) <= not (a and b);
    layer7_outputs(1302) <= a and b;
    layer7_outputs(1303) <= a and b;
    layer7_outputs(1304) <= not a;
    layer7_outputs(1305) <= a;
    layer7_outputs(1306) <= a or b;
    layer7_outputs(1307) <= a;
    layer7_outputs(1308) <= not b;
    layer7_outputs(1309) <= a and not b;
    layer7_outputs(1310) <= a and not b;
    layer7_outputs(1311) <= not b;
    layer7_outputs(1312) <= not a;
    layer7_outputs(1313) <= 1'b0;
    layer7_outputs(1314) <= not a;
    layer7_outputs(1315) <= not a or b;
    layer7_outputs(1316) <= a;
    layer7_outputs(1317) <= a;
    layer7_outputs(1318) <= a and not b;
    layer7_outputs(1319) <= a;
    layer7_outputs(1320) <= a;
    layer7_outputs(1321) <= not b;
    layer7_outputs(1322) <= a or b;
    layer7_outputs(1323) <= not a or b;
    layer7_outputs(1324) <= not a;
    layer7_outputs(1325) <= b and not a;
    layer7_outputs(1326) <= not (a or b);
    layer7_outputs(1327) <= b;
    layer7_outputs(1328) <= not (a or b);
    layer7_outputs(1329) <= b and not a;
    layer7_outputs(1330) <= not a or b;
    layer7_outputs(1331) <= not a or b;
    layer7_outputs(1332) <= a;
    layer7_outputs(1333) <= b;
    layer7_outputs(1334) <= not (a xor b);
    layer7_outputs(1335) <= a and not b;
    layer7_outputs(1336) <= not (a or b);
    layer7_outputs(1337) <= a;
    layer7_outputs(1338) <= not a or b;
    layer7_outputs(1339) <= not a or b;
    layer7_outputs(1340) <= a;
    layer7_outputs(1341) <= not a or b;
    layer7_outputs(1342) <= a and not b;
    layer7_outputs(1343) <= not b;
    layer7_outputs(1344) <= a and not b;
    layer7_outputs(1345) <= not (a and b);
    layer7_outputs(1346) <= a;
    layer7_outputs(1347) <= a;
    layer7_outputs(1348) <= not b;
    layer7_outputs(1349) <= not (a and b);
    layer7_outputs(1350) <= a xor b;
    layer7_outputs(1351) <= b and not a;
    layer7_outputs(1352) <= not a;
    layer7_outputs(1353) <= not (a and b);
    layer7_outputs(1354) <= a;
    layer7_outputs(1355) <= not (a and b);
    layer7_outputs(1356) <= a or b;
    layer7_outputs(1357) <= a;
    layer7_outputs(1358) <= b;
    layer7_outputs(1359) <= not (a or b);
    layer7_outputs(1360) <= a;
    layer7_outputs(1361) <= not a;
    layer7_outputs(1362) <= not a;
    layer7_outputs(1363) <= a;
    layer7_outputs(1364) <= not (a or b);
    layer7_outputs(1365) <= b;
    layer7_outputs(1366) <= 1'b0;
    layer7_outputs(1367) <= not (a and b);
    layer7_outputs(1368) <= not (a or b);
    layer7_outputs(1369) <= a;
    layer7_outputs(1370) <= b;
    layer7_outputs(1371) <= not a;
    layer7_outputs(1372) <= not b;
    layer7_outputs(1373) <= not b or a;
    layer7_outputs(1374) <= a;
    layer7_outputs(1375) <= not (a xor b);
    layer7_outputs(1376) <= not (a and b);
    layer7_outputs(1377) <= a;
    layer7_outputs(1378) <= a or b;
    layer7_outputs(1379) <= b and not a;
    layer7_outputs(1380) <= not b;
    layer7_outputs(1381) <= not a;
    layer7_outputs(1382) <= not a or b;
    layer7_outputs(1383) <= a and not b;
    layer7_outputs(1384) <= a;
    layer7_outputs(1385) <= not a;
    layer7_outputs(1386) <= not b or a;
    layer7_outputs(1387) <= b;
    layer7_outputs(1388) <= not (a and b);
    layer7_outputs(1389) <= not b or a;
    layer7_outputs(1390) <= b;
    layer7_outputs(1391) <= not b or a;
    layer7_outputs(1392) <= 1'b1;
    layer7_outputs(1393) <= not a or b;
    layer7_outputs(1394) <= not b;
    layer7_outputs(1395) <= a and b;
    layer7_outputs(1396) <= a xor b;
    layer7_outputs(1397) <= a xor b;
    layer7_outputs(1398) <= b;
    layer7_outputs(1399) <= a or b;
    layer7_outputs(1400) <= not a;
    layer7_outputs(1401) <= not (a xor b);
    layer7_outputs(1402) <= b;
    layer7_outputs(1403) <= not b;
    layer7_outputs(1404) <= a and b;
    layer7_outputs(1405) <= not b;
    layer7_outputs(1406) <= not (a or b);
    layer7_outputs(1407) <= not b;
    layer7_outputs(1408) <= not a or b;
    layer7_outputs(1409) <= a and b;
    layer7_outputs(1410) <= not a;
    layer7_outputs(1411) <= not a;
    layer7_outputs(1412) <= not b or a;
    layer7_outputs(1413) <= not b or a;
    layer7_outputs(1414) <= a or b;
    layer7_outputs(1415) <= b;
    layer7_outputs(1416) <= b;
    layer7_outputs(1417) <= b and not a;
    layer7_outputs(1418) <= not a;
    layer7_outputs(1419) <= a and b;
    layer7_outputs(1420) <= b;
    layer7_outputs(1421) <= not (a xor b);
    layer7_outputs(1422) <= a;
    layer7_outputs(1423) <= not b or a;
    layer7_outputs(1424) <= a;
    layer7_outputs(1425) <= not a;
    layer7_outputs(1426) <= not b or a;
    layer7_outputs(1427) <= a;
    layer7_outputs(1428) <= not b or a;
    layer7_outputs(1429) <= not b;
    layer7_outputs(1430) <= not b;
    layer7_outputs(1431) <= a and not b;
    layer7_outputs(1432) <= 1'b1;
    layer7_outputs(1433) <= not a or b;
    layer7_outputs(1434) <= b;
    layer7_outputs(1435) <= a and b;
    layer7_outputs(1436) <= not b;
    layer7_outputs(1437) <= a and not b;
    layer7_outputs(1438) <= a and not b;
    layer7_outputs(1439) <= not b;
    layer7_outputs(1440) <= not (a and b);
    layer7_outputs(1441) <= b and not a;
    layer7_outputs(1442) <= not a;
    layer7_outputs(1443) <= a xor b;
    layer7_outputs(1444) <= not a;
    layer7_outputs(1445) <= b;
    layer7_outputs(1446) <= 1'b0;
    layer7_outputs(1447) <= a;
    layer7_outputs(1448) <= a;
    layer7_outputs(1449) <= not a or b;
    layer7_outputs(1450) <= not a;
    layer7_outputs(1451) <= not a or b;
    layer7_outputs(1452) <= not (a xor b);
    layer7_outputs(1453) <= not b;
    layer7_outputs(1454) <= a and not b;
    layer7_outputs(1455) <= not a;
    layer7_outputs(1456) <= a and not b;
    layer7_outputs(1457) <= not b;
    layer7_outputs(1458) <= not a;
    layer7_outputs(1459) <= 1'b0;
    layer7_outputs(1460) <= a or b;
    layer7_outputs(1461) <= b;
    layer7_outputs(1462) <= not b or a;
    layer7_outputs(1463) <= a;
    layer7_outputs(1464) <= not b;
    layer7_outputs(1465) <= b and not a;
    layer7_outputs(1466) <= not a;
    layer7_outputs(1467) <= not a;
    layer7_outputs(1468) <= not a;
    layer7_outputs(1469) <= not a;
    layer7_outputs(1470) <= not (a xor b);
    layer7_outputs(1471) <= a xor b;
    layer7_outputs(1472) <= not a;
    layer7_outputs(1473) <= b;
    layer7_outputs(1474) <= not b;
    layer7_outputs(1475) <= a or b;
    layer7_outputs(1476) <= not a;
    layer7_outputs(1477) <= not b;
    layer7_outputs(1478) <= a or b;
    layer7_outputs(1479) <= 1'b0;
    layer7_outputs(1480) <= a or b;
    layer7_outputs(1481) <= not (a and b);
    layer7_outputs(1482) <= a;
    layer7_outputs(1483) <= a xor b;
    layer7_outputs(1484) <= b;
    layer7_outputs(1485) <= a;
    layer7_outputs(1486) <= a and b;
    layer7_outputs(1487) <= a;
    layer7_outputs(1488) <= not (a xor b);
    layer7_outputs(1489) <= a or b;
    layer7_outputs(1490) <= not (a xor b);
    layer7_outputs(1491) <= a and not b;
    layer7_outputs(1492) <= a and b;
    layer7_outputs(1493) <= not (a and b);
    layer7_outputs(1494) <= b;
    layer7_outputs(1495) <= a and b;
    layer7_outputs(1496) <= b and not a;
    layer7_outputs(1497) <= a or b;
    layer7_outputs(1498) <= not b or a;
    layer7_outputs(1499) <= not a or b;
    layer7_outputs(1500) <= not a or b;
    layer7_outputs(1501) <= not b;
    layer7_outputs(1502) <= not b or a;
    layer7_outputs(1503) <= not b or a;
    layer7_outputs(1504) <= a;
    layer7_outputs(1505) <= a or b;
    layer7_outputs(1506) <= not (a xor b);
    layer7_outputs(1507) <= a and b;
    layer7_outputs(1508) <= a;
    layer7_outputs(1509) <= a;
    layer7_outputs(1510) <= not b or a;
    layer7_outputs(1511) <= not b or a;
    layer7_outputs(1512) <= b and not a;
    layer7_outputs(1513) <= a;
    layer7_outputs(1514) <= not (a and b);
    layer7_outputs(1515) <= not b;
    layer7_outputs(1516) <= a;
    layer7_outputs(1517) <= not b or a;
    layer7_outputs(1518) <= not (a or b);
    layer7_outputs(1519) <= 1'b1;
    layer7_outputs(1520) <= a xor b;
    layer7_outputs(1521) <= not b;
    layer7_outputs(1522) <= b;
    layer7_outputs(1523) <= not (a or b);
    layer7_outputs(1524) <= a or b;
    layer7_outputs(1525) <= a;
    layer7_outputs(1526) <= not a or b;
    layer7_outputs(1527) <= not (a and b);
    layer7_outputs(1528) <= a;
    layer7_outputs(1529) <= a or b;
    layer7_outputs(1530) <= b;
    layer7_outputs(1531) <= 1'b1;
    layer7_outputs(1532) <= a;
    layer7_outputs(1533) <= a;
    layer7_outputs(1534) <= not b or a;
    layer7_outputs(1535) <= a and not b;
    layer7_outputs(1536) <= 1'b0;
    layer7_outputs(1537) <= not a;
    layer7_outputs(1538) <= a;
    layer7_outputs(1539) <= a;
    layer7_outputs(1540) <= not b;
    layer7_outputs(1541) <= a and b;
    layer7_outputs(1542) <= a;
    layer7_outputs(1543) <= a;
    layer7_outputs(1544) <= not b or a;
    layer7_outputs(1545) <= not b;
    layer7_outputs(1546) <= not b;
    layer7_outputs(1547) <= not (a xor b);
    layer7_outputs(1548) <= not a or b;
    layer7_outputs(1549) <= 1'b1;
    layer7_outputs(1550) <= not b or a;
    layer7_outputs(1551) <= not b or a;
    layer7_outputs(1552) <= a;
    layer7_outputs(1553) <= not (a and b);
    layer7_outputs(1554) <= not b;
    layer7_outputs(1555) <= not a;
    layer7_outputs(1556) <= not a;
    layer7_outputs(1557) <= a and not b;
    layer7_outputs(1558) <= not a or b;
    layer7_outputs(1559) <= not b;
    layer7_outputs(1560) <= b and not a;
    layer7_outputs(1561) <= not (a or b);
    layer7_outputs(1562) <= a and not b;
    layer7_outputs(1563) <= a and not b;
    layer7_outputs(1564) <= a and b;
    layer7_outputs(1565) <= a;
    layer7_outputs(1566) <= b and not a;
    layer7_outputs(1567) <= not a or b;
    layer7_outputs(1568) <= b;
    layer7_outputs(1569) <= not (a and b);
    layer7_outputs(1570) <= a and not b;
    layer7_outputs(1571) <= not (a and b);
    layer7_outputs(1572) <= not (a or b);
    layer7_outputs(1573) <= not (a xor b);
    layer7_outputs(1574) <= a and not b;
    layer7_outputs(1575) <= b;
    layer7_outputs(1576) <= b;
    layer7_outputs(1577) <= a;
    layer7_outputs(1578) <= a and b;
    layer7_outputs(1579) <= a and not b;
    layer7_outputs(1580) <= not b;
    layer7_outputs(1581) <= a or b;
    layer7_outputs(1582) <= b and not a;
    layer7_outputs(1583) <= b;
    layer7_outputs(1584) <= not (a and b);
    layer7_outputs(1585) <= not b;
    layer7_outputs(1586) <= not (a xor b);
    layer7_outputs(1587) <= b;
    layer7_outputs(1588) <= not b;
    layer7_outputs(1589) <= not (a and b);
    layer7_outputs(1590) <= a and b;
    layer7_outputs(1591) <= b;
    layer7_outputs(1592) <= a xor b;
    layer7_outputs(1593) <= a;
    layer7_outputs(1594) <= not a;
    layer7_outputs(1595) <= not b;
    layer7_outputs(1596) <= a xor b;
    layer7_outputs(1597) <= not b;
    layer7_outputs(1598) <= a and b;
    layer7_outputs(1599) <= a;
    layer7_outputs(1600) <= b;
    layer7_outputs(1601) <= 1'b1;
    layer7_outputs(1602) <= b;
    layer7_outputs(1603) <= not b;
    layer7_outputs(1604) <= a;
    layer7_outputs(1605) <= a;
    layer7_outputs(1606) <= a or b;
    layer7_outputs(1607) <= a;
    layer7_outputs(1608) <= not (a and b);
    layer7_outputs(1609) <= not (a and b);
    layer7_outputs(1610) <= not (a xor b);
    layer7_outputs(1611) <= b;
    layer7_outputs(1612) <= not b;
    layer7_outputs(1613) <= not a;
    layer7_outputs(1614) <= not a;
    layer7_outputs(1615) <= not b;
    layer7_outputs(1616) <= not a;
    layer7_outputs(1617) <= not a;
    layer7_outputs(1618) <= not b;
    layer7_outputs(1619) <= b and not a;
    layer7_outputs(1620) <= not (a and b);
    layer7_outputs(1621) <= a;
    layer7_outputs(1622) <= not a;
    layer7_outputs(1623) <= not b;
    layer7_outputs(1624) <= b;
    layer7_outputs(1625) <= not b;
    layer7_outputs(1626) <= a xor b;
    layer7_outputs(1627) <= not (a xor b);
    layer7_outputs(1628) <= not b;
    layer7_outputs(1629) <= 1'b1;
    layer7_outputs(1630) <= a and b;
    layer7_outputs(1631) <= a;
    layer7_outputs(1632) <= a and b;
    layer7_outputs(1633) <= not (a or b);
    layer7_outputs(1634) <= b;
    layer7_outputs(1635) <= a;
    layer7_outputs(1636) <= not (a and b);
    layer7_outputs(1637) <= b;
    layer7_outputs(1638) <= not b or a;
    layer7_outputs(1639) <= b;
    layer7_outputs(1640) <= not a or b;
    layer7_outputs(1641) <= a and not b;
    layer7_outputs(1642) <= not (a and b);
    layer7_outputs(1643) <= not (a xor b);
    layer7_outputs(1644) <= not b or a;
    layer7_outputs(1645) <= b and not a;
    layer7_outputs(1646) <= not b;
    layer7_outputs(1647) <= not b;
    layer7_outputs(1648) <= b;
    layer7_outputs(1649) <= not b;
    layer7_outputs(1650) <= a or b;
    layer7_outputs(1651) <= b and not a;
    layer7_outputs(1652) <= not (a and b);
    layer7_outputs(1653) <= b;
    layer7_outputs(1654) <= not (a or b);
    layer7_outputs(1655) <= b and not a;
    layer7_outputs(1656) <= a xor b;
    layer7_outputs(1657) <= not (a and b);
    layer7_outputs(1658) <= a or b;
    layer7_outputs(1659) <= a and not b;
    layer7_outputs(1660) <= not b or a;
    layer7_outputs(1661) <= a and b;
    layer7_outputs(1662) <= b;
    layer7_outputs(1663) <= not a or b;
    layer7_outputs(1664) <= not (a xor b);
    layer7_outputs(1665) <= b and not a;
    layer7_outputs(1666) <= b;
    layer7_outputs(1667) <= b and not a;
    layer7_outputs(1668) <= not b;
    layer7_outputs(1669) <= not a or b;
    layer7_outputs(1670) <= not (a xor b);
    layer7_outputs(1671) <= not a;
    layer7_outputs(1672) <= not a;
    layer7_outputs(1673) <= b;
    layer7_outputs(1674) <= not a;
    layer7_outputs(1675) <= a;
    layer7_outputs(1676) <= not a;
    layer7_outputs(1677) <= a xor b;
    layer7_outputs(1678) <= not b or a;
    layer7_outputs(1679) <= not (a xor b);
    layer7_outputs(1680) <= not b;
    layer7_outputs(1681) <= not b;
    layer7_outputs(1682) <= a and b;
    layer7_outputs(1683) <= not (a xor b);
    layer7_outputs(1684) <= not b;
    layer7_outputs(1685) <= not b;
    layer7_outputs(1686) <= a and not b;
    layer7_outputs(1687) <= a and b;
    layer7_outputs(1688) <= not a;
    layer7_outputs(1689) <= not b;
    layer7_outputs(1690) <= not a;
    layer7_outputs(1691) <= a or b;
    layer7_outputs(1692) <= a;
    layer7_outputs(1693) <= not (a xor b);
    layer7_outputs(1694) <= a and b;
    layer7_outputs(1695) <= a or b;
    layer7_outputs(1696) <= a;
    layer7_outputs(1697) <= not a;
    layer7_outputs(1698) <= not (a xor b);
    layer7_outputs(1699) <= a or b;
    layer7_outputs(1700) <= b;
    layer7_outputs(1701) <= not (a and b);
    layer7_outputs(1702) <= b;
    layer7_outputs(1703) <= not a;
    layer7_outputs(1704) <= a;
    layer7_outputs(1705) <= b;
    layer7_outputs(1706) <= not (a xor b);
    layer7_outputs(1707) <= not b;
    layer7_outputs(1708) <= not a or b;
    layer7_outputs(1709) <= not b;
    layer7_outputs(1710) <= a xor b;
    layer7_outputs(1711) <= a xor b;
    layer7_outputs(1712) <= a xor b;
    layer7_outputs(1713) <= 1'b1;
    layer7_outputs(1714) <= a or b;
    layer7_outputs(1715) <= a or b;
    layer7_outputs(1716) <= b;
    layer7_outputs(1717) <= b and not a;
    layer7_outputs(1718) <= b;
    layer7_outputs(1719) <= not (a and b);
    layer7_outputs(1720) <= b;
    layer7_outputs(1721) <= b;
    layer7_outputs(1722) <= b and not a;
    layer7_outputs(1723) <= b;
    layer7_outputs(1724) <= a;
    layer7_outputs(1725) <= 1'b0;
    layer7_outputs(1726) <= a xor b;
    layer7_outputs(1727) <= a and not b;
    layer7_outputs(1728) <= 1'b0;
    layer7_outputs(1729) <= b;
    layer7_outputs(1730) <= b and not a;
    layer7_outputs(1731) <= b;
    layer7_outputs(1732) <= a and not b;
    layer7_outputs(1733) <= a;
    layer7_outputs(1734) <= not a;
    layer7_outputs(1735) <= a;
    layer7_outputs(1736) <= b;
    layer7_outputs(1737) <= not (a and b);
    layer7_outputs(1738) <= a and not b;
    layer7_outputs(1739) <= b;
    layer7_outputs(1740) <= not b;
    layer7_outputs(1741) <= a;
    layer7_outputs(1742) <= a and not b;
    layer7_outputs(1743) <= not (a or b);
    layer7_outputs(1744) <= a and not b;
    layer7_outputs(1745) <= not (a and b);
    layer7_outputs(1746) <= a;
    layer7_outputs(1747) <= not b or a;
    layer7_outputs(1748) <= not (a or b);
    layer7_outputs(1749) <= 1'b0;
    layer7_outputs(1750) <= a xor b;
    layer7_outputs(1751) <= b and not a;
    layer7_outputs(1752) <= a;
    layer7_outputs(1753) <= a or b;
    layer7_outputs(1754) <= a xor b;
    layer7_outputs(1755) <= a;
    layer7_outputs(1756) <= b and not a;
    layer7_outputs(1757) <= a;
    layer7_outputs(1758) <= not a;
    layer7_outputs(1759) <= not (a and b);
    layer7_outputs(1760) <= not a;
    layer7_outputs(1761) <= not b;
    layer7_outputs(1762) <= not b or a;
    layer7_outputs(1763) <= not b or a;
    layer7_outputs(1764) <= b and not a;
    layer7_outputs(1765) <= not (a xor b);
    layer7_outputs(1766) <= not a;
    layer7_outputs(1767) <= 1'b1;
    layer7_outputs(1768) <= a xor b;
    layer7_outputs(1769) <= not a;
    layer7_outputs(1770) <= not (a and b);
    layer7_outputs(1771) <= a;
    layer7_outputs(1772) <= not b;
    layer7_outputs(1773) <= not b;
    layer7_outputs(1774) <= a xor b;
    layer7_outputs(1775) <= b and not a;
    layer7_outputs(1776) <= a and b;
    layer7_outputs(1777) <= not a;
    layer7_outputs(1778) <= a and b;
    layer7_outputs(1779) <= a or b;
    layer7_outputs(1780) <= not (a xor b);
    layer7_outputs(1781) <= not a;
    layer7_outputs(1782) <= not (a and b);
    layer7_outputs(1783) <= not b;
    layer7_outputs(1784) <= not (a and b);
    layer7_outputs(1785) <= not b or a;
    layer7_outputs(1786) <= a xor b;
    layer7_outputs(1787) <= not b;
    layer7_outputs(1788) <= not (a or b);
    layer7_outputs(1789) <= not a;
    layer7_outputs(1790) <= not a or b;
    layer7_outputs(1791) <= not b;
    layer7_outputs(1792) <= not (a and b);
    layer7_outputs(1793) <= not a;
    layer7_outputs(1794) <= not a or b;
    layer7_outputs(1795) <= a xor b;
    layer7_outputs(1796) <= not a;
    layer7_outputs(1797) <= b;
    layer7_outputs(1798) <= not b;
    layer7_outputs(1799) <= not b or a;
    layer7_outputs(1800) <= a;
    layer7_outputs(1801) <= not a;
    layer7_outputs(1802) <= not b or a;
    layer7_outputs(1803) <= a or b;
    layer7_outputs(1804) <= a and b;
    layer7_outputs(1805) <= a and not b;
    layer7_outputs(1806) <= not b or a;
    layer7_outputs(1807) <= not a;
    layer7_outputs(1808) <= a xor b;
    layer7_outputs(1809) <= not a;
    layer7_outputs(1810) <= not a;
    layer7_outputs(1811) <= a and b;
    layer7_outputs(1812) <= not a;
    layer7_outputs(1813) <= a;
    layer7_outputs(1814) <= not (a or b);
    layer7_outputs(1815) <= a;
    layer7_outputs(1816) <= not (a or b);
    layer7_outputs(1817) <= b;
    layer7_outputs(1818) <= a or b;
    layer7_outputs(1819) <= not (a or b);
    layer7_outputs(1820) <= not b;
    layer7_outputs(1821) <= a or b;
    layer7_outputs(1822) <= not (a and b);
    layer7_outputs(1823) <= a xor b;
    layer7_outputs(1824) <= not a;
    layer7_outputs(1825) <= not (a or b);
    layer7_outputs(1826) <= b;
    layer7_outputs(1827) <= b;
    layer7_outputs(1828) <= a xor b;
    layer7_outputs(1829) <= b and not a;
    layer7_outputs(1830) <= not (a xor b);
    layer7_outputs(1831) <= b;
    layer7_outputs(1832) <= a or b;
    layer7_outputs(1833) <= b and not a;
    layer7_outputs(1834) <= not b or a;
    layer7_outputs(1835) <= not a;
    layer7_outputs(1836) <= not b;
    layer7_outputs(1837) <= not b;
    layer7_outputs(1838) <= a;
    layer7_outputs(1839) <= not a or b;
    layer7_outputs(1840) <= not a;
    layer7_outputs(1841) <= not b;
    layer7_outputs(1842) <= not (a or b);
    layer7_outputs(1843) <= not (a and b);
    layer7_outputs(1844) <= not a or b;
    layer7_outputs(1845) <= not (a xor b);
    layer7_outputs(1846) <= not b;
    layer7_outputs(1847) <= not a;
    layer7_outputs(1848) <= not (a and b);
    layer7_outputs(1849) <= not (a and b);
    layer7_outputs(1850) <= not b;
    layer7_outputs(1851) <= a and not b;
    layer7_outputs(1852) <= a or b;
    layer7_outputs(1853) <= b and not a;
    layer7_outputs(1854) <= not b;
    layer7_outputs(1855) <= a and b;
    layer7_outputs(1856) <= 1'b1;
    layer7_outputs(1857) <= not a or b;
    layer7_outputs(1858) <= not a;
    layer7_outputs(1859) <= not b or a;
    layer7_outputs(1860) <= not b or a;
    layer7_outputs(1861) <= not (a and b);
    layer7_outputs(1862) <= not (a or b);
    layer7_outputs(1863) <= b;
    layer7_outputs(1864) <= not b;
    layer7_outputs(1865) <= a and not b;
    layer7_outputs(1866) <= not b;
    layer7_outputs(1867) <= not a or b;
    layer7_outputs(1868) <= not a;
    layer7_outputs(1869) <= b;
    layer7_outputs(1870) <= not (a or b);
    layer7_outputs(1871) <= not a;
    layer7_outputs(1872) <= not b;
    layer7_outputs(1873) <= not b or a;
    layer7_outputs(1874) <= not b;
    layer7_outputs(1875) <= not (a or b);
    layer7_outputs(1876) <= b;
    layer7_outputs(1877) <= not a or b;
    layer7_outputs(1878) <= not b or a;
    layer7_outputs(1879) <= not a;
    layer7_outputs(1880) <= 1'b0;
    layer7_outputs(1881) <= not a or b;
    layer7_outputs(1882) <= a and b;
    layer7_outputs(1883) <= not a;
    layer7_outputs(1884) <= b;
    layer7_outputs(1885) <= not a or b;
    layer7_outputs(1886) <= a;
    layer7_outputs(1887) <= not a;
    layer7_outputs(1888) <= not a;
    layer7_outputs(1889) <= a and b;
    layer7_outputs(1890) <= b;
    layer7_outputs(1891) <= a;
    layer7_outputs(1892) <= a;
    layer7_outputs(1893) <= not (a or b);
    layer7_outputs(1894) <= a and not b;
    layer7_outputs(1895) <= a;
    layer7_outputs(1896) <= b;
    layer7_outputs(1897) <= a and b;
    layer7_outputs(1898) <= not (a or b);
    layer7_outputs(1899) <= not (a xor b);
    layer7_outputs(1900) <= not b or a;
    layer7_outputs(1901) <= a;
    layer7_outputs(1902) <= not (a and b);
    layer7_outputs(1903) <= not (a xor b);
    layer7_outputs(1904) <= b;
    layer7_outputs(1905) <= not a or b;
    layer7_outputs(1906) <= not a or b;
    layer7_outputs(1907) <= a and not b;
    layer7_outputs(1908) <= a and b;
    layer7_outputs(1909) <= b;
    layer7_outputs(1910) <= a xor b;
    layer7_outputs(1911) <= a and not b;
    layer7_outputs(1912) <= a and b;
    layer7_outputs(1913) <= not (a or b);
    layer7_outputs(1914) <= not b or a;
    layer7_outputs(1915) <= not (a and b);
    layer7_outputs(1916) <= not b or a;
    layer7_outputs(1917) <= b;
    layer7_outputs(1918) <= b and not a;
    layer7_outputs(1919) <= not (a xor b);
    layer7_outputs(1920) <= b and not a;
    layer7_outputs(1921) <= b;
    layer7_outputs(1922) <= not (a or b);
    layer7_outputs(1923) <= not a;
    layer7_outputs(1924) <= not b;
    layer7_outputs(1925) <= not (a and b);
    layer7_outputs(1926) <= not (a xor b);
    layer7_outputs(1927) <= not a;
    layer7_outputs(1928) <= b;
    layer7_outputs(1929) <= a and b;
    layer7_outputs(1930) <= b;
    layer7_outputs(1931) <= a or b;
    layer7_outputs(1932) <= not (a or b);
    layer7_outputs(1933) <= a;
    layer7_outputs(1934) <= not b or a;
    layer7_outputs(1935) <= not a;
    layer7_outputs(1936) <= a or b;
    layer7_outputs(1937) <= not (a xor b);
    layer7_outputs(1938) <= a and not b;
    layer7_outputs(1939) <= not a or b;
    layer7_outputs(1940) <= not a;
    layer7_outputs(1941) <= not b or a;
    layer7_outputs(1942) <= not b;
    layer7_outputs(1943) <= not a;
    layer7_outputs(1944) <= not a;
    layer7_outputs(1945) <= a xor b;
    layer7_outputs(1946) <= not b or a;
    layer7_outputs(1947) <= not b;
    layer7_outputs(1948) <= b;
    layer7_outputs(1949) <= not b or a;
    layer7_outputs(1950) <= not (a and b);
    layer7_outputs(1951) <= b;
    layer7_outputs(1952) <= a or b;
    layer7_outputs(1953) <= b and not a;
    layer7_outputs(1954) <= a and b;
    layer7_outputs(1955) <= a;
    layer7_outputs(1956) <= not a;
    layer7_outputs(1957) <= a and not b;
    layer7_outputs(1958) <= not b;
    layer7_outputs(1959) <= 1'b1;
    layer7_outputs(1960) <= not (a xor b);
    layer7_outputs(1961) <= b;
    layer7_outputs(1962) <= b;
    layer7_outputs(1963) <= a and not b;
    layer7_outputs(1964) <= not a or b;
    layer7_outputs(1965) <= not (a or b);
    layer7_outputs(1966) <= not b;
    layer7_outputs(1967) <= a and b;
    layer7_outputs(1968) <= not b;
    layer7_outputs(1969) <= not (a and b);
    layer7_outputs(1970) <= not a;
    layer7_outputs(1971) <= not b;
    layer7_outputs(1972) <= not a;
    layer7_outputs(1973) <= a;
    layer7_outputs(1974) <= a;
    layer7_outputs(1975) <= a xor b;
    layer7_outputs(1976) <= a;
    layer7_outputs(1977) <= 1'b0;
    layer7_outputs(1978) <= not b or a;
    layer7_outputs(1979) <= not b;
    layer7_outputs(1980) <= a xor b;
    layer7_outputs(1981) <= a and not b;
    layer7_outputs(1982) <= a xor b;
    layer7_outputs(1983) <= not (a or b);
    layer7_outputs(1984) <= a xor b;
    layer7_outputs(1985) <= a or b;
    layer7_outputs(1986) <= not (a xor b);
    layer7_outputs(1987) <= a and b;
    layer7_outputs(1988) <= a and b;
    layer7_outputs(1989) <= b;
    layer7_outputs(1990) <= not (a or b);
    layer7_outputs(1991) <= not b;
    layer7_outputs(1992) <= b;
    layer7_outputs(1993) <= b and not a;
    layer7_outputs(1994) <= not a;
    layer7_outputs(1995) <= not a;
    layer7_outputs(1996) <= not (a xor b);
    layer7_outputs(1997) <= not (a xor b);
    layer7_outputs(1998) <= b;
    layer7_outputs(1999) <= not b or a;
    layer7_outputs(2000) <= a;
    layer7_outputs(2001) <= a or b;
    layer7_outputs(2002) <= not a;
    layer7_outputs(2003) <= b;
    layer7_outputs(2004) <= b;
    layer7_outputs(2005) <= not (a and b);
    layer7_outputs(2006) <= a xor b;
    layer7_outputs(2007) <= not (a or b);
    layer7_outputs(2008) <= a and not b;
    layer7_outputs(2009) <= not (a or b);
    layer7_outputs(2010) <= not a;
    layer7_outputs(2011) <= a xor b;
    layer7_outputs(2012) <= not b;
    layer7_outputs(2013) <= a and b;
    layer7_outputs(2014) <= not b;
    layer7_outputs(2015) <= a;
    layer7_outputs(2016) <= a and not b;
    layer7_outputs(2017) <= not (a or b);
    layer7_outputs(2018) <= b;
    layer7_outputs(2019) <= not (a xor b);
    layer7_outputs(2020) <= a;
    layer7_outputs(2021) <= a xor b;
    layer7_outputs(2022) <= not a or b;
    layer7_outputs(2023) <= not a;
    layer7_outputs(2024) <= not a or b;
    layer7_outputs(2025) <= not b;
    layer7_outputs(2026) <= a and not b;
    layer7_outputs(2027) <= not a;
    layer7_outputs(2028) <= not b;
    layer7_outputs(2029) <= not b;
    layer7_outputs(2030) <= b and not a;
    layer7_outputs(2031) <= not (a and b);
    layer7_outputs(2032) <= a and b;
    layer7_outputs(2033) <= not b;
    layer7_outputs(2034) <= not b;
    layer7_outputs(2035) <= not a or b;
    layer7_outputs(2036) <= not a or b;
    layer7_outputs(2037) <= not b or a;
    layer7_outputs(2038) <= a and b;
    layer7_outputs(2039) <= b and not a;
    layer7_outputs(2040) <= not b;
    layer7_outputs(2041) <= a xor b;
    layer7_outputs(2042) <= not a;
    layer7_outputs(2043) <= a or b;
    layer7_outputs(2044) <= 1'b1;
    layer7_outputs(2045) <= not (a xor b);
    layer7_outputs(2046) <= b;
    layer7_outputs(2047) <= b;
    layer7_outputs(2048) <= not a;
    layer7_outputs(2049) <= not a;
    layer7_outputs(2050) <= not b;
    layer7_outputs(2051) <= b;
    layer7_outputs(2052) <= a or b;
    layer7_outputs(2053) <= not a;
    layer7_outputs(2054) <= not b;
    layer7_outputs(2055) <= not b;
    layer7_outputs(2056) <= a;
    layer7_outputs(2057) <= 1'b1;
    layer7_outputs(2058) <= not a or b;
    layer7_outputs(2059) <= not (a xor b);
    layer7_outputs(2060) <= a or b;
    layer7_outputs(2061) <= not a;
    layer7_outputs(2062) <= not (a or b);
    layer7_outputs(2063) <= a and b;
    layer7_outputs(2064) <= b;
    layer7_outputs(2065) <= not b;
    layer7_outputs(2066) <= not a;
    layer7_outputs(2067) <= a;
    layer7_outputs(2068) <= a or b;
    layer7_outputs(2069) <= not (a and b);
    layer7_outputs(2070) <= not b;
    layer7_outputs(2071) <= b;
    layer7_outputs(2072) <= not b;
    layer7_outputs(2073) <= not b or a;
    layer7_outputs(2074) <= b and not a;
    layer7_outputs(2075) <= a and b;
    layer7_outputs(2076) <= a or b;
    layer7_outputs(2077) <= not a;
    layer7_outputs(2078) <= a;
    layer7_outputs(2079) <= a and not b;
    layer7_outputs(2080) <= not b;
    layer7_outputs(2081) <= 1'b1;
    layer7_outputs(2082) <= not a or b;
    layer7_outputs(2083) <= a or b;
    layer7_outputs(2084) <= not a;
    layer7_outputs(2085) <= a xor b;
    layer7_outputs(2086) <= a and not b;
    layer7_outputs(2087) <= not b or a;
    layer7_outputs(2088) <= not (a and b);
    layer7_outputs(2089) <= b;
    layer7_outputs(2090) <= 1'b0;
    layer7_outputs(2091) <= a or b;
    layer7_outputs(2092) <= not b or a;
    layer7_outputs(2093) <= not a;
    layer7_outputs(2094) <= not a;
    layer7_outputs(2095) <= a and not b;
    layer7_outputs(2096) <= b;
    layer7_outputs(2097) <= not a;
    layer7_outputs(2098) <= not (a or b);
    layer7_outputs(2099) <= a;
    layer7_outputs(2100) <= a and not b;
    layer7_outputs(2101) <= not a;
    layer7_outputs(2102) <= not b;
    layer7_outputs(2103) <= a;
    layer7_outputs(2104) <= not a;
    layer7_outputs(2105) <= not (a xor b);
    layer7_outputs(2106) <= a xor b;
    layer7_outputs(2107) <= not a or b;
    layer7_outputs(2108) <= not b;
    layer7_outputs(2109) <= not (a xor b);
    layer7_outputs(2110) <= 1'b0;
    layer7_outputs(2111) <= not a;
    layer7_outputs(2112) <= b and not a;
    layer7_outputs(2113) <= not (a or b);
    layer7_outputs(2114) <= not (a xor b);
    layer7_outputs(2115) <= not b or a;
    layer7_outputs(2116) <= a and b;
    layer7_outputs(2117) <= a and b;
    layer7_outputs(2118) <= not (a or b);
    layer7_outputs(2119) <= a or b;
    layer7_outputs(2120) <= not a or b;
    layer7_outputs(2121) <= a;
    layer7_outputs(2122) <= not a;
    layer7_outputs(2123) <= not (a xor b);
    layer7_outputs(2124) <= not a;
    layer7_outputs(2125) <= a and not b;
    layer7_outputs(2126) <= b and not a;
    layer7_outputs(2127) <= not b or a;
    layer7_outputs(2128) <= a;
    layer7_outputs(2129) <= a;
    layer7_outputs(2130) <= not b or a;
    layer7_outputs(2131) <= 1'b1;
    layer7_outputs(2132) <= b;
    layer7_outputs(2133) <= a xor b;
    layer7_outputs(2134) <= a;
    layer7_outputs(2135) <= not a;
    layer7_outputs(2136) <= not (a xor b);
    layer7_outputs(2137) <= b;
    layer7_outputs(2138) <= a;
    layer7_outputs(2139) <= not a or b;
    layer7_outputs(2140) <= not (a or b);
    layer7_outputs(2141) <= a xor b;
    layer7_outputs(2142) <= b;
    layer7_outputs(2143) <= a and b;
    layer7_outputs(2144) <= a xor b;
    layer7_outputs(2145) <= not a;
    layer7_outputs(2146) <= b;
    layer7_outputs(2147) <= not b;
    layer7_outputs(2148) <= not (a xor b);
    layer7_outputs(2149) <= b;
    layer7_outputs(2150) <= b;
    layer7_outputs(2151) <= a xor b;
    layer7_outputs(2152) <= a and b;
    layer7_outputs(2153) <= not b;
    layer7_outputs(2154) <= a;
    layer7_outputs(2155) <= a xor b;
    layer7_outputs(2156) <= not b or a;
    layer7_outputs(2157) <= a and not b;
    layer7_outputs(2158) <= not (a xor b);
    layer7_outputs(2159) <= a and not b;
    layer7_outputs(2160) <= a and b;
    layer7_outputs(2161) <= not (a and b);
    layer7_outputs(2162) <= not b or a;
    layer7_outputs(2163) <= not (a and b);
    layer7_outputs(2164) <= not b;
    layer7_outputs(2165) <= not a or b;
    layer7_outputs(2166) <= b;
    layer7_outputs(2167) <= b;
    layer7_outputs(2168) <= 1'b1;
    layer7_outputs(2169) <= not a;
    layer7_outputs(2170) <= a xor b;
    layer7_outputs(2171) <= not (a and b);
    layer7_outputs(2172) <= not b;
    layer7_outputs(2173) <= not a;
    layer7_outputs(2174) <= a xor b;
    layer7_outputs(2175) <= not (a and b);
    layer7_outputs(2176) <= not b or a;
    layer7_outputs(2177) <= not (a xor b);
    layer7_outputs(2178) <= not (a and b);
    layer7_outputs(2179) <= b and not a;
    layer7_outputs(2180) <= not a or b;
    layer7_outputs(2181) <= a xor b;
    layer7_outputs(2182) <= not a or b;
    layer7_outputs(2183) <= a or b;
    layer7_outputs(2184) <= b;
    layer7_outputs(2185) <= b;
    layer7_outputs(2186) <= a xor b;
    layer7_outputs(2187) <= not b;
    layer7_outputs(2188) <= b;
    layer7_outputs(2189) <= b;
    layer7_outputs(2190) <= a;
    layer7_outputs(2191) <= a;
    layer7_outputs(2192) <= a and b;
    layer7_outputs(2193) <= b;
    layer7_outputs(2194) <= a;
    layer7_outputs(2195) <= a or b;
    layer7_outputs(2196) <= a;
    layer7_outputs(2197) <= a;
    layer7_outputs(2198) <= b;
    layer7_outputs(2199) <= b;
    layer7_outputs(2200) <= not a;
    layer7_outputs(2201) <= a and b;
    layer7_outputs(2202) <= 1'b1;
    layer7_outputs(2203) <= a and not b;
    layer7_outputs(2204) <= not (a or b);
    layer7_outputs(2205) <= not (a and b);
    layer7_outputs(2206) <= not a or b;
    layer7_outputs(2207) <= not (a or b);
    layer7_outputs(2208) <= not (a or b);
    layer7_outputs(2209) <= not (a or b);
    layer7_outputs(2210) <= not a;
    layer7_outputs(2211) <= a xor b;
    layer7_outputs(2212) <= a;
    layer7_outputs(2213) <= a xor b;
    layer7_outputs(2214) <= not b or a;
    layer7_outputs(2215) <= a;
    layer7_outputs(2216) <= not b;
    layer7_outputs(2217) <= not a;
    layer7_outputs(2218) <= not (a or b);
    layer7_outputs(2219) <= b;
    layer7_outputs(2220) <= b;
    layer7_outputs(2221) <= b;
    layer7_outputs(2222) <= not b or a;
    layer7_outputs(2223) <= a xor b;
    layer7_outputs(2224) <= b;
    layer7_outputs(2225) <= b;
    layer7_outputs(2226) <= not (a or b);
    layer7_outputs(2227) <= not b;
    layer7_outputs(2228) <= not (a and b);
    layer7_outputs(2229) <= not (a or b);
    layer7_outputs(2230) <= b;
    layer7_outputs(2231) <= a;
    layer7_outputs(2232) <= not (a or b);
    layer7_outputs(2233) <= 1'b1;
    layer7_outputs(2234) <= not b;
    layer7_outputs(2235) <= a;
    layer7_outputs(2236) <= not a or b;
    layer7_outputs(2237) <= b;
    layer7_outputs(2238) <= a and not b;
    layer7_outputs(2239) <= a xor b;
    layer7_outputs(2240) <= a and not b;
    layer7_outputs(2241) <= not b;
    layer7_outputs(2242) <= not b;
    layer7_outputs(2243) <= not a;
    layer7_outputs(2244) <= not b;
    layer7_outputs(2245) <= not b;
    layer7_outputs(2246) <= not a;
    layer7_outputs(2247) <= not b;
    layer7_outputs(2248) <= a xor b;
    layer7_outputs(2249) <= a;
    layer7_outputs(2250) <= a and not b;
    layer7_outputs(2251) <= a and not b;
    layer7_outputs(2252) <= b;
    layer7_outputs(2253) <= not b or a;
    layer7_outputs(2254) <= not (a and b);
    layer7_outputs(2255) <= not a or b;
    layer7_outputs(2256) <= not a;
    layer7_outputs(2257) <= not (a or b);
    layer7_outputs(2258) <= a and not b;
    layer7_outputs(2259) <= not b or a;
    layer7_outputs(2260) <= not (a and b);
    layer7_outputs(2261) <= not b;
    layer7_outputs(2262) <= a;
    layer7_outputs(2263) <= a and b;
    layer7_outputs(2264) <= not b;
    layer7_outputs(2265) <= not b;
    layer7_outputs(2266) <= b and not a;
    layer7_outputs(2267) <= not b;
    layer7_outputs(2268) <= b and not a;
    layer7_outputs(2269) <= not a or b;
    layer7_outputs(2270) <= not a;
    layer7_outputs(2271) <= not a;
    layer7_outputs(2272) <= not (a and b);
    layer7_outputs(2273) <= a and b;
    layer7_outputs(2274) <= a and not b;
    layer7_outputs(2275) <= not a;
    layer7_outputs(2276) <= b and not a;
    layer7_outputs(2277) <= not b;
    layer7_outputs(2278) <= a;
    layer7_outputs(2279) <= a or b;
    layer7_outputs(2280) <= a;
    layer7_outputs(2281) <= not a;
    layer7_outputs(2282) <= a;
    layer7_outputs(2283) <= not (a xor b);
    layer7_outputs(2284) <= a xor b;
    layer7_outputs(2285) <= not (a or b);
    layer7_outputs(2286) <= not a;
    layer7_outputs(2287) <= not a;
    layer7_outputs(2288) <= b;
    layer7_outputs(2289) <= b and not a;
    layer7_outputs(2290) <= a or b;
    layer7_outputs(2291) <= not (a and b);
    layer7_outputs(2292) <= not a;
    layer7_outputs(2293) <= not (a or b);
    layer7_outputs(2294) <= not a or b;
    layer7_outputs(2295) <= a;
    layer7_outputs(2296) <= not (a and b);
    layer7_outputs(2297) <= a;
    layer7_outputs(2298) <= not b;
    layer7_outputs(2299) <= b;
    layer7_outputs(2300) <= not b;
    layer7_outputs(2301) <= a and b;
    layer7_outputs(2302) <= a;
    layer7_outputs(2303) <= not b;
    layer7_outputs(2304) <= not (a xor b);
    layer7_outputs(2305) <= not (a or b);
    layer7_outputs(2306) <= not a or b;
    layer7_outputs(2307) <= not (a and b);
    layer7_outputs(2308) <= a and not b;
    layer7_outputs(2309) <= a and not b;
    layer7_outputs(2310) <= a;
    layer7_outputs(2311) <= a xor b;
    layer7_outputs(2312) <= not b;
    layer7_outputs(2313) <= not (a xor b);
    layer7_outputs(2314) <= b;
    layer7_outputs(2315) <= a;
    layer7_outputs(2316) <= a and not b;
    layer7_outputs(2317) <= not b;
    layer7_outputs(2318) <= a or b;
    layer7_outputs(2319) <= a and b;
    layer7_outputs(2320) <= not b;
    layer7_outputs(2321) <= not a;
    layer7_outputs(2322) <= b;
    layer7_outputs(2323) <= not a or b;
    layer7_outputs(2324) <= not b;
    layer7_outputs(2325) <= b;
    layer7_outputs(2326) <= b;
    layer7_outputs(2327) <= a;
    layer7_outputs(2328) <= a;
    layer7_outputs(2329) <= not a or b;
    layer7_outputs(2330) <= a and not b;
    layer7_outputs(2331) <= a;
    layer7_outputs(2332) <= not (a and b);
    layer7_outputs(2333) <= a or b;
    layer7_outputs(2334) <= not (a xor b);
    layer7_outputs(2335) <= not (a xor b);
    layer7_outputs(2336) <= a;
    layer7_outputs(2337) <= not a;
    layer7_outputs(2338) <= not (a and b);
    layer7_outputs(2339) <= not (a and b);
    layer7_outputs(2340) <= not b or a;
    layer7_outputs(2341) <= a and b;
    layer7_outputs(2342) <= not a;
    layer7_outputs(2343) <= not a;
    layer7_outputs(2344) <= b;
    layer7_outputs(2345) <= not a;
    layer7_outputs(2346) <= b;
    layer7_outputs(2347) <= not b;
    layer7_outputs(2348) <= not (a and b);
    layer7_outputs(2349) <= not a;
    layer7_outputs(2350) <= b and not a;
    layer7_outputs(2351) <= not a or b;
    layer7_outputs(2352) <= not b;
    layer7_outputs(2353) <= a and not b;
    layer7_outputs(2354) <= not b;
    layer7_outputs(2355) <= not (a xor b);
    layer7_outputs(2356) <= not (a or b);
    layer7_outputs(2357) <= not a or b;
    layer7_outputs(2358) <= b;
    layer7_outputs(2359) <= not (a xor b);
    layer7_outputs(2360) <= not a;
    layer7_outputs(2361) <= not b;
    layer7_outputs(2362) <= not a;
    layer7_outputs(2363) <= a;
    layer7_outputs(2364) <= not a;
    layer7_outputs(2365) <= 1'b0;
    layer7_outputs(2366) <= a;
    layer7_outputs(2367) <= b;
    layer7_outputs(2368) <= not a or b;
    layer7_outputs(2369) <= a and b;
    layer7_outputs(2370) <= not a;
    layer7_outputs(2371) <= b;
    layer7_outputs(2372) <= not a;
    layer7_outputs(2373) <= not (a xor b);
    layer7_outputs(2374) <= not b;
    layer7_outputs(2375) <= a;
    layer7_outputs(2376) <= b;
    layer7_outputs(2377) <= not (a or b);
    layer7_outputs(2378) <= not b or a;
    layer7_outputs(2379) <= not a;
    layer7_outputs(2380) <= a and not b;
    layer7_outputs(2381) <= a;
    layer7_outputs(2382) <= not (a and b);
    layer7_outputs(2383) <= not b;
    layer7_outputs(2384) <= not (a or b);
    layer7_outputs(2385) <= not (a and b);
    layer7_outputs(2386) <= not (a and b);
    layer7_outputs(2387) <= not a or b;
    layer7_outputs(2388) <= a and not b;
    layer7_outputs(2389) <= a xor b;
    layer7_outputs(2390) <= not b;
    layer7_outputs(2391) <= a or b;
    layer7_outputs(2392) <= b;
    layer7_outputs(2393) <= a xor b;
    layer7_outputs(2394) <= not (a xor b);
    layer7_outputs(2395) <= not (a xor b);
    layer7_outputs(2396) <= a;
    layer7_outputs(2397) <= b;
    layer7_outputs(2398) <= not (a xor b);
    layer7_outputs(2399) <= a and b;
    layer7_outputs(2400) <= not a;
    layer7_outputs(2401) <= b and not a;
    layer7_outputs(2402) <= a;
    layer7_outputs(2403) <= not (a or b);
    layer7_outputs(2404) <= not a or b;
    layer7_outputs(2405) <= a and not b;
    layer7_outputs(2406) <= not (a xor b);
    layer7_outputs(2407) <= not a or b;
    layer7_outputs(2408) <= b;
    layer7_outputs(2409) <= not b or a;
    layer7_outputs(2410) <= a and not b;
    layer7_outputs(2411) <= b and not a;
    layer7_outputs(2412) <= b and not a;
    layer7_outputs(2413) <= a and not b;
    layer7_outputs(2414) <= not (a or b);
    layer7_outputs(2415) <= not a;
    layer7_outputs(2416) <= not (a or b);
    layer7_outputs(2417) <= not (a or b);
    layer7_outputs(2418) <= not b;
    layer7_outputs(2419) <= a;
    layer7_outputs(2420) <= a or b;
    layer7_outputs(2421) <= a and not b;
    layer7_outputs(2422) <= not (a or b);
    layer7_outputs(2423) <= not b;
    layer7_outputs(2424) <= a xor b;
    layer7_outputs(2425) <= 1'b1;
    layer7_outputs(2426) <= not (a xor b);
    layer7_outputs(2427) <= not (a or b);
    layer7_outputs(2428) <= b;
    layer7_outputs(2429) <= not (a or b);
    layer7_outputs(2430) <= not (a xor b);
    layer7_outputs(2431) <= a;
    layer7_outputs(2432) <= a xor b;
    layer7_outputs(2433) <= b;
    layer7_outputs(2434) <= a xor b;
    layer7_outputs(2435) <= a;
    layer7_outputs(2436) <= b;
    layer7_outputs(2437) <= not b;
    layer7_outputs(2438) <= not a;
    layer7_outputs(2439) <= not a;
    layer7_outputs(2440) <= not a or b;
    layer7_outputs(2441) <= 1'b1;
    layer7_outputs(2442) <= a;
    layer7_outputs(2443) <= not (a or b);
    layer7_outputs(2444) <= not (a and b);
    layer7_outputs(2445) <= not b;
    layer7_outputs(2446) <= not (a and b);
    layer7_outputs(2447) <= not a;
    layer7_outputs(2448) <= not (a xor b);
    layer7_outputs(2449) <= b;
    layer7_outputs(2450) <= not b;
    layer7_outputs(2451) <= a and not b;
    layer7_outputs(2452) <= not b;
    layer7_outputs(2453) <= a;
    layer7_outputs(2454) <= not b;
    layer7_outputs(2455) <= not b;
    layer7_outputs(2456) <= a;
    layer7_outputs(2457) <= 1'b0;
    layer7_outputs(2458) <= a xor b;
    layer7_outputs(2459) <= a and b;
    layer7_outputs(2460) <= not (a and b);
    layer7_outputs(2461) <= a and not b;
    layer7_outputs(2462) <= a xor b;
    layer7_outputs(2463) <= a xor b;
    layer7_outputs(2464) <= not a;
    layer7_outputs(2465) <= a and not b;
    layer7_outputs(2466) <= b;
    layer7_outputs(2467) <= a and not b;
    layer7_outputs(2468) <= not b;
    layer7_outputs(2469) <= not b or a;
    layer7_outputs(2470) <= b;
    layer7_outputs(2471) <= not (a and b);
    layer7_outputs(2472) <= not b or a;
    layer7_outputs(2473) <= not b;
    layer7_outputs(2474) <= a and not b;
    layer7_outputs(2475) <= b;
    layer7_outputs(2476) <= b and not a;
    layer7_outputs(2477) <= not b;
    layer7_outputs(2478) <= not b or a;
    layer7_outputs(2479) <= b and not a;
    layer7_outputs(2480) <= not a or b;
    layer7_outputs(2481) <= not a;
    layer7_outputs(2482) <= a and b;
    layer7_outputs(2483) <= a and b;
    layer7_outputs(2484) <= not (a or b);
    layer7_outputs(2485) <= b;
    layer7_outputs(2486) <= not b or a;
    layer7_outputs(2487) <= not b;
    layer7_outputs(2488) <= not (a or b);
    layer7_outputs(2489) <= b;
    layer7_outputs(2490) <= not (a xor b);
    layer7_outputs(2491) <= not (a or b);
    layer7_outputs(2492) <= a;
    layer7_outputs(2493) <= not a;
    layer7_outputs(2494) <= not b;
    layer7_outputs(2495) <= not (a xor b);
    layer7_outputs(2496) <= not a;
    layer7_outputs(2497) <= not b or a;
    layer7_outputs(2498) <= a xor b;
    layer7_outputs(2499) <= not b;
    layer7_outputs(2500) <= not a;
    layer7_outputs(2501) <= not a;
    layer7_outputs(2502) <= not a;
    layer7_outputs(2503) <= not b;
    layer7_outputs(2504) <= not (a or b);
    layer7_outputs(2505) <= not b or a;
    layer7_outputs(2506) <= not (a and b);
    layer7_outputs(2507) <= not a or b;
    layer7_outputs(2508) <= a xor b;
    layer7_outputs(2509) <= not b or a;
    layer7_outputs(2510) <= b and not a;
    layer7_outputs(2511) <= not a;
    layer7_outputs(2512) <= b;
    layer7_outputs(2513) <= not b;
    layer7_outputs(2514) <= a or b;
    layer7_outputs(2515) <= b;
    layer7_outputs(2516) <= not b or a;
    layer7_outputs(2517) <= b;
    layer7_outputs(2518) <= a or b;
    layer7_outputs(2519) <= not b or a;
    layer7_outputs(2520) <= not (a and b);
    layer7_outputs(2521) <= not a or b;
    layer7_outputs(2522) <= a xor b;
    layer7_outputs(2523) <= not a;
    layer7_outputs(2524) <= b;
    layer7_outputs(2525) <= a and b;
    layer7_outputs(2526) <= a;
    layer7_outputs(2527) <= a;
    layer7_outputs(2528) <= not (a and b);
    layer7_outputs(2529) <= b;
    layer7_outputs(2530) <= a;
    layer7_outputs(2531) <= a;
    layer7_outputs(2532) <= a;
    layer7_outputs(2533) <= a xor b;
    layer7_outputs(2534) <= a;
    layer7_outputs(2535) <= b;
    layer7_outputs(2536) <= not (a or b);
    layer7_outputs(2537) <= a;
    layer7_outputs(2538) <= not a or b;
    layer7_outputs(2539) <= a or b;
    layer7_outputs(2540) <= 1'b0;
    layer7_outputs(2541) <= not b;
    layer7_outputs(2542) <= a and b;
    layer7_outputs(2543) <= not a or b;
    layer7_outputs(2544) <= a;
    layer7_outputs(2545) <= not a;
    layer7_outputs(2546) <= a;
    layer7_outputs(2547) <= not (a xor b);
    layer7_outputs(2548) <= not (a and b);
    layer7_outputs(2549) <= not b;
    layer7_outputs(2550) <= a or b;
    layer7_outputs(2551) <= a xor b;
    layer7_outputs(2552) <= b;
    layer7_outputs(2553) <= not a;
    layer7_outputs(2554) <= not (a or b);
    layer7_outputs(2555) <= b and not a;
    layer7_outputs(2556) <= not b;
    layer7_outputs(2557) <= 1'b1;
    layer7_outputs(2558) <= b;
    layer7_outputs(2559) <= a;
    layer8_outputs(0) <= not b;
    layer8_outputs(1) <= not (a xor b);
    layer8_outputs(2) <= a;
    layer8_outputs(3) <= a or b;
    layer8_outputs(4) <= a;
    layer8_outputs(5) <= a and not b;
    layer8_outputs(6) <= a;
    layer8_outputs(7) <= a xor b;
    layer8_outputs(8) <= not b;
    layer8_outputs(9) <= a and b;
    layer8_outputs(10) <= not (a or b);
    layer8_outputs(11) <= not a;
    layer8_outputs(12) <= b;
    layer8_outputs(13) <= not (a and b);
    layer8_outputs(14) <= not (a xor b);
    layer8_outputs(15) <= 1'b0;
    layer8_outputs(16) <= a;
    layer8_outputs(17) <= not a;
    layer8_outputs(18) <= not (a or b);
    layer8_outputs(19) <= not (a xor b);
    layer8_outputs(20) <= a;
    layer8_outputs(21) <= a or b;
    layer8_outputs(22) <= not (a and b);
    layer8_outputs(23) <= a;
    layer8_outputs(24) <= not b;
    layer8_outputs(25) <= a;
    layer8_outputs(26) <= a or b;
    layer8_outputs(27) <= not b or a;
    layer8_outputs(28) <= a;
    layer8_outputs(29) <= not a;
    layer8_outputs(30) <= a;
    layer8_outputs(31) <= b and not a;
    layer8_outputs(32) <= a and b;
    layer8_outputs(33) <= not b;
    layer8_outputs(34) <= a or b;
    layer8_outputs(35) <= b;
    layer8_outputs(36) <= not b or a;
    layer8_outputs(37) <= b and not a;
    layer8_outputs(38) <= not a or b;
    layer8_outputs(39) <= b;
    layer8_outputs(40) <= not (a xor b);
    layer8_outputs(41) <= a or b;
    layer8_outputs(42) <= not b or a;
    layer8_outputs(43) <= not a;
    layer8_outputs(44) <= b;
    layer8_outputs(45) <= not (a or b);
    layer8_outputs(46) <= a xor b;
    layer8_outputs(47) <= not b or a;
    layer8_outputs(48) <= not (a or b);
    layer8_outputs(49) <= not b;
    layer8_outputs(50) <= b;
    layer8_outputs(51) <= a and b;
    layer8_outputs(52) <= not (a xor b);
    layer8_outputs(53) <= b;
    layer8_outputs(54) <= a xor b;
    layer8_outputs(55) <= b;
    layer8_outputs(56) <= a;
    layer8_outputs(57) <= b and not a;
    layer8_outputs(58) <= not b;
    layer8_outputs(59) <= not b;
    layer8_outputs(60) <= b;
    layer8_outputs(61) <= a xor b;
    layer8_outputs(62) <= a and b;
    layer8_outputs(63) <= a and b;
    layer8_outputs(64) <= not b;
    layer8_outputs(65) <= b and not a;
    layer8_outputs(66) <= b;
    layer8_outputs(67) <= b;
    layer8_outputs(68) <= a xor b;
    layer8_outputs(69) <= not b or a;
    layer8_outputs(70) <= a xor b;
    layer8_outputs(71) <= not b or a;
    layer8_outputs(72) <= not a;
    layer8_outputs(73) <= a;
    layer8_outputs(74) <= b;
    layer8_outputs(75) <= not (a and b);
    layer8_outputs(76) <= a and not b;
    layer8_outputs(77) <= b and not a;
    layer8_outputs(78) <= not (a and b);
    layer8_outputs(79) <= not (a xor b);
    layer8_outputs(80) <= not a or b;
    layer8_outputs(81) <= not b or a;
    layer8_outputs(82) <= a xor b;
    layer8_outputs(83) <= not a or b;
    layer8_outputs(84) <= not a;
    layer8_outputs(85) <= not a or b;
    layer8_outputs(86) <= a or b;
    layer8_outputs(87) <= not (a xor b);
    layer8_outputs(88) <= not a or b;
    layer8_outputs(89) <= a xor b;
    layer8_outputs(90) <= not a or b;
    layer8_outputs(91) <= a xor b;
    layer8_outputs(92) <= b;
    layer8_outputs(93) <= not a;
    layer8_outputs(94) <= a and not b;
    layer8_outputs(95) <= a xor b;
    layer8_outputs(96) <= a or b;
    layer8_outputs(97) <= a;
    layer8_outputs(98) <= b;
    layer8_outputs(99) <= not a or b;
    layer8_outputs(100) <= a;
    layer8_outputs(101) <= not (a and b);
    layer8_outputs(102) <= not (a xor b);
    layer8_outputs(103) <= not a;
    layer8_outputs(104) <= a xor b;
    layer8_outputs(105) <= not b;
    layer8_outputs(106) <= not b;
    layer8_outputs(107) <= a xor b;
    layer8_outputs(108) <= b;
    layer8_outputs(109) <= not b;
    layer8_outputs(110) <= a and b;
    layer8_outputs(111) <= not (a xor b);
    layer8_outputs(112) <= not a;
    layer8_outputs(113) <= b;
    layer8_outputs(114) <= b and not a;
    layer8_outputs(115) <= b and not a;
    layer8_outputs(116) <= a xor b;
    layer8_outputs(117) <= not (a xor b);
    layer8_outputs(118) <= not a;
    layer8_outputs(119) <= not a;
    layer8_outputs(120) <= not a or b;
    layer8_outputs(121) <= not b;
    layer8_outputs(122) <= not a or b;
    layer8_outputs(123) <= b and not a;
    layer8_outputs(124) <= b;
    layer8_outputs(125) <= not b;
    layer8_outputs(126) <= not a;
    layer8_outputs(127) <= not (a xor b);
    layer8_outputs(128) <= a;
    layer8_outputs(129) <= b and not a;
    layer8_outputs(130) <= a and not b;
    layer8_outputs(131) <= 1'b1;
    layer8_outputs(132) <= b;
    layer8_outputs(133) <= not b;
    layer8_outputs(134) <= b;
    layer8_outputs(135) <= not (a xor b);
    layer8_outputs(136) <= a xor b;
    layer8_outputs(137) <= b;
    layer8_outputs(138) <= not a or b;
    layer8_outputs(139) <= a;
    layer8_outputs(140) <= a and not b;
    layer8_outputs(141) <= not b or a;
    layer8_outputs(142) <= not b;
    layer8_outputs(143) <= not b;
    layer8_outputs(144) <= b;
    layer8_outputs(145) <= a;
    layer8_outputs(146) <= b and not a;
    layer8_outputs(147) <= a and not b;
    layer8_outputs(148) <= a xor b;
    layer8_outputs(149) <= not b;
    layer8_outputs(150) <= not a or b;
    layer8_outputs(151) <= not b;
    layer8_outputs(152) <= a and b;
    layer8_outputs(153) <= not (a and b);
    layer8_outputs(154) <= a;
    layer8_outputs(155) <= a xor b;
    layer8_outputs(156) <= not (a xor b);
    layer8_outputs(157) <= not a;
    layer8_outputs(158) <= b;
    layer8_outputs(159) <= not a or b;
    layer8_outputs(160) <= a and not b;
    layer8_outputs(161) <= not b or a;
    layer8_outputs(162) <= b;
    layer8_outputs(163) <= not b or a;
    layer8_outputs(164) <= not (a xor b);
    layer8_outputs(165) <= not (a or b);
    layer8_outputs(166) <= not a;
    layer8_outputs(167) <= not (a and b);
    layer8_outputs(168) <= a and not b;
    layer8_outputs(169) <= not (a xor b);
    layer8_outputs(170) <= not (a xor b);
    layer8_outputs(171) <= not (a and b);
    layer8_outputs(172) <= not b;
    layer8_outputs(173) <= not (a or b);
    layer8_outputs(174) <= not a or b;
    layer8_outputs(175) <= not b;
    layer8_outputs(176) <= not (a xor b);
    layer8_outputs(177) <= a;
    layer8_outputs(178) <= 1'b0;
    layer8_outputs(179) <= not b;
    layer8_outputs(180) <= b and not a;
    layer8_outputs(181) <= a and not b;
    layer8_outputs(182) <= not (a xor b);
    layer8_outputs(183) <= a xor b;
    layer8_outputs(184) <= b;
    layer8_outputs(185) <= b;
    layer8_outputs(186) <= not (a xor b);
    layer8_outputs(187) <= b;
    layer8_outputs(188) <= not b or a;
    layer8_outputs(189) <= not a;
    layer8_outputs(190) <= not a;
    layer8_outputs(191) <= not b or a;
    layer8_outputs(192) <= not b;
    layer8_outputs(193) <= a or b;
    layer8_outputs(194) <= a and b;
    layer8_outputs(195) <= a xor b;
    layer8_outputs(196) <= not a;
    layer8_outputs(197) <= b;
    layer8_outputs(198) <= a and not b;
    layer8_outputs(199) <= not (a or b);
    layer8_outputs(200) <= 1'b1;
    layer8_outputs(201) <= a or b;
    layer8_outputs(202) <= a or b;
    layer8_outputs(203) <= not (a and b);
    layer8_outputs(204) <= 1'b1;
    layer8_outputs(205) <= b and not a;
    layer8_outputs(206) <= not (a and b);
    layer8_outputs(207) <= b and not a;
    layer8_outputs(208) <= a xor b;
    layer8_outputs(209) <= not (a or b);
    layer8_outputs(210) <= b;
    layer8_outputs(211) <= not b;
    layer8_outputs(212) <= 1'b0;
    layer8_outputs(213) <= b;
    layer8_outputs(214) <= not (a or b);
    layer8_outputs(215) <= a and b;
    layer8_outputs(216) <= not a or b;
    layer8_outputs(217) <= a and b;
    layer8_outputs(218) <= a and not b;
    layer8_outputs(219) <= not b;
    layer8_outputs(220) <= not a;
    layer8_outputs(221) <= not a or b;
    layer8_outputs(222) <= not a;
    layer8_outputs(223) <= not b;
    layer8_outputs(224) <= a and not b;
    layer8_outputs(225) <= a;
    layer8_outputs(226) <= a and not b;
    layer8_outputs(227) <= a and not b;
    layer8_outputs(228) <= not (a and b);
    layer8_outputs(229) <= a;
    layer8_outputs(230) <= not (a and b);
    layer8_outputs(231) <= a and not b;
    layer8_outputs(232) <= a or b;
    layer8_outputs(233) <= not a;
    layer8_outputs(234) <= a or b;
    layer8_outputs(235) <= a;
    layer8_outputs(236) <= a xor b;
    layer8_outputs(237) <= b;
    layer8_outputs(238) <= not (a xor b);
    layer8_outputs(239) <= b;
    layer8_outputs(240) <= b and not a;
    layer8_outputs(241) <= a;
    layer8_outputs(242) <= not b or a;
    layer8_outputs(243) <= not b;
    layer8_outputs(244) <= not a;
    layer8_outputs(245) <= b;
    layer8_outputs(246) <= b;
    layer8_outputs(247) <= b;
    layer8_outputs(248) <= not b;
    layer8_outputs(249) <= a and b;
    layer8_outputs(250) <= a xor b;
    layer8_outputs(251) <= not b or a;
    layer8_outputs(252) <= a xor b;
    layer8_outputs(253) <= b;
    layer8_outputs(254) <= not a;
    layer8_outputs(255) <= not (a xor b);
    layer8_outputs(256) <= not a;
    layer8_outputs(257) <= a or b;
    layer8_outputs(258) <= not a or b;
    layer8_outputs(259) <= not (a and b);
    layer8_outputs(260) <= b and not a;
    layer8_outputs(261) <= b;
    layer8_outputs(262) <= not b;
    layer8_outputs(263) <= not b;
    layer8_outputs(264) <= a xor b;
    layer8_outputs(265) <= not (a and b);
    layer8_outputs(266) <= 1'b1;
    layer8_outputs(267) <= not (a xor b);
    layer8_outputs(268) <= not b;
    layer8_outputs(269) <= a and not b;
    layer8_outputs(270) <= not b;
    layer8_outputs(271) <= not b;
    layer8_outputs(272) <= not b or a;
    layer8_outputs(273) <= b;
    layer8_outputs(274) <= not (a or b);
    layer8_outputs(275) <= not (a xor b);
    layer8_outputs(276) <= b and not a;
    layer8_outputs(277) <= a;
    layer8_outputs(278) <= not b or a;
    layer8_outputs(279) <= not a;
    layer8_outputs(280) <= b;
    layer8_outputs(281) <= not (a and b);
    layer8_outputs(282) <= b;
    layer8_outputs(283) <= not b;
    layer8_outputs(284) <= a and b;
    layer8_outputs(285) <= a;
    layer8_outputs(286) <= a xor b;
    layer8_outputs(287) <= b;
    layer8_outputs(288) <= not (a and b);
    layer8_outputs(289) <= a;
    layer8_outputs(290) <= not (a xor b);
    layer8_outputs(291) <= not (a and b);
    layer8_outputs(292) <= not b or a;
    layer8_outputs(293) <= b and not a;
    layer8_outputs(294) <= a;
    layer8_outputs(295) <= not a;
    layer8_outputs(296) <= b and not a;
    layer8_outputs(297) <= a or b;
    layer8_outputs(298) <= 1'b0;
    layer8_outputs(299) <= not b;
    layer8_outputs(300) <= not (a xor b);
    layer8_outputs(301) <= not (a and b);
    layer8_outputs(302) <= a or b;
    layer8_outputs(303) <= b and not a;
    layer8_outputs(304) <= a and not b;
    layer8_outputs(305) <= not (a xor b);
    layer8_outputs(306) <= b;
    layer8_outputs(307) <= 1'b1;
    layer8_outputs(308) <= a;
    layer8_outputs(309) <= not a or b;
    layer8_outputs(310) <= not (a and b);
    layer8_outputs(311) <= not a;
    layer8_outputs(312) <= not (a xor b);
    layer8_outputs(313) <= a;
    layer8_outputs(314) <= not a or b;
    layer8_outputs(315) <= b;
    layer8_outputs(316) <= not b;
    layer8_outputs(317) <= 1'b0;
    layer8_outputs(318) <= b;
    layer8_outputs(319) <= not b or a;
    layer8_outputs(320) <= not (a xor b);
    layer8_outputs(321) <= a or b;
    layer8_outputs(322) <= b;
    layer8_outputs(323) <= not (a and b);
    layer8_outputs(324) <= a;
    layer8_outputs(325) <= a or b;
    layer8_outputs(326) <= a xor b;
    layer8_outputs(327) <= b;
    layer8_outputs(328) <= not (a and b);
    layer8_outputs(329) <= not a or b;
    layer8_outputs(330) <= not a;
    layer8_outputs(331) <= 1'b0;
    layer8_outputs(332) <= a xor b;
    layer8_outputs(333) <= a and b;
    layer8_outputs(334) <= b and not a;
    layer8_outputs(335) <= a;
    layer8_outputs(336) <= a xor b;
    layer8_outputs(337) <= a;
    layer8_outputs(338) <= not a;
    layer8_outputs(339) <= not b;
    layer8_outputs(340) <= a or b;
    layer8_outputs(341) <= b and not a;
    layer8_outputs(342) <= not b or a;
    layer8_outputs(343) <= not (a or b);
    layer8_outputs(344) <= a;
    layer8_outputs(345) <= a;
    layer8_outputs(346) <= not (a and b);
    layer8_outputs(347) <= b;
    layer8_outputs(348) <= a or b;
    layer8_outputs(349) <= a;
    layer8_outputs(350) <= b;
    layer8_outputs(351) <= not (a xor b);
    layer8_outputs(352) <= a and not b;
    layer8_outputs(353) <= not a or b;
    layer8_outputs(354) <= a and not b;
    layer8_outputs(355) <= a;
    layer8_outputs(356) <= a or b;
    layer8_outputs(357) <= not (a or b);
    layer8_outputs(358) <= not b;
    layer8_outputs(359) <= not a;
    layer8_outputs(360) <= not b;
    layer8_outputs(361) <= not a;
    layer8_outputs(362) <= not (a xor b);
    layer8_outputs(363) <= a or b;
    layer8_outputs(364) <= b and not a;
    layer8_outputs(365) <= a xor b;
    layer8_outputs(366) <= a and b;
    layer8_outputs(367) <= a;
    layer8_outputs(368) <= not a;
    layer8_outputs(369) <= not (a or b);
    layer8_outputs(370) <= not (a and b);
    layer8_outputs(371) <= not b;
    layer8_outputs(372) <= a;
    layer8_outputs(373) <= a and not b;
    layer8_outputs(374) <= a;
    layer8_outputs(375) <= a and b;
    layer8_outputs(376) <= a or b;
    layer8_outputs(377) <= not (a xor b);
    layer8_outputs(378) <= not (a xor b);
    layer8_outputs(379) <= a xor b;
    layer8_outputs(380) <= not a;
    layer8_outputs(381) <= not b;
    layer8_outputs(382) <= not a or b;
    layer8_outputs(383) <= not a;
    layer8_outputs(384) <= a or b;
    layer8_outputs(385) <= a and b;
    layer8_outputs(386) <= a and not b;
    layer8_outputs(387) <= a;
    layer8_outputs(388) <= not a;
    layer8_outputs(389) <= not (a or b);
    layer8_outputs(390) <= b;
    layer8_outputs(391) <= a;
    layer8_outputs(392) <= a and not b;
    layer8_outputs(393) <= a and not b;
    layer8_outputs(394) <= not (a xor b);
    layer8_outputs(395) <= a xor b;
    layer8_outputs(396) <= b;
    layer8_outputs(397) <= b;
    layer8_outputs(398) <= b and not a;
    layer8_outputs(399) <= a and not b;
    layer8_outputs(400) <= not a;
    layer8_outputs(401) <= a and b;
    layer8_outputs(402) <= not b;
    layer8_outputs(403) <= not (a or b);
    layer8_outputs(404) <= a;
    layer8_outputs(405) <= not (a and b);
    layer8_outputs(406) <= a;
    layer8_outputs(407) <= not (a and b);
    layer8_outputs(408) <= not b;
    layer8_outputs(409) <= not a;
    layer8_outputs(410) <= not (a xor b);
    layer8_outputs(411) <= not (a xor b);
    layer8_outputs(412) <= a or b;
    layer8_outputs(413) <= a;
    layer8_outputs(414) <= not a or b;
    layer8_outputs(415) <= a or b;
    layer8_outputs(416) <= not (a and b);
    layer8_outputs(417) <= a and b;
    layer8_outputs(418) <= not (a xor b);
    layer8_outputs(419) <= not b;
    layer8_outputs(420) <= a or b;
    layer8_outputs(421) <= not b;
    layer8_outputs(422) <= not b;
    layer8_outputs(423) <= not (a or b);
    layer8_outputs(424) <= b;
    layer8_outputs(425) <= not b;
    layer8_outputs(426) <= not a or b;
    layer8_outputs(427) <= not (a xor b);
    layer8_outputs(428) <= not (a and b);
    layer8_outputs(429) <= a xor b;
    layer8_outputs(430) <= a xor b;
    layer8_outputs(431) <= not b or a;
    layer8_outputs(432) <= not (a or b);
    layer8_outputs(433) <= not a or b;
    layer8_outputs(434) <= a or b;
    layer8_outputs(435) <= a xor b;
    layer8_outputs(436) <= not b;
    layer8_outputs(437) <= not (a and b);
    layer8_outputs(438) <= not (a xor b);
    layer8_outputs(439) <= a and b;
    layer8_outputs(440) <= b;
    layer8_outputs(441) <= not (a xor b);
    layer8_outputs(442) <= a and b;
    layer8_outputs(443) <= a xor b;
    layer8_outputs(444) <= a;
    layer8_outputs(445) <= a;
    layer8_outputs(446) <= b;
    layer8_outputs(447) <= not a;
    layer8_outputs(448) <= b and not a;
    layer8_outputs(449) <= not (a or b);
    layer8_outputs(450) <= not (a and b);
    layer8_outputs(451) <= a and not b;
    layer8_outputs(452) <= b;
    layer8_outputs(453) <= 1'b0;
    layer8_outputs(454) <= a xor b;
    layer8_outputs(455) <= 1'b0;
    layer8_outputs(456) <= a or b;
    layer8_outputs(457) <= not b;
    layer8_outputs(458) <= not (a xor b);
    layer8_outputs(459) <= a;
    layer8_outputs(460) <= a xor b;
    layer8_outputs(461) <= not (a xor b);
    layer8_outputs(462) <= not b;
    layer8_outputs(463) <= not b;
    layer8_outputs(464) <= a and b;
    layer8_outputs(465) <= b;
    layer8_outputs(466) <= a xor b;
    layer8_outputs(467) <= a or b;
    layer8_outputs(468) <= not b;
    layer8_outputs(469) <= not (a and b);
    layer8_outputs(470) <= not b;
    layer8_outputs(471) <= not a;
    layer8_outputs(472) <= a;
    layer8_outputs(473) <= a or b;
    layer8_outputs(474) <= not b or a;
    layer8_outputs(475) <= not b;
    layer8_outputs(476) <= not a or b;
    layer8_outputs(477) <= a;
    layer8_outputs(478) <= a and not b;
    layer8_outputs(479) <= not (a xor b);
    layer8_outputs(480) <= a;
    layer8_outputs(481) <= b;
    layer8_outputs(482) <= a or b;
    layer8_outputs(483) <= not b;
    layer8_outputs(484) <= a xor b;
    layer8_outputs(485) <= a xor b;
    layer8_outputs(486) <= a or b;
    layer8_outputs(487) <= a and b;
    layer8_outputs(488) <= not b;
    layer8_outputs(489) <= not b or a;
    layer8_outputs(490) <= not (a or b);
    layer8_outputs(491) <= not (a xor b);
    layer8_outputs(492) <= b;
    layer8_outputs(493) <= not (a xor b);
    layer8_outputs(494) <= not (a and b);
    layer8_outputs(495) <= a;
    layer8_outputs(496) <= b;
    layer8_outputs(497) <= not (a xor b);
    layer8_outputs(498) <= not (a or b);
    layer8_outputs(499) <= a;
    layer8_outputs(500) <= b;
    layer8_outputs(501) <= a and b;
    layer8_outputs(502) <= a or b;
    layer8_outputs(503) <= not a;
    layer8_outputs(504) <= not b;
    layer8_outputs(505) <= a xor b;
    layer8_outputs(506) <= not b;
    layer8_outputs(507) <= b;
    layer8_outputs(508) <= not b;
    layer8_outputs(509) <= not a or b;
    layer8_outputs(510) <= b;
    layer8_outputs(511) <= 1'b1;
    layer8_outputs(512) <= not (a and b);
    layer8_outputs(513) <= a and not b;
    layer8_outputs(514) <= not (a or b);
    layer8_outputs(515) <= b;
    layer8_outputs(516) <= not b;
    layer8_outputs(517) <= a;
    layer8_outputs(518) <= b and not a;
    layer8_outputs(519) <= not b;
    layer8_outputs(520) <= a and not b;
    layer8_outputs(521) <= not a;
    layer8_outputs(522) <= not (a xor b);
    layer8_outputs(523) <= not b or a;
    layer8_outputs(524) <= not a;
    layer8_outputs(525) <= b and not a;
    layer8_outputs(526) <= a and b;
    layer8_outputs(527) <= not b;
    layer8_outputs(528) <= a and not b;
    layer8_outputs(529) <= not a;
    layer8_outputs(530) <= not (a xor b);
    layer8_outputs(531) <= not b;
    layer8_outputs(532) <= not a;
    layer8_outputs(533) <= not a;
    layer8_outputs(534) <= not (a xor b);
    layer8_outputs(535) <= not a or b;
    layer8_outputs(536) <= not (a or b);
    layer8_outputs(537) <= not a or b;
    layer8_outputs(538) <= a and not b;
    layer8_outputs(539) <= b;
    layer8_outputs(540) <= a;
    layer8_outputs(541) <= b;
    layer8_outputs(542) <= a xor b;
    layer8_outputs(543) <= a xor b;
    layer8_outputs(544) <= not b;
    layer8_outputs(545) <= a;
    layer8_outputs(546) <= not b;
    layer8_outputs(547) <= not (a or b);
    layer8_outputs(548) <= not b;
    layer8_outputs(549) <= a and not b;
    layer8_outputs(550) <= not a or b;
    layer8_outputs(551) <= not (a xor b);
    layer8_outputs(552) <= a and not b;
    layer8_outputs(553) <= a xor b;
    layer8_outputs(554) <= not a or b;
    layer8_outputs(555) <= not b;
    layer8_outputs(556) <= not a;
    layer8_outputs(557) <= not a or b;
    layer8_outputs(558) <= b;
    layer8_outputs(559) <= not b or a;
    layer8_outputs(560) <= not a or b;
    layer8_outputs(561) <= a and not b;
    layer8_outputs(562) <= a;
    layer8_outputs(563) <= a xor b;
    layer8_outputs(564) <= not (a or b);
    layer8_outputs(565) <= a;
    layer8_outputs(566) <= b;
    layer8_outputs(567) <= a or b;
    layer8_outputs(568) <= not b;
    layer8_outputs(569) <= not a;
    layer8_outputs(570) <= not b;
    layer8_outputs(571) <= a xor b;
    layer8_outputs(572) <= b;
    layer8_outputs(573) <= not (a and b);
    layer8_outputs(574) <= not a;
    layer8_outputs(575) <= not a or b;
    layer8_outputs(576) <= a and b;
    layer8_outputs(577) <= b and not a;
    layer8_outputs(578) <= a xor b;
    layer8_outputs(579) <= a;
    layer8_outputs(580) <= not a;
    layer8_outputs(581) <= a and not b;
    layer8_outputs(582) <= not b;
    layer8_outputs(583) <= a xor b;
    layer8_outputs(584) <= b and not a;
    layer8_outputs(585) <= a and not b;
    layer8_outputs(586) <= not a;
    layer8_outputs(587) <= b;
    layer8_outputs(588) <= a;
    layer8_outputs(589) <= not a;
    layer8_outputs(590) <= a;
    layer8_outputs(591) <= not a;
    layer8_outputs(592) <= b;
    layer8_outputs(593) <= a and not b;
    layer8_outputs(594) <= not a;
    layer8_outputs(595) <= a xor b;
    layer8_outputs(596) <= not b;
    layer8_outputs(597) <= not (a xor b);
    layer8_outputs(598) <= not b or a;
    layer8_outputs(599) <= not (a xor b);
    layer8_outputs(600) <= not a;
    layer8_outputs(601) <= a and b;
    layer8_outputs(602) <= not a;
    layer8_outputs(603) <= not (a or b);
    layer8_outputs(604) <= not b;
    layer8_outputs(605) <= a;
    layer8_outputs(606) <= not a or b;
    layer8_outputs(607) <= not b;
    layer8_outputs(608) <= a and not b;
    layer8_outputs(609) <= b;
    layer8_outputs(610) <= not (a xor b);
    layer8_outputs(611) <= not b or a;
    layer8_outputs(612) <= a xor b;
    layer8_outputs(613) <= a or b;
    layer8_outputs(614) <= b;
    layer8_outputs(615) <= a;
    layer8_outputs(616) <= a or b;
    layer8_outputs(617) <= not b;
    layer8_outputs(618) <= not a;
    layer8_outputs(619) <= not (a and b);
    layer8_outputs(620) <= 1'b0;
    layer8_outputs(621) <= b and not a;
    layer8_outputs(622) <= not a;
    layer8_outputs(623) <= a;
    layer8_outputs(624) <= not b or a;
    layer8_outputs(625) <= b;
    layer8_outputs(626) <= not a;
    layer8_outputs(627) <= not (a or b);
    layer8_outputs(628) <= a or b;
    layer8_outputs(629) <= b and not a;
    layer8_outputs(630) <= not (a or b);
    layer8_outputs(631) <= a xor b;
    layer8_outputs(632) <= a;
    layer8_outputs(633) <= a;
    layer8_outputs(634) <= not (a xor b);
    layer8_outputs(635) <= b;
    layer8_outputs(636) <= b;
    layer8_outputs(637) <= not (a and b);
    layer8_outputs(638) <= b;
    layer8_outputs(639) <= not a;
    layer8_outputs(640) <= not (a xor b);
    layer8_outputs(641) <= a or b;
    layer8_outputs(642) <= not b;
    layer8_outputs(643) <= not b;
    layer8_outputs(644) <= a;
    layer8_outputs(645) <= a or b;
    layer8_outputs(646) <= a or b;
    layer8_outputs(647) <= not a or b;
    layer8_outputs(648) <= not a or b;
    layer8_outputs(649) <= b;
    layer8_outputs(650) <= not (a and b);
    layer8_outputs(651) <= b;
    layer8_outputs(652) <= a;
    layer8_outputs(653) <= not a;
    layer8_outputs(654) <= a and not b;
    layer8_outputs(655) <= not (a xor b);
    layer8_outputs(656) <= not a;
    layer8_outputs(657) <= a or b;
    layer8_outputs(658) <= not b;
    layer8_outputs(659) <= not b;
    layer8_outputs(660) <= b;
    layer8_outputs(661) <= b;
    layer8_outputs(662) <= not b or a;
    layer8_outputs(663) <= not b;
    layer8_outputs(664) <= not a;
    layer8_outputs(665) <= not a;
    layer8_outputs(666) <= not a or b;
    layer8_outputs(667) <= not b;
    layer8_outputs(668) <= a xor b;
    layer8_outputs(669) <= not a;
    layer8_outputs(670) <= a and b;
    layer8_outputs(671) <= not (a xor b);
    layer8_outputs(672) <= not b or a;
    layer8_outputs(673) <= not (a or b);
    layer8_outputs(674) <= not a;
    layer8_outputs(675) <= b and not a;
    layer8_outputs(676) <= a and b;
    layer8_outputs(677) <= b and not a;
    layer8_outputs(678) <= not a or b;
    layer8_outputs(679) <= a xor b;
    layer8_outputs(680) <= not b or a;
    layer8_outputs(681) <= not b;
    layer8_outputs(682) <= not a;
    layer8_outputs(683) <= a;
    layer8_outputs(684) <= b;
    layer8_outputs(685) <= not b;
    layer8_outputs(686) <= not a;
    layer8_outputs(687) <= a or b;
    layer8_outputs(688) <= not a;
    layer8_outputs(689) <= a and b;
    layer8_outputs(690) <= a and b;
    layer8_outputs(691) <= not b or a;
    layer8_outputs(692) <= a;
    layer8_outputs(693) <= not b;
    layer8_outputs(694) <= a xor b;
    layer8_outputs(695) <= not a;
    layer8_outputs(696) <= not b or a;
    layer8_outputs(697) <= a;
    layer8_outputs(698) <= a xor b;
    layer8_outputs(699) <= not b;
    layer8_outputs(700) <= not a;
    layer8_outputs(701) <= not b;
    layer8_outputs(702) <= a;
    layer8_outputs(703) <= a or b;
    layer8_outputs(704) <= not b or a;
    layer8_outputs(705) <= not (a or b);
    layer8_outputs(706) <= b;
    layer8_outputs(707) <= a or b;
    layer8_outputs(708) <= not b or a;
    layer8_outputs(709) <= b;
    layer8_outputs(710) <= a and b;
    layer8_outputs(711) <= not a;
    layer8_outputs(712) <= a xor b;
    layer8_outputs(713) <= a and not b;
    layer8_outputs(714) <= a or b;
    layer8_outputs(715) <= not a;
    layer8_outputs(716) <= not (a or b);
    layer8_outputs(717) <= a and b;
    layer8_outputs(718) <= not (a and b);
    layer8_outputs(719) <= not b;
    layer8_outputs(720) <= not (a xor b);
    layer8_outputs(721) <= a or b;
    layer8_outputs(722) <= not a;
    layer8_outputs(723) <= not a;
    layer8_outputs(724) <= not a;
    layer8_outputs(725) <= a;
    layer8_outputs(726) <= a and b;
    layer8_outputs(727) <= not (a xor b);
    layer8_outputs(728) <= a or b;
    layer8_outputs(729) <= a and not b;
    layer8_outputs(730) <= a or b;
    layer8_outputs(731) <= not a or b;
    layer8_outputs(732) <= not a;
    layer8_outputs(733) <= not b or a;
    layer8_outputs(734) <= not (a and b);
    layer8_outputs(735) <= a and not b;
    layer8_outputs(736) <= a and not b;
    layer8_outputs(737) <= not b;
    layer8_outputs(738) <= a xor b;
    layer8_outputs(739) <= a and b;
    layer8_outputs(740) <= a or b;
    layer8_outputs(741) <= not (a and b);
    layer8_outputs(742) <= b;
    layer8_outputs(743) <= not a or b;
    layer8_outputs(744) <= not (a or b);
    layer8_outputs(745) <= not (a and b);
    layer8_outputs(746) <= not a or b;
    layer8_outputs(747) <= b;
    layer8_outputs(748) <= not b;
    layer8_outputs(749) <= a and b;
    layer8_outputs(750) <= b;
    layer8_outputs(751) <= not (a xor b);
    layer8_outputs(752) <= not (a or b);
    layer8_outputs(753) <= not b;
    layer8_outputs(754) <= a;
    layer8_outputs(755) <= b and not a;
    layer8_outputs(756) <= a;
    layer8_outputs(757) <= a and not b;
    layer8_outputs(758) <= a and not b;
    layer8_outputs(759) <= not (a and b);
    layer8_outputs(760) <= b;
    layer8_outputs(761) <= not a;
    layer8_outputs(762) <= not a;
    layer8_outputs(763) <= b;
    layer8_outputs(764) <= not (a xor b);
    layer8_outputs(765) <= not b;
    layer8_outputs(766) <= not a or b;
    layer8_outputs(767) <= not b;
    layer8_outputs(768) <= a or b;
    layer8_outputs(769) <= not (a xor b);
    layer8_outputs(770) <= a xor b;
    layer8_outputs(771) <= a and b;
    layer8_outputs(772) <= not a or b;
    layer8_outputs(773) <= b;
    layer8_outputs(774) <= a;
    layer8_outputs(775) <= not a;
    layer8_outputs(776) <= b and not a;
    layer8_outputs(777) <= not b;
    layer8_outputs(778) <= not b or a;
    layer8_outputs(779) <= not (a xor b);
    layer8_outputs(780) <= b;
    layer8_outputs(781) <= not b;
    layer8_outputs(782) <= not a;
    layer8_outputs(783) <= not b;
    layer8_outputs(784) <= not (a and b);
    layer8_outputs(785) <= a xor b;
    layer8_outputs(786) <= not (a xor b);
    layer8_outputs(787) <= a or b;
    layer8_outputs(788) <= not b;
    layer8_outputs(789) <= b;
    layer8_outputs(790) <= b and not a;
    layer8_outputs(791) <= not b;
    layer8_outputs(792) <= not (a xor b);
    layer8_outputs(793) <= not a or b;
    layer8_outputs(794) <= not a or b;
    layer8_outputs(795) <= b;
    layer8_outputs(796) <= a;
    layer8_outputs(797) <= a xor b;
    layer8_outputs(798) <= not a;
    layer8_outputs(799) <= not a;
    layer8_outputs(800) <= b;
    layer8_outputs(801) <= not a or b;
    layer8_outputs(802) <= b;
    layer8_outputs(803) <= not a;
    layer8_outputs(804) <= not a;
    layer8_outputs(805) <= b;
    layer8_outputs(806) <= a;
    layer8_outputs(807) <= not b;
    layer8_outputs(808) <= not b;
    layer8_outputs(809) <= b and not a;
    layer8_outputs(810) <= a;
    layer8_outputs(811) <= a or b;
    layer8_outputs(812) <= not (a xor b);
    layer8_outputs(813) <= a xor b;
    layer8_outputs(814) <= not b;
    layer8_outputs(815) <= not a or b;
    layer8_outputs(816) <= not (a or b);
    layer8_outputs(817) <= a and not b;
    layer8_outputs(818) <= a and b;
    layer8_outputs(819) <= b;
    layer8_outputs(820) <= not b;
    layer8_outputs(821) <= not b;
    layer8_outputs(822) <= a or b;
    layer8_outputs(823) <= 1'b1;
    layer8_outputs(824) <= a and not b;
    layer8_outputs(825) <= b;
    layer8_outputs(826) <= not (a and b);
    layer8_outputs(827) <= a;
    layer8_outputs(828) <= a or b;
    layer8_outputs(829) <= not (a xor b);
    layer8_outputs(830) <= not b;
    layer8_outputs(831) <= not b;
    layer8_outputs(832) <= not (a xor b);
    layer8_outputs(833) <= not a;
    layer8_outputs(834) <= not b or a;
    layer8_outputs(835) <= not a;
    layer8_outputs(836) <= b;
    layer8_outputs(837) <= not b;
    layer8_outputs(838) <= not a;
    layer8_outputs(839) <= a;
    layer8_outputs(840) <= not b or a;
    layer8_outputs(841) <= a and not b;
    layer8_outputs(842) <= not a or b;
    layer8_outputs(843) <= a and not b;
    layer8_outputs(844) <= b;
    layer8_outputs(845) <= b;
    layer8_outputs(846) <= not (a and b);
    layer8_outputs(847) <= not b;
    layer8_outputs(848) <= not (a or b);
    layer8_outputs(849) <= b;
    layer8_outputs(850) <= not b;
    layer8_outputs(851) <= a xor b;
    layer8_outputs(852) <= not b;
    layer8_outputs(853) <= b and not a;
    layer8_outputs(854) <= b;
    layer8_outputs(855) <= not b;
    layer8_outputs(856) <= not (a and b);
    layer8_outputs(857) <= not b or a;
    layer8_outputs(858) <= a and not b;
    layer8_outputs(859) <= not a;
    layer8_outputs(860) <= not b or a;
    layer8_outputs(861) <= not (a and b);
    layer8_outputs(862) <= a and not b;
    layer8_outputs(863) <= not b;
    layer8_outputs(864) <= not (a xor b);
    layer8_outputs(865) <= a and not b;
    layer8_outputs(866) <= not (a and b);
    layer8_outputs(867) <= a and b;
    layer8_outputs(868) <= b;
    layer8_outputs(869) <= b;
    layer8_outputs(870) <= not b;
    layer8_outputs(871) <= not (a xor b);
    layer8_outputs(872) <= not (a or b);
    layer8_outputs(873) <= b;
    layer8_outputs(874) <= a or b;
    layer8_outputs(875) <= b and not a;
    layer8_outputs(876) <= not (a xor b);
    layer8_outputs(877) <= not b or a;
    layer8_outputs(878) <= 1'b0;
    layer8_outputs(879) <= b;
    layer8_outputs(880) <= not a;
    layer8_outputs(881) <= b and not a;
    layer8_outputs(882) <= not a;
    layer8_outputs(883) <= not b;
    layer8_outputs(884) <= not a;
    layer8_outputs(885) <= not (a and b);
    layer8_outputs(886) <= a xor b;
    layer8_outputs(887) <= b;
    layer8_outputs(888) <= not b;
    layer8_outputs(889) <= not (a or b);
    layer8_outputs(890) <= a xor b;
    layer8_outputs(891) <= a and not b;
    layer8_outputs(892) <= not (a or b);
    layer8_outputs(893) <= not a or b;
    layer8_outputs(894) <= not b;
    layer8_outputs(895) <= a and not b;
    layer8_outputs(896) <= not b or a;
    layer8_outputs(897) <= not a;
    layer8_outputs(898) <= not a;
    layer8_outputs(899) <= a and b;
    layer8_outputs(900) <= not a or b;
    layer8_outputs(901) <= a;
    layer8_outputs(902) <= not b or a;
    layer8_outputs(903) <= a and b;
    layer8_outputs(904) <= not a;
    layer8_outputs(905) <= not a;
    layer8_outputs(906) <= not b;
    layer8_outputs(907) <= a;
    layer8_outputs(908) <= b;
    layer8_outputs(909) <= a or b;
    layer8_outputs(910) <= not (a xor b);
    layer8_outputs(911) <= not b or a;
    layer8_outputs(912) <= a and not b;
    layer8_outputs(913) <= a and not b;
    layer8_outputs(914) <= not (a xor b);
    layer8_outputs(915) <= not b;
    layer8_outputs(916) <= not b;
    layer8_outputs(917) <= not (a and b);
    layer8_outputs(918) <= a xor b;
    layer8_outputs(919) <= not (a xor b);
    layer8_outputs(920) <= not a;
    layer8_outputs(921) <= a and b;
    layer8_outputs(922) <= not (a xor b);
    layer8_outputs(923) <= not (a or b);
    layer8_outputs(924) <= not b;
    layer8_outputs(925) <= a;
    layer8_outputs(926) <= a;
    layer8_outputs(927) <= not b or a;
    layer8_outputs(928) <= not (a xor b);
    layer8_outputs(929) <= not b or a;
    layer8_outputs(930) <= a;
    layer8_outputs(931) <= 1'b1;
    layer8_outputs(932) <= b;
    layer8_outputs(933) <= b and not a;
    layer8_outputs(934) <= a xor b;
    layer8_outputs(935) <= a xor b;
    layer8_outputs(936) <= not a;
    layer8_outputs(937) <= a;
    layer8_outputs(938) <= b;
    layer8_outputs(939) <= not b or a;
    layer8_outputs(940) <= not a or b;
    layer8_outputs(941) <= not (a or b);
    layer8_outputs(942) <= not a;
    layer8_outputs(943) <= 1'b1;
    layer8_outputs(944) <= not (a and b);
    layer8_outputs(945) <= a xor b;
    layer8_outputs(946) <= not a or b;
    layer8_outputs(947) <= not a;
    layer8_outputs(948) <= not (a xor b);
    layer8_outputs(949) <= a xor b;
    layer8_outputs(950) <= b and not a;
    layer8_outputs(951) <= a xor b;
    layer8_outputs(952) <= b and not a;
    layer8_outputs(953) <= not a or b;
    layer8_outputs(954) <= not b or a;
    layer8_outputs(955) <= not b or a;
    layer8_outputs(956) <= a and not b;
    layer8_outputs(957) <= 1'b0;
    layer8_outputs(958) <= not (a and b);
    layer8_outputs(959) <= b and not a;
    layer8_outputs(960) <= not a or b;
    layer8_outputs(961) <= a or b;
    layer8_outputs(962) <= not b;
    layer8_outputs(963) <= a;
    layer8_outputs(964) <= not a;
    layer8_outputs(965) <= not a or b;
    layer8_outputs(966) <= 1'b1;
    layer8_outputs(967) <= b;
    layer8_outputs(968) <= not a;
    layer8_outputs(969) <= a or b;
    layer8_outputs(970) <= not b or a;
    layer8_outputs(971) <= not (a or b);
    layer8_outputs(972) <= not b;
    layer8_outputs(973) <= a or b;
    layer8_outputs(974) <= not (a or b);
    layer8_outputs(975) <= a;
    layer8_outputs(976) <= b and not a;
    layer8_outputs(977) <= not b;
    layer8_outputs(978) <= a;
    layer8_outputs(979) <= not a or b;
    layer8_outputs(980) <= not (a xor b);
    layer8_outputs(981) <= b;
    layer8_outputs(982) <= not a or b;
    layer8_outputs(983) <= not a;
    layer8_outputs(984) <= b;
    layer8_outputs(985) <= a and not b;
    layer8_outputs(986) <= b and not a;
    layer8_outputs(987) <= not b or a;
    layer8_outputs(988) <= b;
    layer8_outputs(989) <= b;
    layer8_outputs(990) <= a and b;
    layer8_outputs(991) <= a;
    layer8_outputs(992) <= b and not a;
    layer8_outputs(993) <= not a;
    layer8_outputs(994) <= not b or a;
    layer8_outputs(995) <= b;
    layer8_outputs(996) <= not a or b;
    layer8_outputs(997) <= not b;
    layer8_outputs(998) <= a;
    layer8_outputs(999) <= a;
    layer8_outputs(1000) <= a;
    layer8_outputs(1001) <= 1'b0;
    layer8_outputs(1002) <= b;
    layer8_outputs(1003) <= b;
    layer8_outputs(1004) <= not (a xor b);
    layer8_outputs(1005) <= a;
    layer8_outputs(1006) <= a;
    layer8_outputs(1007) <= a;
    layer8_outputs(1008) <= b and not a;
    layer8_outputs(1009) <= not a;
    layer8_outputs(1010) <= b and not a;
    layer8_outputs(1011) <= not a;
    layer8_outputs(1012) <= a;
    layer8_outputs(1013) <= a or b;
    layer8_outputs(1014) <= a xor b;
    layer8_outputs(1015) <= not b;
    layer8_outputs(1016) <= not a;
    layer8_outputs(1017) <= not a;
    layer8_outputs(1018) <= a and b;
    layer8_outputs(1019) <= b;
    layer8_outputs(1020) <= not (a xor b);
    layer8_outputs(1021) <= a and b;
    layer8_outputs(1022) <= not b;
    layer8_outputs(1023) <= not b;
    layer8_outputs(1024) <= not b;
    layer8_outputs(1025) <= not a or b;
    layer8_outputs(1026) <= not (a xor b);
    layer8_outputs(1027) <= not b or a;
    layer8_outputs(1028) <= b;
    layer8_outputs(1029) <= not (a and b);
    layer8_outputs(1030) <= not b or a;
    layer8_outputs(1031) <= not (a xor b);
    layer8_outputs(1032) <= b and not a;
    layer8_outputs(1033) <= not (a and b);
    layer8_outputs(1034) <= a;
    layer8_outputs(1035) <= b;
    layer8_outputs(1036) <= a;
    layer8_outputs(1037) <= not (a xor b);
    layer8_outputs(1038) <= not b;
    layer8_outputs(1039) <= b;
    layer8_outputs(1040) <= a xor b;
    layer8_outputs(1041) <= not (a xor b);
    layer8_outputs(1042) <= not a or b;
    layer8_outputs(1043) <= a or b;
    layer8_outputs(1044) <= not (a xor b);
    layer8_outputs(1045) <= not (a and b);
    layer8_outputs(1046) <= not (a xor b);
    layer8_outputs(1047) <= b and not a;
    layer8_outputs(1048) <= b and not a;
    layer8_outputs(1049) <= a xor b;
    layer8_outputs(1050) <= not a;
    layer8_outputs(1051) <= not (a and b);
    layer8_outputs(1052) <= b;
    layer8_outputs(1053) <= not b;
    layer8_outputs(1054) <= not (a xor b);
    layer8_outputs(1055) <= not a;
    layer8_outputs(1056) <= a and not b;
    layer8_outputs(1057) <= not (a xor b);
    layer8_outputs(1058) <= a xor b;
    layer8_outputs(1059) <= a xor b;
    layer8_outputs(1060) <= not b;
    layer8_outputs(1061) <= not a;
    layer8_outputs(1062) <= not (a and b);
    layer8_outputs(1063) <= not b or a;
    layer8_outputs(1064) <= not (a and b);
    layer8_outputs(1065) <= a;
    layer8_outputs(1066) <= not (a and b);
    layer8_outputs(1067) <= a and not b;
    layer8_outputs(1068) <= not a;
    layer8_outputs(1069) <= b;
    layer8_outputs(1070) <= not (a xor b);
    layer8_outputs(1071) <= a and b;
    layer8_outputs(1072) <= not (a or b);
    layer8_outputs(1073) <= not (a or b);
    layer8_outputs(1074) <= a and not b;
    layer8_outputs(1075) <= b;
    layer8_outputs(1076) <= a xor b;
    layer8_outputs(1077) <= a;
    layer8_outputs(1078) <= b;
    layer8_outputs(1079) <= not a;
    layer8_outputs(1080) <= b;
    layer8_outputs(1081) <= a or b;
    layer8_outputs(1082) <= not (a xor b);
    layer8_outputs(1083) <= not (a and b);
    layer8_outputs(1084) <= a and not b;
    layer8_outputs(1085) <= not (a and b);
    layer8_outputs(1086) <= b;
    layer8_outputs(1087) <= not b or a;
    layer8_outputs(1088) <= a or b;
    layer8_outputs(1089) <= a;
    layer8_outputs(1090) <= not b;
    layer8_outputs(1091) <= a;
    layer8_outputs(1092) <= a;
    layer8_outputs(1093) <= a;
    layer8_outputs(1094) <= b and not a;
    layer8_outputs(1095) <= not (a xor b);
    layer8_outputs(1096) <= not (a xor b);
    layer8_outputs(1097) <= not b or a;
    layer8_outputs(1098) <= not a;
    layer8_outputs(1099) <= a;
    layer8_outputs(1100) <= a or b;
    layer8_outputs(1101) <= a and not b;
    layer8_outputs(1102) <= a or b;
    layer8_outputs(1103) <= b;
    layer8_outputs(1104) <= not a;
    layer8_outputs(1105) <= not a;
    layer8_outputs(1106) <= b;
    layer8_outputs(1107) <= a or b;
    layer8_outputs(1108) <= a and b;
    layer8_outputs(1109) <= not (a xor b);
    layer8_outputs(1110) <= b;
    layer8_outputs(1111) <= b;
    layer8_outputs(1112) <= a and not b;
    layer8_outputs(1113) <= not (a and b);
    layer8_outputs(1114) <= not a;
    layer8_outputs(1115) <= not a;
    layer8_outputs(1116) <= not a;
    layer8_outputs(1117) <= b and not a;
    layer8_outputs(1118) <= not (a xor b);
    layer8_outputs(1119) <= not a or b;
    layer8_outputs(1120) <= b;
    layer8_outputs(1121) <= not b or a;
    layer8_outputs(1122) <= not b;
    layer8_outputs(1123) <= a xor b;
    layer8_outputs(1124) <= not (a or b);
    layer8_outputs(1125) <= not (a xor b);
    layer8_outputs(1126) <= b;
    layer8_outputs(1127) <= b and not a;
    layer8_outputs(1128) <= a;
    layer8_outputs(1129) <= a xor b;
    layer8_outputs(1130) <= a;
    layer8_outputs(1131) <= a;
    layer8_outputs(1132) <= not (a and b);
    layer8_outputs(1133) <= not b or a;
    layer8_outputs(1134) <= not (a and b);
    layer8_outputs(1135) <= a xor b;
    layer8_outputs(1136) <= not (a xor b);
    layer8_outputs(1137) <= not a;
    layer8_outputs(1138) <= b;
    layer8_outputs(1139) <= a;
    layer8_outputs(1140) <= a xor b;
    layer8_outputs(1141) <= not (a and b);
    layer8_outputs(1142) <= a;
    layer8_outputs(1143) <= b and not a;
    layer8_outputs(1144) <= not b;
    layer8_outputs(1145) <= a xor b;
    layer8_outputs(1146) <= not b or a;
    layer8_outputs(1147) <= not a or b;
    layer8_outputs(1148) <= not b or a;
    layer8_outputs(1149) <= not b or a;
    layer8_outputs(1150) <= a xor b;
    layer8_outputs(1151) <= not (a xor b);
    layer8_outputs(1152) <= b;
    layer8_outputs(1153) <= b;
    layer8_outputs(1154) <= a and not b;
    layer8_outputs(1155) <= not (a or b);
    layer8_outputs(1156) <= b;
    layer8_outputs(1157) <= b;
    layer8_outputs(1158) <= a xor b;
    layer8_outputs(1159) <= a;
    layer8_outputs(1160) <= not a;
    layer8_outputs(1161) <= not (a or b);
    layer8_outputs(1162) <= b;
    layer8_outputs(1163) <= not a;
    layer8_outputs(1164) <= not b;
    layer8_outputs(1165) <= not (a xor b);
    layer8_outputs(1166) <= a or b;
    layer8_outputs(1167) <= b;
    layer8_outputs(1168) <= a xor b;
    layer8_outputs(1169) <= a xor b;
    layer8_outputs(1170) <= b;
    layer8_outputs(1171) <= b and not a;
    layer8_outputs(1172) <= a;
    layer8_outputs(1173) <= not (a and b);
    layer8_outputs(1174) <= a;
    layer8_outputs(1175) <= not a;
    layer8_outputs(1176) <= a xor b;
    layer8_outputs(1177) <= not (a and b);
    layer8_outputs(1178) <= a;
    layer8_outputs(1179) <= not (a or b);
    layer8_outputs(1180) <= not (a and b);
    layer8_outputs(1181) <= a;
    layer8_outputs(1182) <= not b;
    layer8_outputs(1183) <= a;
    layer8_outputs(1184) <= a;
    layer8_outputs(1185) <= a or b;
    layer8_outputs(1186) <= not (a xor b);
    layer8_outputs(1187) <= not a;
    layer8_outputs(1188) <= a and not b;
    layer8_outputs(1189) <= a xor b;
    layer8_outputs(1190) <= b;
    layer8_outputs(1191) <= not (a xor b);
    layer8_outputs(1192) <= a and b;
    layer8_outputs(1193) <= not (a and b);
    layer8_outputs(1194) <= not (a or b);
    layer8_outputs(1195) <= not (a or b);
    layer8_outputs(1196) <= b;
    layer8_outputs(1197) <= a or b;
    layer8_outputs(1198) <= a;
    layer8_outputs(1199) <= a;
    layer8_outputs(1200) <= a and b;
    layer8_outputs(1201) <= b;
    layer8_outputs(1202) <= not (a xor b);
    layer8_outputs(1203) <= not a;
    layer8_outputs(1204) <= not (a or b);
    layer8_outputs(1205) <= b and not a;
    layer8_outputs(1206) <= b;
    layer8_outputs(1207) <= a or b;
    layer8_outputs(1208) <= not (a or b);
    layer8_outputs(1209) <= not b;
    layer8_outputs(1210) <= b;
    layer8_outputs(1211) <= a;
    layer8_outputs(1212) <= not a;
    layer8_outputs(1213) <= not a or b;
    layer8_outputs(1214) <= not a;
    layer8_outputs(1215) <= not a;
    layer8_outputs(1216) <= not (a xor b);
    layer8_outputs(1217) <= b;
    layer8_outputs(1218) <= not a;
    layer8_outputs(1219) <= not b;
    layer8_outputs(1220) <= a;
    layer8_outputs(1221) <= a xor b;
    layer8_outputs(1222) <= not (a xor b);
    layer8_outputs(1223) <= not (a xor b);
    layer8_outputs(1224) <= not (a xor b);
    layer8_outputs(1225) <= not b;
    layer8_outputs(1226) <= not (a or b);
    layer8_outputs(1227) <= not (a and b);
    layer8_outputs(1228) <= a;
    layer8_outputs(1229) <= a xor b;
    layer8_outputs(1230) <= not a or b;
    layer8_outputs(1231) <= a;
    layer8_outputs(1232) <= a;
    layer8_outputs(1233) <= not b;
    layer8_outputs(1234) <= a and not b;
    layer8_outputs(1235) <= a and b;
    layer8_outputs(1236) <= not b or a;
    layer8_outputs(1237) <= a xor b;
    layer8_outputs(1238) <= not b or a;
    layer8_outputs(1239) <= not (a or b);
    layer8_outputs(1240) <= not a or b;
    layer8_outputs(1241) <= a;
    layer8_outputs(1242) <= a xor b;
    layer8_outputs(1243) <= a;
    layer8_outputs(1244) <= a and not b;
    layer8_outputs(1245) <= not (a xor b);
    layer8_outputs(1246) <= not b;
    layer8_outputs(1247) <= not (a xor b);
    layer8_outputs(1248) <= a and b;
    layer8_outputs(1249) <= not (a and b);
    layer8_outputs(1250) <= not (a and b);
    layer8_outputs(1251) <= not a;
    layer8_outputs(1252) <= not (a or b);
    layer8_outputs(1253) <= not (a xor b);
    layer8_outputs(1254) <= b;
    layer8_outputs(1255) <= not a or b;
    layer8_outputs(1256) <= not (a xor b);
    layer8_outputs(1257) <= not (a or b);
    layer8_outputs(1258) <= b and not a;
    layer8_outputs(1259) <= not a;
    layer8_outputs(1260) <= b and not a;
    layer8_outputs(1261) <= not b;
    layer8_outputs(1262) <= a;
    layer8_outputs(1263) <= b;
    layer8_outputs(1264) <= a and not b;
    layer8_outputs(1265) <= a or b;
    layer8_outputs(1266) <= not (a or b);
    layer8_outputs(1267) <= a xor b;
    layer8_outputs(1268) <= not a or b;
    layer8_outputs(1269) <= not b;
    layer8_outputs(1270) <= not b;
    layer8_outputs(1271) <= not a;
    layer8_outputs(1272) <= not a;
    layer8_outputs(1273) <= not a or b;
    layer8_outputs(1274) <= a;
    layer8_outputs(1275) <= not a;
    layer8_outputs(1276) <= not b;
    layer8_outputs(1277) <= a xor b;
    layer8_outputs(1278) <= not (a or b);
    layer8_outputs(1279) <= not (a xor b);
    layer8_outputs(1280) <= not b;
    layer8_outputs(1281) <= not a;
    layer8_outputs(1282) <= not (a and b);
    layer8_outputs(1283) <= not b;
    layer8_outputs(1284) <= a and b;
    layer8_outputs(1285) <= a xor b;
    layer8_outputs(1286) <= not a;
    layer8_outputs(1287) <= not (a or b);
    layer8_outputs(1288) <= a and b;
    layer8_outputs(1289) <= not (a and b);
    layer8_outputs(1290) <= not a or b;
    layer8_outputs(1291) <= a xor b;
    layer8_outputs(1292) <= not b or a;
    layer8_outputs(1293) <= a and b;
    layer8_outputs(1294) <= a and not b;
    layer8_outputs(1295) <= b;
    layer8_outputs(1296) <= not (a and b);
    layer8_outputs(1297) <= a xor b;
    layer8_outputs(1298) <= b and not a;
    layer8_outputs(1299) <= not (a xor b);
    layer8_outputs(1300) <= b;
    layer8_outputs(1301) <= a;
    layer8_outputs(1302) <= a;
    layer8_outputs(1303) <= not (a xor b);
    layer8_outputs(1304) <= not (a or b);
    layer8_outputs(1305) <= b;
    layer8_outputs(1306) <= a xor b;
    layer8_outputs(1307) <= not b;
    layer8_outputs(1308) <= not a;
    layer8_outputs(1309) <= not (a and b);
    layer8_outputs(1310) <= not a or b;
    layer8_outputs(1311) <= a xor b;
    layer8_outputs(1312) <= not (a xor b);
    layer8_outputs(1313) <= a;
    layer8_outputs(1314) <= not a;
    layer8_outputs(1315) <= a;
    layer8_outputs(1316) <= not (a or b);
    layer8_outputs(1317) <= not b;
    layer8_outputs(1318) <= b;
    layer8_outputs(1319) <= b;
    layer8_outputs(1320) <= b;
    layer8_outputs(1321) <= b and not a;
    layer8_outputs(1322) <= not a;
    layer8_outputs(1323) <= not (a or b);
    layer8_outputs(1324) <= a;
    layer8_outputs(1325) <= a or b;
    layer8_outputs(1326) <= b;
    layer8_outputs(1327) <= a or b;
    layer8_outputs(1328) <= not b or a;
    layer8_outputs(1329) <= not (a or b);
    layer8_outputs(1330) <= not a;
    layer8_outputs(1331) <= a xor b;
    layer8_outputs(1332) <= b;
    layer8_outputs(1333) <= not (a or b);
    layer8_outputs(1334) <= not (a and b);
    layer8_outputs(1335) <= not b or a;
    layer8_outputs(1336) <= not b or a;
    layer8_outputs(1337) <= b and not a;
    layer8_outputs(1338) <= a or b;
    layer8_outputs(1339) <= a and b;
    layer8_outputs(1340) <= a xor b;
    layer8_outputs(1341) <= not a;
    layer8_outputs(1342) <= not a;
    layer8_outputs(1343) <= b and not a;
    layer8_outputs(1344) <= a xor b;
    layer8_outputs(1345) <= a;
    layer8_outputs(1346) <= not b;
    layer8_outputs(1347) <= a xor b;
    layer8_outputs(1348) <= not (a or b);
    layer8_outputs(1349) <= not (a xor b);
    layer8_outputs(1350) <= 1'b0;
    layer8_outputs(1351) <= not a;
    layer8_outputs(1352) <= not b;
    layer8_outputs(1353) <= not a;
    layer8_outputs(1354) <= a and b;
    layer8_outputs(1355) <= a;
    layer8_outputs(1356) <= not b;
    layer8_outputs(1357) <= b;
    layer8_outputs(1358) <= not (a xor b);
    layer8_outputs(1359) <= not (a or b);
    layer8_outputs(1360) <= not (a and b);
    layer8_outputs(1361) <= b and not a;
    layer8_outputs(1362) <= not b;
    layer8_outputs(1363) <= a xor b;
    layer8_outputs(1364) <= a xor b;
    layer8_outputs(1365) <= b;
    layer8_outputs(1366) <= not (a or b);
    layer8_outputs(1367) <= 1'b0;
    layer8_outputs(1368) <= not (a xor b);
    layer8_outputs(1369) <= not b or a;
    layer8_outputs(1370) <= not a;
    layer8_outputs(1371) <= not (a xor b);
    layer8_outputs(1372) <= a and b;
    layer8_outputs(1373) <= a;
    layer8_outputs(1374) <= not a;
    layer8_outputs(1375) <= not b or a;
    layer8_outputs(1376) <= not (a xor b);
    layer8_outputs(1377) <= b;
    layer8_outputs(1378) <= not b or a;
    layer8_outputs(1379) <= b;
    layer8_outputs(1380) <= not a;
    layer8_outputs(1381) <= not b;
    layer8_outputs(1382) <= not a;
    layer8_outputs(1383) <= a or b;
    layer8_outputs(1384) <= not b;
    layer8_outputs(1385) <= not b;
    layer8_outputs(1386) <= a and not b;
    layer8_outputs(1387) <= b;
    layer8_outputs(1388) <= not a;
    layer8_outputs(1389) <= not b or a;
    layer8_outputs(1390) <= not a or b;
    layer8_outputs(1391) <= 1'b1;
    layer8_outputs(1392) <= not a or b;
    layer8_outputs(1393) <= b;
    layer8_outputs(1394) <= not a;
    layer8_outputs(1395) <= not a or b;
    layer8_outputs(1396) <= a and not b;
    layer8_outputs(1397) <= not a;
    layer8_outputs(1398) <= not a;
    layer8_outputs(1399) <= not a;
    layer8_outputs(1400) <= not b;
    layer8_outputs(1401) <= not (a xor b);
    layer8_outputs(1402) <= b and not a;
    layer8_outputs(1403) <= a;
    layer8_outputs(1404) <= not b;
    layer8_outputs(1405) <= a xor b;
    layer8_outputs(1406) <= not b;
    layer8_outputs(1407) <= not a or b;
    layer8_outputs(1408) <= not (a and b);
    layer8_outputs(1409) <= not (a and b);
    layer8_outputs(1410) <= a xor b;
    layer8_outputs(1411) <= not (a or b);
    layer8_outputs(1412) <= not a or b;
    layer8_outputs(1413) <= not b;
    layer8_outputs(1414) <= not a;
    layer8_outputs(1415) <= not a;
    layer8_outputs(1416) <= a or b;
    layer8_outputs(1417) <= not (a or b);
    layer8_outputs(1418) <= b and not a;
    layer8_outputs(1419) <= b;
    layer8_outputs(1420) <= b and not a;
    layer8_outputs(1421) <= not a or b;
    layer8_outputs(1422) <= not b or a;
    layer8_outputs(1423) <= a or b;
    layer8_outputs(1424) <= b and not a;
    layer8_outputs(1425) <= not b;
    layer8_outputs(1426) <= not a;
    layer8_outputs(1427) <= not b;
    layer8_outputs(1428) <= b;
    layer8_outputs(1429) <= a;
    layer8_outputs(1430) <= not a;
    layer8_outputs(1431) <= a and not b;
    layer8_outputs(1432) <= b;
    layer8_outputs(1433) <= not b;
    layer8_outputs(1434) <= b;
    layer8_outputs(1435) <= not b or a;
    layer8_outputs(1436) <= not a;
    layer8_outputs(1437) <= a and b;
    layer8_outputs(1438) <= not b;
    layer8_outputs(1439) <= not b or a;
    layer8_outputs(1440) <= b and not a;
    layer8_outputs(1441) <= a;
    layer8_outputs(1442) <= not a or b;
    layer8_outputs(1443) <= not b;
    layer8_outputs(1444) <= not (a xor b);
    layer8_outputs(1445) <= a and not b;
    layer8_outputs(1446) <= a xor b;
    layer8_outputs(1447) <= not b;
    layer8_outputs(1448) <= not (a or b);
    layer8_outputs(1449) <= not a or b;
    layer8_outputs(1450) <= b and not a;
    layer8_outputs(1451) <= b;
    layer8_outputs(1452) <= not (a xor b);
    layer8_outputs(1453) <= not (a and b);
    layer8_outputs(1454) <= not (a and b);
    layer8_outputs(1455) <= b;
    layer8_outputs(1456) <= not a;
    layer8_outputs(1457) <= not b;
    layer8_outputs(1458) <= not a;
    layer8_outputs(1459) <= not a;
    layer8_outputs(1460) <= a;
    layer8_outputs(1461) <= a and b;
    layer8_outputs(1462) <= b and not a;
    layer8_outputs(1463) <= b;
    layer8_outputs(1464) <= not b;
    layer8_outputs(1465) <= a and b;
    layer8_outputs(1466) <= b;
    layer8_outputs(1467) <= not a;
    layer8_outputs(1468) <= not (a or b);
    layer8_outputs(1469) <= not (a xor b);
    layer8_outputs(1470) <= a;
    layer8_outputs(1471) <= 1'b0;
    layer8_outputs(1472) <= a;
    layer8_outputs(1473) <= not (a xor b);
    layer8_outputs(1474) <= not a or b;
    layer8_outputs(1475) <= a and not b;
    layer8_outputs(1476) <= a and not b;
    layer8_outputs(1477) <= not (a and b);
    layer8_outputs(1478) <= b and not a;
    layer8_outputs(1479) <= not (a xor b);
    layer8_outputs(1480) <= not (a and b);
    layer8_outputs(1481) <= not (a and b);
    layer8_outputs(1482) <= not a;
    layer8_outputs(1483) <= not (a xor b);
    layer8_outputs(1484) <= a and not b;
    layer8_outputs(1485) <= b;
    layer8_outputs(1486) <= not a or b;
    layer8_outputs(1487) <= b;
    layer8_outputs(1488) <= b;
    layer8_outputs(1489) <= b and not a;
    layer8_outputs(1490) <= not b;
    layer8_outputs(1491) <= a xor b;
    layer8_outputs(1492) <= not a;
    layer8_outputs(1493) <= not (a xor b);
    layer8_outputs(1494) <= b;
    layer8_outputs(1495) <= not b;
    layer8_outputs(1496) <= not (a or b);
    layer8_outputs(1497) <= b;
    layer8_outputs(1498) <= a and not b;
    layer8_outputs(1499) <= not (a xor b);
    layer8_outputs(1500) <= not (a and b);
    layer8_outputs(1501) <= a xor b;
    layer8_outputs(1502) <= a;
    layer8_outputs(1503) <= b;
    layer8_outputs(1504) <= a;
    layer8_outputs(1505) <= a xor b;
    layer8_outputs(1506) <= 1'b0;
    layer8_outputs(1507) <= a or b;
    layer8_outputs(1508) <= not (a or b);
    layer8_outputs(1509) <= not a or b;
    layer8_outputs(1510) <= b and not a;
    layer8_outputs(1511) <= b and not a;
    layer8_outputs(1512) <= a or b;
    layer8_outputs(1513) <= b;
    layer8_outputs(1514) <= not a;
    layer8_outputs(1515) <= a;
    layer8_outputs(1516) <= not (a xor b);
    layer8_outputs(1517) <= a and b;
    layer8_outputs(1518) <= not (a and b);
    layer8_outputs(1519) <= not a;
    layer8_outputs(1520) <= 1'b0;
    layer8_outputs(1521) <= not (a xor b);
    layer8_outputs(1522) <= not b;
    layer8_outputs(1523) <= not b;
    layer8_outputs(1524) <= a;
    layer8_outputs(1525) <= a and not b;
    layer8_outputs(1526) <= b;
    layer8_outputs(1527) <= a xor b;
    layer8_outputs(1528) <= a;
    layer8_outputs(1529) <= a and b;
    layer8_outputs(1530) <= not b;
    layer8_outputs(1531) <= not (a xor b);
    layer8_outputs(1532) <= a xor b;
    layer8_outputs(1533) <= not a;
    layer8_outputs(1534) <= not a;
    layer8_outputs(1535) <= b;
    layer8_outputs(1536) <= not a;
    layer8_outputs(1537) <= a or b;
    layer8_outputs(1538) <= a and b;
    layer8_outputs(1539) <= not a or b;
    layer8_outputs(1540) <= not a;
    layer8_outputs(1541) <= not b;
    layer8_outputs(1542) <= not b;
    layer8_outputs(1543) <= a and not b;
    layer8_outputs(1544) <= b and not a;
    layer8_outputs(1545) <= a and b;
    layer8_outputs(1546) <= a and not b;
    layer8_outputs(1547) <= a or b;
    layer8_outputs(1548) <= a;
    layer8_outputs(1549) <= not b or a;
    layer8_outputs(1550) <= not (a xor b);
    layer8_outputs(1551) <= b;
    layer8_outputs(1552) <= not a;
    layer8_outputs(1553) <= not b;
    layer8_outputs(1554) <= a and b;
    layer8_outputs(1555) <= not a;
    layer8_outputs(1556) <= not a;
    layer8_outputs(1557) <= b;
    layer8_outputs(1558) <= a or b;
    layer8_outputs(1559) <= not b or a;
    layer8_outputs(1560) <= not (a xor b);
    layer8_outputs(1561) <= not b or a;
    layer8_outputs(1562) <= not a;
    layer8_outputs(1563) <= not (a xor b);
    layer8_outputs(1564) <= not a;
    layer8_outputs(1565) <= a xor b;
    layer8_outputs(1566) <= b and not a;
    layer8_outputs(1567) <= b and not a;
    layer8_outputs(1568) <= a xor b;
    layer8_outputs(1569) <= not (a or b);
    layer8_outputs(1570) <= a xor b;
    layer8_outputs(1571) <= a and not b;
    layer8_outputs(1572) <= not a or b;
    layer8_outputs(1573) <= 1'b0;
    layer8_outputs(1574) <= b and not a;
    layer8_outputs(1575) <= a and b;
    layer8_outputs(1576) <= b;
    layer8_outputs(1577) <= not a;
    layer8_outputs(1578) <= a xor b;
    layer8_outputs(1579) <= not b;
    layer8_outputs(1580) <= a xor b;
    layer8_outputs(1581) <= not (a xor b);
    layer8_outputs(1582) <= a;
    layer8_outputs(1583) <= b;
    layer8_outputs(1584) <= not a;
    layer8_outputs(1585) <= not (a and b);
    layer8_outputs(1586) <= not (a or b);
    layer8_outputs(1587) <= not (a and b);
    layer8_outputs(1588) <= a xor b;
    layer8_outputs(1589) <= not a or b;
    layer8_outputs(1590) <= not (a xor b);
    layer8_outputs(1591) <= not (a xor b);
    layer8_outputs(1592) <= a and not b;
    layer8_outputs(1593) <= not b;
    layer8_outputs(1594) <= not a;
    layer8_outputs(1595) <= not a or b;
    layer8_outputs(1596) <= a and b;
    layer8_outputs(1597) <= a;
    layer8_outputs(1598) <= not (a xor b);
    layer8_outputs(1599) <= not (a or b);
    layer8_outputs(1600) <= not (a and b);
    layer8_outputs(1601) <= a or b;
    layer8_outputs(1602) <= a xor b;
    layer8_outputs(1603) <= b;
    layer8_outputs(1604) <= not a;
    layer8_outputs(1605) <= b;
    layer8_outputs(1606) <= not a;
    layer8_outputs(1607) <= not a or b;
    layer8_outputs(1608) <= a;
    layer8_outputs(1609) <= not (a or b);
    layer8_outputs(1610) <= b;
    layer8_outputs(1611) <= b;
    layer8_outputs(1612) <= not b or a;
    layer8_outputs(1613) <= not a;
    layer8_outputs(1614) <= not (a xor b);
    layer8_outputs(1615) <= not (a or b);
    layer8_outputs(1616) <= a or b;
    layer8_outputs(1617) <= b;
    layer8_outputs(1618) <= a;
    layer8_outputs(1619) <= not (a and b);
    layer8_outputs(1620) <= a xor b;
    layer8_outputs(1621) <= not b;
    layer8_outputs(1622) <= b and not a;
    layer8_outputs(1623) <= not (a and b);
    layer8_outputs(1624) <= not a;
    layer8_outputs(1625) <= not b or a;
    layer8_outputs(1626) <= b and not a;
    layer8_outputs(1627) <= a xor b;
    layer8_outputs(1628) <= a;
    layer8_outputs(1629) <= not b or a;
    layer8_outputs(1630) <= a;
    layer8_outputs(1631) <= b;
    layer8_outputs(1632) <= a and not b;
    layer8_outputs(1633) <= a;
    layer8_outputs(1634) <= not a;
    layer8_outputs(1635) <= not b;
    layer8_outputs(1636) <= b;
    layer8_outputs(1637) <= b and not a;
    layer8_outputs(1638) <= a and not b;
    layer8_outputs(1639) <= not b or a;
    layer8_outputs(1640) <= b and not a;
    layer8_outputs(1641) <= a xor b;
    layer8_outputs(1642) <= not (a or b);
    layer8_outputs(1643) <= not (a xor b);
    layer8_outputs(1644) <= not a;
    layer8_outputs(1645) <= a;
    layer8_outputs(1646) <= a and b;
    layer8_outputs(1647) <= b;
    layer8_outputs(1648) <= not a;
    layer8_outputs(1649) <= b;
    layer8_outputs(1650) <= not b;
    layer8_outputs(1651) <= a xor b;
    layer8_outputs(1652) <= a xor b;
    layer8_outputs(1653) <= a;
    layer8_outputs(1654) <= not b;
    layer8_outputs(1655) <= not b or a;
    layer8_outputs(1656) <= not a;
    layer8_outputs(1657) <= b;
    layer8_outputs(1658) <= not (a and b);
    layer8_outputs(1659) <= 1'b1;
    layer8_outputs(1660) <= not a or b;
    layer8_outputs(1661) <= not (a or b);
    layer8_outputs(1662) <= not b or a;
    layer8_outputs(1663) <= not (a and b);
    layer8_outputs(1664) <= not a;
    layer8_outputs(1665) <= a and b;
    layer8_outputs(1666) <= a or b;
    layer8_outputs(1667) <= a xor b;
    layer8_outputs(1668) <= not a;
    layer8_outputs(1669) <= b and not a;
    layer8_outputs(1670) <= not b;
    layer8_outputs(1671) <= b and not a;
    layer8_outputs(1672) <= not b or a;
    layer8_outputs(1673) <= not (a or b);
    layer8_outputs(1674) <= not (a xor b);
    layer8_outputs(1675) <= not b;
    layer8_outputs(1676) <= a and not b;
    layer8_outputs(1677) <= a or b;
    layer8_outputs(1678) <= not (a xor b);
    layer8_outputs(1679) <= a and b;
    layer8_outputs(1680) <= a;
    layer8_outputs(1681) <= a and not b;
    layer8_outputs(1682) <= not a;
    layer8_outputs(1683) <= b;
    layer8_outputs(1684) <= not b or a;
    layer8_outputs(1685) <= a and not b;
    layer8_outputs(1686) <= a xor b;
    layer8_outputs(1687) <= not b;
    layer8_outputs(1688) <= a and not b;
    layer8_outputs(1689) <= not b or a;
    layer8_outputs(1690) <= b and not a;
    layer8_outputs(1691) <= not a or b;
    layer8_outputs(1692) <= b;
    layer8_outputs(1693) <= not (a and b);
    layer8_outputs(1694) <= not b or a;
    layer8_outputs(1695) <= b;
    layer8_outputs(1696) <= not (a or b);
    layer8_outputs(1697) <= not b or a;
    layer8_outputs(1698) <= not (a xor b);
    layer8_outputs(1699) <= b;
    layer8_outputs(1700) <= not a;
    layer8_outputs(1701) <= not a or b;
    layer8_outputs(1702) <= a and not b;
    layer8_outputs(1703) <= not a;
    layer8_outputs(1704) <= a;
    layer8_outputs(1705) <= a xor b;
    layer8_outputs(1706) <= b;
    layer8_outputs(1707) <= not (a and b);
    layer8_outputs(1708) <= not a or b;
    layer8_outputs(1709) <= not b;
    layer8_outputs(1710) <= b;
    layer8_outputs(1711) <= not a;
    layer8_outputs(1712) <= b;
    layer8_outputs(1713) <= a;
    layer8_outputs(1714) <= not (a xor b);
    layer8_outputs(1715) <= a xor b;
    layer8_outputs(1716) <= a xor b;
    layer8_outputs(1717) <= a xor b;
    layer8_outputs(1718) <= a xor b;
    layer8_outputs(1719) <= a;
    layer8_outputs(1720) <= not (a xor b);
    layer8_outputs(1721) <= not b or a;
    layer8_outputs(1722) <= not (a or b);
    layer8_outputs(1723) <= not b;
    layer8_outputs(1724) <= b;
    layer8_outputs(1725) <= not b;
    layer8_outputs(1726) <= a xor b;
    layer8_outputs(1727) <= not a;
    layer8_outputs(1728) <= a xor b;
    layer8_outputs(1729) <= a or b;
    layer8_outputs(1730) <= a xor b;
    layer8_outputs(1731) <= b and not a;
    layer8_outputs(1732) <= not a;
    layer8_outputs(1733) <= a;
    layer8_outputs(1734) <= b and not a;
    layer8_outputs(1735) <= not a;
    layer8_outputs(1736) <= a;
    layer8_outputs(1737) <= a and not b;
    layer8_outputs(1738) <= not a;
    layer8_outputs(1739) <= a;
    layer8_outputs(1740) <= a;
    layer8_outputs(1741) <= not (a and b);
    layer8_outputs(1742) <= not a or b;
    layer8_outputs(1743) <= a xor b;
    layer8_outputs(1744) <= not a;
    layer8_outputs(1745) <= a xor b;
    layer8_outputs(1746) <= a and not b;
    layer8_outputs(1747) <= not (a or b);
    layer8_outputs(1748) <= a;
    layer8_outputs(1749) <= not b;
    layer8_outputs(1750) <= b and not a;
    layer8_outputs(1751) <= not (a or b);
    layer8_outputs(1752) <= not (a xor b);
    layer8_outputs(1753) <= not (a and b);
    layer8_outputs(1754) <= not b;
    layer8_outputs(1755) <= a and not b;
    layer8_outputs(1756) <= b;
    layer8_outputs(1757) <= not b;
    layer8_outputs(1758) <= not a;
    layer8_outputs(1759) <= not a or b;
    layer8_outputs(1760) <= not b;
    layer8_outputs(1761) <= not a or b;
    layer8_outputs(1762) <= not (a or b);
    layer8_outputs(1763) <= not a;
    layer8_outputs(1764) <= b;
    layer8_outputs(1765) <= not a;
    layer8_outputs(1766) <= a and not b;
    layer8_outputs(1767) <= not a;
    layer8_outputs(1768) <= not a or b;
    layer8_outputs(1769) <= b;
    layer8_outputs(1770) <= not a or b;
    layer8_outputs(1771) <= not b or a;
    layer8_outputs(1772) <= b and not a;
    layer8_outputs(1773) <= a xor b;
    layer8_outputs(1774) <= not a or b;
    layer8_outputs(1775) <= not a;
    layer8_outputs(1776) <= a or b;
    layer8_outputs(1777) <= a xor b;
    layer8_outputs(1778) <= not b or a;
    layer8_outputs(1779) <= a or b;
    layer8_outputs(1780) <= b;
    layer8_outputs(1781) <= not b;
    layer8_outputs(1782) <= not (a xor b);
    layer8_outputs(1783) <= a;
    layer8_outputs(1784) <= not a;
    layer8_outputs(1785) <= not b;
    layer8_outputs(1786) <= a and b;
    layer8_outputs(1787) <= not (a or b);
    layer8_outputs(1788) <= b;
    layer8_outputs(1789) <= not b;
    layer8_outputs(1790) <= not (a or b);
    layer8_outputs(1791) <= a and b;
    layer8_outputs(1792) <= not b or a;
    layer8_outputs(1793) <= a;
    layer8_outputs(1794) <= a xor b;
    layer8_outputs(1795) <= a or b;
    layer8_outputs(1796) <= 1'b1;
    layer8_outputs(1797) <= a xor b;
    layer8_outputs(1798) <= a or b;
    layer8_outputs(1799) <= b;
    layer8_outputs(1800) <= a;
    layer8_outputs(1801) <= not b or a;
    layer8_outputs(1802) <= a or b;
    layer8_outputs(1803) <= not a;
    layer8_outputs(1804) <= 1'b0;
    layer8_outputs(1805) <= a xor b;
    layer8_outputs(1806) <= not (a or b);
    layer8_outputs(1807) <= not (a xor b);
    layer8_outputs(1808) <= not (a xor b);
    layer8_outputs(1809) <= not a;
    layer8_outputs(1810) <= b;
    layer8_outputs(1811) <= a xor b;
    layer8_outputs(1812) <= a or b;
    layer8_outputs(1813) <= not a;
    layer8_outputs(1814) <= a;
    layer8_outputs(1815) <= not a;
    layer8_outputs(1816) <= not a;
    layer8_outputs(1817) <= b;
    layer8_outputs(1818) <= not b or a;
    layer8_outputs(1819) <= not (a or b);
    layer8_outputs(1820) <= b;
    layer8_outputs(1821) <= a;
    layer8_outputs(1822) <= not a;
    layer8_outputs(1823) <= not a;
    layer8_outputs(1824) <= a;
    layer8_outputs(1825) <= not a or b;
    layer8_outputs(1826) <= not (a xor b);
    layer8_outputs(1827) <= not b or a;
    layer8_outputs(1828) <= not (a xor b);
    layer8_outputs(1829) <= not a;
    layer8_outputs(1830) <= not (a or b);
    layer8_outputs(1831) <= a and not b;
    layer8_outputs(1832) <= b;
    layer8_outputs(1833) <= not a;
    layer8_outputs(1834) <= not b or a;
    layer8_outputs(1835) <= not (a and b);
    layer8_outputs(1836) <= not (a and b);
    layer8_outputs(1837) <= not a;
    layer8_outputs(1838) <= not (a or b);
    layer8_outputs(1839) <= not b;
    layer8_outputs(1840) <= a;
    layer8_outputs(1841) <= a;
    layer8_outputs(1842) <= not (a and b);
    layer8_outputs(1843) <= not a;
    layer8_outputs(1844) <= b;
    layer8_outputs(1845) <= b and not a;
    layer8_outputs(1846) <= not a;
    layer8_outputs(1847) <= not a;
    layer8_outputs(1848) <= not (a and b);
    layer8_outputs(1849) <= not (a or b);
    layer8_outputs(1850) <= not a;
    layer8_outputs(1851) <= a xor b;
    layer8_outputs(1852) <= not (a xor b);
    layer8_outputs(1853) <= not b;
    layer8_outputs(1854) <= not b;
    layer8_outputs(1855) <= not b;
    layer8_outputs(1856) <= a xor b;
    layer8_outputs(1857) <= not b;
    layer8_outputs(1858) <= b;
    layer8_outputs(1859) <= not (a or b);
    layer8_outputs(1860) <= not a;
    layer8_outputs(1861) <= a or b;
    layer8_outputs(1862) <= not (a xor b);
    layer8_outputs(1863) <= not a;
    layer8_outputs(1864) <= a or b;
    layer8_outputs(1865) <= not (a or b);
    layer8_outputs(1866) <= not a or b;
    layer8_outputs(1867) <= a and not b;
    layer8_outputs(1868) <= not (a xor b);
    layer8_outputs(1869) <= a xor b;
    layer8_outputs(1870) <= not b;
    layer8_outputs(1871) <= not (a xor b);
    layer8_outputs(1872) <= a;
    layer8_outputs(1873) <= b;
    layer8_outputs(1874) <= a and not b;
    layer8_outputs(1875) <= not b or a;
    layer8_outputs(1876) <= not b;
    layer8_outputs(1877) <= a xor b;
    layer8_outputs(1878) <= a xor b;
    layer8_outputs(1879) <= not b;
    layer8_outputs(1880) <= not b or a;
    layer8_outputs(1881) <= not a;
    layer8_outputs(1882) <= not b;
    layer8_outputs(1883) <= a or b;
    layer8_outputs(1884) <= a;
    layer8_outputs(1885) <= not (a xor b);
    layer8_outputs(1886) <= not (a xor b);
    layer8_outputs(1887) <= not (a and b);
    layer8_outputs(1888) <= not a or b;
    layer8_outputs(1889) <= a and b;
    layer8_outputs(1890) <= not (a xor b);
    layer8_outputs(1891) <= not (a xor b);
    layer8_outputs(1892) <= not b;
    layer8_outputs(1893) <= a xor b;
    layer8_outputs(1894) <= not a or b;
    layer8_outputs(1895) <= b;
    layer8_outputs(1896) <= not a or b;
    layer8_outputs(1897) <= a and not b;
    layer8_outputs(1898) <= not (a xor b);
    layer8_outputs(1899) <= not b;
    layer8_outputs(1900) <= b;
    layer8_outputs(1901) <= a;
    layer8_outputs(1902) <= not a;
    layer8_outputs(1903) <= not (a or b);
    layer8_outputs(1904) <= not a;
    layer8_outputs(1905) <= a and b;
    layer8_outputs(1906) <= a xor b;
    layer8_outputs(1907) <= a;
    layer8_outputs(1908) <= not b;
    layer8_outputs(1909) <= not b or a;
    layer8_outputs(1910) <= b;
    layer8_outputs(1911) <= not (a xor b);
    layer8_outputs(1912) <= a;
    layer8_outputs(1913) <= not b or a;
    layer8_outputs(1914) <= not b or a;
    layer8_outputs(1915) <= a and b;
    layer8_outputs(1916) <= a xor b;
    layer8_outputs(1917) <= not b or a;
    layer8_outputs(1918) <= not b;
    layer8_outputs(1919) <= not b;
    layer8_outputs(1920) <= not a;
    layer8_outputs(1921) <= a;
    layer8_outputs(1922) <= a xor b;
    layer8_outputs(1923) <= not b or a;
    layer8_outputs(1924) <= not a;
    layer8_outputs(1925) <= not a or b;
    layer8_outputs(1926) <= a and b;
    layer8_outputs(1927) <= not b;
    layer8_outputs(1928) <= a xor b;
    layer8_outputs(1929) <= b;
    layer8_outputs(1930) <= not (a and b);
    layer8_outputs(1931) <= not a;
    layer8_outputs(1932) <= b;
    layer8_outputs(1933) <= not a or b;
    layer8_outputs(1934) <= a;
    layer8_outputs(1935) <= not (a and b);
    layer8_outputs(1936) <= b;
    layer8_outputs(1937) <= b;
    layer8_outputs(1938) <= not a;
    layer8_outputs(1939) <= a;
    layer8_outputs(1940) <= a or b;
    layer8_outputs(1941) <= a and b;
    layer8_outputs(1942) <= b and not a;
    layer8_outputs(1943) <= a;
    layer8_outputs(1944) <= not (a or b);
    layer8_outputs(1945) <= not (a xor b);
    layer8_outputs(1946) <= 1'b0;
    layer8_outputs(1947) <= a;
    layer8_outputs(1948) <= b;
    layer8_outputs(1949) <= not (a xor b);
    layer8_outputs(1950) <= not a;
    layer8_outputs(1951) <= not a;
    layer8_outputs(1952) <= not b;
    layer8_outputs(1953) <= a;
    layer8_outputs(1954) <= not a or b;
    layer8_outputs(1955) <= a xor b;
    layer8_outputs(1956) <= not a;
    layer8_outputs(1957) <= not b or a;
    layer8_outputs(1958) <= b;
    layer8_outputs(1959) <= not a;
    layer8_outputs(1960) <= not (a and b);
    layer8_outputs(1961) <= a and b;
    layer8_outputs(1962) <= b;
    layer8_outputs(1963) <= a;
    layer8_outputs(1964) <= not b or a;
    layer8_outputs(1965) <= a or b;
    layer8_outputs(1966) <= a xor b;
    layer8_outputs(1967) <= b and not a;
    layer8_outputs(1968) <= a;
    layer8_outputs(1969) <= not a or b;
    layer8_outputs(1970) <= a;
    layer8_outputs(1971) <= not b;
    layer8_outputs(1972) <= a xor b;
    layer8_outputs(1973) <= not a or b;
    layer8_outputs(1974) <= not (a and b);
    layer8_outputs(1975) <= not b;
    layer8_outputs(1976) <= not a;
    layer8_outputs(1977) <= b and not a;
    layer8_outputs(1978) <= b;
    layer8_outputs(1979) <= not (a and b);
    layer8_outputs(1980) <= a;
    layer8_outputs(1981) <= 1'b1;
    layer8_outputs(1982) <= not (a and b);
    layer8_outputs(1983) <= a and b;
    layer8_outputs(1984) <= 1'b1;
    layer8_outputs(1985) <= not b;
    layer8_outputs(1986) <= a;
    layer8_outputs(1987) <= not b or a;
    layer8_outputs(1988) <= a and b;
    layer8_outputs(1989) <= not b;
    layer8_outputs(1990) <= not a or b;
    layer8_outputs(1991) <= a;
    layer8_outputs(1992) <= b;
    layer8_outputs(1993) <= not a or b;
    layer8_outputs(1994) <= not b;
    layer8_outputs(1995) <= not b;
    layer8_outputs(1996) <= a;
    layer8_outputs(1997) <= a or b;
    layer8_outputs(1998) <= b;
    layer8_outputs(1999) <= not a or b;
    layer8_outputs(2000) <= b;
    layer8_outputs(2001) <= not a or b;
    layer8_outputs(2002) <= a and b;
    layer8_outputs(2003) <= a;
    layer8_outputs(2004) <= not a or b;
    layer8_outputs(2005) <= not a;
    layer8_outputs(2006) <= a and b;
    layer8_outputs(2007) <= a and not b;
    layer8_outputs(2008) <= a xor b;
    layer8_outputs(2009) <= a;
    layer8_outputs(2010) <= a xor b;
    layer8_outputs(2011) <= not (a or b);
    layer8_outputs(2012) <= a and not b;
    layer8_outputs(2013) <= a and b;
    layer8_outputs(2014) <= b;
    layer8_outputs(2015) <= not a;
    layer8_outputs(2016) <= not (a and b);
    layer8_outputs(2017) <= 1'b1;
    layer8_outputs(2018) <= a;
    layer8_outputs(2019) <= a xor b;
    layer8_outputs(2020) <= a xor b;
    layer8_outputs(2021) <= not a;
    layer8_outputs(2022) <= a;
    layer8_outputs(2023) <= not b;
    layer8_outputs(2024) <= 1'b1;
    layer8_outputs(2025) <= a or b;
    layer8_outputs(2026) <= b and not a;
    layer8_outputs(2027) <= not a;
    layer8_outputs(2028) <= a or b;
    layer8_outputs(2029) <= a and not b;
    layer8_outputs(2030) <= not b or a;
    layer8_outputs(2031) <= not (a xor b);
    layer8_outputs(2032) <= a xor b;
    layer8_outputs(2033) <= a xor b;
    layer8_outputs(2034) <= a;
    layer8_outputs(2035) <= a xor b;
    layer8_outputs(2036) <= not (a xor b);
    layer8_outputs(2037) <= not (a and b);
    layer8_outputs(2038) <= not (a xor b);
    layer8_outputs(2039) <= b;
    layer8_outputs(2040) <= not a;
    layer8_outputs(2041) <= not b;
    layer8_outputs(2042) <= not a;
    layer8_outputs(2043) <= a xor b;
    layer8_outputs(2044) <= b;
    layer8_outputs(2045) <= not b or a;
    layer8_outputs(2046) <= not (a or b);
    layer8_outputs(2047) <= a and b;
    layer8_outputs(2048) <= a xor b;
    layer8_outputs(2049) <= not (a and b);
    layer8_outputs(2050) <= a or b;
    layer8_outputs(2051) <= b;
    layer8_outputs(2052) <= a;
    layer8_outputs(2053) <= not b;
    layer8_outputs(2054) <= b;
    layer8_outputs(2055) <= not a;
    layer8_outputs(2056) <= not a;
    layer8_outputs(2057) <= a and not b;
    layer8_outputs(2058) <= not a;
    layer8_outputs(2059) <= a;
    layer8_outputs(2060) <= not (a xor b);
    layer8_outputs(2061) <= a and not b;
    layer8_outputs(2062) <= not b;
    layer8_outputs(2063) <= b;
    layer8_outputs(2064) <= a xor b;
    layer8_outputs(2065) <= a and b;
    layer8_outputs(2066) <= a and not b;
    layer8_outputs(2067) <= not a or b;
    layer8_outputs(2068) <= not b;
    layer8_outputs(2069) <= not (a xor b);
    layer8_outputs(2070) <= not b or a;
    layer8_outputs(2071) <= a and not b;
    layer8_outputs(2072) <= b and not a;
    layer8_outputs(2073) <= a xor b;
    layer8_outputs(2074) <= not b;
    layer8_outputs(2075) <= 1'b1;
    layer8_outputs(2076) <= a xor b;
    layer8_outputs(2077) <= not (a xor b);
    layer8_outputs(2078) <= a and b;
    layer8_outputs(2079) <= not b or a;
    layer8_outputs(2080) <= not (a and b);
    layer8_outputs(2081) <= 1'b0;
    layer8_outputs(2082) <= a xor b;
    layer8_outputs(2083) <= b;
    layer8_outputs(2084) <= a or b;
    layer8_outputs(2085) <= not b;
    layer8_outputs(2086) <= not a;
    layer8_outputs(2087) <= a;
    layer8_outputs(2088) <= b;
    layer8_outputs(2089) <= a xor b;
    layer8_outputs(2090) <= not (a and b);
    layer8_outputs(2091) <= a or b;
    layer8_outputs(2092) <= not (a or b);
    layer8_outputs(2093) <= a and not b;
    layer8_outputs(2094) <= a and not b;
    layer8_outputs(2095) <= a;
    layer8_outputs(2096) <= a or b;
    layer8_outputs(2097) <= not (a and b);
    layer8_outputs(2098) <= a xor b;
    layer8_outputs(2099) <= b;
    layer8_outputs(2100) <= not a;
    layer8_outputs(2101) <= not b;
    layer8_outputs(2102) <= b and not a;
    layer8_outputs(2103) <= not a;
    layer8_outputs(2104) <= not (a and b);
    layer8_outputs(2105) <= not (a and b);
    layer8_outputs(2106) <= not b;
    layer8_outputs(2107) <= not b or a;
    layer8_outputs(2108) <= a;
    layer8_outputs(2109) <= a or b;
    layer8_outputs(2110) <= not (a and b);
    layer8_outputs(2111) <= not b;
    layer8_outputs(2112) <= a xor b;
    layer8_outputs(2113) <= a and b;
    layer8_outputs(2114) <= b;
    layer8_outputs(2115) <= b;
    layer8_outputs(2116) <= a or b;
    layer8_outputs(2117) <= a xor b;
    layer8_outputs(2118) <= 1'b0;
    layer8_outputs(2119) <= a xor b;
    layer8_outputs(2120) <= not b;
    layer8_outputs(2121) <= b;
    layer8_outputs(2122) <= not (a and b);
    layer8_outputs(2123) <= not b;
    layer8_outputs(2124) <= not b or a;
    layer8_outputs(2125) <= not b;
    layer8_outputs(2126) <= a and not b;
    layer8_outputs(2127) <= not a or b;
    layer8_outputs(2128) <= b;
    layer8_outputs(2129) <= not b;
    layer8_outputs(2130) <= 1'b1;
    layer8_outputs(2131) <= a or b;
    layer8_outputs(2132) <= a xor b;
    layer8_outputs(2133) <= a and not b;
    layer8_outputs(2134) <= 1'b1;
    layer8_outputs(2135) <= a or b;
    layer8_outputs(2136) <= not (a xor b);
    layer8_outputs(2137) <= a;
    layer8_outputs(2138) <= a and not b;
    layer8_outputs(2139) <= not (a xor b);
    layer8_outputs(2140) <= a and b;
    layer8_outputs(2141) <= not (a xor b);
    layer8_outputs(2142) <= a;
    layer8_outputs(2143) <= b;
    layer8_outputs(2144) <= not b;
    layer8_outputs(2145) <= a and not b;
    layer8_outputs(2146) <= a;
    layer8_outputs(2147) <= not (a and b);
    layer8_outputs(2148) <= a and not b;
    layer8_outputs(2149) <= not (a and b);
    layer8_outputs(2150) <= not (a xor b);
    layer8_outputs(2151) <= b;
    layer8_outputs(2152) <= b and not a;
    layer8_outputs(2153) <= b;
    layer8_outputs(2154) <= a and not b;
    layer8_outputs(2155) <= b;
    layer8_outputs(2156) <= a;
    layer8_outputs(2157) <= not b;
    layer8_outputs(2158) <= not (a xor b);
    layer8_outputs(2159) <= not b or a;
    layer8_outputs(2160) <= a xor b;
    layer8_outputs(2161) <= not a or b;
    layer8_outputs(2162) <= not b or a;
    layer8_outputs(2163) <= b and not a;
    layer8_outputs(2164) <= not (a xor b);
    layer8_outputs(2165) <= not (a and b);
    layer8_outputs(2166) <= a;
    layer8_outputs(2167) <= not a;
    layer8_outputs(2168) <= not b;
    layer8_outputs(2169) <= a or b;
    layer8_outputs(2170) <= not b;
    layer8_outputs(2171) <= a xor b;
    layer8_outputs(2172) <= b and not a;
    layer8_outputs(2173) <= not b or a;
    layer8_outputs(2174) <= a and not b;
    layer8_outputs(2175) <= not (a xor b);
    layer8_outputs(2176) <= not b or a;
    layer8_outputs(2177) <= not b;
    layer8_outputs(2178) <= not b;
    layer8_outputs(2179) <= a;
    layer8_outputs(2180) <= a;
    layer8_outputs(2181) <= a;
    layer8_outputs(2182) <= a and b;
    layer8_outputs(2183) <= b;
    layer8_outputs(2184) <= 1'b1;
    layer8_outputs(2185) <= a and b;
    layer8_outputs(2186) <= a;
    layer8_outputs(2187) <= b;
    layer8_outputs(2188) <= not (a and b);
    layer8_outputs(2189) <= a;
    layer8_outputs(2190) <= a;
    layer8_outputs(2191) <= not (a and b);
    layer8_outputs(2192) <= not b;
    layer8_outputs(2193) <= not a;
    layer8_outputs(2194) <= not a;
    layer8_outputs(2195) <= not b;
    layer8_outputs(2196) <= not b;
    layer8_outputs(2197) <= a;
    layer8_outputs(2198) <= not a;
    layer8_outputs(2199) <= b;
    layer8_outputs(2200) <= not (a or b);
    layer8_outputs(2201) <= not a;
    layer8_outputs(2202) <= not (a xor b);
    layer8_outputs(2203) <= a or b;
    layer8_outputs(2204) <= b;
    layer8_outputs(2205) <= not (a xor b);
    layer8_outputs(2206) <= b;
    layer8_outputs(2207) <= a;
    layer8_outputs(2208) <= not b;
    layer8_outputs(2209) <= a and not b;
    layer8_outputs(2210) <= a and not b;
    layer8_outputs(2211) <= not (a or b);
    layer8_outputs(2212) <= not b or a;
    layer8_outputs(2213) <= b;
    layer8_outputs(2214) <= b;
    layer8_outputs(2215) <= a xor b;
    layer8_outputs(2216) <= not b;
    layer8_outputs(2217) <= b;
    layer8_outputs(2218) <= not (a xor b);
    layer8_outputs(2219) <= b and not a;
    layer8_outputs(2220) <= a xor b;
    layer8_outputs(2221) <= not (a or b);
    layer8_outputs(2222) <= not (a and b);
    layer8_outputs(2223) <= a and not b;
    layer8_outputs(2224) <= a;
    layer8_outputs(2225) <= a and b;
    layer8_outputs(2226) <= not (a or b);
    layer8_outputs(2227) <= not a or b;
    layer8_outputs(2228) <= not (a and b);
    layer8_outputs(2229) <= not b or a;
    layer8_outputs(2230) <= a and not b;
    layer8_outputs(2231) <= b and not a;
    layer8_outputs(2232) <= a;
    layer8_outputs(2233) <= a;
    layer8_outputs(2234) <= a;
    layer8_outputs(2235) <= a or b;
    layer8_outputs(2236) <= a;
    layer8_outputs(2237) <= not a or b;
    layer8_outputs(2238) <= a xor b;
    layer8_outputs(2239) <= b and not a;
    layer8_outputs(2240) <= not b;
    layer8_outputs(2241) <= not b;
    layer8_outputs(2242) <= a or b;
    layer8_outputs(2243) <= b;
    layer8_outputs(2244) <= a;
    layer8_outputs(2245) <= a and b;
    layer8_outputs(2246) <= b;
    layer8_outputs(2247) <= not a;
    layer8_outputs(2248) <= not a or b;
    layer8_outputs(2249) <= not b;
    layer8_outputs(2250) <= not a;
    layer8_outputs(2251) <= not b;
    layer8_outputs(2252) <= not b or a;
    layer8_outputs(2253) <= not b;
    layer8_outputs(2254) <= not b or a;
    layer8_outputs(2255) <= not a;
    layer8_outputs(2256) <= b;
    layer8_outputs(2257) <= a or b;
    layer8_outputs(2258) <= not (a xor b);
    layer8_outputs(2259) <= a xor b;
    layer8_outputs(2260) <= not a;
    layer8_outputs(2261) <= b and not a;
    layer8_outputs(2262) <= a xor b;
    layer8_outputs(2263) <= not a;
    layer8_outputs(2264) <= a xor b;
    layer8_outputs(2265) <= a xor b;
    layer8_outputs(2266) <= a;
    layer8_outputs(2267) <= a;
    layer8_outputs(2268) <= a;
    layer8_outputs(2269) <= not b or a;
    layer8_outputs(2270) <= a xor b;
    layer8_outputs(2271) <= b;
    layer8_outputs(2272) <= not b;
    layer8_outputs(2273) <= a and b;
    layer8_outputs(2274) <= not b;
    layer8_outputs(2275) <= not b;
    layer8_outputs(2276) <= not a;
    layer8_outputs(2277) <= a xor b;
    layer8_outputs(2278) <= not a;
    layer8_outputs(2279) <= a;
    layer8_outputs(2280) <= not (a xor b);
    layer8_outputs(2281) <= a xor b;
    layer8_outputs(2282) <= not b;
    layer8_outputs(2283) <= b;
    layer8_outputs(2284) <= a and b;
    layer8_outputs(2285) <= not (a xor b);
    layer8_outputs(2286) <= a and b;
    layer8_outputs(2287) <= a and b;
    layer8_outputs(2288) <= not (a or b);
    layer8_outputs(2289) <= not (a xor b);
    layer8_outputs(2290) <= a xor b;
    layer8_outputs(2291) <= a xor b;
    layer8_outputs(2292) <= b and not a;
    layer8_outputs(2293) <= b;
    layer8_outputs(2294) <= a or b;
    layer8_outputs(2295) <= a xor b;
    layer8_outputs(2296) <= not b;
    layer8_outputs(2297) <= a;
    layer8_outputs(2298) <= not a;
    layer8_outputs(2299) <= b;
    layer8_outputs(2300) <= a xor b;
    layer8_outputs(2301) <= a xor b;
    layer8_outputs(2302) <= b and not a;
    layer8_outputs(2303) <= b;
    layer8_outputs(2304) <= a xor b;
    layer8_outputs(2305) <= not b;
    layer8_outputs(2306) <= b and not a;
    layer8_outputs(2307) <= not a;
    layer8_outputs(2308) <= a;
    layer8_outputs(2309) <= a or b;
    layer8_outputs(2310) <= not a or b;
    layer8_outputs(2311) <= a and not b;
    layer8_outputs(2312) <= a and not b;
    layer8_outputs(2313) <= not (a xor b);
    layer8_outputs(2314) <= a;
    layer8_outputs(2315) <= not (a or b);
    layer8_outputs(2316) <= a;
    layer8_outputs(2317) <= not a or b;
    layer8_outputs(2318) <= not (a or b);
    layer8_outputs(2319) <= a xor b;
    layer8_outputs(2320) <= not (a xor b);
    layer8_outputs(2321) <= a and b;
    layer8_outputs(2322) <= a and b;
    layer8_outputs(2323) <= not (a or b);
    layer8_outputs(2324) <= a xor b;
    layer8_outputs(2325) <= a and not b;
    layer8_outputs(2326) <= not b or a;
    layer8_outputs(2327) <= not (a xor b);
    layer8_outputs(2328) <= a or b;
    layer8_outputs(2329) <= a;
    layer8_outputs(2330) <= a;
    layer8_outputs(2331) <= not (a or b);
    layer8_outputs(2332) <= a xor b;
    layer8_outputs(2333) <= not (a xor b);
    layer8_outputs(2334) <= not b;
    layer8_outputs(2335) <= b;
    layer8_outputs(2336) <= a xor b;
    layer8_outputs(2337) <= not b;
    layer8_outputs(2338) <= b and not a;
    layer8_outputs(2339) <= b;
    layer8_outputs(2340) <= b;
    layer8_outputs(2341) <= a or b;
    layer8_outputs(2342) <= a;
    layer8_outputs(2343) <= a xor b;
    layer8_outputs(2344) <= b;
    layer8_outputs(2345) <= b;
    layer8_outputs(2346) <= not a;
    layer8_outputs(2347) <= a xor b;
    layer8_outputs(2348) <= b and not a;
    layer8_outputs(2349) <= b;
    layer8_outputs(2350) <= not (a and b);
    layer8_outputs(2351) <= not b or a;
    layer8_outputs(2352) <= b and not a;
    layer8_outputs(2353) <= not (a xor b);
    layer8_outputs(2354) <= a and b;
    layer8_outputs(2355) <= a;
    layer8_outputs(2356) <= a and b;
    layer8_outputs(2357) <= not (a and b);
    layer8_outputs(2358) <= a xor b;
    layer8_outputs(2359) <= not b;
    layer8_outputs(2360) <= a;
    layer8_outputs(2361) <= not a or b;
    layer8_outputs(2362) <= a and b;
    layer8_outputs(2363) <= not (a xor b);
    layer8_outputs(2364) <= not a or b;
    layer8_outputs(2365) <= not (a and b);
    layer8_outputs(2366) <= a;
    layer8_outputs(2367) <= not b or a;
    layer8_outputs(2368) <= a;
    layer8_outputs(2369) <= not a;
    layer8_outputs(2370) <= not (a or b);
    layer8_outputs(2371) <= a;
    layer8_outputs(2372) <= not (a xor b);
    layer8_outputs(2373) <= b and not a;
    layer8_outputs(2374) <= b;
    layer8_outputs(2375) <= not b;
    layer8_outputs(2376) <= not a;
    layer8_outputs(2377) <= not b or a;
    layer8_outputs(2378) <= not a;
    layer8_outputs(2379) <= a xor b;
    layer8_outputs(2380) <= a xor b;
    layer8_outputs(2381) <= not (a xor b);
    layer8_outputs(2382) <= a;
    layer8_outputs(2383) <= a and not b;
    layer8_outputs(2384) <= not b;
    layer8_outputs(2385) <= not a;
    layer8_outputs(2386) <= not a or b;
    layer8_outputs(2387) <= not a or b;
    layer8_outputs(2388) <= b and not a;
    layer8_outputs(2389) <= not b;
    layer8_outputs(2390) <= a and b;
    layer8_outputs(2391) <= a xor b;
    layer8_outputs(2392) <= a xor b;
    layer8_outputs(2393) <= a;
    layer8_outputs(2394) <= not (a and b);
    layer8_outputs(2395) <= a;
    layer8_outputs(2396) <= not b;
    layer8_outputs(2397) <= not (a xor b);
    layer8_outputs(2398) <= a;
    layer8_outputs(2399) <= a;
    layer8_outputs(2400) <= not b;
    layer8_outputs(2401) <= not (a and b);
    layer8_outputs(2402) <= not a;
    layer8_outputs(2403) <= not a;
    layer8_outputs(2404) <= not (a and b);
    layer8_outputs(2405) <= not (a and b);
    layer8_outputs(2406) <= not (a xor b);
    layer8_outputs(2407) <= b;
    layer8_outputs(2408) <= a xor b;
    layer8_outputs(2409) <= not b;
    layer8_outputs(2410) <= b;
    layer8_outputs(2411) <= not a or b;
    layer8_outputs(2412) <= a and not b;
    layer8_outputs(2413) <= not (a and b);
    layer8_outputs(2414) <= not (a and b);
    layer8_outputs(2415) <= not b;
    layer8_outputs(2416) <= not (a or b);
    layer8_outputs(2417) <= not b;
    layer8_outputs(2418) <= b;
    layer8_outputs(2419) <= not (a and b);
    layer8_outputs(2420) <= not b;
    layer8_outputs(2421) <= b;
    layer8_outputs(2422) <= not b;
    layer8_outputs(2423) <= b;
    layer8_outputs(2424) <= not (a or b);
    layer8_outputs(2425) <= a xor b;
    layer8_outputs(2426) <= b and not a;
    layer8_outputs(2427) <= not b or a;
    layer8_outputs(2428) <= b and not a;
    layer8_outputs(2429) <= b;
    layer8_outputs(2430) <= not b or a;
    layer8_outputs(2431) <= not b;
    layer8_outputs(2432) <= a or b;
    layer8_outputs(2433) <= not (a or b);
    layer8_outputs(2434) <= not b;
    layer8_outputs(2435) <= not (a or b);
    layer8_outputs(2436) <= not a;
    layer8_outputs(2437) <= a and b;
    layer8_outputs(2438) <= a;
    layer8_outputs(2439) <= not a or b;
    layer8_outputs(2440) <= not (a and b);
    layer8_outputs(2441) <= a xor b;
    layer8_outputs(2442) <= a xor b;
    layer8_outputs(2443) <= not a;
    layer8_outputs(2444) <= a or b;
    layer8_outputs(2445) <= b and not a;
    layer8_outputs(2446) <= not a;
    layer8_outputs(2447) <= b;
    layer8_outputs(2448) <= not a;
    layer8_outputs(2449) <= not a;
    layer8_outputs(2450) <= a;
    layer8_outputs(2451) <= b and not a;
    layer8_outputs(2452) <= not b;
    layer8_outputs(2453) <= not a or b;
    layer8_outputs(2454) <= b and not a;
    layer8_outputs(2455) <= a xor b;
    layer8_outputs(2456) <= b;
    layer8_outputs(2457) <= b and not a;
    layer8_outputs(2458) <= a;
    layer8_outputs(2459) <= not a;
    layer8_outputs(2460) <= not (a and b);
    layer8_outputs(2461) <= not b;
    layer8_outputs(2462) <= a and not b;
    layer8_outputs(2463) <= not (a xor b);
    layer8_outputs(2464) <= b;
    layer8_outputs(2465) <= b;
    layer8_outputs(2466) <= a and not b;
    layer8_outputs(2467) <= a;
    layer8_outputs(2468) <= a;
    layer8_outputs(2469) <= a;
    layer8_outputs(2470) <= a;
    layer8_outputs(2471) <= not (a or b);
    layer8_outputs(2472) <= not b or a;
    layer8_outputs(2473) <= a and not b;
    layer8_outputs(2474) <= b and not a;
    layer8_outputs(2475) <= not b;
    layer8_outputs(2476) <= not (a and b);
    layer8_outputs(2477) <= a and not b;
    layer8_outputs(2478) <= b;
    layer8_outputs(2479) <= a or b;
    layer8_outputs(2480) <= b;
    layer8_outputs(2481) <= a;
    layer8_outputs(2482) <= not a or b;
    layer8_outputs(2483) <= a xor b;
    layer8_outputs(2484) <= not (a xor b);
    layer8_outputs(2485) <= not b;
    layer8_outputs(2486) <= a xor b;
    layer8_outputs(2487) <= not (a or b);
    layer8_outputs(2488) <= a or b;
    layer8_outputs(2489) <= not b or a;
    layer8_outputs(2490) <= not (a or b);
    layer8_outputs(2491) <= b;
    layer8_outputs(2492) <= b and not a;
    layer8_outputs(2493) <= a xor b;
    layer8_outputs(2494) <= a xor b;
    layer8_outputs(2495) <= not a;
    layer8_outputs(2496) <= b and not a;
    layer8_outputs(2497) <= not (a xor b);
    layer8_outputs(2498) <= b and not a;
    layer8_outputs(2499) <= not a;
    layer8_outputs(2500) <= not a or b;
    layer8_outputs(2501) <= b;
    layer8_outputs(2502) <= not (a xor b);
    layer8_outputs(2503) <= a and not b;
    layer8_outputs(2504) <= a and b;
    layer8_outputs(2505) <= a and b;
    layer8_outputs(2506) <= not b;
    layer8_outputs(2507) <= not b or a;
    layer8_outputs(2508) <= b;
    layer8_outputs(2509) <= a and not b;
    layer8_outputs(2510) <= a;
    layer8_outputs(2511) <= not a;
    layer8_outputs(2512) <= not b or a;
    layer8_outputs(2513) <= not (a and b);
    layer8_outputs(2514) <= a;
    layer8_outputs(2515) <= not (a or b);
    layer8_outputs(2516) <= not a;
    layer8_outputs(2517) <= not b;
    layer8_outputs(2518) <= not a or b;
    layer8_outputs(2519) <= not (a xor b);
    layer8_outputs(2520) <= a and b;
    layer8_outputs(2521) <= not a;
    layer8_outputs(2522) <= b;
    layer8_outputs(2523) <= not b or a;
    layer8_outputs(2524) <= b;
    layer8_outputs(2525) <= not a;
    layer8_outputs(2526) <= not b;
    layer8_outputs(2527) <= a xor b;
    layer8_outputs(2528) <= not (a xor b);
    layer8_outputs(2529) <= not (a xor b);
    layer8_outputs(2530) <= b;
    layer8_outputs(2531) <= a;
    layer8_outputs(2532) <= not (a xor b);
    layer8_outputs(2533) <= not (a xor b);
    layer8_outputs(2534) <= b and not a;
    layer8_outputs(2535) <= not a;
    layer8_outputs(2536) <= a;
    layer8_outputs(2537) <= not b;
    layer8_outputs(2538) <= not a or b;
    layer8_outputs(2539) <= not a;
    layer8_outputs(2540) <= a and b;
    layer8_outputs(2541) <= b and not a;
    layer8_outputs(2542) <= a and not b;
    layer8_outputs(2543) <= not b;
    layer8_outputs(2544) <= a and b;
    layer8_outputs(2545) <= a xor b;
    layer8_outputs(2546) <= a or b;
    layer8_outputs(2547) <= not b;
    layer8_outputs(2548) <= a xor b;
    layer8_outputs(2549) <= not (a xor b);
    layer8_outputs(2550) <= not (a and b);
    layer8_outputs(2551) <= not a or b;
    layer8_outputs(2552) <= a xor b;
    layer8_outputs(2553) <= not (a xor b);
    layer8_outputs(2554) <= not a;
    layer8_outputs(2555) <= b;
    layer8_outputs(2556) <= b and not a;
    layer8_outputs(2557) <= not a;
    layer8_outputs(2558) <= a;
    layer8_outputs(2559) <= not b;
    outputs(0) <= a and b;
    outputs(1) <= not (a or b);
    outputs(2) <= a and not b;
    outputs(3) <= a;
    outputs(4) <= not (a xor b);
    outputs(5) <= a;
    outputs(6) <= not (a xor b);
    outputs(7) <= not (a or b);
    outputs(8) <= not b;
    outputs(9) <= not (a or b);
    outputs(10) <= a xor b;
    outputs(11) <= not b;
    outputs(12) <= a and not b;
    outputs(13) <= b;
    outputs(14) <= not a or b;
    outputs(15) <= b;
    outputs(16) <= a;
    outputs(17) <= a;
    outputs(18) <= a and not b;
    outputs(19) <= not (a or b);
    outputs(20) <= a and not b;
    outputs(21) <= a and not b;
    outputs(22) <= a;
    outputs(23) <= a and b;
    outputs(24) <= not a;
    outputs(25) <= a and b;
    outputs(26) <= not b or a;
    outputs(27) <= a and not b;
    outputs(28) <= b;
    outputs(29) <= not b;
    outputs(30) <= not (a xor b);
    outputs(31) <= not (a xor b);
    outputs(32) <= not (a and b);
    outputs(33) <= not b;
    outputs(34) <= a;
    outputs(35) <= a xor b;
    outputs(36) <= a and b;
    outputs(37) <= not (a or b);
    outputs(38) <= a or b;
    outputs(39) <= a;
    outputs(40) <= not (a or b);
    outputs(41) <= a;
    outputs(42) <= not (a xor b);
    outputs(43) <= not (a xor b);
    outputs(44) <= not (a xor b);
    outputs(45) <= not b;
    outputs(46) <= a and b;
    outputs(47) <= a and not b;
    outputs(48) <= a;
    outputs(49) <= a;
    outputs(50) <= b and not a;
    outputs(51) <= a;
    outputs(52) <= not a;
    outputs(53) <= a;
    outputs(54) <= not a;
    outputs(55) <= not a or b;
    outputs(56) <= a xor b;
    outputs(57) <= a;
    outputs(58) <= not (a or b);
    outputs(59) <= a and not b;
    outputs(60) <= not a;
    outputs(61) <= not (a or b);
    outputs(62) <= a;
    outputs(63) <= b;
    outputs(64) <= not a;
    outputs(65) <= b and not a;
    outputs(66) <= not a;
    outputs(67) <= not a;
    outputs(68) <= b and not a;
    outputs(69) <= a;
    outputs(70) <= not a;
    outputs(71) <= a or b;
    outputs(72) <= not (a or b);
    outputs(73) <= a and b;
    outputs(74) <= a and not b;
    outputs(75) <= a;
    outputs(76) <= a xor b;
    outputs(77) <= b and not a;
    outputs(78) <= a xor b;
    outputs(79) <= a xor b;
    outputs(80) <= not b or a;
    outputs(81) <= not (a or b);
    outputs(82) <= a xor b;
    outputs(83) <= a xor b;
    outputs(84) <= not b;
    outputs(85) <= a;
    outputs(86) <= a;
    outputs(87) <= a and b;
    outputs(88) <= not b;
    outputs(89) <= a xor b;
    outputs(90) <= not b;
    outputs(91) <= not a or b;
    outputs(92) <= not b;
    outputs(93) <= b;
    outputs(94) <= not a or b;
    outputs(95) <= not b;
    outputs(96) <= a;
    outputs(97) <= a xor b;
    outputs(98) <= a;
    outputs(99) <= not (a xor b);
    outputs(100) <= not b;
    outputs(101) <= a;
    outputs(102) <= not a;
    outputs(103) <= not b;
    outputs(104) <= b and not a;
    outputs(105) <= b;
    outputs(106) <= not b;
    outputs(107) <= a and not b;
    outputs(108) <= a;
    outputs(109) <= a;
    outputs(110) <= not (a xor b);
    outputs(111) <= a;
    outputs(112) <= not a;
    outputs(113) <= not a;
    outputs(114) <= a and not b;
    outputs(115) <= not a or b;
    outputs(116) <= not b;
    outputs(117) <= a and not b;
    outputs(118) <= b;
    outputs(119) <= a xor b;
    outputs(120) <= b;
    outputs(121) <= not b;
    outputs(122) <= not b;
    outputs(123) <= b;
    outputs(124) <= not (a xor b);
    outputs(125) <= not b;
    outputs(126) <= a xor b;
    outputs(127) <= a and b;
    outputs(128) <= b;
    outputs(129) <= a;
    outputs(130) <= not (a and b);
    outputs(131) <= a and b;
    outputs(132) <= not b;
    outputs(133) <= not b;
    outputs(134) <= not b;
    outputs(135) <= a and not b;
    outputs(136) <= not (a and b);
    outputs(137) <= a xor b;
    outputs(138) <= b and not a;
    outputs(139) <= not a;
    outputs(140) <= b and not a;
    outputs(141) <= a xor b;
    outputs(142) <= not a;
    outputs(143) <= not b;
    outputs(144) <= a;
    outputs(145) <= not a;
    outputs(146) <= not (a xor b);
    outputs(147) <= not b;
    outputs(148) <= a or b;
    outputs(149) <= not (a xor b);
    outputs(150) <= a xor b;
    outputs(151) <= not a;
    outputs(152) <= not b;
    outputs(153) <= not a;
    outputs(154) <= not (a or b);
    outputs(155) <= a xor b;
    outputs(156) <= a xor b;
    outputs(157) <= not (a xor b);
    outputs(158) <= not b;
    outputs(159) <= not a;
    outputs(160) <= not a or b;
    outputs(161) <= not a;
    outputs(162) <= not (a or b);
    outputs(163) <= b and not a;
    outputs(164) <= not (a or b);
    outputs(165) <= b;
    outputs(166) <= not (a or b);
    outputs(167) <= a xor b;
    outputs(168) <= not a;
    outputs(169) <= a xor b;
    outputs(170) <= not (a xor b);
    outputs(171) <= not a;
    outputs(172) <= a xor b;
    outputs(173) <= not a;
    outputs(174) <= b and not a;
    outputs(175) <= b and not a;
    outputs(176) <= b;
    outputs(177) <= b and not a;
    outputs(178) <= b and not a;
    outputs(179) <= a;
    outputs(180) <= not b;
    outputs(181) <= a xor b;
    outputs(182) <= a xor b;
    outputs(183) <= not b;
    outputs(184) <= b and not a;
    outputs(185) <= not (a and b);
    outputs(186) <= a xor b;
    outputs(187) <= a and b;
    outputs(188) <= a xor b;
    outputs(189) <= not (a or b);
    outputs(190) <= b;
    outputs(191) <= a xor b;
    outputs(192) <= not (a xor b);
    outputs(193) <= a and not b;
    outputs(194) <= not (a xor b);
    outputs(195) <= a and b;
    outputs(196) <= a;
    outputs(197) <= not b;
    outputs(198) <= b;
    outputs(199) <= not a;
    outputs(200) <= a xor b;
    outputs(201) <= a or b;
    outputs(202) <= a;
    outputs(203) <= a xor b;
    outputs(204) <= not a;
    outputs(205) <= a;
    outputs(206) <= a;
    outputs(207) <= b and not a;
    outputs(208) <= a and not b;
    outputs(209) <= not a;
    outputs(210) <= a and not b;
    outputs(211) <= a;
    outputs(212) <= not (a or b);
    outputs(213) <= b;
    outputs(214) <= a and b;
    outputs(215) <= not (a or b);
    outputs(216) <= b;
    outputs(217) <= not a;
    outputs(218) <= not (a xor b);
    outputs(219) <= not a;
    outputs(220) <= not (a and b);
    outputs(221) <= a;
    outputs(222) <= not (a xor b);
    outputs(223) <= a and b;
    outputs(224) <= not a;
    outputs(225) <= a and not b;
    outputs(226) <= not b or a;
    outputs(227) <= a xor b;
    outputs(228) <= a and b;
    outputs(229) <= not a;
    outputs(230) <= not b;
    outputs(231) <= not b;
    outputs(232) <= not (a xor b);
    outputs(233) <= b;
    outputs(234) <= b;
    outputs(235) <= a and not b;
    outputs(236) <= not a or b;
    outputs(237) <= b;
    outputs(238) <= not (a xor b);
    outputs(239) <= a;
    outputs(240) <= a and not b;
    outputs(241) <= a;
    outputs(242) <= not a;
    outputs(243) <= b;
    outputs(244) <= a;
    outputs(245) <= not b;
    outputs(246) <= not (a xor b);
    outputs(247) <= not (a or b);
    outputs(248) <= not a;
    outputs(249) <= a;
    outputs(250) <= a;
    outputs(251) <= a and not b;
    outputs(252) <= a and b;
    outputs(253) <= not b;
    outputs(254) <= b;
    outputs(255) <= not b;
    outputs(256) <= a and not b;
    outputs(257) <= not a;
    outputs(258) <= not (a xor b);
    outputs(259) <= a and b;
    outputs(260) <= b and not a;
    outputs(261) <= a xor b;
    outputs(262) <= not b;
    outputs(263) <= a;
    outputs(264) <= b and not a;
    outputs(265) <= b;
    outputs(266) <= b;
    outputs(267) <= not a;
    outputs(268) <= not a;
    outputs(269) <= a and not b;
    outputs(270) <= not b;
    outputs(271) <= b and not a;
    outputs(272) <= a and b;
    outputs(273) <= a and b;
    outputs(274) <= a and b;
    outputs(275) <= a and b;
    outputs(276) <= a;
    outputs(277) <= not a;
    outputs(278) <= not a or b;
    outputs(279) <= a xor b;
    outputs(280) <= not (a or b);
    outputs(281) <= b;
    outputs(282) <= b and not a;
    outputs(283) <= a and not b;
    outputs(284) <= not a;
    outputs(285) <= not a;
    outputs(286) <= not (a or b);
    outputs(287) <= not (a or b);
    outputs(288) <= a xor b;
    outputs(289) <= not a;
    outputs(290) <= b and not a;
    outputs(291) <= not a;
    outputs(292) <= a xor b;
    outputs(293) <= a and not b;
    outputs(294) <= b;
    outputs(295) <= a;
    outputs(296) <= not a;
    outputs(297) <= a;
    outputs(298) <= a xor b;
    outputs(299) <= not (a xor b);
    outputs(300) <= not b;
    outputs(301) <= a and not b;
    outputs(302) <= b;
    outputs(303) <= not a;
    outputs(304) <= a and not b;
    outputs(305) <= a xor b;
    outputs(306) <= a and b;
    outputs(307) <= a;
    outputs(308) <= a xor b;
    outputs(309) <= b and not a;
    outputs(310) <= not a;
    outputs(311) <= not (a or b);
    outputs(312) <= not (a or b);
    outputs(313) <= b;
    outputs(314) <= a;
    outputs(315) <= a;
    outputs(316) <= a and not b;
    outputs(317) <= a xor b;
    outputs(318) <= not b;
    outputs(319) <= a and not b;
    outputs(320) <= a and b;
    outputs(321) <= not (a and b);
    outputs(322) <= not a;
    outputs(323) <= b and not a;
    outputs(324) <= b;
    outputs(325) <= a and b;
    outputs(326) <= a;
    outputs(327) <= b;
    outputs(328) <= b and not a;
    outputs(329) <= a;
    outputs(330) <= b and not a;
    outputs(331) <= a and not b;
    outputs(332) <= a;
    outputs(333) <= not (a or b);
    outputs(334) <= a and not b;
    outputs(335) <= a xor b;
    outputs(336) <= not a;
    outputs(337) <= not (a xor b);
    outputs(338) <= a;
    outputs(339) <= not (a or b);
    outputs(340) <= not a;
    outputs(341) <= not (a or b);
    outputs(342) <= b and not a;
    outputs(343) <= not (a or b);
    outputs(344) <= a xor b;
    outputs(345) <= a;
    outputs(346) <= a;
    outputs(347) <= b and not a;
    outputs(348) <= a and b;
    outputs(349) <= a and not b;
    outputs(350) <= b and not a;
    outputs(351) <= a or b;
    outputs(352) <= b;
    outputs(353) <= a;
    outputs(354) <= a and b;
    outputs(355) <= a and not b;
    outputs(356) <= not b;
    outputs(357) <= a or b;
    outputs(358) <= not a or b;
    outputs(359) <= a and not b;
    outputs(360) <= a and not b;
    outputs(361) <= a xor b;
    outputs(362) <= b;
    outputs(363) <= a;
    outputs(364) <= not (a xor b);
    outputs(365) <= not (a or b);
    outputs(366) <= a and not b;
    outputs(367) <= a;
    outputs(368) <= a and b;
    outputs(369) <= b;
    outputs(370) <= a xor b;
    outputs(371) <= not b;
    outputs(372) <= not (a xor b);
    outputs(373) <= b;
    outputs(374) <= not (a xor b);
    outputs(375) <= not (a or b);
    outputs(376) <= a and not b;
    outputs(377) <= not (a or b);
    outputs(378) <= a and not b;
    outputs(379) <= a and not b;
    outputs(380) <= not b;
    outputs(381) <= a;
    outputs(382) <= a xor b;
    outputs(383) <= not (a or b);
    outputs(384) <= b;
    outputs(385) <= b and not a;
    outputs(386) <= not (a xor b);
    outputs(387) <= a;
    outputs(388) <= a;
    outputs(389) <= not b;
    outputs(390) <= a or b;
    outputs(391) <= not a;
    outputs(392) <= not a;
    outputs(393) <= not a;
    outputs(394) <= not (a xor b);
    outputs(395) <= a and not b;
    outputs(396) <= b and not a;
    outputs(397) <= a and b;
    outputs(398) <= a;
    outputs(399) <= a and b;
    outputs(400) <= not a;
    outputs(401) <= b and not a;
    outputs(402) <= not (a or b);
    outputs(403) <= not a;
    outputs(404) <= b;
    outputs(405) <= not (a or b);
    outputs(406) <= b and not a;
    outputs(407) <= b and not a;
    outputs(408) <= b;
    outputs(409) <= not a;
    outputs(410) <= not (a or b);
    outputs(411) <= not b;
    outputs(412) <= b and not a;
    outputs(413) <= not a;
    outputs(414) <= not b;
    outputs(415) <= a xor b;
    outputs(416) <= not a;
    outputs(417) <= a;
    outputs(418) <= a and not b;
    outputs(419) <= not b;
    outputs(420) <= a and b;
    outputs(421) <= a;
    outputs(422) <= not (a xor b);
    outputs(423) <= a and not b;
    outputs(424) <= a xor b;
    outputs(425) <= a and not b;
    outputs(426) <= a and not b;
    outputs(427) <= not b;
    outputs(428) <= a;
    outputs(429) <= a and b;
    outputs(430) <= b;
    outputs(431) <= a and not b;
    outputs(432) <= b;
    outputs(433) <= a xor b;
    outputs(434) <= not (a or b);
    outputs(435) <= b;
    outputs(436) <= a xor b;
    outputs(437) <= b and not a;
    outputs(438) <= a xor b;
    outputs(439) <= not b;
    outputs(440) <= not (a xor b);
    outputs(441) <= b and not a;
    outputs(442) <= not a;
    outputs(443) <= not a or b;
    outputs(444) <= not (a xor b);
    outputs(445) <= b;
    outputs(446) <= a xor b;
    outputs(447) <= b and not a;
    outputs(448) <= a;
    outputs(449) <= a and b;
    outputs(450) <= a and b;
    outputs(451) <= a and not b;
    outputs(452) <= a;
    outputs(453) <= not a;
    outputs(454) <= a and b;
    outputs(455) <= b and not a;
    outputs(456) <= a xor b;
    outputs(457) <= a xor b;
    outputs(458) <= not b;
    outputs(459) <= not a;
    outputs(460) <= not (a or b);
    outputs(461) <= b;
    outputs(462) <= not (a or b);
    outputs(463) <= b and not a;
    outputs(464) <= a;
    outputs(465) <= not a;
    outputs(466) <= b;
    outputs(467) <= a and b;
    outputs(468) <= a;
    outputs(469) <= a;
    outputs(470) <= not (a or b);
    outputs(471) <= a and b;
    outputs(472) <= a xor b;
    outputs(473) <= a and not b;
    outputs(474) <= a xor b;
    outputs(475) <= a xor b;
    outputs(476) <= not b;
    outputs(477) <= not b;
    outputs(478) <= a and b;
    outputs(479) <= a xor b;
    outputs(480) <= a and not b;
    outputs(481) <= a and b;
    outputs(482) <= not (a xor b);
    outputs(483) <= a xor b;
    outputs(484) <= a;
    outputs(485) <= not (a or b);
    outputs(486) <= a xor b;
    outputs(487) <= not (a or b);
    outputs(488) <= a and not b;
    outputs(489) <= a xor b;
    outputs(490) <= not (a or b);
    outputs(491) <= not b;
    outputs(492) <= b;
    outputs(493) <= not (a or b);
    outputs(494) <= a and b;
    outputs(495) <= not a;
    outputs(496) <= not (a or b);
    outputs(497) <= a and b;
    outputs(498) <= a xor b;
    outputs(499) <= b;
    outputs(500) <= not a;
    outputs(501) <= a and not b;
    outputs(502) <= not b;
    outputs(503) <= a;
    outputs(504) <= not (a xor b);
    outputs(505) <= a and b;
    outputs(506) <= b and not a;
    outputs(507) <= b and not a;
    outputs(508) <= a and b;
    outputs(509) <= b and not a;
    outputs(510) <= not (a or b);
    outputs(511) <= a and not b;
    outputs(512) <= a xor b;
    outputs(513) <= not b;
    outputs(514) <= not (a xor b);
    outputs(515) <= a;
    outputs(516) <= a xor b;
    outputs(517) <= a;
    outputs(518) <= a xor b;
    outputs(519) <= a;
    outputs(520) <= a;
    outputs(521) <= not b;
    outputs(522) <= b;
    outputs(523) <= a and b;
    outputs(524) <= b;
    outputs(525) <= a;
    outputs(526) <= not b or a;
    outputs(527) <= not a;
    outputs(528) <= not (a xor b);
    outputs(529) <= not b;
    outputs(530) <= b;
    outputs(531) <= not (a xor b);
    outputs(532) <= b;
    outputs(533) <= not (a or b);
    outputs(534) <= not b or a;
    outputs(535) <= b;
    outputs(536) <= a;
    outputs(537) <= b;
    outputs(538) <= not b;
    outputs(539) <= b and not a;
    outputs(540) <= not b;
    outputs(541) <= not (a xor b);
    outputs(542) <= not (a xor b);
    outputs(543) <= not (a or b);
    outputs(544) <= b;
    outputs(545) <= a xor b;
    outputs(546) <= not b;
    outputs(547) <= a or b;
    outputs(548) <= a and b;
    outputs(549) <= a xor b;
    outputs(550) <= a xor b;
    outputs(551) <= a;
    outputs(552) <= not (a xor b);
    outputs(553) <= not (a xor b);
    outputs(554) <= b;
    outputs(555) <= not a;
    outputs(556) <= a xor b;
    outputs(557) <= a;
    outputs(558) <= a;
    outputs(559) <= b and not a;
    outputs(560) <= a and not b;
    outputs(561) <= not a;
    outputs(562) <= a or b;
    outputs(563) <= b;
    outputs(564) <= not a;
    outputs(565) <= a xor b;
    outputs(566) <= not (a xor b);
    outputs(567) <= a and not b;
    outputs(568) <= not b or a;
    outputs(569) <= not (a xor b);
    outputs(570) <= not a;
    outputs(571) <= not b;
    outputs(572) <= b and not a;
    outputs(573) <= a and not b;
    outputs(574) <= a;
    outputs(575) <= a xor b;
    outputs(576) <= a and not b;
    outputs(577) <= b and not a;
    outputs(578) <= b;
    outputs(579) <= b and not a;
    outputs(580) <= b;
    outputs(581) <= a;
    outputs(582) <= not (a or b);
    outputs(583) <= not (a xor b);
    outputs(584) <= not (a or b);
    outputs(585) <= not (a xor b);
    outputs(586) <= b;
    outputs(587) <= a;
    outputs(588) <= b;
    outputs(589) <= not a or b;
    outputs(590) <= not a;
    outputs(591) <= not (a or b);
    outputs(592) <= b and not a;
    outputs(593) <= not (a and b);
    outputs(594) <= not a;
    outputs(595) <= not (a or b);
    outputs(596) <= not b;
    outputs(597) <= a;
    outputs(598) <= not a or b;
    outputs(599) <= a;
    outputs(600) <= a;
    outputs(601) <= not b;
    outputs(602) <= a or b;
    outputs(603) <= not a;
    outputs(604) <= not a;
    outputs(605) <= a;
    outputs(606) <= not (a xor b);
    outputs(607) <= a and b;
    outputs(608) <= a xor b;
    outputs(609) <= not a;
    outputs(610) <= not b or a;
    outputs(611) <= not b or a;
    outputs(612) <= a and b;
    outputs(613) <= a;
    outputs(614) <= a xor b;
    outputs(615) <= a or b;
    outputs(616) <= not b or a;
    outputs(617) <= not b;
    outputs(618) <= b and not a;
    outputs(619) <= b;
    outputs(620) <= b;
    outputs(621) <= not b;
    outputs(622) <= not a or b;
    outputs(623) <= a and not b;
    outputs(624) <= b;
    outputs(625) <= not (a and b);
    outputs(626) <= b;
    outputs(627) <= not (a xor b);
    outputs(628) <= not a;
    outputs(629) <= not b;
    outputs(630) <= not b or a;
    outputs(631) <= not a;
    outputs(632) <= b and not a;
    outputs(633) <= not a;
    outputs(634) <= not a;
    outputs(635) <= a and b;
    outputs(636) <= b;
    outputs(637) <= a;
    outputs(638) <= b;
    outputs(639) <= b and not a;
    outputs(640) <= not b or a;
    outputs(641) <= b;
    outputs(642) <= a and b;
    outputs(643) <= a xor b;
    outputs(644) <= not (a xor b);
    outputs(645) <= a or b;
    outputs(646) <= not (a xor b);
    outputs(647) <= b;
    outputs(648) <= not a;
    outputs(649) <= not (a or b);
    outputs(650) <= b;
    outputs(651) <= not b;
    outputs(652) <= not (a xor b);
    outputs(653) <= a and b;
    outputs(654) <= a and b;
    outputs(655) <= not a;
    outputs(656) <= not a or b;
    outputs(657) <= a xor b;
    outputs(658) <= a xor b;
    outputs(659) <= not (a xor b);
    outputs(660) <= b;
    outputs(661) <= a xor b;
    outputs(662) <= not a or b;
    outputs(663) <= a;
    outputs(664) <= not a;
    outputs(665) <= not (a or b);
    outputs(666) <= not a or b;
    outputs(667) <= a and not b;
    outputs(668) <= not a;
    outputs(669) <= b and not a;
    outputs(670) <= b;
    outputs(671) <= b;
    outputs(672) <= not a;
    outputs(673) <= not a;
    outputs(674) <= a;
    outputs(675) <= not (a or b);
    outputs(676) <= not b;
    outputs(677) <= a and b;
    outputs(678) <= not b;
    outputs(679) <= not b;
    outputs(680) <= not (a and b);
    outputs(681) <= not (a xor b);
    outputs(682) <= not (a or b);
    outputs(683) <= not a or b;
    outputs(684) <= not b or a;
    outputs(685) <= a;
    outputs(686) <= b;
    outputs(687) <= b and not a;
    outputs(688) <= not b or a;
    outputs(689) <= not (a or b);
    outputs(690) <= not b;
    outputs(691) <= not b;
    outputs(692) <= a;
    outputs(693) <= not b;
    outputs(694) <= a;
    outputs(695) <= not a;
    outputs(696) <= a and b;
    outputs(697) <= a;
    outputs(698) <= a;
    outputs(699) <= b;
    outputs(700) <= a;
    outputs(701) <= not (a xor b);
    outputs(702) <= a and b;
    outputs(703) <= b and not a;
    outputs(704) <= a;
    outputs(705) <= a and b;
    outputs(706) <= a or b;
    outputs(707) <= not (a xor b);
    outputs(708) <= a and not b;
    outputs(709) <= not (a or b);
    outputs(710) <= a;
    outputs(711) <= a;
    outputs(712) <= not b;
    outputs(713) <= not a;
    outputs(714) <= a and b;
    outputs(715) <= not b;
    outputs(716) <= b and not a;
    outputs(717) <= a and b;
    outputs(718) <= a xor b;
    outputs(719) <= not b;
    outputs(720) <= b;
    outputs(721) <= b;
    outputs(722) <= b;
    outputs(723) <= not a;
    outputs(724) <= not b;
    outputs(725) <= a or b;
    outputs(726) <= not (a or b);
    outputs(727) <= b;
    outputs(728) <= not (a xor b);
    outputs(729) <= not (a and b);
    outputs(730) <= b;
    outputs(731) <= not a;
    outputs(732) <= not b;
    outputs(733) <= not (a xor b);
    outputs(734) <= not b;
    outputs(735) <= not b;
    outputs(736) <= not (a or b);
    outputs(737) <= not (a and b);
    outputs(738) <= a;
    outputs(739) <= a;
    outputs(740) <= a and not b;
    outputs(741) <= not a or b;
    outputs(742) <= b;
    outputs(743) <= b and not a;
    outputs(744) <= not a or b;
    outputs(745) <= b and not a;
    outputs(746) <= a xor b;
    outputs(747) <= not (a xor b);
    outputs(748) <= b;
    outputs(749) <= a xor b;
    outputs(750) <= not a;
    outputs(751) <= a;
    outputs(752) <= not (a or b);
    outputs(753) <= not b;
    outputs(754) <= not a or b;
    outputs(755) <= a and not b;
    outputs(756) <= a;
    outputs(757) <= not a;
    outputs(758) <= b;
    outputs(759) <= b;
    outputs(760) <= not b;
    outputs(761) <= not a or b;
    outputs(762) <= not (a or b);
    outputs(763) <= a and b;
    outputs(764) <= a and not b;
    outputs(765) <= not b or a;
    outputs(766) <= b and not a;
    outputs(767) <= not a;
    outputs(768) <= not b or a;
    outputs(769) <= not a;
    outputs(770) <= not (a or b);
    outputs(771) <= not a or b;
    outputs(772) <= not (a xor b);
    outputs(773) <= not b;
    outputs(774) <= a xor b;
    outputs(775) <= not a;
    outputs(776) <= not b;
    outputs(777) <= b and not a;
    outputs(778) <= a and b;
    outputs(779) <= not a;
    outputs(780) <= b;
    outputs(781) <= not a;
    outputs(782) <= not (a or b);
    outputs(783) <= not a;
    outputs(784) <= a and not b;
    outputs(785) <= a;
    outputs(786) <= not b;
    outputs(787) <= a;
    outputs(788) <= b;
    outputs(789) <= not a or b;
    outputs(790) <= a and b;
    outputs(791) <= a;
    outputs(792) <= not (a or b);
    outputs(793) <= not (a and b);
    outputs(794) <= not (a and b);
    outputs(795) <= not b;
    outputs(796) <= a and not b;
    outputs(797) <= a or b;
    outputs(798) <= a and b;
    outputs(799) <= b and not a;
    outputs(800) <= not (a or b);
    outputs(801) <= not (a xor b);
    outputs(802) <= b;
    outputs(803) <= not a;
    outputs(804) <= a and b;
    outputs(805) <= a and b;
    outputs(806) <= not (a or b);
    outputs(807) <= b and not a;
    outputs(808) <= b;
    outputs(809) <= not (a xor b);
    outputs(810) <= not b;
    outputs(811) <= not b;
    outputs(812) <= not (a xor b);
    outputs(813) <= not b;
    outputs(814) <= not a or b;
    outputs(815) <= a and not b;
    outputs(816) <= not b;
    outputs(817) <= a xor b;
    outputs(818) <= b;
    outputs(819) <= not b;
    outputs(820) <= not a or b;
    outputs(821) <= a;
    outputs(822) <= not a or b;
    outputs(823) <= a and not b;
    outputs(824) <= b;
    outputs(825) <= a and not b;
    outputs(826) <= not a;
    outputs(827) <= b;
    outputs(828) <= not a;
    outputs(829) <= a;
    outputs(830) <= not (a xor b);
    outputs(831) <= a xor b;
    outputs(832) <= a and not b;
    outputs(833) <= a xor b;
    outputs(834) <= not a;
    outputs(835) <= not b;
    outputs(836) <= not (a xor b);
    outputs(837) <= a xor b;
    outputs(838) <= not (a or b);
    outputs(839) <= b;
    outputs(840) <= not (a or b);
    outputs(841) <= a and b;
    outputs(842) <= not a;
    outputs(843) <= a;
    outputs(844) <= not b;
    outputs(845) <= not (a xor b);
    outputs(846) <= b;
    outputs(847) <= a and not b;
    outputs(848) <= not a;
    outputs(849) <= not (a or b);
    outputs(850) <= a and b;
    outputs(851) <= not b;
    outputs(852) <= a xor b;
    outputs(853) <= b;
    outputs(854) <= not (a xor b);
    outputs(855) <= a and b;
    outputs(856) <= a xor b;
    outputs(857) <= b;
    outputs(858) <= not (a xor b);
    outputs(859) <= b and not a;
    outputs(860) <= not (a or b);
    outputs(861) <= a and b;
    outputs(862) <= b;
    outputs(863) <= a or b;
    outputs(864) <= a;
    outputs(865) <= not a;
    outputs(866) <= not (a or b);
    outputs(867) <= not (a or b);
    outputs(868) <= a xor b;
    outputs(869) <= not a;
    outputs(870) <= a and b;
    outputs(871) <= not (a xor b);
    outputs(872) <= b and not a;
    outputs(873) <= not b;
    outputs(874) <= a;
    outputs(875) <= not a;
    outputs(876) <= not a;
    outputs(877) <= a xor b;
    outputs(878) <= a or b;
    outputs(879) <= a and b;
    outputs(880) <= a;
    outputs(881) <= b and not a;
    outputs(882) <= not (a or b);
    outputs(883) <= not (a and b);
    outputs(884) <= not (a or b);
    outputs(885) <= not (a or b);
    outputs(886) <= not a;
    outputs(887) <= b and not a;
    outputs(888) <= not (a xor b);
    outputs(889) <= a and b;
    outputs(890) <= b and not a;
    outputs(891) <= a and not b;
    outputs(892) <= not a or b;
    outputs(893) <= not a or b;
    outputs(894) <= a and b;
    outputs(895) <= not a;
    outputs(896) <= not b;
    outputs(897) <= b;
    outputs(898) <= not (a xor b);
    outputs(899) <= a xor b;
    outputs(900) <= not (a and b);
    outputs(901) <= not (a or b);
    outputs(902) <= a and not b;
    outputs(903) <= not (a or b);
    outputs(904) <= not b;
    outputs(905) <= a xor b;
    outputs(906) <= not (a or b);
    outputs(907) <= a xor b;
    outputs(908) <= a and b;
    outputs(909) <= not (a or b);
    outputs(910) <= not b;
    outputs(911) <= not a;
    outputs(912) <= a and not b;
    outputs(913) <= b;
    outputs(914) <= not a;
    outputs(915) <= a xor b;
    outputs(916) <= not (a xor b);
    outputs(917) <= not a;
    outputs(918) <= a and b;
    outputs(919) <= a xor b;
    outputs(920) <= not (a or b);
    outputs(921) <= not a or b;
    outputs(922) <= b;
    outputs(923) <= not (a or b);
    outputs(924) <= not a;
    outputs(925) <= a or b;
    outputs(926) <= not a;
    outputs(927) <= not a;
    outputs(928) <= not a;
    outputs(929) <= b;
    outputs(930) <= a and b;
    outputs(931) <= b;
    outputs(932) <= not (a and b);
    outputs(933) <= not (a xor b);
    outputs(934) <= not (a xor b);
    outputs(935) <= a xor b;
    outputs(936) <= a xor b;
    outputs(937) <= b;
    outputs(938) <= a;
    outputs(939) <= not b;
    outputs(940) <= b and not a;
    outputs(941) <= not a;
    outputs(942) <= a and not b;
    outputs(943) <= a;
    outputs(944) <= a;
    outputs(945) <= not b;
    outputs(946) <= a and b;
    outputs(947) <= a and b;
    outputs(948) <= a xor b;
    outputs(949) <= a;
    outputs(950) <= not (a or b);
    outputs(951) <= b;
    outputs(952) <= a and b;
    outputs(953) <= not (a xor b);
    outputs(954) <= a or b;
    outputs(955) <= not b;
    outputs(956) <= not (a or b);
    outputs(957) <= not b or a;
    outputs(958) <= b;
    outputs(959) <= not (a xor b);
    outputs(960) <= a;
    outputs(961) <= not b;
    outputs(962) <= not (a or b);
    outputs(963) <= b;
    outputs(964) <= not a or b;
    outputs(965) <= b and not a;
    outputs(966) <= a or b;
    outputs(967) <= b;
    outputs(968) <= not (a and b);
    outputs(969) <= a and b;
    outputs(970) <= not (a xor b);
    outputs(971) <= not a;
    outputs(972) <= b and not a;
    outputs(973) <= b;
    outputs(974) <= b and not a;
    outputs(975) <= not b;
    outputs(976) <= not b;
    outputs(977) <= not (a or b);
    outputs(978) <= b and not a;
    outputs(979) <= a and not b;
    outputs(980) <= not (a xor b);
    outputs(981) <= not (a xor b);
    outputs(982) <= not a or b;
    outputs(983) <= b;
    outputs(984) <= b;
    outputs(985) <= not b;
    outputs(986) <= a xor b;
    outputs(987) <= b;
    outputs(988) <= not a;
    outputs(989) <= a xor b;
    outputs(990) <= a xor b;
    outputs(991) <= not b;
    outputs(992) <= b and not a;
    outputs(993) <= b and not a;
    outputs(994) <= not a;
    outputs(995) <= b;
    outputs(996) <= not a;
    outputs(997) <= a or b;
    outputs(998) <= not b;
    outputs(999) <= not (a xor b);
    outputs(1000) <= not a;
    outputs(1001) <= not b;
    outputs(1002) <= not b;
    outputs(1003) <= a and not b;
    outputs(1004) <= not b;
    outputs(1005) <= b;
    outputs(1006) <= b;
    outputs(1007) <= a;
    outputs(1008) <= b;
    outputs(1009) <= not a;
    outputs(1010) <= b;
    outputs(1011) <= a xor b;
    outputs(1012) <= a and b;
    outputs(1013) <= not a;
    outputs(1014) <= a xor b;
    outputs(1015) <= a and not b;
    outputs(1016) <= not (a xor b);
    outputs(1017) <= a and b;
    outputs(1018) <= not (a xor b);
    outputs(1019) <= not b;
    outputs(1020) <= not (a or b);
    outputs(1021) <= b and not a;
    outputs(1022) <= a;
    outputs(1023) <= a;
    outputs(1024) <= a xor b;
    outputs(1025) <= not (a and b);
    outputs(1026) <= a and not b;
    outputs(1027) <= a;
    outputs(1028) <= a xor b;
    outputs(1029) <= not a or b;
    outputs(1030) <= not (a xor b);
    outputs(1031) <= b;
    outputs(1032) <= a xor b;
    outputs(1033) <= not (a xor b);
    outputs(1034) <= b;
    outputs(1035) <= not (a or b);
    outputs(1036) <= b;
    outputs(1037) <= not a;
    outputs(1038) <= b and not a;
    outputs(1039) <= a or b;
    outputs(1040) <= not a or b;
    outputs(1041) <= b;
    outputs(1042) <= not a;
    outputs(1043) <= a and not b;
    outputs(1044) <= not a;
    outputs(1045) <= not b or a;
    outputs(1046) <= a;
    outputs(1047) <= a xor b;
    outputs(1048) <= b and not a;
    outputs(1049) <= b;
    outputs(1050) <= b;
    outputs(1051) <= a and b;
    outputs(1052) <= not b;
    outputs(1053) <= not b;
    outputs(1054) <= a;
    outputs(1055) <= a and b;
    outputs(1056) <= a xor b;
    outputs(1057) <= b;
    outputs(1058) <= not a;
    outputs(1059) <= b;
    outputs(1060) <= a and not b;
    outputs(1061) <= a xor b;
    outputs(1062) <= b;
    outputs(1063) <= a and not b;
    outputs(1064) <= a and not b;
    outputs(1065) <= a xor b;
    outputs(1066) <= not b;
    outputs(1067) <= a or b;
    outputs(1068) <= not (a xor b);
    outputs(1069) <= not b;
    outputs(1070) <= not b;
    outputs(1071) <= b and not a;
    outputs(1072) <= a;
    outputs(1073) <= a and b;
    outputs(1074) <= a xor b;
    outputs(1075) <= not (a and b);
    outputs(1076) <= not (a xor b);
    outputs(1077) <= a and not b;
    outputs(1078) <= not b or a;
    outputs(1079) <= a and not b;
    outputs(1080) <= a xor b;
    outputs(1081) <= not a;
    outputs(1082) <= a or b;
    outputs(1083) <= not b;
    outputs(1084) <= not b;
    outputs(1085) <= not a;
    outputs(1086) <= not a;
    outputs(1087) <= not (a or b);
    outputs(1088) <= not a or b;
    outputs(1089) <= b;
    outputs(1090) <= not b;
    outputs(1091) <= a and b;
    outputs(1092) <= not b;
    outputs(1093) <= not (a xor b);
    outputs(1094) <= b;
    outputs(1095) <= not (a or b);
    outputs(1096) <= not a;
    outputs(1097) <= not a;
    outputs(1098) <= a xor b;
    outputs(1099) <= a and not b;
    outputs(1100) <= b and not a;
    outputs(1101) <= a and b;
    outputs(1102) <= not b;
    outputs(1103) <= not b;
    outputs(1104) <= b;
    outputs(1105) <= b;
    outputs(1106) <= b and not a;
    outputs(1107) <= not a;
    outputs(1108) <= a xor b;
    outputs(1109) <= a and b;
    outputs(1110) <= b;
    outputs(1111) <= b;
    outputs(1112) <= not a;
    outputs(1113) <= not a;
    outputs(1114) <= not b;
    outputs(1115) <= not a;
    outputs(1116) <= a;
    outputs(1117) <= a;
    outputs(1118) <= a and b;
    outputs(1119) <= not a;
    outputs(1120) <= not a;
    outputs(1121) <= b;
    outputs(1122) <= a xor b;
    outputs(1123) <= not (a xor b);
    outputs(1124) <= a and b;
    outputs(1125) <= a and b;
    outputs(1126) <= a and not b;
    outputs(1127) <= not a;
    outputs(1128) <= not (a xor b);
    outputs(1129) <= a xor b;
    outputs(1130) <= a;
    outputs(1131) <= b and not a;
    outputs(1132) <= b and not a;
    outputs(1133) <= b;
    outputs(1134) <= a and not b;
    outputs(1135) <= a and not b;
    outputs(1136) <= b and not a;
    outputs(1137) <= not b;
    outputs(1138) <= not a;
    outputs(1139) <= a;
    outputs(1140) <= b;
    outputs(1141) <= not b;
    outputs(1142) <= b and not a;
    outputs(1143) <= a xor b;
    outputs(1144) <= b and not a;
    outputs(1145) <= not b;
    outputs(1146) <= a and b;
    outputs(1147) <= b and not a;
    outputs(1148) <= not b;
    outputs(1149) <= b;
    outputs(1150) <= not (a or b);
    outputs(1151) <= a xor b;
    outputs(1152) <= not a;
    outputs(1153) <= a;
    outputs(1154) <= b;
    outputs(1155) <= b;
    outputs(1156) <= not (a or b);
    outputs(1157) <= not a;
    outputs(1158) <= a;
    outputs(1159) <= not a;
    outputs(1160) <= not b;
    outputs(1161) <= b;
    outputs(1162) <= not b;
    outputs(1163) <= not a;
    outputs(1164) <= not b;
    outputs(1165) <= a;
    outputs(1166) <= a and b;
    outputs(1167) <= not b;
    outputs(1168) <= a;
    outputs(1169) <= not a;
    outputs(1170) <= a;
    outputs(1171) <= b;
    outputs(1172) <= a;
    outputs(1173) <= not b or a;
    outputs(1174) <= b and not a;
    outputs(1175) <= b;
    outputs(1176) <= not (a xor b);
    outputs(1177) <= a;
    outputs(1178) <= not b;
    outputs(1179) <= not b;
    outputs(1180) <= not (a or b);
    outputs(1181) <= not b;
    outputs(1182) <= b and not a;
    outputs(1183) <= a xor b;
    outputs(1184) <= not (a xor b);
    outputs(1185) <= a and b;
    outputs(1186) <= not (a or b);
    outputs(1187) <= not (a xor b);
    outputs(1188) <= a xor b;
    outputs(1189) <= a;
    outputs(1190) <= not b;
    outputs(1191) <= a;
    outputs(1192) <= a xor b;
    outputs(1193) <= not (a or b);
    outputs(1194) <= a xor b;
    outputs(1195) <= a xor b;
    outputs(1196) <= a or b;
    outputs(1197) <= a;
    outputs(1198) <= not b;
    outputs(1199) <= a and not b;
    outputs(1200) <= not b;
    outputs(1201) <= a;
    outputs(1202) <= a xor b;
    outputs(1203) <= not (a and b);
    outputs(1204) <= a;
    outputs(1205) <= b and not a;
    outputs(1206) <= a and b;
    outputs(1207) <= not b;
    outputs(1208) <= a;
    outputs(1209) <= not a;
    outputs(1210) <= not b;
    outputs(1211) <= not b;
    outputs(1212) <= a and b;
    outputs(1213) <= not b;
    outputs(1214) <= a and b;
    outputs(1215) <= a;
    outputs(1216) <= a and not b;
    outputs(1217) <= not a;
    outputs(1218) <= a and not b;
    outputs(1219) <= not (a xor b);
    outputs(1220) <= a and not b;
    outputs(1221) <= a xor b;
    outputs(1222) <= not (a xor b);
    outputs(1223) <= not a;
    outputs(1224) <= a xor b;
    outputs(1225) <= a and not b;
    outputs(1226) <= not (a xor b);
    outputs(1227) <= b and not a;
    outputs(1228) <= a xor b;
    outputs(1229) <= b;
    outputs(1230) <= a xor b;
    outputs(1231) <= a or b;
    outputs(1232) <= a xor b;
    outputs(1233) <= a and b;
    outputs(1234) <= a and not b;
    outputs(1235) <= b;
    outputs(1236) <= a and b;
    outputs(1237) <= not (a xor b);
    outputs(1238) <= a and b;
    outputs(1239) <= a xor b;
    outputs(1240) <= not (a xor b);
    outputs(1241) <= a;
    outputs(1242) <= b and not a;
    outputs(1243) <= a xor b;
    outputs(1244) <= not (a xor b);
    outputs(1245) <= a and b;
    outputs(1246) <= a xor b;
    outputs(1247) <= not b;
    outputs(1248) <= not a;
    outputs(1249) <= a;
    outputs(1250) <= a xor b;
    outputs(1251) <= b;
    outputs(1252) <= a and not b;
    outputs(1253) <= not (a xor b);
    outputs(1254) <= a xor b;
    outputs(1255) <= not (a or b);
    outputs(1256) <= not (a or b);
    outputs(1257) <= not (a xor b);
    outputs(1258) <= a;
    outputs(1259) <= a or b;
    outputs(1260) <= a or b;
    outputs(1261) <= a xor b;
    outputs(1262) <= not a;
    outputs(1263) <= not (a xor b);
    outputs(1264) <= b and not a;
    outputs(1265) <= not a;
    outputs(1266) <= a and not b;
    outputs(1267) <= not b;
    outputs(1268) <= not b;
    outputs(1269) <= a;
    outputs(1270) <= not b;
    outputs(1271) <= a;
    outputs(1272) <= b;
    outputs(1273) <= not a;
    outputs(1274) <= not b;
    outputs(1275) <= a;
    outputs(1276) <= not b;
    outputs(1277) <= a and b;
    outputs(1278) <= not b;
    outputs(1279) <= a and not b;
    outputs(1280) <= a;
    outputs(1281) <= b and not a;
    outputs(1282) <= b;
    outputs(1283) <= not a;
    outputs(1284) <= not (a xor b);
    outputs(1285) <= b and not a;
    outputs(1286) <= not b;
    outputs(1287) <= a and not b;
    outputs(1288) <= b and not a;
    outputs(1289) <= a xor b;
    outputs(1290) <= b and not a;
    outputs(1291) <= b;
    outputs(1292) <= a and b;
    outputs(1293) <= a;
    outputs(1294) <= a;
    outputs(1295) <= a and b;
    outputs(1296) <= not a;
    outputs(1297) <= not (a and b);
    outputs(1298) <= a and b;
    outputs(1299) <= b;
    outputs(1300) <= b;
    outputs(1301) <= not b;
    outputs(1302) <= a and b;
    outputs(1303) <= not b;
    outputs(1304) <= a;
    outputs(1305) <= not (a or b);
    outputs(1306) <= not b;
    outputs(1307) <= a;
    outputs(1308) <= not b;
    outputs(1309) <= not b;
    outputs(1310) <= a and b;
    outputs(1311) <= b and not a;
    outputs(1312) <= b;
    outputs(1313) <= not (a or b);
    outputs(1314) <= a;
    outputs(1315) <= not (a xor b);
    outputs(1316) <= not a or b;
    outputs(1317) <= not b;
    outputs(1318) <= not a;
    outputs(1319) <= a;
    outputs(1320) <= not a or b;
    outputs(1321) <= b;
    outputs(1322) <= a and not b;
    outputs(1323) <= a;
    outputs(1324) <= not a;
    outputs(1325) <= a and not b;
    outputs(1326) <= b;
    outputs(1327) <= a xor b;
    outputs(1328) <= not (a and b);
    outputs(1329) <= not b;
    outputs(1330) <= a xor b;
    outputs(1331) <= not b;
    outputs(1332) <= a and not b;
    outputs(1333) <= b;
    outputs(1334) <= not a;
    outputs(1335) <= not (a xor b);
    outputs(1336) <= a xor b;
    outputs(1337) <= not (a xor b);
    outputs(1338) <= not (a xor b);
    outputs(1339) <= a xor b;
    outputs(1340) <= not b;
    outputs(1341) <= not (a xor b);
    outputs(1342) <= a;
    outputs(1343) <= not b or a;
    outputs(1344) <= a xor b;
    outputs(1345) <= not (a xor b);
    outputs(1346) <= b and not a;
    outputs(1347) <= not b;
    outputs(1348) <= not b;
    outputs(1349) <= not b;
    outputs(1350) <= not (a xor b);
    outputs(1351) <= not a;
    outputs(1352) <= not (a or b);
    outputs(1353) <= not (a xor b);
    outputs(1354) <= a xor b;
    outputs(1355) <= a and b;
    outputs(1356) <= a xor b;
    outputs(1357) <= b;
    outputs(1358) <= a or b;
    outputs(1359) <= a;
    outputs(1360) <= not a or b;
    outputs(1361) <= b;
    outputs(1362) <= b;
    outputs(1363) <= b and not a;
    outputs(1364) <= b and not a;
    outputs(1365) <= a xor b;
    outputs(1366) <= not (a and b);
    outputs(1367) <= not a;
    outputs(1368) <= not a;
    outputs(1369) <= a and b;
    outputs(1370) <= not (a xor b);
    outputs(1371) <= a;
    outputs(1372) <= a and b;
    outputs(1373) <= b;
    outputs(1374) <= not b or a;
    outputs(1375) <= not a;
    outputs(1376) <= not b;
    outputs(1377) <= not b;
    outputs(1378) <= a;
    outputs(1379) <= b;
    outputs(1380) <= b;
    outputs(1381) <= b;
    outputs(1382) <= not b;
    outputs(1383) <= b and not a;
    outputs(1384) <= not b;
    outputs(1385) <= a and b;
    outputs(1386) <= b;
    outputs(1387) <= not b;
    outputs(1388) <= not (a or b);
    outputs(1389) <= not a;
    outputs(1390) <= a xor b;
    outputs(1391) <= a xor b;
    outputs(1392) <= a or b;
    outputs(1393) <= b;
    outputs(1394) <= not b;
    outputs(1395) <= not (a and b);
    outputs(1396) <= a xor b;
    outputs(1397) <= b and not a;
    outputs(1398) <= a;
    outputs(1399) <= b;
    outputs(1400) <= b;
    outputs(1401) <= b and not a;
    outputs(1402) <= not b;
    outputs(1403) <= not (a and b);
    outputs(1404) <= a xor b;
    outputs(1405) <= not (a and b);
    outputs(1406) <= b;
    outputs(1407) <= a xor b;
    outputs(1408) <= a xor b;
    outputs(1409) <= not (a xor b);
    outputs(1410) <= not b or a;
    outputs(1411) <= not a or b;
    outputs(1412) <= b;
    outputs(1413) <= not a;
    outputs(1414) <= not (a xor b);
    outputs(1415) <= a xor b;
    outputs(1416) <= not (a xor b);
    outputs(1417) <= a or b;
    outputs(1418) <= a or b;
    outputs(1419) <= b;
    outputs(1420) <= a xor b;
    outputs(1421) <= not b or a;
    outputs(1422) <= not a;
    outputs(1423) <= not a;
    outputs(1424) <= not (a or b);
    outputs(1425) <= not a;
    outputs(1426) <= not a;
    outputs(1427) <= not (a xor b);
    outputs(1428) <= not (a and b);
    outputs(1429) <= not b;
    outputs(1430) <= not a;
    outputs(1431) <= not (a or b);
    outputs(1432) <= b and not a;
    outputs(1433) <= not (a xor b);
    outputs(1434) <= not a;
    outputs(1435) <= a;
    outputs(1436) <= not (a xor b);
    outputs(1437) <= not a;
    outputs(1438) <= b and not a;
    outputs(1439) <= not b;
    outputs(1440) <= a;
    outputs(1441) <= not a;
    outputs(1442) <= b;
    outputs(1443) <= a xor b;
    outputs(1444) <= not (a xor b);
    outputs(1445) <= b;
    outputs(1446) <= b;
    outputs(1447) <= a;
    outputs(1448) <= not a;
    outputs(1449) <= a;
    outputs(1450) <= b and not a;
    outputs(1451) <= not (a or b);
    outputs(1452) <= not a;
    outputs(1453) <= not b;
    outputs(1454) <= a and not b;
    outputs(1455) <= b;
    outputs(1456) <= not (a xor b);
    outputs(1457) <= b;
    outputs(1458) <= a;
    outputs(1459) <= a xor b;
    outputs(1460) <= a xor b;
    outputs(1461) <= a and not b;
    outputs(1462) <= not (a or b);
    outputs(1463) <= not a;
    outputs(1464) <= not a or b;
    outputs(1465) <= a;
    outputs(1466) <= a xor b;
    outputs(1467) <= not b or a;
    outputs(1468) <= a;
    outputs(1469) <= not (a xor b);
    outputs(1470) <= a xor b;
    outputs(1471) <= not a;
    outputs(1472) <= not a or b;
    outputs(1473) <= a;
    outputs(1474) <= not a;
    outputs(1475) <= a;
    outputs(1476) <= not (a or b);
    outputs(1477) <= not (a xor b);
    outputs(1478) <= b and not a;
    outputs(1479) <= b;
    outputs(1480) <= not a or b;
    outputs(1481) <= b and not a;
    outputs(1482) <= b and not a;
    outputs(1483) <= not a;
    outputs(1484) <= not a;
    outputs(1485) <= not (a xor b);
    outputs(1486) <= b;
    outputs(1487) <= not b;
    outputs(1488) <= b and not a;
    outputs(1489) <= not (a or b);
    outputs(1490) <= a xor b;
    outputs(1491) <= not (a xor b);
    outputs(1492) <= b;
    outputs(1493) <= not b;
    outputs(1494) <= not b;
    outputs(1495) <= a;
    outputs(1496) <= a and not b;
    outputs(1497) <= a and b;
    outputs(1498) <= a and b;
    outputs(1499) <= not b;
    outputs(1500) <= not a;
    outputs(1501) <= not (a and b);
    outputs(1502) <= a or b;
    outputs(1503) <= b;
    outputs(1504) <= not (a xor b);
    outputs(1505) <= not a;
    outputs(1506) <= a;
    outputs(1507) <= a xor b;
    outputs(1508) <= not (a xor b);
    outputs(1509) <= not (a or b);
    outputs(1510) <= a xor b;
    outputs(1511) <= not (a xor b);
    outputs(1512) <= not b or a;
    outputs(1513) <= b;
    outputs(1514) <= not b;
    outputs(1515) <= a xor b;
    outputs(1516) <= not b;
    outputs(1517) <= not b;
    outputs(1518) <= a xor b;
    outputs(1519) <= a xor b;
    outputs(1520) <= not (a xor b);
    outputs(1521) <= a;
    outputs(1522) <= not b or a;
    outputs(1523) <= not (a or b);
    outputs(1524) <= not a;
    outputs(1525) <= a and not b;
    outputs(1526) <= a xor b;
    outputs(1527) <= b and not a;
    outputs(1528) <= a or b;
    outputs(1529) <= a xor b;
    outputs(1530) <= not (a xor b);
    outputs(1531) <= a xor b;
    outputs(1532) <= not (a xor b);
    outputs(1533) <= a and b;
    outputs(1534) <= not a;
    outputs(1535) <= not (a or b);
    outputs(1536) <= a xor b;
    outputs(1537) <= not a;
    outputs(1538) <= not b;
    outputs(1539) <= a xor b;
    outputs(1540) <= not b;
    outputs(1541) <= a xor b;
    outputs(1542) <= not (a xor b);
    outputs(1543) <= not a;
    outputs(1544) <= not b;
    outputs(1545) <= a;
    outputs(1546) <= not (a or b);
    outputs(1547) <= not (a or b);
    outputs(1548) <= b;
    outputs(1549) <= a xor b;
    outputs(1550) <= a;
    outputs(1551) <= not a;
    outputs(1552) <= a;
    outputs(1553) <= a xor b;
    outputs(1554) <= not (a xor b);
    outputs(1555) <= a and not b;
    outputs(1556) <= not (a or b);
    outputs(1557) <= not b;
    outputs(1558) <= not a;
    outputs(1559) <= not a;
    outputs(1560) <= a xor b;
    outputs(1561) <= a xor b;
    outputs(1562) <= a xor b;
    outputs(1563) <= a xor b;
    outputs(1564) <= not (a xor b);
    outputs(1565) <= b;
    outputs(1566) <= b and not a;
    outputs(1567) <= a and not b;
    outputs(1568) <= not b;
    outputs(1569) <= not a;
    outputs(1570) <= not (a or b);
    outputs(1571) <= b;
    outputs(1572) <= a and not b;
    outputs(1573) <= not b;
    outputs(1574) <= not (a xor b);
    outputs(1575) <= a xor b;
    outputs(1576) <= a;
    outputs(1577) <= b;
    outputs(1578) <= b;
    outputs(1579) <= b;
    outputs(1580) <= not a;
    outputs(1581) <= not a;
    outputs(1582) <= a and b;
    outputs(1583) <= not b;
    outputs(1584) <= a xor b;
    outputs(1585) <= not (a and b);
    outputs(1586) <= not a;
    outputs(1587) <= not a or b;
    outputs(1588) <= a;
    outputs(1589) <= not b;
    outputs(1590) <= b;
    outputs(1591) <= not (a xor b);
    outputs(1592) <= not a;
    outputs(1593) <= not b;
    outputs(1594) <= not (a xor b);
    outputs(1595) <= not (a or b);
    outputs(1596) <= not b;
    outputs(1597) <= a and not b;
    outputs(1598) <= b;
    outputs(1599) <= a;
    outputs(1600) <= b;
    outputs(1601) <= not a;
    outputs(1602) <= a xor b;
    outputs(1603) <= not (a xor b);
    outputs(1604) <= b;
    outputs(1605) <= not a;
    outputs(1606) <= a xor b;
    outputs(1607) <= a and not b;
    outputs(1608) <= not a;
    outputs(1609) <= a and b;
    outputs(1610) <= not a;
    outputs(1611) <= not a;
    outputs(1612) <= a and not b;
    outputs(1613) <= not (a and b);
    outputs(1614) <= a;
    outputs(1615) <= a xor b;
    outputs(1616) <= a xor b;
    outputs(1617) <= a;
    outputs(1618) <= not (a or b);
    outputs(1619) <= not b;
    outputs(1620) <= a and not b;
    outputs(1621) <= not (a xor b);
    outputs(1622) <= not (a xor b);
    outputs(1623) <= not b;
    outputs(1624) <= b;
    outputs(1625) <= not b;
    outputs(1626) <= not b;
    outputs(1627) <= not b;
    outputs(1628) <= a;
    outputs(1629) <= a or b;
    outputs(1630) <= a and b;
    outputs(1631) <= a;
    outputs(1632) <= not b;
    outputs(1633) <= b;
    outputs(1634) <= a;
    outputs(1635) <= not a;
    outputs(1636) <= not a or b;
    outputs(1637) <= a xor b;
    outputs(1638) <= a;
    outputs(1639) <= b and not a;
    outputs(1640) <= a xor b;
    outputs(1641) <= not (a xor b);
    outputs(1642) <= a;
    outputs(1643) <= a and not b;
    outputs(1644) <= not a;
    outputs(1645) <= not (a xor b);
    outputs(1646) <= b;
    outputs(1647) <= not a;
    outputs(1648) <= not b;
    outputs(1649) <= a and not b;
    outputs(1650) <= a;
    outputs(1651) <= a and not b;
    outputs(1652) <= a xor b;
    outputs(1653) <= a xor b;
    outputs(1654) <= b and not a;
    outputs(1655) <= not a;
    outputs(1656) <= a;
    outputs(1657) <= a xor b;
    outputs(1658) <= not (a or b);
    outputs(1659) <= b;
    outputs(1660) <= b and not a;
    outputs(1661) <= a;
    outputs(1662) <= not b;
    outputs(1663) <= a and not b;
    outputs(1664) <= b and not a;
    outputs(1665) <= a and b;
    outputs(1666) <= not (a and b);
    outputs(1667) <= not (a or b);
    outputs(1668) <= not b;
    outputs(1669) <= not a;
    outputs(1670) <= not (a or b);
    outputs(1671) <= a xor b;
    outputs(1672) <= a xor b;
    outputs(1673) <= b;
    outputs(1674) <= a xor b;
    outputs(1675) <= not b;
    outputs(1676) <= b;
    outputs(1677) <= a and b;
    outputs(1678) <= a or b;
    outputs(1679) <= not (a and b);
    outputs(1680) <= a xor b;
    outputs(1681) <= not a;
    outputs(1682) <= not (a xor b);
    outputs(1683) <= not a;
    outputs(1684) <= a xor b;
    outputs(1685) <= b;
    outputs(1686) <= b;
    outputs(1687) <= not a;
    outputs(1688) <= not (a xor b);
    outputs(1689) <= not (a or b);
    outputs(1690) <= not (a xor b);
    outputs(1691) <= b;
    outputs(1692) <= not b or a;
    outputs(1693) <= not (a or b);
    outputs(1694) <= not a;
    outputs(1695) <= a or b;
    outputs(1696) <= not (a or b);
    outputs(1697) <= not (a xor b);
    outputs(1698) <= b;
    outputs(1699) <= b and not a;
    outputs(1700) <= a xor b;
    outputs(1701) <= b;
    outputs(1702) <= a;
    outputs(1703) <= not (a or b);
    outputs(1704) <= a;
    outputs(1705) <= a xor b;
    outputs(1706) <= a xor b;
    outputs(1707) <= not b;
    outputs(1708) <= not a;
    outputs(1709) <= a xor b;
    outputs(1710) <= not a;
    outputs(1711) <= not b;
    outputs(1712) <= not a;
    outputs(1713) <= not b;
    outputs(1714) <= not b or a;
    outputs(1715) <= a xor b;
    outputs(1716) <= a xor b;
    outputs(1717) <= a;
    outputs(1718) <= b;
    outputs(1719) <= not b;
    outputs(1720) <= not (a xor b);
    outputs(1721) <= not a;
    outputs(1722) <= b;
    outputs(1723) <= a;
    outputs(1724) <= b;
    outputs(1725) <= not a;
    outputs(1726) <= not (a xor b);
    outputs(1727) <= not (a xor b);
    outputs(1728) <= a and b;
    outputs(1729) <= not (a xor b);
    outputs(1730) <= not a;
    outputs(1731) <= not (a xor b);
    outputs(1732) <= not a;
    outputs(1733) <= a;
    outputs(1734) <= not (a and b);
    outputs(1735) <= not a;
    outputs(1736) <= a and not b;
    outputs(1737) <= a;
    outputs(1738) <= a xor b;
    outputs(1739) <= not b;
    outputs(1740) <= not b;
    outputs(1741) <= a xor b;
    outputs(1742) <= a;
    outputs(1743) <= not b;
    outputs(1744) <= not b;
    outputs(1745) <= not (a xor b);
    outputs(1746) <= not (a xor b);
    outputs(1747) <= not (a xor b);
    outputs(1748) <= a xor b;
    outputs(1749) <= a xor b;
    outputs(1750) <= a;
    outputs(1751) <= not b or a;
    outputs(1752) <= b and not a;
    outputs(1753) <= b and not a;
    outputs(1754) <= not (a xor b);
    outputs(1755) <= not b;
    outputs(1756) <= not (a xor b);
    outputs(1757) <= a xor b;
    outputs(1758) <= not (a or b);
    outputs(1759) <= a xor b;
    outputs(1760) <= a;
    outputs(1761) <= a;
    outputs(1762) <= b and not a;
    outputs(1763) <= not a;
    outputs(1764) <= b and not a;
    outputs(1765) <= a xor b;
    outputs(1766) <= not b;
    outputs(1767) <= not (a or b);
    outputs(1768) <= not b;
    outputs(1769) <= a xor b;
    outputs(1770) <= not (a xor b);
    outputs(1771) <= not b or a;
    outputs(1772) <= b;
    outputs(1773) <= a xor b;
    outputs(1774) <= a xor b;
    outputs(1775) <= not a;
    outputs(1776) <= b and not a;
    outputs(1777) <= a xor b;
    outputs(1778) <= a;
    outputs(1779) <= not (a and b);
    outputs(1780) <= a or b;
    outputs(1781) <= not (a and b);
    outputs(1782) <= a and b;
    outputs(1783) <= a and b;
    outputs(1784) <= a or b;
    outputs(1785) <= not a;
    outputs(1786) <= a and b;
    outputs(1787) <= not (a and b);
    outputs(1788) <= not (a and b);
    outputs(1789) <= not (a or b);
    outputs(1790) <= not (a xor b);
    outputs(1791) <= a;
    outputs(1792) <= a and not b;
    outputs(1793) <= not (a xor b);
    outputs(1794) <= a;
    outputs(1795) <= not b;
    outputs(1796) <= b;
    outputs(1797) <= not b;
    outputs(1798) <= a;
    outputs(1799) <= not a;
    outputs(1800) <= not (a or b);
    outputs(1801) <= not (a xor b);
    outputs(1802) <= not a;
    outputs(1803) <= not a;
    outputs(1804) <= b and not a;
    outputs(1805) <= not (a xor b);
    outputs(1806) <= a and b;
    outputs(1807) <= not a;
    outputs(1808) <= a;
    outputs(1809) <= a;
    outputs(1810) <= a;
    outputs(1811) <= b;
    outputs(1812) <= not b;
    outputs(1813) <= not b;
    outputs(1814) <= not b;
    outputs(1815) <= b;
    outputs(1816) <= not (a or b);
    outputs(1817) <= a;
    outputs(1818) <= a and not b;
    outputs(1819) <= not (a xor b);
    outputs(1820) <= b;
    outputs(1821) <= a xor b;
    outputs(1822) <= a and not b;
    outputs(1823) <= not a;
    outputs(1824) <= b and not a;
    outputs(1825) <= a and b;
    outputs(1826) <= b;
    outputs(1827) <= not a;
    outputs(1828) <= not (a xor b);
    outputs(1829) <= not b;
    outputs(1830) <= not b or a;
    outputs(1831) <= a xor b;
    outputs(1832) <= b;
    outputs(1833) <= a;
    outputs(1834) <= not (a or b);
    outputs(1835) <= a and not b;
    outputs(1836) <= not a;
    outputs(1837) <= not a;
    outputs(1838) <= b;
    outputs(1839) <= b;
    outputs(1840) <= not a;
    outputs(1841) <= not a;
    outputs(1842) <= b;
    outputs(1843) <= not (a xor b);
    outputs(1844) <= a;
    outputs(1845) <= b;
    outputs(1846) <= not b;
    outputs(1847) <= a;
    outputs(1848) <= not (a xor b);
    outputs(1849) <= a and b;
    outputs(1850) <= a;
    outputs(1851) <= not (a or b);
    outputs(1852) <= not a or b;
    outputs(1853) <= not a;
    outputs(1854) <= a and b;
    outputs(1855) <= not a;
    outputs(1856) <= a xor b;
    outputs(1857) <= a and b;
    outputs(1858) <= a xor b;
    outputs(1859) <= b and not a;
    outputs(1860) <= b;
    outputs(1861) <= a xor b;
    outputs(1862) <= not (a or b);
    outputs(1863) <= a or b;
    outputs(1864) <= a;
    outputs(1865) <= b and not a;
    outputs(1866) <= a xor b;
    outputs(1867) <= a;
    outputs(1868) <= not b or a;
    outputs(1869) <= not b;
    outputs(1870) <= b;
    outputs(1871) <= a xor b;
    outputs(1872) <= not (a or b);
    outputs(1873) <= b;
    outputs(1874) <= not (a xor b);
    outputs(1875) <= not a;
    outputs(1876) <= b and not a;
    outputs(1877) <= not b;
    outputs(1878) <= a;
    outputs(1879) <= b;
    outputs(1880) <= a and not b;
    outputs(1881) <= not a;
    outputs(1882) <= b;
    outputs(1883) <= not (a xor b);
    outputs(1884) <= not (a or b);
    outputs(1885) <= not a;
    outputs(1886) <= not a;
    outputs(1887) <= b;
    outputs(1888) <= not (a xor b);
    outputs(1889) <= not a;
    outputs(1890) <= b;
    outputs(1891) <= not (a xor b);
    outputs(1892) <= not (a or b);
    outputs(1893) <= a;
    outputs(1894) <= a and b;
    outputs(1895) <= a;
    outputs(1896) <= a;
    outputs(1897) <= not b;
    outputs(1898) <= a xor b;
    outputs(1899) <= not a;
    outputs(1900) <= a and b;
    outputs(1901) <= a and b;
    outputs(1902) <= a;
    outputs(1903) <= a;
    outputs(1904) <= not (a xor b);
    outputs(1905) <= not (a or b);
    outputs(1906) <= not a or b;
    outputs(1907) <= a xor b;
    outputs(1908) <= not (a or b);
    outputs(1909) <= not a;
    outputs(1910) <= a xor b;
    outputs(1911) <= a xor b;
    outputs(1912) <= not (a or b);
    outputs(1913) <= not (a xor b);
    outputs(1914) <= a;
    outputs(1915) <= b and not a;
    outputs(1916) <= a and not b;
    outputs(1917) <= b;
    outputs(1918) <= a;
    outputs(1919) <= a xor b;
    outputs(1920) <= not (a or b);
    outputs(1921) <= b and not a;
    outputs(1922) <= a;
    outputs(1923) <= a and not b;
    outputs(1924) <= b and not a;
    outputs(1925) <= a;
    outputs(1926) <= a and not b;
    outputs(1927) <= a xor b;
    outputs(1928) <= not a or b;
    outputs(1929) <= a and b;
    outputs(1930) <= not b;
    outputs(1931) <= a xor b;
    outputs(1932) <= b;
    outputs(1933) <= not b;
    outputs(1934) <= b;
    outputs(1935) <= b and not a;
    outputs(1936) <= not a;
    outputs(1937) <= not a;
    outputs(1938) <= not (a xor b);
    outputs(1939) <= a;
    outputs(1940) <= not b;
    outputs(1941) <= not b;
    outputs(1942) <= a;
    outputs(1943) <= a and b;
    outputs(1944) <= not a;
    outputs(1945) <= a xor b;
    outputs(1946) <= a and not b;
    outputs(1947) <= a and b;
    outputs(1948) <= b;
    outputs(1949) <= not (a and b);
    outputs(1950) <= not b;
    outputs(1951) <= not b;
    outputs(1952) <= not b;
    outputs(1953) <= not a;
    outputs(1954) <= b;
    outputs(1955) <= a xor b;
    outputs(1956) <= not a;
    outputs(1957) <= a;
    outputs(1958) <= not a;
    outputs(1959) <= a;
    outputs(1960) <= not (a xor b);
    outputs(1961) <= a xor b;
    outputs(1962) <= b and not a;
    outputs(1963) <= not (a or b);
    outputs(1964) <= b;
    outputs(1965) <= not (a xor b);
    outputs(1966) <= b;
    outputs(1967) <= a;
    outputs(1968) <= a and not b;
    outputs(1969) <= a and not b;
    outputs(1970) <= a;
    outputs(1971) <= not a or b;
    outputs(1972) <= a;
    outputs(1973) <= a xor b;
    outputs(1974) <= a xor b;
    outputs(1975) <= b;
    outputs(1976) <= not (a xor b);
    outputs(1977) <= not a;
    outputs(1978) <= not b;
    outputs(1979) <= a xor b;
    outputs(1980) <= a and b;
    outputs(1981) <= not a;
    outputs(1982) <= a and b;
    outputs(1983) <= b;
    outputs(1984) <= not a;
    outputs(1985) <= a;
    outputs(1986) <= a or b;
    outputs(1987) <= not a;
    outputs(1988) <= a;
    outputs(1989) <= not b;
    outputs(1990) <= a xor b;
    outputs(1991) <= not a;
    outputs(1992) <= a and not b;
    outputs(1993) <= not a or b;
    outputs(1994) <= a and b;
    outputs(1995) <= not b;
    outputs(1996) <= not a;
    outputs(1997) <= a xor b;
    outputs(1998) <= a and not b;
    outputs(1999) <= not a;
    outputs(2000) <= not a;
    outputs(2001) <= a xor b;
    outputs(2002) <= not (a xor b);
    outputs(2003) <= a;
    outputs(2004) <= not a;
    outputs(2005) <= a xor b;
    outputs(2006) <= a and not b;
    outputs(2007) <= not (a xor b);
    outputs(2008) <= not a or b;
    outputs(2009) <= b;
    outputs(2010) <= not (a xor b);
    outputs(2011) <= a and b;
    outputs(2012) <= a and b;
    outputs(2013) <= a;
    outputs(2014) <= not b;
    outputs(2015) <= a;
    outputs(2016) <= a and not b;
    outputs(2017) <= not (a xor b);
    outputs(2018) <= not (a xor b);
    outputs(2019) <= not (a and b);
    outputs(2020) <= b;
    outputs(2021) <= a and b;
    outputs(2022) <= b and not a;
    outputs(2023) <= not (a xor b);
    outputs(2024) <= not (a or b);
    outputs(2025) <= a and b;
    outputs(2026) <= not b;
    outputs(2027) <= a and not b;
    outputs(2028) <= a xor b;
    outputs(2029) <= not b;
    outputs(2030) <= a and not b;
    outputs(2031) <= b;
    outputs(2032) <= not (a or b);
    outputs(2033) <= a;
    outputs(2034) <= b and not a;
    outputs(2035) <= a;
    outputs(2036) <= a xor b;
    outputs(2037) <= not (a xor b);
    outputs(2038) <= b and not a;
    outputs(2039) <= b;
    outputs(2040) <= b;
    outputs(2041) <= not (a or b);
    outputs(2042) <= not (a or b);
    outputs(2043) <= not b;
    outputs(2044) <= b and not a;
    outputs(2045) <= a;
    outputs(2046) <= a xor b;
    outputs(2047) <= not (a xor b);
    outputs(2048) <= not (a and b);
    outputs(2049) <= a and not b;
    outputs(2050) <= not (a xor b);
    outputs(2051) <= a;
    outputs(2052) <= b and not a;
    outputs(2053) <= b and not a;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= a xor b;
    outputs(2056) <= b and not a;
    outputs(2057) <= b;
    outputs(2058) <= a;
    outputs(2059) <= not a;
    outputs(2060) <= a or b;
    outputs(2061) <= a;
    outputs(2062) <= not a;
    outputs(2063) <= a xor b;
    outputs(2064) <= a;
    outputs(2065) <= not (a or b);
    outputs(2066) <= a and not b;
    outputs(2067) <= not b;
    outputs(2068) <= not a;
    outputs(2069) <= not b;
    outputs(2070) <= a xor b;
    outputs(2071) <= a xor b;
    outputs(2072) <= b;
    outputs(2073) <= not (a xor b);
    outputs(2074) <= not a or b;
    outputs(2075) <= b and not a;
    outputs(2076) <= a and b;
    outputs(2077) <= not (a xor b);
    outputs(2078) <= not (a xor b);
    outputs(2079) <= not (a or b);
    outputs(2080) <= b;
    outputs(2081) <= not a;
    outputs(2082) <= b and not a;
    outputs(2083) <= not (a and b);
    outputs(2084) <= b;
    outputs(2085) <= not b;
    outputs(2086) <= not (a and b);
    outputs(2087) <= not b or a;
    outputs(2088) <= not a;
    outputs(2089) <= a;
    outputs(2090) <= b and not a;
    outputs(2091) <= not (a and b);
    outputs(2092) <= not a or b;
    outputs(2093) <= b;
    outputs(2094) <= not b;
    outputs(2095) <= a xor b;
    outputs(2096) <= not b;
    outputs(2097) <= a and b;
    outputs(2098) <= not (a or b);
    outputs(2099) <= not (a xor b);
    outputs(2100) <= not a;
    outputs(2101) <= a and b;
    outputs(2102) <= not (a xor b);
    outputs(2103) <= a xor b;
    outputs(2104) <= not b;
    outputs(2105) <= not a;
    outputs(2106) <= a xor b;
    outputs(2107) <= not (a or b);
    outputs(2108) <= b;
    outputs(2109) <= a xor b;
    outputs(2110) <= b and not a;
    outputs(2111) <= b and not a;
    outputs(2112) <= b and not a;
    outputs(2113) <= a and not b;
    outputs(2114) <= a and not b;
    outputs(2115) <= b;
    outputs(2116) <= not a;
    outputs(2117) <= not (a xor b);
    outputs(2118) <= a and not b;
    outputs(2119) <= b;
    outputs(2120) <= a xor b;
    outputs(2121) <= not (a or b);
    outputs(2122) <= b;
    outputs(2123) <= not b;
    outputs(2124) <= a and b;
    outputs(2125) <= not (a or b);
    outputs(2126) <= a xor b;
    outputs(2127) <= a xor b;
    outputs(2128) <= a or b;
    outputs(2129) <= b and not a;
    outputs(2130) <= not (a xor b);
    outputs(2131) <= not (a xor b);
    outputs(2132) <= a and not b;
    outputs(2133) <= not (a xor b);
    outputs(2134) <= b;
    outputs(2135) <= a;
    outputs(2136) <= not (a and b);
    outputs(2137) <= not a;
    outputs(2138) <= not a;
    outputs(2139) <= b and not a;
    outputs(2140) <= not (a xor b);
    outputs(2141) <= not a;
    outputs(2142) <= b;
    outputs(2143) <= b and not a;
    outputs(2144) <= not (a xor b);
    outputs(2145) <= not (a xor b);
    outputs(2146) <= a and b;
    outputs(2147) <= not b;
    outputs(2148) <= a and b;
    outputs(2149) <= a;
    outputs(2150) <= a xor b;
    outputs(2151) <= not (a xor b);
    outputs(2152) <= not b;
    outputs(2153) <= b;
    outputs(2154) <= not (a xor b);
    outputs(2155) <= not (a xor b);
    outputs(2156) <= not (a or b);
    outputs(2157) <= not b;
    outputs(2158) <= a xor b;
    outputs(2159) <= a xor b;
    outputs(2160) <= a;
    outputs(2161) <= a;
    outputs(2162) <= a and not b;
    outputs(2163) <= not a;
    outputs(2164) <= not b;
    outputs(2165) <= a;
    outputs(2166) <= not (a xor b);
    outputs(2167) <= not (a or b);
    outputs(2168) <= a xor b;
    outputs(2169) <= b;
    outputs(2170) <= not (a xor b);
    outputs(2171) <= a xor b;
    outputs(2172) <= not a;
    outputs(2173) <= b;
    outputs(2174) <= not b;
    outputs(2175) <= a xor b;
    outputs(2176) <= a and not b;
    outputs(2177) <= not (a and b);
    outputs(2178) <= not a;
    outputs(2179) <= not (a xor b);
    outputs(2180) <= a xor b;
    outputs(2181) <= not (a xor b);
    outputs(2182) <= a xor b;
    outputs(2183) <= not (a or b);
    outputs(2184) <= a xor b;
    outputs(2185) <= a xor b;
    outputs(2186) <= b;
    outputs(2187) <= b and not a;
    outputs(2188) <= not (a xor b);
    outputs(2189) <= a and b;
    outputs(2190) <= b;
    outputs(2191) <= not b or a;
    outputs(2192) <= not a;
    outputs(2193) <= a xor b;
    outputs(2194) <= a xor b;
    outputs(2195) <= not a;
    outputs(2196) <= b and not a;
    outputs(2197) <= a;
    outputs(2198) <= not b;
    outputs(2199) <= not (a or b);
    outputs(2200) <= b;
    outputs(2201) <= not (a xor b);
    outputs(2202) <= a and b;
    outputs(2203) <= not b;
    outputs(2204) <= not a;
    outputs(2205) <= a xor b;
    outputs(2206) <= not (a xor b);
    outputs(2207) <= not (a or b);
    outputs(2208) <= a and b;
    outputs(2209) <= not (a xor b);
    outputs(2210) <= not (a xor b);
    outputs(2211) <= not a;
    outputs(2212) <= b and not a;
    outputs(2213) <= a xor b;
    outputs(2214) <= a and b;
    outputs(2215) <= not (a xor b);
    outputs(2216) <= not b;
    outputs(2217) <= not a;
    outputs(2218) <= a;
    outputs(2219) <= not (a xor b);
    outputs(2220) <= not a;
    outputs(2221) <= b;
    outputs(2222) <= a and b;
    outputs(2223) <= a and b;
    outputs(2224) <= not b;
    outputs(2225) <= a;
    outputs(2226) <= a;
    outputs(2227) <= a and not b;
    outputs(2228) <= a and b;
    outputs(2229) <= a and b;
    outputs(2230) <= a xor b;
    outputs(2231) <= not (a or b);
    outputs(2232) <= not (a and b);
    outputs(2233) <= not a;
    outputs(2234) <= not (a xor b);
    outputs(2235) <= not (a and b);
    outputs(2236) <= b;
    outputs(2237) <= b and not a;
    outputs(2238) <= a xor b;
    outputs(2239) <= b;
    outputs(2240) <= a and not b;
    outputs(2241) <= b and not a;
    outputs(2242) <= not (a or b);
    outputs(2243) <= not b;
    outputs(2244) <= a and b;
    outputs(2245) <= a xor b;
    outputs(2246) <= not (a and b);
    outputs(2247) <= b;
    outputs(2248) <= a xor b;
    outputs(2249) <= b;
    outputs(2250) <= a and not b;
    outputs(2251) <= b;
    outputs(2252) <= not a;
    outputs(2253) <= a and b;
    outputs(2254) <= b and not a;
    outputs(2255) <= b and not a;
    outputs(2256) <= b and not a;
    outputs(2257) <= not b;
    outputs(2258) <= a;
    outputs(2259) <= not a;
    outputs(2260) <= not a;
    outputs(2261) <= not (a xor b);
    outputs(2262) <= not (a xor b);
    outputs(2263) <= not (a xor b);
    outputs(2264) <= not b;
    outputs(2265) <= a and b;
    outputs(2266) <= not (a or b);
    outputs(2267) <= not a;
    outputs(2268) <= a and not b;
    outputs(2269) <= b and not a;
    outputs(2270) <= not a;
    outputs(2271) <= a and not b;
    outputs(2272) <= a and b;
    outputs(2273) <= not a;
    outputs(2274) <= not (a and b);
    outputs(2275) <= a and b;
    outputs(2276) <= not (a xor b);
    outputs(2277) <= a and not b;
    outputs(2278) <= a xor b;
    outputs(2279) <= a and not b;
    outputs(2280) <= not a;
    outputs(2281) <= a;
    outputs(2282) <= b;
    outputs(2283) <= not (a xor b);
    outputs(2284) <= not b;
    outputs(2285) <= a and not b;
    outputs(2286) <= not b or a;
    outputs(2287) <= a xor b;
    outputs(2288) <= not a;
    outputs(2289) <= not (a xor b);
    outputs(2290) <= b;
    outputs(2291) <= a or b;
    outputs(2292) <= a and not b;
    outputs(2293) <= not (a or b);
    outputs(2294) <= not a or b;
    outputs(2295) <= not a;
    outputs(2296) <= not b or a;
    outputs(2297) <= not (a or b);
    outputs(2298) <= a xor b;
    outputs(2299) <= not a;
    outputs(2300) <= not b;
    outputs(2301) <= not a or b;
    outputs(2302) <= a;
    outputs(2303) <= not (a xor b);
    outputs(2304) <= a and b;
    outputs(2305) <= not (a xor b);
    outputs(2306) <= not (a xor b);
    outputs(2307) <= not b or a;
    outputs(2308) <= a xor b;
    outputs(2309) <= b and not a;
    outputs(2310) <= not a;
    outputs(2311) <= not a;
    outputs(2312) <= not (a or b);
    outputs(2313) <= not b;
    outputs(2314) <= not b;
    outputs(2315) <= not b;
    outputs(2316) <= a or b;
    outputs(2317) <= not a;
    outputs(2318) <= not b;
    outputs(2319) <= a or b;
    outputs(2320) <= b;
    outputs(2321) <= b and not a;
    outputs(2322) <= a and not b;
    outputs(2323) <= a and not b;
    outputs(2324) <= a;
    outputs(2325) <= a;
    outputs(2326) <= not a;
    outputs(2327) <= not b;
    outputs(2328) <= not b or a;
    outputs(2329) <= a xor b;
    outputs(2330) <= b;
    outputs(2331) <= b and not a;
    outputs(2332) <= not (a xor b);
    outputs(2333) <= a and not b;
    outputs(2334) <= not (a xor b);
    outputs(2335) <= a and not b;
    outputs(2336) <= a;
    outputs(2337) <= not b;
    outputs(2338) <= a xor b;
    outputs(2339) <= b;
    outputs(2340) <= not (a and b);
    outputs(2341) <= a and b;
    outputs(2342) <= not b or a;
    outputs(2343) <= not b;
    outputs(2344) <= not a or b;
    outputs(2345) <= a;
    outputs(2346) <= b;
    outputs(2347) <= not a;
    outputs(2348) <= a and b;
    outputs(2349) <= a xor b;
    outputs(2350) <= a xor b;
    outputs(2351) <= b;
    outputs(2352) <= not b;
    outputs(2353) <= a and b;
    outputs(2354) <= a;
    outputs(2355) <= b;
    outputs(2356) <= a;
    outputs(2357) <= not b;
    outputs(2358) <= not b or a;
    outputs(2359) <= a;
    outputs(2360) <= not a;
    outputs(2361) <= not (a xor b);
    outputs(2362) <= not a;
    outputs(2363) <= a;
    outputs(2364) <= b;
    outputs(2365) <= a;
    outputs(2366) <= b and not a;
    outputs(2367) <= a and b;
    outputs(2368) <= not (a or b);
    outputs(2369) <= b;
    outputs(2370) <= not (a or b);
    outputs(2371) <= b and not a;
    outputs(2372) <= not (a xor b);
    outputs(2373) <= not (a xor b);
    outputs(2374) <= not a;
    outputs(2375) <= not b;
    outputs(2376) <= b and not a;
    outputs(2377) <= b;
    outputs(2378) <= a and b;
    outputs(2379) <= a and b;
    outputs(2380) <= a and b;
    outputs(2381) <= b and not a;
    outputs(2382) <= a and not b;
    outputs(2383) <= a xor b;
    outputs(2384) <= b and not a;
    outputs(2385) <= b;
    outputs(2386) <= b;
    outputs(2387) <= a;
    outputs(2388) <= not b or a;
    outputs(2389) <= a xor b;
    outputs(2390) <= b and not a;
    outputs(2391) <= not (a xor b);
    outputs(2392) <= a or b;
    outputs(2393) <= not (a xor b);
    outputs(2394) <= not a;
    outputs(2395) <= not (a or b);
    outputs(2396) <= b;
    outputs(2397) <= not b;
    outputs(2398) <= not a or b;
    outputs(2399) <= a xor b;
    outputs(2400) <= a and b;
    outputs(2401) <= not b;
    outputs(2402) <= not (a or b);
    outputs(2403) <= not a;
    outputs(2404) <= a xor b;
    outputs(2405) <= a xor b;
    outputs(2406) <= a xor b;
    outputs(2407) <= b and not a;
    outputs(2408) <= b;
    outputs(2409) <= a xor b;
    outputs(2410) <= not (a xor b);
    outputs(2411) <= not a;
    outputs(2412) <= not b or a;
    outputs(2413) <= not a;
    outputs(2414) <= a;
    outputs(2415) <= b and not a;
    outputs(2416) <= a or b;
    outputs(2417) <= not b;
    outputs(2418) <= b;
    outputs(2419) <= a;
    outputs(2420) <= a and not b;
    outputs(2421) <= a and b;
    outputs(2422) <= a xor b;
    outputs(2423) <= a and not b;
    outputs(2424) <= b and not a;
    outputs(2425) <= b;
    outputs(2426) <= not (a or b);
    outputs(2427) <= a;
    outputs(2428) <= not (a or b);
    outputs(2429) <= not b or a;
    outputs(2430) <= not b;
    outputs(2431) <= not (a xor b);
    outputs(2432) <= a xor b;
    outputs(2433) <= b and not a;
    outputs(2434) <= b;
    outputs(2435) <= a;
    outputs(2436) <= not a;
    outputs(2437) <= b;
    outputs(2438) <= b and not a;
    outputs(2439) <= not b or a;
    outputs(2440) <= a and b;
    outputs(2441) <= b;
    outputs(2442) <= b;
    outputs(2443) <= a xor b;
    outputs(2444) <= not (a xor b);
    outputs(2445) <= not (a xor b);
    outputs(2446) <= not (a xor b);
    outputs(2447) <= a and not b;
    outputs(2448) <= not b;
    outputs(2449) <= not (a xor b);
    outputs(2450) <= a xor b;
    outputs(2451) <= b;
    outputs(2452) <= b and not a;
    outputs(2453) <= a;
    outputs(2454) <= b;
    outputs(2455) <= a or b;
    outputs(2456) <= not a;
    outputs(2457) <= a and b;
    outputs(2458) <= not (a and b);
    outputs(2459) <= a xor b;
    outputs(2460) <= a xor b;
    outputs(2461) <= not b;
    outputs(2462) <= a and not b;
    outputs(2463) <= a and not b;
    outputs(2464) <= a and b;
    outputs(2465) <= a and b;
    outputs(2466) <= not (a or b);
    outputs(2467) <= not (a xor b);
    outputs(2468) <= not (a xor b);
    outputs(2469) <= not a or b;
    outputs(2470) <= not (a xor b);
    outputs(2471) <= b;
    outputs(2472) <= b;
    outputs(2473) <= not a;
    outputs(2474) <= a xor b;
    outputs(2475) <= b and not a;
    outputs(2476) <= not b;
    outputs(2477) <= not b;
    outputs(2478) <= not (a and b);
    outputs(2479) <= a or b;
    outputs(2480) <= b;
    outputs(2481) <= a and not b;
    outputs(2482) <= not b;
    outputs(2483) <= b;
    outputs(2484) <= not (a or b);
    outputs(2485) <= a or b;
    outputs(2486) <= not (a xor b);
    outputs(2487) <= not (a or b);
    outputs(2488) <= a or b;
    outputs(2489) <= not b;
    outputs(2490) <= not b;
    outputs(2491) <= a and b;
    outputs(2492) <= not b;
    outputs(2493) <= not b;
    outputs(2494) <= not a;
    outputs(2495) <= a;
    outputs(2496) <= a and b;
    outputs(2497) <= not (a xor b);
    outputs(2498) <= not a;
    outputs(2499) <= a and b;
    outputs(2500) <= a and not b;
    outputs(2501) <= a;
    outputs(2502) <= a xor b;
    outputs(2503) <= a and not b;
    outputs(2504) <= b and not a;
    outputs(2505) <= not b;
    outputs(2506) <= not a;
    outputs(2507) <= a and b;
    outputs(2508) <= not a;
    outputs(2509) <= a and b;
    outputs(2510) <= not b;
    outputs(2511) <= a and b;
    outputs(2512) <= b;
    outputs(2513) <= not (a and b);
    outputs(2514) <= not a;
    outputs(2515) <= not (a or b);
    outputs(2516) <= not a;
    outputs(2517) <= b and not a;
    outputs(2518) <= a xor b;
    outputs(2519) <= a and b;
    outputs(2520) <= not b;
    outputs(2521) <= a xor b;
    outputs(2522) <= not (a xor b);
    outputs(2523) <= b and not a;
    outputs(2524) <= not (a or b);
    outputs(2525) <= a and b;
    outputs(2526) <= not (a xor b);
    outputs(2527) <= a xor b;
    outputs(2528) <= not a;
    outputs(2529) <= not (a or b);
    outputs(2530) <= a and b;
    outputs(2531) <= not b;
    outputs(2532) <= a xor b;
    outputs(2533) <= b;
    outputs(2534) <= not (a xor b);
    outputs(2535) <= b and not a;
    outputs(2536) <= a xor b;
    outputs(2537) <= b and not a;
    outputs(2538) <= not b;
    outputs(2539) <= a;
    outputs(2540) <= b;
    outputs(2541) <= a xor b;
    outputs(2542) <= a and not b;
    outputs(2543) <= not (a or b);
    outputs(2544) <= not (a or b);
    outputs(2545) <= b;
    outputs(2546) <= not (a or b);
    outputs(2547) <= b;
    outputs(2548) <= b;
    outputs(2549) <= b and not a;
    outputs(2550) <= a;
    outputs(2551) <= a xor b;
    outputs(2552) <= not b or a;
    outputs(2553) <= not (a or b);
    outputs(2554) <= b;
    outputs(2555) <= a and b;
    outputs(2556) <= not (a xor b);
    outputs(2557) <= a and b;
    outputs(2558) <= a and b;
    outputs(2559) <= a and b;
end Behavioral;
