library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(5119 downto 0);
    signal layer1_outputs: std_logic_vector(5119 downto 0);
    signal layer2_outputs: std_logic_vector(5119 downto 0);
    signal layer3_outputs: std_logic_vector(5119 downto 0);
    signal layer4_outputs: std_logic_vector(5119 downto 0);

begin
    layer0_outputs(0) <= b;
    layer0_outputs(1) <= a xor b;
    layer0_outputs(2) <= not (a or b);
    layer0_outputs(3) <= not a or b;
    layer0_outputs(4) <= not b or a;
    layer0_outputs(5) <= '0';
    layer0_outputs(6) <= not a or b;
    layer0_outputs(7) <= '0';
    layer0_outputs(8) <= not a or b;
    layer0_outputs(9) <= not (a xor b);
    layer0_outputs(10) <= not a or b;
    layer0_outputs(11) <= '0';
    layer0_outputs(12) <= not (a xor b);
    layer0_outputs(13) <= b and not a;
    layer0_outputs(14) <= b;
    layer0_outputs(15) <= not (a or b);
    layer0_outputs(16) <= not a or b;
    layer0_outputs(17) <= b and not a;
    layer0_outputs(18) <= not (a or b);
    layer0_outputs(19) <= not (a and b);
    layer0_outputs(20) <= b and not a;
    layer0_outputs(21) <= a xor b;
    layer0_outputs(22) <= b;
    layer0_outputs(23) <= not a or b;
    layer0_outputs(24) <= a;
    layer0_outputs(25) <= a;
    layer0_outputs(26) <= not (a or b);
    layer0_outputs(27) <= a or b;
    layer0_outputs(28) <= not a;
    layer0_outputs(29) <= not (a and b);
    layer0_outputs(30) <= b;
    layer0_outputs(31) <= not a or b;
    layer0_outputs(32) <= b;
    layer0_outputs(33) <= a or b;
    layer0_outputs(34) <= not (a or b);
    layer0_outputs(35) <= a;
    layer0_outputs(36) <= a;
    layer0_outputs(37) <= not (a and b);
    layer0_outputs(38) <= a;
    layer0_outputs(39) <= a and not b;
    layer0_outputs(40) <= not (a and b);
    layer0_outputs(41) <= not (a and b);
    layer0_outputs(42) <= a or b;
    layer0_outputs(43) <= not (a or b);
    layer0_outputs(44) <= not a;
    layer0_outputs(45) <= b and not a;
    layer0_outputs(46) <= a and b;
    layer0_outputs(47) <= '0';
    layer0_outputs(48) <= b and not a;
    layer0_outputs(49) <= a and not b;
    layer0_outputs(50) <= not (a and b);
    layer0_outputs(51) <= a or b;
    layer0_outputs(52) <= not a;
    layer0_outputs(53) <= not (a or b);
    layer0_outputs(54) <= not b;
    layer0_outputs(55) <= not (a xor b);
    layer0_outputs(56) <= b and not a;
    layer0_outputs(57) <= b;
    layer0_outputs(58) <= a or b;
    layer0_outputs(59) <= a or b;
    layer0_outputs(60) <= not (a or b);
    layer0_outputs(61) <= '1';
    layer0_outputs(62) <= a or b;
    layer0_outputs(63) <= not (a or b);
    layer0_outputs(64) <= b;
    layer0_outputs(65) <= b;
    layer0_outputs(66) <= not (a and b);
    layer0_outputs(67) <= a;
    layer0_outputs(68) <= '1';
    layer0_outputs(69) <= a and b;
    layer0_outputs(70) <= b;
    layer0_outputs(71) <= '1';
    layer0_outputs(72) <= '0';
    layer0_outputs(73) <= a or b;
    layer0_outputs(74) <= a or b;
    layer0_outputs(75) <= not b;
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= not b or a;
    layer0_outputs(78) <= not b or a;
    layer0_outputs(79) <= a or b;
    layer0_outputs(80) <= b and not a;
    layer0_outputs(81) <= a or b;
    layer0_outputs(82) <= a and not b;
    layer0_outputs(83) <= not a;
    layer0_outputs(84) <= not b;
    layer0_outputs(85) <= a;
    layer0_outputs(86) <= not b;
    layer0_outputs(87) <= not (a or b);
    layer0_outputs(88) <= '1';
    layer0_outputs(89) <= not a or b;
    layer0_outputs(90) <= not b;
    layer0_outputs(91) <= not a;
    layer0_outputs(92) <= b;
    layer0_outputs(93) <= not (a or b);
    layer0_outputs(94) <= not (a xor b);
    layer0_outputs(95) <= not (a or b);
    layer0_outputs(96) <= a and not b;
    layer0_outputs(97) <= a;
    layer0_outputs(98) <= '0';
    layer0_outputs(99) <= b;
    layer0_outputs(100) <= a or b;
    layer0_outputs(101) <= not (a xor b);
    layer0_outputs(102) <= b and not a;
    layer0_outputs(103) <= a;
    layer0_outputs(104) <= b and not a;
    layer0_outputs(105) <= b;
    layer0_outputs(106) <= b and not a;
    layer0_outputs(107) <= a or b;
    layer0_outputs(108) <= a xor b;
    layer0_outputs(109) <= not (a or b);
    layer0_outputs(110) <= a or b;
    layer0_outputs(111) <= not a or b;
    layer0_outputs(112) <= not a;
    layer0_outputs(113) <= not a or b;
    layer0_outputs(114) <= not b or a;
    layer0_outputs(115) <= '0';
    layer0_outputs(116) <= b;
    layer0_outputs(117) <= a and not b;
    layer0_outputs(118) <= a or b;
    layer0_outputs(119) <= not (a or b);
    layer0_outputs(120) <= not b;
    layer0_outputs(121) <= b;
    layer0_outputs(122) <= a xor b;
    layer0_outputs(123) <= not (a or b);
    layer0_outputs(124) <= not b or a;
    layer0_outputs(125) <= not (a xor b);
    layer0_outputs(126) <= not (a or b);
    layer0_outputs(127) <= '1';
    layer0_outputs(128) <= not a or b;
    layer0_outputs(129) <= not a or b;
    layer0_outputs(130) <= not b or a;
    layer0_outputs(131) <= a or b;
    layer0_outputs(132) <= not a;
    layer0_outputs(133) <= not (a or b);
    layer0_outputs(134) <= not b;
    layer0_outputs(135) <= a and not b;
    layer0_outputs(136) <= b;
    layer0_outputs(137) <= b and not a;
    layer0_outputs(138) <= a;
    layer0_outputs(139) <= not (a and b);
    layer0_outputs(140) <= not a;
    layer0_outputs(141) <= a or b;
    layer0_outputs(142) <= a or b;
    layer0_outputs(143) <= '0';
    layer0_outputs(144) <= '0';
    layer0_outputs(145) <= b and not a;
    layer0_outputs(146) <= not a or b;
    layer0_outputs(147) <= b;
    layer0_outputs(148) <= a;
    layer0_outputs(149) <= not a;
    layer0_outputs(150) <= '1';
    layer0_outputs(151) <= b and not a;
    layer0_outputs(152) <= not b or a;
    layer0_outputs(153) <= not (a xor b);
    layer0_outputs(154) <= not a;
    layer0_outputs(155) <= b and not a;
    layer0_outputs(156) <= not a or b;
    layer0_outputs(157) <= not (a or b);
    layer0_outputs(158) <= a or b;
    layer0_outputs(159) <= not (a and b);
    layer0_outputs(160) <= not b or a;
    layer0_outputs(161) <= '0';
    layer0_outputs(162) <= not a or b;
    layer0_outputs(163) <= not a or b;
    layer0_outputs(164) <= not b or a;
    layer0_outputs(165) <= b;
    layer0_outputs(166) <= b and not a;
    layer0_outputs(167) <= a or b;
    layer0_outputs(168) <= not b;
    layer0_outputs(169) <= a or b;
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= not a;
    layer0_outputs(172) <= a or b;
    layer0_outputs(173) <= not b;
    layer0_outputs(174) <= a and not b;
    layer0_outputs(175) <= a or b;
    layer0_outputs(176) <= not (a xor b);
    layer0_outputs(177) <= not (a or b);
    layer0_outputs(178) <= a;
    layer0_outputs(179) <= not a or b;
    layer0_outputs(180) <= not a or b;
    layer0_outputs(181) <= b and not a;
    layer0_outputs(182) <= not (a or b);
    layer0_outputs(183) <= not a or b;
    layer0_outputs(184) <= b and not a;
    layer0_outputs(185) <= not a;
    layer0_outputs(186) <= b;
    layer0_outputs(187) <= not b or a;
    layer0_outputs(188) <= a and not b;
    layer0_outputs(189) <= not (a and b);
    layer0_outputs(190) <= '1';
    layer0_outputs(191) <= b and not a;
    layer0_outputs(192) <= not (a xor b);
    layer0_outputs(193) <= not a or b;
    layer0_outputs(194) <= not b;
    layer0_outputs(195) <= b;
    layer0_outputs(196) <= a and not b;
    layer0_outputs(197) <= a;
    layer0_outputs(198) <= not b;
    layer0_outputs(199) <= not b or a;
    layer0_outputs(200) <= not b or a;
    layer0_outputs(201) <= not (a or b);
    layer0_outputs(202) <= not a;
    layer0_outputs(203) <= a and not b;
    layer0_outputs(204) <= a;
    layer0_outputs(205) <= not (a or b);
    layer0_outputs(206) <= not b;
    layer0_outputs(207) <= '1';
    layer0_outputs(208) <= a;
    layer0_outputs(209) <= a or b;
    layer0_outputs(210) <= a;
    layer0_outputs(211) <= a or b;
    layer0_outputs(212) <= '0';
    layer0_outputs(213) <= a or b;
    layer0_outputs(214) <= '0';
    layer0_outputs(215) <= b;
    layer0_outputs(216) <= a;
    layer0_outputs(217) <= not (a or b);
    layer0_outputs(218) <= '1';
    layer0_outputs(219) <= a;
    layer0_outputs(220) <= a or b;
    layer0_outputs(221) <= not b or a;
    layer0_outputs(222) <= not b;
    layer0_outputs(223) <= not a;
    layer0_outputs(224) <= a and not b;
    layer0_outputs(225) <= b;
    layer0_outputs(226) <= not (a or b);
    layer0_outputs(227) <= not a;
    layer0_outputs(228) <= not (a or b);
    layer0_outputs(229) <= not a or b;
    layer0_outputs(230) <= not (a or b);
    layer0_outputs(231) <= a xor b;
    layer0_outputs(232) <= not a or b;
    layer0_outputs(233) <= not b;
    layer0_outputs(234) <= a;
    layer0_outputs(235) <= b;
    layer0_outputs(236) <= a;
    layer0_outputs(237) <= a xor b;
    layer0_outputs(238) <= a or b;
    layer0_outputs(239) <= a or b;
    layer0_outputs(240) <= b and not a;
    layer0_outputs(241) <= not (a and b);
    layer0_outputs(242) <= not a;
    layer0_outputs(243) <= not b;
    layer0_outputs(244) <= '0';
    layer0_outputs(245) <= a and b;
    layer0_outputs(246) <= not a;
    layer0_outputs(247) <= a xor b;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= not (a or b);
    layer0_outputs(250) <= a and not b;
    layer0_outputs(251) <= not (a or b);
    layer0_outputs(252) <= not b;
    layer0_outputs(253) <= not a;
    layer0_outputs(254) <= a and b;
    layer0_outputs(255) <= not b;
    layer0_outputs(256) <= '1';
    layer0_outputs(257) <= not (a and b);
    layer0_outputs(258) <= not b;
    layer0_outputs(259) <= '1';
    layer0_outputs(260) <= not b or a;
    layer0_outputs(261) <= not a or b;
    layer0_outputs(262) <= b and not a;
    layer0_outputs(263) <= not a or b;
    layer0_outputs(264) <= a or b;
    layer0_outputs(265) <= b;
    layer0_outputs(266) <= not (a and b);
    layer0_outputs(267) <= a and not b;
    layer0_outputs(268) <= b;
    layer0_outputs(269) <= a and b;
    layer0_outputs(270) <= a or b;
    layer0_outputs(271) <= '0';
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= b and not a;
    layer0_outputs(274) <= not (a or b);
    layer0_outputs(275) <= not (a or b);
    layer0_outputs(276) <= b and not a;
    layer0_outputs(277) <= not (a or b);
    layer0_outputs(278) <= a or b;
    layer0_outputs(279) <= not (a or b);
    layer0_outputs(280) <= a xor b;
    layer0_outputs(281) <= b;
    layer0_outputs(282) <= b and not a;
    layer0_outputs(283) <= not (a or b);
    layer0_outputs(284) <= not (a and b);
    layer0_outputs(285) <= not a or b;
    layer0_outputs(286) <= a or b;
    layer0_outputs(287) <= not (a or b);
    layer0_outputs(288) <= not a;
    layer0_outputs(289) <= not b;
    layer0_outputs(290) <= b;
    layer0_outputs(291) <= not a;
    layer0_outputs(292) <= b and not a;
    layer0_outputs(293) <= a or b;
    layer0_outputs(294) <= a and not b;
    layer0_outputs(295) <= not (a or b);
    layer0_outputs(296) <= '1';
    layer0_outputs(297) <= a;
    layer0_outputs(298) <= not (a or b);
    layer0_outputs(299) <= b and not a;
    layer0_outputs(300) <= a xor b;
    layer0_outputs(301) <= a or b;
    layer0_outputs(302) <= not b or a;
    layer0_outputs(303) <= not a;
    layer0_outputs(304) <= a xor b;
    layer0_outputs(305) <= not a;
    layer0_outputs(306) <= not (a xor b);
    layer0_outputs(307) <= a and b;
    layer0_outputs(308) <= not a;
    layer0_outputs(309) <= b and not a;
    layer0_outputs(310) <= b and not a;
    layer0_outputs(311) <= not (a or b);
    layer0_outputs(312) <= not b;
    layer0_outputs(313) <= not b;
    layer0_outputs(314) <= b and not a;
    layer0_outputs(315) <= a xor b;
    layer0_outputs(316) <= not b or a;
    layer0_outputs(317) <= b and not a;
    layer0_outputs(318) <= a and not b;
    layer0_outputs(319) <= not b;
    layer0_outputs(320) <= not b;
    layer0_outputs(321) <= '1';
    layer0_outputs(322) <= not (a or b);
    layer0_outputs(323) <= b and not a;
    layer0_outputs(324) <= not a;
    layer0_outputs(325) <= '0';
    layer0_outputs(326) <= a or b;
    layer0_outputs(327) <= b and not a;
    layer0_outputs(328) <= not a or b;
    layer0_outputs(329) <= not a;
    layer0_outputs(330) <= '1';
    layer0_outputs(331) <= '0';
    layer0_outputs(332) <= not b;
    layer0_outputs(333) <= not a;
    layer0_outputs(334) <= not (a xor b);
    layer0_outputs(335) <= not (a xor b);
    layer0_outputs(336) <= a or b;
    layer0_outputs(337) <= not a or b;
    layer0_outputs(338) <= '1';
    layer0_outputs(339) <= '1';
    layer0_outputs(340) <= a;
    layer0_outputs(341) <= '1';
    layer0_outputs(342) <= b;
    layer0_outputs(343) <= a and not b;
    layer0_outputs(344) <= a and b;
    layer0_outputs(345) <= not b;
    layer0_outputs(346) <= not (a or b);
    layer0_outputs(347) <= a and not b;
    layer0_outputs(348) <= not (a or b);
    layer0_outputs(349) <= a and b;
    layer0_outputs(350) <= not b;
    layer0_outputs(351) <= not b or a;
    layer0_outputs(352) <= a or b;
    layer0_outputs(353) <= b;
    layer0_outputs(354) <= a or b;
    layer0_outputs(355) <= not (a xor b);
    layer0_outputs(356) <= not (a xor b);
    layer0_outputs(357) <= b;
    layer0_outputs(358) <= not (a or b);
    layer0_outputs(359) <= a and not b;
    layer0_outputs(360) <= not (a xor b);
    layer0_outputs(361) <= a and b;
    layer0_outputs(362) <= not a;
    layer0_outputs(363) <= a and b;
    layer0_outputs(364) <= '0';
    layer0_outputs(365) <= a xor b;
    layer0_outputs(366) <= a xor b;
    layer0_outputs(367) <= not (a xor b);
    layer0_outputs(368) <= not a or b;
    layer0_outputs(369) <= not (a xor b);
    layer0_outputs(370) <= a;
    layer0_outputs(371) <= not b;
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= not a;
    layer0_outputs(374) <= not (a and b);
    layer0_outputs(375) <= a and b;
    layer0_outputs(376) <= a xor b;
    layer0_outputs(377) <= a or b;
    layer0_outputs(378) <= not a;
    layer0_outputs(379) <= b;
    layer0_outputs(380) <= a or b;
    layer0_outputs(381) <= not a or b;
    layer0_outputs(382) <= not (a xor b);
    layer0_outputs(383) <= '0';
    layer0_outputs(384) <= not b;
    layer0_outputs(385) <= not b or a;
    layer0_outputs(386) <= not a;
    layer0_outputs(387) <= not (a xor b);
    layer0_outputs(388) <= not a;
    layer0_outputs(389) <= a;
    layer0_outputs(390) <= not (a xor b);
    layer0_outputs(391) <= '1';
    layer0_outputs(392) <= a;
    layer0_outputs(393) <= not (a and b);
    layer0_outputs(394) <= not b;
    layer0_outputs(395) <= '1';
    layer0_outputs(396) <= not b or a;
    layer0_outputs(397) <= not b or a;
    layer0_outputs(398) <= not b;
    layer0_outputs(399) <= not (a or b);
    layer0_outputs(400) <= b;
    layer0_outputs(401) <= b;
    layer0_outputs(402) <= a;
    layer0_outputs(403) <= a;
    layer0_outputs(404) <= not b;
    layer0_outputs(405) <= a or b;
    layer0_outputs(406) <= a;
    layer0_outputs(407) <= a and not b;
    layer0_outputs(408) <= '1';
    layer0_outputs(409) <= not (a or b);
    layer0_outputs(410) <= not (a or b);
    layer0_outputs(411) <= not (a or b);
    layer0_outputs(412) <= not a or b;
    layer0_outputs(413) <= '0';
    layer0_outputs(414) <= '1';
    layer0_outputs(415) <= '0';
    layer0_outputs(416) <= a or b;
    layer0_outputs(417) <= not b;
    layer0_outputs(418) <= b and not a;
    layer0_outputs(419) <= not b or a;
    layer0_outputs(420) <= a;
    layer0_outputs(421) <= a or b;
    layer0_outputs(422) <= not a or b;
    layer0_outputs(423) <= '1';
    layer0_outputs(424) <= not b;
    layer0_outputs(425) <= b;
    layer0_outputs(426) <= not b or a;
    layer0_outputs(427) <= not (a xor b);
    layer0_outputs(428) <= not b or a;
    layer0_outputs(429) <= not a or b;
    layer0_outputs(430) <= '1';
    layer0_outputs(431) <= not b or a;
    layer0_outputs(432) <= b and not a;
    layer0_outputs(433) <= b;
    layer0_outputs(434) <= b;
    layer0_outputs(435) <= a;
    layer0_outputs(436) <= not b;
    layer0_outputs(437) <= a and b;
    layer0_outputs(438) <= a or b;
    layer0_outputs(439) <= not b or a;
    layer0_outputs(440) <= not b or a;
    layer0_outputs(441) <= a and not b;
    layer0_outputs(442) <= b and not a;
    layer0_outputs(443) <= a or b;
    layer0_outputs(444) <= a or b;
    layer0_outputs(445) <= a;
    layer0_outputs(446) <= a and not b;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= not a;
    layer0_outputs(449) <= not b or a;
    layer0_outputs(450) <= a;
    layer0_outputs(451) <= not b;
    layer0_outputs(452) <= a xor b;
    layer0_outputs(453) <= not (a or b);
    layer0_outputs(454) <= b and not a;
    layer0_outputs(455) <= a;
    layer0_outputs(456) <= not (a or b);
    layer0_outputs(457) <= '1';
    layer0_outputs(458) <= a and not b;
    layer0_outputs(459) <= a or b;
    layer0_outputs(460) <= a or b;
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= b and not a;
    layer0_outputs(463) <= not (a and b);
    layer0_outputs(464) <= not a or b;
    layer0_outputs(465) <= b and not a;
    layer0_outputs(466) <= not a;
    layer0_outputs(467) <= b and not a;
    layer0_outputs(468) <= a or b;
    layer0_outputs(469) <= a and not b;
    layer0_outputs(470) <= b and not a;
    layer0_outputs(471) <= not a;
    layer0_outputs(472) <= not (a xor b);
    layer0_outputs(473) <= a xor b;
    layer0_outputs(474) <= b and not a;
    layer0_outputs(475) <= not b or a;
    layer0_outputs(476) <= not a;
    layer0_outputs(477) <= not (a or b);
    layer0_outputs(478) <= a;
    layer0_outputs(479) <= a and b;
    layer0_outputs(480) <= not (a and b);
    layer0_outputs(481) <= not b or a;
    layer0_outputs(482) <= a and b;
    layer0_outputs(483) <= not b;
    layer0_outputs(484) <= not (a xor b);
    layer0_outputs(485) <= not (a xor b);
    layer0_outputs(486) <= a or b;
    layer0_outputs(487) <= not a;
    layer0_outputs(488) <= not a;
    layer0_outputs(489) <= a;
    layer0_outputs(490) <= a or b;
    layer0_outputs(491) <= a and not b;
    layer0_outputs(492) <= not b;
    layer0_outputs(493) <= a xor b;
    layer0_outputs(494) <= a and not b;
    layer0_outputs(495) <= a;
    layer0_outputs(496) <= b;
    layer0_outputs(497) <= not b;
    layer0_outputs(498) <= b and not a;
    layer0_outputs(499) <= not b;
    layer0_outputs(500) <= b;
    layer0_outputs(501) <= a and b;
    layer0_outputs(502) <= not b;
    layer0_outputs(503) <= b;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= a or b;
    layer0_outputs(506) <= not a;
    layer0_outputs(507) <= not (a and b);
    layer0_outputs(508) <= b and not a;
    layer0_outputs(509) <= not b;
    layer0_outputs(510) <= not (a and b);
    layer0_outputs(511) <= not (a and b);
    layer0_outputs(512) <= b;
    layer0_outputs(513) <= b;
    layer0_outputs(514) <= a;
    layer0_outputs(515) <= a or b;
    layer0_outputs(516) <= not (a or b);
    layer0_outputs(517) <= a and not b;
    layer0_outputs(518) <= '0';
    layer0_outputs(519) <= b;
    layer0_outputs(520) <= not b;
    layer0_outputs(521) <= a xor b;
    layer0_outputs(522) <= not (a and b);
    layer0_outputs(523) <= '1';
    layer0_outputs(524) <= b;
    layer0_outputs(525) <= a xor b;
    layer0_outputs(526) <= '0';
    layer0_outputs(527) <= '0';
    layer0_outputs(528) <= a;
    layer0_outputs(529) <= not b or a;
    layer0_outputs(530) <= not (a and b);
    layer0_outputs(531) <= a and not b;
    layer0_outputs(532) <= b;
    layer0_outputs(533) <= a;
    layer0_outputs(534) <= b;
    layer0_outputs(535) <= not (a or b);
    layer0_outputs(536) <= b;
    layer0_outputs(537) <= not (a or b);
    layer0_outputs(538) <= a or b;
    layer0_outputs(539) <= not (a xor b);
    layer0_outputs(540) <= '1';
    layer0_outputs(541) <= '0';
    layer0_outputs(542) <= not a or b;
    layer0_outputs(543) <= b;
    layer0_outputs(544) <= a;
    layer0_outputs(545) <= a and not b;
    layer0_outputs(546) <= not b or a;
    layer0_outputs(547) <= a;
    layer0_outputs(548) <= a xor b;
    layer0_outputs(549) <= not a;
    layer0_outputs(550) <= not b;
    layer0_outputs(551) <= not a or b;
    layer0_outputs(552) <= not a;
    layer0_outputs(553) <= a and not b;
    layer0_outputs(554) <= a and not b;
    layer0_outputs(555) <= not b or a;
    layer0_outputs(556) <= not (a or b);
    layer0_outputs(557) <= not (a or b);
    layer0_outputs(558) <= not (a and b);
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= a;
    layer0_outputs(561) <= not (a or b);
    layer0_outputs(562) <= not (a xor b);
    layer0_outputs(563) <= b and not a;
    layer0_outputs(564) <= not (a xor b);
    layer0_outputs(565) <= a and b;
    layer0_outputs(566) <= a or b;
    layer0_outputs(567) <= not (a xor b);
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= a and not b;
    layer0_outputs(570) <= a and not b;
    layer0_outputs(571) <= '1';
    layer0_outputs(572) <= not (a xor b);
    layer0_outputs(573) <= a and not b;
    layer0_outputs(574) <= a xor b;
    layer0_outputs(575) <= a or b;
    layer0_outputs(576) <= a;
    layer0_outputs(577) <= '0';
    layer0_outputs(578) <= not b;
    layer0_outputs(579) <= a;
    layer0_outputs(580) <= a or b;
    layer0_outputs(581) <= b;
    layer0_outputs(582) <= not b or a;
    layer0_outputs(583) <= not b or a;
    layer0_outputs(584) <= not (a or b);
    layer0_outputs(585) <= b and not a;
    layer0_outputs(586) <= not b or a;
    layer0_outputs(587) <= a and not b;
    layer0_outputs(588) <= not (a and b);
    layer0_outputs(589) <= a and not b;
    layer0_outputs(590) <= not a;
    layer0_outputs(591) <= not b or a;
    layer0_outputs(592) <= a or b;
    layer0_outputs(593) <= '1';
    layer0_outputs(594) <= not b;
    layer0_outputs(595) <= a xor b;
    layer0_outputs(596) <= not a or b;
    layer0_outputs(597) <= a and not b;
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= a or b;
    layer0_outputs(600) <= not b or a;
    layer0_outputs(601) <= not b;
    layer0_outputs(602) <= a or b;
    layer0_outputs(603) <= not (a or b);
    layer0_outputs(604) <= not a or b;
    layer0_outputs(605) <= not b;
    layer0_outputs(606) <= '1';
    layer0_outputs(607) <= b and not a;
    layer0_outputs(608) <= a and b;
    layer0_outputs(609) <= not (a and b);
    layer0_outputs(610) <= b and not a;
    layer0_outputs(611) <= a;
    layer0_outputs(612) <= '1';
    layer0_outputs(613) <= not b;
    layer0_outputs(614) <= not b;
    layer0_outputs(615) <= a;
    layer0_outputs(616) <= a or b;
    layer0_outputs(617) <= a and b;
    layer0_outputs(618) <= not b or a;
    layer0_outputs(619) <= not b;
    layer0_outputs(620) <= not (a or b);
    layer0_outputs(621) <= a and not b;
    layer0_outputs(622) <= a and not b;
    layer0_outputs(623) <= a and not b;
    layer0_outputs(624) <= not a or b;
    layer0_outputs(625) <= not (a xor b);
    layer0_outputs(626) <= not (a xor b);
    layer0_outputs(627) <= '0';
    layer0_outputs(628) <= not (a xor b);
    layer0_outputs(629) <= a or b;
    layer0_outputs(630) <= a;
    layer0_outputs(631) <= '1';
    layer0_outputs(632) <= '0';
    layer0_outputs(633) <= not b or a;
    layer0_outputs(634) <= a or b;
    layer0_outputs(635) <= '0';
    layer0_outputs(636) <= a or b;
    layer0_outputs(637) <= b and not a;
    layer0_outputs(638) <= not b or a;
    layer0_outputs(639) <= not b or a;
    layer0_outputs(640) <= '1';
    layer0_outputs(641) <= a;
    layer0_outputs(642) <= not (a xor b);
    layer0_outputs(643) <= a xor b;
    layer0_outputs(644) <= not b or a;
    layer0_outputs(645) <= b;
    layer0_outputs(646) <= not (a xor b);
    layer0_outputs(647) <= b;
    layer0_outputs(648) <= a or b;
    layer0_outputs(649) <= b;
    layer0_outputs(650) <= not (a xor b);
    layer0_outputs(651) <= a and b;
    layer0_outputs(652) <= b;
    layer0_outputs(653) <= not a;
    layer0_outputs(654) <= not a;
    layer0_outputs(655) <= a and not b;
    layer0_outputs(656) <= '1';
    layer0_outputs(657) <= b and not a;
    layer0_outputs(658) <= not (a xor b);
    layer0_outputs(659) <= not (a or b);
    layer0_outputs(660) <= b;
    layer0_outputs(661) <= not b;
    layer0_outputs(662) <= not b;
    layer0_outputs(663) <= a xor b;
    layer0_outputs(664) <= b;
    layer0_outputs(665) <= not a;
    layer0_outputs(666) <= a or b;
    layer0_outputs(667) <= b and not a;
    layer0_outputs(668) <= a;
    layer0_outputs(669) <= a xor b;
    layer0_outputs(670) <= '1';
    layer0_outputs(671) <= not a or b;
    layer0_outputs(672) <= b;
    layer0_outputs(673) <= not (a or b);
    layer0_outputs(674) <= not (a and b);
    layer0_outputs(675) <= not a;
    layer0_outputs(676) <= not b or a;
    layer0_outputs(677) <= b and not a;
    layer0_outputs(678) <= not (a or b);
    layer0_outputs(679) <= not a;
    layer0_outputs(680) <= b and not a;
    layer0_outputs(681) <= b;
    layer0_outputs(682) <= b;
    layer0_outputs(683) <= a or b;
    layer0_outputs(684) <= not (a or b);
    layer0_outputs(685) <= a xor b;
    layer0_outputs(686) <= a xor b;
    layer0_outputs(687) <= not b;
    layer0_outputs(688) <= b and not a;
    layer0_outputs(689) <= b and not a;
    layer0_outputs(690) <= not (a or b);
    layer0_outputs(691) <= not a or b;
    layer0_outputs(692) <= not (a or b);
    layer0_outputs(693) <= not a;
    layer0_outputs(694) <= a or b;
    layer0_outputs(695) <= not a or b;
    layer0_outputs(696) <= not (a or b);
    layer0_outputs(697) <= not b;
    layer0_outputs(698) <= not a;
    layer0_outputs(699) <= b and not a;
    layer0_outputs(700) <= not (a xor b);
    layer0_outputs(701) <= a or b;
    layer0_outputs(702) <= b;
    layer0_outputs(703) <= a xor b;
    layer0_outputs(704) <= a and b;
    layer0_outputs(705) <= b;
    layer0_outputs(706) <= not a;
    layer0_outputs(707) <= a xor b;
    layer0_outputs(708) <= not a;
    layer0_outputs(709) <= b;
    layer0_outputs(710) <= a and b;
    layer0_outputs(711) <= a;
    layer0_outputs(712) <= a and not b;
    layer0_outputs(713) <= '1';
    layer0_outputs(714) <= not b;
    layer0_outputs(715) <= not b;
    layer0_outputs(716) <= b;
    layer0_outputs(717) <= a xor b;
    layer0_outputs(718) <= not b or a;
    layer0_outputs(719) <= not (a or b);
    layer0_outputs(720) <= not (a or b);
    layer0_outputs(721) <= '0';
    layer0_outputs(722) <= '0';
    layer0_outputs(723) <= a and b;
    layer0_outputs(724) <= a or b;
    layer0_outputs(725) <= '1';
    layer0_outputs(726) <= not b or a;
    layer0_outputs(727) <= not a or b;
    layer0_outputs(728) <= a and not b;
    layer0_outputs(729) <= a or b;
    layer0_outputs(730) <= a xor b;
    layer0_outputs(731) <= not (a or b);
    layer0_outputs(732) <= b and not a;
    layer0_outputs(733) <= a or b;
    layer0_outputs(734) <= a and not b;
    layer0_outputs(735) <= not b;
    layer0_outputs(736) <= not (a xor b);
    layer0_outputs(737) <= not b or a;
    layer0_outputs(738) <= b and not a;
    layer0_outputs(739) <= not a;
    layer0_outputs(740) <= not (a or b);
    layer0_outputs(741) <= not a;
    layer0_outputs(742) <= '1';
    layer0_outputs(743) <= not b or a;
    layer0_outputs(744) <= b;
    layer0_outputs(745) <= a or b;
    layer0_outputs(746) <= a or b;
    layer0_outputs(747) <= a and b;
    layer0_outputs(748) <= not (a or b);
    layer0_outputs(749) <= a xor b;
    layer0_outputs(750) <= b and not a;
    layer0_outputs(751) <= b and not a;
    layer0_outputs(752) <= not a or b;
    layer0_outputs(753) <= a or b;
    layer0_outputs(754) <= b;
    layer0_outputs(755) <= b;
    layer0_outputs(756) <= a or b;
    layer0_outputs(757) <= not a or b;
    layer0_outputs(758) <= a or b;
    layer0_outputs(759) <= b;
    layer0_outputs(760) <= not b or a;
    layer0_outputs(761) <= not (a or b);
    layer0_outputs(762) <= a and not b;
    layer0_outputs(763) <= a;
    layer0_outputs(764) <= not (a or b);
    layer0_outputs(765) <= b;
    layer0_outputs(766) <= '1';
    layer0_outputs(767) <= b and not a;
    layer0_outputs(768) <= '1';
    layer0_outputs(769) <= a xor b;
    layer0_outputs(770) <= not a;
    layer0_outputs(771) <= a and b;
    layer0_outputs(772) <= not (a or b);
    layer0_outputs(773) <= a or b;
    layer0_outputs(774) <= a and not b;
    layer0_outputs(775) <= not a or b;
    layer0_outputs(776) <= not b;
    layer0_outputs(777) <= not (a or b);
    layer0_outputs(778) <= b and not a;
    layer0_outputs(779) <= not b or a;
    layer0_outputs(780) <= b;
    layer0_outputs(781) <= not (a xor b);
    layer0_outputs(782) <= not b;
    layer0_outputs(783) <= not b;
    layer0_outputs(784) <= a and not b;
    layer0_outputs(785) <= not (a or b);
    layer0_outputs(786) <= not a or b;
    layer0_outputs(787) <= not b;
    layer0_outputs(788) <= a;
    layer0_outputs(789) <= not a;
    layer0_outputs(790) <= not (a or b);
    layer0_outputs(791) <= '1';
    layer0_outputs(792) <= not (a xor b);
    layer0_outputs(793) <= not b;
    layer0_outputs(794) <= a or b;
    layer0_outputs(795) <= a xor b;
    layer0_outputs(796) <= not (a or b);
    layer0_outputs(797) <= b;
    layer0_outputs(798) <= not a;
    layer0_outputs(799) <= not a or b;
    layer0_outputs(800) <= b;
    layer0_outputs(801) <= a and b;
    layer0_outputs(802) <= a;
    layer0_outputs(803) <= not (a or b);
    layer0_outputs(804) <= a;
    layer0_outputs(805) <= a xor b;
    layer0_outputs(806) <= a or b;
    layer0_outputs(807) <= a or b;
    layer0_outputs(808) <= a and not b;
    layer0_outputs(809) <= not (a or b);
    layer0_outputs(810) <= a or b;
    layer0_outputs(811) <= a;
    layer0_outputs(812) <= not b;
    layer0_outputs(813) <= a and not b;
    layer0_outputs(814) <= a or b;
    layer0_outputs(815) <= not a;
    layer0_outputs(816) <= '1';
    layer0_outputs(817) <= '0';
    layer0_outputs(818) <= not (a xor b);
    layer0_outputs(819) <= not a;
    layer0_outputs(820) <= not (a or b);
    layer0_outputs(821) <= not (a xor b);
    layer0_outputs(822) <= not a or b;
    layer0_outputs(823) <= a or b;
    layer0_outputs(824) <= a;
    layer0_outputs(825) <= b;
    layer0_outputs(826) <= '0';
    layer0_outputs(827) <= a xor b;
    layer0_outputs(828) <= b;
    layer0_outputs(829) <= a or b;
    layer0_outputs(830) <= a and not b;
    layer0_outputs(831) <= not a;
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= b;
    layer0_outputs(834) <= not a or b;
    layer0_outputs(835) <= a or b;
    layer0_outputs(836) <= a and not b;
    layer0_outputs(837) <= not (a or b);
    layer0_outputs(838) <= a or b;
    layer0_outputs(839) <= not (a or b);
    layer0_outputs(840) <= not b;
    layer0_outputs(841) <= '1';
    layer0_outputs(842) <= a xor b;
    layer0_outputs(843) <= not (a and b);
    layer0_outputs(844) <= a;
    layer0_outputs(845) <= a or b;
    layer0_outputs(846) <= a or b;
    layer0_outputs(847) <= b and not a;
    layer0_outputs(848) <= not (a and b);
    layer0_outputs(849) <= not (a or b);
    layer0_outputs(850) <= not a;
    layer0_outputs(851) <= b;
    layer0_outputs(852) <= not b;
    layer0_outputs(853) <= not a or b;
    layer0_outputs(854) <= b and not a;
    layer0_outputs(855) <= '1';
    layer0_outputs(856) <= b and not a;
    layer0_outputs(857) <= not (a xor b);
    layer0_outputs(858) <= a or b;
    layer0_outputs(859) <= b;
    layer0_outputs(860) <= b;
    layer0_outputs(861) <= a and not b;
    layer0_outputs(862) <= b;
    layer0_outputs(863) <= a xor b;
    layer0_outputs(864) <= a and not b;
    layer0_outputs(865) <= not b;
    layer0_outputs(866) <= not a or b;
    layer0_outputs(867) <= a and not b;
    layer0_outputs(868) <= not b;
    layer0_outputs(869) <= '0';
    layer0_outputs(870) <= not (a or b);
    layer0_outputs(871) <= not b or a;
    layer0_outputs(872) <= '0';
    layer0_outputs(873) <= not (a or b);
    layer0_outputs(874) <= not (a xor b);
    layer0_outputs(875) <= a or b;
    layer0_outputs(876) <= b;
    layer0_outputs(877) <= not (a and b);
    layer0_outputs(878) <= not (a and b);
    layer0_outputs(879) <= '1';
    layer0_outputs(880) <= a;
    layer0_outputs(881) <= a and b;
    layer0_outputs(882) <= a or b;
    layer0_outputs(883) <= not b or a;
    layer0_outputs(884) <= not (a xor b);
    layer0_outputs(885) <= not (a or b);
    layer0_outputs(886) <= not (a or b);
    layer0_outputs(887) <= not b or a;
    layer0_outputs(888) <= not b or a;
    layer0_outputs(889) <= b and not a;
    layer0_outputs(890) <= not (a or b);
    layer0_outputs(891) <= not b;
    layer0_outputs(892) <= a or b;
    layer0_outputs(893) <= b and not a;
    layer0_outputs(894) <= not b or a;
    layer0_outputs(895) <= '1';
    layer0_outputs(896) <= not b;
    layer0_outputs(897) <= not (a or b);
    layer0_outputs(898) <= a and not b;
    layer0_outputs(899) <= b and not a;
    layer0_outputs(900) <= a and not b;
    layer0_outputs(901) <= not b;
    layer0_outputs(902) <= a;
    layer0_outputs(903) <= not (a or b);
    layer0_outputs(904) <= a;
    layer0_outputs(905) <= not a;
    layer0_outputs(906) <= b and not a;
    layer0_outputs(907) <= not (a or b);
    layer0_outputs(908) <= not (a or b);
    layer0_outputs(909) <= not (a or b);
    layer0_outputs(910) <= not a;
    layer0_outputs(911) <= a;
    layer0_outputs(912) <= not b or a;
    layer0_outputs(913) <= not (a or b);
    layer0_outputs(914) <= a or b;
    layer0_outputs(915) <= b;
    layer0_outputs(916) <= b and not a;
    layer0_outputs(917) <= not (a or b);
    layer0_outputs(918) <= not (a or b);
    layer0_outputs(919) <= not b;
    layer0_outputs(920) <= not (a xor b);
    layer0_outputs(921) <= not (a or b);
    layer0_outputs(922) <= not a;
    layer0_outputs(923) <= not b;
    layer0_outputs(924) <= not a or b;
    layer0_outputs(925) <= not (a or b);
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= b and not a;
    layer0_outputs(928) <= a and b;
    layer0_outputs(929) <= not (a or b);
    layer0_outputs(930) <= not (a xor b);
    layer0_outputs(931) <= not a or b;
    layer0_outputs(932) <= not a or b;
    layer0_outputs(933) <= a or b;
    layer0_outputs(934) <= b;
    layer0_outputs(935) <= a;
    layer0_outputs(936) <= not (a and b);
    layer0_outputs(937) <= not b or a;
    layer0_outputs(938) <= b;
    layer0_outputs(939) <= a;
    layer0_outputs(940) <= b;
    layer0_outputs(941) <= not b;
    layer0_outputs(942) <= not (a or b);
    layer0_outputs(943) <= not (a and b);
    layer0_outputs(944) <= not b or a;
    layer0_outputs(945) <= a and not b;
    layer0_outputs(946) <= not (a or b);
    layer0_outputs(947) <= not (a or b);
    layer0_outputs(948) <= not a;
    layer0_outputs(949) <= a;
    layer0_outputs(950) <= '0';
    layer0_outputs(951) <= a xor b;
    layer0_outputs(952) <= '1';
    layer0_outputs(953) <= '1';
    layer0_outputs(954) <= '1';
    layer0_outputs(955) <= b and not a;
    layer0_outputs(956) <= not a or b;
    layer0_outputs(957) <= not b;
    layer0_outputs(958) <= not (a xor b);
    layer0_outputs(959) <= b and not a;
    layer0_outputs(960) <= not b or a;
    layer0_outputs(961) <= a xor b;
    layer0_outputs(962) <= '0';
    layer0_outputs(963) <= not (a or b);
    layer0_outputs(964) <= a xor b;
    layer0_outputs(965) <= a;
    layer0_outputs(966) <= not (a xor b);
    layer0_outputs(967) <= not a or b;
    layer0_outputs(968) <= a or b;
    layer0_outputs(969) <= a xor b;
    layer0_outputs(970) <= not b or a;
    layer0_outputs(971) <= a and b;
    layer0_outputs(972) <= b and not a;
    layer0_outputs(973) <= b;
    layer0_outputs(974) <= b and not a;
    layer0_outputs(975) <= not (a or b);
    layer0_outputs(976) <= a xor b;
    layer0_outputs(977) <= a and b;
    layer0_outputs(978) <= '1';
    layer0_outputs(979) <= a and b;
    layer0_outputs(980) <= not b;
    layer0_outputs(981) <= not b;
    layer0_outputs(982) <= not a;
    layer0_outputs(983) <= not a;
    layer0_outputs(984) <= not (a or b);
    layer0_outputs(985) <= b;
    layer0_outputs(986) <= not (a xor b);
    layer0_outputs(987) <= a or b;
    layer0_outputs(988) <= a and b;
    layer0_outputs(989) <= not (a or b);
    layer0_outputs(990) <= not (a and b);
    layer0_outputs(991) <= '0';
    layer0_outputs(992) <= not b;
    layer0_outputs(993) <= a xor b;
    layer0_outputs(994) <= a or b;
    layer0_outputs(995) <= a and b;
    layer0_outputs(996) <= not a;
    layer0_outputs(997) <= a or b;
    layer0_outputs(998) <= b and not a;
    layer0_outputs(999) <= not (a or b);
    layer0_outputs(1000) <= not b;
    layer0_outputs(1001) <= not a;
    layer0_outputs(1002) <= a xor b;
    layer0_outputs(1003) <= a or b;
    layer0_outputs(1004) <= not (a or b);
    layer0_outputs(1005) <= not b;
    layer0_outputs(1006) <= '1';
    layer0_outputs(1007) <= not b or a;
    layer0_outputs(1008) <= b;
    layer0_outputs(1009) <= '1';
    layer0_outputs(1010) <= a or b;
    layer0_outputs(1011) <= a and b;
    layer0_outputs(1012) <= b;
    layer0_outputs(1013) <= b and not a;
    layer0_outputs(1014) <= a or b;
    layer0_outputs(1015) <= not a;
    layer0_outputs(1016) <= '0';
    layer0_outputs(1017) <= a or b;
    layer0_outputs(1018) <= '1';
    layer0_outputs(1019) <= '1';
    layer0_outputs(1020) <= not b or a;
    layer0_outputs(1021) <= not a;
    layer0_outputs(1022) <= a xor b;
    layer0_outputs(1023) <= a and not b;
    layer0_outputs(1024) <= not a;
    layer0_outputs(1025) <= not a;
    layer0_outputs(1026) <= not (a or b);
    layer0_outputs(1027) <= not (a or b);
    layer0_outputs(1028) <= not (a or b);
    layer0_outputs(1029) <= b and not a;
    layer0_outputs(1030) <= a;
    layer0_outputs(1031) <= a or b;
    layer0_outputs(1032) <= not a;
    layer0_outputs(1033) <= not (a or b);
    layer0_outputs(1034) <= not b;
    layer0_outputs(1035) <= a xor b;
    layer0_outputs(1036) <= not (a and b);
    layer0_outputs(1037) <= not a or b;
    layer0_outputs(1038) <= not (a or b);
    layer0_outputs(1039) <= a and b;
    layer0_outputs(1040) <= a or b;
    layer0_outputs(1041) <= a;
    layer0_outputs(1042) <= not b or a;
    layer0_outputs(1043) <= not a;
    layer0_outputs(1044) <= not b or a;
    layer0_outputs(1045) <= a or b;
    layer0_outputs(1046) <= a xor b;
    layer0_outputs(1047) <= '1';
    layer0_outputs(1048) <= not a or b;
    layer0_outputs(1049) <= '0';
    layer0_outputs(1050) <= a and not b;
    layer0_outputs(1051) <= a and not b;
    layer0_outputs(1052) <= a or b;
    layer0_outputs(1053) <= a;
    layer0_outputs(1054) <= not a;
    layer0_outputs(1055) <= b and not a;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= not a;
    layer0_outputs(1058) <= not (a or b);
    layer0_outputs(1059) <= a xor b;
    layer0_outputs(1060) <= not b or a;
    layer0_outputs(1061) <= not (a or b);
    layer0_outputs(1062) <= a xor b;
    layer0_outputs(1063) <= a and not b;
    layer0_outputs(1064) <= not (a or b);
    layer0_outputs(1065) <= not a;
    layer0_outputs(1066) <= not b;
    layer0_outputs(1067) <= not a;
    layer0_outputs(1068) <= b;
    layer0_outputs(1069) <= '0';
    layer0_outputs(1070) <= not b;
    layer0_outputs(1071) <= b and not a;
    layer0_outputs(1072) <= a;
    layer0_outputs(1073) <= not (a or b);
    layer0_outputs(1074) <= not (a and b);
    layer0_outputs(1075) <= not b or a;
    layer0_outputs(1076) <= not a or b;
    layer0_outputs(1077) <= not a or b;
    layer0_outputs(1078) <= not (a xor b);
    layer0_outputs(1079) <= a xor b;
    layer0_outputs(1080) <= a and b;
    layer0_outputs(1081) <= '1';
    layer0_outputs(1082) <= a and b;
    layer0_outputs(1083) <= a and b;
    layer0_outputs(1084) <= a or b;
    layer0_outputs(1085) <= not (a or b);
    layer0_outputs(1086) <= not b;
    layer0_outputs(1087) <= not b;
    layer0_outputs(1088) <= not a;
    layer0_outputs(1089) <= not b;
    layer0_outputs(1090) <= '0';
    layer0_outputs(1091) <= b and not a;
    layer0_outputs(1092) <= not (a or b);
    layer0_outputs(1093) <= b;
    layer0_outputs(1094) <= a or b;
    layer0_outputs(1095) <= a or b;
    layer0_outputs(1096) <= not a;
    layer0_outputs(1097) <= b and not a;
    layer0_outputs(1098) <= not (a or b);
    layer0_outputs(1099) <= '0';
    layer0_outputs(1100) <= a xor b;
    layer0_outputs(1101) <= not (a or b);
    layer0_outputs(1102) <= not (a or b);
    layer0_outputs(1103) <= not b;
    layer0_outputs(1104) <= not (a or b);
    layer0_outputs(1105) <= not b;
    layer0_outputs(1106) <= not b;
    layer0_outputs(1107) <= not (a or b);
    layer0_outputs(1108) <= not (a xor b);
    layer0_outputs(1109) <= a or b;
    layer0_outputs(1110) <= b;
    layer0_outputs(1111) <= a or b;
    layer0_outputs(1112) <= not (a or b);
    layer0_outputs(1113) <= a;
    layer0_outputs(1114) <= a and not b;
    layer0_outputs(1115) <= not (a xor b);
    layer0_outputs(1116) <= not a or b;
    layer0_outputs(1117) <= a;
    layer0_outputs(1118) <= not a;
    layer0_outputs(1119) <= a or b;
    layer0_outputs(1120) <= not b;
    layer0_outputs(1121) <= a or b;
    layer0_outputs(1122) <= not (a xor b);
    layer0_outputs(1123) <= not b or a;
    layer0_outputs(1124) <= '1';
    layer0_outputs(1125) <= not b;
    layer0_outputs(1126) <= a xor b;
    layer0_outputs(1127) <= not a or b;
    layer0_outputs(1128) <= a and not b;
    layer0_outputs(1129) <= a or b;
    layer0_outputs(1130) <= not (a or b);
    layer0_outputs(1131) <= not b or a;
    layer0_outputs(1132) <= not a or b;
    layer0_outputs(1133) <= b and not a;
    layer0_outputs(1134) <= not a;
    layer0_outputs(1135) <= a and not b;
    layer0_outputs(1136) <= a;
    layer0_outputs(1137) <= not b or a;
    layer0_outputs(1138) <= not a;
    layer0_outputs(1139) <= '1';
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= '1';
    layer0_outputs(1142) <= b;
    layer0_outputs(1143) <= a xor b;
    layer0_outputs(1144) <= a;
    layer0_outputs(1145) <= not (a and b);
    layer0_outputs(1146) <= not a;
    layer0_outputs(1147) <= a or b;
    layer0_outputs(1148) <= not (a or b);
    layer0_outputs(1149) <= a;
    layer0_outputs(1150) <= a or b;
    layer0_outputs(1151) <= a and b;
    layer0_outputs(1152) <= not a or b;
    layer0_outputs(1153) <= '0';
    layer0_outputs(1154) <= a xor b;
    layer0_outputs(1155) <= '1';
    layer0_outputs(1156) <= b and not a;
    layer0_outputs(1157) <= not b or a;
    layer0_outputs(1158) <= not b or a;
    layer0_outputs(1159) <= not a;
    layer0_outputs(1160) <= a and not b;
    layer0_outputs(1161) <= a;
    layer0_outputs(1162) <= a and not b;
    layer0_outputs(1163) <= a or b;
    layer0_outputs(1164) <= b;
    layer0_outputs(1165) <= not (a and b);
    layer0_outputs(1166) <= '0';
    layer0_outputs(1167) <= a or b;
    layer0_outputs(1168) <= a or b;
    layer0_outputs(1169) <= b;
    layer0_outputs(1170) <= '1';
    layer0_outputs(1171) <= a and not b;
    layer0_outputs(1172) <= not b;
    layer0_outputs(1173) <= '0';
    layer0_outputs(1174) <= a or b;
    layer0_outputs(1175) <= a xor b;
    layer0_outputs(1176) <= not (a or b);
    layer0_outputs(1177) <= not (a or b);
    layer0_outputs(1178) <= a and not b;
    layer0_outputs(1179) <= a;
    layer0_outputs(1180) <= b;
    layer0_outputs(1181) <= not (a or b);
    layer0_outputs(1182) <= not (a or b);
    layer0_outputs(1183) <= '1';
    layer0_outputs(1184) <= not a or b;
    layer0_outputs(1185) <= not (a or b);
    layer0_outputs(1186) <= a or b;
    layer0_outputs(1187) <= not a or b;
    layer0_outputs(1188) <= not (a or b);
    layer0_outputs(1189) <= not (a or b);
    layer0_outputs(1190) <= not a;
    layer0_outputs(1191) <= '0';
    layer0_outputs(1192) <= b;
    layer0_outputs(1193) <= not a or b;
    layer0_outputs(1194) <= not a or b;
    layer0_outputs(1195) <= a or b;
    layer0_outputs(1196) <= not (a xor b);
    layer0_outputs(1197) <= not b;
    layer0_outputs(1198) <= not b;
    layer0_outputs(1199) <= b and not a;
    layer0_outputs(1200) <= not a or b;
    layer0_outputs(1201) <= a or b;
    layer0_outputs(1202) <= not (a or b);
    layer0_outputs(1203) <= not (a or b);
    layer0_outputs(1204) <= b;
    layer0_outputs(1205) <= not a or b;
    layer0_outputs(1206) <= a xor b;
    layer0_outputs(1207) <= '0';
    layer0_outputs(1208) <= not a;
    layer0_outputs(1209) <= not b;
    layer0_outputs(1210) <= not (a and b);
    layer0_outputs(1211) <= a and b;
    layer0_outputs(1212) <= '0';
    layer0_outputs(1213) <= a xor b;
    layer0_outputs(1214) <= a;
    layer0_outputs(1215) <= not a;
    layer0_outputs(1216) <= not (a xor b);
    layer0_outputs(1217) <= a;
    layer0_outputs(1218) <= not a or b;
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= a and b;
    layer0_outputs(1221) <= not a or b;
    layer0_outputs(1222) <= a;
    layer0_outputs(1223) <= not b;
    layer0_outputs(1224) <= a or b;
    layer0_outputs(1225) <= b and not a;
    layer0_outputs(1226) <= a or b;
    layer0_outputs(1227) <= a and b;
    layer0_outputs(1228) <= not b;
    layer0_outputs(1229) <= b and not a;
    layer0_outputs(1230) <= not a;
    layer0_outputs(1231) <= not a;
    layer0_outputs(1232) <= not (a and b);
    layer0_outputs(1233) <= a xor b;
    layer0_outputs(1234) <= not (a xor b);
    layer0_outputs(1235) <= a and not b;
    layer0_outputs(1236) <= b;
    layer0_outputs(1237) <= not b or a;
    layer0_outputs(1238) <= not b or a;
    layer0_outputs(1239) <= a;
    layer0_outputs(1240) <= b;
    layer0_outputs(1241) <= a and not b;
    layer0_outputs(1242) <= not b or a;
    layer0_outputs(1243) <= not b or a;
    layer0_outputs(1244) <= not b or a;
    layer0_outputs(1245) <= '0';
    layer0_outputs(1246) <= not (a and b);
    layer0_outputs(1247) <= a;
    layer0_outputs(1248) <= not b;
    layer0_outputs(1249) <= b and not a;
    layer0_outputs(1250) <= not b or a;
    layer0_outputs(1251) <= not a;
    layer0_outputs(1252) <= not a;
    layer0_outputs(1253) <= not b;
    layer0_outputs(1254) <= not b;
    layer0_outputs(1255) <= not (a or b);
    layer0_outputs(1256) <= '1';
    layer0_outputs(1257) <= a or b;
    layer0_outputs(1258) <= not b;
    layer0_outputs(1259) <= a and b;
    layer0_outputs(1260) <= a or b;
    layer0_outputs(1261) <= not a or b;
    layer0_outputs(1262) <= a xor b;
    layer0_outputs(1263) <= not b;
    layer0_outputs(1264) <= not b or a;
    layer0_outputs(1265) <= b;
    layer0_outputs(1266) <= a xor b;
    layer0_outputs(1267) <= a and not b;
    layer0_outputs(1268) <= not (a or b);
    layer0_outputs(1269) <= '0';
    layer0_outputs(1270) <= a and not b;
    layer0_outputs(1271) <= not a or b;
    layer0_outputs(1272) <= not b;
    layer0_outputs(1273) <= b;
    layer0_outputs(1274) <= not b or a;
    layer0_outputs(1275) <= b and not a;
    layer0_outputs(1276) <= '0';
    layer0_outputs(1277) <= a;
    layer0_outputs(1278) <= not (a xor b);
    layer0_outputs(1279) <= not b or a;
    layer0_outputs(1280) <= not a;
    layer0_outputs(1281) <= a or b;
    layer0_outputs(1282) <= a;
    layer0_outputs(1283) <= not b or a;
    layer0_outputs(1284) <= b and not a;
    layer0_outputs(1285) <= not a or b;
    layer0_outputs(1286) <= not (a and b);
    layer0_outputs(1287) <= not (a or b);
    layer0_outputs(1288) <= not (a and b);
    layer0_outputs(1289) <= a;
    layer0_outputs(1290) <= a and not b;
    layer0_outputs(1291) <= '1';
    layer0_outputs(1292) <= a xor b;
    layer0_outputs(1293) <= not a;
    layer0_outputs(1294) <= not b;
    layer0_outputs(1295) <= b;
    layer0_outputs(1296) <= a and not b;
    layer0_outputs(1297) <= a or b;
    layer0_outputs(1298) <= not b;
    layer0_outputs(1299) <= not (a or b);
    layer0_outputs(1300) <= b;
    layer0_outputs(1301) <= not a;
    layer0_outputs(1302) <= b and not a;
    layer0_outputs(1303) <= '0';
    layer0_outputs(1304) <= not a or b;
    layer0_outputs(1305) <= not (a or b);
    layer0_outputs(1306) <= not (a xor b);
    layer0_outputs(1307) <= not (a or b);
    layer0_outputs(1308) <= '0';
    layer0_outputs(1309) <= a and not b;
    layer0_outputs(1310) <= not (a or b);
    layer0_outputs(1311) <= a or b;
    layer0_outputs(1312) <= a and not b;
    layer0_outputs(1313) <= a and b;
    layer0_outputs(1314) <= not b;
    layer0_outputs(1315) <= a xor b;
    layer0_outputs(1316) <= a and not b;
    layer0_outputs(1317) <= not b or a;
    layer0_outputs(1318) <= not (a and b);
    layer0_outputs(1319) <= not a;
    layer0_outputs(1320) <= not (a xor b);
    layer0_outputs(1321) <= not a;
    layer0_outputs(1322) <= not (a or b);
    layer0_outputs(1323) <= not b;
    layer0_outputs(1324) <= '1';
    layer0_outputs(1325) <= not (a or b);
    layer0_outputs(1326) <= not (a xor b);
    layer0_outputs(1327) <= not (a xor b);
    layer0_outputs(1328) <= a or b;
    layer0_outputs(1329) <= not b;
    layer0_outputs(1330) <= not a;
    layer0_outputs(1331) <= not (a or b);
    layer0_outputs(1332) <= not a or b;
    layer0_outputs(1333) <= not a;
    layer0_outputs(1334) <= b;
    layer0_outputs(1335) <= not a or b;
    layer0_outputs(1336) <= '0';
    layer0_outputs(1337) <= not a;
    layer0_outputs(1338) <= not (a and b);
    layer0_outputs(1339) <= a;
    layer0_outputs(1340) <= b;
    layer0_outputs(1341) <= a or b;
    layer0_outputs(1342) <= not b or a;
    layer0_outputs(1343) <= b;
    layer0_outputs(1344) <= not a or b;
    layer0_outputs(1345) <= not b or a;
    layer0_outputs(1346) <= a;
    layer0_outputs(1347) <= not (a or b);
    layer0_outputs(1348) <= not a or b;
    layer0_outputs(1349) <= '1';
    layer0_outputs(1350) <= a xor b;
    layer0_outputs(1351) <= a xor b;
    layer0_outputs(1352) <= not b;
    layer0_outputs(1353) <= b and not a;
    layer0_outputs(1354) <= a and not b;
    layer0_outputs(1355) <= a xor b;
    layer0_outputs(1356) <= a or b;
    layer0_outputs(1357) <= not a or b;
    layer0_outputs(1358) <= b;
    layer0_outputs(1359) <= a;
    layer0_outputs(1360) <= a;
    layer0_outputs(1361) <= a xor b;
    layer0_outputs(1362) <= a and not b;
    layer0_outputs(1363) <= '1';
    layer0_outputs(1364) <= not (a or b);
    layer0_outputs(1365) <= not b;
    layer0_outputs(1366) <= a xor b;
    layer0_outputs(1367) <= b;
    layer0_outputs(1368) <= a;
    layer0_outputs(1369) <= a xor b;
    layer0_outputs(1370) <= a or b;
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= not (a xor b);
    layer0_outputs(1373) <= not b or a;
    layer0_outputs(1374) <= b;
    layer0_outputs(1375) <= b;
    layer0_outputs(1376) <= not b;
    layer0_outputs(1377) <= '0';
    layer0_outputs(1378) <= not b;
    layer0_outputs(1379) <= b;
    layer0_outputs(1380) <= not b;
    layer0_outputs(1381) <= '1';
    layer0_outputs(1382) <= not (a or b);
    layer0_outputs(1383) <= a xor b;
    layer0_outputs(1384) <= a and not b;
    layer0_outputs(1385) <= b and not a;
    layer0_outputs(1386) <= '0';
    layer0_outputs(1387) <= a;
    layer0_outputs(1388) <= '0';
    layer0_outputs(1389) <= not b;
    layer0_outputs(1390) <= a and not b;
    layer0_outputs(1391) <= not (a or b);
    layer0_outputs(1392) <= not a;
    layer0_outputs(1393) <= not (a xor b);
    layer0_outputs(1394) <= not (a xor b);
    layer0_outputs(1395) <= not (a or b);
    layer0_outputs(1396) <= not b or a;
    layer0_outputs(1397) <= not (a and b);
    layer0_outputs(1398) <= b and not a;
    layer0_outputs(1399) <= not (a xor b);
    layer0_outputs(1400) <= b and not a;
    layer0_outputs(1401) <= not a;
    layer0_outputs(1402) <= not (a or b);
    layer0_outputs(1403) <= not (a xor b);
    layer0_outputs(1404) <= not (a xor b);
    layer0_outputs(1405) <= a and not b;
    layer0_outputs(1406) <= not b;
    layer0_outputs(1407) <= a and not b;
    layer0_outputs(1408) <= a xor b;
    layer0_outputs(1409) <= b;
    layer0_outputs(1410) <= b and not a;
    layer0_outputs(1411) <= a or b;
    layer0_outputs(1412) <= not b or a;
    layer0_outputs(1413) <= not (a or b);
    layer0_outputs(1414) <= '0';
    layer0_outputs(1415) <= not a or b;
    layer0_outputs(1416) <= b and not a;
    layer0_outputs(1417) <= a or b;
    layer0_outputs(1418) <= not (a or b);
    layer0_outputs(1419) <= a xor b;
    layer0_outputs(1420) <= not (a or b);
    layer0_outputs(1421) <= not (a or b);
    layer0_outputs(1422) <= not a;
    layer0_outputs(1423) <= b and not a;
    layer0_outputs(1424) <= a;
    layer0_outputs(1425) <= a xor b;
    layer0_outputs(1426) <= a or b;
    layer0_outputs(1427) <= a or b;
    layer0_outputs(1428) <= a;
    layer0_outputs(1429) <= b and not a;
    layer0_outputs(1430) <= not (a xor b);
    layer0_outputs(1431) <= a or b;
    layer0_outputs(1432) <= a;
    layer0_outputs(1433) <= not (a and b);
    layer0_outputs(1434) <= not (a or b);
    layer0_outputs(1435) <= not (a or b);
    layer0_outputs(1436) <= not (a and b);
    layer0_outputs(1437) <= a;
    layer0_outputs(1438) <= a or b;
    layer0_outputs(1439) <= not (a or b);
    layer0_outputs(1440) <= a or b;
    layer0_outputs(1441) <= a;
    layer0_outputs(1442) <= not a or b;
    layer0_outputs(1443) <= b and not a;
    layer0_outputs(1444) <= b and not a;
    layer0_outputs(1445) <= not (a and b);
    layer0_outputs(1446) <= not a;
    layer0_outputs(1447) <= '1';
    layer0_outputs(1448) <= a xor b;
    layer0_outputs(1449) <= a;
    layer0_outputs(1450) <= a xor b;
    layer0_outputs(1451) <= b and not a;
    layer0_outputs(1452) <= not (a or b);
    layer0_outputs(1453) <= not (a or b);
    layer0_outputs(1454) <= a and b;
    layer0_outputs(1455) <= '0';
    layer0_outputs(1456) <= not (a xor b);
    layer0_outputs(1457) <= a or b;
    layer0_outputs(1458) <= b;
    layer0_outputs(1459) <= a and not b;
    layer0_outputs(1460) <= not (a xor b);
    layer0_outputs(1461) <= b and not a;
    layer0_outputs(1462) <= a;
    layer0_outputs(1463) <= not b;
    layer0_outputs(1464) <= a xor b;
    layer0_outputs(1465) <= a and b;
    layer0_outputs(1466) <= b;
    layer0_outputs(1467) <= b;
    layer0_outputs(1468) <= not b;
    layer0_outputs(1469) <= b and not a;
    layer0_outputs(1470) <= '0';
    layer0_outputs(1471) <= a and not b;
    layer0_outputs(1472) <= a or b;
    layer0_outputs(1473) <= a;
    layer0_outputs(1474) <= not b or a;
    layer0_outputs(1475) <= not (a or b);
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= a;
    layer0_outputs(1478) <= a and not b;
    layer0_outputs(1479) <= a and not b;
    layer0_outputs(1480) <= not a;
    layer0_outputs(1481) <= not a;
    layer0_outputs(1482) <= '1';
    layer0_outputs(1483) <= not b;
    layer0_outputs(1484) <= not (a or b);
    layer0_outputs(1485) <= a or b;
    layer0_outputs(1486) <= a;
    layer0_outputs(1487) <= not a or b;
    layer0_outputs(1488) <= a and not b;
    layer0_outputs(1489) <= a and not b;
    layer0_outputs(1490) <= b;
    layer0_outputs(1491) <= b;
    layer0_outputs(1492) <= not b or a;
    layer0_outputs(1493) <= not a;
    layer0_outputs(1494) <= not (a xor b);
    layer0_outputs(1495) <= not a or b;
    layer0_outputs(1496) <= not (a or b);
    layer0_outputs(1497) <= a xor b;
    layer0_outputs(1498) <= '0';
    layer0_outputs(1499) <= b;
    layer0_outputs(1500) <= not b or a;
    layer0_outputs(1501) <= '1';
    layer0_outputs(1502) <= a and b;
    layer0_outputs(1503) <= not (a or b);
    layer0_outputs(1504) <= not a or b;
    layer0_outputs(1505) <= not (a and b);
    layer0_outputs(1506) <= not a;
    layer0_outputs(1507) <= a or b;
    layer0_outputs(1508) <= not (a xor b);
    layer0_outputs(1509) <= a and b;
    layer0_outputs(1510) <= b;
    layer0_outputs(1511) <= a or b;
    layer0_outputs(1512) <= not a;
    layer0_outputs(1513) <= a and not b;
    layer0_outputs(1514) <= '1';
    layer0_outputs(1515) <= b;
    layer0_outputs(1516) <= a or b;
    layer0_outputs(1517) <= not (a and b);
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= b and not a;
    layer0_outputs(1520) <= a and not b;
    layer0_outputs(1521) <= not a or b;
    layer0_outputs(1522) <= a or b;
    layer0_outputs(1523) <= a or b;
    layer0_outputs(1524) <= b and not a;
    layer0_outputs(1525) <= not b;
    layer0_outputs(1526) <= b and not a;
    layer0_outputs(1527) <= '0';
    layer0_outputs(1528) <= a;
    layer0_outputs(1529) <= b and not a;
    layer0_outputs(1530) <= a or b;
    layer0_outputs(1531) <= b and not a;
    layer0_outputs(1532) <= not (a or b);
    layer0_outputs(1533) <= a or b;
    layer0_outputs(1534) <= a or b;
    layer0_outputs(1535) <= '0';
    layer0_outputs(1536) <= not a;
    layer0_outputs(1537) <= not a;
    layer0_outputs(1538) <= a or b;
    layer0_outputs(1539) <= not (a or b);
    layer0_outputs(1540) <= not (a xor b);
    layer0_outputs(1541) <= a;
    layer0_outputs(1542) <= a and not b;
    layer0_outputs(1543) <= not b or a;
    layer0_outputs(1544) <= not b or a;
    layer0_outputs(1545) <= not (a or b);
    layer0_outputs(1546) <= not b or a;
    layer0_outputs(1547) <= a and b;
    layer0_outputs(1548) <= a;
    layer0_outputs(1549) <= not (a or b);
    layer0_outputs(1550) <= not b;
    layer0_outputs(1551) <= a or b;
    layer0_outputs(1552) <= not a or b;
    layer0_outputs(1553) <= a or b;
    layer0_outputs(1554) <= b;
    layer0_outputs(1555) <= a and b;
    layer0_outputs(1556) <= not b;
    layer0_outputs(1557) <= '0';
    layer0_outputs(1558) <= b;
    layer0_outputs(1559) <= b;
    layer0_outputs(1560) <= not (a xor b);
    layer0_outputs(1561) <= a and b;
    layer0_outputs(1562) <= b;
    layer0_outputs(1563) <= not a;
    layer0_outputs(1564) <= not b or a;
    layer0_outputs(1565) <= a and b;
    layer0_outputs(1566) <= b and not a;
    layer0_outputs(1567) <= not (a and b);
    layer0_outputs(1568) <= a or b;
    layer0_outputs(1569) <= not a;
    layer0_outputs(1570) <= a and b;
    layer0_outputs(1571) <= a;
    layer0_outputs(1572) <= a or b;
    layer0_outputs(1573) <= b and not a;
    layer0_outputs(1574) <= not b or a;
    layer0_outputs(1575) <= a;
    layer0_outputs(1576) <= a;
    layer0_outputs(1577) <= a or b;
    layer0_outputs(1578) <= a or b;
    layer0_outputs(1579) <= a and b;
    layer0_outputs(1580) <= a and not b;
    layer0_outputs(1581) <= '1';
    layer0_outputs(1582) <= b and not a;
    layer0_outputs(1583) <= not b;
    layer0_outputs(1584) <= not b or a;
    layer0_outputs(1585) <= not b;
    layer0_outputs(1586) <= b and not a;
    layer0_outputs(1587) <= not b;
    layer0_outputs(1588) <= not (a xor b);
    layer0_outputs(1589) <= not a;
    layer0_outputs(1590) <= not a or b;
    layer0_outputs(1591) <= b and not a;
    layer0_outputs(1592) <= b and not a;
    layer0_outputs(1593) <= a and b;
    layer0_outputs(1594) <= not (a or b);
    layer0_outputs(1595) <= a and b;
    layer0_outputs(1596) <= b;
    layer0_outputs(1597) <= a and not b;
    layer0_outputs(1598) <= not b;
    layer0_outputs(1599) <= b and not a;
    layer0_outputs(1600) <= not a or b;
    layer0_outputs(1601) <= a or b;
    layer0_outputs(1602) <= not (a or b);
    layer0_outputs(1603) <= not (a or b);
    layer0_outputs(1604) <= b and not a;
    layer0_outputs(1605) <= a or b;
    layer0_outputs(1606) <= a and b;
    layer0_outputs(1607) <= '1';
    layer0_outputs(1608) <= not (a xor b);
    layer0_outputs(1609) <= not (a and b);
    layer0_outputs(1610) <= a and not b;
    layer0_outputs(1611) <= b;
    layer0_outputs(1612) <= not a or b;
    layer0_outputs(1613) <= not a;
    layer0_outputs(1614) <= a;
    layer0_outputs(1615) <= b;
    layer0_outputs(1616) <= not (a or b);
    layer0_outputs(1617) <= not b or a;
    layer0_outputs(1618) <= not (a and b);
    layer0_outputs(1619) <= a and not b;
    layer0_outputs(1620) <= not (a and b);
    layer0_outputs(1621) <= not b;
    layer0_outputs(1622) <= a and not b;
    layer0_outputs(1623) <= not b or a;
    layer0_outputs(1624) <= not (a xor b);
    layer0_outputs(1625) <= b and not a;
    layer0_outputs(1626) <= not b or a;
    layer0_outputs(1627) <= b;
    layer0_outputs(1628) <= not (a or b);
    layer0_outputs(1629) <= not a or b;
    layer0_outputs(1630) <= not (a or b);
    layer0_outputs(1631) <= a;
    layer0_outputs(1632) <= not b or a;
    layer0_outputs(1633) <= '1';
    layer0_outputs(1634) <= not (a xor b);
    layer0_outputs(1635) <= b;
    layer0_outputs(1636) <= a and b;
    layer0_outputs(1637) <= b and not a;
    layer0_outputs(1638) <= a or b;
    layer0_outputs(1639) <= not b;
    layer0_outputs(1640) <= a or b;
    layer0_outputs(1641) <= a;
    layer0_outputs(1642) <= a or b;
    layer0_outputs(1643) <= not a;
    layer0_outputs(1644) <= not b;
    layer0_outputs(1645) <= a or b;
    layer0_outputs(1646) <= a and b;
    layer0_outputs(1647) <= not a;
    layer0_outputs(1648) <= not (a xor b);
    layer0_outputs(1649) <= a or b;
    layer0_outputs(1650) <= a;
    layer0_outputs(1651) <= a and not b;
    layer0_outputs(1652) <= '0';
    layer0_outputs(1653) <= b;
    layer0_outputs(1654) <= not a;
    layer0_outputs(1655) <= not (a and b);
    layer0_outputs(1656) <= not b or a;
    layer0_outputs(1657) <= not a or b;
    layer0_outputs(1658) <= not (a xor b);
    layer0_outputs(1659) <= a or b;
    layer0_outputs(1660) <= b and not a;
    layer0_outputs(1661) <= not (a xor b);
    layer0_outputs(1662) <= not (a or b);
    layer0_outputs(1663) <= not (a or b);
    layer0_outputs(1664) <= not b or a;
    layer0_outputs(1665) <= a or b;
    layer0_outputs(1666) <= not (a and b);
    layer0_outputs(1667) <= a or b;
    layer0_outputs(1668) <= a or b;
    layer0_outputs(1669) <= not a or b;
    layer0_outputs(1670) <= b;
    layer0_outputs(1671) <= '1';
    layer0_outputs(1672) <= a;
    layer0_outputs(1673) <= not (a xor b);
    layer0_outputs(1674) <= b and not a;
    layer0_outputs(1675) <= b and not a;
    layer0_outputs(1676) <= not a;
    layer0_outputs(1677) <= not b;
    layer0_outputs(1678) <= not b or a;
    layer0_outputs(1679) <= a and not b;
    layer0_outputs(1680) <= a or b;
    layer0_outputs(1681) <= a and b;
    layer0_outputs(1682) <= a;
    layer0_outputs(1683) <= '0';
    layer0_outputs(1684) <= not b or a;
    layer0_outputs(1685) <= not b or a;
    layer0_outputs(1686) <= a;
    layer0_outputs(1687) <= not b;
    layer0_outputs(1688) <= not a or b;
    layer0_outputs(1689) <= not (a xor b);
    layer0_outputs(1690) <= not b;
    layer0_outputs(1691) <= a;
    layer0_outputs(1692) <= b and not a;
    layer0_outputs(1693) <= not (a xor b);
    layer0_outputs(1694) <= not (a or b);
    layer0_outputs(1695) <= a or b;
    layer0_outputs(1696) <= a or b;
    layer0_outputs(1697) <= '0';
    layer0_outputs(1698) <= not b;
    layer0_outputs(1699) <= not (a or b);
    layer0_outputs(1700) <= not (a and b);
    layer0_outputs(1701) <= not (a xor b);
    layer0_outputs(1702) <= not (a or b);
    layer0_outputs(1703) <= not (a or b);
    layer0_outputs(1704) <= not a or b;
    layer0_outputs(1705) <= not a;
    layer0_outputs(1706) <= b;
    layer0_outputs(1707) <= a xor b;
    layer0_outputs(1708) <= b and not a;
    layer0_outputs(1709) <= not (a and b);
    layer0_outputs(1710) <= a;
    layer0_outputs(1711) <= not (a xor b);
    layer0_outputs(1712) <= a or b;
    layer0_outputs(1713) <= a or b;
    layer0_outputs(1714) <= a xor b;
    layer0_outputs(1715) <= not b;
    layer0_outputs(1716) <= a xor b;
    layer0_outputs(1717) <= not b or a;
    layer0_outputs(1718) <= not a or b;
    layer0_outputs(1719) <= not a or b;
    layer0_outputs(1720) <= a xor b;
    layer0_outputs(1721) <= b and not a;
    layer0_outputs(1722) <= a or b;
    layer0_outputs(1723) <= b;
    layer0_outputs(1724) <= '0';
    layer0_outputs(1725) <= a and not b;
    layer0_outputs(1726) <= '0';
    layer0_outputs(1727) <= not (a or b);
    layer0_outputs(1728) <= not a or b;
    layer0_outputs(1729) <= not b or a;
    layer0_outputs(1730) <= a and not b;
    layer0_outputs(1731) <= not (a or b);
    layer0_outputs(1732) <= not b;
    layer0_outputs(1733) <= b and not a;
    layer0_outputs(1734) <= a and b;
    layer0_outputs(1735) <= '1';
    layer0_outputs(1736) <= not a;
    layer0_outputs(1737) <= a or b;
    layer0_outputs(1738) <= not (a xor b);
    layer0_outputs(1739) <= a;
    layer0_outputs(1740) <= a;
    layer0_outputs(1741) <= not b;
    layer0_outputs(1742) <= a or b;
    layer0_outputs(1743) <= b and not a;
    layer0_outputs(1744) <= not (a or b);
    layer0_outputs(1745) <= not (a or b);
    layer0_outputs(1746) <= a xor b;
    layer0_outputs(1747) <= not a or b;
    layer0_outputs(1748) <= not b or a;
    layer0_outputs(1749) <= a and not b;
    layer0_outputs(1750) <= b and not a;
    layer0_outputs(1751) <= a xor b;
    layer0_outputs(1752) <= a xor b;
    layer0_outputs(1753) <= '1';
    layer0_outputs(1754) <= a or b;
    layer0_outputs(1755) <= not (a or b);
    layer0_outputs(1756) <= not (a or b);
    layer0_outputs(1757) <= not (a or b);
    layer0_outputs(1758) <= not a or b;
    layer0_outputs(1759) <= a or b;
    layer0_outputs(1760) <= b;
    layer0_outputs(1761) <= b;
    layer0_outputs(1762) <= not (a or b);
    layer0_outputs(1763) <= a or b;
    layer0_outputs(1764) <= not a;
    layer0_outputs(1765) <= not (a and b);
    layer0_outputs(1766) <= not a;
    layer0_outputs(1767) <= b;
    layer0_outputs(1768) <= not a or b;
    layer0_outputs(1769) <= not (a or b);
    layer0_outputs(1770) <= b;
    layer0_outputs(1771) <= not a or b;
    layer0_outputs(1772) <= not a or b;
    layer0_outputs(1773) <= a and not b;
    layer0_outputs(1774) <= a or b;
    layer0_outputs(1775) <= not (a or b);
    layer0_outputs(1776) <= not (a or b);
    layer0_outputs(1777) <= not a or b;
    layer0_outputs(1778) <= b;
    layer0_outputs(1779) <= not b;
    layer0_outputs(1780) <= b and not a;
    layer0_outputs(1781) <= a or b;
    layer0_outputs(1782) <= not (a or b);
    layer0_outputs(1783) <= a or b;
    layer0_outputs(1784) <= b;
    layer0_outputs(1785) <= a and not b;
    layer0_outputs(1786) <= a or b;
    layer0_outputs(1787) <= a;
    layer0_outputs(1788) <= not (a xor b);
    layer0_outputs(1789) <= not (a or b);
    layer0_outputs(1790) <= a xor b;
    layer0_outputs(1791) <= a and b;
    layer0_outputs(1792) <= a and not b;
    layer0_outputs(1793) <= not a;
    layer0_outputs(1794) <= a xor b;
    layer0_outputs(1795) <= a or b;
    layer0_outputs(1796) <= b;
    layer0_outputs(1797) <= not b;
    layer0_outputs(1798) <= b;
    layer0_outputs(1799) <= b;
    layer0_outputs(1800) <= not b or a;
    layer0_outputs(1801) <= a or b;
    layer0_outputs(1802) <= a;
    layer0_outputs(1803) <= '1';
    layer0_outputs(1804) <= a xor b;
    layer0_outputs(1805) <= not (a or b);
    layer0_outputs(1806) <= b and not a;
    layer0_outputs(1807) <= b;
    layer0_outputs(1808) <= a and not b;
    layer0_outputs(1809) <= b;
    layer0_outputs(1810) <= not a or b;
    layer0_outputs(1811) <= not (a xor b);
    layer0_outputs(1812) <= b;
    layer0_outputs(1813) <= not b or a;
    layer0_outputs(1814) <= not (a or b);
    layer0_outputs(1815) <= not (a or b);
    layer0_outputs(1816) <= b;
    layer0_outputs(1817) <= not (a xor b);
    layer0_outputs(1818) <= a xor b;
    layer0_outputs(1819) <= a;
    layer0_outputs(1820) <= not b or a;
    layer0_outputs(1821) <= a xor b;
    layer0_outputs(1822) <= a;
    layer0_outputs(1823) <= a;
    layer0_outputs(1824) <= b and not a;
    layer0_outputs(1825) <= not a;
    layer0_outputs(1826) <= a and b;
    layer0_outputs(1827) <= a xor b;
    layer0_outputs(1828) <= a and not b;
    layer0_outputs(1829) <= '0';
    layer0_outputs(1830) <= not a or b;
    layer0_outputs(1831) <= a xor b;
    layer0_outputs(1832) <= '1';
    layer0_outputs(1833) <= not (a xor b);
    layer0_outputs(1834) <= not a or b;
    layer0_outputs(1835) <= '1';
    layer0_outputs(1836) <= not b;
    layer0_outputs(1837) <= not b;
    layer0_outputs(1838) <= a or b;
    layer0_outputs(1839) <= not (a or b);
    layer0_outputs(1840) <= not b or a;
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= not b;
    layer0_outputs(1843) <= b and not a;
    layer0_outputs(1844) <= a;
    layer0_outputs(1845) <= not a;
    layer0_outputs(1846) <= not (a or b);
    layer0_outputs(1847) <= not b;
    layer0_outputs(1848) <= not b or a;
    layer0_outputs(1849) <= not (a or b);
    layer0_outputs(1850) <= not (a or b);
    layer0_outputs(1851) <= not (a and b);
    layer0_outputs(1852) <= not b or a;
    layer0_outputs(1853) <= not a or b;
    layer0_outputs(1854) <= not (a or b);
    layer0_outputs(1855) <= not b;
    layer0_outputs(1856) <= not (a or b);
    layer0_outputs(1857) <= a or b;
    layer0_outputs(1858) <= a or b;
    layer0_outputs(1859) <= b;
    layer0_outputs(1860) <= not b or a;
    layer0_outputs(1861) <= '1';
    layer0_outputs(1862) <= a and not b;
    layer0_outputs(1863) <= a or b;
    layer0_outputs(1864) <= not b or a;
    layer0_outputs(1865) <= a xor b;
    layer0_outputs(1866) <= not (a or b);
    layer0_outputs(1867) <= not b;
    layer0_outputs(1868) <= b;
    layer0_outputs(1869) <= not (a or b);
    layer0_outputs(1870) <= a or b;
    layer0_outputs(1871) <= a or b;
    layer0_outputs(1872) <= not a;
    layer0_outputs(1873) <= not a;
    layer0_outputs(1874) <= not b;
    layer0_outputs(1875) <= not b or a;
    layer0_outputs(1876) <= not b;
    layer0_outputs(1877) <= not b or a;
    layer0_outputs(1878) <= not (a or b);
    layer0_outputs(1879) <= not b;
    layer0_outputs(1880) <= not (a and b);
    layer0_outputs(1881) <= not a or b;
    layer0_outputs(1882) <= not b or a;
    layer0_outputs(1883) <= a;
    layer0_outputs(1884) <= a and not b;
    layer0_outputs(1885) <= not b or a;
    layer0_outputs(1886) <= not (a or b);
    layer0_outputs(1887) <= a;
    layer0_outputs(1888) <= not b or a;
    layer0_outputs(1889) <= not b;
    layer0_outputs(1890) <= a or b;
    layer0_outputs(1891) <= not b;
    layer0_outputs(1892) <= a or b;
    layer0_outputs(1893) <= a;
    layer0_outputs(1894) <= a or b;
    layer0_outputs(1895) <= b;
    layer0_outputs(1896) <= a;
    layer0_outputs(1897) <= not a;
    layer0_outputs(1898) <= not b or a;
    layer0_outputs(1899) <= a and not b;
    layer0_outputs(1900) <= b and not a;
    layer0_outputs(1901) <= a;
    layer0_outputs(1902) <= b and not a;
    layer0_outputs(1903) <= '0';
    layer0_outputs(1904) <= a or b;
    layer0_outputs(1905) <= not b;
    layer0_outputs(1906) <= a and b;
    layer0_outputs(1907) <= '0';
    layer0_outputs(1908) <= not b;
    layer0_outputs(1909) <= b and not a;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= not (a and b);
    layer0_outputs(1912) <= a xor b;
    layer0_outputs(1913) <= b;
    layer0_outputs(1914) <= not a or b;
    layer0_outputs(1915) <= not (a or b);
    layer0_outputs(1916) <= a and b;
    layer0_outputs(1917) <= not b;
    layer0_outputs(1918) <= a;
    layer0_outputs(1919) <= b and not a;
    layer0_outputs(1920) <= b;
    layer0_outputs(1921) <= b;
    layer0_outputs(1922) <= not (a or b);
    layer0_outputs(1923) <= not b;
    layer0_outputs(1924) <= not (a xor b);
    layer0_outputs(1925) <= not a;
    layer0_outputs(1926) <= not a or b;
    layer0_outputs(1927) <= a;
    layer0_outputs(1928) <= a xor b;
    layer0_outputs(1929) <= '0';
    layer0_outputs(1930) <= not b;
    layer0_outputs(1931) <= not (a xor b);
    layer0_outputs(1932) <= b;
    layer0_outputs(1933) <= not (a xor b);
    layer0_outputs(1934) <= a or b;
    layer0_outputs(1935) <= a xor b;
    layer0_outputs(1936) <= b and not a;
    layer0_outputs(1937) <= b;
    layer0_outputs(1938) <= a;
    layer0_outputs(1939) <= a or b;
    layer0_outputs(1940) <= not a;
    layer0_outputs(1941) <= b and not a;
    layer0_outputs(1942) <= a and b;
    layer0_outputs(1943) <= not (a or b);
    layer0_outputs(1944) <= not a or b;
    layer0_outputs(1945) <= a and not b;
    layer0_outputs(1946) <= a and not b;
    layer0_outputs(1947) <= a or b;
    layer0_outputs(1948) <= b;
    layer0_outputs(1949) <= a;
    layer0_outputs(1950) <= not b;
    layer0_outputs(1951) <= a and not b;
    layer0_outputs(1952) <= not (a or b);
    layer0_outputs(1953) <= not b;
    layer0_outputs(1954) <= not b or a;
    layer0_outputs(1955) <= not a;
    layer0_outputs(1956) <= a or b;
    layer0_outputs(1957) <= not b;
    layer0_outputs(1958) <= a xor b;
    layer0_outputs(1959) <= a xor b;
    layer0_outputs(1960) <= not (a and b);
    layer0_outputs(1961) <= not b or a;
    layer0_outputs(1962) <= a or b;
    layer0_outputs(1963) <= a and b;
    layer0_outputs(1964) <= a or b;
    layer0_outputs(1965) <= not b or a;
    layer0_outputs(1966) <= not (a xor b);
    layer0_outputs(1967) <= not a;
    layer0_outputs(1968) <= not b;
    layer0_outputs(1969) <= a;
    layer0_outputs(1970) <= a or b;
    layer0_outputs(1971) <= '1';
    layer0_outputs(1972) <= not a;
    layer0_outputs(1973) <= not (a and b);
    layer0_outputs(1974) <= not b;
    layer0_outputs(1975) <= a xor b;
    layer0_outputs(1976) <= not (a or b);
    layer0_outputs(1977) <= b and not a;
    layer0_outputs(1978) <= not a or b;
    layer0_outputs(1979) <= a;
    layer0_outputs(1980) <= a or b;
    layer0_outputs(1981) <= not a or b;
    layer0_outputs(1982) <= a xor b;
    layer0_outputs(1983) <= not (a xor b);
    layer0_outputs(1984) <= '0';
    layer0_outputs(1985) <= b;
    layer0_outputs(1986) <= a;
    layer0_outputs(1987) <= not a;
    layer0_outputs(1988) <= a or b;
    layer0_outputs(1989) <= a;
    layer0_outputs(1990) <= a and not b;
    layer0_outputs(1991) <= not a;
    layer0_outputs(1992) <= b and not a;
    layer0_outputs(1993) <= '0';
    layer0_outputs(1994) <= not b or a;
    layer0_outputs(1995) <= b and not a;
    layer0_outputs(1996) <= not b or a;
    layer0_outputs(1997) <= a and not b;
    layer0_outputs(1998) <= '1';
    layer0_outputs(1999) <= not (a xor b);
    layer0_outputs(2000) <= b;
    layer0_outputs(2001) <= a xor b;
    layer0_outputs(2002) <= b;
    layer0_outputs(2003) <= not a or b;
    layer0_outputs(2004) <= not (a xor b);
    layer0_outputs(2005) <= a xor b;
    layer0_outputs(2006) <= a and not b;
    layer0_outputs(2007) <= b;
    layer0_outputs(2008) <= not b;
    layer0_outputs(2009) <= a and b;
    layer0_outputs(2010) <= not b;
    layer0_outputs(2011) <= not b;
    layer0_outputs(2012) <= a;
    layer0_outputs(2013) <= b and not a;
    layer0_outputs(2014) <= a and not b;
    layer0_outputs(2015) <= not a or b;
    layer0_outputs(2016) <= a xor b;
    layer0_outputs(2017) <= not a;
    layer0_outputs(2018) <= not a;
    layer0_outputs(2019) <= not (a xor b);
    layer0_outputs(2020) <= not a;
    layer0_outputs(2021) <= not b or a;
    layer0_outputs(2022) <= a and not b;
    layer0_outputs(2023) <= not (a or b);
    layer0_outputs(2024) <= not (a and b);
    layer0_outputs(2025) <= '1';
    layer0_outputs(2026) <= a or b;
    layer0_outputs(2027) <= a;
    layer0_outputs(2028) <= a or b;
    layer0_outputs(2029) <= b;
    layer0_outputs(2030) <= b and not a;
    layer0_outputs(2031) <= '1';
    layer0_outputs(2032) <= not (a xor b);
    layer0_outputs(2033) <= a xor b;
    layer0_outputs(2034) <= not a or b;
    layer0_outputs(2035) <= a xor b;
    layer0_outputs(2036) <= not a;
    layer0_outputs(2037) <= '0';
    layer0_outputs(2038) <= b;
    layer0_outputs(2039) <= not b or a;
    layer0_outputs(2040) <= '1';
    layer0_outputs(2041) <= '0';
    layer0_outputs(2042) <= not (a or b);
    layer0_outputs(2043) <= a and not b;
    layer0_outputs(2044) <= not a;
    layer0_outputs(2045) <= a and not b;
    layer0_outputs(2046) <= a and not b;
    layer0_outputs(2047) <= not a or b;
    layer0_outputs(2048) <= b;
    layer0_outputs(2049) <= not (a xor b);
    layer0_outputs(2050) <= not (a xor b);
    layer0_outputs(2051) <= not (a or b);
    layer0_outputs(2052) <= not (a and b);
    layer0_outputs(2053) <= not (a or b);
    layer0_outputs(2054) <= b;
    layer0_outputs(2055) <= not b or a;
    layer0_outputs(2056) <= a and b;
    layer0_outputs(2057) <= b and not a;
    layer0_outputs(2058) <= a and not b;
    layer0_outputs(2059) <= a;
    layer0_outputs(2060) <= a;
    layer0_outputs(2061) <= not a or b;
    layer0_outputs(2062) <= not (a xor b);
    layer0_outputs(2063) <= a or b;
    layer0_outputs(2064) <= a or b;
    layer0_outputs(2065) <= '0';
    layer0_outputs(2066) <= b and not a;
    layer0_outputs(2067) <= b and not a;
    layer0_outputs(2068) <= a or b;
    layer0_outputs(2069) <= b and not a;
    layer0_outputs(2070) <= a;
    layer0_outputs(2071) <= not (a or b);
    layer0_outputs(2072) <= '1';
    layer0_outputs(2073) <= b and not a;
    layer0_outputs(2074) <= a xor b;
    layer0_outputs(2075) <= b;
    layer0_outputs(2076) <= not (a or b);
    layer0_outputs(2077) <= not a or b;
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= not (a or b);
    layer0_outputs(2080) <= not b;
    layer0_outputs(2081) <= a or b;
    layer0_outputs(2082) <= a or b;
    layer0_outputs(2083) <= a and b;
    layer0_outputs(2084) <= a xor b;
    layer0_outputs(2085) <= not b;
    layer0_outputs(2086) <= a xor b;
    layer0_outputs(2087) <= '0';
    layer0_outputs(2088) <= not (a xor b);
    layer0_outputs(2089) <= a and b;
    layer0_outputs(2090) <= a or b;
    layer0_outputs(2091) <= a and not b;
    layer0_outputs(2092) <= not (a xor b);
    layer0_outputs(2093) <= not (a or b);
    layer0_outputs(2094) <= b;
    layer0_outputs(2095) <= a xor b;
    layer0_outputs(2096) <= not (a and b);
    layer0_outputs(2097) <= a xor b;
    layer0_outputs(2098) <= not (a or b);
    layer0_outputs(2099) <= b;
    layer0_outputs(2100) <= not a;
    layer0_outputs(2101) <= a and not b;
    layer0_outputs(2102) <= not b;
    layer0_outputs(2103) <= not a or b;
    layer0_outputs(2104) <= not (a or b);
    layer0_outputs(2105) <= not b or a;
    layer0_outputs(2106) <= not b or a;
    layer0_outputs(2107) <= b and not a;
    layer0_outputs(2108) <= b;
    layer0_outputs(2109) <= not (a and b);
    layer0_outputs(2110) <= a and b;
    layer0_outputs(2111) <= a or b;
    layer0_outputs(2112) <= not b;
    layer0_outputs(2113) <= not (a or b);
    layer0_outputs(2114) <= not b;
    layer0_outputs(2115) <= a or b;
    layer0_outputs(2116) <= a and not b;
    layer0_outputs(2117) <= not a or b;
    layer0_outputs(2118) <= a and b;
    layer0_outputs(2119) <= a xor b;
    layer0_outputs(2120) <= not a or b;
    layer0_outputs(2121) <= not a;
    layer0_outputs(2122) <= a;
    layer0_outputs(2123) <= not a;
    layer0_outputs(2124) <= not a;
    layer0_outputs(2125) <= not b;
    layer0_outputs(2126) <= not (a xor b);
    layer0_outputs(2127) <= a or b;
    layer0_outputs(2128) <= b;
    layer0_outputs(2129) <= '1';
    layer0_outputs(2130) <= a xor b;
    layer0_outputs(2131) <= a xor b;
    layer0_outputs(2132) <= not (a or b);
    layer0_outputs(2133) <= a and b;
    layer0_outputs(2134) <= a and b;
    layer0_outputs(2135) <= b and not a;
    layer0_outputs(2136) <= a and not b;
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= a and not b;
    layer0_outputs(2139) <= '0';
    layer0_outputs(2140) <= b and not a;
    layer0_outputs(2141) <= a xor b;
    layer0_outputs(2142) <= not (a xor b);
    layer0_outputs(2143) <= not (a or b);
    layer0_outputs(2144) <= a and not b;
    layer0_outputs(2145) <= '1';
    layer0_outputs(2146) <= not a;
    layer0_outputs(2147) <= not (a or b);
    layer0_outputs(2148) <= not b or a;
    layer0_outputs(2149) <= b;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= not (a xor b);
    layer0_outputs(2152) <= b and not a;
    layer0_outputs(2153) <= a xor b;
    layer0_outputs(2154) <= not b;
    layer0_outputs(2155) <= not b or a;
    layer0_outputs(2156) <= not a or b;
    layer0_outputs(2157) <= b;
    layer0_outputs(2158) <= not a or b;
    layer0_outputs(2159) <= a xor b;
    layer0_outputs(2160) <= not (a or b);
    layer0_outputs(2161) <= a or b;
    layer0_outputs(2162) <= not (a xor b);
    layer0_outputs(2163) <= not b;
    layer0_outputs(2164) <= '0';
    layer0_outputs(2165) <= not b;
    layer0_outputs(2166) <= a;
    layer0_outputs(2167) <= not a or b;
    layer0_outputs(2168) <= not a;
    layer0_outputs(2169) <= a and not b;
    layer0_outputs(2170) <= a;
    layer0_outputs(2171) <= a and not b;
    layer0_outputs(2172) <= not (a or b);
    layer0_outputs(2173) <= a or b;
    layer0_outputs(2174) <= not b;
    layer0_outputs(2175) <= not (a and b);
    layer0_outputs(2176) <= a and not b;
    layer0_outputs(2177) <= '1';
    layer0_outputs(2178) <= not (a xor b);
    layer0_outputs(2179) <= not (a xor b);
    layer0_outputs(2180) <= b;
    layer0_outputs(2181) <= a and b;
    layer0_outputs(2182) <= not (a or b);
    layer0_outputs(2183) <= a xor b;
    layer0_outputs(2184) <= not (a or b);
    layer0_outputs(2185) <= a and not b;
    layer0_outputs(2186) <= a and b;
    layer0_outputs(2187) <= a xor b;
    layer0_outputs(2188) <= b;
    layer0_outputs(2189) <= a xor b;
    layer0_outputs(2190) <= not b;
    layer0_outputs(2191) <= a xor b;
    layer0_outputs(2192) <= a and b;
    layer0_outputs(2193) <= b and not a;
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= '1';
    layer0_outputs(2196) <= b and not a;
    layer0_outputs(2197) <= a;
    layer0_outputs(2198) <= a and not b;
    layer0_outputs(2199) <= '0';
    layer0_outputs(2200) <= not a;
    layer0_outputs(2201) <= b;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= not (a or b);
    layer0_outputs(2204) <= '0';
    layer0_outputs(2205) <= a and not b;
    layer0_outputs(2206) <= '0';
    layer0_outputs(2207) <= not (a or b);
    layer0_outputs(2208) <= b;
    layer0_outputs(2209) <= not a or b;
    layer0_outputs(2210) <= a and b;
    layer0_outputs(2211) <= not (a xor b);
    layer0_outputs(2212) <= a and b;
    layer0_outputs(2213) <= a or b;
    layer0_outputs(2214) <= not b;
    layer0_outputs(2215) <= a or b;
    layer0_outputs(2216) <= not a or b;
    layer0_outputs(2217) <= b;
    layer0_outputs(2218) <= not (a or b);
    layer0_outputs(2219) <= not b or a;
    layer0_outputs(2220) <= a or b;
    layer0_outputs(2221) <= not b;
    layer0_outputs(2222) <= not (a or b);
    layer0_outputs(2223) <= not a;
    layer0_outputs(2224) <= not (a or b);
    layer0_outputs(2225) <= '0';
    layer0_outputs(2226) <= a;
    layer0_outputs(2227) <= '1';
    layer0_outputs(2228) <= a and not b;
    layer0_outputs(2229) <= not (a or b);
    layer0_outputs(2230) <= a or b;
    layer0_outputs(2231) <= a xor b;
    layer0_outputs(2232) <= a and not b;
    layer0_outputs(2233) <= not (a xor b);
    layer0_outputs(2234) <= a;
    layer0_outputs(2235) <= not (a or b);
    layer0_outputs(2236) <= not b or a;
    layer0_outputs(2237) <= a xor b;
    layer0_outputs(2238) <= a xor b;
    layer0_outputs(2239) <= '1';
    layer0_outputs(2240) <= '1';
    layer0_outputs(2241) <= not a or b;
    layer0_outputs(2242) <= not (a xor b);
    layer0_outputs(2243) <= not a;
    layer0_outputs(2244) <= not (a or b);
    layer0_outputs(2245) <= a;
    layer0_outputs(2246) <= a and not b;
    layer0_outputs(2247) <= not b;
    layer0_outputs(2248) <= not a or b;
    layer0_outputs(2249) <= not a or b;
    layer0_outputs(2250) <= b;
    layer0_outputs(2251) <= a and b;
    layer0_outputs(2252) <= a and not b;
    layer0_outputs(2253) <= not (a or b);
    layer0_outputs(2254) <= not a;
    layer0_outputs(2255) <= not a or b;
    layer0_outputs(2256) <= b and not a;
    layer0_outputs(2257) <= not (a or b);
    layer0_outputs(2258) <= a or b;
    layer0_outputs(2259) <= not (a or b);
    layer0_outputs(2260) <= a xor b;
    layer0_outputs(2261) <= not a;
    layer0_outputs(2262) <= not (a or b);
    layer0_outputs(2263) <= not b;
    layer0_outputs(2264) <= b;
    layer0_outputs(2265) <= not a;
    layer0_outputs(2266) <= b;
    layer0_outputs(2267) <= b and not a;
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= a or b;
    layer0_outputs(2270) <= not (a or b);
    layer0_outputs(2271) <= not (a or b);
    layer0_outputs(2272) <= not (a and b);
    layer0_outputs(2273) <= not (a or b);
    layer0_outputs(2274) <= '1';
    layer0_outputs(2275) <= not b;
    layer0_outputs(2276) <= not a;
    layer0_outputs(2277) <= b;
    layer0_outputs(2278) <= not a;
    layer0_outputs(2279) <= not (a and b);
    layer0_outputs(2280) <= a or b;
    layer0_outputs(2281) <= b;
    layer0_outputs(2282) <= b and not a;
    layer0_outputs(2283) <= a or b;
    layer0_outputs(2284) <= '0';
    layer0_outputs(2285) <= a or b;
    layer0_outputs(2286) <= a or b;
    layer0_outputs(2287) <= not a or b;
    layer0_outputs(2288) <= a xor b;
    layer0_outputs(2289) <= not a;
    layer0_outputs(2290) <= not b;
    layer0_outputs(2291) <= a or b;
    layer0_outputs(2292) <= '1';
    layer0_outputs(2293) <= b and not a;
    layer0_outputs(2294) <= not a;
    layer0_outputs(2295) <= b and not a;
    layer0_outputs(2296) <= a;
    layer0_outputs(2297) <= not b or a;
    layer0_outputs(2298) <= not a or b;
    layer0_outputs(2299) <= b and not a;
    layer0_outputs(2300) <= not b;
    layer0_outputs(2301) <= not b;
    layer0_outputs(2302) <= not a or b;
    layer0_outputs(2303) <= a or b;
    layer0_outputs(2304) <= '0';
    layer0_outputs(2305) <= not (a and b);
    layer0_outputs(2306) <= not (a xor b);
    layer0_outputs(2307) <= b and not a;
    layer0_outputs(2308) <= not a or b;
    layer0_outputs(2309) <= not (a and b);
    layer0_outputs(2310) <= not b;
    layer0_outputs(2311) <= '1';
    layer0_outputs(2312) <= not (a or b);
    layer0_outputs(2313) <= a and b;
    layer0_outputs(2314) <= '1';
    layer0_outputs(2315) <= not (a or b);
    layer0_outputs(2316) <= b and not a;
    layer0_outputs(2317) <= not (a or b);
    layer0_outputs(2318) <= not b or a;
    layer0_outputs(2319) <= a and not b;
    layer0_outputs(2320) <= a and not b;
    layer0_outputs(2321) <= not (a or b);
    layer0_outputs(2322) <= not (a or b);
    layer0_outputs(2323) <= not b;
    layer0_outputs(2324) <= a or b;
    layer0_outputs(2325) <= a xor b;
    layer0_outputs(2326) <= not (a or b);
    layer0_outputs(2327) <= '1';
    layer0_outputs(2328) <= a xor b;
    layer0_outputs(2329) <= b;
    layer0_outputs(2330) <= not a;
    layer0_outputs(2331) <= not (a or b);
    layer0_outputs(2332) <= b;
    layer0_outputs(2333) <= not a or b;
    layer0_outputs(2334) <= not b;
    layer0_outputs(2335) <= not a or b;
    layer0_outputs(2336) <= b;
    layer0_outputs(2337) <= not b or a;
    layer0_outputs(2338) <= a xor b;
    layer0_outputs(2339) <= a or b;
    layer0_outputs(2340) <= a or b;
    layer0_outputs(2341) <= a and b;
    layer0_outputs(2342) <= '1';
    layer0_outputs(2343) <= not (a or b);
    layer0_outputs(2344) <= '0';
    layer0_outputs(2345) <= not a or b;
    layer0_outputs(2346) <= not (a xor b);
    layer0_outputs(2347) <= not (a xor b);
    layer0_outputs(2348) <= a and not b;
    layer0_outputs(2349) <= not b;
    layer0_outputs(2350) <= not b or a;
    layer0_outputs(2351) <= a;
    layer0_outputs(2352) <= '1';
    layer0_outputs(2353) <= not b;
    layer0_outputs(2354) <= b and not a;
    layer0_outputs(2355) <= not (a or b);
    layer0_outputs(2356) <= a or b;
    layer0_outputs(2357) <= a xor b;
    layer0_outputs(2358) <= not (a xor b);
    layer0_outputs(2359) <= a or b;
    layer0_outputs(2360) <= a and b;
    layer0_outputs(2361) <= b;
    layer0_outputs(2362) <= a xor b;
    layer0_outputs(2363) <= a or b;
    layer0_outputs(2364) <= not (a xor b);
    layer0_outputs(2365) <= not (a xor b);
    layer0_outputs(2366) <= not (a xor b);
    layer0_outputs(2367) <= a or b;
    layer0_outputs(2368) <= '1';
    layer0_outputs(2369) <= not b;
    layer0_outputs(2370) <= not b;
    layer0_outputs(2371) <= b and not a;
    layer0_outputs(2372) <= not (a or b);
    layer0_outputs(2373) <= a and not b;
    layer0_outputs(2374) <= a;
    layer0_outputs(2375) <= a or b;
    layer0_outputs(2376) <= b;
    layer0_outputs(2377) <= not (a xor b);
    layer0_outputs(2378) <= not b or a;
    layer0_outputs(2379) <= not (a xor b);
    layer0_outputs(2380) <= not b;
    layer0_outputs(2381) <= not a or b;
    layer0_outputs(2382) <= a or b;
    layer0_outputs(2383) <= not a or b;
    layer0_outputs(2384) <= a;
    layer0_outputs(2385) <= a xor b;
    layer0_outputs(2386) <= not a;
    layer0_outputs(2387) <= a or b;
    layer0_outputs(2388) <= a and not b;
    layer0_outputs(2389) <= b;
    layer0_outputs(2390) <= a;
    layer0_outputs(2391) <= a xor b;
    layer0_outputs(2392) <= a xor b;
    layer0_outputs(2393) <= a;
    layer0_outputs(2394) <= '1';
    layer0_outputs(2395) <= not (a or b);
    layer0_outputs(2396) <= a xor b;
    layer0_outputs(2397) <= b;
    layer0_outputs(2398) <= a or b;
    layer0_outputs(2399) <= b;
    layer0_outputs(2400) <= '1';
    layer0_outputs(2401) <= a and not b;
    layer0_outputs(2402) <= a and not b;
    layer0_outputs(2403) <= a and not b;
    layer0_outputs(2404) <= not a;
    layer0_outputs(2405) <= b;
    layer0_outputs(2406) <= not (a xor b);
    layer0_outputs(2407) <= not b or a;
    layer0_outputs(2408) <= a and not b;
    layer0_outputs(2409) <= not a;
    layer0_outputs(2410) <= not (a or b);
    layer0_outputs(2411) <= not b or a;
    layer0_outputs(2412) <= '1';
    layer0_outputs(2413) <= not b or a;
    layer0_outputs(2414) <= not a;
    layer0_outputs(2415) <= a xor b;
    layer0_outputs(2416) <= not b;
    layer0_outputs(2417) <= a;
    layer0_outputs(2418) <= not (a and b);
    layer0_outputs(2419) <= not a or b;
    layer0_outputs(2420) <= not b;
    layer0_outputs(2421) <= not b;
    layer0_outputs(2422) <= not a;
    layer0_outputs(2423) <= a xor b;
    layer0_outputs(2424) <= not b;
    layer0_outputs(2425) <= a xor b;
    layer0_outputs(2426) <= a;
    layer0_outputs(2427) <= a;
    layer0_outputs(2428) <= not b or a;
    layer0_outputs(2429) <= a or b;
    layer0_outputs(2430) <= a and not b;
    layer0_outputs(2431) <= not a or b;
    layer0_outputs(2432) <= not a;
    layer0_outputs(2433) <= not (a xor b);
    layer0_outputs(2434) <= a or b;
    layer0_outputs(2435) <= a or b;
    layer0_outputs(2436) <= not b or a;
    layer0_outputs(2437) <= '1';
    layer0_outputs(2438) <= '0';
    layer0_outputs(2439) <= b and not a;
    layer0_outputs(2440) <= a;
    layer0_outputs(2441) <= a;
    layer0_outputs(2442) <= a or b;
    layer0_outputs(2443) <= not a;
    layer0_outputs(2444) <= not b;
    layer0_outputs(2445) <= not (a xor b);
    layer0_outputs(2446) <= b and not a;
    layer0_outputs(2447) <= not a or b;
    layer0_outputs(2448) <= not (a xor b);
    layer0_outputs(2449) <= a and b;
    layer0_outputs(2450) <= not (a or b);
    layer0_outputs(2451) <= b;
    layer0_outputs(2452) <= not a;
    layer0_outputs(2453) <= b and not a;
    layer0_outputs(2454) <= a and not b;
    layer0_outputs(2455) <= not b or a;
    layer0_outputs(2456) <= not (a or b);
    layer0_outputs(2457) <= a or b;
    layer0_outputs(2458) <= b and not a;
    layer0_outputs(2459) <= not (a xor b);
    layer0_outputs(2460) <= b and not a;
    layer0_outputs(2461) <= a;
    layer0_outputs(2462) <= not (a or b);
    layer0_outputs(2463) <= not (a or b);
    layer0_outputs(2464) <= a or b;
    layer0_outputs(2465) <= not (a and b);
    layer0_outputs(2466) <= not (a xor b);
    layer0_outputs(2467) <= a or b;
    layer0_outputs(2468) <= not (a or b);
    layer0_outputs(2469) <= '1';
    layer0_outputs(2470) <= b;
    layer0_outputs(2471) <= not a;
    layer0_outputs(2472) <= '0';
    layer0_outputs(2473) <= b;
    layer0_outputs(2474) <= not (a xor b);
    layer0_outputs(2475) <= not a;
    layer0_outputs(2476) <= a and not b;
    layer0_outputs(2477) <= a xor b;
    layer0_outputs(2478) <= b and not a;
    layer0_outputs(2479) <= a xor b;
    layer0_outputs(2480) <= not a;
    layer0_outputs(2481) <= a;
    layer0_outputs(2482) <= a or b;
    layer0_outputs(2483) <= a or b;
    layer0_outputs(2484) <= a;
    layer0_outputs(2485) <= a;
    layer0_outputs(2486) <= a or b;
    layer0_outputs(2487) <= a xor b;
    layer0_outputs(2488) <= a or b;
    layer0_outputs(2489) <= not a or b;
    layer0_outputs(2490) <= not b;
    layer0_outputs(2491) <= not (a or b);
    layer0_outputs(2492) <= not (a and b);
    layer0_outputs(2493) <= not b or a;
    layer0_outputs(2494) <= not a or b;
    layer0_outputs(2495) <= a xor b;
    layer0_outputs(2496) <= a or b;
    layer0_outputs(2497) <= not a;
    layer0_outputs(2498) <= a and not b;
    layer0_outputs(2499) <= not (a or b);
    layer0_outputs(2500) <= not (a or b);
    layer0_outputs(2501) <= b;
    layer0_outputs(2502) <= a and not b;
    layer0_outputs(2503) <= not a or b;
    layer0_outputs(2504) <= '0';
    layer0_outputs(2505) <= not a;
    layer0_outputs(2506) <= a xor b;
    layer0_outputs(2507) <= not a;
    layer0_outputs(2508) <= b and not a;
    layer0_outputs(2509) <= not (a or b);
    layer0_outputs(2510) <= not (a or b);
    layer0_outputs(2511) <= b and not a;
    layer0_outputs(2512) <= not a or b;
    layer0_outputs(2513) <= not (a or b);
    layer0_outputs(2514) <= b;
    layer0_outputs(2515) <= '1';
    layer0_outputs(2516) <= b;
    layer0_outputs(2517) <= not a;
    layer0_outputs(2518) <= a;
    layer0_outputs(2519) <= '1';
    layer0_outputs(2520) <= '0';
    layer0_outputs(2521) <= a;
    layer0_outputs(2522) <= a and not b;
    layer0_outputs(2523) <= '1';
    layer0_outputs(2524) <= not b;
    layer0_outputs(2525) <= not a;
    layer0_outputs(2526) <= a or b;
    layer0_outputs(2527) <= b and not a;
    layer0_outputs(2528) <= '0';
    layer0_outputs(2529) <= not a or b;
    layer0_outputs(2530) <= b;
    layer0_outputs(2531) <= '0';
    layer0_outputs(2532) <= a or b;
    layer0_outputs(2533) <= a and b;
    layer0_outputs(2534) <= a and b;
    layer0_outputs(2535) <= b;
    layer0_outputs(2536) <= a or b;
    layer0_outputs(2537) <= not a;
    layer0_outputs(2538) <= b and not a;
    layer0_outputs(2539) <= not (a or b);
    layer0_outputs(2540) <= not (a or b);
    layer0_outputs(2541) <= a or b;
    layer0_outputs(2542) <= b and not a;
    layer0_outputs(2543) <= a or b;
    layer0_outputs(2544) <= '1';
    layer0_outputs(2545) <= b;
    layer0_outputs(2546) <= a;
    layer0_outputs(2547) <= not b;
    layer0_outputs(2548) <= '0';
    layer0_outputs(2549) <= not (a xor b);
    layer0_outputs(2550) <= a or b;
    layer0_outputs(2551) <= a and b;
    layer0_outputs(2552) <= not a;
    layer0_outputs(2553) <= not b or a;
    layer0_outputs(2554) <= a xor b;
    layer0_outputs(2555) <= not (a or b);
    layer0_outputs(2556) <= a;
    layer0_outputs(2557) <= a xor b;
    layer0_outputs(2558) <= a xor b;
    layer0_outputs(2559) <= not (a or b);
    layer0_outputs(2560) <= not (a xor b);
    layer0_outputs(2561) <= not a or b;
    layer0_outputs(2562) <= not a;
    layer0_outputs(2563) <= '0';
    layer0_outputs(2564) <= '0';
    layer0_outputs(2565) <= not a or b;
    layer0_outputs(2566) <= not a or b;
    layer0_outputs(2567) <= b and not a;
    layer0_outputs(2568) <= not b or a;
    layer0_outputs(2569) <= a and not b;
    layer0_outputs(2570) <= not b or a;
    layer0_outputs(2571) <= not a or b;
    layer0_outputs(2572) <= a or b;
    layer0_outputs(2573) <= not b or a;
    layer0_outputs(2574) <= not (a and b);
    layer0_outputs(2575) <= a;
    layer0_outputs(2576) <= not b or a;
    layer0_outputs(2577) <= a;
    layer0_outputs(2578) <= a or b;
    layer0_outputs(2579) <= a and b;
    layer0_outputs(2580) <= b;
    layer0_outputs(2581) <= a or b;
    layer0_outputs(2582) <= not b or a;
    layer0_outputs(2583) <= b and not a;
    layer0_outputs(2584) <= b;
    layer0_outputs(2585) <= a or b;
    layer0_outputs(2586) <= not a or b;
    layer0_outputs(2587) <= a and b;
    layer0_outputs(2588) <= a xor b;
    layer0_outputs(2589) <= not a;
    layer0_outputs(2590) <= not b or a;
    layer0_outputs(2591) <= not b or a;
    layer0_outputs(2592) <= b and not a;
    layer0_outputs(2593) <= not (a or b);
    layer0_outputs(2594) <= not b;
    layer0_outputs(2595) <= not a;
    layer0_outputs(2596) <= a xor b;
    layer0_outputs(2597) <= not a;
    layer0_outputs(2598) <= not (a and b);
    layer0_outputs(2599) <= not (a and b);
    layer0_outputs(2600) <= a or b;
    layer0_outputs(2601) <= not b;
    layer0_outputs(2602) <= not b;
    layer0_outputs(2603) <= not (a xor b);
    layer0_outputs(2604) <= b;
    layer0_outputs(2605) <= a and b;
    layer0_outputs(2606) <= a or b;
    layer0_outputs(2607) <= not (a xor b);
    layer0_outputs(2608) <= not (a xor b);
    layer0_outputs(2609) <= not (a and b);
    layer0_outputs(2610) <= a xor b;
    layer0_outputs(2611) <= a or b;
    layer0_outputs(2612) <= '1';
    layer0_outputs(2613) <= a or b;
    layer0_outputs(2614) <= a and b;
    layer0_outputs(2615) <= '0';
    layer0_outputs(2616) <= not (a or b);
    layer0_outputs(2617) <= not (a and b);
    layer0_outputs(2618) <= a;
    layer0_outputs(2619) <= b and not a;
    layer0_outputs(2620) <= a;
    layer0_outputs(2621) <= a;
    layer0_outputs(2622) <= a xor b;
    layer0_outputs(2623) <= '0';
    layer0_outputs(2624) <= not (a or b);
    layer0_outputs(2625) <= not a;
    layer0_outputs(2626) <= a;
    layer0_outputs(2627) <= not b;
    layer0_outputs(2628) <= not b;
    layer0_outputs(2629) <= not (a xor b);
    layer0_outputs(2630) <= not (a xor b);
    layer0_outputs(2631) <= not (a xor b);
    layer0_outputs(2632) <= a;
    layer0_outputs(2633) <= b and not a;
    layer0_outputs(2634) <= a or b;
    layer0_outputs(2635) <= a and not b;
    layer0_outputs(2636) <= a and b;
    layer0_outputs(2637) <= a or b;
    layer0_outputs(2638) <= a;
    layer0_outputs(2639) <= not a;
    layer0_outputs(2640) <= b;
    layer0_outputs(2641) <= not a or b;
    layer0_outputs(2642) <= a and b;
    layer0_outputs(2643) <= a or b;
    layer0_outputs(2644) <= b;
    layer0_outputs(2645) <= not b or a;
    layer0_outputs(2646) <= a;
    layer0_outputs(2647) <= not b;
    layer0_outputs(2648) <= a xor b;
    layer0_outputs(2649) <= not (a or b);
    layer0_outputs(2650) <= not (a xor b);
    layer0_outputs(2651) <= '1';
    layer0_outputs(2652) <= not (a or b);
    layer0_outputs(2653) <= not a or b;
    layer0_outputs(2654) <= not a or b;
    layer0_outputs(2655) <= a;
    layer0_outputs(2656) <= b and not a;
    layer0_outputs(2657) <= not a;
    layer0_outputs(2658) <= '0';
    layer0_outputs(2659) <= not b or a;
    layer0_outputs(2660) <= a or b;
    layer0_outputs(2661) <= not (a and b);
    layer0_outputs(2662) <= not a;
    layer0_outputs(2663) <= not (a or b);
    layer0_outputs(2664) <= not b;
    layer0_outputs(2665) <= a xor b;
    layer0_outputs(2666) <= not (a xor b);
    layer0_outputs(2667) <= '1';
    layer0_outputs(2668) <= b;
    layer0_outputs(2669) <= a or b;
    layer0_outputs(2670) <= a;
    layer0_outputs(2671) <= a and not b;
    layer0_outputs(2672) <= not a;
    layer0_outputs(2673) <= a and not b;
    layer0_outputs(2674) <= not a;
    layer0_outputs(2675) <= a and not b;
    layer0_outputs(2676) <= a or b;
    layer0_outputs(2677) <= '0';
    layer0_outputs(2678) <= a or b;
    layer0_outputs(2679) <= a;
    layer0_outputs(2680) <= not (a or b);
    layer0_outputs(2681) <= a xor b;
    layer0_outputs(2682) <= a;
    layer0_outputs(2683) <= '1';
    layer0_outputs(2684) <= a and b;
    layer0_outputs(2685) <= not b or a;
    layer0_outputs(2686) <= b and not a;
    layer0_outputs(2687) <= not (a or b);
    layer0_outputs(2688) <= not (a or b);
    layer0_outputs(2689) <= not (a or b);
    layer0_outputs(2690) <= not (a or b);
    layer0_outputs(2691) <= b and not a;
    layer0_outputs(2692) <= not a;
    layer0_outputs(2693) <= '1';
    layer0_outputs(2694) <= '0';
    layer0_outputs(2695) <= not a or b;
    layer0_outputs(2696) <= not a;
    layer0_outputs(2697) <= not (a xor b);
    layer0_outputs(2698) <= '0';
    layer0_outputs(2699) <= not a;
    layer0_outputs(2700) <= '1';
    layer0_outputs(2701) <= '1';
    layer0_outputs(2702) <= not (a or b);
    layer0_outputs(2703) <= not a;
    layer0_outputs(2704) <= a and b;
    layer0_outputs(2705) <= not (a or b);
    layer0_outputs(2706) <= a;
    layer0_outputs(2707) <= a or b;
    layer0_outputs(2708) <= not (a xor b);
    layer0_outputs(2709) <= a and b;
    layer0_outputs(2710) <= not a;
    layer0_outputs(2711) <= a or b;
    layer0_outputs(2712) <= a;
    layer0_outputs(2713) <= a;
    layer0_outputs(2714) <= not b;
    layer0_outputs(2715) <= not a or b;
    layer0_outputs(2716) <= not (a xor b);
    layer0_outputs(2717) <= not (a or b);
    layer0_outputs(2718) <= '1';
    layer0_outputs(2719) <= '1';
    layer0_outputs(2720) <= not a;
    layer0_outputs(2721) <= not a;
    layer0_outputs(2722) <= not a;
    layer0_outputs(2723) <= not b or a;
    layer0_outputs(2724) <= a and not b;
    layer0_outputs(2725) <= not a or b;
    layer0_outputs(2726) <= b;
    layer0_outputs(2727) <= '0';
    layer0_outputs(2728) <= b and not a;
    layer0_outputs(2729) <= b and not a;
    layer0_outputs(2730) <= '1';
    layer0_outputs(2731) <= not (a or b);
    layer0_outputs(2732) <= b;
    layer0_outputs(2733) <= not a;
    layer0_outputs(2734) <= b;
    layer0_outputs(2735) <= b and not a;
    layer0_outputs(2736) <= not a;
    layer0_outputs(2737) <= a or b;
    layer0_outputs(2738) <= b;
    layer0_outputs(2739) <= a;
    layer0_outputs(2740) <= not a;
    layer0_outputs(2741) <= not b;
    layer0_outputs(2742) <= a;
    layer0_outputs(2743) <= b and not a;
    layer0_outputs(2744) <= a and not b;
    layer0_outputs(2745) <= not (a and b);
    layer0_outputs(2746) <= not b or a;
    layer0_outputs(2747) <= a xor b;
    layer0_outputs(2748) <= a;
    layer0_outputs(2749) <= not (a or b);
    layer0_outputs(2750) <= not b or a;
    layer0_outputs(2751) <= b;
    layer0_outputs(2752) <= not b;
    layer0_outputs(2753) <= not (a or b);
    layer0_outputs(2754) <= b and not a;
    layer0_outputs(2755) <= b;
    layer0_outputs(2756) <= not b;
    layer0_outputs(2757) <= b and not a;
    layer0_outputs(2758) <= '1';
    layer0_outputs(2759) <= not a;
    layer0_outputs(2760) <= a;
    layer0_outputs(2761) <= b;
    layer0_outputs(2762) <= not a or b;
    layer0_outputs(2763) <= not a or b;
    layer0_outputs(2764) <= not a or b;
    layer0_outputs(2765) <= not (a or b);
    layer0_outputs(2766) <= b;
    layer0_outputs(2767) <= not (a or b);
    layer0_outputs(2768) <= not a;
    layer0_outputs(2769) <= b;
    layer0_outputs(2770) <= a and b;
    layer0_outputs(2771) <= b and not a;
    layer0_outputs(2772) <= a and not b;
    layer0_outputs(2773) <= not b;
    layer0_outputs(2774) <= a;
    layer0_outputs(2775) <= a or b;
    layer0_outputs(2776) <= not b;
    layer0_outputs(2777) <= a and b;
    layer0_outputs(2778) <= not (a or b);
    layer0_outputs(2779) <= not a;
    layer0_outputs(2780) <= b and not a;
    layer0_outputs(2781) <= not (a or b);
    layer0_outputs(2782) <= '0';
    layer0_outputs(2783) <= '1';
    layer0_outputs(2784) <= a or b;
    layer0_outputs(2785) <= not a;
    layer0_outputs(2786) <= not b;
    layer0_outputs(2787) <= not (a or b);
    layer0_outputs(2788) <= not b or a;
    layer0_outputs(2789) <= not b or a;
    layer0_outputs(2790) <= not b or a;
    layer0_outputs(2791) <= a and not b;
    layer0_outputs(2792) <= b;
    layer0_outputs(2793) <= not b;
    layer0_outputs(2794) <= not (a and b);
    layer0_outputs(2795) <= a and not b;
    layer0_outputs(2796) <= not b;
    layer0_outputs(2797) <= b;
    layer0_outputs(2798) <= '1';
    layer0_outputs(2799) <= not b;
    layer0_outputs(2800) <= a or b;
    layer0_outputs(2801) <= not (a xor b);
    layer0_outputs(2802) <= not (a and b);
    layer0_outputs(2803) <= not b or a;
    layer0_outputs(2804) <= not a or b;
    layer0_outputs(2805) <= a or b;
    layer0_outputs(2806) <= not (a or b);
    layer0_outputs(2807) <= not b;
    layer0_outputs(2808) <= not (a or b);
    layer0_outputs(2809) <= a or b;
    layer0_outputs(2810) <= a;
    layer0_outputs(2811) <= a;
    layer0_outputs(2812) <= '1';
    layer0_outputs(2813) <= a or b;
    layer0_outputs(2814) <= not (a or b);
    layer0_outputs(2815) <= b;
    layer0_outputs(2816) <= not a;
    layer0_outputs(2817) <= b;
    layer0_outputs(2818) <= a xor b;
    layer0_outputs(2819) <= a;
    layer0_outputs(2820) <= not (a xor b);
    layer0_outputs(2821) <= not (a and b);
    layer0_outputs(2822) <= not (a or b);
    layer0_outputs(2823) <= not (a or b);
    layer0_outputs(2824) <= not b;
    layer0_outputs(2825) <= a;
    layer0_outputs(2826) <= a xor b;
    layer0_outputs(2827) <= not a or b;
    layer0_outputs(2828) <= a or b;
    layer0_outputs(2829) <= not b or a;
    layer0_outputs(2830) <= b;
    layer0_outputs(2831) <= not (a xor b);
    layer0_outputs(2832) <= b;
    layer0_outputs(2833) <= a and b;
    layer0_outputs(2834) <= b and not a;
    layer0_outputs(2835) <= a or b;
    layer0_outputs(2836) <= not (a or b);
    layer0_outputs(2837) <= a or b;
    layer0_outputs(2838) <= not (a or b);
    layer0_outputs(2839) <= not (a or b);
    layer0_outputs(2840) <= not b or a;
    layer0_outputs(2841) <= not a;
    layer0_outputs(2842) <= a and not b;
    layer0_outputs(2843) <= not a;
    layer0_outputs(2844) <= not a or b;
    layer0_outputs(2845) <= not a or b;
    layer0_outputs(2846) <= not a;
    layer0_outputs(2847) <= a or b;
    layer0_outputs(2848) <= a;
    layer0_outputs(2849) <= a;
    layer0_outputs(2850) <= '0';
    layer0_outputs(2851) <= not (a xor b);
    layer0_outputs(2852) <= a and b;
    layer0_outputs(2853) <= b;
    layer0_outputs(2854) <= b and not a;
    layer0_outputs(2855) <= not (a xor b);
    layer0_outputs(2856) <= b;
    layer0_outputs(2857) <= a and not b;
    layer0_outputs(2858) <= not (a or b);
    layer0_outputs(2859) <= b;
    layer0_outputs(2860) <= a or b;
    layer0_outputs(2861) <= '1';
    layer0_outputs(2862) <= a and not b;
    layer0_outputs(2863) <= a or b;
    layer0_outputs(2864) <= not (a xor b);
    layer0_outputs(2865) <= a and not b;
    layer0_outputs(2866) <= a xor b;
    layer0_outputs(2867) <= a or b;
    layer0_outputs(2868) <= a xor b;
    layer0_outputs(2869) <= not a;
    layer0_outputs(2870) <= not (a and b);
    layer0_outputs(2871) <= not b;
    layer0_outputs(2872) <= not a;
    layer0_outputs(2873) <= a and b;
    layer0_outputs(2874) <= b;
    layer0_outputs(2875) <= not b;
    layer0_outputs(2876) <= b;
    layer0_outputs(2877) <= a and b;
    layer0_outputs(2878) <= a or b;
    layer0_outputs(2879) <= a xor b;
    layer0_outputs(2880) <= not (a or b);
    layer0_outputs(2881) <= b and not a;
    layer0_outputs(2882) <= '0';
    layer0_outputs(2883) <= a;
    layer0_outputs(2884) <= a xor b;
    layer0_outputs(2885) <= not (a or b);
    layer0_outputs(2886) <= not b;
    layer0_outputs(2887) <= b and not a;
    layer0_outputs(2888) <= not (a and b);
    layer0_outputs(2889) <= not (a xor b);
    layer0_outputs(2890) <= '0';
    layer0_outputs(2891) <= not a;
    layer0_outputs(2892) <= not (a xor b);
    layer0_outputs(2893) <= '0';
    layer0_outputs(2894) <= not (a xor b);
    layer0_outputs(2895) <= not (a or b);
    layer0_outputs(2896) <= a or b;
    layer0_outputs(2897) <= not (a xor b);
    layer0_outputs(2898) <= not (a and b);
    layer0_outputs(2899) <= not b or a;
    layer0_outputs(2900) <= a or b;
    layer0_outputs(2901) <= b and not a;
    layer0_outputs(2902) <= a or b;
    layer0_outputs(2903) <= a and b;
    layer0_outputs(2904) <= b and not a;
    layer0_outputs(2905) <= a or b;
    layer0_outputs(2906) <= b;
    layer0_outputs(2907) <= not b;
    layer0_outputs(2908) <= a or b;
    layer0_outputs(2909) <= not (a xor b);
    layer0_outputs(2910) <= '0';
    layer0_outputs(2911) <= a or b;
    layer0_outputs(2912) <= '1';
    layer0_outputs(2913) <= a or b;
    layer0_outputs(2914) <= '1';
    layer0_outputs(2915) <= not b or a;
    layer0_outputs(2916) <= not (a or b);
    layer0_outputs(2917) <= not a;
    layer0_outputs(2918) <= not b or a;
    layer0_outputs(2919) <= not a or b;
    layer0_outputs(2920) <= a and b;
    layer0_outputs(2921) <= not a or b;
    layer0_outputs(2922) <= b;
    layer0_outputs(2923) <= a or b;
    layer0_outputs(2924) <= a xor b;
    layer0_outputs(2925) <= a or b;
    layer0_outputs(2926) <= a or b;
    layer0_outputs(2927) <= not b or a;
    layer0_outputs(2928) <= not a or b;
    layer0_outputs(2929) <= a or b;
    layer0_outputs(2930) <= a or b;
    layer0_outputs(2931) <= not (a xor b);
    layer0_outputs(2932) <= a;
    layer0_outputs(2933) <= not (a or b);
    layer0_outputs(2934) <= not a or b;
    layer0_outputs(2935) <= a and not b;
    layer0_outputs(2936) <= a;
    layer0_outputs(2937) <= b;
    layer0_outputs(2938) <= not b;
    layer0_outputs(2939) <= a or b;
    layer0_outputs(2940) <= not (a xor b);
    layer0_outputs(2941) <= not (a and b);
    layer0_outputs(2942) <= '0';
    layer0_outputs(2943) <= a or b;
    layer0_outputs(2944) <= not a;
    layer0_outputs(2945) <= not a;
    layer0_outputs(2946) <= not a;
    layer0_outputs(2947) <= '0';
    layer0_outputs(2948) <= a xor b;
    layer0_outputs(2949) <= not (a or b);
    layer0_outputs(2950) <= a;
    layer0_outputs(2951) <= not (a or b);
    layer0_outputs(2952) <= not (a or b);
    layer0_outputs(2953) <= '0';
    layer0_outputs(2954) <= b and not a;
    layer0_outputs(2955) <= not (a xor b);
    layer0_outputs(2956) <= not b;
    layer0_outputs(2957) <= b and not a;
    layer0_outputs(2958) <= '1';
    layer0_outputs(2959) <= a and b;
    layer0_outputs(2960) <= not (a xor b);
    layer0_outputs(2961) <= b;
    layer0_outputs(2962) <= not a;
    layer0_outputs(2963) <= not (a and b);
    layer0_outputs(2964) <= not b or a;
    layer0_outputs(2965) <= not (a and b);
    layer0_outputs(2966) <= not (a xor b);
    layer0_outputs(2967) <= a and b;
    layer0_outputs(2968) <= a and b;
    layer0_outputs(2969) <= b;
    layer0_outputs(2970) <= not b;
    layer0_outputs(2971) <= not a;
    layer0_outputs(2972) <= not b;
    layer0_outputs(2973) <= a and b;
    layer0_outputs(2974) <= not b or a;
    layer0_outputs(2975) <= a or b;
    layer0_outputs(2976) <= not (a or b);
    layer0_outputs(2977) <= not b or a;
    layer0_outputs(2978) <= a and b;
    layer0_outputs(2979) <= b and not a;
    layer0_outputs(2980) <= b and not a;
    layer0_outputs(2981) <= not (a or b);
    layer0_outputs(2982) <= a;
    layer0_outputs(2983) <= a xor b;
    layer0_outputs(2984) <= a xor b;
    layer0_outputs(2985) <= b;
    layer0_outputs(2986) <= not a;
    layer0_outputs(2987) <= b;
    layer0_outputs(2988) <= not b;
    layer0_outputs(2989) <= not (a and b);
    layer0_outputs(2990) <= not a or b;
    layer0_outputs(2991) <= not (a xor b);
    layer0_outputs(2992) <= not b or a;
    layer0_outputs(2993) <= b and not a;
    layer0_outputs(2994) <= b and not a;
    layer0_outputs(2995) <= '0';
    layer0_outputs(2996) <= '1';
    layer0_outputs(2997) <= a;
    layer0_outputs(2998) <= b and not a;
    layer0_outputs(2999) <= not a or b;
    layer0_outputs(3000) <= not a or b;
    layer0_outputs(3001) <= b;
    layer0_outputs(3002) <= b;
    layer0_outputs(3003) <= '0';
    layer0_outputs(3004) <= not (a xor b);
    layer0_outputs(3005) <= not b;
    layer0_outputs(3006) <= not (a xor b);
    layer0_outputs(3007) <= b;
    layer0_outputs(3008) <= a;
    layer0_outputs(3009) <= b;
    layer0_outputs(3010) <= not a;
    layer0_outputs(3011) <= '0';
    layer0_outputs(3012) <= not a or b;
    layer0_outputs(3013) <= not (a or b);
    layer0_outputs(3014) <= b and not a;
    layer0_outputs(3015) <= not b or a;
    layer0_outputs(3016) <= a or b;
    layer0_outputs(3017) <= not (a or b);
    layer0_outputs(3018) <= not b or a;
    layer0_outputs(3019) <= not a or b;
    layer0_outputs(3020) <= b;
    layer0_outputs(3021) <= not a;
    layer0_outputs(3022) <= a;
    layer0_outputs(3023) <= not (a and b);
    layer0_outputs(3024) <= a or b;
    layer0_outputs(3025) <= not a or b;
    layer0_outputs(3026) <= not (a or b);
    layer0_outputs(3027) <= a or b;
    layer0_outputs(3028) <= a or b;
    layer0_outputs(3029) <= b and not a;
    layer0_outputs(3030) <= not (a and b);
    layer0_outputs(3031) <= not a or b;
    layer0_outputs(3032) <= not (a xor b);
    layer0_outputs(3033) <= a;
    layer0_outputs(3034) <= not (a or b);
    layer0_outputs(3035) <= a or b;
    layer0_outputs(3036) <= b;
    layer0_outputs(3037) <= a and b;
    layer0_outputs(3038) <= not (a xor b);
    layer0_outputs(3039) <= a or b;
    layer0_outputs(3040) <= not b or a;
    layer0_outputs(3041) <= not b or a;
    layer0_outputs(3042) <= not (a xor b);
    layer0_outputs(3043) <= not a or b;
    layer0_outputs(3044) <= a and not b;
    layer0_outputs(3045) <= not b;
    layer0_outputs(3046) <= a or b;
    layer0_outputs(3047) <= '0';
    layer0_outputs(3048) <= not a;
    layer0_outputs(3049) <= a and not b;
    layer0_outputs(3050) <= not a;
    layer0_outputs(3051) <= not b;
    layer0_outputs(3052) <= a or b;
    layer0_outputs(3053) <= b;
    layer0_outputs(3054) <= a or b;
    layer0_outputs(3055) <= not (a or b);
    layer0_outputs(3056) <= not (a or b);
    layer0_outputs(3057) <= not (a and b);
    layer0_outputs(3058) <= not b;
    layer0_outputs(3059) <= a and not b;
    layer0_outputs(3060) <= a;
    layer0_outputs(3061) <= not a or b;
    layer0_outputs(3062) <= not (a xor b);
    layer0_outputs(3063) <= '1';
    layer0_outputs(3064) <= a or b;
    layer0_outputs(3065) <= not (a or b);
    layer0_outputs(3066) <= a;
    layer0_outputs(3067) <= b;
    layer0_outputs(3068) <= not a or b;
    layer0_outputs(3069) <= not (a or b);
    layer0_outputs(3070) <= not b;
    layer0_outputs(3071) <= not (a or b);
    layer0_outputs(3072) <= a xor b;
    layer0_outputs(3073) <= a or b;
    layer0_outputs(3074) <= not (a or b);
    layer0_outputs(3075) <= not (a xor b);
    layer0_outputs(3076) <= not (a xor b);
    layer0_outputs(3077) <= a or b;
    layer0_outputs(3078) <= not a;
    layer0_outputs(3079) <= a xor b;
    layer0_outputs(3080) <= a or b;
    layer0_outputs(3081) <= a and b;
    layer0_outputs(3082) <= a;
    layer0_outputs(3083) <= a xor b;
    layer0_outputs(3084) <= not b;
    layer0_outputs(3085) <= a or b;
    layer0_outputs(3086) <= b;
    layer0_outputs(3087) <= b and not a;
    layer0_outputs(3088) <= not b or a;
    layer0_outputs(3089) <= b;
    layer0_outputs(3090) <= '1';
    layer0_outputs(3091) <= a and b;
    layer0_outputs(3092) <= a;
    layer0_outputs(3093) <= a or b;
    layer0_outputs(3094) <= a or b;
    layer0_outputs(3095) <= a or b;
    layer0_outputs(3096) <= b and not a;
    layer0_outputs(3097) <= not b;
    layer0_outputs(3098) <= not (a xor b);
    layer0_outputs(3099) <= a and b;
    layer0_outputs(3100) <= a xor b;
    layer0_outputs(3101) <= b;
    layer0_outputs(3102) <= b and not a;
    layer0_outputs(3103) <= a;
    layer0_outputs(3104) <= a and not b;
    layer0_outputs(3105) <= not (a xor b);
    layer0_outputs(3106) <= a;
    layer0_outputs(3107) <= not a;
    layer0_outputs(3108) <= not a or b;
    layer0_outputs(3109) <= not (a or b);
    layer0_outputs(3110) <= b;
    layer0_outputs(3111) <= not (a or b);
    layer0_outputs(3112) <= not a or b;
    layer0_outputs(3113) <= a or b;
    layer0_outputs(3114) <= a or b;
    layer0_outputs(3115) <= not a;
    layer0_outputs(3116) <= '1';
    layer0_outputs(3117) <= '1';
    layer0_outputs(3118) <= not (a xor b);
    layer0_outputs(3119) <= a or b;
    layer0_outputs(3120) <= '1';
    layer0_outputs(3121) <= a xor b;
    layer0_outputs(3122) <= b;
    layer0_outputs(3123) <= not (a or b);
    layer0_outputs(3124) <= not (a xor b);
    layer0_outputs(3125) <= not a;
    layer0_outputs(3126) <= a;
    layer0_outputs(3127) <= not a;
    layer0_outputs(3128) <= a;
    layer0_outputs(3129) <= '1';
    layer0_outputs(3130) <= not (a or b);
    layer0_outputs(3131) <= b;
    layer0_outputs(3132) <= not (a or b);
    layer0_outputs(3133) <= a and not b;
    layer0_outputs(3134) <= not a;
    layer0_outputs(3135) <= a or b;
    layer0_outputs(3136) <= b and not a;
    layer0_outputs(3137) <= a xor b;
    layer0_outputs(3138) <= not a or b;
    layer0_outputs(3139) <= not b;
    layer0_outputs(3140) <= not (a or b);
    layer0_outputs(3141) <= not (a xor b);
    layer0_outputs(3142) <= a and b;
    layer0_outputs(3143) <= not b;
    layer0_outputs(3144) <= not a;
    layer0_outputs(3145) <= b and not a;
    layer0_outputs(3146) <= b and not a;
    layer0_outputs(3147) <= a and b;
    layer0_outputs(3148) <= b and not a;
    layer0_outputs(3149) <= not (a or b);
    layer0_outputs(3150) <= a or b;
    layer0_outputs(3151) <= not b;
    layer0_outputs(3152) <= a or b;
    layer0_outputs(3153) <= not (a or b);
    layer0_outputs(3154) <= not b;
    layer0_outputs(3155) <= a and b;
    layer0_outputs(3156) <= a;
    layer0_outputs(3157) <= a and not b;
    layer0_outputs(3158) <= b;
    layer0_outputs(3159) <= '0';
    layer0_outputs(3160) <= not b;
    layer0_outputs(3161) <= a;
    layer0_outputs(3162) <= not b or a;
    layer0_outputs(3163) <= not (a or b);
    layer0_outputs(3164) <= a;
    layer0_outputs(3165) <= not a or b;
    layer0_outputs(3166) <= not (a and b);
    layer0_outputs(3167) <= b;
    layer0_outputs(3168) <= a and not b;
    layer0_outputs(3169) <= a;
    layer0_outputs(3170) <= not a;
    layer0_outputs(3171) <= not b or a;
    layer0_outputs(3172) <= a or b;
    layer0_outputs(3173) <= b;
    layer0_outputs(3174) <= not a or b;
    layer0_outputs(3175) <= a xor b;
    layer0_outputs(3176) <= not a or b;
    layer0_outputs(3177) <= not (a or b);
    layer0_outputs(3178) <= not (a or b);
    layer0_outputs(3179) <= not a;
    layer0_outputs(3180) <= a or b;
    layer0_outputs(3181) <= not (a or b);
    layer0_outputs(3182) <= a xor b;
    layer0_outputs(3183) <= not a or b;
    layer0_outputs(3184) <= not b;
    layer0_outputs(3185) <= not b or a;
    layer0_outputs(3186) <= a xor b;
    layer0_outputs(3187) <= not (a xor b);
    layer0_outputs(3188) <= not b;
    layer0_outputs(3189) <= not (a xor b);
    layer0_outputs(3190) <= not (a or b);
    layer0_outputs(3191) <= not b;
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= not (a or b);
    layer0_outputs(3194) <= not a or b;
    layer0_outputs(3195) <= not a;
    layer0_outputs(3196) <= b;
    layer0_outputs(3197) <= a;
    layer0_outputs(3198) <= '0';
    layer0_outputs(3199) <= a and b;
    layer0_outputs(3200) <= not (a or b);
    layer0_outputs(3201) <= '1';
    layer0_outputs(3202) <= a or b;
    layer0_outputs(3203) <= not b;
    layer0_outputs(3204) <= a or b;
    layer0_outputs(3205) <= not b or a;
    layer0_outputs(3206) <= b and not a;
    layer0_outputs(3207) <= not b;
    layer0_outputs(3208) <= not a;
    layer0_outputs(3209) <= b and not a;
    layer0_outputs(3210) <= not b;
    layer0_outputs(3211) <= a and not b;
    layer0_outputs(3212) <= a or b;
    layer0_outputs(3213) <= not (a or b);
    layer0_outputs(3214) <= not a or b;
    layer0_outputs(3215) <= a and not b;
    layer0_outputs(3216) <= not (a or b);
    layer0_outputs(3217) <= a xor b;
    layer0_outputs(3218) <= not b or a;
    layer0_outputs(3219) <= b;
    layer0_outputs(3220) <= a or b;
    layer0_outputs(3221) <= a or b;
    layer0_outputs(3222) <= a;
    layer0_outputs(3223) <= not (a xor b);
    layer0_outputs(3224) <= a xor b;
    layer0_outputs(3225) <= not b or a;
    layer0_outputs(3226) <= not b or a;
    layer0_outputs(3227) <= not (a or b);
    layer0_outputs(3228) <= a;
    layer0_outputs(3229) <= a;
    layer0_outputs(3230) <= b;
    layer0_outputs(3231) <= a xor b;
    layer0_outputs(3232) <= not (a and b);
    layer0_outputs(3233) <= a or b;
    layer0_outputs(3234) <= not b;
    layer0_outputs(3235) <= not b or a;
    layer0_outputs(3236) <= a;
    layer0_outputs(3237) <= a xor b;
    layer0_outputs(3238) <= not (a xor b);
    layer0_outputs(3239) <= a and b;
    layer0_outputs(3240) <= not a;
    layer0_outputs(3241) <= not (a xor b);
    layer0_outputs(3242) <= a or b;
    layer0_outputs(3243) <= a or b;
    layer0_outputs(3244) <= not (a xor b);
    layer0_outputs(3245) <= not (a xor b);
    layer0_outputs(3246) <= not a;
    layer0_outputs(3247) <= not a or b;
    layer0_outputs(3248) <= not a or b;
    layer0_outputs(3249) <= not b;
    layer0_outputs(3250) <= a and not b;
    layer0_outputs(3251) <= a;
    layer0_outputs(3252) <= not b or a;
    layer0_outputs(3253) <= not b or a;
    layer0_outputs(3254) <= not (a or b);
    layer0_outputs(3255) <= a and not b;
    layer0_outputs(3256) <= a or b;
    layer0_outputs(3257) <= not (a xor b);
    layer0_outputs(3258) <= a;
    layer0_outputs(3259) <= not b or a;
    layer0_outputs(3260) <= a and b;
    layer0_outputs(3261) <= not a or b;
    layer0_outputs(3262) <= a and b;
    layer0_outputs(3263) <= not (a or b);
    layer0_outputs(3264) <= a;
    layer0_outputs(3265) <= a or b;
    layer0_outputs(3266) <= a or b;
    layer0_outputs(3267) <= '1';
    layer0_outputs(3268) <= a or b;
    layer0_outputs(3269) <= '1';
    layer0_outputs(3270) <= a or b;
    layer0_outputs(3271) <= not a;
    layer0_outputs(3272) <= a;
    layer0_outputs(3273) <= not (a or b);
    layer0_outputs(3274) <= not b;
    layer0_outputs(3275) <= a and not b;
    layer0_outputs(3276) <= not (a xor b);
    layer0_outputs(3277) <= a and not b;
    layer0_outputs(3278) <= not (a or b);
    layer0_outputs(3279) <= '0';
    layer0_outputs(3280) <= not (a or b);
    layer0_outputs(3281) <= '0';
    layer0_outputs(3282) <= not a or b;
    layer0_outputs(3283) <= a or b;
    layer0_outputs(3284) <= not (a xor b);
    layer0_outputs(3285) <= a or b;
    layer0_outputs(3286) <= not (a or b);
    layer0_outputs(3287) <= not a;
    layer0_outputs(3288) <= not a or b;
    layer0_outputs(3289) <= a and not b;
    layer0_outputs(3290) <= b;
    layer0_outputs(3291) <= b;
    layer0_outputs(3292) <= not (a xor b);
    layer0_outputs(3293) <= '0';
    layer0_outputs(3294) <= a and not b;
    layer0_outputs(3295) <= not a or b;
    layer0_outputs(3296) <= b and not a;
    layer0_outputs(3297) <= '1';
    layer0_outputs(3298) <= not a;
    layer0_outputs(3299) <= b and not a;
    layer0_outputs(3300) <= not (a xor b);
    layer0_outputs(3301) <= b and not a;
    layer0_outputs(3302) <= a xor b;
    layer0_outputs(3303) <= not b or a;
    layer0_outputs(3304) <= b;
    layer0_outputs(3305) <= not (a or b);
    layer0_outputs(3306) <= not a;
    layer0_outputs(3307) <= b;
    layer0_outputs(3308) <= not (a or b);
    layer0_outputs(3309) <= '1';
    layer0_outputs(3310) <= not a or b;
    layer0_outputs(3311) <= not b or a;
    layer0_outputs(3312) <= a xor b;
    layer0_outputs(3313) <= a and not b;
    layer0_outputs(3314) <= '0';
    layer0_outputs(3315) <= a;
    layer0_outputs(3316) <= not a;
    layer0_outputs(3317) <= not a;
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= a and not b;
    layer0_outputs(3320) <= not a or b;
    layer0_outputs(3321) <= not a;
    layer0_outputs(3322) <= a xor b;
    layer0_outputs(3323) <= not (a or b);
    layer0_outputs(3324) <= not b;
    layer0_outputs(3325) <= a or b;
    layer0_outputs(3326) <= not a;
    layer0_outputs(3327) <= not (a and b);
    layer0_outputs(3328) <= not b or a;
    layer0_outputs(3329) <= not a;
    layer0_outputs(3330) <= not a or b;
    layer0_outputs(3331) <= not b or a;
    layer0_outputs(3332) <= not (a or b);
    layer0_outputs(3333) <= b and not a;
    layer0_outputs(3334) <= not b;
    layer0_outputs(3335) <= a;
    layer0_outputs(3336) <= a or b;
    layer0_outputs(3337) <= a and b;
    layer0_outputs(3338) <= a and not b;
    layer0_outputs(3339) <= not b or a;
    layer0_outputs(3340) <= not a;
    layer0_outputs(3341) <= '1';
    layer0_outputs(3342) <= not (a xor b);
    layer0_outputs(3343) <= not b or a;
    layer0_outputs(3344) <= b;
    layer0_outputs(3345) <= not a or b;
    layer0_outputs(3346) <= a or b;
    layer0_outputs(3347) <= a and not b;
    layer0_outputs(3348) <= a and b;
    layer0_outputs(3349) <= a xor b;
    layer0_outputs(3350) <= not (a xor b);
    layer0_outputs(3351) <= not b;
    layer0_outputs(3352) <= not b;
    layer0_outputs(3353) <= not (a xor b);
    layer0_outputs(3354) <= not a;
    layer0_outputs(3355) <= not (a or b);
    layer0_outputs(3356) <= a or b;
    layer0_outputs(3357) <= a;
    layer0_outputs(3358) <= a;
    layer0_outputs(3359) <= not a;
    layer0_outputs(3360) <= '1';
    layer0_outputs(3361) <= not b;
    layer0_outputs(3362) <= a xor b;
    layer0_outputs(3363) <= b;
    layer0_outputs(3364) <= not (a or b);
    layer0_outputs(3365) <= not b or a;
    layer0_outputs(3366) <= a xor b;
    layer0_outputs(3367) <= '1';
    layer0_outputs(3368) <= not b or a;
    layer0_outputs(3369) <= not a or b;
    layer0_outputs(3370) <= a;
    layer0_outputs(3371) <= '1';
    layer0_outputs(3372) <= not (a and b);
    layer0_outputs(3373) <= a or b;
    layer0_outputs(3374) <= b;
    layer0_outputs(3375) <= not (a or b);
    layer0_outputs(3376) <= not (a or b);
    layer0_outputs(3377) <= b and not a;
    layer0_outputs(3378) <= '0';
    layer0_outputs(3379) <= not (a or b);
    layer0_outputs(3380) <= a;
    layer0_outputs(3381) <= a;
    layer0_outputs(3382) <= a xor b;
    layer0_outputs(3383) <= b;
    layer0_outputs(3384) <= b;
    layer0_outputs(3385) <= a xor b;
    layer0_outputs(3386) <= b;
    layer0_outputs(3387) <= b;
    layer0_outputs(3388) <= not (a or b);
    layer0_outputs(3389) <= not b or a;
    layer0_outputs(3390) <= a or b;
    layer0_outputs(3391) <= not (a or b);
    layer0_outputs(3392) <= not a or b;
    layer0_outputs(3393) <= b;
    layer0_outputs(3394) <= b and not a;
    layer0_outputs(3395) <= not a or b;
    layer0_outputs(3396) <= not (a and b);
    layer0_outputs(3397) <= b and not a;
    layer0_outputs(3398) <= '1';
    layer0_outputs(3399) <= not a or b;
    layer0_outputs(3400) <= a;
    layer0_outputs(3401) <= not (a xor b);
    layer0_outputs(3402) <= a or b;
    layer0_outputs(3403) <= a;
    layer0_outputs(3404) <= a or b;
    layer0_outputs(3405) <= not b;
    layer0_outputs(3406) <= not (a and b);
    layer0_outputs(3407) <= not a;
    layer0_outputs(3408) <= b;
    layer0_outputs(3409) <= not b;
    layer0_outputs(3410) <= not b or a;
    layer0_outputs(3411) <= a or b;
    layer0_outputs(3412) <= not (a xor b);
    layer0_outputs(3413) <= a xor b;
    layer0_outputs(3414) <= a or b;
    layer0_outputs(3415) <= '0';
    layer0_outputs(3416) <= not (a xor b);
    layer0_outputs(3417) <= not a;
    layer0_outputs(3418) <= not (a or b);
    layer0_outputs(3419) <= a or b;
    layer0_outputs(3420) <= not a;
    layer0_outputs(3421) <= '1';
    layer0_outputs(3422) <= not (a or b);
    layer0_outputs(3423) <= not a;
    layer0_outputs(3424) <= a;
    layer0_outputs(3425) <= a;
    layer0_outputs(3426) <= b and not a;
    layer0_outputs(3427) <= not (a or b);
    layer0_outputs(3428) <= a xor b;
    layer0_outputs(3429) <= b and not a;
    layer0_outputs(3430) <= a or b;
    layer0_outputs(3431) <= b;
    layer0_outputs(3432) <= not b;
    layer0_outputs(3433) <= a;
    layer0_outputs(3434) <= '1';
    layer0_outputs(3435) <= not (a or b);
    layer0_outputs(3436) <= not a or b;
    layer0_outputs(3437) <= not a;
    layer0_outputs(3438) <= b and not a;
    layer0_outputs(3439) <= not (a or b);
    layer0_outputs(3440) <= not (a and b);
    layer0_outputs(3441) <= b;
    layer0_outputs(3442) <= not b or a;
    layer0_outputs(3443) <= not (a xor b);
    layer0_outputs(3444) <= a or b;
    layer0_outputs(3445) <= a;
    layer0_outputs(3446) <= b and not a;
    layer0_outputs(3447) <= not (a and b);
    layer0_outputs(3448) <= not b;
    layer0_outputs(3449) <= not b or a;
    layer0_outputs(3450) <= a;
    layer0_outputs(3451) <= not a or b;
    layer0_outputs(3452) <= not a;
    layer0_outputs(3453) <= not a or b;
    layer0_outputs(3454) <= not a;
    layer0_outputs(3455) <= b;
    layer0_outputs(3456) <= not a or b;
    layer0_outputs(3457) <= a xor b;
    layer0_outputs(3458) <= a;
    layer0_outputs(3459) <= not (a or b);
    layer0_outputs(3460) <= b;
    layer0_outputs(3461) <= b and not a;
    layer0_outputs(3462) <= a and not b;
    layer0_outputs(3463) <= not b or a;
    layer0_outputs(3464) <= not a;
    layer0_outputs(3465) <= not a;
    layer0_outputs(3466) <= a or b;
    layer0_outputs(3467) <= a;
    layer0_outputs(3468) <= not b or a;
    layer0_outputs(3469) <= not a;
    layer0_outputs(3470) <= '1';
    layer0_outputs(3471) <= '0';
    layer0_outputs(3472) <= not (a or b);
    layer0_outputs(3473) <= a;
    layer0_outputs(3474) <= not (a or b);
    layer0_outputs(3475) <= a and not b;
    layer0_outputs(3476) <= not (a and b);
    layer0_outputs(3477) <= not a;
    layer0_outputs(3478) <= b;
    layer0_outputs(3479) <= '0';
    layer0_outputs(3480) <= not (a or b);
    layer0_outputs(3481) <= not a or b;
    layer0_outputs(3482) <= a xor b;
    layer0_outputs(3483) <= b and not a;
    layer0_outputs(3484) <= not (a and b);
    layer0_outputs(3485) <= not (a xor b);
    layer0_outputs(3486) <= not b;
    layer0_outputs(3487) <= not (a or b);
    layer0_outputs(3488) <= not b or a;
    layer0_outputs(3489) <= not b;
    layer0_outputs(3490) <= not b or a;
    layer0_outputs(3491) <= a xor b;
    layer0_outputs(3492) <= not b or a;
    layer0_outputs(3493) <= b;
    layer0_outputs(3494) <= a or b;
    layer0_outputs(3495) <= not b or a;
    layer0_outputs(3496) <= not a;
    layer0_outputs(3497) <= a xor b;
    layer0_outputs(3498) <= a xor b;
    layer0_outputs(3499) <= not (a or b);
    layer0_outputs(3500) <= a;
    layer0_outputs(3501) <= a and b;
    layer0_outputs(3502) <= b and not a;
    layer0_outputs(3503) <= not (a and b);
    layer0_outputs(3504) <= not a or b;
    layer0_outputs(3505) <= a or b;
    layer0_outputs(3506) <= a and b;
    layer0_outputs(3507) <= a;
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= a or b;
    layer0_outputs(3510) <= a;
    layer0_outputs(3511) <= a and b;
    layer0_outputs(3512) <= not b or a;
    layer0_outputs(3513) <= a xor b;
    layer0_outputs(3514) <= not (a or b);
    layer0_outputs(3515) <= not b or a;
    layer0_outputs(3516) <= '0';
    layer0_outputs(3517) <= b and not a;
    layer0_outputs(3518) <= not b or a;
    layer0_outputs(3519) <= a;
    layer0_outputs(3520) <= not (a xor b);
    layer0_outputs(3521) <= not b;
    layer0_outputs(3522) <= a or b;
    layer0_outputs(3523) <= '1';
    layer0_outputs(3524) <= b;
    layer0_outputs(3525) <= b and not a;
    layer0_outputs(3526) <= not b or a;
    layer0_outputs(3527) <= not b;
    layer0_outputs(3528) <= a;
    layer0_outputs(3529) <= not b or a;
    layer0_outputs(3530) <= a or b;
    layer0_outputs(3531) <= '1';
    layer0_outputs(3532) <= a;
    layer0_outputs(3533) <= b and not a;
    layer0_outputs(3534) <= not b;
    layer0_outputs(3535) <= not a;
    layer0_outputs(3536) <= not (a and b);
    layer0_outputs(3537) <= not a;
    layer0_outputs(3538) <= a or b;
    layer0_outputs(3539) <= not a;
    layer0_outputs(3540) <= a;
    layer0_outputs(3541) <= a xor b;
    layer0_outputs(3542) <= not a;
    layer0_outputs(3543) <= a;
    layer0_outputs(3544) <= not (a and b);
    layer0_outputs(3545) <= b and not a;
    layer0_outputs(3546) <= b and not a;
    layer0_outputs(3547) <= not (a xor b);
    layer0_outputs(3548) <= not b;
    layer0_outputs(3549) <= not (a and b);
    layer0_outputs(3550) <= b and not a;
    layer0_outputs(3551) <= a and not b;
    layer0_outputs(3552) <= b;
    layer0_outputs(3553) <= not (a or b);
    layer0_outputs(3554) <= not (a or b);
    layer0_outputs(3555) <= not (a or b);
    layer0_outputs(3556) <= not (a xor b);
    layer0_outputs(3557) <= not a or b;
    layer0_outputs(3558) <= not a or b;
    layer0_outputs(3559) <= not a;
    layer0_outputs(3560) <= not (a xor b);
    layer0_outputs(3561) <= not b or a;
    layer0_outputs(3562) <= '1';
    layer0_outputs(3563) <= not b;
    layer0_outputs(3564) <= not b;
    layer0_outputs(3565) <= a;
    layer0_outputs(3566) <= a or b;
    layer0_outputs(3567) <= not b or a;
    layer0_outputs(3568) <= a or b;
    layer0_outputs(3569) <= not (a and b);
    layer0_outputs(3570) <= a xor b;
    layer0_outputs(3571) <= '0';
    layer0_outputs(3572) <= '0';
    layer0_outputs(3573) <= b;
    layer0_outputs(3574) <= not (a or b);
    layer0_outputs(3575) <= not (a or b);
    layer0_outputs(3576) <= b;
    layer0_outputs(3577) <= not (a xor b);
    layer0_outputs(3578) <= a and not b;
    layer0_outputs(3579) <= not a;
    layer0_outputs(3580) <= not (a or b);
    layer0_outputs(3581) <= not b or a;
    layer0_outputs(3582) <= not a or b;
    layer0_outputs(3583) <= not (a or b);
    layer0_outputs(3584) <= b;
    layer0_outputs(3585) <= a or b;
    layer0_outputs(3586) <= b and not a;
    layer0_outputs(3587) <= b;
    layer0_outputs(3588) <= b and not a;
    layer0_outputs(3589) <= '1';
    layer0_outputs(3590) <= not a or b;
    layer0_outputs(3591) <= a;
    layer0_outputs(3592) <= not b or a;
    layer0_outputs(3593) <= b and not a;
    layer0_outputs(3594) <= a and not b;
    layer0_outputs(3595) <= a xor b;
    layer0_outputs(3596) <= not (a xor b);
    layer0_outputs(3597) <= a;
    layer0_outputs(3598) <= a xor b;
    layer0_outputs(3599) <= not (a and b);
    layer0_outputs(3600) <= not (a or b);
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= not b or a;
    layer0_outputs(3603) <= not a or b;
    layer0_outputs(3604) <= not b or a;
    layer0_outputs(3605) <= not (a xor b);
    layer0_outputs(3606) <= a or b;
    layer0_outputs(3607) <= not (a and b);
    layer0_outputs(3608) <= a and not b;
    layer0_outputs(3609) <= not (a or b);
    layer0_outputs(3610) <= not b or a;
    layer0_outputs(3611) <= b and not a;
    layer0_outputs(3612) <= a and not b;
    layer0_outputs(3613) <= b;
    layer0_outputs(3614) <= a and not b;
    layer0_outputs(3615) <= a xor b;
    layer0_outputs(3616) <= a and not b;
    layer0_outputs(3617) <= a;
    layer0_outputs(3618) <= not b;
    layer0_outputs(3619) <= a xor b;
    layer0_outputs(3620) <= a xor b;
    layer0_outputs(3621) <= b and not a;
    layer0_outputs(3622) <= a and b;
    layer0_outputs(3623) <= not a or b;
    layer0_outputs(3624) <= '1';
    layer0_outputs(3625) <= not b;
    layer0_outputs(3626) <= not a;
    layer0_outputs(3627) <= not a;
    layer0_outputs(3628) <= '0';
    layer0_outputs(3629) <= b and not a;
    layer0_outputs(3630) <= not (a xor b);
    layer0_outputs(3631) <= not b or a;
    layer0_outputs(3632) <= a;
    layer0_outputs(3633) <= not b;
    layer0_outputs(3634) <= not b;
    layer0_outputs(3635) <= '0';
    layer0_outputs(3636) <= not b;
    layer0_outputs(3637) <= not b;
    layer0_outputs(3638) <= a and not b;
    layer0_outputs(3639) <= a or b;
    layer0_outputs(3640) <= a and not b;
    layer0_outputs(3641) <= a and b;
    layer0_outputs(3642) <= '1';
    layer0_outputs(3643) <= b;
    layer0_outputs(3644) <= a xor b;
    layer0_outputs(3645) <= a and b;
    layer0_outputs(3646) <= not a;
    layer0_outputs(3647) <= a xor b;
    layer0_outputs(3648) <= not (a or b);
    layer0_outputs(3649) <= b and not a;
    layer0_outputs(3650) <= '0';
    layer0_outputs(3651) <= a and not b;
    layer0_outputs(3652) <= not a;
    layer0_outputs(3653) <= not (a and b);
    layer0_outputs(3654) <= b;
    layer0_outputs(3655) <= not (a xor b);
    layer0_outputs(3656) <= not (a or b);
    layer0_outputs(3657) <= not (a or b);
    layer0_outputs(3658) <= a xor b;
    layer0_outputs(3659) <= not (a xor b);
    layer0_outputs(3660) <= '1';
    layer0_outputs(3661) <= not (a or b);
    layer0_outputs(3662) <= a and not b;
    layer0_outputs(3663) <= not (a xor b);
    layer0_outputs(3664) <= '0';
    layer0_outputs(3665) <= a xor b;
    layer0_outputs(3666) <= a xor b;
    layer0_outputs(3667) <= not a;
    layer0_outputs(3668) <= not b;
    layer0_outputs(3669) <= not a;
    layer0_outputs(3670) <= not (a xor b);
    layer0_outputs(3671) <= not (a or b);
    layer0_outputs(3672) <= not (a and b);
    layer0_outputs(3673) <= '1';
    layer0_outputs(3674) <= b;
    layer0_outputs(3675) <= not a or b;
    layer0_outputs(3676) <= '0';
    layer0_outputs(3677) <= not (a and b);
    layer0_outputs(3678) <= not b;
    layer0_outputs(3679) <= a;
    layer0_outputs(3680) <= not (a or b);
    layer0_outputs(3681) <= not (a or b);
    layer0_outputs(3682) <= a or b;
    layer0_outputs(3683) <= '1';
    layer0_outputs(3684) <= a xor b;
    layer0_outputs(3685) <= a xor b;
    layer0_outputs(3686) <= a and b;
    layer0_outputs(3687) <= a;
    layer0_outputs(3688) <= not a or b;
    layer0_outputs(3689) <= a xor b;
    layer0_outputs(3690) <= not (a or b);
    layer0_outputs(3691) <= '0';
    layer0_outputs(3692) <= b;
    layer0_outputs(3693) <= '0';
    layer0_outputs(3694) <= a and not b;
    layer0_outputs(3695) <= not b or a;
    layer0_outputs(3696) <= not (a and b);
    layer0_outputs(3697) <= a;
    layer0_outputs(3698) <= not b;
    layer0_outputs(3699) <= not b;
    layer0_outputs(3700) <= not b or a;
    layer0_outputs(3701) <= b;
    layer0_outputs(3702) <= a;
    layer0_outputs(3703) <= a or b;
    layer0_outputs(3704) <= b;
    layer0_outputs(3705) <= a;
    layer0_outputs(3706) <= b and not a;
    layer0_outputs(3707) <= b and not a;
    layer0_outputs(3708) <= not a;
    layer0_outputs(3709) <= not (a or b);
    layer0_outputs(3710) <= a;
    layer0_outputs(3711) <= b;
    layer0_outputs(3712) <= not a or b;
    layer0_outputs(3713) <= a or b;
    layer0_outputs(3714) <= not a or b;
    layer0_outputs(3715) <= a xor b;
    layer0_outputs(3716) <= a and b;
    layer0_outputs(3717) <= not b or a;
    layer0_outputs(3718) <= b and not a;
    layer0_outputs(3719) <= not b or a;
    layer0_outputs(3720) <= a;
    layer0_outputs(3721) <= not b;
    layer0_outputs(3722) <= a or b;
    layer0_outputs(3723) <= a or b;
    layer0_outputs(3724) <= a;
    layer0_outputs(3725) <= a or b;
    layer0_outputs(3726) <= not a;
    layer0_outputs(3727) <= a or b;
    layer0_outputs(3728) <= b and not a;
    layer0_outputs(3729) <= b and not a;
    layer0_outputs(3730) <= not b or a;
    layer0_outputs(3731) <= '0';
    layer0_outputs(3732) <= a or b;
    layer0_outputs(3733) <= not b or a;
    layer0_outputs(3734) <= not a;
    layer0_outputs(3735) <= a and b;
    layer0_outputs(3736) <= not b;
    layer0_outputs(3737) <= a and not b;
    layer0_outputs(3738) <= not b;
    layer0_outputs(3739) <= not a or b;
    layer0_outputs(3740) <= b and not a;
    layer0_outputs(3741) <= b;
    layer0_outputs(3742) <= a xor b;
    layer0_outputs(3743) <= not (a xor b);
    layer0_outputs(3744) <= not b;
    layer0_outputs(3745) <= a or b;
    layer0_outputs(3746) <= a and not b;
    layer0_outputs(3747) <= not (a or b);
    layer0_outputs(3748) <= not (a and b);
    layer0_outputs(3749) <= a and not b;
    layer0_outputs(3750) <= a;
    layer0_outputs(3751) <= b and not a;
    layer0_outputs(3752) <= not (a xor b);
    layer0_outputs(3753) <= a or b;
    layer0_outputs(3754) <= a and not b;
    layer0_outputs(3755) <= not (a or b);
    layer0_outputs(3756) <= a or b;
    layer0_outputs(3757) <= not b;
    layer0_outputs(3758) <= not (a or b);
    layer0_outputs(3759) <= a xor b;
    layer0_outputs(3760) <= '1';
    layer0_outputs(3761) <= b;
    layer0_outputs(3762) <= a and not b;
    layer0_outputs(3763) <= not b;
    layer0_outputs(3764) <= not (a xor b);
    layer0_outputs(3765) <= b and not a;
    layer0_outputs(3766) <= b;
    layer0_outputs(3767) <= not a or b;
    layer0_outputs(3768) <= not b;
    layer0_outputs(3769) <= b and not a;
    layer0_outputs(3770) <= b and not a;
    layer0_outputs(3771) <= not b or a;
    layer0_outputs(3772) <= not (a or b);
    layer0_outputs(3773) <= not (a xor b);
    layer0_outputs(3774) <= not b or a;
    layer0_outputs(3775) <= a xor b;
    layer0_outputs(3776) <= a or b;
    layer0_outputs(3777) <= not (a xor b);
    layer0_outputs(3778) <= a or b;
    layer0_outputs(3779) <= '0';
    layer0_outputs(3780) <= a or b;
    layer0_outputs(3781) <= not b;
    layer0_outputs(3782) <= b and not a;
    layer0_outputs(3783) <= not b;
    layer0_outputs(3784) <= a or b;
    layer0_outputs(3785) <= not b;
    layer0_outputs(3786) <= not b or a;
    layer0_outputs(3787) <= a and not b;
    layer0_outputs(3788) <= a or b;
    layer0_outputs(3789) <= a or b;
    layer0_outputs(3790) <= not b or a;
    layer0_outputs(3791) <= a and not b;
    layer0_outputs(3792) <= not (a or b);
    layer0_outputs(3793) <= not b or a;
    layer0_outputs(3794) <= not a;
    layer0_outputs(3795) <= a or b;
    layer0_outputs(3796) <= a;
    layer0_outputs(3797) <= not (a or b);
    layer0_outputs(3798) <= b and not a;
    layer0_outputs(3799) <= a or b;
    layer0_outputs(3800) <= not b or a;
    layer0_outputs(3801) <= not b or a;
    layer0_outputs(3802) <= b;
    layer0_outputs(3803) <= not (a xor b);
    layer0_outputs(3804) <= b and not a;
    layer0_outputs(3805) <= '1';
    layer0_outputs(3806) <= b;
    layer0_outputs(3807) <= a and b;
    layer0_outputs(3808) <= not a;
    layer0_outputs(3809) <= not (a xor b);
    layer0_outputs(3810) <= a or b;
    layer0_outputs(3811) <= not b;
    layer0_outputs(3812) <= not a or b;
    layer0_outputs(3813) <= a or b;
    layer0_outputs(3814) <= '1';
    layer0_outputs(3815) <= a or b;
    layer0_outputs(3816) <= a;
    layer0_outputs(3817) <= b and not a;
    layer0_outputs(3818) <= not a or b;
    layer0_outputs(3819) <= not (a or b);
    layer0_outputs(3820) <= a;
    layer0_outputs(3821) <= not (a or b);
    layer0_outputs(3822) <= a xor b;
    layer0_outputs(3823) <= not b or a;
    layer0_outputs(3824) <= not a or b;
    layer0_outputs(3825) <= a;
    layer0_outputs(3826) <= a or b;
    layer0_outputs(3827) <= a and b;
    layer0_outputs(3828) <= a or b;
    layer0_outputs(3829) <= not b or a;
    layer0_outputs(3830) <= a;
    layer0_outputs(3831) <= not a or b;
    layer0_outputs(3832) <= a;
    layer0_outputs(3833) <= a xor b;
    layer0_outputs(3834) <= not a;
    layer0_outputs(3835) <= not (a and b);
    layer0_outputs(3836) <= a or b;
    layer0_outputs(3837) <= a;
    layer0_outputs(3838) <= not b or a;
    layer0_outputs(3839) <= a or b;
    layer0_outputs(3840) <= '0';
    layer0_outputs(3841) <= not a or b;
    layer0_outputs(3842) <= a or b;
    layer0_outputs(3843) <= not (a or b);
    layer0_outputs(3844) <= not a or b;
    layer0_outputs(3845) <= a;
    layer0_outputs(3846) <= a or b;
    layer0_outputs(3847) <= a or b;
    layer0_outputs(3848) <= not (a or b);
    layer0_outputs(3849) <= a or b;
    layer0_outputs(3850) <= b;
    layer0_outputs(3851) <= not (a and b);
    layer0_outputs(3852) <= a or b;
    layer0_outputs(3853) <= '1';
    layer0_outputs(3854) <= not b;
    layer0_outputs(3855) <= a xor b;
    layer0_outputs(3856) <= b;
    layer0_outputs(3857) <= a or b;
    layer0_outputs(3858) <= not (a or b);
    layer0_outputs(3859) <= a and not b;
    layer0_outputs(3860) <= not b or a;
    layer0_outputs(3861) <= not a or b;
    layer0_outputs(3862) <= a and not b;
    layer0_outputs(3863) <= a;
    layer0_outputs(3864) <= a;
    layer0_outputs(3865) <= not a or b;
    layer0_outputs(3866) <= a;
    layer0_outputs(3867) <= a xor b;
    layer0_outputs(3868) <= not (a or b);
    layer0_outputs(3869) <= not (a or b);
    layer0_outputs(3870) <= not b;
    layer0_outputs(3871) <= not b or a;
    layer0_outputs(3872) <= a and b;
    layer0_outputs(3873) <= not a or b;
    layer0_outputs(3874) <= a or b;
    layer0_outputs(3875) <= not b or a;
    layer0_outputs(3876) <= not a;
    layer0_outputs(3877) <= a;
    layer0_outputs(3878) <= not (a xor b);
    layer0_outputs(3879) <= a or b;
    layer0_outputs(3880) <= '0';
    layer0_outputs(3881) <= not b;
    layer0_outputs(3882) <= not b or a;
    layer0_outputs(3883) <= b;
    layer0_outputs(3884) <= b;
    layer0_outputs(3885) <= not b;
    layer0_outputs(3886) <= a xor b;
    layer0_outputs(3887) <= a and not b;
    layer0_outputs(3888) <= a or b;
    layer0_outputs(3889) <= '1';
    layer0_outputs(3890) <= not (a xor b);
    layer0_outputs(3891) <= not b;
    layer0_outputs(3892) <= not a or b;
    layer0_outputs(3893) <= a and b;
    layer0_outputs(3894) <= a xor b;
    layer0_outputs(3895) <= not b or a;
    layer0_outputs(3896) <= a and not b;
    layer0_outputs(3897) <= not (a and b);
    layer0_outputs(3898) <= '1';
    layer0_outputs(3899) <= a or b;
    layer0_outputs(3900) <= not a;
    layer0_outputs(3901) <= not (a or b);
    layer0_outputs(3902) <= a;
    layer0_outputs(3903) <= '0';
    layer0_outputs(3904) <= b;
    layer0_outputs(3905) <= a or b;
    layer0_outputs(3906) <= a xor b;
    layer0_outputs(3907) <= not a;
    layer0_outputs(3908) <= b and not a;
    layer0_outputs(3909) <= not b;
    layer0_outputs(3910) <= not (a and b);
    layer0_outputs(3911) <= b;
    layer0_outputs(3912) <= not (a xor b);
    layer0_outputs(3913) <= not (a or b);
    layer0_outputs(3914) <= a;
    layer0_outputs(3915) <= b;
    layer0_outputs(3916) <= not a or b;
    layer0_outputs(3917) <= a or b;
    layer0_outputs(3918) <= b and not a;
    layer0_outputs(3919) <= b;
    layer0_outputs(3920) <= not (a or b);
    layer0_outputs(3921) <= not b;
    layer0_outputs(3922) <= not (a or b);
    layer0_outputs(3923) <= not a or b;
    layer0_outputs(3924) <= a;
    layer0_outputs(3925) <= not b;
    layer0_outputs(3926) <= not (a or b);
    layer0_outputs(3927) <= not b;
    layer0_outputs(3928) <= not b;
    layer0_outputs(3929) <= a or b;
    layer0_outputs(3930) <= not b or a;
    layer0_outputs(3931) <= not a or b;
    layer0_outputs(3932) <= a or b;
    layer0_outputs(3933) <= b;
    layer0_outputs(3934) <= not b;
    layer0_outputs(3935) <= not a or b;
    layer0_outputs(3936) <= a;
    layer0_outputs(3937) <= not a or b;
    layer0_outputs(3938) <= a or b;
    layer0_outputs(3939) <= not (a or b);
    layer0_outputs(3940) <= b;
    layer0_outputs(3941) <= '0';
    layer0_outputs(3942) <= a;
    layer0_outputs(3943) <= not a;
    layer0_outputs(3944) <= a xor b;
    layer0_outputs(3945) <= not b or a;
    layer0_outputs(3946) <= a xor b;
    layer0_outputs(3947) <= a or b;
    layer0_outputs(3948) <= a;
    layer0_outputs(3949) <= b;
    layer0_outputs(3950) <= not (a xor b);
    layer0_outputs(3951) <= a or b;
    layer0_outputs(3952) <= not (a or b);
    layer0_outputs(3953) <= not a;
    layer0_outputs(3954) <= '0';
    layer0_outputs(3955) <= '0';
    layer0_outputs(3956) <= not b;
    layer0_outputs(3957) <= b;
    layer0_outputs(3958) <= a;
    layer0_outputs(3959) <= not (a or b);
    layer0_outputs(3960) <= a and not b;
    layer0_outputs(3961) <= not a or b;
    layer0_outputs(3962) <= b and not a;
    layer0_outputs(3963) <= a and b;
    layer0_outputs(3964) <= not a or b;
    layer0_outputs(3965) <= a;
    layer0_outputs(3966) <= not a;
    layer0_outputs(3967) <= not a or b;
    layer0_outputs(3968) <= not a;
    layer0_outputs(3969) <= not (a and b);
    layer0_outputs(3970) <= not (a xor b);
    layer0_outputs(3971) <= a;
    layer0_outputs(3972) <= '1';
    layer0_outputs(3973) <= '0';
    layer0_outputs(3974) <= a or b;
    layer0_outputs(3975) <= b;
    layer0_outputs(3976) <= '1';
    layer0_outputs(3977) <= a and not b;
    layer0_outputs(3978) <= b and not a;
    layer0_outputs(3979) <= not a or b;
    layer0_outputs(3980) <= not (a or b);
    layer0_outputs(3981) <= a xor b;
    layer0_outputs(3982) <= not (a or b);
    layer0_outputs(3983) <= not (a and b);
    layer0_outputs(3984) <= a or b;
    layer0_outputs(3985) <= b and not a;
    layer0_outputs(3986) <= a and not b;
    layer0_outputs(3987) <= a xor b;
    layer0_outputs(3988) <= a xor b;
    layer0_outputs(3989) <= not a or b;
    layer0_outputs(3990) <= a;
    layer0_outputs(3991) <= a or b;
    layer0_outputs(3992) <= not a;
    layer0_outputs(3993) <= b;
    layer0_outputs(3994) <= not (a or b);
    layer0_outputs(3995) <= b and not a;
    layer0_outputs(3996) <= not a or b;
    layer0_outputs(3997) <= not (a or b);
    layer0_outputs(3998) <= a or b;
    layer0_outputs(3999) <= b and not a;
    layer0_outputs(4000) <= not a or b;
    layer0_outputs(4001) <= a or b;
    layer0_outputs(4002) <= '0';
    layer0_outputs(4003) <= b and not a;
    layer0_outputs(4004) <= b;
    layer0_outputs(4005) <= not (a or b);
    layer0_outputs(4006) <= b;
    layer0_outputs(4007) <= not (a xor b);
    layer0_outputs(4008) <= b;
    layer0_outputs(4009) <= not b;
    layer0_outputs(4010) <= '1';
    layer0_outputs(4011) <= b and not a;
    layer0_outputs(4012) <= b and not a;
    layer0_outputs(4013) <= not b;
    layer0_outputs(4014) <= a and not b;
    layer0_outputs(4015) <= not (a and b);
    layer0_outputs(4016) <= a or b;
    layer0_outputs(4017) <= not b;
    layer0_outputs(4018) <= a and b;
    layer0_outputs(4019) <= not b;
    layer0_outputs(4020) <= a or b;
    layer0_outputs(4021) <= not b or a;
    layer0_outputs(4022) <= a or b;
    layer0_outputs(4023) <= not a;
    layer0_outputs(4024) <= a or b;
    layer0_outputs(4025) <= '0';
    layer0_outputs(4026) <= '0';
    layer0_outputs(4027) <= not (a or b);
    layer0_outputs(4028) <= not b or a;
    layer0_outputs(4029) <= b and not a;
    layer0_outputs(4030) <= a xor b;
    layer0_outputs(4031) <= not b or a;
    layer0_outputs(4032) <= not a or b;
    layer0_outputs(4033) <= not a;
    layer0_outputs(4034) <= not a or b;
    layer0_outputs(4035) <= a;
    layer0_outputs(4036) <= a or b;
    layer0_outputs(4037) <= b;
    layer0_outputs(4038) <= not (a and b);
    layer0_outputs(4039) <= not b;
    layer0_outputs(4040) <= not (a or b);
    layer0_outputs(4041) <= not a or b;
    layer0_outputs(4042) <= '0';
    layer0_outputs(4043) <= a xor b;
    layer0_outputs(4044) <= not (a xor b);
    layer0_outputs(4045) <= b;
    layer0_outputs(4046) <= not (a and b);
    layer0_outputs(4047) <= b;
    layer0_outputs(4048) <= a xor b;
    layer0_outputs(4049) <= a and b;
    layer0_outputs(4050) <= not (a xor b);
    layer0_outputs(4051) <= '1';
    layer0_outputs(4052) <= not b;
    layer0_outputs(4053) <= b;
    layer0_outputs(4054) <= not b or a;
    layer0_outputs(4055) <= b;
    layer0_outputs(4056) <= b and not a;
    layer0_outputs(4057) <= not (a or b);
    layer0_outputs(4058) <= a;
    layer0_outputs(4059) <= not b or a;
    layer0_outputs(4060) <= a;
    layer0_outputs(4061) <= not a;
    layer0_outputs(4062) <= not a;
    layer0_outputs(4063) <= a;
    layer0_outputs(4064) <= '0';
    layer0_outputs(4065) <= b and not a;
    layer0_outputs(4066) <= b and not a;
    layer0_outputs(4067) <= not (a or b);
    layer0_outputs(4068) <= not (a and b);
    layer0_outputs(4069) <= a;
    layer0_outputs(4070) <= b and not a;
    layer0_outputs(4071) <= a and b;
    layer0_outputs(4072) <= not b or a;
    layer0_outputs(4073) <= a xor b;
    layer0_outputs(4074) <= not (a xor b);
    layer0_outputs(4075) <= a;
    layer0_outputs(4076) <= not (a or b);
    layer0_outputs(4077) <= '0';
    layer0_outputs(4078) <= not (a or b);
    layer0_outputs(4079) <= not a or b;
    layer0_outputs(4080) <= not (a and b);
    layer0_outputs(4081) <= not (a or b);
    layer0_outputs(4082) <= a and not b;
    layer0_outputs(4083) <= not b or a;
    layer0_outputs(4084) <= a xor b;
    layer0_outputs(4085) <= a xor b;
    layer0_outputs(4086) <= a and b;
    layer0_outputs(4087) <= a;
    layer0_outputs(4088) <= a and b;
    layer0_outputs(4089) <= not (a or b);
    layer0_outputs(4090) <= not a;
    layer0_outputs(4091) <= '0';
    layer0_outputs(4092) <= a and b;
    layer0_outputs(4093) <= not a;
    layer0_outputs(4094) <= a and b;
    layer0_outputs(4095) <= b;
    layer0_outputs(4096) <= a or b;
    layer0_outputs(4097) <= not b;
    layer0_outputs(4098) <= a or b;
    layer0_outputs(4099) <= a xor b;
    layer0_outputs(4100) <= not a or b;
    layer0_outputs(4101) <= not (a xor b);
    layer0_outputs(4102) <= a xor b;
    layer0_outputs(4103) <= b and not a;
    layer0_outputs(4104) <= not (a or b);
    layer0_outputs(4105) <= b;
    layer0_outputs(4106) <= b;
    layer0_outputs(4107) <= not b;
    layer0_outputs(4108) <= a xor b;
    layer0_outputs(4109) <= a or b;
    layer0_outputs(4110) <= not a;
    layer0_outputs(4111) <= not (a xor b);
    layer0_outputs(4112) <= not a or b;
    layer0_outputs(4113) <= not b or a;
    layer0_outputs(4114) <= not (a xor b);
    layer0_outputs(4115) <= a and not b;
    layer0_outputs(4116) <= not a;
    layer0_outputs(4117) <= a and not b;
    layer0_outputs(4118) <= a;
    layer0_outputs(4119) <= not (a xor b);
    layer0_outputs(4120) <= a xor b;
    layer0_outputs(4121) <= a or b;
    layer0_outputs(4122) <= not b;
    layer0_outputs(4123) <= b;
    layer0_outputs(4124) <= b;
    layer0_outputs(4125) <= not a;
    layer0_outputs(4126) <= not a;
    layer0_outputs(4127) <= not (a xor b);
    layer0_outputs(4128) <= not a or b;
    layer0_outputs(4129) <= a;
    layer0_outputs(4130) <= a or b;
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= a and b;
    layer0_outputs(4133) <= not b;
    layer0_outputs(4134) <= '0';
    layer0_outputs(4135) <= a or b;
    layer0_outputs(4136) <= not (a or b);
    layer0_outputs(4137) <= a and b;
    layer0_outputs(4138) <= not b;
    layer0_outputs(4139) <= not a or b;
    layer0_outputs(4140) <= not a or b;
    layer0_outputs(4141) <= a xor b;
    layer0_outputs(4142) <= '1';
    layer0_outputs(4143) <= '0';
    layer0_outputs(4144) <= b and not a;
    layer0_outputs(4145) <= a and not b;
    layer0_outputs(4146) <= not b;
    layer0_outputs(4147) <= not (a and b);
    layer0_outputs(4148) <= '1';
    layer0_outputs(4149) <= not b;
    layer0_outputs(4150) <= not (a xor b);
    layer0_outputs(4151) <= a and b;
    layer0_outputs(4152) <= not b or a;
    layer0_outputs(4153) <= not a;
    layer0_outputs(4154) <= not a or b;
    layer0_outputs(4155) <= a or b;
    layer0_outputs(4156) <= '0';
    layer0_outputs(4157) <= not (a or b);
    layer0_outputs(4158) <= not a;
    layer0_outputs(4159) <= not a or b;
    layer0_outputs(4160) <= b and not a;
    layer0_outputs(4161) <= not (a or b);
    layer0_outputs(4162) <= a xor b;
    layer0_outputs(4163) <= not a;
    layer0_outputs(4164) <= not b or a;
    layer0_outputs(4165) <= not (a xor b);
    layer0_outputs(4166) <= b;
    layer0_outputs(4167) <= not (a or b);
    layer0_outputs(4168) <= not (a xor b);
    layer0_outputs(4169) <= not a or b;
    layer0_outputs(4170) <= not a or b;
    layer0_outputs(4171) <= a or b;
    layer0_outputs(4172) <= b;
    layer0_outputs(4173) <= not (a xor b);
    layer0_outputs(4174) <= not (a or b);
    layer0_outputs(4175) <= not (a or b);
    layer0_outputs(4176) <= not a or b;
    layer0_outputs(4177) <= a and b;
    layer0_outputs(4178) <= a and not b;
    layer0_outputs(4179) <= not (a or b);
    layer0_outputs(4180) <= b;
    layer0_outputs(4181) <= not a or b;
    layer0_outputs(4182) <= b;
    layer0_outputs(4183) <= not (a and b);
    layer0_outputs(4184) <= not b or a;
    layer0_outputs(4185) <= '1';
    layer0_outputs(4186) <= a and b;
    layer0_outputs(4187) <= a;
    layer0_outputs(4188) <= a or b;
    layer0_outputs(4189) <= a and b;
    layer0_outputs(4190) <= a xor b;
    layer0_outputs(4191) <= not (a or b);
    layer0_outputs(4192) <= not a;
    layer0_outputs(4193) <= not (a or b);
    layer0_outputs(4194) <= a or b;
    layer0_outputs(4195) <= a and b;
    layer0_outputs(4196) <= not (a or b);
    layer0_outputs(4197) <= b;
    layer0_outputs(4198) <= not b;
    layer0_outputs(4199) <= a or b;
    layer0_outputs(4200) <= a and not b;
    layer0_outputs(4201) <= a;
    layer0_outputs(4202) <= not (a or b);
    layer0_outputs(4203) <= a and not b;
    layer0_outputs(4204) <= a and b;
    layer0_outputs(4205) <= a and not b;
    layer0_outputs(4206) <= not a or b;
    layer0_outputs(4207) <= a;
    layer0_outputs(4208) <= a and b;
    layer0_outputs(4209) <= a or b;
    layer0_outputs(4210) <= not b or a;
    layer0_outputs(4211) <= a xor b;
    layer0_outputs(4212) <= a or b;
    layer0_outputs(4213) <= a or b;
    layer0_outputs(4214) <= a;
    layer0_outputs(4215) <= b and not a;
    layer0_outputs(4216) <= a or b;
    layer0_outputs(4217) <= not (a or b);
    layer0_outputs(4218) <= not (a xor b);
    layer0_outputs(4219) <= a and not b;
    layer0_outputs(4220) <= a or b;
    layer0_outputs(4221) <= not (a xor b);
    layer0_outputs(4222) <= not a;
    layer0_outputs(4223) <= a xor b;
    layer0_outputs(4224) <= not a or b;
    layer0_outputs(4225) <= a or b;
    layer0_outputs(4226) <= a xor b;
    layer0_outputs(4227) <= b and not a;
    layer0_outputs(4228) <= b;
    layer0_outputs(4229) <= a and not b;
    layer0_outputs(4230) <= not (a xor b);
    layer0_outputs(4231) <= b;
    layer0_outputs(4232) <= not (a or b);
    layer0_outputs(4233) <= a and not b;
    layer0_outputs(4234) <= not a or b;
    layer0_outputs(4235) <= not b or a;
    layer0_outputs(4236) <= a;
    layer0_outputs(4237) <= '0';
    layer0_outputs(4238) <= b and not a;
    layer0_outputs(4239) <= not (a or b);
    layer0_outputs(4240) <= not a or b;
    layer0_outputs(4241) <= '0';
    layer0_outputs(4242) <= a;
    layer0_outputs(4243) <= not (a or b);
    layer0_outputs(4244) <= not b or a;
    layer0_outputs(4245) <= not (a or b);
    layer0_outputs(4246) <= b;
    layer0_outputs(4247) <= b;
    layer0_outputs(4248) <= a or b;
    layer0_outputs(4249) <= b;
    layer0_outputs(4250) <= not b or a;
    layer0_outputs(4251) <= not (a and b);
    layer0_outputs(4252) <= not a;
    layer0_outputs(4253) <= not a or b;
    layer0_outputs(4254) <= not b;
    layer0_outputs(4255) <= not (a xor b);
    layer0_outputs(4256) <= not (a and b);
    layer0_outputs(4257) <= b;
    layer0_outputs(4258) <= b and not a;
    layer0_outputs(4259) <= not (a xor b);
    layer0_outputs(4260) <= not (a xor b);
    layer0_outputs(4261) <= a and not b;
    layer0_outputs(4262) <= b;
    layer0_outputs(4263) <= not (a or b);
    layer0_outputs(4264) <= not (a or b);
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= not b or a;
    layer0_outputs(4267) <= not (a and b);
    layer0_outputs(4268) <= not b;
    layer0_outputs(4269) <= not b;
    layer0_outputs(4270) <= a;
    layer0_outputs(4271) <= not b;
    layer0_outputs(4272) <= b;
    layer0_outputs(4273) <= '0';
    layer0_outputs(4274) <= not a;
    layer0_outputs(4275) <= '1';
    layer0_outputs(4276) <= a;
    layer0_outputs(4277) <= '1';
    layer0_outputs(4278) <= a or b;
    layer0_outputs(4279) <= b and not a;
    layer0_outputs(4280) <= a or b;
    layer0_outputs(4281) <= a or b;
    layer0_outputs(4282) <= not (a or b);
    layer0_outputs(4283) <= a;
    layer0_outputs(4284) <= not a;
    layer0_outputs(4285) <= a;
    layer0_outputs(4286) <= not (a and b);
    layer0_outputs(4287) <= not a or b;
    layer0_outputs(4288) <= a and not b;
    layer0_outputs(4289) <= a;
    layer0_outputs(4290) <= a xor b;
    layer0_outputs(4291) <= a or b;
    layer0_outputs(4292) <= not b;
    layer0_outputs(4293) <= a or b;
    layer0_outputs(4294) <= a;
    layer0_outputs(4295) <= a or b;
    layer0_outputs(4296) <= not a or b;
    layer0_outputs(4297) <= not (a and b);
    layer0_outputs(4298) <= a or b;
    layer0_outputs(4299) <= b;
    layer0_outputs(4300) <= not (a or b);
    layer0_outputs(4301) <= b;
    layer0_outputs(4302) <= b and not a;
    layer0_outputs(4303) <= a and not b;
    layer0_outputs(4304) <= a and not b;
    layer0_outputs(4305) <= not b or a;
    layer0_outputs(4306) <= a xor b;
    layer0_outputs(4307) <= a;
    layer0_outputs(4308) <= a xor b;
    layer0_outputs(4309) <= a or b;
    layer0_outputs(4310) <= a xor b;
    layer0_outputs(4311) <= a;
    layer0_outputs(4312) <= not a;
    layer0_outputs(4313) <= not (a xor b);
    layer0_outputs(4314) <= a xor b;
    layer0_outputs(4315) <= not (a and b);
    layer0_outputs(4316) <= b;
    layer0_outputs(4317) <= not b or a;
    layer0_outputs(4318) <= a or b;
    layer0_outputs(4319) <= a;
    layer0_outputs(4320) <= not b;
    layer0_outputs(4321) <= b;
    layer0_outputs(4322) <= not (a xor b);
    layer0_outputs(4323) <= a or b;
    layer0_outputs(4324) <= a;
    layer0_outputs(4325) <= '1';
    layer0_outputs(4326) <= not b or a;
    layer0_outputs(4327) <= not b;
    layer0_outputs(4328) <= not b;
    layer0_outputs(4329) <= b;
    layer0_outputs(4330) <= not a or b;
    layer0_outputs(4331) <= not b or a;
    layer0_outputs(4332) <= not b;
    layer0_outputs(4333) <= a or b;
    layer0_outputs(4334) <= a and not b;
    layer0_outputs(4335) <= a xor b;
    layer0_outputs(4336) <= not b or a;
    layer0_outputs(4337) <= not a or b;
    layer0_outputs(4338) <= not a;
    layer0_outputs(4339) <= not b;
    layer0_outputs(4340) <= a or b;
    layer0_outputs(4341) <= not a;
    layer0_outputs(4342) <= not (a and b);
    layer0_outputs(4343) <= not (a and b);
    layer0_outputs(4344) <= not b or a;
    layer0_outputs(4345) <= b;
    layer0_outputs(4346) <= not (a or b);
    layer0_outputs(4347) <= not b;
    layer0_outputs(4348) <= not (a or b);
    layer0_outputs(4349) <= not (a xor b);
    layer0_outputs(4350) <= not (a xor b);
    layer0_outputs(4351) <= not b or a;
    layer0_outputs(4352) <= a xor b;
    layer0_outputs(4353) <= not b;
    layer0_outputs(4354) <= a xor b;
    layer0_outputs(4355) <= a and not b;
    layer0_outputs(4356) <= a or b;
    layer0_outputs(4357) <= not (a or b);
    layer0_outputs(4358) <= '1';
    layer0_outputs(4359) <= not b;
    layer0_outputs(4360) <= a xor b;
    layer0_outputs(4361) <= not b;
    layer0_outputs(4362) <= b;
    layer0_outputs(4363) <= a and not b;
    layer0_outputs(4364) <= a or b;
    layer0_outputs(4365) <= a and not b;
    layer0_outputs(4366) <= not b;
    layer0_outputs(4367) <= a xor b;
    layer0_outputs(4368) <= not a or b;
    layer0_outputs(4369) <= b;
    layer0_outputs(4370) <= not a or b;
    layer0_outputs(4371) <= a or b;
    layer0_outputs(4372) <= not a;
    layer0_outputs(4373) <= not a or b;
    layer0_outputs(4374) <= a or b;
    layer0_outputs(4375) <= not a or b;
    layer0_outputs(4376) <= a and not b;
    layer0_outputs(4377) <= not (a xor b);
    layer0_outputs(4378) <= not (a xor b);
    layer0_outputs(4379) <= a xor b;
    layer0_outputs(4380) <= not (a xor b);
    layer0_outputs(4381) <= not a;
    layer0_outputs(4382) <= a or b;
    layer0_outputs(4383) <= not (a or b);
    layer0_outputs(4384) <= not (a or b);
    layer0_outputs(4385) <= a or b;
    layer0_outputs(4386) <= '1';
    layer0_outputs(4387) <= a or b;
    layer0_outputs(4388) <= a xor b;
    layer0_outputs(4389) <= a or b;
    layer0_outputs(4390) <= a or b;
    layer0_outputs(4391) <= not (a xor b);
    layer0_outputs(4392) <= not (a xor b);
    layer0_outputs(4393) <= a and not b;
    layer0_outputs(4394) <= not b;
    layer0_outputs(4395) <= not a or b;
    layer0_outputs(4396) <= not (a xor b);
    layer0_outputs(4397) <= a xor b;
    layer0_outputs(4398) <= not (a xor b);
    layer0_outputs(4399) <= not b;
    layer0_outputs(4400) <= not b or a;
    layer0_outputs(4401) <= not (a and b);
    layer0_outputs(4402) <= a or b;
    layer0_outputs(4403) <= not (a or b);
    layer0_outputs(4404) <= a or b;
    layer0_outputs(4405) <= b;
    layer0_outputs(4406) <= not (a xor b);
    layer0_outputs(4407) <= a;
    layer0_outputs(4408) <= not (a or b);
    layer0_outputs(4409) <= a or b;
    layer0_outputs(4410) <= a and not b;
    layer0_outputs(4411) <= not a;
    layer0_outputs(4412) <= not (a xor b);
    layer0_outputs(4413) <= not a or b;
    layer0_outputs(4414) <= not a or b;
    layer0_outputs(4415) <= not a or b;
    layer0_outputs(4416) <= not a;
    layer0_outputs(4417) <= not b or a;
    layer0_outputs(4418) <= not a or b;
    layer0_outputs(4419) <= '0';
    layer0_outputs(4420) <= not (a or b);
    layer0_outputs(4421) <= b and not a;
    layer0_outputs(4422) <= not a;
    layer0_outputs(4423) <= a xor b;
    layer0_outputs(4424) <= not b;
    layer0_outputs(4425) <= a or b;
    layer0_outputs(4426) <= a or b;
    layer0_outputs(4427) <= not (a or b);
    layer0_outputs(4428) <= a and b;
    layer0_outputs(4429) <= a or b;
    layer0_outputs(4430) <= a;
    layer0_outputs(4431) <= b and not a;
    layer0_outputs(4432) <= not (a xor b);
    layer0_outputs(4433) <= '0';
    layer0_outputs(4434) <= not a;
    layer0_outputs(4435) <= b;
    layer0_outputs(4436) <= a and b;
    layer0_outputs(4437) <= a and not b;
    layer0_outputs(4438) <= '1';
    layer0_outputs(4439) <= not b or a;
    layer0_outputs(4440) <= not a;
    layer0_outputs(4441) <= '0';
    layer0_outputs(4442) <= a or b;
    layer0_outputs(4443) <= not (a or b);
    layer0_outputs(4444) <= a xor b;
    layer0_outputs(4445) <= not (a or b);
    layer0_outputs(4446) <= a and b;
    layer0_outputs(4447) <= a or b;
    layer0_outputs(4448) <= not (a and b);
    layer0_outputs(4449) <= not (a or b);
    layer0_outputs(4450) <= '0';
    layer0_outputs(4451) <= not b or a;
    layer0_outputs(4452) <= a and not b;
    layer0_outputs(4453) <= a and not b;
    layer0_outputs(4454) <= not (a or b);
    layer0_outputs(4455) <= not (a or b);
    layer0_outputs(4456) <= a;
    layer0_outputs(4457) <= a or b;
    layer0_outputs(4458) <= a and not b;
    layer0_outputs(4459) <= b and not a;
    layer0_outputs(4460) <= not (a or b);
    layer0_outputs(4461) <= a;
    layer0_outputs(4462) <= not a;
    layer0_outputs(4463) <= not a;
    layer0_outputs(4464) <= a;
    layer0_outputs(4465) <= '0';
    layer0_outputs(4466) <= not b;
    layer0_outputs(4467) <= '0';
    layer0_outputs(4468) <= '1';
    layer0_outputs(4469) <= not (a or b);
    layer0_outputs(4470) <= b;
    layer0_outputs(4471) <= not a or b;
    layer0_outputs(4472) <= a or b;
    layer0_outputs(4473) <= a and b;
    layer0_outputs(4474) <= b and not a;
    layer0_outputs(4475) <= b;
    layer0_outputs(4476) <= a;
    layer0_outputs(4477) <= b and not a;
    layer0_outputs(4478) <= not a;
    layer0_outputs(4479) <= a xor b;
    layer0_outputs(4480) <= b;
    layer0_outputs(4481) <= not b;
    layer0_outputs(4482) <= a and not b;
    layer0_outputs(4483) <= a;
    layer0_outputs(4484) <= not a or b;
    layer0_outputs(4485) <= not b;
    layer0_outputs(4486) <= a and b;
    layer0_outputs(4487) <= not b;
    layer0_outputs(4488) <= b and not a;
    layer0_outputs(4489) <= not b;
    layer0_outputs(4490) <= a and b;
    layer0_outputs(4491) <= a and not b;
    layer0_outputs(4492) <= a xor b;
    layer0_outputs(4493) <= not (a xor b);
    layer0_outputs(4494) <= a or b;
    layer0_outputs(4495) <= not (a or b);
    layer0_outputs(4496) <= not (a xor b);
    layer0_outputs(4497) <= a and not b;
    layer0_outputs(4498) <= a and b;
    layer0_outputs(4499) <= b;
    layer0_outputs(4500) <= not (a xor b);
    layer0_outputs(4501) <= '1';
    layer0_outputs(4502) <= not a;
    layer0_outputs(4503) <= not (a xor b);
    layer0_outputs(4504) <= a and not b;
    layer0_outputs(4505) <= b;
    layer0_outputs(4506) <= not (a or b);
    layer0_outputs(4507) <= a or b;
    layer0_outputs(4508) <= a xor b;
    layer0_outputs(4509) <= a or b;
    layer0_outputs(4510) <= not (a xor b);
    layer0_outputs(4511) <= not (a or b);
    layer0_outputs(4512) <= not (a and b);
    layer0_outputs(4513) <= a or b;
    layer0_outputs(4514) <= '1';
    layer0_outputs(4515) <= a;
    layer0_outputs(4516) <= a xor b;
    layer0_outputs(4517) <= not (a xor b);
    layer0_outputs(4518) <= a xor b;
    layer0_outputs(4519) <= not (a xor b);
    layer0_outputs(4520) <= not (a or b);
    layer0_outputs(4521) <= not a;
    layer0_outputs(4522) <= a or b;
    layer0_outputs(4523) <= not (a xor b);
    layer0_outputs(4524) <= '0';
    layer0_outputs(4525) <= not b or a;
    layer0_outputs(4526) <= not (a and b);
    layer0_outputs(4527) <= not (a or b);
    layer0_outputs(4528) <= a;
    layer0_outputs(4529) <= a;
    layer0_outputs(4530) <= a;
    layer0_outputs(4531) <= a;
    layer0_outputs(4532) <= b;
    layer0_outputs(4533) <= not (a or b);
    layer0_outputs(4534) <= not (a xor b);
    layer0_outputs(4535) <= b;
    layer0_outputs(4536) <= not a or b;
    layer0_outputs(4537) <= not (a xor b);
    layer0_outputs(4538) <= b;
    layer0_outputs(4539) <= a or b;
    layer0_outputs(4540) <= a xor b;
    layer0_outputs(4541) <= not a;
    layer0_outputs(4542) <= b;
    layer0_outputs(4543) <= b;
    layer0_outputs(4544) <= not (a or b);
    layer0_outputs(4545) <= not (a xor b);
    layer0_outputs(4546) <= a xor b;
    layer0_outputs(4547) <= not (a or b);
    layer0_outputs(4548) <= not a;
    layer0_outputs(4549) <= b and not a;
    layer0_outputs(4550) <= a xor b;
    layer0_outputs(4551) <= a;
    layer0_outputs(4552) <= b and not a;
    layer0_outputs(4553) <= a and not b;
    layer0_outputs(4554) <= not a or b;
    layer0_outputs(4555) <= a and b;
    layer0_outputs(4556) <= a;
    layer0_outputs(4557) <= not (a or b);
    layer0_outputs(4558) <= not b or a;
    layer0_outputs(4559) <= a;
    layer0_outputs(4560) <= not b or a;
    layer0_outputs(4561) <= b;
    layer0_outputs(4562) <= a;
    layer0_outputs(4563) <= a or b;
    layer0_outputs(4564) <= not b or a;
    layer0_outputs(4565) <= a or b;
    layer0_outputs(4566) <= not (a or b);
    layer0_outputs(4567) <= not (a xor b);
    layer0_outputs(4568) <= a xor b;
    layer0_outputs(4569) <= a xor b;
    layer0_outputs(4570) <= not b;
    layer0_outputs(4571) <= a or b;
    layer0_outputs(4572) <= b;
    layer0_outputs(4573) <= a and not b;
    layer0_outputs(4574) <= not a or b;
    layer0_outputs(4575) <= a xor b;
    layer0_outputs(4576) <= '1';
    layer0_outputs(4577) <= not (a or b);
    layer0_outputs(4578) <= not a or b;
    layer0_outputs(4579) <= not a;
    layer0_outputs(4580) <= not a;
    layer0_outputs(4581) <= not (a or b);
    layer0_outputs(4582) <= not b;
    layer0_outputs(4583) <= b and not a;
    layer0_outputs(4584) <= a or b;
    layer0_outputs(4585) <= not (a or b);
    layer0_outputs(4586) <= not a;
    layer0_outputs(4587) <= a;
    layer0_outputs(4588) <= '0';
    layer0_outputs(4589) <= a xor b;
    layer0_outputs(4590) <= not (a and b);
    layer0_outputs(4591) <= b;
    layer0_outputs(4592) <= a or b;
    layer0_outputs(4593) <= a or b;
    layer0_outputs(4594) <= a or b;
    layer0_outputs(4595) <= not a;
    layer0_outputs(4596) <= not b;
    layer0_outputs(4597) <= not b;
    layer0_outputs(4598) <= not (a or b);
    layer0_outputs(4599) <= a;
    layer0_outputs(4600) <= b;
    layer0_outputs(4601) <= a xor b;
    layer0_outputs(4602) <= not (a or b);
    layer0_outputs(4603) <= not (a or b);
    layer0_outputs(4604) <= not a;
    layer0_outputs(4605) <= not (a or b);
    layer0_outputs(4606) <= '1';
    layer0_outputs(4607) <= a or b;
    layer0_outputs(4608) <= not b;
    layer0_outputs(4609) <= a and not b;
    layer0_outputs(4610) <= '0';
    layer0_outputs(4611) <= '1';
    layer0_outputs(4612) <= not (a xor b);
    layer0_outputs(4613) <= not (a xor b);
    layer0_outputs(4614) <= not (a and b);
    layer0_outputs(4615) <= b and not a;
    layer0_outputs(4616) <= not a or b;
    layer0_outputs(4617) <= not b or a;
    layer0_outputs(4618) <= not (a or b);
    layer0_outputs(4619) <= not (a or b);
    layer0_outputs(4620) <= not b;
    layer0_outputs(4621) <= a or b;
    layer0_outputs(4622) <= not (a or b);
    layer0_outputs(4623) <= '0';
    layer0_outputs(4624) <= not (a or b);
    layer0_outputs(4625) <= not (a xor b);
    layer0_outputs(4626) <= a;
    layer0_outputs(4627) <= not b or a;
    layer0_outputs(4628) <= a;
    layer0_outputs(4629) <= a;
    layer0_outputs(4630) <= not a or b;
    layer0_outputs(4631) <= a xor b;
    layer0_outputs(4632) <= not a or b;
    layer0_outputs(4633) <= not (a or b);
    layer0_outputs(4634) <= not (a or b);
    layer0_outputs(4635) <= not (a or b);
    layer0_outputs(4636) <= not (a or b);
    layer0_outputs(4637) <= not a or b;
    layer0_outputs(4638) <= a and not b;
    layer0_outputs(4639) <= not a;
    layer0_outputs(4640) <= not a;
    layer0_outputs(4641) <= not a;
    layer0_outputs(4642) <= not (a or b);
    layer0_outputs(4643) <= not (a and b);
    layer0_outputs(4644) <= a xor b;
    layer0_outputs(4645) <= b and not a;
    layer0_outputs(4646) <= not b;
    layer0_outputs(4647) <= b;
    layer0_outputs(4648) <= a and not b;
    layer0_outputs(4649) <= a xor b;
    layer0_outputs(4650) <= a xor b;
    layer0_outputs(4651) <= a and not b;
    layer0_outputs(4652) <= a and not b;
    layer0_outputs(4653) <= a and b;
    layer0_outputs(4654) <= not b or a;
    layer0_outputs(4655) <= not (a or b);
    layer0_outputs(4656) <= a and not b;
    layer0_outputs(4657) <= a and not b;
    layer0_outputs(4658) <= not (a or b);
    layer0_outputs(4659) <= a xor b;
    layer0_outputs(4660) <= b;
    layer0_outputs(4661) <= not (a xor b);
    layer0_outputs(4662) <= not (a xor b);
    layer0_outputs(4663) <= a;
    layer0_outputs(4664) <= a and not b;
    layer0_outputs(4665) <= a or b;
    layer0_outputs(4666) <= not (a or b);
    layer0_outputs(4667) <= not b;
    layer0_outputs(4668) <= not a or b;
    layer0_outputs(4669) <= a and not b;
    layer0_outputs(4670) <= not b;
    layer0_outputs(4671) <= b;
    layer0_outputs(4672) <= a or b;
    layer0_outputs(4673) <= b and not a;
    layer0_outputs(4674) <= '1';
    layer0_outputs(4675) <= a xor b;
    layer0_outputs(4676) <= b and not a;
    layer0_outputs(4677) <= b and not a;
    layer0_outputs(4678) <= not (a or b);
    layer0_outputs(4679) <= a and not b;
    layer0_outputs(4680) <= a xor b;
    layer0_outputs(4681) <= '1';
    layer0_outputs(4682) <= b;
    layer0_outputs(4683) <= a and not b;
    layer0_outputs(4684) <= b and not a;
    layer0_outputs(4685) <= a xor b;
    layer0_outputs(4686) <= b and not a;
    layer0_outputs(4687) <= a;
    layer0_outputs(4688) <= a;
    layer0_outputs(4689) <= a or b;
    layer0_outputs(4690) <= not (a and b);
    layer0_outputs(4691) <= a or b;
    layer0_outputs(4692) <= not b or a;
    layer0_outputs(4693) <= not (a xor b);
    layer0_outputs(4694) <= b and not a;
    layer0_outputs(4695) <= not a or b;
    layer0_outputs(4696) <= a and not b;
    layer0_outputs(4697) <= a and not b;
    layer0_outputs(4698) <= not (a or b);
    layer0_outputs(4699) <= a or b;
    layer0_outputs(4700) <= not (a xor b);
    layer0_outputs(4701) <= not (a or b);
    layer0_outputs(4702) <= not (a or b);
    layer0_outputs(4703) <= not (a or b);
    layer0_outputs(4704) <= not (a and b);
    layer0_outputs(4705) <= '0';
    layer0_outputs(4706) <= a;
    layer0_outputs(4707) <= a;
    layer0_outputs(4708) <= not (a or b);
    layer0_outputs(4709) <= a or b;
    layer0_outputs(4710) <= '0';
    layer0_outputs(4711) <= not b or a;
    layer0_outputs(4712) <= '1';
    layer0_outputs(4713) <= not (a xor b);
    layer0_outputs(4714) <= '0';
    layer0_outputs(4715) <= a or b;
    layer0_outputs(4716) <= not a or b;
    layer0_outputs(4717) <= not (a or b);
    layer0_outputs(4718) <= a and not b;
    layer0_outputs(4719) <= not b;
    layer0_outputs(4720) <= not b;
    layer0_outputs(4721) <= not (a or b);
    layer0_outputs(4722) <= '1';
    layer0_outputs(4723) <= not b;
    layer0_outputs(4724) <= a or b;
    layer0_outputs(4725) <= a or b;
    layer0_outputs(4726) <= not b;
    layer0_outputs(4727) <= b and not a;
    layer0_outputs(4728) <= '1';
    layer0_outputs(4729) <= not a or b;
    layer0_outputs(4730) <= '1';
    layer0_outputs(4731) <= not (a or b);
    layer0_outputs(4732) <= b and not a;
    layer0_outputs(4733) <= '0';
    layer0_outputs(4734) <= not b or a;
    layer0_outputs(4735) <= a and not b;
    layer0_outputs(4736) <= not b;
    layer0_outputs(4737) <= not (a or b);
    layer0_outputs(4738) <= not (a xor b);
    layer0_outputs(4739) <= a and not b;
    layer0_outputs(4740) <= a xor b;
    layer0_outputs(4741) <= a and not b;
    layer0_outputs(4742) <= b;
    layer0_outputs(4743) <= not a or b;
    layer0_outputs(4744) <= a or b;
    layer0_outputs(4745) <= a and not b;
    layer0_outputs(4746) <= not (a xor b);
    layer0_outputs(4747) <= b and not a;
    layer0_outputs(4748) <= '0';
    layer0_outputs(4749) <= not a;
    layer0_outputs(4750) <= a and not b;
    layer0_outputs(4751) <= not b;
    layer0_outputs(4752) <= not b or a;
    layer0_outputs(4753) <= a and not b;
    layer0_outputs(4754) <= '0';
    layer0_outputs(4755) <= not a;
    layer0_outputs(4756) <= not a;
    layer0_outputs(4757) <= a;
    layer0_outputs(4758) <= a or b;
    layer0_outputs(4759) <= a or b;
    layer0_outputs(4760) <= '0';
    layer0_outputs(4761) <= a xor b;
    layer0_outputs(4762) <= not (a or b);
    layer0_outputs(4763) <= a;
    layer0_outputs(4764) <= a and not b;
    layer0_outputs(4765) <= not b;
    layer0_outputs(4766) <= a xor b;
    layer0_outputs(4767) <= not (a or b);
    layer0_outputs(4768) <= a and b;
    layer0_outputs(4769) <= not (a or b);
    layer0_outputs(4770) <= a xor b;
    layer0_outputs(4771) <= a or b;
    layer0_outputs(4772) <= b and not a;
    layer0_outputs(4773) <= not b or a;
    layer0_outputs(4774) <= b and not a;
    layer0_outputs(4775) <= a;
    layer0_outputs(4776) <= not (a and b);
    layer0_outputs(4777) <= a or b;
    layer0_outputs(4778) <= not a or b;
    layer0_outputs(4779) <= b and not a;
    layer0_outputs(4780) <= not (a xor b);
    layer0_outputs(4781) <= b;
    layer0_outputs(4782) <= b and not a;
    layer0_outputs(4783) <= b;
    layer0_outputs(4784) <= a xor b;
    layer0_outputs(4785) <= b;
    layer0_outputs(4786) <= b and not a;
    layer0_outputs(4787) <= not (a or b);
    layer0_outputs(4788) <= '1';
    layer0_outputs(4789) <= a and not b;
    layer0_outputs(4790) <= a or b;
    layer0_outputs(4791) <= not a;
    layer0_outputs(4792) <= not a;
    layer0_outputs(4793) <= a xor b;
    layer0_outputs(4794) <= '1';
    layer0_outputs(4795) <= '1';
    layer0_outputs(4796) <= a xor b;
    layer0_outputs(4797) <= b and not a;
    layer0_outputs(4798) <= a and b;
    layer0_outputs(4799) <= not b;
    layer0_outputs(4800) <= a or b;
    layer0_outputs(4801) <= not b;
    layer0_outputs(4802) <= b and not a;
    layer0_outputs(4803) <= not b or a;
    layer0_outputs(4804) <= not a;
    layer0_outputs(4805) <= b;
    layer0_outputs(4806) <= '1';
    layer0_outputs(4807) <= not b;
    layer0_outputs(4808) <= not (a xor b);
    layer0_outputs(4809) <= not b;
    layer0_outputs(4810) <= a and not b;
    layer0_outputs(4811) <= '0';
    layer0_outputs(4812) <= '1';
    layer0_outputs(4813) <= not b or a;
    layer0_outputs(4814) <= not b;
    layer0_outputs(4815) <= '0';
    layer0_outputs(4816) <= not (a xor b);
    layer0_outputs(4817) <= a;
    layer0_outputs(4818) <= not (a or b);
    layer0_outputs(4819) <= not (a or b);
    layer0_outputs(4820) <= a or b;
    layer0_outputs(4821) <= not b;
    layer0_outputs(4822) <= a;
    layer0_outputs(4823) <= not (a or b);
    layer0_outputs(4824) <= a or b;
    layer0_outputs(4825) <= not (a xor b);
    layer0_outputs(4826) <= not a;
    layer0_outputs(4827) <= not (a and b);
    layer0_outputs(4828) <= not a;
    layer0_outputs(4829) <= a;
    layer0_outputs(4830) <= not (a xor b);
    layer0_outputs(4831) <= not a or b;
    layer0_outputs(4832) <= not (a or b);
    layer0_outputs(4833) <= a xor b;
    layer0_outputs(4834) <= not (a xor b);
    layer0_outputs(4835) <= a and not b;
    layer0_outputs(4836) <= not (a or b);
    layer0_outputs(4837) <= '0';
    layer0_outputs(4838) <= not a;
    layer0_outputs(4839) <= a or b;
    layer0_outputs(4840) <= not b or a;
    layer0_outputs(4841) <= not (a or b);
    layer0_outputs(4842) <= a or b;
    layer0_outputs(4843) <= a;
    layer0_outputs(4844) <= b;
    layer0_outputs(4845) <= b;
    layer0_outputs(4846) <= not b;
    layer0_outputs(4847) <= a or b;
    layer0_outputs(4848) <= not (a or b);
    layer0_outputs(4849) <= b and not a;
    layer0_outputs(4850) <= not (a or b);
    layer0_outputs(4851) <= a and not b;
    layer0_outputs(4852) <= not (a xor b);
    layer0_outputs(4853) <= b;
    layer0_outputs(4854) <= a and not b;
    layer0_outputs(4855) <= not a;
    layer0_outputs(4856) <= not b or a;
    layer0_outputs(4857) <= not a or b;
    layer0_outputs(4858) <= not (a or b);
    layer0_outputs(4859) <= a;
    layer0_outputs(4860) <= a and b;
    layer0_outputs(4861) <= a xor b;
    layer0_outputs(4862) <= a xor b;
    layer0_outputs(4863) <= not a or b;
    layer0_outputs(4864) <= a and b;
    layer0_outputs(4865) <= not a or b;
    layer0_outputs(4866) <= not a;
    layer0_outputs(4867) <= not a or b;
    layer0_outputs(4868) <= not b or a;
    layer0_outputs(4869) <= a or b;
    layer0_outputs(4870) <= not b or a;
    layer0_outputs(4871) <= a or b;
    layer0_outputs(4872) <= a or b;
    layer0_outputs(4873) <= a or b;
    layer0_outputs(4874) <= a or b;
    layer0_outputs(4875) <= a or b;
    layer0_outputs(4876) <= not b;
    layer0_outputs(4877) <= not a or b;
    layer0_outputs(4878) <= a;
    layer0_outputs(4879) <= not a;
    layer0_outputs(4880) <= a;
    layer0_outputs(4881) <= a and not b;
    layer0_outputs(4882) <= a xor b;
    layer0_outputs(4883) <= not a or b;
    layer0_outputs(4884) <= b and not a;
    layer0_outputs(4885) <= not a or b;
    layer0_outputs(4886) <= b and not a;
    layer0_outputs(4887) <= b and not a;
    layer0_outputs(4888) <= '1';
    layer0_outputs(4889) <= '0';
    layer0_outputs(4890) <= a or b;
    layer0_outputs(4891) <= not (a or b);
    layer0_outputs(4892) <= not a;
    layer0_outputs(4893) <= not (a or b);
    layer0_outputs(4894) <= not b or a;
    layer0_outputs(4895) <= '1';
    layer0_outputs(4896) <= a xor b;
    layer0_outputs(4897) <= b;
    layer0_outputs(4898) <= not b;
    layer0_outputs(4899) <= a xor b;
    layer0_outputs(4900) <= b;
    layer0_outputs(4901) <= not (a and b);
    layer0_outputs(4902) <= a or b;
    layer0_outputs(4903) <= b and not a;
    layer0_outputs(4904) <= not (a or b);
    layer0_outputs(4905) <= b;
    layer0_outputs(4906) <= '0';
    layer0_outputs(4907) <= not b;
    layer0_outputs(4908) <= not (a or b);
    layer0_outputs(4909) <= a xor b;
    layer0_outputs(4910) <= a and b;
    layer0_outputs(4911) <= a xor b;
    layer0_outputs(4912) <= a;
    layer0_outputs(4913) <= a;
    layer0_outputs(4914) <= not (a xor b);
    layer0_outputs(4915) <= not b;
    layer0_outputs(4916) <= not (a xor b);
    layer0_outputs(4917) <= not b or a;
    layer0_outputs(4918) <= a;
    layer0_outputs(4919) <= not (a xor b);
    layer0_outputs(4920) <= not (a or b);
    layer0_outputs(4921) <= not (a xor b);
    layer0_outputs(4922) <= a or b;
    layer0_outputs(4923) <= a and not b;
    layer0_outputs(4924) <= '0';
    layer0_outputs(4925) <= not b or a;
    layer0_outputs(4926) <= not (a xor b);
    layer0_outputs(4927) <= a or b;
    layer0_outputs(4928) <= b and not a;
    layer0_outputs(4929) <= a and not b;
    layer0_outputs(4930) <= not a;
    layer0_outputs(4931) <= not a;
    layer0_outputs(4932) <= not b or a;
    layer0_outputs(4933) <= '1';
    layer0_outputs(4934) <= b;
    layer0_outputs(4935) <= a or b;
    layer0_outputs(4936) <= a xor b;
    layer0_outputs(4937) <= not (a or b);
    layer0_outputs(4938) <= '1';
    layer0_outputs(4939) <= a and b;
    layer0_outputs(4940) <= a;
    layer0_outputs(4941) <= not b or a;
    layer0_outputs(4942) <= not (a or b);
    layer0_outputs(4943) <= not b;
    layer0_outputs(4944) <= b and not a;
    layer0_outputs(4945) <= a or b;
    layer0_outputs(4946) <= a xor b;
    layer0_outputs(4947) <= a;
    layer0_outputs(4948) <= '1';
    layer0_outputs(4949) <= '0';
    layer0_outputs(4950) <= b and not a;
    layer0_outputs(4951) <= not a;
    layer0_outputs(4952) <= a or b;
    layer0_outputs(4953) <= not a or b;
    layer0_outputs(4954) <= not a or b;
    layer0_outputs(4955) <= not (a xor b);
    layer0_outputs(4956) <= not (a or b);
    layer0_outputs(4957) <= b;
    layer0_outputs(4958) <= not (a xor b);
    layer0_outputs(4959) <= b and not a;
    layer0_outputs(4960) <= a or b;
    layer0_outputs(4961) <= not (a or b);
    layer0_outputs(4962) <= a xor b;
    layer0_outputs(4963) <= a or b;
    layer0_outputs(4964) <= a;
    layer0_outputs(4965) <= a and b;
    layer0_outputs(4966) <= not b;
    layer0_outputs(4967) <= '0';
    layer0_outputs(4968) <= not a;
    layer0_outputs(4969) <= not (a or b);
    layer0_outputs(4970) <= '1';
    layer0_outputs(4971) <= not (a or b);
    layer0_outputs(4972) <= not b;
    layer0_outputs(4973) <= '1';
    layer0_outputs(4974) <= b and not a;
    layer0_outputs(4975) <= a and not b;
    layer0_outputs(4976) <= b and not a;
    layer0_outputs(4977) <= not a or b;
    layer0_outputs(4978) <= a or b;
    layer0_outputs(4979) <= a;
    layer0_outputs(4980) <= a and b;
    layer0_outputs(4981) <= b and not a;
    layer0_outputs(4982) <= not b or a;
    layer0_outputs(4983) <= a and b;
    layer0_outputs(4984) <= a;
    layer0_outputs(4985) <= not b or a;
    layer0_outputs(4986) <= b and not a;
    layer0_outputs(4987) <= not (a or b);
    layer0_outputs(4988) <= not (a or b);
    layer0_outputs(4989) <= b;
    layer0_outputs(4990) <= not b or a;
    layer0_outputs(4991) <= not (a or b);
    layer0_outputs(4992) <= b and not a;
    layer0_outputs(4993) <= not (a and b);
    layer0_outputs(4994) <= not b or a;
    layer0_outputs(4995) <= not (a and b);
    layer0_outputs(4996) <= a and not b;
    layer0_outputs(4997) <= not b or a;
    layer0_outputs(4998) <= a or b;
    layer0_outputs(4999) <= b and not a;
    layer0_outputs(5000) <= not b or a;
    layer0_outputs(5001) <= a or b;
    layer0_outputs(5002) <= not b or a;
    layer0_outputs(5003) <= a xor b;
    layer0_outputs(5004) <= a xor b;
    layer0_outputs(5005) <= not b or a;
    layer0_outputs(5006) <= '1';
    layer0_outputs(5007) <= not (a or b);
    layer0_outputs(5008) <= not a or b;
    layer0_outputs(5009) <= not b;
    layer0_outputs(5010) <= b;
    layer0_outputs(5011) <= '1';
    layer0_outputs(5012) <= '1';
    layer0_outputs(5013) <= not (a or b);
    layer0_outputs(5014) <= not a or b;
    layer0_outputs(5015) <= a;
    layer0_outputs(5016) <= not (a xor b);
    layer0_outputs(5017) <= a;
    layer0_outputs(5018) <= not (a or b);
    layer0_outputs(5019) <= b and not a;
    layer0_outputs(5020) <= a or b;
    layer0_outputs(5021) <= a and b;
    layer0_outputs(5022) <= not b;
    layer0_outputs(5023) <= not (a xor b);
    layer0_outputs(5024) <= '0';
    layer0_outputs(5025) <= not a or b;
    layer0_outputs(5026) <= a and not b;
    layer0_outputs(5027) <= a and b;
    layer0_outputs(5028) <= not (a or b);
    layer0_outputs(5029) <= '0';
    layer0_outputs(5030) <= not b;
    layer0_outputs(5031) <= a or b;
    layer0_outputs(5032) <= not (a xor b);
    layer0_outputs(5033) <= b and not a;
    layer0_outputs(5034) <= not (a and b);
    layer0_outputs(5035) <= not b or a;
    layer0_outputs(5036) <= not a or b;
    layer0_outputs(5037) <= a and not b;
    layer0_outputs(5038) <= not (a or b);
    layer0_outputs(5039) <= a;
    layer0_outputs(5040) <= not (a or b);
    layer0_outputs(5041) <= a and not b;
    layer0_outputs(5042) <= a and b;
    layer0_outputs(5043) <= a or b;
    layer0_outputs(5044) <= a and b;
    layer0_outputs(5045) <= not b or a;
    layer0_outputs(5046) <= b and not a;
    layer0_outputs(5047) <= b and not a;
    layer0_outputs(5048) <= not b or a;
    layer0_outputs(5049) <= '1';
    layer0_outputs(5050) <= a or b;
    layer0_outputs(5051) <= not a;
    layer0_outputs(5052) <= not (a xor b);
    layer0_outputs(5053) <= b;
    layer0_outputs(5054) <= a;
    layer0_outputs(5055) <= a and not b;
    layer0_outputs(5056) <= not (a or b);
    layer0_outputs(5057) <= a xor b;
    layer0_outputs(5058) <= not (a or b);
    layer0_outputs(5059) <= not a or b;
    layer0_outputs(5060) <= a and not b;
    layer0_outputs(5061) <= '1';
    layer0_outputs(5062) <= b;
    layer0_outputs(5063) <= '0';
    layer0_outputs(5064) <= not a;
    layer0_outputs(5065) <= b;
    layer0_outputs(5066) <= a and not b;
    layer0_outputs(5067) <= '1';
    layer0_outputs(5068) <= a or b;
    layer0_outputs(5069) <= a or b;
    layer0_outputs(5070) <= not a;
    layer0_outputs(5071) <= b and not a;
    layer0_outputs(5072) <= not (a xor b);
    layer0_outputs(5073) <= not a;
    layer0_outputs(5074) <= a;
    layer0_outputs(5075) <= not a or b;
    layer0_outputs(5076) <= not (a or b);
    layer0_outputs(5077) <= a and not b;
    layer0_outputs(5078) <= not (a or b);
    layer0_outputs(5079) <= not a;
    layer0_outputs(5080) <= '1';
    layer0_outputs(5081) <= not a or b;
    layer0_outputs(5082) <= not b;
    layer0_outputs(5083) <= not (a or b);
    layer0_outputs(5084) <= a and b;
    layer0_outputs(5085) <= a and not b;
    layer0_outputs(5086) <= not (a and b);
    layer0_outputs(5087) <= not a or b;
    layer0_outputs(5088) <= a and b;
    layer0_outputs(5089) <= a;
    layer0_outputs(5090) <= a and not b;
    layer0_outputs(5091) <= b and not a;
    layer0_outputs(5092) <= a xor b;
    layer0_outputs(5093) <= b and not a;
    layer0_outputs(5094) <= a xor b;
    layer0_outputs(5095) <= b;
    layer0_outputs(5096) <= not a;
    layer0_outputs(5097) <= b;
    layer0_outputs(5098) <= '1';
    layer0_outputs(5099) <= not (a or b);
    layer0_outputs(5100) <= not (a or b);
    layer0_outputs(5101) <= b and not a;
    layer0_outputs(5102) <= a and not b;
    layer0_outputs(5103) <= not b;
    layer0_outputs(5104) <= not (a or b);
    layer0_outputs(5105) <= a or b;
    layer0_outputs(5106) <= not b;
    layer0_outputs(5107) <= a and not b;
    layer0_outputs(5108) <= b;
    layer0_outputs(5109) <= not a;
    layer0_outputs(5110) <= not (a or b);
    layer0_outputs(5111) <= not a;
    layer0_outputs(5112) <= b;
    layer0_outputs(5113) <= not (a or b);
    layer0_outputs(5114) <= b and not a;
    layer0_outputs(5115) <= not (a and b);
    layer0_outputs(5116) <= a;
    layer0_outputs(5117) <= not (a xor b);
    layer0_outputs(5118) <= a or b;
    layer0_outputs(5119) <= not (a or b);
    layer1_outputs(0) <= not (a or b);
    layer1_outputs(1) <= not (a and b);
    layer1_outputs(2) <= not (a xor b);
    layer1_outputs(3) <= a;
    layer1_outputs(4) <= b;
    layer1_outputs(5) <= not b or a;
    layer1_outputs(6) <= a and not b;
    layer1_outputs(7) <= a or b;
    layer1_outputs(8) <= b and not a;
    layer1_outputs(9) <= not (a and b);
    layer1_outputs(10) <= not b;
    layer1_outputs(11) <= not (a and b);
    layer1_outputs(12) <= a and b;
    layer1_outputs(13) <= a;
    layer1_outputs(14) <= b;
    layer1_outputs(15) <= '1';
    layer1_outputs(16) <= not b;
    layer1_outputs(17) <= not (a and b);
    layer1_outputs(18) <= a;
    layer1_outputs(19) <= a or b;
    layer1_outputs(20) <= b;
    layer1_outputs(21) <= not (a xor b);
    layer1_outputs(22) <= not b or a;
    layer1_outputs(23) <= a and b;
    layer1_outputs(24) <= b and not a;
    layer1_outputs(25) <= not b;
    layer1_outputs(26) <= not b;
    layer1_outputs(27) <= not a;
    layer1_outputs(28) <= b;
    layer1_outputs(29) <= a and b;
    layer1_outputs(30) <= '1';
    layer1_outputs(31) <= a or b;
    layer1_outputs(32) <= a or b;
    layer1_outputs(33) <= a;
    layer1_outputs(34) <= not a or b;
    layer1_outputs(35) <= not b or a;
    layer1_outputs(36) <= not (a or b);
    layer1_outputs(37) <= not (a and b);
    layer1_outputs(38) <= a xor b;
    layer1_outputs(39) <= a and not b;
    layer1_outputs(40) <= a;
    layer1_outputs(41) <= not (a and b);
    layer1_outputs(42) <= not (a or b);
    layer1_outputs(43) <= a and not b;
    layer1_outputs(44) <= b and not a;
    layer1_outputs(45) <= a and not b;
    layer1_outputs(46) <= not (a xor b);
    layer1_outputs(47) <= not a;
    layer1_outputs(48) <= not b or a;
    layer1_outputs(49) <= '0';
    layer1_outputs(50) <= a and not b;
    layer1_outputs(51) <= a or b;
    layer1_outputs(52) <= b and not a;
    layer1_outputs(53) <= not b;
    layer1_outputs(54) <= a or b;
    layer1_outputs(55) <= b and not a;
    layer1_outputs(56) <= not b;
    layer1_outputs(57) <= not (a and b);
    layer1_outputs(58) <= not b;
    layer1_outputs(59) <= a and not b;
    layer1_outputs(60) <= a and not b;
    layer1_outputs(61) <= not b;
    layer1_outputs(62) <= b;
    layer1_outputs(63) <= not (a and b);
    layer1_outputs(64) <= not a;
    layer1_outputs(65) <= not a or b;
    layer1_outputs(66) <= a;
    layer1_outputs(67) <= not a;
    layer1_outputs(68) <= not (a and b);
    layer1_outputs(69) <= not (a and b);
    layer1_outputs(70) <= not b;
    layer1_outputs(71) <= '1';
    layer1_outputs(72) <= not (a or b);
    layer1_outputs(73) <= not b;
    layer1_outputs(74) <= '0';
    layer1_outputs(75) <= a and b;
    layer1_outputs(76) <= not b or a;
    layer1_outputs(77) <= b;
    layer1_outputs(78) <= b and not a;
    layer1_outputs(79) <= a and not b;
    layer1_outputs(80) <= '0';
    layer1_outputs(81) <= not b or a;
    layer1_outputs(82) <= not b;
    layer1_outputs(83) <= not (a xor b);
    layer1_outputs(84) <= a and not b;
    layer1_outputs(85) <= not (a or b);
    layer1_outputs(86) <= b and not a;
    layer1_outputs(87) <= a and b;
    layer1_outputs(88) <= not b;
    layer1_outputs(89) <= a and b;
    layer1_outputs(90) <= not (a or b);
    layer1_outputs(91) <= b;
    layer1_outputs(92) <= a;
    layer1_outputs(93) <= not b;
    layer1_outputs(94) <= not (a and b);
    layer1_outputs(95) <= '1';
    layer1_outputs(96) <= a and b;
    layer1_outputs(97) <= b;
    layer1_outputs(98) <= a xor b;
    layer1_outputs(99) <= a;
    layer1_outputs(100) <= a and not b;
    layer1_outputs(101) <= b and not a;
    layer1_outputs(102) <= not a;
    layer1_outputs(103) <= a;
    layer1_outputs(104) <= not (a and b);
    layer1_outputs(105) <= not a or b;
    layer1_outputs(106) <= b;
    layer1_outputs(107) <= not a or b;
    layer1_outputs(108) <= a and b;
    layer1_outputs(109) <= a and b;
    layer1_outputs(110) <= a and b;
    layer1_outputs(111) <= b;
    layer1_outputs(112) <= '1';
    layer1_outputs(113) <= not b;
    layer1_outputs(114) <= b;
    layer1_outputs(115) <= a;
    layer1_outputs(116) <= not b or a;
    layer1_outputs(117) <= not a;
    layer1_outputs(118) <= not (a xor b);
    layer1_outputs(119) <= a and not b;
    layer1_outputs(120) <= b and not a;
    layer1_outputs(121) <= a xor b;
    layer1_outputs(122) <= not a;
    layer1_outputs(123) <= a and b;
    layer1_outputs(124) <= not a;
    layer1_outputs(125) <= a and not b;
    layer1_outputs(126) <= not b;
    layer1_outputs(127) <= not b;
    layer1_outputs(128) <= a and b;
    layer1_outputs(129) <= a and b;
    layer1_outputs(130) <= not a;
    layer1_outputs(131) <= a xor b;
    layer1_outputs(132) <= a or b;
    layer1_outputs(133) <= not b;
    layer1_outputs(134) <= b and not a;
    layer1_outputs(135) <= a;
    layer1_outputs(136) <= b and not a;
    layer1_outputs(137) <= a or b;
    layer1_outputs(138) <= not a or b;
    layer1_outputs(139) <= not b;
    layer1_outputs(140) <= not (a and b);
    layer1_outputs(141) <= not a;
    layer1_outputs(142) <= b;
    layer1_outputs(143) <= a and not b;
    layer1_outputs(144) <= b and not a;
    layer1_outputs(145) <= a and b;
    layer1_outputs(146) <= '0';
    layer1_outputs(147) <= a;
    layer1_outputs(148) <= a and not b;
    layer1_outputs(149) <= '0';
    layer1_outputs(150) <= not a or b;
    layer1_outputs(151) <= a and not b;
    layer1_outputs(152) <= not b;
    layer1_outputs(153) <= a or b;
    layer1_outputs(154) <= a;
    layer1_outputs(155) <= not (a xor b);
    layer1_outputs(156) <= a xor b;
    layer1_outputs(157) <= a or b;
    layer1_outputs(158) <= '0';
    layer1_outputs(159) <= a and b;
    layer1_outputs(160) <= a and b;
    layer1_outputs(161) <= not b;
    layer1_outputs(162) <= a and b;
    layer1_outputs(163) <= not a or b;
    layer1_outputs(164) <= not a;
    layer1_outputs(165) <= a;
    layer1_outputs(166) <= not a;
    layer1_outputs(167) <= a and b;
    layer1_outputs(168) <= '0';
    layer1_outputs(169) <= not a;
    layer1_outputs(170) <= not b;
    layer1_outputs(171) <= b;
    layer1_outputs(172) <= not (a or b);
    layer1_outputs(173) <= not b or a;
    layer1_outputs(174) <= not b;
    layer1_outputs(175) <= not a or b;
    layer1_outputs(176) <= not b or a;
    layer1_outputs(177) <= not b;
    layer1_outputs(178) <= b and not a;
    layer1_outputs(179) <= a;
    layer1_outputs(180) <= not b or a;
    layer1_outputs(181) <= b;
    layer1_outputs(182) <= a and b;
    layer1_outputs(183) <= a or b;
    layer1_outputs(184) <= not b or a;
    layer1_outputs(185) <= a xor b;
    layer1_outputs(186) <= a or b;
    layer1_outputs(187) <= a;
    layer1_outputs(188) <= a;
    layer1_outputs(189) <= not b;
    layer1_outputs(190) <= not a or b;
    layer1_outputs(191) <= a and not b;
    layer1_outputs(192) <= not (a and b);
    layer1_outputs(193) <= a;
    layer1_outputs(194) <= a xor b;
    layer1_outputs(195) <= not a;
    layer1_outputs(196) <= '1';
    layer1_outputs(197) <= not a;
    layer1_outputs(198) <= b and not a;
    layer1_outputs(199) <= not (a and b);
    layer1_outputs(200) <= a or b;
    layer1_outputs(201) <= not (a and b);
    layer1_outputs(202) <= not b;
    layer1_outputs(203) <= b;
    layer1_outputs(204) <= b and not a;
    layer1_outputs(205) <= not a or b;
    layer1_outputs(206) <= not a;
    layer1_outputs(207) <= not a;
    layer1_outputs(208) <= not (a or b);
    layer1_outputs(209) <= not a;
    layer1_outputs(210) <= b;
    layer1_outputs(211) <= a xor b;
    layer1_outputs(212) <= not a;
    layer1_outputs(213) <= not b;
    layer1_outputs(214) <= a and not b;
    layer1_outputs(215) <= a or b;
    layer1_outputs(216) <= a xor b;
    layer1_outputs(217) <= '0';
    layer1_outputs(218) <= b;
    layer1_outputs(219) <= b and not a;
    layer1_outputs(220) <= b;
    layer1_outputs(221) <= not a;
    layer1_outputs(222) <= a and not b;
    layer1_outputs(223) <= b;
    layer1_outputs(224) <= not a or b;
    layer1_outputs(225) <= a;
    layer1_outputs(226) <= b;
    layer1_outputs(227) <= a and not b;
    layer1_outputs(228) <= not a or b;
    layer1_outputs(229) <= b and not a;
    layer1_outputs(230) <= a;
    layer1_outputs(231) <= a and b;
    layer1_outputs(232) <= a and b;
    layer1_outputs(233) <= not a;
    layer1_outputs(234) <= a;
    layer1_outputs(235) <= not (a and b);
    layer1_outputs(236) <= a and b;
    layer1_outputs(237) <= not a or b;
    layer1_outputs(238) <= a;
    layer1_outputs(239) <= a;
    layer1_outputs(240) <= not (a xor b);
    layer1_outputs(241) <= b;
    layer1_outputs(242) <= a;
    layer1_outputs(243) <= not a;
    layer1_outputs(244) <= a or b;
    layer1_outputs(245) <= not b or a;
    layer1_outputs(246) <= b;
    layer1_outputs(247) <= a and b;
    layer1_outputs(248) <= a or b;
    layer1_outputs(249) <= b;
    layer1_outputs(250) <= a and not b;
    layer1_outputs(251) <= not (a or b);
    layer1_outputs(252) <= b;
    layer1_outputs(253) <= not a;
    layer1_outputs(254) <= b;
    layer1_outputs(255) <= not a;
    layer1_outputs(256) <= not a or b;
    layer1_outputs(257) <= not (a and b);
    layer1_outputs(258) <= a xor b;
    layer1_outputs(259) <= a and b;
    layer1_outputs(260) <= b;
    layer1_outputs(261) <= not (a xor b);
    layer1_outputs(262) <= not b;
    layer1_outputs(263) <= not (a and b);
    layer1_outputs(264) <= not b;
    layer1_outputs(265) <= not (a or b);
    layer1_outputs(266) <= not (a or b);
    layer1_outputs(267) <= a and b;
    layer1_outputs(268) <= a;
    layer1_outputs(269) <= not a;
    layer1_outputs(270) <= b and not a;
    layer1_outputs(271) <= not b;
    layer1_outputs(272) <= a xor b;
    layer1_outputs(273) <= b;
    layer1_outputs(274) <= a and b;
    layer1_outputs(275) <= a and not b;
    layer1_outputs(276) <= '0';
    layer1_outputs(277) <= b;
    layer1_outputs(278) <= a;
    layer1_outputs(279) <= a;
    layer1_outputs(280) <= a or b;
    layer1_outputs(281) <= not a or b;
    layer1_outputs(282) <= not (a and b);
    layer1_outputs(283) <= not a or b;
    layer1_outputs(284) <= b;
    layer1_outputs(285) <= a and not b;
    layer1_outputs(286) <= b and not a;
    layer1_outputs(287) <= b;
    layer1_outputs(288) <= not b or a;
    layer1_outputs(289) <= not a;
    layer1_outputs(290) <= b and not a;
    layer1_outputs(291) <= not (a and b);
    layer1_outputs(292) <= a or b;
    layer1_outputs(293) <= a or b;
    layer1_outputs(294) <= a and not b;
    layer1_outputs(295) <= not b;
    layer1_outputs(296) <= a or b;
    layer1_outputs(297) <= '1';
    layer1_outputs(298) <= b and not a;
    layer1_outputs(299) <= not b or a;
    layer1_outputs(300) <= not (a and b);
    layer1_outputs(301) <= a xor b;
    layer1_outputs(302) <= a or b;
    layer1_outputs(303) <= not b;
    layer1_outputs(304) <= not (a xor b);
    layer1_outputs(305) <= not (a or b);
    layer1_outputs(306) <= not (a or b);
    layer1_outputs(307) <= not a;
    layer1_outputs(308) <= not (a xor b);
    layer1_outputs(309) <= a and not b;
    layer1_outputs(310) <= a;
    layer1_outputs(311) <= '0';
    layer1_outputs(312) <= not (a or b);
    layer1_outputs(313) <= not a;
    layer1_outputs(314) <= not b;
    layer1_outputs(315) <= not a;
    layer1_outputs(316) <= not (a and b);
    layer1_outputs(317) <= b;
    layer1_outputs(318) <= not b or a;
    layer1_outputs(319) <= not b;
    layer1_outputs(320) <= not b;
    layer1_outputs(321) <= not b;
    layer1_outputs(322) <= b and not a;
    layer1_outputs(323) <= a or b;
    layer1_outputs(324) <= a;
    layer1_outputs(325) <= b and not a;
    layer1_outputs(326) <= not (a and b);
    layer1_outputs(327) <= not b or a;
    layer1_outputs(328) <= not b;
    layer1_outputs(329) <= a;
    layer1_outputs(330) <= '1';
    layer1_outputs(331) <= a;
    layer1_outputs(332) <= not a;
    layer1_outputs(333) <= a and b;
    layer1_outputs(334) <= a and b;
    layer1_outputs(335) <= not b;
    layer1_outputs(336) <= b;
    layer1_outputs(337) <= not b;
    layer1_outputs(338) <= a and not b;
    layer1_outputs(339) <= b;
    layer1_outputs(340) <= a;
    layer1_outputs(341) <= a and not b;
    layer1_outputs(342) <= b;
    layer1_outputs(343) <= a or b;
    layer1_outputs(344) <= '0';
    layer1_outputs(345) <= '0';
    layer1_outputs(346) <= a and not b;
    layer1_outputs(347) <= b and not a;
    layer1_outputs(348) <= not (a and b);
    layer1_outputs(349) <= not b or a;
    layer1_outputs(350) <= b and not a;
    layer1_outputs(351) <= not a or b;
    layer1_outputs(352) <= not b;
    layer1_outputs(353) <= not b;
    layer1_outputs(354) <= not (a xor b);
    layer1_outputs(355) <= not (a and b);
    layer1_outputs(356) <= '1';
    layer1_outputs(357) <= b;
    layer1_outputs(358) <= a or b;
    layer1_outputs(359) <= a;
    layer1_outputs(360) <= b and not a;
    layer1_outputs(361) <= '1';
    layer1_outputs(362) <= a or b;
    layer1_outputs(363) <= a;
    layer1_outputs(364) <= b and not a;
    layer1_outputs(365) <= a and not b;
    layer1_outputs(366) <= a;
    layer1_outputs(367) <= a xor b;
    layer1_outputs(368) <= a;
    layer1_outputs(369) <= not a or b;
    layer1_outputs(370) <= not b;
    layer1_outputs(371) <= b and not a;
    layer1_outputs(372) <= not a;
    layer1_outputs(373) <= not a or b;
    layer1_outputs(374) <= not b;
    layer1_outputs(375) <= not a;
    layer1_outputs(376) <= a;
    layer1_outputs(377) <= a and b;
    layer1_outputs(378) <= a;
    layer1_outputs(379) <= a and not b;
    layer1_outputs(380) <= not b or a;
    layer1_outputs(381) <= not a;
    layer1_outputs(382) <= b and not a;
    layer1_outputs(383) <= not b;
    layer1_outputs(384) <= b;
    layer1_outputs(385) <= not b;
    layer1_outputs(386) <= a;
    layer1_outputs(387) <= b;
    layer1_outputs(388) <= not b or a;
    layer1_outputs(389) <= a or b;
    layer1_outputs(390) <= b;
    layer1_outputs(391) <= not b or a;
    layer1_outputs(392) <= a and not b;
    layer1_outputs(393) <= a and not b;
    layer1_outputs(394) <= a and b;
    layer1_outputs(395) <= not b;
    layer1_outputs(396) <= not (a and b);
    layer1_outputs(397) <= not a or b;
    layer1_outputs(398) <= not (a xor b);
    layer1_outputs(399) <= a;
    layer1_outputs(400) <= not (a and b);
    layer1_outputs(401) <= a and not b;
    layer1_outputs(402) <= '0';
    layer1_outputs(403) <= '1';
    layer1_outputs(404) <= not (a and b);
    layer1_outputs(405) <= not b;
    layer1_outputs(406) <= a or b;
    layer1_outputs(407) <= a xor b;
    layer1_outputs(408) <= not b;
    layer1_outputs(409) <= a xor b;
    layer1_outputs(410) <= a or b;
    layer1_outputs(411) <= not (a and b);
    layer1_outputs(412) <= not (a and b);
    layer1_outputs(413) <= not a or b;
    layer1_outputs(414) <= a and b;
    layer1_outputs(415) <= '0';
    layer1_outputs(416) <= not (a and b);
    layer1_outputs(417) <= '0';
    layer1_outputs(418) <= b and not a;
    layer1_outputs(419) <= not b or a;
    layer1_outputs(420) <= a and not b;
    layer1_outputs(421) <= not a or b;
    layer1_outputs(422) <= not a;
    layer1_outputs(423) <= not (a xor b);
    layer1_outputs(424) <= not a;
    layer1_outputs(425) <= b;
    layer1_outputs(426) <= a;
    layer1_outputs(427) <= not (a or b);
    layer1_outputs(428) <= a and b;
    layer1_outputs(429) <= not a;
    layer1_outputs(430) <= a and not b;
    layer1_outputs(431) <= b;
    layer1_outputs(432) <= not (a or b);
    layer1_outputs(433) <= b;
    layer1_outputs(434) <= b and not a;
    layer1_outputs(435) <= b;
    layer1_outputs(436) <= b and not a;
    layer1_outputs(437) <= b;
    layer1_outputs(438) <= not a or b;
    layer1_outputs(439) <= a and not b;
    layer1_outputs(440) <= b;
    layer1_outputs(441) <= not (a and b);
    layer1_outputs(442) <= a and b;
    layer1_outputs(443) <= b and not a;
    layer1_outputs(444) <= not (a and b);
    layer1_outputs(445) <= '0';
    layer1_outputs(446) <= not (a or b);
    layer1_outputs(447) <= b and not a;
    layer1_outputs(448) <= not b or a;
    layer1_outputs(449) <= not b;
    layer1_outputs(450) <= b and not a;
    layer1_outputs(451) <= a and b;
    layer1_outputs(452) <= b and not a;
    layer1_outputs(453) <= not a;
    layer1_outputs(454) <= '1';
    layer1_outputs(455) <= b;
    layer1_outputs(456) <= a xor b;
    layer1_outputs(457) <= not a;
    layer1_outputs(458) <= not (a or b);
    layer1_outputs(459) <= not a or b;
    layer1_outputs(460) <= a and not b;
    layer1_outputs(461) <= b and not a;
    layer1_outputs(462) <= a or b;
    layer1_outputs(463) <= a or b;
    layer1_outputs(464) <= not (a and b);
    layer1_outputs(465) <= not a;
    layer1_outputs(466) <= not (a and b);
    layer1_outputs(467) <= b;
    layer1_outputs(468) <= not a;
    layer1_outputs(469) <= a;
    layer1_outputs(470) <= not b;
    layer1_outputs(471) <= b;
    layer1_outputs(472) <= a and b;
    layer1_outputs(473) <= not b;
    layer1_outputs(474) <= '1';
    layer1_outputs(475) <= not a or b;
    layer1_outputs(476) <= not (a and b);
    layer1_outputs(477) <= a;
    layer1_outputs(478) <= b;
    layer1_outputs(479) <= a xor b;
    layer1_outputs(480) <= not a or b;
    layer1_outputs(481) <= not a;
    layer1_outputs(482) <= not b;
    layer1_outputs(483) <= a and b;
    layer1_outputs(484) <= b;
    layer1_outputs(485) <= not (a or b);
    layer1_outputs(486) <= b and not a;
    layer1_outputs(487) <= a and b;
    layer1_outputs(488) <= not a;
    layer1_outputs(489) <= b;
    layer1_outputs(490) <= not b;
    layer1_outputs(491) <= not (a and b);
    layer1_outputs(492) <= b and not a;
    layer1_outputs(493) <= '1';
    layer1_outputs(494) <= a or b;
    layer1_outputs(495) <= not b;
    layer1_outputs(496) <= not (a xor b);
    layer1_outputs(497) <= not (a and b);
    layer1_outputs(498) <= a or b;
    layer1_outputs(499) <= a;
    layer1_outputs(500) <= not a;
    layer1_outputs(501) <= a and not b;
    layer1_outputs(502) <= b;
    layer1_outputs(503) <= a;
    layer1_outputs(504) <= a xor b;
    layer1_outputs(505) <= not a or b;
    layer1_outputs(506) <= not b;
    layer1_outputs(507) <= b;
    layer1_outputs(508) <= a or b;
    layer1_outputs(509) <= not a;
    layer1_outputs(510) <= '0';
    layer1_outputs(511) <= not a or b;
    layer1_outputs(512) <= a and b;
    layer1_outputs(513) <= not a;
    layer1_outputs(514) <= a;
    layer1_outputs(515) <= not (a and b);
    layer1_outputs(516) <= not (a xor b);
    layer1_outputs(517) <= b;
    layer1_outputs(518) <= b;
    layer1_outputs(519) <= not b or a;
    layer1_outputs(520) <= '0';
    layer1_outputs(521) <= not b;
    layer1_outputs(522) <= a and not b;
    layer1_outputs(523) <= a;
    layer1_outputs(524) <= b and not a;
    layer1_outputs(525) <= b;
    layer1_outputs(526) <= not b;
    layer1_outputs(527) <= a or b;
    layer1_outputs(528) <= not b or a;
    layer1_outputs(529) <= '0';
    layer1_outputs(530) <= not b;
    layer1_outputs(531) <= not b or a;
    layer1_outputs(532) <= a and b;
    layer1_outputs(533) <= not b or a;
    layer1_outputs(534) <= not (a and b);
    layer1_outputs(535) <= b and not a;
    layer1_outputs(536) <= b;
    layer1_outputs(537) <= not b or a;
    layer1_outputs(538) <= '1';
    layer1_outputs(539) <= a;
    layer1_outputs(540) <= b;
    layer1_outputs(541) <= b;
    layer1_outputs(542) <= a and not b;
    layer1_outputs(543) <= not b or a;
    layer1_outputs(544) <= a xor b;
    layer1_outputs(545) <= a or b;
    layer1_outputs(546) <= '0';
    layer1_outputs(547) <= a and not b;
    layer1_outputs(548) <= b;
    layer1_outputs(549) <= a;
    layer1_outputs(550) <= b and not a;
    layer1_outputs(551) <= not (a and b);
    layer1_outputs(552) <= not (a xor b);
    layer1_outputs(553) <= a or b;
    layer1_outputs(554) <= '0';
    layer1_outputs(555) <= not a;
    layer1_outputs(556) <= b;
    layer1_outputs(557) <= not (a xor b);
    layer1_outputs(558) <= b;
    layer1_outputs(559) <= not (a xor b);
    layer1_outputs(560) <= not (a xor b);
    layer1_outputs(561) <= not a or b;
    layer1_outputs(562) <= a or b;
    layer1_outputs(563) <= b;
    layer1_outputs(564) <= b;
    layer1_outputs(565) <= a xor b;
    layer1_outputs(566) <= '1';
    layer1_outputs(567) <= b and not a;
    layer1_outputs(568) <= '0';
    layer1_outputs(569) <= '0';
    layer1_outputs(570) <= not b;
    layer1_outputs(571) <= a and b;
    layer1_outputs(572) <= a;
    layer1_outputs(573) <= not b;
    layer1_outputs(574) <= not b or a;
    layer1_outputs(575) <= not (a xor b);
    layer1_outputs(576) <= not a;
    layer1_outputs(577) <= b and not a;
    layer1_outputs(578) <= b;
    layer1_outputs(579) <= not a;
    layer1_outputs(580) <= '1';
    layer1_outputs(581) <= a or b;
    layer1_outputs(582) <= not (a and b);
    layer1_outputs(583) <= b and not a;
    layer1_outputs(584) <= not (a or b);
    layer1_outputs(585) <= a or b;
    layer1_outputs(586) <= not (a xor b);
    layer1_outputs(587) <= not (a or b);
    layer1_outputs(588) <= not b or a;
    layer1_outputs(589) <= not (a xor b);
    layer1_outputs(590) <= not b;
    layer1_outputs(591) <= not a;
    layer1_outputs(592) <= b;
    layer1_outputs(593) <= b and not a;
    layer1_outputs(594) <= not b;
    layer1_outputs(595) <= not (a or b);
    layer1_outputs(596) <= a and not b;
    layer1_outputs(597) <= '1';
    layer1_outputs(598) <= b;
    layer1_outputs(599) <= not (a and b);
    layer1_outputs(600) <= not (a xor b);
    layer1_outputs(601) <= a and b;
    layer1_outputs(602) <= not a or b;
    layer1_outputs(603) <= a;
    layer1_outputs(604) <= not b or a;
    layer1_outputs(605) <= a;
    layer1_outputs(606) <= a and not b;
    layer1_outputs(607) <= a and not b;
    layer1_outputs(608) <= a or b;
    layer1_outputs(609) <= '1';
    layer1_outputs(610) <= b;
    layer1_outputs(611) <= a and not b;
    layer1_outputs(612) <= a and b;
    layer1_outputs(613) <= not b or a;
    layer1_outputs(614) <= a and not b;
    layer1_outputs(615) <= not a;
    layer1_outputs(616) <= a and not b;
    layer1_outputs(617) <= not a;
    layer1_outputs(618) <= not a or b;
    layer1_outputs(619) <= b and not a;
    layer1_outputs(620) <= b;
    layer1_outputs(621) <= not (a or b);
    layer1_outputs(622) <= not b;
    layer1_outputs(623) <= not (a or b);
    layer1_outputs(624) <= not (a and b);
    layer1_outputs(625) <= '0';
    layer1_outputs(626) <= '0';
    layer1_outputs(627) <= not b;
    layer1_outputs(628) <= b;
    layer1_outputs(629) <= not a;
    layer1_outputs(630) <= not b;
    layer1_outputs(631) <= not a;
    layer1_outputs(632) <= a and b;
    layer1_outputs(633) <= not a or b;
    layer1_outputs(634) <= b and not a;
    layer1_outputs(635) <= a and b;
    layer1_outputs(636) <= a;
    layer1_outputs(637) <= not b;
    layer1_outputs(638) <= a or b;
    layer1_outputs(639) <= not (a and b);
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= not (a and b);
    layer1_outputs(642) <= not a or b;
    layer1_outputs(643) <= not a;
    layer1_outputs(644) <= b and not a;
    layer1_outputs(645) <= b;
    layer1_outputs(646) <= not b;
    layer1_outputs(647) <= a;
    layer1_outputs(648) <= not b;
    layer1_outputs(649) <= not b or a;
    layer1_outputs(650) <= '0';
    layer1_outputs(651) <= not (a xor b);
    layer1_outputs(652) <= not b or a;
    layer1_outputs(653) <= a;
    layer1_outputs(654) <= a or b;
    layer1_outputs(655) <= a or b;
    layer1_outputs(656) <= not a or b;
    layer1_outputs(657) <= a;
    layer1_outputs(658) <= not b;
    layer1_outputs(659) <= not (a xor b);
    layer1_outputs(660) <= a and b;
    layer1_outputs(661) <= not b or a;
    layer1_outputs(662) <= a and not b;
    layer1_outputs(663) <= a or b;
    layer1_outputs(664) <= '0';
    layer1_outputs(665) <= a xor b;
    layer1_outputs(666) <= b;
    layer1_outputs(667) <= not b or a;
    layer1_outputs(668) <= not a;
    layer1_outputs(669) <= b and not a;
    layer1_outputs(670) <= not a;
    layer1_outputs(671) <= b;
    layer1_outputs(672) <= not a or b;
    layer1_outputs(673) <= not b or a;
    layer1_outputs(674) <= a;
    layer1_outputs(675) <= not (a or b);
    layer1_outputs(676) <= a and b;
    layer1_outputs(677) <= not (a or b);
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= '1';
    layer1_outputs(680) <= b;
    layer1_outputs(681) <= b and not a;
    layer1_outputs(682) <= a;
    layer1_outputs(683) <= not (a and b);
    layer1_outputs(684) <= not b or a;
    layer1_outputs(685) <= not (a xor b);
    layer1_outputs(686) <= a and not b;
    layer1_outputs(687) <= b and not a;
    layer1_outputs(688) <= not (a xor b);
    layer1_outputs(689) <= not a or b;
    layer1_outputs(690) <= not b;
    layer1_outputs(691) <= a;
    layer1_outputs(692) <= b and not a;
    layer1_outputs(693) <= a;
    layer1_outputs(694) <= a and not b;
    layer1_outputs(695) <= b and not a;
    layer1_outputs(696) <= not b;
    layer1_outputs(697) <= not (a xor b);
    layer1_outputs(698) <= a and not b;
    layer1_outputs(699) <= a and not b;
    layer1_outputs(700) <= not (a and b);
    layer1_outputs(701) <= not a;
    layer1_outputs(702) <= b and not a;
    layer1_outputs(703) <= not b;
    layer1_outputs(704) <= '0';
    layer1_outputs(705) <= a;
    layer1_outputs(706) <= not (a or b);
    layer1_outputs(707) <= not b or a;
    layer1_outputs(708) <= not (a xor b);
    layer1_outputs(709) <= a or b;
    layer1_outputs(710) <= not (a or b);
    layer1_outputs(711) <= a xor b;
    layer1_outputs(712) <= b and not a;
    layer1_outputs(713) <= a and b;
    layer1_outputs(714) <= not (a xor b);
    layer1_outputs(715) <= a;
    layer1_outputs(716) <= b;
    layer1_outputs(717) <= b;
    layer1_outputs(718) <= not a or b;
    layer1_outputs(719) <= not b or a;
    layer1_outputs(720) <= not (a and b);
    layer1_outputs(721) <= not b;
    layer1_outputs(722) <= b;
    layer1_outputs(723) <= not (a or b);
    layer1_outputs(724) <= not (a xor b);
    layer1_outputs(725) <= not b or a;
    layer1_outputs(726) <= not b;
    layer1_outputs(727) <= a or b;
    layer1_outputs(728) <= '0';
    layer1_outputs(729) <= not a or b;
    layer1_outputs(730) <= not (a and b);
    layer1_outputs(731) <= not a;
    layer1_outputs(732) <= a;
    layer1_outputs(733) <= not (a or b);
    layer1_outputs(734) <= b;
    layer1_outputs(735) <= a and not b;
    layer1_outputs(736) <= a or b;
    layer1_outputs(737) <= b;
    layer1_outputs(738) <= not a;
    layer1_outputs(739) <= not b or a;
    layer1_outputs(740) <= not (a or b);
    layer1_outputs(741) <= not a;
    layer1_outputs(742) <= b;
    layer1_outputs(743) <= a and not b;
    layer1_outputs(744) <= b;
    layer1_outputs(745) <= b and not a;
    layer1_outputs(746) <= not (a xor b);
    layer1_outputs(747) <= not b;
    layer1_outputs(748) <= not (a or b);
    layer1_outputs(749) <= b and not a;
    layer1_outputs(750) <= a;
    layer1_outputs(751) <= not (a or b);
    layer1_outputs(752) <= not b;
    layer1_outputs(753) <= b and not a;
    layer1_outputs(754) <= not b;
    layer1_outputs(755) <= b;
    layer1_outputs(756) <= not b;
    layer1_outputs(757) <= not a;
    layer1_outputs(758) <= a xor b;
    layer1_outputs(759) <= a and b;
    layer1_outputs(760) <= not b;
    layer1_outputs(761) <= not (a xor b);
    layer1_outputs(762) <= not (a or b);
    layer1_outputs(763) <= b and not a;
    layer1_outputs(764) <= not (a or b);
    layer1_outputs(765) <= not (a xor b);
    layer1_outputs(766) <= b;
    layer1_outputs(767) <= not b;
    layer1_outputs(768) <= a;
    layer1_outputs(769) <= b;
    layer1_outputs(770) <= not a;
    layer1_outputs(771) <= not b or a;
    layer1_outputs(772) <= '0';
    layer1_outputs(773) <= a or b;
    layer1_outputs(774) <= not b or a;
    layer1_outputs(775) <= a or b;
    layer1_outputs(776) <= a;
    layer1_outputs(777) <= a and not b;
    layer1_outputs(778) <= not b;
    layer1_outputs(779) <= '0';
    layer1_outputs(780) <= a or b;
    layer1_outputs(781) <= a;
    layer1_outputs(782) <= not b or a;
    layer1_outputs(783) <= a or b;
    layer1_outputs(784) <= a and not b;
    layer1_outputs(785) <= b and not a;
    layer1_outputs(786) <= b;
    layer1_outputs(787) <= a;
    layer1_outputs(788) <= not (a or b);
    layer1_outputs(789) <= not b;
    layer1_outputs(790) <= not b;
    layer1_outputs(791) <= not a;
    layer1_outputs(792) <= b and not a;
    layer1_outputs(793) <= not a or b;
    layer1_outputs(794) <= a or b;
    layer1_outputs(795) <= a or b;
    layer1_outputs(796) <= a;
    layer1_outputs(797) <= b;
    layer1_outputs(798) <= not a or b;
    layer1_outputs(799) <= not (a and b);
    layer1_outputs(800) <= b and not a;
    layer1_outputs(801) <= b;
    layer1_outputs(802) <= not a or b;
    layer1_outputs(803) <= not (a or b);
    layer1_outputs(804) <= a or b;
    layer1_outputs(805) <= not b or a;
    layer1_outputs(806) <= b;
    layer1_outputs(807) <= not (a xor b);
    layer1_outputs(808) <= not b or a;
    layer1_outputs(809) <= a or b;
    layer1_outputs(810) <= not a or b;
    layer1_outputs(811) <= not b or a;
    layer1_outputs(812) <= '0';
    layer1_outputs(813) <= b and not a;
    layer1_outputs(814) <= b;
    layer1_outputs(815) <= not (a xor b);
    layer1_outputs(816) <= '1';
    layer1_outputs(817) <= b;
    layer1_outputs(818) <= not b;
    layer1_outputs(819) <= not a or b;
    layer1_outputs(820) <= b and not a;
    layer1_outputs(821) <= a;
    layer1_outputs(822) <= b;
    layer1_outputs(823) <= a and not b;
    layer1_outputs(824) <= not a or b;
    layer1_outputs(825) <= a xor b;
    layer1_outputs(826) <= a and not b;
    layer1_outputs(827) <= b;
    layer1_outputs(828) <= a;
    layer1_outputs(829) <= not (a and b);
    layer1_outputs(830) <= a and not b;
    layer1_outputs(831) <= '1';
    layer1_outputs(832) <= a or b;
    layer1_outputs(833) <= a;
    layer1_outputs(834) <= not (a or b);
    layer1_outputs(835) <= not a or b;
    layer1_outputs(836) <= a xor b;
    layer1_outputs(837) <= not b or a;
    layer1_outputs(838) <= not b or a;
    layer1_outputs(839) <= not a;
    layer1_outputs(840) <= not b or a;
    layer1_outputs(841) <= not (a and b);
    layer1_outputs(842) <= b;
    layer1_outputs(843) <= not b or a;
    layer1_outputs(844) <= not (a and b);
    layer1_outputs(845) <= '1';
    layer1_outputs(846) <= a xor b;
    layer1_outputs(847) <= not a;
    layer1_outputs(848) <= b;
    layer1_outputs(849) <= a and not b;
    layer1_outputs(850) <= '1';
    layer1_outputs(851) <= a and b;
    layer1_outputs(852) <= not a or b;
    layer1_outputs(853) <= not a or b;
    layer1_outputs(854) <= b;
    layer1_outputs(855) <= b;
    layer1_outputs(856) <= a and b;
    layer1_outputs(857) <= a and b;
    layer1_outputs(858) <= not a;
    layer1_outputs(859) <= not a;
    layer1_outputs(860) <= not a;
    layer1_outputs(861) <= not (a and b);
    layer1_outputs(862) <= a;
    layer1_outputs(863) <= not a;
    layer1_outputs(864) <= not a;
    layer1_outputs(865) <= a or b;
    layer1_outputs(866) <= not a or b;
    layer1_outputs(867) <= a xor b;
    layer1_outputs(868) <= not a or b;
    layer1_outputs(869) <= b;
    layer1_outputs(870) <= not (a xor b);
    layer1_outputs(871) <= not (a or b);
    layer1_outputs(872) <= a;
    layer1_outputs(873) <= not (a or b);
    layer1_outputs(874) <= not (a xor b);
    layer1_outputs(875) <= not (a or b);
    layer1_outputs(876) <= a and b;
    layer1_outputs(877) <= '1';
    layer1_outputs(878) <= a or b;
    layer1_outputs(879) <= a and not b;
    layer1_outputs(880) <= a and not b;
    layer1_outputs(881) <= b;
    layer1_outputs(882) <= a or b;
    layer1_outputs(883) <= a or b;
    layer1_outputs(884) <= a xor b;
    layer1_outputs(885) <= a or b;
    layer1_outputs(886) <= a or b;
    layer1_outputs(887) <= not a;
    layer1_outputs(888) <= not (a or b);
    layer1_outputs(889) <= '1';
    layer1_outputs(890) <= not (a or b);
    layer1_outputs(891) <= a;
    layer1_outputs(892) <= '1';
    layer1_outputs(893) <= not b or a;
    layer1_outputs(894) <= not a or b;
    layer1_outputs(895) <= a or b;
    layer1_outputs(896) <= not b or a;
    layer1_outputs(897) <= a;
    layer1_outputs(898) <= a or b;
    layer1_outputs(899) <= '1';
    layer1_outputs(900) <= a;
    layer1_outputs(901) <= a or b;
    layer1_outputs(902) <= not b or a;
    layer1_outputs(903) <= not a;
    layer1_outputs(904) <= a or b;
    layer1_outputs(905) <= not b or a;
    layer1_outputs(906) <= b and not a;
    layer1_outputs(907) <= not (a and b);
    layer1_outputs(908) <= not a;
    layer1_outputs(909) <= a;
    layer1_outputs(910) <= not b;
    layer1_outputs(911) <= not (a and b);
    layer1_outputs(912) <= b and not a;
    layer1_outputs(913) <= not (a or b);
    layer1_outputs(914) <= a;
    layer1_outputs(915) <= not b or a;
    layer1_outputs(916) <= not b;
    layer1_outputs(917) <= b;
    layer1_outputs(918) <= a and b;
    layer1_outputs(919) <= not (a or b);
    layer1_outputs(920) <= not b or a;
    layer1_outputs(921) <= not (a and b);
    layer1_outputs(922) <= a and b;
    layer1_outputs(923) <= not (a xor b);
    layer1_outputs(924) <= not a;
    layer1_outputs(925) <= not b;
    layer1_outputs(926) <= not (a and b);
    layer1_outputs(927) <= '0';
    layer1_outputs(928) <= not (a or b);
    layer1_outputs(929) <= a and b;
    layer1_outputs(930) <= not a;
    layer1_outputs(931) <= not a;
    layer1_outputs(932) <= not a;
    layer1_outputs(933) <= a xor b;
    layer1_outputs(934) <= a or b;
    layer1_outputs(935) <= not a or b;
    layer1_outputs(936) <= a;
    layer1_outputs(937) <= a and not b;
    layer1_outputs(938) <= b and not a;
    layer1_outputs(939) <= a or b;
    layer1_outputs(940) <= not (a or b);
    layer1_outputs(941) <= b;
    layer1_outputs(942) <= not (a and b);
    layer1_outputs(943) <= b and not a;
    layer1_outputs(944) <= not a;
    layer1_outputs(945) <= a or b;
    layer1_outputs(946) <= not b;
    layer1_outputs(947) <= a and not b;
    layer1_outputs(948) <= a xor b;
    layer1_outputs(949) <= a;
    layer1_outputs(950) <= not b;
    layer1_outputs(951) <= not (a and b);
    layer1_outputs(952) <= not b;
    layer1_outputs(953) <= not (a or b);
    layer1_outputs(954) <= b;
    layer1_outputs(955) <= not b;
    layer1_outputs(956) <= not (a and b);
    layer1_outputs(957) <= not a;
    layer1_outputs(958) <= a or b;
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= not a or b;
    layer1_outputs(961) <= not (a and b);
    layer1_outputs(962) <= not a or b;
    layer1_outputs(963) <= a or b;
    layer1_outputs(964) <= not (a and b);
    layer1_outputs(965) <= b;
    layer1_outputs(966) <= not a or b;
    layer1_outputs(967) <= b;
    layer1_outputs(968) <= not b;
    layer1_outputs(969) <= not a or b;
    layer1_outputs(970) <= not a;
    layer1_outputs(971) <= not b or a;
    layer1_outputs(972) <= not (a and b);
    layer1_outputs(973) <= a and b;
    layer1_outputs(974) <= a xor b;
    layer1_outputs(975) <= b and not a;
    layer1_outputs(976) <= not b;
    layer1_outputs(977) <= not a;
    layer1_outputs(978) <= a xor b;
    layer1_outputs(979) <= not a;
    layer1_outputs(980) <= not b or a;
    layer1_outputs(981) <= not a or b;
    layer1_outputs(982) <= a or b;
    layer1_outputs(983) <= b and not a;
    layer1_outputs(984) <= not a or b;
    layer1_outputs(985) <= not (a and b);
    layer1_outputs(986) <= b;
    layer1_outputs(987) <= not a or b;
    layer1_outputs(988) <= '1';
    layer1_outputs(989) <= not (a and b);
    layer1_outputs(990) <= not a or b;
    layer1_outputs(991) <= a xor b;
    layer1_outputs(992) <= b;
    layer1_outputs(993) <= not b or a;
    layer1_outputs(994) <= a and not b;
    layer1_outputs(995) <= a;
    layer1_outputs(996) <= not b or a;
    layer1_outputs(997) <= not (a and b);
    layer1_outputs(998) <= '1';
    layer1_outputs(999) <= not a;
    layer1_outputs(1000) <= not b or a;
    layer1_outputs(1001) <= a or b;
    layer1_outputs(1002) <= not (a and b);
    layer1_outputs(1003) <= not (a and b);
    layer1_outputs(1004) <= a or b;
    layer1_outputs(1005) <= a;
    layer1_outputs(1006) <= not b or a;
    layer1_outputs(1007) <= a or b;
    layer1_outputs(1008) <= not b;
    layer1_outputs(1009) <= not (a xor b);
    layer1_outputs(1010) <= b;
    layer1_outputs(1011) <= not (a or b);
    layer1_outputs(1012) <= b and not a;
    layer1_outputs(1013) <= not b;
    layer1_outputs(1014) <= b and not a;
    layer1_outputs(1015) <= not (a or b);
    layer1_outputs(1016) <= not b;
    layer1_outputs(1017) <= not b;
    layer1_outputs(1018) <= b and not a;
    layer1_outputs(1019) <= not a or b;
    layer1_outputs(1020) <= a xor b;
    layer1_outputs(1021) <= not b;
    layer1_outputs(1022) <= a and b;
    layer1_outputs(1023) <= b;
    layer1_outputs(1024) <= a xor b;
    layer1_outputs(1025) <= b;
    layer1_outputs(1026) <= not (a xor b);
    layer1_outputs(1027) <= not (a or b);
    layer1_outputs(1028) <= not a;
    layer1_outputs(1029) <= not a;
    layer1_outputs(1030) <= not a;
    layer1_outputs(1031) <= not a or b;
    layer1_outputs(1032) <= not a;
    layer1_outputs(1033) <= a or b;
    layer1_outputs(1034) <= not (a and b);
    layer1_outputs(1035) <= b;
    layer1_outputs(1036) <= b;
    layer1_outputs(1037) <= not a;
    layer1_outputs(1038) <= not b;
    layer1_outputs(1039) <= not (a or b);
    layer1_outputs(1040) <= not (a or b);
    layer1_outputs(1041) <= not a or b;
    layer1_outputs(1042) <= '1';
    layer1_outputs(1043) <= not a;
    layer1_outputs(1044) <= not a;
    layer1_outputs(1045) <= not a;
    layer1_outputs(1046) <= not (a and b);
    layer1_outputs(1047) <= a;
    layer1_outputs(1048) <= a;
    layer1_outputs(1049) <= not b;
    layer1_outputs(1050) <= not b or a;
    layer1_outputs(1051) <= not b or a;
    layer1_outputs(1052) <= b and not a;
    layer1_outputs(1053) <= a or b;
    layer1_outputs(1054) <= a or b;
    layer1_outputs(1055) <= not a or b;
    layer1_outputs(1056) <= b and not a;
    layer1_outputs(1057) <= b;
    layer1_outputs(1058) <= not (a or b);
    layer1_outputs(1059) <= '0';
    layer1_outputs(1060) <= not b;
    layer1_outputs(1061) <= a;
    layer1_outputs(1062) <= '0';
    layer1_outputs(1063) <= not (a and b);
    layer1_outputs(1064) <= a and b;
    layer1_outputs(1065) <= b;
    layer1_outputs(1066) <= not a or b;
    layer1_outputs(1067) <= a or b;
    layer1_outputs(1068) <= a or b;
    layer1_outputs(1069) <= not a or b;
    layer1_outputs(1070) <= not b or a;
    layer1_outputs(1071) <= not (a or b);
    layer1_outputs(1072) <= a and b;
    layer1_outputs(1073) <= not b or a;
    layer1_outputs(1074) <= a xor b;
    layer1_outputs(1075) <= not a;
    layer1_outputs(1076) <= a and b;
    layer1_outputs(1077) <= b;
    layer1_outputs(1078) <= a and b;
    layer1_outputs(1079) <= a and b;
    layer1_outputs(1080) <= a xor b;
    layer1_outputs(1081) <= a;
    layer1_outputs(1082) <= not a;
    layer1_outputs(1083) <= b;
    layer1_outputs(1084) <= not a or b;
    layer1_outputs(1085) <= not a or b;
    layer1_outputs(1086) <= not b;
    layer1_outputs(1087) <= not b;
    layer1_outputs(1088) <= '1';
    layer1_outputs(1089) <= not (a xor b);
    layer1_outputs(1090) <= not a;
    layer1_outputs(1091) <= b;
    layer1_outputs(1092) <= a or b;
    layer1_outputs(1093) <= a;
    layer1_outputs(1094) <= not b or a;
    layer1_outputs(1095) <= not a;
    layer1_outputs(1096) <= '1';
    layer1_outputs(1097) <= a and not b;
    layer1_outputs(1098) <= not (a and b);
    layer1_outputs(1099) <= b;
    layer1_outputs(1100) <= b and not a;
    layer1_outputs(1101) <= a or b;
    layer1_outputs(1102) <= not (a or b);
    layer1_outputs(1103) <= not b or a;
    layer1_outputs(1104) <= a and b;
    layer1_outputs(1105) <= not a;
    layer1_outputs(1106) <= not (a and b);
    layer1_outputs(1107) <= b;
    layer1_outputs(1108) <= a;
    layer1_outputs(1109) <= b and not a;
    layer1_outputs(1110) <= a and not b;
    layer1_outputs(1111) <= '1';
    layer1_outputs(1112) <= not (a xor b);
    layer1_outputs(1113) <= a xor b;
    layer1_outputs(1114) <= a and b;
    layer1_outputs(1115) <= a and not b;
    layer1_outputs(1116) <= '0';
    layer1_outputs(1117) <= not (a and b);
    layer1_outputs(1118) <= not a or b;
    layer1_outputs(1119) <= a and b;
    layer1_outputs(1120) <= a and not b;
    layer1_outputs(1121) <= a;
    layer1_outputs(1122) <= not (a and b);
    layer1_outputs(1123) <= b and not a;
    layer1_outputs(1124) <= a;
    layer1_outputs(1125) <= b;
    layer1_outputs(1126) <= b;
    layer1_outputs(1127) <= b and not a;
    layer1_outputs(1128) <= a xor b;
    layer1_outputs(1129) <= not (a and b);
    layer1_outputs(1130) <= a and not b;
    layer1_outputs(1131) <= not b or a;
    layer1_outputs(1132) <= a xor b;
    layer1_outputs(1133) <= not b or a;
    layer1_outputs(1134) <= a or b;
    layer1_outputs(1135) <= a and b;
    layer1_outputs(1136) <= a;
    layer1_outputs(1137) <= not (a or b);
    layer1_outputs(1138) <= not a or b;
    layer1_outputs(1139) <= b and not a;
    layer1_outputs(1140) <= a;
    layer1_outputs(1141) <= a or b;
    layer1_outputs(1142) <= '0';
    layer1_outputs(1143) <= a;
    layer1_outputs(1144) <= not (a and b);
    layer1_outputs(1145) <= not a;
    layer1_outputs(1146) <= not (a and b);
    layer1_outputs(1147) <= a and b;
    layer1_outputs(1148) <= not b;
    layer1_outputs(1149) <= not b;
    layer1_outputs(1150) <= not b or a;
    layer1_outputs(1151) <= a and not b;
    layer1_outputs(1152) <= not (a and b);
    layer1_outputs(1153) <= b and not a;
    layer1_outputs(1154) <= b;
    layer1_outputs(1155) <= a xor b;
    layer1_outputs(1156) <= not b or a;
    layer1_outputs(1157) <= a and b;
    layer1_outputs(1158) <= b and not a;
    layer1_outputs(1159) <= not b;
    layer1_outputs(1160) <= not b or a;
    layer1_outputs(1161) <= a xor b;
    layer1_outputs(1162) <= not a or b;
    layer1_outputs(1163) <= b and not a;
    layer1_outputs(1164) <= a and b;
    layer1_outputs(1165) <= b and not a;
    layer1_outputs(1166) <= b;
    layer1_outputs(1167) <= not a;
    layer1_outputs(1168) <= not (a and b);
    layer1_outputs(1169) <= not a;
    layer1_outputs(1170) <= '1';
    layer1_outputs(1171) <= not a;
    layer1_outputs(1172) <= b;
    layer1_outputs(1173) <= not (a and b);
    layer1_outputs(1174) <= b and not a;
    layer1_outputs(1175) <= a or b;
    layer1_outputs(1176) <= not a or b;
    layer1_outputs(1177) <= a and not b;
    layer1_outputs(1178) <= a xor b;
    layer1_outputs(1179) <= a or b;
    layer1_outputs(1180) <= not b or a;
    layer1_outputs(1181) <= not b or a;
    layer1_outputs(1182) <= not (a or b);
    layer1_outputs(1183) <= not b or a;
    layer1_outputs(1184) <= a and not b;
    layer1_outputs(1185) <= '0';
    layer1_outputs(1186) <= not (a and b);
    layer1_outputs(1187) <= not (a and b);
    layer1_outputs(1188) <= a and not b;
    layer1_outputs(1189) <= b;
    layer1_outputs(1190) <= not a or b;
    layer1_outputs(1191) <= '1';
    layer1_outputs(1192) <= not (a and b);
    layer1_outputs(1193) <= not (a and b);
    layer1_outputs(1194) <= b;
    layer1_outputs(1195) <= '0';
    layer1_outputs(1196) <= not a;
    layer1_outputs(1197) <= not (a and b);
    layer1_outputs(1198) <= a;
    layer1_outputs(1199) <= a xor b;
    layer1_outputs(1200) <= not b;
    layer1_outputs(1201) <= not b or a;
    layer1_outputs(1202) <= not (a or b);
    layer1_outputs(1203) <= not b or a;
    layer1_outputs(1204) <= b;
    layer1_outputs(1205) <= a or b;
    layer1_outputs(1206) <= not b;
    layer1_outputs(1207) <= a xor b;
    layer1_outputs(1208) <= not a or b;
    layer1_outputs(1209) <= not b or a;
    layer1_outputs(1210) <= a;
    layer1_outputs(1211) <= not b or a;
    layer1_outputs(1212) <= not b or a;
    layer1_outputs(1213) <= a;
    layer1_outputs(1214) <= not a;
    layer1_outputs(1215) <= '0';
    layer1_outputs(1216) <= not a;
    layer1_outputs(1217) <= a and not b;
    layer1_outputs(1218) <= a or b;
    layer1_outputs(1219) <= a;
    layer1_outputs(1220) <= a;
    layer1_outputs(1221) <= '1';
    layer1_outputs(1222) <= not a;
    layer1_outputs(1223) <= not (a and b);
    layer1_outputs(1224) <= b and not a;
    layer1_outputs(1225) <= not (a and b);
    layer1_outputs(1226) <= not b or a;
    layer1_outputs(1227) <= a;
    layer1_outputs(1228) <= not (a xor b);
    layer1_outputs(1229) <= not a;
    layer1_outputs(1230) <= b;
    layer1_outputs(1231) <= not (a and b);
    layer1_outputs(1232) <= b;
    layer1_outputs(1233) <= a and not b;
    layer1_outputs(1234) <= not (a or b);
    layer1_outputs(1235) <= a and not b;
    layer1_outputs(1236) <= a or b;
    layer1_outputs(1237) <= a and b;
    layer1_outputs(1238) <= not b;
    layer1_outputs(1239) <= not b;
    layer1_outputs(1240) <= a and b;
    layer1_outputs(1241) <= not b;
    layer1_outputs(1242) <= b and not a;
    layer1_outputs(1243) <= not (a and b);
    layer1_outputs(1244) <= not (a or b);
    layer1_outputs(1245) <= not (a or b);
    layer1_outputs(1246) <= a;
    layer1_outputs(1247) <= not a or b;
    layer1_outputs(1248) <= a or b;
    layer1_outputs(1249) <= a and b;
    layer1_outputs(1250) <= not b;
    layer1_outputs(1251) <= '1';
    layer1_outputs(1252) <= not b or a;
    layer1_outputs(1253) <= a or b;
    layer1_outputs(1254) <= not a;
    layer1_outputs(1255) <= b;
    layer1_outputs(1256) <= not a;
    layer1_outputs(1257) <= b;
    layer1_outputs(1258) <= a and b;
    layer1_outputs(1259) <= a xor b;
    layer1_outputs(1260) <= not b or a;
    layer1_outputs(1261) <= not a;
    layer1_outputs(1262) <= a;
    layer1_outputs(1263) <= a or b;
    layer1_outputs(1264) <= not b;
    layer1_outputs(1265) <= not (a and b);
    layer1_outputs(1266) <= b;
    layer1_outputs(1267) <= b and not a;
    layer1_outputs(1268) <= a and not b;
    layer1_outputs(1269) <= not (a or b);
    layer1_outputs(1270) <= not b or a;
    layer1_outputs(1271) <= b;
    layer1_outputs(1272) <= not (a or b);
    layer1_outputs(1273) <= not a;
    layer1_outputs(1274) <= a xor b;
    layer1_outputs(1275) <= b;
    layer1_outputs(1276) <= a;
    layer1_outputs(1277) <= b and not a;
    layer1_outputs(1278) <= not (a and b);
    layer1_outputs(1279) <= not (a or b);
    layer1_outputs(1280) <= not b or a;
    layer1_outputs(1281) <= not a or b;
    layer1_outputs(1282) <= a and not b;
    layer1_outputs(1283) <= b and not a;
    layer1_outputs(1284) <= not a;
    layer1_outputs(1285) <= a;
    layer1_outputs(1286) <= a;
    layer1_outputs(1287) <= not b;
    layer1_outputs(1288) <= not b or a;
    layer1_outputs(1289) <= not (a or b);
    layer1_outputs(1290) <= b and not a;
    layer1_outputs(1291) <= a and not b;
    layer1_outputs(1292) <= a xor b;
    layer1_outputs(1293) <= a and b;
    layer1_outputs(1294) <= not (a or b);
    layer1_outputs(1295) <= b;
    layer1_outputs(1296) <= not b or a;
    layer1_outputs(1297) <= not b or a;
    layer1_outputs(1298) <= b and not a;
    layer1_outputs(1299) <= '0';
    layer1_outputs(1300) <= a or b;
    layer1_outputs(1301) <= '0';
    layer1_outputs(1302) <= not b;
    layer1_outputs(1303) <= not (a and b);
    layer1_outputs(1304) <= not a;
    layer1_outputs(1305) <= not (a or b);
    layer1_outputs(1306) <= '1';
    layer1_outputs(1307) <= a;
    layer1_outputs(1308) <= not (a and b);
    layer1_outputs(1309) <= not b;
    layer1_outputs(1310) <= '1';
    layer1_outputs(1311) <= a xor b;
    layer1_outputs(1312) <= not b;
    layer1_outputs(1313) <= b;
    layer1_outputs(1314) <= a and not b;
    layer1_outputs(1315) <= a and not b;
    layer1_outputs(1316) <= b and not a;
    layer1_outputs(1317) <= not (a and b);
    layer1_outputs(1318) <= not a;
    layer1_outputs(1319) <= a and b;
    layer1_outputs(1320) <= not b;
    layer1_outputs(1321) <= a;
    layer1_outputs(1322) <= not b or a;
    layer1_outputs(1323) <= not a or b;
    layer1_outputs(1324) <= not a;
    layer1_outputs(1325) <= '0';
    layer1_outputs(1326) <= a;
    layer1_outputs(1327) <= not a or b;
    layer1_outputs(1328) <= not (a or b);
    layer1_outputs(1329) <= '1';
    layer1_outputs(1330) <= '0';
    layer1_outputs(1331) <= not a;
    layer1_outputs(1332) <= a xor b;
    layer1_outputs(1333) <= not a;
    layer1_outputs(1334) <= not (a xor b);
    layer1_outputs(1335) <= not a or b;
    layer1_outputs(1336) <= not a;
    layer1_outputs(1337) <= a and b;
    layer1_outputs(1338) <= '1';
    layer1_outputs(1339) <= a and b;
    layer1_outputs(1340) <= '1';
    layer1_outputs(1341) <= not b;
    layer1_outputs(1342) <= not (a and b);
    layer1_outputs(1343) <= not (a or b);
    layer1_outputs(1344) <= not b;
    layer1_outputs(1345) <= not b;
    layer1_outputs(1346) <= b;
    layer1_outputs(1347) <= '1';
    layer1_outputs(1348) <= not (a xor b);
    layer1_outputs(1349) <= a and not b;
    layer1_outputs(1350) <= not a or b;
    layer1_outputs(1351) <= '0';
    layer1_outputs(1352) <= a or b;
    layer1_outputs(1353) <= not a or b;
    layer1_outputs(1354) <= b and not a;
    layer1_outputs(1355) <= a xor b;
    layer1_outputs(1356) <= a;
    layer1_outputs(1357) <= not a or b;
    layer1_outputs(1358) <= not b;
    layer1_outputs(1359) <= not b;
    layer1_outputs(1360) <= not (a and b);
    layer1_outputs(1361) <= not (a or b);
    layer1_outputs(1362) <= '1';
    layer1_outputs(1363) <= not b;
    layer1_outputs(1364) <= not b;
    layer1_outputs(1365) <= not (a xor b);
    layer1_outputs(1366) <= not (a and b);
    layer1_outputs(1367) <= not a;
    layer1_outputs(1368) <= a;
    layer1_outputs(1369) <= not a;
    layer1_outputs(1370) <= not a;
    layer1_outputs(1371) <= a or b;
    layer1_outputs(1372) <= b;
    layer1_outputs(1373) <= not b;
    layer1_outputs(1374) <= not (a and b);
    layer1_outputs(1375) <= not a or b;
    layer1_outputs(1376) <= not (a and b);
    layer1_outputs(1377) <= not b or a;
    layer1_outputs(1378) <= a and not b;
    layer1_outputs(1379) <= a xor b;
    layer1_outputs(1380) <= a xor b;
    layer1_outputs(1381) <= not a or b;
    layer1_outputs(1382) <= b and not a;
    layer1_outputs(1383) <= a;
    layer1_outputs(1384) <= b;
    layer1_outputs(1385) <= b;
    layer1_outputs(1386) <= b and not a;
    layer1_outputs(1387) <= a and not b;
    layer1_outputs(1388) <= '1';
    layer1_outputs(1389) <= not b;
    layer1_outputs(1390) <= a and b;
    layer1_outputs(1391) <= not a;
    layer1_outputs(1392) <= a;
    layer1_outputs(1393) <= b;
    layer1_outputs(1394) <= a or b;
    layer1_outputs(1395) <= b;
    layer1_outputs(1396) <= not (a or b);
    layer1_outputs(1397) <= a and b;
    layer1_outputs(1398) <= b;
    layer1_outputs(1399) <= not (a xor b);
    layer1_outputs(1400) <= b and not a;
    layer1_outputs(1401) <= not (a xor b);
    layer1_outputs(1402) <= not a;
    layer1_outputs(1403) <= '1';
    layer1_outputs(1404) <= not b or a;
    layer1_outputs(1405) <= a or b;
    layer1_outputs(1406) <= b;
    layer1_outputs(1407) <= a and not b;
    layer1_outputs(1408) <= not (a xor b);
    layer1_outputs(1409) <= a and not b;
    layer1_outputs(1410) <= not b;
    layer1_outputs(1411) <= not b or a;
    layer1_outputs(1412) <= not (a or b);
    layer1_outputs(1413) <= not a or b;
    layer1_outputs(1414) <= not b or a;
    layer1_outputs(1415) <= not (a or b);
    layer1_outputs(1416) <= not (a or b);
    layer1_outputs(1417) <= a xor b;
    layer1_outputs(1418) <= not b;
    layer1_outputs(1419) <= not a or b;
    layer1_outputs(1420) <= not (a or b);
    layer1_outputs(1421) <= a and not b;
    layer1_outputs(1422) <= a;
    layer1_outputs(1423) <= not (a and b);
    layer1_outputs(1424) <= not a or b;
    layer1_outputs(1425) <= a;
    layer1_outputs(1426) <= not (a and b);
    layer1_outputs(1427) <= b and not a;
    layer1_outputs(1428) <= '1';
    layer1_outputs(1429) <= a and not b;
    layer1_outputs(1430) <= a and not b;
    layer1_outputs(1431) <= not b;
    layer1_outputs(1432) <= a or b;
    layer1_outputs(1433) <= not (a or b);
    layer1_outputs(1434) <= not a;
    layer1_outputs(1435) <= '0';
    layer1_outputs(1436) <= a or b;
    layer1_outputs(1437) <= b and not a;
    layer1_outputs(1438) <= not (a and b);
    layer1_outputs(1439) <= not b;
    layer1_outputs(1440) <= a;
    layer1_outputs(1441) <= not a or b;
    layer1_outputs(1442) <= not (a xor b);
    layer1_outputs(1443) <= b and not a;
    layer1_outputs(1444) <= not b;
    layer1_outputs(1445) <= not b;
    layer1_outputs(1446) <= b and not a;
    layer1_outputs(1447) <= not (a and b);
    layer1_outputs(1448) <= not a;
    layer1_outputs(1449) <= not b;
    layer1_outputs(1450) <= a and not b;
    layer1_outputs(1451) <= a and b;
    layer1_outputs(1452) <= a and not b;
    layer1_outputs(1453) <= not a;
    layer1_outputs(1454) <= a;
    layer1_outputs(1455) <= not a or b;
    layer1_outputs(1456) <= not (a xor b);
    layer1_outputs(1457) <= not b or a;
    layer1_outputs(1458) <= a;
    layer1_outputs(1459) <= not a or b;
    layer1_outputs(1460) <= not a or b;
    layer1_outputs(1461) <= a and b;
    layer1_outputs(1462) <= a or b;
    layer1_outputs(1463) <= a and not b;
    layer1_outputs(1464) <= '1';
    layer1_outputs(1465) <= '0';
    layer1_outputs(1466) <= not b or a;
    layer1_outputs(1467) <= b and not a;
    layer1_outputs(1468) <= a and b;
    layer1_outputs(1469) <= '0';
    layer1_outputs(1470) <= not (a or b);
    layer1_outputs(1471) <= a xor b;
    layer1_outputs(1472) <= b;
    layer1_outputs(1473) <= not a;
    layer1_outputs(1474) <= a or b;
    layer1_outputs(1475) <= '0';
    layer1_outputs(1476) <= b and not a;
    layer1_outputs(1477) <= '0';
    layer1_outputs(1478) <= a or b;
    layer1_outputs(1479) <= '1';
    layer1_outputs(1480) <= '1';
    layer1_outputs(1481) <= a xor b;
    layer1_outputs(1482) <= not a;
    layer1_outputs(1483) <= not (a and b);
    layer1_outputs(1484) <= b;
    layer1_outputs(1485) <= b;
    layer1_outputs(1486) <= a or b;
    layer1_outputs(1487) <= not a;
    layer1_outputs(1488) <= a;
    layer1_outputs(1489) <= not a;
    layer1_outputs(1490) <= not a;
    layer1_outputs(1491) <= not a or b;
    layer1_outputs(1492) <= a;
    layer1_outputs(1493) <= a xor b;
    layer1_outputs(1494) <= not a;
    layer1_outputs(1495) <= not a or b;
    layer1_outputs(1496) <= not (a xor b);
    layer1_outputs(1497) <= '1';
    layer1_outputs(1498) <= not (a and b);
    layer1_outputs(1499) <= not a;
    layer1_outputs(1500) <= not a;
    layer1_outputs(1501) <= a and b;
    layer1_outputs(1502) <= not b;
    layer1_outputs(1503) <= not b;
    layer1_outputs(1504) <= not a;
    layer1_outputs(1505) <= '1';
    layer1_outputs(1506) <= '1';
    layer1_outputs(1507) <= a and not b;
    layer1_outputs(1508) <= b;
    layer1_outputs(1509) <= not a or b;
    layer1_outputs(1510) <= a and not b;
    layer1_outputs(1511) <= a and b;
    layer1_outputs(1512) <= not a;
    layer1_outputs(1513) <= not a or b;
    layer1_outputs(1514) <= not a;
    layer1_outputs(1515) <= not a;
    layer1_outputs(1516) <= a xor b;
    layer1_outputs(1517) <= not (a xor b);
    layer1_outputs(1518) <= a;
    layer1_outputs(1519) <= not (a or b);
    layer1_outputs(1520) <= not a or b;
    layer1_outputs(1521) <= a or b;
    layer1_outputs(1522) <= b and not a;
    layer1_outputs(1523) <= not (a xor b);
    layer1_outputs(1524) <= a xor b;
    layer1_outputs(1525) <= not b or a;
    layer1_outputs(1526) <= not a or b;
    layer1_outputs(1527) <= a and b;
    layer1_outputs(1528) <= a;
    layer1_outputs(1529) <= b and not a;
    layer1_outputs(1530) <= a;
    layer1_outputs(1531) <= not (a or b);
    layer1_outputs(1532) <= b and not a;
    layer1_outputs(1533) <= not (a or b);
    layer1_outputs(1534) <= not a or b;
    layer1_outputs(1535) <= not b or a;
    layer1_outputs(1536) <= not a;
    layer1_outputs(1537) <= a or b;
    layer1_outputs(1538) <= a;
    layer1_outputs(1539) <= b;
    layer1_outputs(1540) <= b and not a;
    layer1_outputs(1541) <= not (a xor b);
    layer1_outputs(1542) <= not (a and b);
    layer1_outputs(1543) <= not (a and b);
    layer1_outputs(1544) <= not b;
    layer1_outputs(1545) <= b;
    layer1_outputs(1546) <= not a;
    layer1_outputs(1547) <= not b;
    layer1_outputs(1548) <= not (a or b);
    layer1_outputs(1549) <= a or b;
    layer1_outputs(1550) <= b and not a;
    layer1_outputs(1551) <= b and not a;
    layer1_outputs(1552) <= a xor b;
    layer1_outputs(1553) <= not b;
    layer1_outputs(1554) <= not (a xor b);
    layer1_outputs(1555) <= '0';
    layer1_outputs(1556) <= a xor b;
    layer1_outputs(1557) <= not a;
    layer1_outputs(1558) <= not (a xor b);
    layer1_outputs(1559) <= b;
    layer1_outputs(1560) <= not b or a;
    layer1_outputs(1561) <= a and b;
    layer1_outputs(1562) <= a or b;
    layer1_outputs(1563) <= a or b;
    layer1_outputs(1564) <= a and not b;
    layer1_outputs(1565) <= not b or a;
    layer1_outputs(1566) <= not a;
    layer1_outputs(1567) <= a and not b;
    layer1_outputs(1568) <= b;
    layer1_outputs(1569) <= '0';
    layer1_outputs(1570) <= not b;
    layer1_outputs(1571) <= a or b;
    layer1_outputs(1572) <= a and b;
    layer1_outputs(1573) <= not b;
    layer1_outputs(1574) <= not (a or b);
    layer1_outputs(1575) <= a;
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= b;
    layer1_outputs(1578) <= a or b;
    layer1_outputs(1579) <= not (a and b);
    layer1_outputs(1580) <= not a or b;
    layer1_outputs(1581) <= a or b;
    layer1_outputs(1582) <= a and not b;
    layer1_outputs(1583) <= not b or a;
    layer1_outputs(1584) <= b and not a;
    layer1_outputs(1585) <= b and not a;
    layer1_outputs(1586) <= not a or b;
    layer1_outputs(1587) <= not (a or b);
    layer1_outputs(1588) <= '1';
    layer1_outputs(1589) <= a and b;
    layer1_outputs(1590) <= not (a and b);
    layer1_outputs(1591) <= not b or a;
    layer1_outputs(1592) <= not b;
    layer1_outputs(1593) <= not (a and b);
    layer1_outputs(1594) <= a and not b;
    layer1_outputs(1595) <= b and not a;
    layer1_outputs(1596) <= a and not b;
    layer1_outputs(1597) <= a and not b;
    layer1_outputs(1598) <= a;
    layer1_outputs(1599) <= a xor b;
    layer1_outputs(1600) <= '0';
    layer1_outputs(1601) <= a;
    layer1_outputs(1602) <= not a;
    layer1_outputs(1603) <= not b or a;
    layer1_outputs(1604) <= b;
    layer1_outputs(1605) <= a and not b;
    layer1_outputs(1606) <= not a;
    layer1_outputs(1607) <= a xor b;
    layer1_outputs(1608) <= a and not b;
    layer1_outputs(1609) <= a xor b;
    layer1_outputs(1610) <= not a or b;
    layer1_outputs(1611) <= a or b;
    layer1_outputs(1612) <= a or b;
    layer1_outputs(1613) <= a and b;
    layer1_outputs(1614) <= a and not b;
    layer1_outputs(1615) <= not b;
    layer1_outputs(1616) <= not b or a;
    layer1_outputs(1617) <= not a;
    layer1_outputs(1618) <= not (a xor b);
    layer1_outputs(1619) <= a;
    layer1_outputs(1620) <= not (a or b);
    layer1_outputs(1621) <= not b or a;
    layer1_outputs(1622) <= b and not a;
    layer1_outputs(1623) <= b and not a;
    layer1_outputs(1624) <= a and not b;
    layer1_outputs(1625) <= a or b;
    layer1_outputs(1626) <= a;
    layer1_outputs(1627) <= not a;
    layer1_outputs(1628) <= a xor b;
    layer1_outputs(1629) <= a or b;
    layer1_outputs(1630) <= b and not a;
    layer1_outputs(1631) <= not a;
    layer1_outputs(1632) <= not b or a;
    layer1_outputs(1633) <= not (a and b);
    layer1_outputs(1634) <= not (a xor b);
    layer1_outputs(1635) <= not (a or b);
    layer1_outputs(1636) <= a and b;
    layer1_outputs(1637) <= b and not a;
    layer1_outputs(1638) <= '0';
    layer1_outputs(1639) <= a and not b;
    layer1_outputs(1640) <= not b or a;
    layer1_outputs(1641) <= not b;
    layer1_outputs(1642) <= not b or a;
    layer1_outputs(1643) <= not (a and b);
    layer1_outputs(1644) <= a and not b;
    layer1_outputs(1645) <= a and not b;
    layer1_outputs(1646) <= a and not b;
    layer1_outputs(1647) <= not b;
    layer1_outputs(1648) <= not a;
    layer1_outputs(1649) <= a xor b;
    layer1_outputs(1650) <= a and b;
    layer1_outputs(1651) <= a and not b;
    layer1_outputs(1652) <= not (a and b);
    layer1_outputs(1653) <= not b;
    layer1_outputs(1654) <= not b or a;
    layer1_outputs(1655) <= b;
    layer1_outputs(1656) <= '0';
    layer1_outputs(1657) <= not b;
    layer1_outputs(1658) <= a;
    layer1_outputs(1659) <= not b;
    layer1_outputs(1660) <= a xor b;
    layer1_outputs(1661) <= a and not b;
    layer1_outputs(1662) <= b;
    layer1_outputs(1663) <= not b;
    layer1_outputs(1664) <= not (a or b);
    layer1_outputs(1665) <= a or b;
    layer1_outputs(1666) <= a and not b;
    layer1_outputs(1667) <= not a;
    layer1_outputs(1668) <= not (a or b);
    layer1_outputs(1669) <= a;
    layer1_outputs(1670) <= a;
    layer1_outputs(1671) <= a;
    layer1_outputs(1672) <= b;
    layer1_outputs(1673) <= a;
    layer1_outputs(1674) <= not b or a;
    layer1_outputs(1675) <= not a or b;
    layer1_outputs(1676) <= not b;
    layer1_outputs(1677) <= a and b;
    layer1_outputs(1678) <= a and not b;
    layer1_outputs(1679) <= not a;
    layer1_outputs(1680) <= not (a and b);
    layer1_outputs(1681) <= not b;
    layer1_outputs(1682) <= b and not a;
    layer1_outputs(1683) <= not (a or b);
    layer1_outputs(1684) <= '0';
    layer1_outputs(1685) <= not a;
    layer1_outputs(1686) <= b and not a;
    layer1_outputs(1687) <= not b or a;
    layer1_outputs(1688) <= a or b;
    layer1_outputs(1689) <= '0';
    layer1_outputs(1690) <= b;
    layer1_outputs(1691) <= not (a xor b);
    layer1_outputs(1692) <= not a or b;
    layer1_outputs(1693) <= not b or a;
    layer1_outputs(1694) <= not a;
    layer1_outputs(1695) <= not (a and b);
    layer1_outputs(1696) <= '1';
    layer1_outputs(1697) <= not a;
    layer1_outputs(1698) <= a and not b;
    layer1_outputs(1699) <= not (a xor b);
    layer1_outputs(1700) <= a and not b;
    layer1_outputs(1701) <= b;
    layer1_outputs(1702) <= not a or b;
    layer1_outputs(1703) <= a;
    layer1_outputs(1704) <= not (a and b);
    layer1_outputs(1705) <= not b or a;
    layer1_outputs(1706) <= not b;
    layer1_outputs(1707) <= a and not b;
    layer1_outputs(1708) <= a;
    layer1_outputs(1709) <= not (a or b);
    layer1_outputs(1710) <= '0';
    layer1_outputs(1711) <= b;
    layer1_outputs(1712) <= b and not a;
    layer1_outputs(1713) <= b;
    layer1_outputs(1714) <= not (a xor b);
    layer1_outputs(1715) <= not a;
    layer1_outputs(1716) <= not b or a;
    layer1_outputs(1717) <= b and not a;
    layer1_outputs(1718) <= not a;
    layer1_outputs(1719) <= not a;
    layer1_outputs(1720) <= b;
    layer1_outputs(1721) <= b;
    layer1_outputs(1722) <= b and not a;
    layer1_outputs(1723) <= a;
    layer1_outputs(1724) <= not a;
    layer1_outputs(1725) <= b;
    layer1_outputs(1726) <= a and b;
    layer1_outputs(1727) <= a and not b;
    layer1_outputs(1728) <= not (a xor b);
    layer1_outputs(1729) <= a and b;
    layer1_outputs(1730) <= not b or a;
    layer1_outputs(1731) <= b and not a;
    layer1_outputs(1732) <= not a or b;
    layer1_outputs(1733) <= not (a and b);
    layer1_outputs(1734) <= not b;
    layer1_outputs(1735) <= not b;
    layer1_outputs(1736) <= a;
    layer1_outputs(1737) <= a;
    layer1_outputs(1738) <= b;
    layer1_outputs(1739) <= a and not b;
    layer1_outputs(1740) <= a and not b;
    layer1_outputs(1741) <= '1';
    layer1_outputs(1742) <= a and b;
    layer1_outputs(1743) <= not a or b;
    layer1_outputs(1744) <= '1';
    layer1_outputs(1745) <= not a or b;
    layer1_outputs(1746) <= a or b;
    layer1_outputs(1747) <= a and b;
    layer1_outputs(1748) <= not b;
    layer1_outputs(1749) <= not a or b;
    layer1_outputs(1750) <= a;
    layer1_outputs(1751) <= not a;
    layer1_outputs(1752) <= b and not a;
    layer1_outputs(1753) <= a xor b;
    layer1_outputs(1754) <= '1';
    layer1_outputs(1755) <= b;
    layer1_outputs(1756) <= b and not a;
    layer1_outputs(1757) <= b and not a;
    layer1_outputs(1758) <= a and b;
    layer1_outputs(1759) <= not a or b;
    layer1_outputs(1760) <= not (a xor b);
    layer1_outputs(1761) <= a and not b;
    layer1_outputs(1762) <= not a or b;
    layer1_outputs(1763) <= a;
    layer1_outputs(1764) <= not (a and b);
    layer1_outputs(1765) <= a and not b;
    layer1_outputs(1766) <= not a;
    layer1_outputs(1767) <= b and not a;
    layer1_outputs(1768) <= b;
    layer1_outputs(1769) <= a and not b;
    layer1_outputs(1770) <= not (a and b);
    layer1_outputs(1771) <= not a;
    layer1_outputs(1772) <= a and not b;
    layer1_outputs(1773) <= a xor b;
    layer1_outputs(1774) <= not a;
    layer1_outputs(1775) <= not a;
    layer1_outputs(1776) <= '0';
    layer1_outputs(1777) <= a and b;
    layer1_outputs(1778) <= not b or a;
    layer1_outputs(1779) <= b;
    layer1_outputs(1780) <= not b or a;
    layer1_outputs(1781) <= a;
    layer1_outputs(1782) <= a;
    layer1_outputs(1783) <= not a;
    layer1_outputs(1784) <= not b;
    layer1_outputs(1785) <= b;
    layer1_outputs(1786) <= not a or b;
    layer1_outputs(1787) <= not (a and b);
    layer1_outputs(1788) <= a and not b;
    layer1_outputs(1789) <= b and not a;
    layer1_outputs(1790) <= b and not a;
    layer1_outputs(1791) <= '0';
    layer1_outputs(1792) <= a;
    layer1_outputs(1793) <= b and not a;
    layer1_outputs(1794) <= not (a and b);
    layer1_outputs(1795) <= a and b;
    layer1_outputs(1796) <= not a;
    layer1_outputs(1797) <= not a or b;
    layer1_outputs(1798) <= not (a and b);
    layer1_outputs(1799) <= a or b;
    layer1_outputs(1800) <= '0';
    layer1_outputs(1801) <= a xor b;
    layer1_outputs(1802) <= a and b;
    layer1_outputs(1803) <= not a or b;
    layer1_outputs(1804) <= b;
    layer1_outputs(1805) <= '1';
    layer1_outputs(1806) <= not a or b;
    layer1_outputs(1807) <= not (a or b);
    layer1_outputs(1808) <= a xor b;
    layer1_outputs(1809) <= not a;
    layer1_outputs(1810) <= a and b;
    layer1_outputs(1811) <= '1';
    layer1_outputs(1812) <= '0';
    layer1_outputs(1813) <= a and b;
    layer1_outputs(1814) <= '0';
    layer1_outputs(1815) <= not (a or b);
    layer1_outputs(1816) <= not (a and b);
    layer1_outputs(1817) <= not (a or b);
    layer1_outputs(1818) <= not a;
    layer1_outputs(1819) <= b;
    layer1_outputs(1820) <= a and not b;
    layer1_outputs(1821) <= a or b;
    layer1_outputs(1822) <= a and not b;
    layer1_outputs(1823) <= a and b;
    layer1_outputs(1824) <= b;
    layer1_outputs(1825) <= not (a and b);
    layer1_outputs(1826) <= not a;
    layer1_outputs(1827) <= a and b;
    layer1_outputs(1828) <= b and not a;
    layer1_outputs(1829) <= a or b;
    layer1_outputs(1830) <= '0';
    layer1_outputs(1831) <= b and not a;
    layer1_outputs(1832) <= not b;
    layer1_outputs(1833) <= not a or b;
    layer1_outputs(1834) <= a and b;
    layer1_outputs(1835) <= a;
    layer1_outputs(1836) <= b;
    layer1_outputs(1837) <= a xor b;
    layer1_outputs(1838) <= not a;
    layer1_outputs(1839) <= not (a and b);
    layer1_outputs(1840) <= not (a and b);
    layer1_outputs(1841) <= b;
    layer1_outputs(1842) <= not b;
    layer1_outputs(1843) <= b;
    layer1_outputs(1844) <= not (a xor b);
    layer1_outputs(1845) <= b;
    layer1_outputs(1846) <= b;
    layer1_outputs(1847) <= not (a xor b);
    layer1_outputs(1848) <= a xor b;
    layer1_outputs(1849) <= a and b;
    layer1_outputs(1850) <= not (a and b);
    layer1_outputs(1851) <= a;
    layer1_outputs(1852) <= not (a or b);
    layer1_outputs(1853) <= not b;
    layer1_outputs(1854) <= b and not a;
    layer1_outputs(1855) <= a or b;
    layer1_outputs(1856) <= not (a and b);
    layer1_outputs(1857) <= not a;
    layer1_outputs(1858) <= not (a or b);
    layer1_outputs(1859) <= '1';
    layer1_outputs(1860) <= not a;
    layer1_outputs(1861) <= not a;
    layer1_outputs(1862) <= not (a or b);
    layer1_outputs(1863) <= b and not a;
    layer1_outputs(1864) <= a and b;
    layer1_outputs(1865) <= a;
    layer1_outputs(1866) <= a and not b;
    layer1_outputs(1867) <= not a;
    layer1_outputs(1868) <= a or b;
    layer1_outputs(1869) <= not b or a;
    layer1_outputs(1870) <= a;
    layer1_outputs(1871) <= not b or a;
    layer1_outputs(1872) <= a and b;
    layer1_outputs(1873) <= a or b;
    layer1_outputs(1874) <= a and b;
    layer1_outputs(1875) <= not a or b;
    layer1_outputs(1876) <= a and b;
    layer1_outputs(1877) <= not (a xor b);
    layer1_outputs(1878) <= not a;
    layer1_outputs(1879) <= '1';
    layer1_outputs(1880) <= a or b;
    layer1_outputs(1881) <= a or b;
    layer1_outputs(1882) <= '0';
    layer1_outputs(1883) <= not a;
    layer1_outputs(1884) <= not (a xor b);
    layer1_outputs(1885) <= a and b;
    layer1_outputs(1886) <= a;
    layer1_outputs(1887) <= not b or a;
    layer1_outputs(1888) <= not b;
    layer1_outputs(1889) <= a or b;
    layer1_outputs(1890) <= not b or a;
    layer1_outputs(1891) <= not a;
    layer1_outputs(1892) <= '0';
    layer1_outputs(1893) <= '0';
    layer1_outputs(1894) <= not b;
    layer1_outputs(1895) <= a and not b;
    layer1_outputs(1896) <= not (a and b);
    layer1_outputs(1897) <= not a;
    layer1_outputs(1898) <= a and not b;
    layer1_outputs(1899) <= not (a and b);
    layer1_outputs(1900) <= a and b;
    layer1_outputs(1901) <= a;
    layer1_outputs(1902) <= a and not b;
    layer1_outputs(1903) <= b;
    layer1_outputs(1904) <= b;
    layer1_outputs(1905) <= not (a xor b);
    layer1_outputs(1906) <= a;
    layer1_outputs(1907) <= a or b;
    layer1_outputs(1908) <= not (a xor b);
    layer1_outputs(1909) <= not b or a;
    layer1_outputs(1910) <= not b;
    layer1_outputs(1911) <= not (a or b);
    layer1_outputs(1912) <= not b;
    layer1_outputs(1913) <= not (a and b);
    layer1_outputs(1914) <= a;
    layer1_outputs(1915) <= a;
    layer1_outputs(1916) <= a and b;
    layer1_outputs(1917) <= b and not a;
    layer1_outputs(1918) <= not (a and b);
    layer1_outputs(1919) <= a and b;
    layer1_outputs(1920) <= a and b;
    layer1_outputs(1921) <= not (a or b);
    layer1_outputs(1922) <= not a;
    layer1_outputs(1923) <= not b or a;
    layer1_outputs(1924) <= a and b;
    layer1_outputs(1925) <= a xor b;
    layer1_outputs(1926) <= not (a or b);
    layer1_outputs(1927) <= b and not a;
    layer1_outputs(1928) <= b;
    layer1_outputs(1929) <= '0';
    layer1_outputs(1930) <= '0';
    layer1_outputs(1931) <= b and not a;
    layer1_outputs(1932) <= not a;
    layer1_outputs(1933) <= not a or b;
    layer1_outputs(1934) <= b and not a;
    layer1_outputs(1935) <= b;
    layer1_outputs(1936) <= b and not a;
    layer1_outputs(1937) <= a;
    layer1_outputs(1938) <= not b or a;
    layer1_outputs(1939) <= not (a or b);
    layer1_outputs(1940) <= a xor b;
    layer1_outputs(1941) <= a;
    layer1_outputs(1942) <= not a or b;
    layer1_outputs(1943) <= b;
    layer1_outputs(1944) <= a and b;
    layer1_outputs(1945) <= a;
    layer1_outputs(1946) <= not (a and b);
    layer1_outputs(1947) <= b and not a;
    layer1_outputs(1948) <= '0';
    layer1_outputs(1949) <= not (a or b);
    layer1_outputs(1950) <= not a or b;
    layer1_outputs(1951) <= a or b;
    layer1_outputs(1952) <= a and not b;
    layer1_outputs(1953) <= b;
    layer1_outputs(1954) <= a;
    layer1_outputs(1955) <= not (a and b);
    layer1_outputs(1956) <= b;
    layer1_outputs(1957) <= not (a and b);
    layer1_outputs(1958) <= not b;
    layer1_outputs(1959) <= not a or b;
    layer1_outputs(1960) <= b;
    layer1_outputs(1961) <= '0';
    layer1_outputs(1962) <= b;
    layer1_outputs(1963) <= b;
    layer1_outputs(1964) <= not a or b;
    layer1_outputs(1965) <= not a or b;
    layer1_outputs(1966) <= a xor b;
    layer1_outputs(1967) <= not b or a;
    layer1_outputs(1968) <= b;
    layer1_outputs(1969) <= a or b;
    layer1_outputs(1970) <= not (a and b);
    layer1_outputs(1971) <= not b;
    layer1_outputs(1972) <= a or b;
    layer1_outputs(1973) <= not b;
    layer1_outputs(1974) <= not a;
    layer1_outputs(1975) <= not (a xor b);
    layer1_outputs(1976) <= a;
    layer1_outputs(1977) <= a;
    layer1_outputs(1978) <= a and b;
    layer1_outputs(1979) <= a xor b;
    layer1_outputs(1980) <= b and not a;
    layer1_outputs(1981) <= a;
    layer1_outputs(1982) <= a;
    layer1_outputs(1983) <= '1';
    layer1_outputs(1984) <= a and not b;
    layer1_outputs(1985) <= not b;
    layer1_outputs(1986) <= not (a and b);
    layer1_outputs(1987) <= not b or a;
    layer1_outputs(1988) <= a or b;
    layer1_outputs(1989) <= not a or b;
    layer1_outputs(1990) <= not b or a;
    layer1_outputs(1991) <= b and not a;
    layer1_outputs(1992) <= a and b;
    layer1_outputs(1993) <= a and not b;
    layer1_outputs(1994) <= a and b;
    layer1_outputs(1995) <= a;
    layer1_outputs(1996) <= b and not a;
    layer1_outputs(1997) <= not b or a;
    layer1_outputs(1998) <= not b or a;
    layer1_outputs(1999) <= not a;
    layer1_outputs(2000) <= not b;
    layer1_outputs(2001) <= not b or a;
    layer1_outputs(2002) <= a or b;
    layer1_outputs(2003) <= not (a and b);
    layer1_outputs(2004) <= not (a xor b);
    layer1_outputs(2005) <= '1';
    layer1_outputs(2006) <= b;
    layer1_outputs(2007) <= '0';
    layer1_outputs(2008) <= '0';
    layer1_outputs(2009) <= a or b;
    layer1_outputs(2010) <= not a;
    layer1_outputs(2011) <= not b;
    layer1_outputs(2012) <= b;
    layer1_outputs(2013) <= not b;
    layer1_outputs(2014) <= a and not b;
    layer1_outputs(2015) <= not a or b;
    layer1_outputs(2016) <= a and not b;
    layer1_outputs(2017) <= a;
    layer1_outputs(2018) <= a or b;
    layer1_outputs(2019) <= not b;
    layer1_outputs(2020) <= not (a or b);
    layer1_outputs(2021) <= not b;
    layer1_outputs(2022) <= a or b;
    layer1_outputs(2023) <= not (a and b);
    layer1_outputs(2024) <= not a or b;
    layer1_outputs(2025) <= not b or a;
    layer1_outputs(2026) <= not a or b;
    layer1_outputs(2027) <= not b;
    layer1_outputs(2028) <= a or b;
    layer1_outputs(2029) <= a or b;
    layer1_outputs(2030) <= not a;
    layer1_outputs(2031) <= b;
    layer1_outputs(2032) <= not (a xor b);
    layer1_outputs(2033) <= not b;
    layer1_outputs(2034) <= not a or b;
    layer1_outputs(2035) <= a and not b;
    layer1_outputs(2036) <= not a;
    layer1_outputs(2037) <= a;
    layer1_outputs(2038) <= b and not a;
    layer1_outputs(2039) <= not b or a;
    layer1_outputs(2040) <= a xor b;
    layer1_outputs(2041) <= not b or a;
    layer1_outputs(2042) <= not a;
    layer1_outputs(2043) <= not a or b;
    layer1_outputs(2044) <= not a;
    layer1_outputs(2045) <= not a;
    layer1_outputs(2046) <= not (a and b);
    layer1_outputs(2047) <= not (a or b);
    layer1_outputs(2048) <= a and b;
    layer1_outputs(2049) <= a;
    layer1_outputs(2050) <= not b or a;
    layer1_outputs(2051) <= a and b;
    layer1_outputs(2052) <= not (a and b);
    layer1_outputs(2053) <= not b;
    layer1_outputs(2054) <= not (a and b);
    layer1_outputs(2055) <= '0';
    layer1_outputs(2056) <= b and not a;
    layer1_outputs(2057) <= not a;
    layer1_outputs(2058) <= a xor b;
    layer1_outputs(2059) <= a;
    layer1_outputs(2060) <= b;
    layer1_outputs(2061) <= not (a and b);
    layer1_outputs(2062) <= not a;
    layer1_outputs(2063) <= not a;
    layer1_outputs(2064) <= a or b;
    layer1_outputs(2065) <= not (a and b);
    layer1_outputs(2066) <= not b or a;
    layer1_outputs(2067) <= b;
    layer1_outputs(2068) <= a and not b;
    layer1_outputs(2069) <= not (a or b);
    layer1_outputs(2070) <= a or b;
    layer1_outputs(2071) <= a and not b;
    layer1_outputs(2072) <= a;
    layer1_outputs(2073) <= not a or b;
    layer1_outputs(2074) <= a and b;
    layer1_outputs(2075) <= not a or b;
    layer1_outputs(2076) <= not a;
    layer1_outputs(2077) <= not a;
    layer1_outputs(2078) <= not (a or b);
    layer1_outputs(2079) <= not b or a;
    layer1_outputs(2080) <= not (a and b);
    layer1_outputs(2081) <= not (a and b);
    layer1_outputs(2082) <= not b or a;
    layer1_outputs(2083) <= not a;
    layer1_outputs(2084) <= not (a and b);
    layer1_outputs(2085) <= b;
    layer1_outputs(2086) <= not b;
    layer1_outputs(2087) <= a xor b;
    layer1_outputs(2088) <= a;
    layer1_outputs(2089) <= a;
    layer1_outputs(2090) <= not a;
    layer1_outputs(2091) <= b and not a;
    layer1_outputs(2092) <= b;
    layer1_outputs(2093) <= not b or a;
    layer1_outputs(2094) <= b and not a;
    layer1_outputs(2095) <= b;
    layer1_outputs(2096) <= not b;
    layer1_outputs(2097) <= b;
    layer1_outputs(2098) <= b;
    layer1_outputs(2099) <= b;
    layer1_outputs(2100) <= not a;
    layer1_outputs(2101) <= a and not b;
    layer1_outputs(2102) <= a and not b;
    layer1_outputs(2103) <= not a;
    layer1_outputs(2104) <= not a;
    layer1_outputs(2105) <= a;
    layer1_outputs(2106) <= not (a xor b);
    layer1_outputs(2107) <= not (a and b);
    layer1_outputs(2108) <= '0';
    layer1_outputs(2109) <= not a;
    layer1_outputs(2110) <= a and not b;
    layer1_outputs(2111) <= not (a or b);
    layer1_outputs(2112) <= b;
    layer1_outputs(2113) <= a and not b;
    layer1_outputs(2114) <= a and b;
    layer1_outputs(2115) <= not a or b;
    layer1_outputs(2116) <= not (a or b);
    layer1_outputs(2117) <= not (a or b);
    layer1_outputs(2118) <= not b or a;
    layer1_outputs(2119) <= a and b;
    layer1_outputs(2120) <= b and not a;
    layer1_outputs(2121) <= not a;
    layer1_outputs(2122) <= not (a or b);
    layer1_outputs(2123) <= a and not b;
    layer1_outputs(2124) <= not (a xor b);
    layer1_outputs(2125) <= not b;
    layer1_outputs(2126) <= b and not a;
    layer1_outputs(2127) <= not a or b;
    layer1_outputs(2128) <= not a;
    layer1_outputs(2129) <= a and not b;
    layer1_outputs(2130) <= not a;
    layer1_outputs(2131) <= not b;
    layer1_outputs(2132) <= b and not a;
    layer1_outputs(2133) <= a;
    layer1_outputs(2134) <= b;
    layer1_outputs(2135) <= b;
    layer1_outputs(2136) <= '0';
    layer1_outputs(2137) <= a and b;
    layer1_outputs(2138) <= '0';
    layer1_outputs(2139) <= '0';
    layer1_outputs(2140) <= a and b;
    layer1_outputs(2141) <= b and not a;
    layer1_outputs(2142) <= a or b;
    layer1_outputs(2143) <= not (a and b);
    layer1_outputs(2144) <= a and b;
    layer1_outputs(2145) <= not b;
    layer1_outputs(2146) <= a or b;
    layer1_outputs(2147) <= a and not b;
    layer1_outputs(2148) <= a and b;
    layer1_outputs(2149) <= not (a or b);
    layer1_outputs(2150) <= a or b;
    layer1_outputs(2151) <= not b or a;
    layer1_outputs(2152) <= a and not b;
    layer1_outputs(2153) <= a;
    layer1_outputs(2154) <= b;
    layer1_outputs(2155) <= not a or b;
    layer1_outputs(2156) <= '1';
    layer1_outputs(2157) <= b and not a;
    layer1_outputs(2158) <= not a or b;
    layer1_outputs(2159) <= not a or b;
    layer1_outputs(2160) <= b and not a;
    layer1_outputs(2161) <= a and not b;
    layer1_outputs(2162) <= not (a and b);
    layer1_outputs(2163) <= '0';
    layer1_outputs(2164) <= not b or a;
    layer1_outputs(2165) <= a;
    layer1_outputs(2166) <= not b or a;
    layer1_outputs(2167) <= b and not a;
    layer1_outputs(2168) <= not a or b;
    layer1_outputs(2169) <= a;
    layer1_outputs(2170) <= b;
    layer1_outputs(2171) <= a or b;
    layer1_outputs(2172) <= a and not b;
    layer1_outputs(2173) <= not b or a;
    layer1_outputs(2174) <= not b or a;
    layer1_outputs(2175) <= not a or b;
    layer1_outputs(2176) <= not a or b;
    layer1_outputs(2177) <= not a;
    layer1_outputs(2178) <= not (a xor b);
    layer1_outputs(2179) <= not a;
    layer1_outputs(2180) <= b;
    layer1_outputs(2181) <= b;
    layer1_outputs(2182) <= '1';
    layer1_outputs(2183) <= b;
    layer1_outputs(2184) <= a xor b;
    layer1_outputs(2185) <= not a or b;
    layer1_outputs(2186) <= not a;
    layer1_outputs(2187) <= not (a or b);
    layer1_outputs(2188) <= a and b;
    layer1_outputs(2189) <= a and b;
    layer1_outputs(2190) <= b;
    layer1_outputs(2191) <= a and not b;
    layer1_outputs(2192) <= not b or a;
    layer1_outputs(2193) <= not (a or b);
    layer1_outputs(2194) <= a and b;
    layer1_outputs(2195) <= b and not a;
    layer1_outputs(2196) <= a xor b;
    layer1_outputs(2197) <= a;
    layer1_outputs(2198) <= not (a or b);
    layer1_outputs(2199) <= a or b;
    layer1_outputs(2200) <= b and not a;
    layer1_outputs(2201) <= a;
    layer1_outputs(2202) <= a xor b;
    layer1_outputs(2203) <= not a;
    layer1_outputs(2204) <= not a or b;
    layer1_outputs(2205) <= not b;
    layer1_outputs(2206) <= not a;
    layer1_outputs(2207) <= not (a or b);
    layer1_outputs(2208) <= b and not a;
    layer1_outputs(2209) <= not a or b;
    layer1_outputs(2210) <= a;
    layer1_outputs(2211) <= not b;
    layer1_outputs(2212) <= not a;
    layer1_outputs(2213) <= a;
    layer1_outputs(2214) <= a or b;
    layer1_outputs(2215) <= not a;
    layer1_outputs(2216) <= a xor b;
    layer1_outputs(2217) <= '0';
    layer1_outputs(2218) <= a;
    layer1_outputs(2219) <= not (a and b);
    layer1_outputs(2220) <= a and b;
    layer1_outputs(2221) <= '1';
    layer1_outputs(2222) <= not (a and b);
    layer1_outputs(2223) <= a and not b;
    layer1_outputs(2224) <= not b or a;
    layer1_outputs(2225) <= not a;
    layer1_outputs(2226) <= a or b;
    layer1_outputs(2227) <= not a;
    layer1_outputs(2228) <= a and b;
    layer1_outputs(2229) <= b and not a;
    layer1_outputs(2230) <= not (a and b);
    layer1_outputs(2231) <= a xor b;
    layer1_outputs(2232) <= not b or a;
    layer1_outputs(2233) <= not (a and b);
    layer1_outputs(2234) <= a;
    layer1_outputs(2235) <= a and b;
    layer1_outputs(2236) <= a and b;
    layer1_outputs(2237) <= a or b;
    layer1_outputs(2238) <= b;
    layer1_outputs(2239) <= b and not a;
    layer1_outputs(2240) <= a and not b;
    layer1_outputs(2241) <= b and not a;
    layer1_outputs(2242) <= a;
    layer1_outputs(2243) <= a and b;
    layer1_outputs(2244) <= not (a xor b);
    layer1_outputs(2245) <= not a or b;
    layer1_outputs(2246) <= not (a or b);
    layer1_outputs(2247) <= not a;
    layer1_outputs(2248) <= not a;
    layer1_outputs(2249) <= b;
    layer1_outputs(2250) <= not (a xor b);
    layer1_outputs(2251) <= '0';
    layer1_outputs(2252) <= a and not b;
    layer1_outputs(2253) <= not (a or b);
    layer1_outputs(2254) <= not b;
    layer1_outputs(2255) <= a and b;
    layer1_outputs(2256) <= not a or b;
    layer1_outputs(2257) <= '0';
    layer1_outputs(2258) <= not a or b;
    layer1_outputs(2259) <= not (a and b);
    layer1_outputs(2260) <= a or b;
    layer1_outputs(2261) <= a and b;
    layer1_outputs(2262) <= '0';
    layer1_outputs(2263) <= not b;
    layer1_outputs(2264) <= b and not a;
    layer1_outputs(2265) <= a;
    layer1_outputs(2266) <= not b or a;
    layer1_outputs(2267) <= not b;
    layer1_outputs(2268) <= not b;
    layer1_outputs(2269) <= b;
    layer1_outputs(2270) <= a xor b;
    layer1_outputs(2271) <= a;
    layer1_outputs(2272) <= not a;
    layer1_outputs(2273) <= a and b;
    layer1_outputs(2274) <= '0';
    layer1_outputs(2275) <= not b or a;
    layer1_outputs(2276) <= not a;
    layer1_outputs(2277) <= not b;
    layer1_outputs(2278) <= b;
    layer1_outputs(2279) <= not b;
    layer1_outputs(2280) <= not (a and b);
    layer1_outputs(2281) <= not (a or b);
    layer1_outputs(2282) <= not (a and b);
    layer1_outputs(2283) <= '1';
    layer1_outputs(2284) <= '0';
    layer1_outputs(2285) <= not a;
    layer1_outputs(2286) <= not a;
    layer1_outputs(2287) <= a xor b;
    layer1_outputs(2288) <= not (a and b);
    layer1_outputs(2289) <= a;
    layer1_outputs(2290) <= a or b;
    layer1_outputs(2291) <= '1';
    layer1_outputs(2292) <= a xor b;
    layer1_outputs(2293) <= a or b;
    layer1_outputs(2294) <= not a;
    layer1_outputs(2295) <= '0';
    layer1_outputs(2296) <= a and b;
    layer1_outputs(2297) <= a and b;
    layer1_outputs(2298) <= '1';
    layer1_outputs(2299) <= not b;
    layer1_outputs(2300) <= not a;
    layer1_outputs(2301) <= a;
    layer1_outputs(2302) <= not (a and b);
    layer1_outputs(2303) <= a xor b;
    layer1_outputs(2304) <= a and b;
    layer1_outputs(2305) <= a;
    layer1_outputs(2306) <= a;
    layer1_outputs(2307) <= b and not a;
    layer1_outputs(2308) <= not b;
    layer1_outputs(2309) <= a;
    layer1_outputs(2310) <= a and not b;
    layer1_outputs(2311) <= not (a and b);
    layer1_outputs(2312) <= a;
    layer1_outputs(2313) <= '1';
    layer1_outputs(2314) <= a;
    layer1_outputs(2315) <= not b;
    layer1_outputs(2316) <= not b;
    layer1_outputs(2317) <= a;
    layer1_outputs(2318) <= a and b;
    layer1_outputs(2319) <= not a or b;
    layer1_outputs(2320) <= b and not a;
    layer1_outputs(2321) <= not a or b;
    layer1_outputs(2322) <= not (a xor b);
    layer1_outputs(2323) <= not (a and b);
    layer1_outputs(2324) <= not (a or b);
    layer1_outputs(2325) <= a;
    layer1_outputs(2326) <= '1';
    layer1_outputs(2327) <= a and b;
    layer1_outputs(2328) <= not a;
    layer1_outputs(2329) <= a and b;
    layer1_outputs(2330) <= not a;
    layer1_outputs(2331) <= a xor b;
    layer1_outputs(2332) <= not b;
    layer1_outputs(2333) <= a;
    layer1_outputs(2334) <= not (a and b);
    layer1_outputs(2335) <= not a;
    layer1_outputs(2336) <= not (a or b);
    layer1_outputs(2337) <= not (a and b);
    layer1_outputs(2338) <= a or b;
    layer1_outputs(2339) <= not (a and b);
    layer1_outputs(2340) <= a;
    layer1_outputs(2341) <= a;
    layer1_outputs(2342) <= not (a or b);
    layer1_outputs(2343) <= not b;
    layer1_outputs(2344) <= '0';
    layer1_outputs(2345) <= not (a or b);
    layer1_outputs(2346) <= not a or b;
    layer1_outputs(2347) <= not a or b;
    layer1_outputs(2348) <= not a;
    layer1_outputs(2349) <= '0';
    layer1_outputs(2350) <= '0';
    layer1_outputs(2351) <= a xor b;
    layer1_outputs(2352) <= b;
    layer1_outputs(2353) <= b and not a;
    layer1_outputs(2354) <= a and b;
    layer1_outputs(2355) <= a or b;
    layer1_outputs(2356) <= a or b;
    layer1_outputs(2357) <= b and not a;
    layer1_outputs(2358) <= not a or b;
    layer1_outputs(2359) <= '0';
    layer1_outputs(2360) <= not (a or b);
    layer1_outputs(2361) <= not (a xor b);
    layer1_outputs(2362) <= b;
    layer1_outputs(2363) <= '1';
    layer1_outputs(2364) <= a;
    layer1_outputs(2365) <= b;
    layer1_outputs(2366) <= a;
    layer1_outputs(2367) <= a or b;
    layer1_outputs(2368) <= '1';
    layer1_outputs(2369) <= a and b;
    layer1_outputs(2370) <= not (a and b);
    layer1_outputs(2371) <= not a;
    layer1_outputs(2372) <= not (a and b);
    layer1_outputs(2373) <= not a or b;
    layer1_outputs(2374) <= not b;
    layer1_outputs(2375) <= '1';
    layer1_outputs(2376) <= not (a or b);
    layer1_outputs(2377) <= not (a and b);
    layer1_outputs(2378) <= not b;
    layer1_outputs(2379) <= a;
    layer1_outputs(2380) <= '1';
    layer1_outputs(2381) <= b and not a;
    layer1_outputs(2382) <= not b;
    layer1_outputs(2383) <= a and not b;
    layer1_outputs(2384) <= a;
    layer1_outputs(2385) <= b and not a;
    layer1_outputs(2386) <= not b or a;
    layer1_outputs(2387) <= not a or b;
    layer1_outputs(2388) <= '1';
    layer1_outputs(2389) <= not (a or b);
    layer1_outputs(2390) <= a xor b;
    layer1_outputs(2391) <= b;
    layer1_outputs(2392) <= not b;
    layer1_outputs(2393) <= a or b;
    layer1_outputs(2394) <= not b;
    layer1_outputs(2395) <= not b or a;
    layer1_outputs(2396) <= a and not b;
    layer1_outputs(2397) <= not a or b;
    layer1_outputs(2398) <= not a;
    layer1_outputs(2399) <= not a;
    layer1_outputs(2400) <= a and b;
    layer1_outputs(2401) <= b;
    layer1_outputs(2402) <= '0';
    layer1_outputs(2403) <= '0';
    layer1_outputs(2404) <= not a;
    layer1_outputs(2405) <= not (a or b);
    layer1_outputs(2406) <= not (a or b);
    layer1_outputs(2407) <= a and not b;
    layer1_outputs(2408) <= a and not b;
    layer1_outputs(2409) <= not (a and b);
    layer1_outputs(2410) <= b;
    layer1_outputs(2411) <= a or b;
    layer1_outputs(2412) <= not (a and b);
    layer1_outputs(2413) <= not a;
    layer1_outputs(2414) <= not (a and b);
    layer1_outputs(2415) <= b and not a;
    layer1_outputs(2416) <= b;
    layer1_outputs(2417) <= a;
    layer1_outputs(2418) <= not a;
    layer1_outputs(2419) <= b and not a;
    layer1_outputs(2420) <= not a or b;
    layer1_outputs(2421) <= not b;
    layer1_outputs(2422) <= a or b;
    layer1_outputs(2423) <= not b;
    layer1_outputs(2424) <= '0';
    layer1_outputs(2425) <= a;
    layer1_outputs(2426) <= b and not a;
    layer1_outputs(2427) <= not a;
    layer1_outputs(2428) <= a;
    layer1_outputs(2429) <= a;
    layer1_outputs(2430) <= not a;
    layer1_outputs(2431) <= a and not b;
    layer1_outputs(2432) <= a xor b;
    layer1_outputs(2433) <= '1';
    layer1_outputs(2434) <= not b;
    layer1_outputs(2435) <= not (a or b);
    layer1_outputs(2436) <= '0';
    layer1_outputs(2437) <= b and not a;
    layer1_outputs(2438) <= b and not a;
    layer1_outputs(2439) <= not (a or b);
    layer1_outputs(2440) <= not a;
    layer1_outputs(2441) <= b and not a;
    layer1_outputs(2442) <= not b or a;
    layer1_outputs(2443) <= not (a xor b);
    layer1_outputs(2444) <= not (a xor b);
    layer1_outputs(2445) <= not (a and b);
    layer1_outputs(2446) <= a or b;
    layer1_outputs(2447) <= not (a or b);
    layer1_outputs(2448) <= a;
    layer1_outputs(2449) <= not a or b;
    layer1_outputs(2450) <= a and not b;
    layer1_outputs(2451) <= b;
    layer1_outputs(2452) <= a;
    layer1_outputs(2453) <= a and b;
    layer1_outputs(2454) <= a;
    layer1_outputs(2455) <= b;
    layer1_outputs(2456) <= b;
    layer1_outputs(2457) <= not b or a;
    layer1_outputs(2458) <= not b or a;
    layer1_outputs(2459) <= not a or b;
    layer1_outputs(2460) <= b and not a;
    layer1_outputs(2461) <= b and not a;
    layer1_outputs(2462) <= '0';
    layer1_outputs(2463) <= b;
    layer1_outputs(2464) <= a and b;
    layer1_outputs(2465) <= not a;
    layer1_outputs(2466) <= a or b;
    layer1_outputs(2467) <= b;
    layer1_outputs(2468) <= not (a or b);
    layer1_outputs(2469) <= not (a or b);
    layer1_outputs(2470) <= not (a and b);
    layer1_outputs(2471) <= a and not b;
    layer1_outputs(2472) <= a;
    layer1_outputs(2473) <= not b;
    layer1_outputs(2474) <= not a;
    layer1_outputs(2475) <= b;
    layer1_outputs(2476) <= a or b;
    layer1_outputs(2477) <= not a;
    layer1_outputs(2478) <= not b;
    layer1_outputs(2479) <= not (a xor b);
    layer1_outputs(2480) <= a and not b;
    layer1_outputs(2481) <= not b or a;
    layer1_outputs(2482) <= a and not b;
    layer1_outputs(2483) <= b;
    layer1_outputs(2484) <= b;
    layer1_outputs(2485) <= '0';
    layer1_outputs(2486) <= a and b;
    layer1_outputs(2487) <= a and b;
    layer1_outputs(2488) <= a and b;
    layer1_outputs(2489) <= b;
    layer1_outputs(2490) <= not b or a;
    layer1_outputs(2491) <= b and not a;
    layer1_outputs(2492) <= not a or b;
    layer1_outputs(2493) <= a and not b;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= a;
    layer1_outputs(2496) <= '0';
    layer1_outputs(2497) <= b;
    layer1_outputs(2498) <= not a;
    layer1_outputs(2499) <= not b;
    layer1_outputs(2500) <= a and not b;
    layer1_outputs(2501) <= b and not a;
    layer1_outputs(2502) <= a;
    layer1_outputs(2503) <= not (a xor b);
    layer1_outputs(2504) <= b;
    layer1_outputs(2505) <= not (a xor b);
    layer1_outputs(2506) <= not b or a;
    layer1_outputs(2507) <= b;
    layer1_outputs(2508) <= a;
    layer1_outputs(2509) <= a xor b;
    layer1_outputs(2510) <= not (a xor b);
    layer1_outputs(2511) <= a and b;
    layer1_outputs(2512) <= not b;
    layer1_outputs(2513) <= a and not b;
    layer1_outputs(2514) <= b and not a;
    layer1_outputs(2515) <= '0';
    layer1_outputs(2516) <= b and not a;
    layer1_outputs(2517) <= a xor b;
    layer1_outputs(2518) <= a and b;
    layer1_outputs(2519) <= not a or b;
    layer1_outputs(2520) <= a;
    layer1_outputs(2521) <= not a or b;
    layer1_outputs(2522) <= not b;
    layer1_outputs(2523) <= b and not a;
    layer1_outputs(2524) <= not b or a;
    layer1_outputs(2525) <= a;
    layer1_outputs(2526) <= a xor b;
    layer1_outputs(2527) <= not (a or b);
    layer1_outputs(2528) <= not a or b;
    layer1_outputs(2529) <= not a or b;
    layer1_outputs(2530) <= not b or a;
    layer1_outputs(2531) <= b;
    layer1_outputs(2532) <= a xor b;
    layer1_outputs(2533) <= not a;
    layer1_outputs(2534) <= not a;
    layer1_outputs(2535) <= a;
    layer1_outputs(2536) <= not (a and b);
    layer1_outputs(2537) <= not a or b;
    layer1_outputs(2538) <= a and b;
    layer1_outputs(2539) <= b and not a;
    layer1_outputs(2540) <= not b or a;
    layer1_outputs(2541) <= not b;
    layer1_outputs(2542) <= not a or b;
    layer1_outputs(2543) <= a xor b;
    layer1_outputs(2544) <= not (a xor b);
    layer1_outputs(2545) <= not a or b;
    layer1_outputs(2546) <= b;
    layer1_outputs(2547) <= not a or b;
    layer1_outputs(2548) <= not a or b;
    layer1_outputs(2549) <= not b or a;
    layer1_outputs(2550) <= not a;
    layer1_outputs(2551) <= a and not b;
    layer1_outputs(2552) <= a;
    layer1_outputs(2553) <= b and not a;
    layer1_outputs(2554) <= '1';
    layer1_outputs(2555) <= not (a or b);
    layer1_outputs(2556) <= a or b;
    layer1_outputs(2557) <= '0';
    layer1_outputs(2558) <= not b;
    layer1_outputs(2559) <= a and not b;
    layer1_outputs(2560) <= not (a and b);
    layer1_outputs(2561) <= b;
    layer1_outputs(2562) <= a and not b;
    layer1_outputs(2563) <= a;
    layer1_outputs(2564) <= a;
    layer1_outputs(2565) <= not (a or b);
    layer1_outputs(2566) <= not a or b;
    layer1_outputs(2567) <= b and not a;
    layer1_outputs(2568) <= a;
    layer1_outputs(2569) <= a;
    layer1_outputs(2570) <= b;
    layer1_outputs(2571) <= not b or a;
    layer1_outputs(2572) <= b;
    layer1_outputs(2573) <= a and b;
    layer1_outputs(2574) <= not (a and b);
    layer1_outputs(2575) <= b;
    layer1_outputs(2576) <= not b or a;
    layer1_outputs(2577) <= not a;
    layer1_outputs(2578) <= not (a and b);
    layer1_outputs(2579) <= not a;
    layer1_outputs(2580) <= not b;
    layer1_outputs(2581) <= a;
    layer1_outputs(2582) <= a and not b;
    layer1_outputs(2583) <= not b;
    layer1_outputs(2584) <= not b or a;
    layer1_outputs(2585) <= a;
    layer1_outputs(2586) <= not b or a;
    layer1_outputs(2587) <= a xor b;
    layer1_outputs(2588) <= not (a and b);
    layer1_outputs(2589) <= a or b;
    layer1_outputs(2590) <= not (a and b);
    layer1_outputs(2591) <= a or b;
    layer1_outputs(2592) <= not b or a;
    layer1_outputs(2593) <= a xor b;
    layer1_outputs(2594) <= not b;
    layer1_outputs(2595) <= not a;
    layer1_outputs(2596) <= not b;
    layer1_outputs(2597) <= a or b;
    layer1_outputs(2598) <= not (a or b);
    layer1_outputs(2599) <= b and not a;
    layer1_outputs(2600) <= b and not a;
    layer1_outputs(2601) <= a and b;
    layer1_outputs(2602) <= a xor b;
    layer1_outputs(2603) <= not a or b;
    layer1_outputs(2604) <= b and not a;
    layer1_outputs(2605) <= b and not a;
    layer1_outputs(2606) <= a and not b;
    layer1_outputs(2607) <= a and b;
    layer1_outputs(2608) <= a and b;
    layer1_outputs(2609) <= a or b;
    layer1_outputs(2610) <= not a;
    layer1_outputs(2611) <= not a or b;
    layer1_outputs(2612) <= a;
    layer1_outputs(2613) <= a xor b;
    layer1_outputs(2614) <= b and not a;
    layer1_outputs(2615) <= not a;
    layer1_outputs(2616) <= not (a or b);
    layer1_outputs(2617) <= not (a and b);
    layer1_outputs(2618) <= not (a xor b);
    layer1_outputs(2619) <= not b;
    layer1_outputs(2620) <= a and not b;
    layer1_outputs(2621) <= not b;
    layer1_outputs(2622) <= not b or a;
    layer1_outputs(2623) <= not b;
    layer1_outputs(2624) <= '0';
    layer1_outputs(2625) <= a and b;
    layer1_outputs(2626) <= b;
    layer1_outputs(2627) <= a xor b;
    layer1_outputs(2628) <= not a;
    layer1_outputs(2629) <= '0';
    layer1_outputs(2630) <= not (a or b);
    layer1_outputs(2631) <= a xor b;
    layer1_outputs(2632) <= not a or b;
    layer1_outputs(2633) <= a or b;
    layer1_outputs(2634) <= not a;
    layer1_outputs(2635) <= not (a or b);
    layer1_outputs(2636) <= a xor b;
    layer1_outputs(2637) <= not (a or b);
    layer1_outputs(2638) <= b and not a;
    layer1_outputs(2639) <= not (a and b);
    layer1_outputs(2640) <= not (a or b);
    layer1_outputs(2641) <= b and not a;
    layer1_outputs(2642) <= not b;
    layer1_outputs(2643) <= b and not a;
    layer1_outputs(2644) <= a;
    layer1_outputs(2645) <= a;
    layer1_outputs(2646) <= not b or a;
    layer1_outputs(2647) <= b;
    layer1_outputs(2648) <= a and b;
    layer1_outputs(2649) <= a and not b;
    layer1_outputs(2650) <= not a or b;
    layer1_outputs(2651) <= '1';
    layer1_outputs(2652) <= b;
    layer1_outputs(2653) <= b;
    layer1_outputs(2654) <= '0';
    layer1_outputs(2655) <= not b or a;
    layer1_outputs(2656) <= b and not a;
    layer1_outputs(2657) <= not b or a;
    layer1_outputs(2658) <= a;
    layer1_outputs(2659) <= '0';
    layer1_outputs(2660) <= a;
    layer1_outputs(2661) <= '0';
    layer1_outputs(2662) <= not a;
    layer1_outputs(2663) <= not (a or b);
    layer1_outputs(2664) <= '1';
    layer1_outputs(2665) <= a;
    layer1_outputs(2666) <= a;
    layer1_outputs(2667) <= a or b;
    layer1_outputs(2668) <= a and b;
    layer1_outputs(2669) <= a;
    layer1_outputs(2670) <= a;
    layer1_outputs(2671) <= a and b;
    layer1_outputs(2672) <= not b or a;
    layer1_outputs(2673) <= not a;
    layer1_outputs(2674) <= a and b;
    layer1_outputs(2675) <= b;
    layer1_outputs(2676) <= not a or b;
    layer1_outputs(2677) <= not (a and b);
    layer1_outputs(2678) <= '0';
    layer1_outputs(2679) <= not (a xor b);
    layer1_outputs(2680) <= not (a xor b);
    layer1_outputs(2681) <= not b;
    layer1_outputs(2682) <= not a;
    layer1_outputs(2683) <= a;
    layer1_outputs(2684) <= '1';
    layer1_outputs(2685) <= a;
    layer1_outputs(2686) <= a;
    layer1_outputs(2687) <= b;
    layer1_outputs(2688) <= not b or a;
    layer1_outputs(2689) <= a;
    layer1_outputs(2690) <= not (a and b);
    layer1_outputs(2691) <= not (a or b);
    layer1_outputs(2692) <= not a or b;
    layer1_outputs(2693) <= b;
    layer1_outputs(2694) <= b;
    layer1_outputs(2695) <= not (a and b);
    layer1_outputs(2696) <= not a;
    layer1_outputs(2697) <= not (a xor b);
    layer1_outputs(2698) <= not a;
    layer1_outputs(2699) <= not b;
    layer1_outputs(2700) <= b and not a;
    layer1_outputs(2701) <= not b or a;
    layer1_outputs(2702) <= a xor b;
    layer1_outputs(2703) <= not (a and b);
    layer1_outputs(2704) <= not b;
    layer1_outputs(2705) <= b and not a;
    layer1_outputs(2706) <= a and not b;
    layer1_outputs(2707) <= a and not b;
    layer1_outputs(2708) <= not b or a;
    layer1_outputs(2709) <= b;
    layer1_outputs(2710) <= a;
    layer1_outputs(2711) <= a;
    layer1_outputs(2712) <= a and not b;
    layer1_outputs(2713) <= not b;
    layer1_outputs(2714) <= not b;
    layer1_outputs(2715) <= not a;
    layer1_outputs(2716) <= b;
    layer1_outputs(2717) <= not (a xor b);
    layer1_outputs(2718) <= b;
    layer1_outputs(2719) <= not a or b;
    layer1_outputs(2720) <= a or b;
    layer1_outputs(2721) <= a xor b;
    layer1_outputs(2722) <= not (a or b);
    layer1_outputs(2723) <= not a or b;
    layer1_outputs(2724) <= a and not b;
    layer1_outputs(2725) <= not a or b;
    layer1_outputs(2726) <= a and b;
    layer1_outputs(2727) <= a or b;
    layer1_outputs(2728) <= not b;
    layer1_outputs(2729) <= not b or a;
    layer1_outputs(2730) <= not (a or b);
    layer1_outputs(2731) <= b;
    layer1_outputs(2732) <= a and b;
    layer1_outputs(2733) <= not a or b;
    layer1_outputs(2734) <= not a;
    layer1_outputs(2735) <= a or b;
    layer1_outputs(2736) <= not (a and b);
    layer1_outputs(2737) <= a and b;
    layer1_outputs(2738) <= b and not a;
    layer1_outputs(2739) <= b and not a;
    layer1_outputs(2740) <= b;
    layer1_outputs(2741) <= not b;
    layer1_outputs(2742) <= a and not b;
    layer1_outputs(2743) <= b;
    layer1_outputs(2744) <= a;
    layer1_outputs(2745) <= a and b;
    layer1_outputs(2746) <= not b;
    layer1_outputs(2747) <= not (a or b);
    layer1_outputs(2748) <= a xor b;
    layer1_outputs(2749) <= not a;
    layer1_outputs(2750) <= '1';
    layer1_outputs(2751) <= a and b;
    layer1_outputs(2752) <= not b or a;
    layer1_outputs(2753) <= not (a and b);
    layer1_outputs(2754) <= not a or b;
    layer1_outputs(2755) <= a or b;
    layer1_outputs(2756) <= not a;
    layer1_outputs(2757) <= a;
    layer1_outputs(2758) <= not b;
    layer1_outputs(2759) <= a and b;
    layer1_outputs(2760) <= not a or b;
    layer1_outputs(2761) <= not b or a;
    layer1_outputs(2762) <= a xor b;
    layer1_outputs(2763) <= b;
    layer1_outputs(2764) <= a or b;
    layer1_outputs(2765) <= a and b;
    layer1_outputs(2766) <= a;
    layer1_outputs(2767) <= a;
    layer1_outputs(2768) <= a or b;
    layer1_outputs(2769) <= not a or b;
    layer1_outputs(2770) <= '0';
    layer1_outputs(2771) <= a or b;
    layer1_outputs(2772) <= b and not a;
    layer1_outputs(2773) <= a or b;
    layer1_outputs(2774) <= not a;
    layer1_outputs(2775) <= not b;
    layer1_outputs(2776) <= not a;
    layer1_outputs(2777) <= not (a or b);
    layer1_outputs(2778) <= not b or a;
    layer1_outputs(2779) <= not a or b;
    layer1_outputs(2780) <= not (a xor b);
    layer1_outputs(2781) <= not b;
    layer1_outputs(2782) <= not a;
    layer1_outputs(2783) <= not (a xor b);
    layer1_outputs(2784) <= not a;
    layer1_outputs(2785) <= b;
    layer1_outputs(2786) <= not b;
    layer1_outputs(2787) <= a and not b;
    layer1_outputs(2788) <= not b;
    layer1_outputs(2789) <= a and not b;
    layer1_outputs(2790) <= a and b;
    layer1_outputs(2791) <= '0';
    layer1_outputs(2792) <= not (a or b);
    layer1_outputs(2793) <= not (a and b);
    layer1_outputs(2794) <= not a;
    layer1_outputs(2795) <= b;
    layer1_outputs(2796) <= b and not a;
    layer1_outputs(2797) <= b;
    layer1_outputs(2798) <= b;
    layer1_outputs(2799) <= b and not a;
    layer1_outputs(2800) <= a xor b;
    layer1_outputs(2801) <= a;
    layer1_outputs(2802) <= not (a or b);
    layer1_outputs(2803) <= not a;
    layer1_outputs(2804) <= not a;
    layer1_outputs(2805) <= b;
    layer1_outputs(2806) <= '1';
    layer1_outputs(2807) <= a and not b;
    layer1_outputs(2808) <= not (a or b);
    layer1_outputs(2809) <= not (a or b);
    layer1_outputs(2810) <= b and not a;
    layer1_outputs(2811) <= a and not b;
    layer1_outputs(2812) <= a or b;
    layer1_outputs(2813) <= not a;
    layer1_outputs(2814) <= '1';
    layer1_outputs(2815) <= not a;
    layer1_outputs(2816) <= not a;
    layer1_outputs(2817) <= not (a xor b);
    layer1_outputs(2818) <= a and not b;
    layer1_outputs(2819) <= a and not b;
    layer1_outputs(2820) <= a xor b;
    layer1_outputs(2821) <= '0';
    layer1_outputs(2822) <= not b or a;
    layer1_outputs(2823) <= not b or a;
    layer1_outputs(2824) <= a and not b;
    layer1_outputs(2825) <= not (a and b);
    layer1_outputs(2826) <= not (a and b);
    layer1_outputs(2827) <= a and b;
    layer1_outputs(2828) <= a and not b;
    layer1_outputs(2829) <= a and not b;
    layer1_outputs(2830) <= not a;
    layer1_outputs(2831) <= a xor b;
    layer1_outputs(2832) <= a;
    layer1_outputs(2833) <= not (a xor b);
    layer1_outputs(2834) <= a and b;
    layer1_outputs(2835) <= b;
    layer1_outputs(2836) <= not (a or b);
    layer1_outputs(2837) <= a;
    layer1_outputs(2838) <= '1';
    layer1_outputs(2839) <= '0';
    layer1_outputs(2840) <= '0';
    layer1_outputs(2841) <= not (a or b);
    layer1_outputs(2842) <= not (a and b);
    layer1_outputs(2843) <= not b or a;
    layer1_outputs(2844) <= not (a and b);
    layer1_outputs(2845) <= a and b;
    layer1_outputs(2846) <= a and not b;
    layer1_outputs(2847) <= not (a and b);
    layer1_outputs(2848) <= b;
    layer1_outputs(2849) <= a or b;
    layer1_outputs(2850) <= a and b;
    layer1_outputs(2851) <= not (a and b);
    layer1_outputs(2852) <= not (a or b);
    layer1_outputs(2853) <= a;
    layer1_outputs(2854) <= not (a and b);
    layer1_outputs(2855) <= '0';
    layer1_outputs(2856) <= a or b;
    layer1_outputs(2857) <= a;
    layer1_outputs(2858) <= b;
    layer1_outputs(2859) <= a and b;
    layer1_outputs(2860) <= a;
    layer1_outputs(2861) <= not a;
    layer1_outputs(2862) <= '1';
    layer1_outputs(2863) <= a;
    layer1_outputs(2864) <= b;
    layer1_outputs(2865) <= not b or a;
    layer1_outputs(2866) <= b and not a;
    layer1_outputs(2867) <= not (a or b);
    layer1_outputs(2868) <= not (a xor b);
    layer1_outputs(2869) <= b;
    layer1_outputs(2870) <= b;
    layer1_outputs(2871) <= not b or a;
    layer1_outputs(2872) <= not (a or b);
    layer1_outputs(2873) <= not (a and b);
    layer1_outputs(2874) <= not a or b;
    layer1_outputs(2875) <= a xor b;
    layer1_outputs(2876) <= a and b;
    layer1_outputs(2877) <= a or b;
    layer1_outputs(2878) <= a xor b;
    layer1_outputs(2879) <= b and not a;
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= b;
    layer1_outputs(2882) <= b;
    layer1_outputs(2883) <= not b;
    layer1_outputs(2884) <= '1';
    layer1_outputs(2885) <= not a;
    layer1_outputs(2886) <= b;
    layer1_outputs(2887) <= '0';
    layer1_outputs(2888) <= not b or a;
    layer1_outputs(2889) <= not a or b;
    layer1_outputs(2890) <= not b or a;
    layer1_outputs(2891) <= a or b;
    layer1_outputs(2892) <= b and not a;
    layer1_outputs(2893) <= a;
    layer1_outputs(2894) <= not b;
    layer1_outputs(2895) <= not b;
    layer1_outputs(2896) <= not a;
    layer1_outputs(2897) <= b;
    layer1_outputs(2898) <= not a;
    layer1_outputs(2899) <= not (a xor b);
    layer1_outputs(2900) <= a or b;
    layer1_outputs(2901) <= not b;
    layer1_outputs(2902) <= a or b;
    layer1_outputs(2903) <= not (a or b);
    layer1_outputs(2904) <= a or b;
    layer1_outputs(2905) <= a and b;
    layer1_outputs(2906) <= not b;
    layer1_outputs(2907) <= a or b;
    layer1_outputs(2908) <= not a or b;
    layer1_outputs(2909) <= not b;
    layer1_outputs(2910) <= not b or a;
    layer1_outputs(2911) <= b;
    layer1_outputs(2912) <= b and not a;
    layer1_outputs(2913) <= not (a xor b);
    layer1_outputs(2914) <= not a or b;
    layer1_outputs(2915) <= '0';
    layer1_outputs(2916) <= a;
    layer1_outputs(2917) <= not b;
    layer1_outputs(2918) <= not (a and b);
    layer1_outputs(2919) <= not a;
    layer1_outputs(2920) <= a xor b;
    layer1_outputs(2921) <= not a;
    layer1_outputs(2922) <= '0';
    layer1_outputs(2923) <= a and b;
    layer1_outputs(2924) <= not b;
    layer1_outputs(2925) <= not a;
    layer1_outputs(2926) <= not a or b;
    layer1_outputs(2927) <= b;
    layer1_outputs(2928) <= not (a xor b);
    layer1_outputs(2929) <= a;
    layer1_outputs(2930) <= not (a xor b);
    layer1_outputs(2931) <= a or b;
    layer1_outputs(2932) <= a;
    layer1_outputs(2933) <= a or b;
    layer1_outputs(2934) <= not b;
    layer1_outputs(2935) <= b and not a;
    layer1_outputs(2936) <= a and b;
    layer1_outputs(2937) <= b and not a;
    layer1_outputs(2938) <= not b or a;
    layer1_outputs(2939) <= not a;
    layer1_outputs(2940) <= not a;
    layer1_outputs(2941) <= b;
    layer1_outputs(2942) <= a and b;
    layer1_outputs(2943) <= not a;
    layer1_outputs(2944) <= a and not b;
    layer1_outputs(2945) <= not (a and b);
    layer1_outputs(2946) <= a and b;
    layer1_outputs(2947) <= not (a xor b);
    layer1_outputs(2948) <= '0';
    layer1_outputs(2949) <= not b;
    layer1_outputs(2950) <= a and b;
    layer1_outputs(2951) <= not (a xor b);
    layer1_outputs(2952) <= '1';
    layer1_outputs(2953) <= not a or b;
    layer1_outputs(2954) <= not b or a;
    layer1_outputs(2955) <= not b or a;
    layer1_outputs(2956) <= not b or a;
    layer1_outputs(2957) <= a or b;
    layer1_outputs(2958) <= not b;
    layer1_outputs(2959) <= a and not b;
    layer1_outputs(2960) <= '0';
    layer1_outputs(2961) <= not (a and b);
    layer1_outputs(2962) <= b;
    layer1_outputs(2963) <= b;
    layer1_outputs(2964) <= a and not b;
    layer1_outputs(2965) <= not (a or b);
    layer1_outputs(2966) <= b and not a;
    layer1_outputs(2967) <= a xor b;
    layer1_outputs(2968) <= not (a xor b);
    layer1_outputs(2969) <= a or b;
    layer1_outputs(2970) <= '0';
    layer1_outputs(2971) <= b;
    layer1_outputs(2972) <= a and not b;
    layer1_outputs(2973) <= a and not b;
    layer1_outputs(2974) <= a and not b;
    layer1_outputs(2975) <= not a;
    layer1_outputs(2976) <= a;
    layer1_outputs(2977) <= not b;
    layer1_outputs(2978) <= '1';
    layer1_outputs(2979) <= not a;
    layer1_outputs(2980) <= '1';
    layer1_outputs(2981) <= not (a or b);
    layer1_outputs(2982) <= b;
    layer1_outputs(2983) <= a and not b;
    layer1_outputs(2984) <= a xor b;
    layer1_outputs(2985) <= b and not a;
    layer1_outputs(2986) <= '0';
    layer1_outputs(2987) <= not b or a;
    layer1_outputs(2988) <= not a;
    layer1_outputs(2989) <= a and not b;
    layer1_outputs(2990) <= not b;
    layer1_outputs(2991) <= a;
    layer1_outputs(2992) <= not (a and b);
    layer1_outputs(2993) <= '0';
    layer1_outputs(2994) <= '0';
    layer1_outputs(2995) <= not a;
    layer1_outputs(2996) <= '0';
    layer1_outputs(2997) <= not a;
    layer1_outputs(2998) <= not (a or b);
    layer1_outputs(2999) <= a;
    layer1_outputs(3000) <= not a;
    layer1_outputs(3001) <= not a;
    layer1_outputs(3002) <= a;
    layer1_outputs(3003) <= not b;
    layer1_outputs(3004) <= not a;
    layer1_outputs(3005) <= not (a or b);
    layer1_outputs(3006) <= '1';
    layer1_outputs(3007) <= '0';
    layer1_outputs(3008) <= a and not b;
    layer1_outputs(3009) <= a;
    layer1_outputs(3010) <= b;
    layer1_outputs(3011) <= not b;
    layer1_outputs(3012) <= not (a or b);
    layer1_outputs(3013) <= not b or a;
    layer1_outputs(3014) <= b;
    layer1_outputs(3015) <= b and not a;
    layer1_outputs(3016) <= not (a xor b);
    layer1_outputs(3017) <= b;
    layer1_outputs(3018) <= a;
    layer1_outputs(3019) <= not b or a;
    layer1_outputs(3020) <= not b or a;
    layer1_outputs(3021) <= '0';
    layer1_outputs(3022) <= not (a or b);
    layer1_outputs(3023) <= a and not b;
    layer1_outputs(3024) <= b and not a;
    layer1_outputs(3025) <= b;
    layer1_outputs(3026) <= a;
    layer1_outputs(3027) <= not a;
    layer1_outputs(3028) <= not (a or b);
    layer1_outputs(3029) <= not (a xor b);
    layer1_outputs(3030) <= b;
    layer1_outputs(3031) <= '0';
    layer1_outputs(3032) <= not b or a;
    layer1_outputs(3033) <= not (a or b);
    layer1_outputs(3034) <= a and not b;
    layer1_outputs(3035) <= a;
    layer1_outputs(3036) <= not (a and b);
    layer1_outputs(3037) <= not b or a;
    layer1_outputs(3038) <= a and not b;
    layer1_outputs(3039) <= not a or b;
    layer1_outputs(3040) <= a or b;
    layer1_outputs(3041) <= not b or a;
    layer1_outputs(3042) <= not (a and b);
    layer1_outputs(3043) <= not (a or b);
    layer1_outputs(3044) <= not a;
    layer1_outputs(3045) <= '0';
    layer1_outputs(3046) <= not (a or b);
    layer1_outputs(3047) <= a;
    layer1_outputs(3048) <= a or b;
    layer1_outputs(3049) <= not (a and b);
    layer1_outputs(3050) <= a and not b;
    layer1_outputs(3051) <= b;
    layer1_outputs(3052) <= not a or b;
    layer1_outputs(3053) <= a and not b;
    layer1_outputs(3054) <= b and not a;
    layer1_outputs(3055) <= b and not a;
    layer1_outputs(3056) <= not a;
    layer1_outputs(3057) <= not a;
    layer1_outputs(3058) <= not (a or b);
    layer1_outputs(3059) <= a or b;
    layer1_outputs(3060) <= not (a or b);
    layer1_outputs(3061) <= not (a or b);
    layer1_outputs(3062) <= not b or a;
    layer1_outputs(3063) <= not (a or b);
    layer1_outputs(3064) <= a and b;
    layer1_outputs(3065) <= not (a and b);
    layer1_outputs(3066) <= '1';
    layer1_outputs(3067) <= b and not a;
    layer1_outputs(3068) <= '1';
    layer1_outputs(3069) <= b;
    layer1_outputs(3070) <= b;
    layer1_outputs(3071) <= not a or b;
    layer1_outputs(3072) <= not a;
    layer1_outputs(3073) <= a or b;
    layer1_outputs(3074) <= not a;
    layer1_outputs(3075) <= '0';
    layer1_outputs(3076) <= b;
    layer1_outputs(3077) <= b;
    layer1_outputs(3078) <= not b or a;
    layer1_outputs(3079) <= a and b;
    layer1_outputs(3080) <= not a or b;
    layer1_outputs(3081) <= b and not a;
    layer1_outputs(3082) <= a;
    layer1_outputs(3083) <= not a;
    layer1_outputs(3084) <= a xor b;
    layer1_outputs(3085) <= not a or b;
    layer1_outputs(3086) <= not (a or b);
    layer1_outputs(3087) <= not (a and b);
    layer1_outputs(3088) <= not a;
    layer1_outputs(3089) <= a and b;
    layer1_outputs(3090) <= not a or b;
    layer1_outputs(3091) <= b;
    layer1_outputs(3092) <= not (a and b);
    layer1_outputs(3093) <= not b;
    layer1_outputs(3094) <= a and not b;
    layer1_outputs(3095) <= a;
    layer1_outputs(3096) <= b and not a;
    layer1_outputs(3097) <= not (a or b);
    layer1_outputs(3098) <= not (a and b);
    layer1_outputs(3099) <= a and b;
    layer1_outputs(3100) <= b and not a;
    layer1_outputs(3101) <= '0';
    layer1_outputs(3102) <= not (a xor b);
    layer1_outputs(3103) <= not b or a;
    layer1_outputs(3104) <= a xor b;
    layer1_outputs(3105) <= a or b;
    layer1_outputs(3106) <= not (a xor b);
    layer1_outputs(3107) <= a and b;
    layer1_outputs(3108) <= a and b;
    layer1_outputs(3109) <= a;
    layer1_outputs(3110) <= a;
    layer1_outputs(3111) <= not a or b;
    layer1_outputs(3112) <= a xor b;
    layer1_outputs(3113) <= a and not b;
    layer1_outputs(3114) <= a and b;
    layer1_outputs(3115) <= b and not a;
    layer1_outputs(3116) <= '0';
    layer1_outputs(3117) <= a or b;
    layer1_outputs(3118) <= not (a and b);
    layer1_outputs(3119) <= not (a and b);
    layer1_outputs(3120) <= b;
    layer1_outputs(3121) <= a;
    layer1_outputs(3122) <= not b;
    layer1_outputs(3123) <= not (a or b);
    layer1_outputs(3124) <= not a;
    layer1_outputs(3125) <= not (a and b);
    layer1_outputs(3126) <= b;
    layer1_outputs(3127) <= b;
    layer1_outputs(3128) <= not (a xor b);
    layer1_outputs(3129) <= a;
    layer1_outputs(3130) <= not (a and b);
    layer1_outputs(3131) <= b;
    layer1_outputs(3132) <= '1';
    layer1_outputs(3133) <= not (a xor b);
    layer1_outputs(3134) <= a or b;
    layer1_outputs(3135) <= b and not a;
    layer1_outputs(3136) <= not (a xor b);
    layer1_outputs(3137) <= a xor b;
    layer1_outputs(3138) <= a and not b;
    layer1_outputs(3139) <= not a;
    layer1_outputs(3140) <= a or b;
    layer1_outputs(3141) <= '0';
    layer1_outputs(3142) <= not a;
    layer1_outputs(3143) <= a and b;
    layer1_outputs(3144) <= a and not b;
    layer1_outputs(3145) <= a;
    layer1_outputs(3146) <= a xor b;
    layer1_outputs(3147) <= '1';
    layer1_outputs(3148) <= a and not b;
    layer1_outputs(3149) <= b;
    layer1_outputs(3150) <= a;
    layer1_outputs(3151) <= not a or b;
    layer1_outputs(3152) <= a xor b;
    layer1_outputs(3153) <= a;
    layer1_outputs(3154) <= not (a and b);
    layer1_outputs(3155) <= '1';
    layer1_outputs(3156) <= a;
    layer1_outputs(3157) <= b and not a;
    layer1_outputs(3158) <= not b or a;
    layer1_outputs(3159) <= not (a xor b);
    layer1_outputs(3160) <= not a;
    layer1_outputs(3161) <= not b or a;
    layer1_outputs(3162) <= a or b;
    layer1_outputs(3163) <= not (a or b);
    layer1_outputs(3164) <= not (a xor b);
    layer1_outputs(3165) <= not b or a;
    layer1_outputs(3166) <= a and not b;
    layer1_outputs(3167) <= a or b;
    layer1_outputs(3168) <= a and b;
    layer1_outputs(3169) <= not b;
    layer1_outputs(3170) <= not b or a;
    layer1_outputs(3171) <= '1';
    layer1_outputs(3172) <= '0';
    layer1_outputs(3173) <= not a or b;
    layer1_outputs(3174) <= a and b;
    layer1_outputs(3175) <= not a or b;
    layer1_outputs(3176) <= a;
    layer1_outputs(3177) <= not (a xor b);
    layer1_outputs(3178) <= a;
    layer1_outputs(3179) <= not b;
    layer1_outputs(3180) <= a xor b;
    layer1_outputs(3181) <= a and not b;
    layer1_outputs(3182) <= not (a or b);
    layer1_outputs(3183) <= not (a and b);
    layer1_outputs(3184) <= not b;
    layer1_outputs(3185) <= not (a xor b);
    layer1_outputs(3186) <= not (a and b);
    layer1_outputs(3187) <= b and not a;
    layer1_outputs(3188) <= not (a and b);
    layer1_outputs(3189) <= b and not a;
    layer1_outputs(3190) <= not (a or b);
    layer1_outputs(3191) <= a xor b;
    layer1_outputs(3192) <= b;
    layer1_outputs(3193) <= not a or b;
    layer1_outputs(3194) <= b;
    layer1_outputs(3195) <= a;
    layer1_outputs(3196) <= b;
    layer1_outputs(3197) <= not (a or b);
    layer1_outputs(3198) <= b and not a;
    layer1_outputs(3199) <= not b or a;
    layer1_outputs(3200) <= not a or b;
    layer1_outputs(3201) <= a and not b;
    layer1_outputs(3202) <= a;
    layer1_outputs(3203) <= not a;
    layer1_outputs(3204) <= a;
    layer1_outputs(3205) <= b;
    layer1_outputs(3206) <= not b or a;
    layer1_outputs(3207) <= not a or b;
    layer1_outputs(3208) <= a and b;
    layer1_outputs(3209) <= not b;
    layer1_outputs(3210) <= not a;
    layer1_outputs(3211) <= a;
    layer1_outputs(3212) <= a and not b;
    layer1_outputs(3213) <= not b or a;
    layer1_outputs(3214) <= not (a or b);
    layer1_outputs(3215) <= a and b;
    layer1_outputs(3216) <= not b or a;
    layer1_outputs(3217) <= a;
    layer1_outputs(3218) <= b and not a;
    layer1_outputs(3219) <= b;
    layer1_outputs(3220) <= b;
    layer1_outputs(3221) <= b;
    layer1_outputs(3222) <= not b or a;
    layer1_outputs(3223) <= not b or a;
    layer1_outputs(3224) <= a xor b;
    layer1_outputs(3225) <= a;
    layer1_outputs(3226) <= not a or b;
    layer1_outputs(3227) <= not b or a;
    layer1_outputs(3228) <= a or b;
    layer1_outputs(3229) <= a;
    layer1_outputs(3230) <= not b or a;
    layer1_outputs(3231) <= b;
    layer1_outputs(3232) <= not a;
    layer1_outputs(3233) <= b;
    layer1_outputs(3234) <= a and not b;
    layer1_outputs(3235) <= b and not a;
    layer1_outputs(3236) <= '0';
    layer1_outputs(3237) <= not b or a;
    layer1_outputs(3238) <= not b;
    layer1_outputs(3239) <= not (a and b);
    layer1_outputs(3240) <= a and not b;
    layer1_outputs(3241) <= not b;
    layer1_outputs(3242) <= not (a or b);
    layer1_outputs(3243) <= '0';
    layer1_outputs(3244) <= b;
    layer1_outputs(3245) <= '0';
    layer1_outputs(3246) <= a;
    layer1_outputs(3247) <= a and not b;
    layer1_outputs(3248) <= not (a or b);
    layer1_outputs(3249) <= a and b;
    layer1_outputs(3250) <= not a or b;
    layer1_outputs(3251) <= not (a xor b);
    layer1_outputs(3252) <= a and not b;
    layer1_outputs(3253) <= not (a and b);
    layer1_outputs(3254) <= a and not b;
    layer1_outputs(3255) <= not b or a;
    layer1_outputs(3256) <= a xor b;
    layer1_outputs(3257) <= a and not b;
    layer1_outputs(3258) <= b;
    layer1_outputs(3259) <= not b or a;
    layer1_outputs(3260) <= not (a and b);
    layer1_outputs(3261) <= a and not b;
    layer1_outputs(3262) <= not (a and b);
    layer1_outputs(3263) <= a and not b;
    layer1_outputs(3264) <= a and not b;
    layer1_outputs(3265) <= not (a and b);
    layer1_outputs(3266) <= a and b;
    layer1_outputs(3267) <= not a;
    layer1_outputs(3268) <= not (a xor b);
    layer1_outputs(3269) <= not b or a;
    layer1_outputs(3270) <= a xor b;
    layer1_outputs(3271) <= '1';
    layer1_outputs(3272) <= not (a or b);
    layer1_outputs(3273) <= b and not a;
    layer1_outputs(3274) <= a and not b;
    layer1_outputs(3275) <= not b;
    layer1_outputs(3276) <= a or b;
    layer1_outputs(3277) <= a and b;
    layer1_outputs(3278) <= a and b;
    layer1_outputs(3279) <= a and b;
    layer1_outputs(3280) <= '0';
    layer1_outputs(3281) <= a xor b;
    layer1_outputs(3282) <= a or b;
    layer1_outputs(3283) <= a and b;
    layer1_outputs(3284) <= a and not b;
    layer1_outputs(3285) <= not (a and b);
    layer1_outputs(3286) <= a and b;
    layer1_outputs(3287) <= b and not a;
    layer1_outputs(3288) <= a;
    layer1_outputs(3289) <= a or b;
    layer1_outputs(3290) <= a or b;
    layer1_outputs(3291) <= not b;
    layer1_outputs(3292) <= '0';
    layer1_outputs(3293) <= not a;
    layer1_outputs(3294) <= not b or a;
    layer1_outputs(3295) <= not (a xor b);
    layer1_outputs(3296) <= b;
    layer1_outputs(3297) <= a;
    layer1_outputs(3298) <= not b;
    layer1_outputs(3299) <= a and b;
    layer1_outputs(3300) <= not (a or b);
    layer1_outputs(3301) <= not a;
    layer1_outputs(3302) <= not (a and b);
    layer1_outputs(3303) <= not b or a;
    layer1_outputs(3304) <= a or b;
    layer1_outputs(3305) <= '0';
    layer1_outputs(3306) <= not b or a;
    layer1_outputs(3307) <= a and not b;
    layer1_outputs(3308) <= b and not a;
    layer1_outputs(3309) <= a and b;
    layer1_outputs(3310) <= not b or a;
    layer1_outputs(3311) <= not b;
    layer1_outputs(3312) <= a;
    layer1_outputs(3313) <= not b or a;
    layer1_outputs(3314) <= '0';
    layer1_outputs(3315) <= not a;
    layer1_outputs(3316) <= a;
    layer1_outputs(3317) <= not a;
    layer1_outputs(3318) <= a;
    layer1_outputs(3319) <= a;
    layer1_outputs(3320) <= not (a or b);
    layer1_outputs(3321) <= a and not b;
    layer1_outputs(3322) <= a and not b;
    layer1_outputs(3323) <= '1';
    layer1_outputs(3324) <= a;
    layer1_outputs(3325) <= not b;
    layer1_outputs(3326) <= '0';
    layer1_outputs(3327) <= not b or a;
    layer1_outputs(3328) <= '0';
    layer1_outputs(3329) <= a;
    layer1_outputs(3330) <= b;
    layer1_outputs(3331) <= not b or a;
    layer1_outputs(3332) <= a;
    layer1_outputs(3333) <= not a or b;
    layer1_outputs(3334) <= b;
    layer1_outputs(3335) <= b;
    layer1_outputs(3336) <= not (a and b);
    layer1_outputs(3337) <= a;
    layer1_outputs(3338) <= a and not b;
    layer1_outputs(3339) <= b and not a;
    layer1_outputs(3340) <= a and b;
    layer1_outputs(3341) <= a or b;
    layer1_outputs(3342) <= a xor b;
    layer1_outputs(3343) <= not a or b;
    layer1_outputs(3344) <= b;
    layer1_outputs(3345) <= not (a and b);
    layer1_outputs(3346) <= not a;
    layer1_outputs(3347) <= not a or b;
    layer1_outputs(3348) <= not (a or b);
    layer1_outputs(3349) <= not (a and b);
    layer1_outputs(3350) <= '1';
    layer1_outputs(3351) <= not b;
    layer1_outputs(3352) <= not a or b;
    layer1_outputs(3353) <= a and not b;
    layer1_outputs(3354) <= a xor b;
    layer1_outputs(3355) <= a xor b;
    layer1_outputs(3356) <= a;
    layer1_outputs(3357) <= a or b;
    layer1_outputs(3358) <= not b or a;
    layer1_outputs(3359) <= not (a or b);
    layer1_outputs(3360) <= a and b;
    layer1_outputs(3361) <= not b;
    layer1_outputs(3362) <= b and not a;
    layer1_outputs(3363) <= a or b;
    layer1_outputs(3364) <= not (a or b);
    layer1_outputs(3365) <= a or b;
    layer1_outputs(3366) <= not b or a;
    layer1_outputs(3367) <= a and b;
    layer1_outputs(3368) <= not b or a;
    layer1_outputs(3369) <= a or b;
    layer1_outputs(3370) <= '1';
    layer1_outputs(3371) <= a and b;
    layer1_outputs(3372) <= not a;
    layer1_outputs(3373) <= a or b;
    layer1_outputs(3374) <= b;
    layer1_outputs(3375) <= a or b;
    layer1_outputs(3376) <= not b;
    layer1_outputs(3377) <= a or b;
    layer1_outputs(3378) <= not b or a;
    layer1_outputs(3379) <= not a;
    layer1_outputs(3380) <= not b or a;
    layer1_outputs(3381) <= a and not b;
    layer1_outputs(3382) <= a;
    layer1_outputs(3383) <= not a;
    layer1_outputs(3384) <= a and not b;
    layer1_outputs(3385) <= '0';
    layer1_outputs(3386) <= a and b;
    layer1_outputs(3387) <= a;
    layer1_outputs(3388) <= a;
    layer1_outputs(3389) <= a xor b;
    layer1_outputs(3390) <= not b;
    layer1_outputs(3391) <= a;
    layer1_outputs(3392) <= not (a or b);
    layer1_outputs(3393) <= not (a and b);
    layer1_outputs(3394) <= b;
    layer1_outputs(3395) <= a;
    layer1_outputs(3396) <= '1';
    layer1_outputs(3397) <= not a;
    layer1_outputs(3398) <= '0';
    layer1_outputs(3399) <= a and b;
    layer1_outputs(3400) <= not (a and b);
    layer1_outputs(3401) <= not a;
    layer1_outputs(3402) <= not b or a;
    layer1_outputs(3403) <= not b or a;
    layer1_outputs(3404) <= b;
    layer1_outputs(3405) <= not (a xor b);
    layer1_outputs(3406) <= not b;
    layer1_outputs(3407) <= not a or b;
    layer1_outputs(3408) <= not b;
    layer1_outputs(3409) <= not a or b;
    layer1_outputs(3410) <= not a or b;
    layer1_outputs(3411) <= '0';
    layer1_outputs(3412) <= not (a or b);
    layer1_outputs(3413) <= not b;
    layer1_outputs(3414) <= '1';
    layer1_outputs(3415) <= '1';
    layer1_outputs(3416) <= not b;
    layer1_outputs(3417) <= a;
    layer1_outputs(3418) <= a and b;
    layer1_outputs(3419) <= a or b;
    layer1_outputs(3420) <= not b or a;
    layer1_outputs(3421) <= a and b;
    layer1_outputs(3422) <= not (a xor b);
    layer1_outputs(3423) <= a and b;
    layer1_outputs(3424) <= not b;
    layer1_outputs(3425) <= a and not b;
    layer1_outputs(3426) <= a or b;
    layer1_outputs(3427) <= not (a or b);
    layer1_outputs(3428) <= not a;
    layer1_outputs(3429) <= a or b;
    layer1_outputs(3430) <= not (a or b);
    layer1_outputs(3431) <= a and not b;
    layer1_outputs(3432) <= not b;
    layer1_outputs(3433) <= a and not b;
    layer1_outputs(3434) <= a and b;
    layer1_outputs(3435) <= not (a xor b);
    layer1_outputs(3436) <= a or b;
    layer1_outputs(3437) <= not (a and b);
    layer1_outputs(3438) <= not (a and b);
    layer1_outputs(3439) <= not (a or b);
    layer1_outputs(3440) <= b;
    layer1_outputs(3441) <= '0';
    layer1_outputs(3442) <= b and not a;
    layer1_outputs(3443) <= not a;
    layer1_outputs(3444) <= not (a or b);
    layer1_outputs(3445) <= '1';
    layer1_outputs(3446) <= not b;
    layer1_outputs(3447) <= not (a and b);
    layer1_outputs(3448) <= not b or a;
    layer1_outputs(3449) <= not a or b;
    layer1_outputs(3450) <= not (a and b);
    layer1_outputs(3451) <= not (a or b);
    layer1_outputs(3452) <= a and not b;
    layer1_outputs(3453) <= not b or a;
    layer1_outputs(3454) <= a and b;
    layer1_outputs(3455) <= '0';
    layer1_outputs(3456) <= not (a or b);
    layer1_outputs(3457) <= a;
    layer1_outputs(3458) <= a and b;
    layer1_outputs(3459) <= a or b;
    layer1_outputs(3460) <= b and not a;
    layer1_outputs(3461) <= not (a and b);
    layer1_outputs(3462) <= a and b;
    layer1_outputs(3463) <= b and not a;
    layer1_outputs(3464) <= not (a xor b);
    layer1_outputs(3465) <= b and not a;
    layer1_outputs(3466) <= not (a or b);
    layer1_outputs(3467) <= a and b;
    layer1_outputs(3468) <= not b or a;
    layer1_outputs(3469) <= a;
    layer1_outputs(3470) <= not b or a;
    layer1_outputs(3471) <= a or b;
    layer1_outputs(3472) <= b and not a;
    layer1_outputs(3473) <= b;
    layer1_outputs(3474) <= not b;
    layer1_outputs(3475) <= not (a or b);
    layer1_outputs(3476) <= '1';
    layer1_outputs(3477) <= b;
    layer1_outputs(3478) <= a or b;
    layer1_outputs(3479) <= not b;
    layer1_outputs(3480) <= not (a or b);
    layer1_outputs(3481) <= not a or b;
    layer1_outputs(3482) <= a;
    layer1_outputs(3483) <= not (a and b);
    layer1_outputs(3484) <= b;
    layer1_outputs(3485) <= not b;
    layer1_outputs(3486) <= not b;
    layer1_outputs(3487) <= not (a and b);
    layer1_outputs(3488) <= not (a or b);
    layer1_outputs(3489) <= b;
    layer1_outputs(3490) <= not a;
    layer1_outputs(3491) <= not (a or b);
    layer1_outputs(3492) <= b;
    layer1_outputs(3493) <= not a or b;
    layer1_outputs(3494) <= not (a and b);
    layer1_outputs(3495) <= not b;
    layer1_outputs(3496) <= not a or b;
    layer1_outputs(3497) <= b;
    layer1_outputs(3498) <= b;
    layer1_outputs(3499) <= a and b;
    layer1_outputs(3500) <= not a or b;
    layer1_outputs(3501) <= a;
    layer1_outputs(3502) <= not b;
    layer1_outputs(3503) <= not (a and b);
    layer1_outputs(3504) <= a and not b;
    layer1_outputs(3505) <= b and not a;
    layer1_outputs(3506) <= a;
    layer1_outputs(3507) <= a;
    layer1_outputs(3508) <= a or b;
    layer1_outputs(3509) <= '0';
    layer1_outputs(3510) <= a and b;
    layer1_outputs(3511) <= not a;
    layer1_outputs(3512) <= not (a or b);
    layer1_outputs(3513) <= b;
    layer1_outputs(3514) <= b;
    layer1_outputs(3515) <= not a;
    layer1_outputs(3516) <= not b;
    layer1_outputs(3517) <= not (a or b);
    layer1_outputs(3518) <= not a or b;
    layer1_outputs(3519) <= not a or b;
    layer1_outputs(3520) <= not (a xor b);
    layer1_outputs(3521) <= not a or b;
    layer1_outputs(3522) <= not (a and b);
    layer1_outputs(3523) <= not (a or b);
    layer1_outputs(3524) <= b;
    layer1_outputs(3525) <= a and b;
    layer1_outputs(3526) <= a xor b;
    layer1_outputs(3527) <= not b;
    layer1_outputs(3528) <= a or b;
    layer1_outputs(3529) <= b and not a;
    layer1_outputs(3530) <= b and not a;
    layer1_outputs(3531) <= '0';
    layer1_outputs(3532) <= not b;
    layer1_outputs(3533) <= a and b;
    layer1_outputs(3534) <= not b;
    layer1_outputs(3535) <= a and not b;
    layer1_outputs(3536) <= not a;
    layer1_outputs(3537) <= '1';
    layer1_outputs(3538) <= not (a xor b);
    layer1_outputs(3539) <= not (a or b);
    layer1_outputs(3540) <= a and not b;
    layer1_outputs(3541) <= b and not a;
    layer1_outputs(3542) <= not a or b;
    layer1_outputs(3543) <= a or b;
    layer1_outputs(3544) <= not b or a;
    layer1_outputs(3545) <= a;
    layer1_outputs(3546) <= not b;
    layer1_outputs(3547) <= not a;
    layer1_outputs(3548) <= a;
    layer1_outputs(3549) <= b;
    layer1_outputs(3550) <= a;
    layer1_outputs(3551) <= '1';
    layer1_outputs(3552) <= not (a and b);
    layer1_outputs(3553) <= not a;
    layer1_outputs(3554) <= a or b;
    layer1_outputs(3555) <= not b or a;
    layer1_outputs(3556) <= b;
    layer1_outputs(3557) <= not a;
    layer1_outputs(3558) <= not b or a;
    layer1_outputs(3559) <= a;
    layer1_outputs(3560) <= a or b;
    layer1_outputs(3561) <= not (a and b);
    layer1_outputs(3562) <= b and not a;
    layer1_outputs(3563) <= b and not a;
    layer1_outputs(3564) <= not b or a;
    layer1_outputs(3565) <= b;
    layer1_outputs(3566) <= a and not b;
    layer1_outputs(3567) <= not (a xor b);
    layer1_outputs(3568) <= '1';
    layer1_outputs(3569) <= not (a and b);
    layer1_outputs(3570) <= a or b;
    layer1_outputs(3571) <= a or b;
    layer1_outputs(3572) <= a and b;
    layer1_outputs(3573) <= a and b;
    layer1_outputs(3574) <= b and not a;
    layer1_outputs(3575) <= not a;
    layer1_outputs(3576) <= a and b;
    layer1_outputs(3577) <= not a or b;
    layer1_outputs(3578) <= b;
    layer1_outputs(3579) <= not b;
    layer1_outputs(3580) <= a;
    layer1_outputs(3581) <= b and not a;
    layer1_outputs(3582) <= not (a or b);
    layer1_outputs(3583) <= a;
    layer1_outputs(3584) <= a and b;
    layer1_outputs(3585) <= a and not b;
    layer1_outputs(3586) <= a and not b;
    layer1_outputs(3587) <= not a;
    layer1_outputs(3588) <= not (a or b);
    layer1_outputs(3589) <= not b;
    layer1_outputs(3590) <= a;
    layer1_outputs(3591) <= not (a and b);
    layer1_outputs(3592) <= not a;
    layer1_outputs(3593) <= b and not a;
    layer1_outputs(3594) <= not (a and b);
    layer1_outputs(3595) <= not a or b;
    layer1_outputs(3596) <= b and not a;
    layer1_outputs(3597) <= not (a or b);
    layer1_outputs(3598) <= a;
    layer1_outputs(3599) <= not b;
    layer1_outputs(3600) <= a and not b;
    layer1_outputs(3601) <= not (a and b);
    layer1_outputs(3602) <= b;
    layer1_outputs(3603) <= b;
    layer1_outputs(3604) <= not (a or b);
    layer1_outputs(3605) <= not a or b;
    layer1_outputs(3606) <= not b or a;
    layer1_outputs(3607) <= not b;
    layer1_outputs(3608) <= a and not b;
    layer1_outputs(3609) <= a;
    layer1_outputs(3610) <= not (a and b);
    layer1_outputs(3611) <= a and not b;
    layer1_outputs(3612) <= a and b;
    layer1_outputs(3613) <= not a;
    layer1_outputs(3614) <= '0';
    layer1_outputs(3615) <= not b or a;
    layer1_outputs(3616) <= b and not a;
    layer1_outputs(3617) <= a and b;
    layer1_outputs(3618) <= not (a or b);
    layer1_outputs(3619) <= b and not a;
    layer1_outputs(3620) <= '0';
    layer1_outputs(3621) <= a;
    layer1_outputs(3622) <= a xor b;
    layer1_outputs(3623) <= not b or a;
    layer1_outputs(3624) <= b and not a;
    layer1_outputs(3625) <= b and not a;
    layer1_outputs(3626) <= not (a or b);
    layer1_outputs(3627) <= a and b;
    layer1_outputs(3628) <= '1';
    layer1_outputs(3629) <= not b or a;
    layer1_outputs(3630) <= a or b;
    layer1_outputs(3631) <= a and b;
    layer1_outputs(3632) <= b;
    layer1_outputs(3633) <= a and b;
    layer1_outputs(3634) <= a and b;
    layer1_outputs(3635) <= not (a xor b);
    layer1_outputs(3636) <= '1';
    layer1_outputs(3637) <= not b;
    layer1_outputs(3638) <= '0';
    layer1_outputs(3639) <= not a or b;
    layer1_outputs(3640) <= not b;
    layer1_outputs(3641) <= a and b;
    layer1_outputs(3642) <= not b or a;
    layer1_outputs(3643) <= a and b;
    layer1_outputs(3644) <= a or b;
    layer1_outputs(3645) <= a or b;
    layer1_outputs(3646) <= not b;
    layer1_outputs(3647) <= not b;
    layer1_outputs(3648) <= a and not b;
    layer1_outputs(3649) <= a or b;
    layer1_outputs(3650) <= '1';
    layer1_outputs(3651) <= a;
    layer1_outputs(3652) <= a;
    layer1_outputs(3653) <= not b;
    layer1_outputs(3654) <= not (a and b);
    layer1_outputs(3655) <= not a or b;
    layer1_outputs(3656) <= not (a and b);
    layer1_outputs(3657) <= not b or a;
    layer1_outputs(3658) <= not (a xor b);
    layer1_outputs(3659) <= a;
    layer1_outputs(3660) <= b and not a;
    layer1_outputs(3661) <= not (a or b);
    layer1_outputs(3662) <= not b;
    layer1_outputs(3663) <= a and not b;
    layer1_outputs(3664) <= not a;
    layer1_outputs(3665) <= b and not a;
    layer1_outputs(3666) <= not a or b;
    layer1_outputs(3667) <= not a;
    layer1_outputs(3668) <= a and b;
    layer1_outputs(3669) <= a and not b;
    layer1_outputs(3670) <= a xor b;
    layer1_outputs(3671) <= not a;
    layer1_outputs(3672) <= not a;
    layer1_outputs(3673) <= b;
    layer1_outputs(3674) <= not (a xor b);
    layer1_outputs(3675) <= b and not a;
    layer1_outputs(3676) <= a or b;
    layer1_outputs(3677) <= '1';
    layer1_outputs(3678) <= not (a xor b);
    layer1_outputs(3679) <= not b;
    layer1_outputs(3680) <= a and b;
    layer1_outputs(3681) <= a xor b;
    layer1_outputs(3682) <= a and b;
    layer1_outputs(3683) <= a and not b;
    layer1_outputs(3684) <= a and b;
    layer1_outputs(3685) <= not b or a;
    layer1_outputs(3686) <= b and not a;
    layer1_outputs(3687) <= not a or b;
    layer1_outputs(3688) <= a and not b;
    layer1_outputs(3689) <= b and not a;
    layer1_outputs(3690) <= not (a xor b);
    layer1_outputs(3691) <= not (a and b);
    layer1_outputs(3692) <= '1';
    layer1_outputs(3693) <= a;
    layer1_outputs(3694) <= not b or a;
    layer1_outputs(3695) <= a xor b;
    layer1_outputs(3696) <= a and b;
    layer1_outputs(3697) <= not (a or b);
    layer1_outputs(3698) <= b;
    layer1_outputs(3699) <= a;
    layer1_outputs(3700) <= not (a or b);
    layer1_outputs(3701) <= a and not b;
    layer1_outputs(3702) <= a and b;
    layer1_outputs(3703) <= b;
    layer1_outputs(3704) <= b and not a;
    layer1_outputs(3705) <= not a;
    layer1_outputs(3706) <= a;
    layer1_outputs(3707) <= not (a xor b);
    layer1_outputs(3708) <= a and b;
    layer1_outputs(3709) <= not a;
    layer1_outputs(3710) <= not (a and b);
    layer1_outputs(3711) <= not a or b;
    layer1_outputs(3712) <= not a or b;
    layer1_outputs(3713) <= not b;
    layer1_outputs(3714) <= a;
    layer1_outputs(3715) <= a and not b;
    layer1_outputs(3716) <= not a;
    layer1_outputs(3717) <= not b or a;
    layer1_outputs(3718) <= a;
    layer1_outputs(3719) <= not (a and b);
    layer1_outputs(3720) <= not a;
    layer1_outputs(3721) <= not (a and b);
    layer1_outputs(3722) <= a and b;
    layer1_outputs(3723) <= not (a or b);
    layer1_outputs(3724) <= not a;
    layer1_outputs(3725) <= a;
    layer1_outputs(3726) <= a;
    layer1_outputs(3727) <= b;
    layer1_outputs(3728) <= a or b;
    layer1_outputs(3729) <= not (a and b);
    layer1_outputs(3730) <= '1';
    layer1_outputs(3731) <= b;
    layer1_outputs(3732) <= not a;
    layer1_outputs(3733) <= not (a or b);
    layer1_outputs(3734) <= a or b;
    layer1_outputs(3735) <= not b or a;
    layer1_outputs(3736) <= a and b;
    layer1_outputs(3737) <= not b or a;
    layer1_outputs(3738) <= a xor b;
    layer1_outputs(3739) <= b;
    layer1_outputs(3740) <= not (a or b);
    layer1_outputs(3741) <= b and not a;
    layer1_outputs(3742) <= not b or a;
    layer1_outputs(3743) <= a xor b;
    layer1_outputs(3744) <= not (a or b);
    layer1_outputs(3745) <= not (a and b);
    layer1_outputs(3746) <= a xor b;
    layer1_outputs(3747) <= not a;
    layer1_outputs(3748) <= not a;
    layer1_outputs(3749) <= a;
    layer1_outputs(3750) <= a;
    layer1_outputs(3751) <= a or b;
    layer1_outputs(3752) <= not a;
    layer1_outputs(3753) <= a;
    layer1_outputs(3754) <= not b;
    layer1_outputs(3755) <= not a or b;
    layer1_outputs(3756) <= '0';
    layer1_outputs(3757) <= not (a and b);
    layer1_outputs(3758) <= b;
    layer1_outputs(3759) <= not (a or b);
    layer1_outputs(3760) <= b;
    layer1_outputs(3761) <= a or b;
    layer1_outputs(3762) <= b and not a;
    layer1_outputs(3763) <= a or b;
    layer1_outputs(3764) <= '0';
    layer1_outputs(3765) <= not (a xor b);
    layer1_outputs(3766) <= not b;
    layer1_outputs(3767) <= a and not b;
    layer1_outputs(3768) <= a;
    layer1_outputs(3769) <= a xor b;
    layer1_outputs(3770) <= b and not a;
    layer1_outputs(3771) <= a or b;
    layer1_outputs(3772) <= not b;
    layer1_outputs(3773) <= not (a and b);
    layer1_outputs(3774) <= not a or b;
    layer1_outputs(3775) <= '1';
    layer1_outputs(3776) <= a or b;
    layer1_outputs(3777) <= '1';
    layer1_outputs(3778) <= b and not a;
    layer1_outputs(3779) <= b;
    layer1_outputs(3780) <= not a or b;
    layer1_outputs(3781) <= not b;
    layer1_outputs(3782) <= a xor b;
    layer1_outputs(3783) <= a;
    layer1_outputs(3784) <= a;
    layer1_outputs(3785) <= not b or a;
    layer1_outputs(3786) <= a or b;
    layer1_outputs(3787) <= a and b;
    layer1_outputs(3788) <= not a;
    layer1_outputs(3789) <= b and not a;
    layer1_outputs(3790) <= a or b;
    layer1_outputs(3791) <= a and not b;
    layer1_outputs(3792) <= not a;
    layer1_outputs(3793) <= a xor b;
    layer1_outputs(3794) <= not b or a;
    layer1_outputs(3795) <= '0';
    layer1_outputs(3796) <= not a;
    layer1_outputs(3797) <= not (a and b);
    layer1_outputs(3798) <= '1';
    layer1_outputs(3799) <= b and not a;
    layer1_outputs(3800) <= b;
    layer1_outputs(3801) <= a and not b;
    layer1_outputs(3802) <= b and not a;
    layer1_outputs(3803) <= not a;
    layer1_outputs(3804) <= a;
    layer1_outputs(3805) <= not b or a;
    layer1_outputs(3806) <= not a or b;
    layer1_outputs(3807) <= not b;
    layer1_outputs(3808) <= not (a and b);
    layer1_outputs(3809) <= '1';
    layer1_outputs(3810) <= a;
    layer1_outputs(3811) <= not (a and b);
    layer1_outputs(3812) <= b and not a;
    layer1_outputs(3813) <= not b or a;
    layer1_outputs(3814) <= not b;
    layer1_outputs(3815) <= not (a xor b);
    layer1_outputs(3816) <= not b;
    layer1_outputs(3817) <= b;
    layer1_outputs(3818) <= b;
    layer1_outputs(3819) <= not a or b;
    layer1_outputs(3820) <= not (a xor b);
    layer1_outputs(3821) <= not (a xor b);
    layer1_outputs(3822) <= not a or b;
    layer1_outputs(3823) <= not (a or b);
    layer1_outputs(3824) <= a and not b;
    layer1_outputs(3825) <= not b;
    layer1_outputs(3826) <= not b;
    layer1_outputs(3827) <= a;
    layer1_outputs(3828) <= a;
    layer1_outputs(3829) <= a;
    layer1_outputs(3830) <= b and not a;
    layer1_outputs(3831) <= a and b;
    layer1_outputs(3832) <= not b or a;
    layer1_outputs(3833) <= '0';
    layer1_outputs(3834) <= not a;
    layer1_outputs(3835) <= a and not b;
    layer1_outputs(3836) <= b;
    layer1_outputs(3837) <= a xor b;
    layer1_outputs(3838) <= '1';
    layer1_outputs(3839) <= a;
    layer1_outputs(3840) <= b;
    layer1_outputs(3841) <= not b or a;
    layer1_outputs(3842) <= not a or b;
    layer1_outputs(3843) <= b;
    layer1_outputs(3844) <= not (a or b);
    layer1_outputs(3845) <= not a or b;
    layer1_outputs(3846) <= '1';
    layer1_outputs(3847) <= not b;
    layer1_outputs(3848) <= not b or a;
    layer1_outputs(3849) <= not a or b;
    layer1_outputs(3850) <= b and not a;
    layer1_outputs(3851) <= a and not b;
    layer1_outputs(3852) <= a and not b;
    layer1_outputs(3853) <= not (a and b);
    layer1_outputs(3854) <= not a;
    layer1_outputs(3855) <= a;
    layer1_outputs(3856) <= a and not b;
    layer1_outputs(3857) <= a or b;
    layer1_outputs(3858) <= b and not a;
    layer1_outputs(3859) <= a;
    layer1_outputs(3860) <= a or b;
    layer1_outputs(3861) <= b;
    layer1_outputs(3862) <= not b;
    layer1_outputs(3863) <= not a or b;
    layer1_outputs(3864) <= a xor b;
    layer1_outputs(3865) <= not a or b;
    layer1_outputs(3866) <= not b;
    layer1_outputs(3867) <= not a or b;
    layer1_outputs(3868) <= a or b;
    layer1_outputs(3869) <= not a;
    layer1_outputs(3870) <= not (a xor b);
    layer1_outputs(3871) <= not (a and b);
    layer1_outputs(3872) <= a and b;
    layer1_outputs(3873) <= a and b;
    layer1_outputs(3874) <= not (a and b);
    layer1_outputs(3875) <= '1';
    layer1_outputs(3876) <= '1';
    layer1_outputs(3877) <= '0';
    layer1_outputs(3878) <= a and not b;
    layer1_outputs(3879) <= b;
    layer1_outputs(3880) <= not (a and b);
    layer1_outputs(3881) <= b;
    layer1_outputs(3882) <= not (a or b);
    layer1_outputs(3883) <= a and not b;
    layer1_outputs(3884) <= not (a xor b);
    layer1_outputs(3885) <= a or b;
    layer1_outputs(3886) <= a;
    layer1_outputs(3887) <= not (a or b);
    layer1_outputs(3888) <= not a;
    layer1_outputs(3889) <= not (a xor b);
    layer1_outputs(3890) <= a;
    layer1_outputs(3891) <= not (a xor b);
    layer1_outputs(3892) <= not a or b;
    layer1_outputs(3893) <= b and not a;
    layer1_outputs(3894) <= not b;
    layer1_outputs(3895) <= b;
    layer1_outputs(3896) <= a or b;
    layer1_outputs(3897) <= a and not b;
    layer1_outputs(3898) <= a and b;
    layer1_outputs(3899) <= not a;
    layer1_outputs(3900) <= b;
    layer1_outputs(3901) <= '0';
    layer1_outputs(3902) <= b;
    layer1_outputs(3903) <= not b;
    layer1_outputs(3904) <= not b;
    layer1_outputs(3905) <= a;
    layer1_outputs(3906) <= a;
    layer1_outputs(3907) <= not a;
    layer1_outputs(3908) <= not a or b;
    layer1_outputs(3909) <= a and b;
    layer1_outputs(3910) <= not a or b;
    layer1_outputs(3911) <= not a or b;
    layer1_outputs(3912) <= not b;
    layer1_outputs(3913) <= not (a and b);
    layer1_outputs(3914) <= a;
    layer1_outputs(3915) <= not (a or b);
    layer1_outputs(3916) <= not a;
    layer1_outputs(3917) <= not b;
    layer1_outputs(3918) <= a;
    layer1_outputs(3919) <= b and not a;
    layer1_outputs(3920) <= not b or a;
    layer1_outputs(3921) <= not b;
    layer1_outputs(3922) <= not a;
    layer1_outputs(3923) <= a or b;
    layer1_outputs(3924) <= not b or a;
    layer1_outputs(3925) <= b;
    layer1_outputs(3926) <= a and b;
    layer1_outputs(3927) <= not a;
    layer1_outputs(3928) <= a;
    layer1_outputs(3929) <= not (a and b);
    layer1_outputs(3930) <= not b;
    layer1_outputs(3931) <= a;
    layer1_outputs(3932) <= a or b;
    layer1_outputs(3933) <= not b;
    layer1_outputs(3934) <= '1';
    layer1_outputs(3935) <= a or b;
    layer1_outputs(3936) <= b;
    layer1_outputs(3937) <= not a or b;
    layer1_outputs(3938) <= a or b;
    layer1_outputs(3939) <= not a;
    layer1_outputs(3940) <= b;
    layer1_outputs(3941) <= b and not a;
    layer1_outputs(3942) <= not a or b;
    layer1_outputs(3943) <= not a or b;
    layer1_outputs(3944) <= not (a or b);
    layer1_outputs(3945) <= a or b;
    layer1_outputs(3946) <= not b or a;
    layer1_outputs(3947) <= not (a or b);
    layer1_outputs(3948) <= not b;
    layer1_outputs(3949) <= not (a xor b);
    layer1_outputs(3950) <= a;
    layer1_outputs(3951) <= not a;
    layer1_outputs(3952) <= not a or b;
    layer1_outputs(3953) <= not a;
    layer1_outputs(3954) <= not b;
    layer1_outputs(3955) <= not a or b;
    layer1_outputs(3956) <= not b;
    layer1_outputs(3957) <= '1';
    layer1_outputs(3958) <= a;
    layer1_outputs(3959) <= not a;
    layer1_outputs(3960) <= not (a or b);
    layer1_outputs(3961) <= b and not a;
    layer1_outputs(3962) <= '1';
    layer1_outputs(3963) <= not b;
    layer1_outputs(3964) <= not b or a;
    layer1_outputs(3965) <= not a or b;
    layer1_outputs(3966) <= not a or b;
    layer1_outputs(3967) <= a;
    layer1_outputs(3968) <= a or b;
    layer1_outputs(3969) <= a;
    layer1_outputs(3970) <= '1';
    layer1_outputs(3971) <= not b;
    layer1_outputs(3972) <= b and not a;
    layer1_outputs(3973) <= not (a and b);
    layer1_outputs(3974) <= a or b;
    layer1_outputs(3975) <= not a or b;
    layer1_outputs(3976) <= not (a or b);
    layer1_outputs(3977) <= b;
    layer1_outputs(3978) <= a and not b;
    layer1_outputs(3979) <= b;
    layer1_outputs(3980) <= a and b;
    layer1_outputs(3981) <= not b;
    layer1_outputs(3982) <= a xor b;
    layer1_outputs(3983) <= '1';
    layer1_outputs(3984) <= a and b;
    layer1_outputs(3985) <= a;
    layer1_outputs(3986) <= a;
    layer1_outputs(3987) <= not a;
    layer1_outputs(3988) <= not b;
    layer1_outputs(3989) <= not (a and b);
    layer1_outputs(3990) <= a xor b;
    layer1_outputs(3991) <= a;
    layer1_outputs(3992) <= not (a or b);
    layer1_outputs(3993) <= b and not a;
    layer1_outputs(3994) <= a;
    layer1_outputs(3995) <= '0';
    layer1_outputs(3996) <= not b or a;
    layer1_outputs(3997) <= not (a or b);
    layer1_outputs(3998) <= not a or b;
    layer1_outputs(3999) <= a;
    layer1_outputs(4000) <= a or b;
    layer1_outputs(4001) <= a;
    layer1_outputs(4002) <= not b or a;
    layer1_outputs(4003) <= not (a or b);
    layer1_outputs(4004) <= b and not a;
    layer1_outputs(4005) <= not a;
    layer1_outputs(4006) <= '1';
    layer1_outputs(4007) <= b;
    layer1_outputs(4008) <= a and b;
    layer1_outputs(4009) <= not a or b;
    layer1_outputs(4010) <= not a or b;
    layer1_outputs(4011) <= not (a or b);
    layer1_outputs(4012) <= a or b;
    layer1_outputs(4013) <= a;
    layer1_outputs(4014) <= b and not a;
    layer1_outputs(4015) <= a xor b;
    layer1_outputs(4016) <= b;
    layer1_outputs(4017) <= not b;
    layer1_outputs(4018) <= a;
    layer1_outputs(4019) <= a;
    layer1_outputs(4020) <= b and not a;
    layer1_outputs(4021) <= not (a xor b);
    layer1_outputs(4022) <= a;
    layer1_outputs(4023) <= not a;
    layer1_outputs(4024) <= b;
    layer1_outputs(4025) <= a;
    layer1_outputs(4026) <= not (a and b);
    layer1_outputs(4027) <= a and b;
    layer1_outputs(4028) <= not b or a;
    layer1_outputs(4029) <= not (a or b);
    layer1_outputs(4030) <= b and not a;
    layer1_outputs(4031) <= b;
    layer1_outputs(4032) <= a and not b;
    layer1_outputs(4033) <= not (a and b);
    layer1_outputs(4034) <= not b or a;
    layer1_outputs(4035) <= a or b;
    layer1_outputs(4036) <= not a or b;
    layer1_outputs(4037) <= a and not b;
    layer1_outputs(4038) <= a;
    layer1_outputs(4039) <= not b;
    layer1_outputs(4040) <= a and b;
    layer1_outputs(4041) <= a and b;
    layer1_outputs(4042) <= not b or a;
    layer1_outputs(4043) <= not b;
    layer1_outputs(4044) <= not b;
    layer1_outputs(4045) <= not b or a;
    layer1_outputs(4046) <= a or b;
    layer1_outputs(4047) <= a and b;
    layer1_outputs(4048) <= b and not a;
    layer1_outputs(4049) <= a and not b;
    layer1_outputs(4050) <= not (a or b);
    layer1_outputs(4051) <= not b or a;
    layer1_outputs(4052) <= not b;
    layer1_outputs(4053) <= not (a or b);
    layer1_outputs(4054) <= a and b;
    layer1_outputs(4055) <= not (a or b);
    layer1_outputs(4056) <= a and not b;
    layer1_outputs(4057) <= not a;
    layer1_outputs(4058) <= b and not a;
    layer1_outputs(4059) <= b and not a;
    layer1_outputs(4060) <= b;
    layer1_outputs(4061) <= a and not b;
    layer1_outputs(4062) <= a;
    layer1_outputs(4063) <= b and not a;
    layer1_outputs(4064) <= a or b;
    layer1_outputs(4065) <= not b or a;
    layer1_outputs(4066) <= a and not b;
    layer1_outputs(4067) <= not b;
    layer1_outputs(4068) <= b;
    layer1_outputs(4069) <= a and not b;
    layer1_outputs(4070) <= a or b;
    layer1_outputs(4071) <= not b;
    layer1_outputs(4072) <= b and not a;
    layer1_outputs(4073) <= not (a or b);
    layer1_outputs(4074) <= b and not a;
    layer1_outputs(4075) <= '0';
    layer1_outputs(4076) <= a or b;
    layer1_outputs(4077) <= a or b;
    layer1_outputs(4078) <= b;
    layer1_outputs(4079) <= not a;
    layer1_outputs(4080) <= '0';
    layer1_outputs(4081) <= '1';
    layer1_outputs(4082) <= not (a or b);
    layer1_outputs(4083) <= a and not b;
    layer1_outputs(4084) <= a and b;
    layer1_outputs(4085) <= a;
    layer1_outputs(4086) <= a and b;
    layer1_outputs(4087) <= not (a or b);
    layer1_outputs(4088) <= not (a and b);
    layer1_outputs(4089) <= b and not a;
    layer1_outputs(4090) <= b;
    layer1_outputs(4091) <= a;
    layer1_outputs(4092) <= not (a xor b);
    layer1_outputs(4093) <= a;
    layer1_outputs(4094) <= a and not b;
    layer1_outputs(4095) <= a and not b;
    layer1_outputs(4096) <= a;
    layer1_outputs(4097) <= a or b;
    layer1_outputs(4098) <= not b or a;
    layer1_outputs(4099) <= a or b;
    layer1_outputs(4100) <= not b;
    layer1_outputs(4101) <= not a;
    layer1_outputs(4102) <= not (a xor b);
    layer1_outputs(4103) <= not (a and b);
    layer1_outputs(4104) <= not b;
    layer1_outputs(4105) <= not (a or b);
    layer1_outputs(4106) <= not a;
    layer1_outputs(4107) <= not a;
    layer1_outputs(4108) <= not a or b;
    layer1_outputs(4109) <= not a;
    layer1_outputs(4110) <= not (a xor b);
    layer1_outputs(4111) <= not a or b;
    layer1_outputs(4112) <= a xor b;
    layer1_outputs(4113) <= not (a and b);
    layer1_outputs(4114) <= not b;
    layer1_outputs(4115) <= b;
    layer1_outputs(4116) <= not a;
    layer1_outputs(4117) <= a and not b;
    layer1_outputs(4118) <= not b;
    layer1_outputs(4119) <= a;
    layer1_outputs(4120) <= a;
    layer1_outputs(4121) <= not (a or b);
    layer1_outputs(4122) <= not a;
    layer1_outputs(4123) <= a;
    layer1_outputs(4124) <= b and not a;
    layer1_outputs(4125) <= a;
    layer1_outputs(4126) <= a and not b;
    layer1_outputs(4127) <= '0';
    layer1_outputs(4128) <= a or b;
    layer1_outputs(4129) <= not b;
    layer1_outputs(4130) <= not a;
    layer1_outputs(4131) <= not a or b;
    layer1_outputs(4132) <= a or b;
    layer1_outputs(4133) <= not a or b;
    layer1_outputs(4134) <= not a;
    layer1_outputs(4135) <= b;
    layer1_outputs(4136) <= '0';
    layer1_outputs(4137) <= a and b;
    layer1_outputs(4138) <= not (a or b);
    layer1_outputs(4139) <= not b or a;
    layer1_outputs(4140) <= a or b;
    layer1_outputs(4141) <= b;
    layer1_outputs(4142) <= not (a or b);
    layer1_outputs(4143) <= b;
    layer1_outputs(4144) <= not (a and b);
    layer1_outputs(4145) <= '0';
    layer1_outputs(4146) <= a or b;
    layer1_outputs(4147) <= not b;
    layer1_outputs(4148) <= b and not a;
    layer1_outputs(4149) <= not b or a;
    layer1_outputs(4150) <= not b or a;
    layer1_outputs(4151) <= not a or b;
    layer1_outputs(4152) <= not b;
    layer1_outputs(4153) <= not a;
    layer1_outputs(4154) <= '0';
    layer1_outputs(4155) <= b and not a;
    layer1_outputs(4156) <= a xor b;
    layer1_outputs(4157) <= a;
    layer1_outputs(4158) <= not b or a;
    layer1_outputs(4159) <= not (a and b);
    layer1_outputs(4160) <= a;
    layer1_outputs(4161) <= '1';
    layer1_outputs(4162) <= not b;
    layer1_outputs(4163) <= b and not a;
    layer1_outputs(4164) <= a and b;
    layer1_outputs(4165) <= b;
    layer1_outputs(4166) <= not (a xor b);
    layer1_outputs(4167) <= not (a xor b);
    layer1_outputs(4168) <= '0';
    layer1_outputs(4169) <= a or b;
    layer1_outputs(4170) <= b and not a;
    layer1_outputs(4171) <= not (a and b);
    layer1_outputs(4172) <= a;
    layer1_outputs(4173) <= b;
    layer1_outputs(4174) <= not a;
    layer1_outputs(4175) <= not (a and b);
    layer1_outputs(4176) <= not a or b;
    layer1_outputs(4177) <= not (a and b);
    layer1_outputs(4178) <= not (a xor b);
    layer1_outputs(4179) <= a or b;
    layer1_outputs(4180) <= a or b;
    layer1_outputs(4181) <= b;
    layer1_outputs(4182) <= a;
    layer1_outputs(4183) <= not b or a;
    layer1_outputs(4184) <= a and b;
    layer1_outputs(4185) <= not (a or b);
    layer1_outputs(4186) <= not (a and b);
    layer1_outputs(4187) <= not b or a;
    layer1_outputs(4188) <= b;
    layer1_outputs(4189) <= '0';
    layer1_outputs(4190) <= a or b;
    layer1_outputs(4191) <= not a;
    layer1_outputs(4192) <= not a;
    layer1_outputs(4193) <= a;
    layer1_outputs(4194) <= b and not a;
    layer1_outputs(4195) <= not a;
    layer1_outputs(4196) <= a xor b;
    layer1_outputs(4197) <= b;
    layer1_outputs(4198) <= not (a xor b);
    layer1_outputs(4199) <= not b or a;
    layer1_outputs(4200) <= not a;
    layer1_outputs(4201) <= '0';
    layer1_outputs(4202) <= not a or b;
    layer1_outputs(4203) <= '1';
    layer1_outputs(4204) <= a and b;
    layer1_outputs(4205) <= not (a or b);
    layer1_outputs(4206) <= b;
    layer1_outputs(4207) <= a or b;
    layer1_outputs(4208) <= a xor b;
    layer1_outputs(4209) <= a and not b;
    layer1_outputs(4210) <= not (a or b);
    layer1_outputs(4211) <= b;
    layer1_outputs(4212) <= a xor b;
    layer1_outputs(4213) <= a and not b;
    layer1_outputs(4214) <= b;
    layer1_outputs(4215) <= not b;
    layer1_outputs(4216) <= not a;
    layer1_outputs(4217) <= not b or a;
    layer1_outputs(4218) <= a xor b;
    layer1_outputs(4219) <= a or b;
    layer1_outputs(4220) <= a xor b;
    layer1_outputs(4221) <= not (a or b);
    layer1_outputs(4222) <= a xor b;
    layer1_outputs(4223) <= a and b;
    layer1_outputs(4224) <= b;
    layer1_outputs(4225) <= a and b;
    layer1_outputs(4226) <= not a or b;
    layer1_outputs(4227) <= b;
    layer1_outputs(4228) <= '0';
    layer1_outputs(4229) <= not (a or b);
    layer1_outputs(4230) <= b;
    layer1_outputs(4231) <= a and not b;
    layer1_outputs(4232) <= not b;
    layer1_outputs(4233) <= '1';
    layer1_outputs(4234) <= b and not a;
    layer1_outputs(4235) <= a;
    layer1_outputs(4236) <= not b or a;
    layer1_outputs(4237) <= not (a xor b);
    layer1_outputs(4238) <= not a or b;
    layer1_outputs(4239) <= a and not b;
    layer1_outputs(4240) <= '0';
    layer1_outputs(4241) <= b and not a;
    layer1_outputs(4242) <= not (a and b);
    layer1_outputs(4243) <= not (a and b);
    layer1_outputs(4244) <= not b or a;
    layer1_outputs(4245) <= a xor b;
    layer1_outputs(4246) <= not a;
    layer1_outputs(4247) <= b;
    layer1_outputs(4248) <= a and not b;
    layer1_outputs(4249) <= a;
    layer1_outputs(4250) <= '0';
    layer1_outputs(4251) <= not (a or b);
    layer1_outputs(4252) <= not (a or b);
    layer1_outputs(4253) <= '0';
    layer1_outputs(4254) <= not a;
    layer1_outputs(4255) <= a;
    layer1_outputs(4256) <= '0';
    layer1_outputs(4257) <= not a;
    layer1_outputs(4258) <= not (a and b);
    layer1_outputs(4259) <= a;
    layer1_outputs(4260) <= not a;
    layer1_outputs(4261) <= a;
    layer1_outputs(4262) <= b;
    layer1_outputs(4263) <= b;
    layer1_outputs(4264) <= not a;
    layer1_outputs(4265) <= not (a xor b);
    layer1_outputs(4266) <= not a;
    layer1_outputs(4267) <= a xor b;
    layer1_outputs(4268) <= b;
    layer1_outputs(4269) <= not (a and b);
    layer1_outputs(4270) <= not (a or b);
    layer1_outputs(4271) <= a;
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= not b or a;
    layer1_outputs(4274) <= a;
    layer1_outputs(4275) <= '1';
    layer1_outputs(4276) <= a or b;
    layer1_outputs(4277) <= not (a and b);
    layer1_outputs(4278) <= not (a or b);
    layer1_outputs(4279) <= not a or b;
    layer1_outputs(4280) <= b;
    layer1_outputs(4281) <= b and not a;
    layer1_outputs(4282) <= not a or b;
    layer1_outputs(4283) <= b;
    layer1_outputs(4284) <= b;
    layer1_outputs(4285) <= a;
    layer1_outputs(4286) <= not b;
    layer1_outputs(4287) <= a or b;
    layer1_outputs(4288) <= a and not b;
    layer1_outputs(4289) <= not b;
    layer1_outputs(4290) <= not b or a;
    layer1_outputs(4291) <= not b;
    layer1_outputs(4292) <= not b or a;
    layer1_outputs(4293) <= b;
    layer1_outputs(4294) <= a and b;
    layer1_outputs(4295) <= a and not b;
    layer1_outputs(4296) <= not a;
    layer1_outputs(4297) <= not b or a;
    layer1_outputs(4298) <= not b or a;
    layer1_outputs(4299) <= a and not b;
    layer1_outputs(4300) <= b;
    layer1_outputs(4301) <= not a or b;
    layer1_outputs(4302) <= b and not a;
    layer1_outputs(4303) <= a and b;
    layer1_outputs(4304) <= not b or a;
    layer1_outputs(4305) <= b;
    layer1_outputs(4306) <= '1';
    layer1_outputs(4307) <= not b or a;
    layer1_outputs(4308) <= '1';
    layer1_outputs(4309) <= not (a or b);
    layer1_outputs(4310) <= not (a and b);
    layer1_outputs(4311) <= not a;
    layer1_outputs(4312) <= not a or b;
    layer1_outputs(4313) <= '0';
    layer1_outputs(4314) <= not b or a;
    layer1_outputs(4315) <= a;
    layer1_outputs(4316) <= not a or b;
    layer1_outputs(4317) <= not b;
    layer1_outputs(4318) <= '1';
    layer1_outputs(4319) <= a or b;
    layer1_outputs(4320) <= not (a and b);
    layer1_outputs(4321) <= b;
    layer1_outputs(4322) <= a xor b;
    layer1_outputs(4323) <= a or b;
    layer1_outputs(4324) <= b and not a;
    layer1_outputs(4325) <= b and not a;
    layer1_outputs(4326) <= '1';
    layer1_outputs(4327) <= a;
    layer1_outputs(4328) <= a and b;
    layer1_outputs(4329) <= not (a xor b);
    layer1_outputs(4330) <= a;
    layer1_outputs(4331) <= not b;
    layer1_outputs(4332) <= b;
    layer1_outputs(4333) <= not b;
    layer1_outputs(4334) <= b and not a;
    layer1_outputs(4335) <= '0';
    layer1_outputs(4336) <= a or b;
    layer1_outputs(4337) <= a;
    layer1_outputs(4338) <= not b or a;
    layer1_outputs(4339) <= not (a xor b);
    layer1_outputs(4340) <= not (a or b);
    layer1_outputs(4341) <= not (a xor b);
    layer1_outputs(4342) <= not a;
    layer1_outputs(4343) <= a and not b;
    layer1_outputs(4344) <= b and not a;
    layer1_outputs(4345) <= b;
    layer1_outputs(4346) <= '1';
    layer1_outputs(4347) <= '1';
    layer1_outputs(4348) <= a and b;
    layer1_outputs(4349) <= b;
    layer1_outputs(4350) <= a;
    layer1_outputs(4351) <= not b or a;
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= b and not a;
    layer1_outputs(4354) <= not a or b;
    layer1_outputs(4355) <= not a;
    layer1_outputs(4356) <= a or b;
    layer1_outputs(4357) <= not b;
    layer1_outputs(4358) <= a or b;
    layer1_outputs(4359) <= a and not b;
    layer1_outputs(4360) <= not (a or b);
    layer1_outputs(4361) <= not (a or b);
    layer1_outputs(4362) <= not b;
    layer1_outputs(4363) <= not b;
    layer1_outputs(4364) <= b and not a;
    layer1_outputs(4365) <= not (a and b);
    layer1_outputs(4366) <= not b;
    layer1_outputs(4367) <= not b;
    layer1_outputs(4368) <= not b;
    layer1_outputs(4369) <= a;
    layer1_outputs(4370) <= not (a or b);
    layer1_outputs(4371) <= not a or b;
    layer1_outputs(4372) <= not a;
    layer1_outputs(4373) <= not b or a;
    layer1_outputs(4374) <= a and b;
    layer1_outputs(4375) <= a and b;
    layer1_outputs(4376) <= b and not a;
    layer1_outputs(4377) <= a and not b;
    layer1_outputs(4378) <= not (a xor b);
    layer1_outputs(4379) <= a;
    layer1_outputs(4380) <= '0';
    layer1_outputs(4381) <= b;
    layer1_outputs(4382) <= not a or b;
    layer1_outputs(4383) <= a and not b;
    layer1_outputs(4384) <= b;
    layer1_outputs(4385) <= not a or b;
    layer1_outputs(4386) <= a;
    layer1_outputs(4387) <= b;
    layer1_outputs(4388) <= a;
    layer1_outputs(4389) <= a or b;
    layer1_outputs(4390) <= not (a or b);
    layer1_outputs(4391) <= b;
    layer1_outputs(4392) <= a or b;
    layer1_outputs(4393) <= not (a and b);
    layer1_outputs(4394) <= not (a or b);
    layer1_outputs(4395) <= not (a xor b);
    layer1_outputs(4396) <= b and not a;
    layer1_outputs(4397) <= '0';
    layer1_outputs(4398) <= a and b;
    layer1_outputs(4399) <= not (a xor b);
    layer1_outputs(4400) <= '0';
    layer1_outputs(4401) <= not b or a;
    layer1_outputs(4402) <= not (a and b);
    layer1_outputs(4403) <= not a;
    layer1_outputs(4404) <= a;
    layer1_outputs(4405) <= not (a xor b);
    layer1_outputs(4406) <= a xor b;
    layer1_outputs(4407) <= not b;
    layer1_outputs(4408) <= not b;
    layer1_outputs(4409) <= b;
    layer1_outputs(4410) <= not (a and b);
    layer1_outputs(4411) <= not a;
    layer1_outputs(4412) <= not b;
    layer1_outputs(4413) <= not (a xor b);
    layer1_outputs(4414) <= not a or b;
    layer1_outputs(4415) <= a or b;
    layer1_outputs(4416) <= not a;
    layer1_outputs(4417) <= not (a or b);
    layer1_outputs(4418) <= a and b;
    layer1_outputs(4419) <= a or b;
    layer1_outputs(4420) <= not b;
    layer1_outputs(4421) <= not (a or b);
    layer1_outputs(4422) <= not (a or b);
    layer1_outputs(4423) <= not b or a;
    layer1_outputs(4424) <= a or b;
    layer1_outputs(4425) <= not b;
    layer1_outputs(4426) <= not a;
    layer1_outputs(4427) <= not a or b;
    layer1_outputs(4428) <= '1';
    layer1_outputs(4429) <= a and b;
    layer1_outputs(4430) <= a;
    layer1_outputs(4431) <= not b;
    layer1_outputs(4432) <= not b or a;
    layer1_outputs(4433) <= not (a xor b);
    layer1_outputs(4434) <= a or b;
    layer1_outputs(4435) <= not b or a;
    layer1_outputs(4436) <= b;
    layer1_outputs(4437) <= a and b;
    layer1_outputs(4438) <= b and not a;
    layer1_outputs(4439) <= not b or a;
    layer1_outputs(4440) <= b and not a;
    layer1_outputs(4441) <= not (a xor b);
    layer1_outputs(4442) <= a;
    layer1_outputs(4443) <= not b or a;
    layer1_outputs(4444) <= a and b;
    layer1_outputs(4445) <= a and b;
    layer1_outputs(4446) <= not (a or b);
    layer1_outputs(4447) <= not (a or b);
    layer1_outputs(4448) <= a and not b;
    layer1_outputs(4449) <= a;
    layer1_outputs(4450) <= a or b;
    layer1_outputs(4451) <= not (a and b);
    layer1_outputs(4452) <= a or b;
    layer1_outputs(4453) <= not (a or b);
    layer1_outputs(4454) <= not a or b;
    layer1_outputs(4455) <= a and b;
    layer1_outputs(4456) <= '0';
    layer1_outputs(4457) <= not (a and b);
    layer1_outputs(4458) <= a and not b;
    layer1_outputs(4459) <= not b;
    layer1_outputs(4460) <= not a or b;
    layer1_outputs(4461) <= not a or b;
    layer1_outputs(4462) <= a and b;
    layer1_outputs(4463) <= not a;
    layer1_outputs(4464) <= a or b;
    layer1_outputs(4465) <= b;
    layer1_outputs(4466) <= not (a xor b);
    layer1_outputs(4467) <= a or b;
    layer1_outputs(4468) <= a and b;
    layer1_outputs(4469) <= a and b;
    layer1_outputs(4470) <= not (a or b);
    layer1_outputs(4471) <= '0';
    layer1_outputs(4472) <= a and not b;
    layer1_outputs(4473) <= '0';
    layer1_outputs(4474) <= b;
    layer1_outputs(4475) <= a or b;
    layer1_outputs(4476) <= not (a and b);
    layer1_outputs(4477) <= b and not a;
    layer1_outputs(4478) <= a or b;
    layer1_outputs(4479) <= not (a and b);
    layer1_outputs(4480) <= a and not b;
    layer1_outputs(4481) <= a and not b;
    layer1_outputs(4482) <= a and not b;
    layer1_outputs(4483) <= '1';
    layer1_outputs(4484) <= not (a or b);
    layer1_outputs(4485) <= b;
    layer1_outputs(4486) <= '0';
    layer1_outputs(4487) <= a and not b;
    layer1_outputs(4488) <= a or b;
    layer1_outputs(4489) <= not (a or b);
    layer1_outputs(4490) <= a and b;
    layer1_outputs(4491) <= not b or a;
    layer1_outputs(4492) <= not a;
    layer1_outputs(4493) <= a xor b;
    layer1_outputs(4494) <= not a or b;
    layer1_outputs(4495) <= a and b;
    layer1_outputs(4496) <= a or b;
    layer1_outputs(4497) <= a and b;
    layer1_outputs(4498) <= not (a and b);
    layer1_outputs(4499) <= b and not a;
    layer1_outputs(4500) <= not a or b;
    layer1_outputs(4501) <= a and not b;
    layer1_outputs(4502) <= not (a or b);
    layer1_outputs(4503) <= not (a or b);
    layer1_outputs(4504) <= b;
    layer1_outputs(4505) <= a and b;
    layer1_outputs(4506) <= a and b;
    layer1_outputs(4507) <= b;
    layer1_outputs(4508) <= not b or a;
    layer1_outputs(4509) <= not a or b;
    layer1_outputs(4510) <= not a;
    layer1_outputs(4511) <= a and b;
    layer1_outputs(4512) <= b;
    layer1_outputs(4513) <= a;
    layer1_outputs(4514) <= b and not a;
    layer1_outputs(4515) <= '1';
    layer1_outputs(4516) <= a;
    layer1_outputs(4517) <= b and not a;
    layer1_outputs(4518) <= b and not a;
    layer1_outputs(4519) <= not b;
    layer1_outputs(4520) <= not b or a;
    layer1_outputs(4521) <= not (a and b);
    layer1_outputs(4522) <= b;
    layer1_outputs(4523) <= not (a and b);
    layer1_outputs(4524) <= b;
    layer1_outputs(4525) <= not (a and b);
    layer1_outputs(4526) <= not b;
    layer1_outputs(4527) <= not b or a;
    layer1_outputs(4528) <= b and not a;
    layer1_outputs(4529) <= a;
    layer1_outputs(4530) <= not b;
    layer1_outputs(4531) <= a;
    layer1_outputs(4532) <= a and b;
    layer1_outputs(4533) <= b;
    layer1_outputs(4534) <= b and not a;
    layer1_outputs(4535) <= not a;
    layer1_outputs(4536) <= not (a or b);
    layer1_outputs(4537) <= b;
    layer1_outputs(4538) <= b;
    layer1_outputs(4539) <= not a;
    layer1_outputs(4540) <= a;
    layer1_outputs(4541) <= not b;
    layer1_outputs(4542) <= a and not b;
    layer1_outputs(4543) <= a and b;
    layer1_outputs(4544) <= b;
    layer1_outputs(4545) <= not a;
    layer1_outputs(4546) <= b;
    layer1_outputs(4547) <= not a;
    layer1_outputs(4548) <= a;
    layer1_outputs(4549) <= not (a or b);
    layer1_outputs(4550) <= b and not a;
    layer1_outputs(4551) <= not b;
    layer1_outputs(4552) <= '1';
    layer1_outputs(4553) <= not b;
    layer1_outputs(4554) <= not a;
    layer1_outputs(4555) <= b and not a;
    layer1_outputs(4556) <= not a or b;
    layer1_outputs(4557) <= a;
    layer1_outputs(4558) <= a;
    layer1_outputs(4559) <= b and not a;
    layer1_outputs(4560) <= not b;
    layer1_outputs(4561) <= not a;
    layer1_outputs(4562) <= not b;
    layer1_outputs(4563) <= not (a or b);
    layer1_outputs(4564) <= a;
    layer1_outputs(4565) <= not a;
    layer1_outputs(4566) <= a and not b;
    layer1_outputs(4567) <= a and not b;
    layer1_outputs(4568) <= a and not b;
    layer1_outputs(4569) <= b and not a;
    layer1_outputs(4570) <= not a or b;
    layer1_outputs(4571) <= not (a and b);
    layer1_outputs(4572) <= not b;
    layer1_outputs(4573) <= not b;
    layer1_outputs(4574) <= not a;
    layer1_outputs(4575) <= '1';
    layer1_outputs(4576) <= not a;
    layer1_outputs(4577) <= not b or a;
    layer1_outputs(4578) <= a and b;
    layer1_outputs(4579) <= b and not a;
    layer1_outputs(4580) <= '1';
    layer1_outputs(4581) <= a and b;
    layer1_outputs(4582) <= b and not a;
    layer1_outputs(4583) <= not (a xor b);
    layer1_outputs(4584) <= not b or a;
    layer1_outputs(4585) <= b and not a;
    layer1_outputs(4586) <= a and not b;
    layer1_outputs(4587) <= a;
    layer1_outputs(4588) <= not (a or b);
    layer1_outputs(4589) <= '0';
    layer1_outputs(4590) <= not a;
    layer1_outputs(4591) <= b and not a;
    layer1_outputs(4592) <= not (a and b);
    layer1_outputs(4593) <= a and not b;
    layer1_outputs(4594) <= not a or b;
    layer1_outputs(4595) <= not (a or b);
    layer1_outputs(4596) <= not (a xor b);
    layer1_outputs(4597) <= a;
    layer1_outputs(4598) <= not (a or b);
    layer1_outputs(4599) <= not b or a;
    layer1_outputs(4600) <= not (a and b);
    layer1_outputs(4601) <= a or b;
    layer1_outputs(4602) <= not b;
    layer1_outputs(4603) <= a or b;
    layer1_outputs(4604) <= not (a and b);
    layer1_outputs(4605) <= not a;
    layer1_outputs(4606) <= a xor b;
    layer1_outputs(4607) <= not b;
    layer1_outputs(4608) <= a;
    layer1_outputs(4609) <= not (a xor b);
    layer1_outputs(4610) <= a and b;
    layer1_outputs(4611) <= a and b;
    layer1_outputs(4612) <= a;
    layer1_outputs(4613) <= not b or a;
    layer1_outputs(4614) <= a;
    layer1_outputs(4615) <= not b;
    layer1_outputs(4616) <= '1';
    layer1_outputs(4617) <= not (a or b);
    layer1_outputs(4618) <= not b or a;
    layer1_outputs(4619) <= not b or a;
    layer1_outputs(4620) <= a xor b;
    layer1_outputs(4621) <= '1';
    layer1_outputs(4622) <= not (a xor b);
    layer1_outputs(4623) <= not a or b;
    layer1_outputs(4624) <= b;
    layer1_outputs(4625) <= b;
    layer1_outputs(4626) <= b and not a;
    layer1_outputs(4627) <= not (a or b);
    layer1_outputs(4628) <= not b or a;
    layer1_outputs(4629) <= '0';
    layer1_outputs(4630) <= a and not b;
    layer1_outputs(4631) <= not b or a;
    layer1_outputs(4632) <= not a or b;
    layer1_outputs(4633) <= b;
    layer1_outputs(4634) <= a;
    layer1_outputs(4635) <= '0';
    layer1_outputs(4636) <= not b;
    layer1_outputs(4637) <= b and not a;
    layer1_outputs(4638) <= not (a or b);
    layer1_outputs(4639) <= not a;
    layer1_outputs(4640) <= a or b;
    layer1_outputs(4641) <= b;
    layer1_outputs(4642) <= a;
    layer1_outputs(4643) <= not a or b;
    layer1_outputs(4644) <= a and b;
    layer1_outputs(4645) <= not b;
    layer1_outputs(4646) <= not b;
    layer1_outputs(4647) <= not (a or b);
    layer1_outputs(4648) <= a;
    layer1_outputs(4649) <= not b or a;
    layer1_outputs(4650) <= not b or a;
    layer1_outputs(4651) <= a;
    layer1_outputs(4652) <= a or b;
    layer1_outputs(4653) <= not b;
    layer1_outputs(4654) <= a and b;
    layer1_outputs(4655) <= not b;
    layer1_outputs(4656) <= a;
    layer1_outputs(4657) <= a and b;
    layer1_outputs(4658) <= b and not a;
    layer1_outputs(4659) <= not a;
    layer1_outputs(4660) <= not (a xor b);
    layer1_outputs(4661) <= a and not b;
    layer1_outputs(4662) <= not a;
    layer1_outputs(4663) <= a;
    layer1_outputs(4664) <= not a;
    layer1_outputs(4665) <= not (a and b);
    layer1_outputs(4666) <= a or b;
    layer1_outputs(4667) <= not b;
    layer1_outputs(4668) <= not b;
    layer1_outputs(4669) <= not a or b;
    layer1_outputs(4670) <= a xor b;
    layer1_outputs(4671) <= a xor b;
    layer1_outputs(4672) <= not a or b;
    layer1_outputs(4673) <= not b or a;
    layer1_outputs(4674) <= not a;
    layer1_outputs(4675) <= a;
    layer1_outputs(4676) <= '0';
    layer1_outputs(4677) <= not b;
    layer1_outputs(4678) <= '1';
    layer1_outputs(4679) <= a;
    layer1_outputs(4680) <= b;
    layer1_outputs(4681) <= '1';
    layer1_outputs(4682) <= not b;
    layer1_outputs(4683) <= not b or a;
    layer1_outputs(4684) <= not (a or b);
    layer1_outputs(4685) <= not b or a;
    layer1_outputs(4686) <= not (a and b);
    layer1_outputs(4687) <= a and not b;
    layer1_outputs(4688) <= a xor b;
    layer1_outputs(4689) <= not b;
    layer1_outputs(4690) <= '0';
    layer1_outputs(4691) <= b and not a;
    layer1_outputs(4692) <= not (a or b);
    layer1_outputs(4693) <= b;
    layer1_outputs(4694) <= not a or b;
    layer1_outputs(4695) <= a and not b;
    layer1_outputs(4696) <= not b or a;
    layer1_outputs(4697) <= b;
    layer1_outputs(4698) <= not a;
    layer1_outputs(4699) <= a and b;
    layer1_outputs(4700) <= a and not b;
    layer1_outputs(4701) <= not (a and b);
    layer1_outputs(4702) <= a and b;
    layer1_outputs(4703) <= '1';
    layer1_outputs(4704) <= a or b;
    layer1_outputs(4705) <= b;
    layer1_outputs(4706) <= a and not b;
    layer1_outputs(4707) <= a or b;
    layer1_outputs(4708) <= '0';
    layer1_outputs(4709) <= a and not b;
    layer1_outputs(4710) <= a and not b;
    layer1_outputs(4711) <= a;
    layer1_outputs(4712) <= a;
    layer1_outputs(4713) <= not (a or b);
    layer1_outputs(4714) <= not b or a;
    layer1_outputs(4715) <= b and not a;
    layer1_outputs(4716) <= b and not a;
    layer1_outputs(4717) <= a and b;
    layer1_outputs(4718) <= not b or a;
    layer1_outputs(4719) <= not (a or b);
    layer1_outputs(4720) <= not (a xor b);
    layer1_outputs(4721) <= a and not b;
    layer1_outputs(4722) <= not b;
    layer1_outputs(4723) <= a and not b;
    layer1_outputs(4724) <= not (a xor b);
    layer1_outputs(4725) <= b and not a;
    layer1_outputs(4726) <= not a;
    layer1_outputs(4727) <= a and not b;
    layer1_outputs(4728) <= b and not a;
    layer1_outputs(4729) <= b;
    layer1_outputs(4730) <= b and not a;
    layer1_outputs(4731) <= not (a and b);
    layer1_outputs(4732) <= a or b;
    layer1_outputs(4733) <= '1';
    layer1_outputs(4734) <= not b;
    layer1_outputs(4735) <= not (a and b);
    layer1_outputs(4736) <= b and not a;
    layer1_outputs(4737) <= not a;
    layer1_outputs(4738) <= not b;
    layer1_outputs(4739) <= not (a xor b);
    layer1_outputs(4740) <= not a or b;
    layer1_outputs(4741) <= a and not b;
    layer1_outputs(4742) <= not b or a;
    layer1_outputs(4743) <= not b;
    layer1_outputs(4744) <= not b;
    layer1_outputs(4745) <= a and b;
    layer1_outputs(4746) <= a and b;
    layer1_outputs(4747) <= b;
    layer1_outputs(4748) <= not (a and b);
    layer1_outputs(4749) <= not (a and b);
    layer1_outputs(4750) <= '1';
    layer1_outputs(4751) <= not a;
    layer1_outputs(4752) <= not a or b;
    layer1_outputs(4753) <= b;
    layer1_outputs(4754) <= not b or a;
    layer1_outputs(4755) <= a xor b;
    layer1_outputs(4756) <= not a;
    layer1_outputs(4757) <= a;
    layer1_outputs(4758) <= not (a and b);
    layer1_outputs(4759) <= not b;
    layer1_outputs(4760) <= a or b;
    layer1_outputs(4761) <= not b or a;
    layer1_outputs(4762) <= not b;
    layer1_outputs(4763) <= b and not a;
    layer1_outputs(4764) <= not (a and b);
    layer1_outputs(4765) <= '1';
    layer1_outputs(4766) <= not a;
    layer1_outputs(4767) <= b;
    layer1_outputs(4768) <= b;
    layer1_outputs(4769) <= a and not b;
    layer1_outputs(4770) <= not (a xor b);
    layer1_outputs(4771) <= a and not b;
    layer1_outputs(4772) <= not (a or b);
    layer1_outputs(4773) <= a and not b;
    layer1_outputs(4774) <= a or b;
    layer1_outputs(4775) <= not (a or b);
    layer1_outputs(4776) <= b;
    layer1_outputs(4777) <= a and b;
    layer1_outputs(4778) <= not b or a;
    layer1_outputs(4779) <= b;
    layer1_outputs(4780) <= not b or a;
    layer1_outputs(4781) <= '1';
    layer1_outputs(4782) <= b;
    layer1_outputs(4783) <= not a;
    layer1_outputs(4784) <= not (a and b);
    layer1_outputs(4785) <= a;
    layer1_outputs(4786) <= not (a and b);
    layer1_outputs(4787) <= b;
    layer1_outputs(4788) <= not b;
    layer1_outputs(4789) <= '0';
    layer1_outputs(4790) <= a;
    layer1_outputs(4791) <= not b or a;
    layer1_outputs(4792) <= not a;
    layer1_outputs(4793) <= not b or a;
    layer1_outputs(4794) <= b and not a;
    layer1_outputs(4795) <= a or b;
    layer1_outputs(4796) <= not a;
    layer1_outputs(4797) <= not (a and b);
    layer1_outputs(4798) <= not (a and b);
    layer1_outputs(4799) <= not b;
    layer1_outputs(4800) <= b;
    layer1_outputs(4801) <= not b;
    layer1_outputs(4802) <= not a or b;
    layer1_outputs(4803) <= b;
    layer1_outputs(4804) <= a;
    layer1_outputs(4805) <= not b;
    layer1_outputs(4806) <= not (a and b);
    layer1_outputs(4807) <= '1';
    layer1_outputs(4808) <= not a or b;
    layer1_outputs(4809) <= not (a and b);
    layer1_outputs(4810) <= a xor b;
    layer1_outputs(4811) <= a and b;
    layer1_outputs(4812) <= a and not b;
    layer1_outputs(4813) <= a and b;
    layer1_outputs(4814) <= '0';
    layer1_outputs(4815) <= not (a and b);
    layer1_outputs(4816) <= not a or b;
    layer1_outputs(4817) <= b;
    layer1_outputs(4818) <= not a;
    layer1_outputs(4819) <= a or b;
    layer1_outputs(4820) <= not (a xor b);
    layer1_outputs(4821) <= '1';
    layer1_outputs(4822) <= not b or a;
    layer1_outputs(4823) <= '1';
    layer1_outputs(4824) <= a and b;
    layer1_outputs(4825) <= not b;
    layer1_outputs(4826) <= a;
    layer1_outputs(4827) <= not (a or b);
    layer1_outputs(4828) <= not a or b;
    layer1_outputs(4829) <= b;
    layer1_outputs(4830) <= a and b;
    layer1_outputs(4831) <= a;
    layer1_outputs(4832) <= b;
    layer1_outputs(4833) <= '1';
    layer1_outputs(4834) <= a xor b;
    layer1_outputs(4835) <= not b;
    layer1_outputs(4836) <= not b;
    layer1_outputs(4837) <= b and not a;
    layer1_outputs(4838) <= not b;
    layer1_outputs(4839) <= b and not a;
    layer1_outputs(4840) <= not b or a;
    layer1_outputs(4841) <= not b or a;
    layer1_outputs(4842) <= not a;
    layer1_outputs(4843) <= a and b;
    layer1_outputs(4844) <= a;
    layer1_outputs(4845) <= not a;
    layer1_outputs(4846) <= not b or a;
    layer1_outputs(4847) <= a and b;
    layer1_outputs(4848) <= not a;
    layer1_outputs(4849) <= b;
    layer1_outputs(4850) <= a and not b;
    layer1_outputs(4851) <= a xor b;
    layer1_outputs(4852) <= b;
    layer1_outputs(4853) <= b;
    layer1_outputs(4854) <= a;
    layer1_outputs(4855) <= not b;
    layer1_outputs(4856) <= a and b;
    layer1_outputs(4857) <= a;
    layer1_outputs(4858) <= '1';
    layer1_outputs(4859) <= not a;
    layer1_outputs(4860) <= not (a and b);
    layer1_outputs(4861) <= a xor b;
    layer1_outputs(4862) <= not (a or b);
    layer1_outputs(4863) <= not (a xor b);
    layer1_outputs(4864) <= a and not b;
    layer1_outputs(4865) <= not a;
    layer1_outputs(4866) <= not b;
    layer1_outputs(4867) <= b and not a;
    layer1_outputs(4868) <= not a;
    layer1_outputs(4869) <= a and not b;
    layer1_outputs(4870) <= b;
    layer1_outputs(4871) <= not b;
    layer1_outputs(4872) <= a xor b;
    layer1_outputs(4873) <= a or b;
    layer1_outputs(4874) <= not b or a;
    layer1_outputs(4875) <= a or b;
    layer1_outputs(4876) <= a;
    layer1_outputs(4877) <= not (a xor b);
    layer1_outputs(4878) <= not a or b;
    layer1_outputs(4879) <= a and b;
    layer1_outputs(4880) <= a;
    layer1_outputs(4881) <= not b;
    layer1_outputs(4882) <= a and not b;
    layer1_outputs(4883) <= '1';
    layer1_outputs(4884) <= not (a or b);
    layer1_outputs(4885) <= not b;
    layer1_outputs(4886) <= not (a and b);
    layer1_outputs(4887) <= b;
    layer1_outputs(4888) <= b;
    layer1_outputs(4889) <= not b;
    layer1_outputs(4890) <= not a;
    layer1_outputs(4891) <= b and not a;
    layer1_outputs(4892) <= '0';
    layer1_outputs(4893) <= a and not b;
    layer1_outputs(4894) <= not a;
    layer1_outputs(4895) <= '0';
    layer1_outputs(4896) <= not a or b;
    layer1_outputs(4897) <= not a;
    layer1_outputs(4898) <= '0';
    layer1_outputs(4899) <= b and not a;
    layer1_outputs(4900) <= a and not b;
    layer1_outputs(4901) <= not a;
    layer1_outputs(4902) <= '1';
    layer1_outputs(4903) <= a or b;
    layer1_outputs(4904) <= a;
    layer1_outputs(4905) <= a and b;
    layer1_outputs(4906) <= not b;
    layer1_outputs(4907) <= a and b;
    layer1_outputs(4908) <= not a or b;
    layer1_outputs(4909) <= not (a or b);
    layer1_outputs(4910) <= not b;
    layer1_outputs(4911) <= not (a and b);
    layer1_outputs(4912) <= not (a xor b);
    layer1_outputs(4913) <= not (a and b);
    layer1_outputs(4914) <= not (a xor b);
    layer1_outputs(4915) <= b and not a;
    layer1_outputs(4916) <= not b or a;
    layer1_outputs(4917) <= a and not b;
    layer1_outputs(4918) <= b;
    layer1_outputs(4919) <= not b or a;
    layer1_outputs(4920) <= '1';
    layer1_outputs(4921) <= not a or b;
    layer1_outputs(4922) <= not (a or b);
    layer1_outputs(4923) <= a;
    layer1_outputs(4924) <= '0';
    layer1_outputs(4925) <= not (a or b);
    layer1_outputs(4926) <= b;
    layer1_outputs(4927) <= not (a and b);
    layer1_outputs(4928) <= b;
    layer1_outputs(4929) <= not a;
    layer1_outputs(4930) <= a;
    layer1_outputs(4931) <= not (a and b);
    layer1_outputs(4932) <= '1';
    layer1_outputs(4933) <= b;
    layer1_outputs(4934) <= a or b;
    layer1_outputs(4935) <= a xor b;
    layer1_outputs(4936) <= a and not b;
    layer1_outputs(4937) <= not (a and b);
    layer1_outputs(4938) <= not (a xor b);
    layer1_outputs(4939) <= a and not b;
    layer1_outputs(4940) <= a and b;
    layer1_outputs(4941) <= a and not b;
    layer1_outputs(4942) <= not a or b;
    layer1_outputs(4943) <= a and not b;
    layer1_outputs(4944) <= not a;
    layer1_outputs(4945) <= '0';
    layer1_outputs(4946) <= not b or a;
    layer1_outputs(4947) <= not a;
    layer1_outputs(4948) <= not (a xor b);
    layer1_outputs(4949) <= not b or a;
    layer1_outputs(4950) <= b and not a;
    layer1_outputs(4951) <= a;
    layer1_outputs(4952) <= a and not b;
    layer1_outputs(4953) <= a and b;
    layer1_outputs(4954) <= not (a and b);
    layer1_outputs(4955) <= not a;
    layer1_outputs(4956) <= '0';
    layer1_outputs(4957) <= b;
    layer1_outputs(4958) <= a and b;
    layer1_outputs(4959) <= '0';
    layer1_outputs(4960) <= '0';
    layer1_outputs(4961) <= a and not b;
    layer1_outputs(4962) <= a and not b;
    layer1_outputs(4963) <= not a or b;
    layer1_outputs(4964) <= not (a and b);
    layer1_outputs(4965) <= b and not a;
    layer1_outputs(4966) <= not a or b;
    layer1_outputs(4967) <= not (a and b);
    layer1_outputs(4968) <= not a;
    layer1_outputs(4969) <= not b;
    layer1_outputs(4970) <= a or b;
    layer1_outputs(4971) <= not (a and b);
    layer1_outputs(4972) <= not (a and b);
    layer1_outputs(4973) <= not a or b;
    layer1_outputs(4974) <= b and not a;
    layer1_outputs(4975) <= not (a and b);
    layer1_outputs(4976) <= not a or b;
    layer1_outputs(4977) <= a;
    layer1_outputs(4978) <= a;
    layer1_outputs(4979) <= a xor b;
    layer1_outputs(4980) <= a and not b;
    layer1_outputs(4981) <= a or b;
    layer1_outputs(4982) <= b;
    layer1_outputs(4983) <= a and not b;
    layer1_outputs(4984) <= not (a or b);
    layer1_outputs(4985) <= a and b;
    layer1_outputs(4986) <= a;
    layer1_outputs(4987) <= a;
    layer1_outputs(4988) <= not b;
    layer1_outputs(4989) <= a;
    layer1_outputs(4990) <= not b;
    layer1_outputs(4991) <= not b;
    layer1_outputs(4992) <= b and not a;
    layer1_outputs(4993) <= not (a and b);
    layer1_outputs(4994) <= b;
    layer1_outputs(4995) <= a and not b;
    layer1_outputs(4996) <= a;
    layer1_outputs(4997) <= a;
    layer1_outputs(4998) <= a and not b;
    layer1_outputs(4999) <= a;
    layer1_outputs(5000) <= b and not a;
    layer1_outputs(5001) <= not a;
    layer1_outputs(5002) <= not b;
    layer1_outputs(5003) <= not a or b;
    layer1_outputs(5004) <= not (a xor b);
    layer1_outputs(5005) <= a;
    layer1_outputs(5006) <= a or b;
    layer1_outputs(5007) <= a;
    layer1_outputs(5008) <= not a;
    layer1_outputs(5009) <= not b;
    layer1_outputs(5010) <= '0';
    layer1_outputs(5011) <= a and b;
    layer1_outputs(5012) <= not b or a;
    layer1_outputs(5013) <= a;
    layer1_outputs(5014) <= not b or a;
    layer1_outputs(5015) <= not b or a;
    layer1_outputs(5016) <= not a;
    layer1_outputs(5017) <= '0';
    layer1_outputs(5018) <= b and not a;
    layer1_outputs(5019) <= a;
    layer1_outputs(5020) <= not a or b;
    layer1_outputs(5021) <= a and b;
    layer1_outputs(5022) <= not b;
    layer1_outputs(5023) <= b and not a;
    layer1_outputs(5024) <= b and not a;
    layer1_outputs(5025) <= a or b;
    layer1_outputs(5026) <= '0';
    layer1_outputs(5027) <= b and not a;
    layer1_outputs(5028) <= a and b;
    layer1_outputs(5029) <= '0';
    layer1_outputs(5030) <= a;
    layer1_outputs(5031) <= not (a xor b);
    layer1_outputs(5032) <= a;
    layer1_outputs(5033) <= a and b;
    layer1_outputs(5034) <= not (a or b);
    layer1_outputs(5035) <= b;
    layer1_outputs(5036) <= not (a and b);
    layer1_outputs(5037) <= not (a or b);
    layer1_outputs(5038) <= a and b;
    layer1_outputs(5039) <= '0';
    layer1_outputs(5040) <= not b;
    layer1_outputs(5041) <= not (a and b);
    layer1_outputs(5042) <= not a or b;
    layer1_outputs(5043) <= a and not b;
    layer1_outputs(5044) <= not b;
    layer1_outputs(5045) <= a and not b;
    layer1_outputs(5046) <= a and not b;
    layer1_outputs(5047) <= a;
    layer1_outputs(5048) <= b;
    layer1_outputs(5049) <= b and not a;
    layer1_outputs(5050) <= '0';
    layer1_outputs(5051) <= a and b;
    layer1_outputs(5052) <= not (a and b);
    layer1_outputs(5053) <= not (a xor b);
    layer1_outputs(5054) <= not (a or b);
    layer1_outputs(5055) <= a and not b;
    layer1_outputs(5056) <= b and not a;
    layer1_outputs(5057) <= a and b;
    layer1_outputs(5058) <= a or b;
    layer1_outputs(5059) <= not b;
    layer1_outputs(5060) <= not (a or b);
    layer1_outputs(5061) <= not b;
    layer1_outputs(5062) <= a xor b;
    layer1_outputs(5063) <= not a;
    layer1_outputs(5064) <= not (a or b);
    layer1_outputs(5065) <= a;
    layer1_outputs(5066) <= not b or a;
    layer1_outputs(5067) <= not b;
    layer1_outputs(5068) <= a or b;
    layer1_outputs(5069) <= not (a and b);
    layer1_outputs(5070) <= not a or b;
    layer1_outputs(5071) <= not a;
    layer1_outputs(5072) <= not a or b;
    layer1_outputs(5073) <= not (a or b);
    layer1_outputs(5074) <= a and b;
    layer1_outputs(5075) <= '1';
    layer1_outputs(5076) <= b;
    layer1_outputs(5077) <= not b;
    layer1_outputs(5078) <= a and b;
    layer1_outputs(5079) <= a;
    layer1_outputs(5080) <= not b or a;
    layer1_outputs(5081) <= b and not a;
    layer1_outputs(5082) <= b;
    layer1_outputs(5083) <= a and b;
    layer1_outputs(5084) <= a or b;
    layer1_outputs(5085) <= not a;
    layer1_outputs(5086) <= a;
    layer1_outputs(5087) <= a and not b;
    layer1_outputs(5088) <= b;
    layer1_outputs(5089) <= a xor b;
    layer1_outputs(5090) <= a;
    layer1_outputs(5091) <= not b or a;
    layer1_outputs(5092) <= a;
    layer1_outputs(5093) <= not b or a;
    layer1_outputs(5094) <= a and not b;
    layer1_outputs(5095) <= not a or b;
    layer1_outputs(5096) <= not b;
    layer1_outputs(5097) <= a or b;
    layer1_outputs(5098) <= not (a or b);
    layer1_outputs(5099) <= a and not b;
    layer1_outputs(5100) <= a and b;
    layer1_outputs(5101) <= a xor b;
    layer1_outputs(5102) <= not b;
    layer1_outputs(5103) <= a or b;
    layer1_outputs(5104) <= '1';
    layer1_outputs(5105) <= a and not b;
    layer1_outputs(5106) <= a;
    layer1_outputs(5107) <= a and not b;
    layer1_outputs(5108) <= not (a and b);
    layer1_outputs(5109) <= b;
    layer1_outputs(5110) <= b;
    layer1_outputs(5111) <= not (a or b);
    layer1_outputs(5112) <= not a or b;
    layer1_outputs(5113) <= not (a and b);
    layer1_outputs(5114) <= not a;
    layer1_outputs(5115) <= not b or a;
    layer1_outputs(5116) <= b and not a;
    layer1_outputs(5117) <= '1';
    layer1_outputs(5118) <= not a or b;
    layer1_outputs(5119) <= '0';
    layer2_outputs(0) <= not a;
    layer2_outputs(1) <= b;
    layer2_outputs(2) <= '1';
    layer2_outputs(3) <= not b or a;
    layer2_outputs(4) <= a;
    layer2_outputs(5) <= b and not a;
    layer2_outputs(6) <= b and not a;
    layer2_outputs(7) <= b and not a;
    layer2_outputs(8) <= not b;
    layer2_outputs(9) <= not a;
    layer2_outputs(10) <= not b;
    layer2_outputs(11) <= a or b;
    layer2_outputs(12) <= not a;
    layer2_outputs(13) <= not a;
    layer2_outputs(14) <= not a or b;
    layer2_outputs(15) <= a;
    layer2_outputs(16) <= not (a and b);
    layer2_outputs(17) <= not a;
    layer2_outputs(18) <= a xor b;
    layer2_outputs(19) <= a;
    layer2_outputs(20) <= not (a or b);
    layer2_outputs(21) <= not (a or b);
    layer2_outputs(22) <= a and not b;
    layer2_outputs(23) <= b;
    layer2_outputs(24) <= not a or b;
    layer2_outputs(25) <= not (a xor b);
    layer2_outputs(26) <= '0';
    layer2_outputs(27) <= not (a or b);
    layer2_outputs(28) <= a xor b;
    layer2_outputs(29) <= b;
    layer2_outputs(30) <= a and not b;
    layer2_outputs(31) <= not (a and b);
    layer2_outputs(32) <= a or b;
    layer2_outputs(33) <= a;
    layer2_outputs(34) <= a;
    layer2_outputs(35) <= a and b;
    layer2_outputs(36) <= not (a and b);
    layer2_outputs(37) <= not b or a;
    layer2_outputs(38) <= not a;
    layer2_outputs(39) <= not b or a;
    layer2_outputs(40) <= not (a xor b);
    layer2_outputs(41) <= not a;
    layer2_outputs(42) <= a;
    layer2_outputs(43) <= not a or b;
    layer2_outputs(44) <= a and b;
    layer2_outputs(45) <= b;
    layer2_outputs(46) <= not a;
    layer2_outputs(47) <= not (a or b);
    layer2_outputs(48) <= a and not b;
    layer2_outputs(49) <= not b;
    layer2_outputs(50) <= not (a or b);
    layer2_outputs(51) <= not b or a;
    layer2_outputs(52) <= a;
    layer2_outputs(53) <= not (a and b);
    layer2_outputs(54) <= a;
    layer2_outputs(55) <= not (a xor b);
    layer2_outputs(56) <= not a or b;
    layer2_outputs(57) <= not a;
    layer2_outputs(58) <= b;
    layer2_outputs(59) <= a and b;
    layer2_outputs(60) <= b;
    layer2_outputs(61) <= a and b;
    layer2_outputs(62) <= not b or a;
    layer2_outputs(63) <= not (a or b);
    layer2_outputs(64) <= not b or a;
    layer2_outputs(65) <= a and not b;
    layer2_outputs(66) <= not (a and b);
    layer2_outputs(67) <= a;
    layer2_outputs(68) <= not b;
    layer2_outputs(69) <= b and not a;
    layer2_outputs(70) <= '0';
    layer2_outputs(71) <= not (a or b);
    layer2_outputs(72) <= a;
    layer2_outputs(73) <= b;
    layer2_outputs(74) <= '0';
    layer2_outputs(75) <= not b;
    layer2_outputs(76) <= not b;
    layer2_outputs(77) <= not b or a;
    layer2_outputs(78) <= a;
    layer2_outputs(79) <= a or b;
    layer2_outputs(80) <= b;
    layer2_outputs(81) <= b;
    layer2_outputs(82) <= a or b;
    layer2_outputs(83) <= not a or b;
    layer2_outputs(84) <= b;
    layer2_outputs(85) <= not b;
    layer2_outputs(86) <= a;
    layer2_outputs(87) <= not (a or b);
    layer2_outputs(88) <= a;
    layer2_outputs(89) <= b;
    layer2_outputs(90) <= a;
    layer2_outputs(91) <= not b;
    layer2_outputs(92) <= a;
    layer2_outputs(93) <= not (a or b);
    layer2_outputs(94) <= a xor b;
    layer2_outputs(95) <= not a or b;
    layer2_outputs(96) <= b;
    layer2_outputs(97) <= a xor b;
    layer2_outputs(98) <= b;
    layer2_outputs(99) <= a;
    layer2_outputs(100) <= a and not b;
    layer2_outputs(101) <= not b;
    layer2_outputs(102) <= not (a or b);
    layer2_outputs(103) <= not a;
    layer2_outputs(104) <= a or b;
    layer2_outputs(105) <= not a or b;
    layer2_outputs(106) <= not a or b;
    layer2_outputs(107) <= '1';
    layer2_outputs(108) <= b and not a;
    layer2_outputs(109) <= not b;
    layer2_outputs(110) <= not a;
    layer2_outputs(111) <= not (a and b);
    layer2_outputs(112) <= a;
    layer2_outputs(113) <= a;
    layer2_outputs(114) <= a or b;
    layer2_outputs(115) <= a;
    layer2_outputs(116) <= a xor b;
    layer2_outputs(117) <= not a or b;
    layer2_outputs(118) <= a and not b;
    layer2_outputs(119) <= a and not b;
    layer2_outputs(120) <= b;
    layer2_outputs(121) <= a and not b;
    layer2_outputs(122) <= b;
    layer2_outputs(123) <= not b or a;
    layer2_outputs(124) <= not b or a;
    layer2_outputs(125) <= not b;
    layer2_outputs(126) <= b and not a;
    layer2_outputs(127) <= b;
    layer2_outputs(128) <= a xor b;
    layer2_outputs(129) <= a;
    layer2_outputs(130) <= not (a xor b);
    layer2_outputs(131) <= not a or b;
    layer2_outputs(132) <= a xor b;
    layer2_outputs(133) <= a and not b;
    layer2_outputs(134) <= b;
    layer2_outputs(135) <= not b or a;
    layer2_outputs(136) <= not a;
    layer2_outputs(137) <= b and not a;
    layer2_outputs(138) <= not b;
    layer2_outputs(139) <= a;
    layer2_outputs(140) <= a and not b;
    layer2_outputs(141) <= a xor b;
    layer2_outputs(142) <= a;
    layer2_outputs(143) <= not a;
    layer2_outputs(144) <= not b;
    layer2_outputs(145) <= a and b;
    layer2_outputs(146) <= b;
    layer2_outputs(147) <= not b;
    layer2_outputs(148) <= a xor b;
    layer2_outputs(149) <= not b;
    layer2_outputs(150) <= not b;
    layer2_outputs(151) <= not (a xor b);
    layer2_outputs(152) <= not b or a;
    layer2_outputs(153) <= not (a or b);
    layer2_outputs(154) <= '1';
    layer2_outputs(155) <= a and b;
    layer2_outputs(156) <= a or b;
    layer2_outputs(157) <= a xor b;
    layer2_outputs(158) <= a or b;
    layer2_outputs(159) <= a and b;
    layer2_outputs(160) <= not a;
    layer2_outputs(161) <= a or b;
    layer2_outputs(162) <= b;
    layer2_outputs(163) <= not (a xor b);
    layer2_outputs(164) <= b;
    layer2_outputs(165) <= not (a and b);
    layer2_outputs(166) <= not (a and b);
    layer2_outputs(167) <= a;
    layer2_outputs(168) <= a or b;
    layer2_outputs(169) <= b and not a;
    layer2_outputs(170) <= not (a and b);
    layer2_outputs(171) <= a;
    layer2_outputs(172) <= not (a or b);
    layer2_outputs(173) <= not a or b;
    layer2_outputs(174) <= a;
    layer2_outputs(175) <= a or b;
    layer2_outputs(176) <= a or b;
    layer2_outputs(177) <= not a;
    layer2_outputs(178) <= b and not a;
    layer2_outputs(179) <= b;
    layer2_outputs(180) <= not a;
    layer2_outputs(181) <= b;
    layer2_outputs(182) <= not b or a;
    layer2_outputs(183) <= not (a or b);
    layer2_outputs(184) <= b;
    layer2_outputs(185) <= a;
    layer2_outputs(186) <= not (a or b);
    layer2_outputs(187) <= not a;
    layer2_outputs(188) <= not (a and b);
    layer2_outputs(189) <= a and not b;
    layer2_outputs(190) <= not b;
    layer2_outputs(191) <= not (a and b);
    layer2_outputs(192) <= not (a and b);
    layer2_outputs(193) <= a or b;
    layer2_outputs(194) <= not (a and b);
    layer2_outputs(195) <= b;
    layer2_outputs(196) <= not b or a;
    layer2_outputs(197) <= a;
    layer2_outputs(198) <= not (a or b);
    layer2_outputs(199) <= a;
    layer2_outputs(200) <= not a or b;
    layer2_outputs(201) <= b and not a;
    layer2_outputs(202) <= not a;
    layer2_outputs(203) <= not b;
    layer2_outputs(204) <= not (a and b);
    layer2_outputs(205) <= a and not b;
    layer2_outputs(206) <= not b or a;
    layer2_outputs(207) <= a;
    layer2_outputs(208) <= a and b;
    layer2_outputs(209) <= not a;
    layer2_outputs(210) <= not a or b;
    layer2_outputs(211) <= not b or a;
    layer2_outputs(212) <= a and not b;
    layer2_outputs(213) <= not b or a;
    layer2_outputs(214) <= b and not a;
    layer2_outputs(215) <= a;
    layer2_outputs(216) <= not a;
    layer2_outputs(217) <= a;
    layer2_outputs(218) <= a;
    layer2_outputs(219) <= b;
    layer2_outputs(220) <= not b;
    layer2_outputs(221) <= '1';
    layer2_outputs(222) <= b;
    layer2_outputs(223) <= not (a and b);
    layer2_outputs(224) <= b;
    layer2_outputs(225) <= a;
    layer2_outputs(226) <= a xor b;
    layer2_outputs(227) <= not (a and b);
    layer2_outputs(228) <= a and b;
    layer2_outputs(229) <= not a;
    layer2_outputs(230) <= not (a or b);
    layer2_outputs(231) <= not a or b;
    layer2_outputs(232) <= not (a or b);
    layer2_outputs(233) <= b;
    layer2_outputs(234) <= b;
    layer2_outputs(235) <= not b;
    layer2_outputs(236) <= a xor b;
    layer2_outputs(237) <= not a;
    layer2_outputs(238) <= not a;
    layer2_outputs(239) <= not a;
    layer2_outputs(240) <= not a;
    layer2_outputs(241) <= not a;
    layer2_outputs(242) <= not (a or b);
    layer2_outputs(243) <= b;
    layer2_outputs(244) <= a xor b;
    layer2_outputs(245) <= not b or a;
    layer2_outputs(246) <= not b;
    layer2_outputs(247) <= not (a and b);
    layer2_outputs(248) <= a;
    layer2_outputs(249) <= not b or a;
    layer2_outputs(250) <= not b;
    layer2_outputs(251) <= not (a and b);
    layer2_outputs(252) <= a;
    layer2_outputs(253) <= not (a or b);
    layer2_outputs(254) <= a xor b;
    layer2_outputs(255) <= a;
    layer2_outputs(256) <= not (a or b);
    layer2_outputs(257) <= a or b;
    layer2_outputs(258) <= a or b;
    layer2_outputs(259) <= a or b;
    layer2_outputs(260) <= a;
    layer2_outputs(261) <= not a or b;
    layer2_outputs(262) <= a xor b;
    layer2_outputs(263) <= not b or a;
    layer2_outputs(264) <= b;
    layer2_outputs(265) <= a and not b;
    layer2_outputs(266) <= not b;
    layer2_outputs(267) <= a and b;
    layer2_outputs(268) <= not b;
    layer2_outputs(269) <= a and b;
    layer2_outputs(270) <= not b;
    layer2_outputs(271) <= not b;
    layer2_outputs(272) <= not a or b;
    layer2_outputs(273) <= b and not a;
    layer2_outputs(274) <= not (a and b);
    layer2_outputs(275) <= b;
    layer2_outputs(276) <= a;
    layer2_outputs(277) <= not (a and b);
    layer2_outputs(278) <= not (a or b);
    layer2_outputs(279) <= a;
    layer2_outputs(280) <= not b;
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= a xor b;
    layer2_outputs(283) <= not b or a;
    layer2_outputs(284) <= a or b;
    layer2_outputs(285) <= not b or a;
    layer2_outputs(286) <= not a or b;
    layer2_outputs(287) <= b and not a;
    layer2_outputs(288) <= not (a xor b);
    layer2_outputs(289) <= b and not a;
    layer2_outputs(290) <= not b;
    layer2_outputs(291) <= not a;
    layer2_outputs(292) <= a;
    layer2_outputs(293) <= not a or b;
    layer2_outputs(294) <= not a or b;
    layer2_outputs(295) <= not b;
    layer2_outputs(296) <= not b;
    layer2_outputs(297) <= '0';
    layer2_outputs(298) <= a;
    layer2_outputs(299) <= not (a and b);
    layer2_outputs(300) <= not (a xor b);
    layer2_outputs(301) <= not a or b;
    layer2_outputs(302) <= b;
    layer2_outputs(303) <= not (a or b);
    layer2_outputs(304) <= not (a xor b);
    layer2_outputs(305) <= a and not b;
    layer2_outputs(306) <= not a;
    layer2_outputs(307) <= not a;
    layer2_outputs(308) <= not (a and b);
    layer2_outputs(309) <= b;
    layer2_outputs(310) <= a or b;
    layer2_outputs(311) <= not b;
    layer2_outputs(312) <= not a;
    layer2_outputs(313) <= not b or a;
    layer2_outputs(314) <= not (a and b);
    layer2_outputs(315) <= a;
    layer2_outputs(316) <= not a;
    layer2_outputs(317) <= a or b;
    layer2_outputs(318) <= not b or a;
    layer2_outputs(319) <= not (a and b);
    layer2_outputs(320) <= not (a or b);
    layer2_outputs(321) <= not a;
    layer2_outputs(322) <= a;
    layer2_outputs(323) <= b and not a;
    layer2_outputs(324) <= not a or b;
    layer2_outputs(325) <= not b or a;
    layer2_outputs(326) <= not (a or b);
    layer2_outputs(327) <= a and not b;
    layer2_outputs(328) <= not b;
    layer2_outputs(329) <= not (a or b);
    layer2_outputs(330) <= b;
    layer2_outputs(331) <= b and not a;
    layer2_outputs(332) <= b;
    layer2_outputs(333) <= not (a and b);
    layer2_outputs(334) <= not a;
    layer2_outputs(335) <= a and b;
    layer2_outputs(336) <= not b;
    layer2_outputs(337) <= not a;
    layer2_outputs(338) <= not b;
    layer2_outputs(339) <= not (a or b);
    layer2_outputs(340) <= b and not a;
    layer2_outputs(341) <= not b or a;
    layer2_outputs(342) <= a and not b;
    layer2_outputs(343) <= b;
    layer2_outputs(344) <= '1';
    layer2_outputs(345) <= a or b;
    layer2_outputs(346) <= not b;
    layer2_outputs(347) <= not (a xor b);
    layer2_outputs(348) <= b;
    layer2_outputs(349) <= not b;
    layer2_outputs(350) <= not a or b;
    layer2_outputs(351) <= '1';
    layer2_outputs(352) <= not b or a;
    layer2_outputs(353) <= not (a or b);
    layer2_outputs(354) <= not b;
    layer2_outputs(355) <= not b;
    layer2_outputs(356) <= a and not b;
    layer2_outputs(357) <= b;
    layer2_outputs(358) <= a and b;
    layer2_outputs(359) <= not b or a;
    layer2_outputs(360) <= not a or b;
    layer2_outputs(361) <= not a or b;
    layer2_outputs(362) <= a;
    layer2_outputs(363) <= not a or b;
    layer2_outputs(364) <= b;
    layer2_outputs(365) <= not (a and b);
    layer2_outputs(366) <= '1';
    layer2_outputs(367) <= a or b;
    layer2_outputs(368) <= not a or b;
    layer2_outputs(369) <= '1';
    layer2_outputs(370) <= not (a and b);
    layer2_outputs(371) <= not b;
    layer2_outputs(372) <= a and not b;
    layer2_outputs(373) <= not (a xor b);
    layer2_outputs(374) <= not b;
    layer2_outputs(375) <= not a;
    layer2_outputs(376) <= not b;
    layer2_outputs(377) <= b;
    layer2_outputs(378) <= not b or a;
    layer2_outputs(379) <= b and not a;
    layer2_outputs(380) <= a or b;
    layer2_outputs(381) <= not (a or b);
    layer2_outputs(382) <= not a;
    layer2_outputs(383) <= a;
    layer2_outputs(384) <= not a;
    layer2_outputs(385) <= not a;
    layer2_outputs(386) <= a xor b;
    layer2_outputs(387) <= not a or b;
    layer2_outputs(388) <= b and not a;
    layer2_outputs(389) <= not a;
    layer2_outputs(390) <= b and not a;
    layer2_outputs(391) <= a;
    layer2_outputs(392) <= '1';
    layer2_outputs(393) <= a or b;
    layer2_outputs(394) <= a;
    layer2_outputs(395) <= not (a xor b);
    layer2_outputs(396) <= not a;
    layer2_outputs(397) <= a;
    layer2_outputs(398) <= a and b;
    layer2_outputs(399) <= not b;
    layer2_outputs(400) <= not (a or b);
    layer2_outputs(401) <= not b or a;
    layer2_outputs(402) <= b;
    layer2_outputs(403) <= a and not b;
    layer2_outputs(404) <= b;
    layer2_outputs(405) <= b;
    layer2_outputs(406) <= '0';
    layer2_outputs(407) <= not a;
    layer2_outputs(408) <= not (a or b);
    layer2_outputs(409) <= a and not b;
    layer2_outputs(410) <= not a or b;
    layer2_outputs(411) <= not a;
    layer2_outputs(412) <= not a or b;
    layer2_outputs(413) <= not b;
    layer2_outputs(414) <= not (a or b);
    layer2_outputs(415) <= b;
    layer2_outputs(416) <= not a;
    layer2_outputs(417) <= not (a or b);
    layer2_outputs(418) <= a or b;
    layer2_outputs(419) <= not b or a;
    layer2_outputs(420) <= b;
    layer2_outputs(421) <= not b or a;
    layer2_outputs(422) <= not a or b;
    layer2_outputs(423) <= b;
    layer2_outputs(424) <= a or b;
    layer2_outputs(425) <= '1';
    layer2_outputs(426) <= '1';
    layer2_outputs(427) <= a and not b;
    layer2_outputs(428) <= '1';
    layer2_outputs(429) <= a or b;
    layer2_outputs(430) <= b;
    layer2_outputs(431) <= '0';
    layer2_outputs(432) <= not a or b;
    layer2_outputs(433) <= a and b;
    layer2_outputs(434) <= a or b;
    layer2_outputs(435) <= a and b;
    layer2_outputs(436) <= a;
    layer2_outputs(437) <= a and not b;
    layer2_outputs(438) <= not (a and b);
    layer2_outputs(439) <= not b or a;
    layer2_outputs(440) <= a or b;
    layer2_outputs(441) <= a and not b;
    layer2_outputs(442) <= a and b;
    layer2_outputs(443) <= a;
    layer2_outputs(444) <= not a or b;
    layer2_outputs(445) <= not (a xor b);
    layer2_outputs(446) <= not b;
    layer2_outputs(447) <= not a;
    layer2_outputs(448) <= '0';
    layer2_outputs(449) <= not (a and b);
    layer2_outputs(450) <= not b;
    layer2_outputs(451) <= a;
    layer2_outputs(452) <= a and not b;
    layer2_outputs(453) <= not b;
    layer2_outputs(454) <= a or b;
    layer2_outputs(455) <= a;
    layer2_outputs(456) <= a and not b;
    layer2_outputs(457) <= a and b;
    layer2_outputs(458) <= not a or b;
    layer2_outputs(459) <= a and not b;
    layer2_outputs(460) <= a and b;
    layer2_outputs(461) <= not a or b;
    layer2_outputs(462) <= not b;
    layer2_outputs(463) <= not (a and b);
    layer2_outputs(464) <= not (a or b);
    layer2_outputs(465) <= not b;
    layer2_outputs(466) <= a or b;
    layer2_outputs(467) <= not (a xor b);
    layer2_outputs(468) <= not a or b;
    layer2_outputs(469) <= '0';
    layer2_outputs(470) <= not a or b;
    layer2_outputs(471) <= a;
    layer2_outputs(472) <= not (a or b);
    layer2_outputs(473) <= a and not b;
    layer2_outputs(474) <= a;
    layer2_outputs(475) <= not (a and b);
    layer2_outputs(476) <= a and b;
    layer2_outputs(477) <= not b;
    layer2_outputs(478) <= b and not a;
    layer2_outputs(479) <= '0';
    layer2_outputs(480) <= not (a or b);
    layer2_outputs(481) <= a and not b;
    layer2_outputs(482) <= b;
    layer2_outputs(483) <= a;
    layer2_outputs(484) <= not (a and b);
    layer2_outputs(485) <= a and not b;
    layer2_outputs(486) <= not a or b;
    layer2_outputs(487) <= '1';
    layer2_outputs(488) <= a and not b;
    layer2_outputs(489) <= a and b;
    layer2_outputs(490) <= b and not a;
    layer2_outputs(491) <= b and not a;
    layer2_outputs(492) <= a and b;
    layer2_outputs(493) <= not a;
    layer2_outputs(494) <= not b;
    layer2_outputs(495) <= a;
    layer2_outputs(496) <= b and not a;
    layer2_outputs(497) <= a or b;
    layer2_outputs(498) <= b;
    layer2_outputs(499) <= a and b;
    layer2_outputs(500) <= a or b;
    layer2_outputs(501) <= '1';
    layer2_outputs(502) <= not a;
    layer2_outputs(503) <= not (a and b);
    layer2_outputs(504) <= not a;
    layer2_outputs(505) <= not b;
    layer2_outputs(506) <= not a or b;
    layer2_outputs(507) <= b;
    layer2_outputs(508) <= not b;
    layer2_outputs(509) <= not b;
    layer2_outputs(510) <= a or b;
    layer2_outputs(511) <= b;
    layer2_outputs(512) <= a or b;
    layer2_outputs(513) <= a and b;
    layer2_outputs(514) <= a xor b;
    layer2_outputs(515) <= '1';
    layer2_outputs(516) <= not a;
    layer2_outputs(517) <= b;
    layer2_outputs(518) <= not a or b;
    layer2_outputs(519) <= '0';
    layer2_outputs(520) <= not (a and b);
    layer2_outputs(521) <= not (a or b);
    layer2_outputs(522) <= b and not a;
    layer2_outputs(523) <= b;
    layer2_outputs(524) <= not (a and b);
    layer2_outputs(525) <= a or b;
    layer2_outputs(526) <= not a or b;
    layer2_outputs(527) <= '1';
    layer2_outputs(528) <= b;
    layer2_outputs(529) <= not (a or b);
    layer2_outputs(530) <= not b or a;
    layer2_outputs(531) <= b;
    layer2_outputs(532) <= not (a and b);
    layer2_outputs(533) <= not (a and b);
    layer2_outputs(534) <= a;
    layer2_outputs(535) <= not (a xor b);
    layer2_outputs(536) <= a or b;
    layer2_outputs(537) <= not a;
    layer2_outputs(538) <= '0';
    layer2_outputs(539) <= not a or b;
    layer2_outputs(540) <= a;
    layer2_outputs(541) <= not (a and b);
    layer2_outputs(542) <= b and not a;
    layer2_outputs(543) <= not (a or b);
    layer2_outputs(544) <= a;
    layer2_outputs(545) <= a and b;
    layer2_outputs(546) <= not (a xor b);
    layer2_outputs(547) <= b;
    layer2_outputs(548) <= b;
    layer2_outputs(549) <= b;
    layer2_outputs(550) <= a and b;
    layer2_outputs(551) <= a and not b;
    layer2_outputs(552) <= not a;
    layer2_outputs(553) <= a or b;
    layer2_outputs(554) <= not b;
    layer2_outputs(555) <= not (a or b);
    layer2_outputs(556) <= b;
    layer2_outputs(557) <= a or b;
    layer2_outputs(558) <= not a;
    layer2_outputs(559) <= b;
    layer2_outputs(560) <= not a or b;
    layer2_outputs(561) <= not (a or b);
    layer2_outputs(562) <= a;
    layer2_outputs(563) <= b;
    layer2_outputs(564) <= b;
    layer2_outputs(565) <= not b or a;
    layer2_outputs(566) <= not b or a;
    layer2_outputs(567) <= not b;
    layer2_outputs(568) <= '1';
    layer2_outputs(569) <= a and not b;
    layer2_outputs(570) <= not (a xor b);
    layer2_outputs(571) <= not (a or b);
    layer2_outputs(572) <= not a or b;
    layer2_outputs(573) <= not (a xor b);
    layer2_outputs(574) <= a and not b;
    layer2_outputs(575) <= a;
    layer2_outputs(576) <= not b;
    layer2_outputs(577) <= a or b;
    layer2_outputs(578) <= b;
    layer2_outputs(579) <= not b or a;
    layer2_outputs(580) <= b and not a;
    layer2_outputs(581) <= a and not b;
    layer2_outputs(582) <= not a;
    layer2_outputs(583) <= '0';
    layer2_outputs(584) <= not (a or b);
    layer2_outputs(585) <= '1';
    layer2_outputs(586) <= '0';
    layer2_outputs(587) <= b and not a;
    layer2_outputs(588) <= not a;
    layer2_outputs(589) <= a or b;
    layer2_outputs(590) <= not a;
    layer2_outputs(591) <= '1';
    layer2_outputs(592) <= not (a or b);
    layer2_outputs(593) <= b and not a;
    layer2_outputs(594) <= a and b;
    layer2_outputs(595) <= not (a and b);
    layer2_outputs(596) <= not b;
    layer2_outputs(597) <= not a or b;
    layer2_outputs(598) <= '0';
    layer2_outputs(599) <= a and not b;
    layer2_outputs(600) <= '0';
    layer2_outputs(601) <= a and not b;
    layer2_outputs(602) <= a;
    layer2_outputs(603) <= b and not a;
    layer2_outputs(604) <= not (a or b);
    layer2_outputs(605) <= b;
    layer2_outputs(606) <= '0';
    layer2_outputs(607) <= '0';
    layer2_outputs(608) <= a xor b;
    layer2_outputs(609) <= not (a and b);
    layer2_outputs(610) <= a or b;
    layer2_outputs(611) <= not (a xor b);
    layer2_outputs(612) <= a and not b;
    layer2_outputs(613) <= a and not b;
    layer2_outputs(614) <= not (a and b);
    layer2_outputs(615) <= not (a xor b);
    layer2_outputs(616) <= not a or b;
    layer2_outputs(617) <= not (a and b);
    layer2_outputs(618) <= not b or a;
    layer2_outputs(619) <= a or b;
    layer2_outputs(620) <= a and b;
    layer2_outputs(621) <= b;
    layer2_outputs(622) <= not a or b;
    layer2_outputs(623) <= b;
    layer2_outputs(624) <= not (a xor b);
    layer2_outputs(625) <= not a;
    layer2_outputs(626) <= '1';
    layer2_outputs(627) <= not a or b;
    layer2_outputs(628) <= not (a or b);
    layer2_outputs(629) <= a and not b;
    layer2_outputs(630) <= b;
    layer2_outputs(631) <= not a;
    layer2_outputs(632) <= a or b;
    layer2_outputs(633) <= not b;
    layer2_outputs(634) <= a;
    layer2_outputs(635) <= a and b;
    layer2_outputs(636) <= not a or b;
    layer2_outputs(637) <= not a;
    layer2_outputs(638) <= a;
    layer2_outputs(639) <= a and not b;
    layer2_outputs(640) <= not b or a;
    layer2_outputs(641) <= b;
    layer2_outputs(642) <= b;
    layer2_outputs(643) <= not a or b;
    layer2_outputs(644) <= b and not a;
    layer2_outputs(645) <= not b or a;
    layer2_outputs(646) <= a and b;
    layer2_outputs(647) <= '0';
    layer2_outputs(648) <= not b;
    layer2_outputs(649) <= a or b;
    layer2_outputs(650) <= not a or b;
    layer2_outputs(651) <= b;
    layer2_outputs(652) <= a and not b;
    layer2_outputs(653) <= not a;
    layer2_outputs(654) <= not (a xor b);
    layer2_outputs(655) <= not a;
    layer2_outputs(656) <= not a or b;
    layer2_outputs(657) <= not b;
    layer2_outputs(658) <= '0';
    layer2_outputs(659) <= a and not b;
    layer2_outputs(660) <= b;
    layer2_outputs(661) <= a;
    layer2_outputs(662) <= b;
    layer2_outputs(663) <= a and not b;
    layer2_outputs(664) <= not (a or b);
    layer2_outputs(665) <= a and not b;
    layer2_outputs(666) <= a and b;
    layer2_outputs(667) <= a and not b;
    layer2_outputs(668) <= not a;
    layer2_outputs(669) <= not (a and b);
    layer2_outputs(670) <= not (a and b);
    layer2_outputs(671) <= b;
    layer2_outputs(672) <= not a;
    layer2_outputs(673) <= not a or b;
    layer2_outputs(674) <= not a or b;
    layer2_outputs(675) <= not a or b;
    layer2_outputs(676) <= not a;
    layer2_outputs(677) <= a and b;
    layer2_outputs(678) <= b;
    layer2_outputs(679) <= a or b;
    layer2_outputs(680) <= b;
    layer2_outputs(681) <= a or b;
    layer2_outputs(682) <= a and b;
    layer2_outputs(683) <= a;
    layer2_outputs(684) <= b;
    layer2_outputs(685) <= not (a and b);
    layer2_outputs(686) <= not b;
    layer2_outputs(687) <= a;
    layer2_outputs(688) <= b and not a;
    layer2_outputs(689) <= not b;
    layer2_outputs(690) <= a or b;
    layer2_outputs(691) <= not a;
    layer2_outputs(692) <= a and not b;
    layer2_outputs(693) <= not b;
    layer2_outputs(694) <= a and b;
    layer2_outputs(695) <= a and not b;
    layer2_outputs(696) <= not b;
    layer2_outputs(697) <= not (a or b);
    layer2_outputs(698) <= a or b;
    layer2_outputs(699) <= '0';
    layer2_outputs(700) <= '0';
    layer2_outputs(701) <= not (a and b);
    layer2_outputs(702) <= not a or b;
    layer2_outputs(703) <= not (a xor b);
    layer2_outputs(704) <= b;
    layer2_outputs(705) <= not a;
    layer2_outputs(706) <= not b or a;
    layer2_outputs(707) <= a or b;
    layer2_outputs(708) <= a or b;
    layer2_outputs(709) <= a and b;
    layer2_outputs(710) <= a and b;
    layer2_outputs(711) <= b;
    layer2_outputs(712) <= not (a and b);
    layer2_outputs(713) <= b;
    layer2_outputs(714) <= b and not a;
    layer2_outputs(715) <= a and b;
    layer2_outputs(716) <= not b;
    layer2_outputs(717) <= '1';
    layer2_outputs(718) <= a and b;
    layer2_outputs(719) <= a and not b;
    layer2_outputs(720) <= not (a and b);
    layer2_outputs(721) <= a or b;
    layer2_outputs(722) <= a and not b;
    layer2_outputs(723) <= a and b;
    layer2_outputs(724) <= not b or a;
    layer2_outputs(725) <= a;
    layer2_outputs(726) <= not (a xor b);
    layer2_outputs(727) <= not b;
    layer2_outputs(728) <= not (a and b);
    layer2_outputs(729) <= a;
    layer2_outputs(730) <= not (a or b);
    layer2_outputs(731) <= not (a or b);
    layer2_outputs(732) <= a xor b;
    layer2_outputs(733) <= not b;
    layer2_outputs(734) <= b;
    layer2_outputs(735) <= not (a xor b);
    layer2_outputs(736) <= not a;
    layer2_outputs(737) <= '1';
    layer2_outputs(738) <= b;
    layer2_outputs(739) <= not (a and b);
    layer2_outputs(740) <= a and not b;
    layer2_outputs(741) <= not a or b;
    layer2_outputs(742) <= not b;
    layer2_outputs(743) <= a;
    layer2_outputs(744) <= not a;
    layer2_outputs(745) <= not b;
    layer2_outputs(746) <= a and b;
    layer2_outputs(747) <= not a;
    layer2_outputs(748) <= b and not a;
    layer2_outputs(749) <= not a;
    layer2_outputs(750) <= b and not a;
    layer2_outputs(751) <= not (a or b);
    layer2_outputs(752) <= not (a and b);
    layer2_outputs(753) <= not (a xor b);
    layer2_outputs(754) <= not b or a;
    layer2_outputs(755) <= b and not a;
    layer2_outputs(756) <= '1';
    layer2_outputs(757) <= not b;
    layer2_outputs(758) <= not a;
    layer2_outputs(759) <= not (a or b);
    layer2_outputs(760) <= a;
    layer2_outputs(761) <= b and not a;
    layer2_outputs(762) <= b;
    layer2_outputs(763) <= a and not b;
    layer2_outputs(764) <= not b or a;
    layer2_outputs(765) <= a;
    layer2_outputs(766) <= a;
    layer2_outputs(767) <= b;
    layer2_outputs(768) <= b and not a;
    layer2_outputs(769) <= '1';
    layer2_outputs(770) <= a or b;
    layer2_outputs(771) <= not b or a;
    layer2_outputs(772) <= not (a xor b);
    layer2_outputs(773) <= not (a xor b);
    layer2_outputs(774) <= not (a xor b);
    layer2_outputs(775) <= not (a xor b);
    layer2_outputs(776) <= not a;
    layer2_outputs(777) <= a;
    layer2_outputs(778) <= a or b;
    layer2_outputs(779) <= not a;
    layer2_outputs(780) <= not b or a;
    layer2_outputs(781) <= a and b;
    layer2_outputs(782) <= not (a and b);
    layer2_outputs(783) <= b;
    layer2_outputs(784) <= a or b;
    layer2_outputs(785) <= b;
    layer2_outputs(786) <= a and not b;
    layer2_outputs(787) <= not (a and b);
    layer2_outputs(788) <= a xor b;
    layer2_outputs(789) <= not a;
    layer2_outputs(790) <= not (a and b);
    layer2_outputs(791) <= not a;
    layer2_outputs(792) <= a and b;
    layer2_outputs(793) <= not (a xor b);
    layer2_outputs(794) <= not (a and b);
    layer2_outputs(795) <= not b;
    layer2_outputs(796) <= not b or a;
    layer2_outputs(797) <= a and not b;
    layer2_outputs(798) <= '0';
    layer2_outputs(799) <= not a;
    layer2_outputs(800) <= b and not a;
    layer2_outputs(801) <= a;
    layer2_outputs(802) <= not a or b;
    layer2_outputs(803) <= not (a xor b);
    layer2_outputs(804) <= a and b;
    layer2_outputs(805) <= a or b;
    layer2_outputs(806) <= b;
    layer2_outputs(807) <= a;
    layer2_outputs(808) <= '0';
    layer2_outputs(809) <= not (a xor b);
    layer2_outputs(810) <= a;
    layer2_outputs(811) <= not (a and b);
    layer2_outputs(812) <= a xor b;
    layer2_outputs(813) <= not (a or b);
    layer2_outputs(814) <= a and not b;
    layer2_outputs(815) <= b;
    layer2_outputs(816) <= b;
    layer2_outputs(817) <= b and not a;
    layer2_outputs(818) <= not b or a;
    layer2_outputs(819) <= not (a xor b);
    layer2_outputs(820) <= not (a xor b);
    layer2_outputs(821) <= not a;
    layer2_outputs(822) <= a or b;
    layer2_outputs(823) <= not b or a;
    layer2_outputs(824) <= not a or b;
    layer2_outputs(825) <= '0';
    layer2_outputs(826) <= not b or a;
    layer2_outputs(827) <= a;
    layer2_outputs(828) <= b;
    layer2_outputs(829) <= a and not b;
    layer2_outputs(830) <= b and not a;
    layer2_outputs(831) <= not b;
    layer2_outputs(832) <= not (a or b);
    layer2_outputs(833) <= '0';
    layer2_outputs(834) <= a;
    layer2_outputs(835) <= b;
    layer2_outputs(836) <= not a;
    layer2_outputs(837) <= not b or a;
    layer2_outputs(838) <= not (a or b);
    layer2_outputs(839) <= not (a or b);
    layer2_outputs(840) <= not a or b;
    layer2_outputs(841) <= not (a and b);
    layer2_outputs(842) <= b;
    layer2_outputs(843) <= b and not a;
    layer2_outputs(844) <= not (a or b);
    layer2_outputs(845) <= a and not b;
    layer2_outputs(846) <= a or b;
    layer2_outputs(847) <= b;
    layer2_outputs(848) <= not a or b;
    layer2_outputs(849) <= a and not b;
    layer2_outputs(850) <= b and not a;
    layer2_outputs(851) <= a and not b;
    layer2_outputs(852) <= not b or a;
    layer2_outputs(853) <= a;
    layer2_outputs(854) <= not b or a;
    layer2_outputs(855) <= b and not a;
    layer2_outputs(856) <= not (a or b);
    layer2_outputs(857) <= a and b;
    layer2_outputs(858) <= a and b;
    layer2_outputs(859) <= not (a and b);
    layer2_outputs(860) <= b;
    layer2_outputs(861) <= a and b;
    layer2_outputs(862) <= not (a xor b);
    layer2_outputs(863) <= b;
    layer2_outputs(864) <= b and not a;
    layer2_outputs(865) <= b;
    layer2_outputs(866) <= not (a or b);
    layer2_outputs(867) <= b and not a;
    layer2_outputs(868) <= a xor b;
    layer2_outputs(869) <= not a;
    layer2_outputs(870) <= b and not a;
    layer2_outputs(871) <= b;
    layer2_outputs(872) <= not a;
    layer2_outputs(873) <= b;
    layer2_outputs(874) <= a or b;
    layer2_outputs(875) <= a and not b;
    layer2_outputs(876) <= not a or b;
    layer2_outputs(877) <= b;
    layer2_outputs(878) <= not a;
    layer2_outputs(879) <= b and not a;
    layer2_outputs(880) <= a xor b;
    layer2_outputs(881) <= a or b;
    layer2_outputs(882) <= a;
    layer2_outputs(883) <= a or b;
    layer2_outputs(884) <= a xor b;
    layer2_outputs(885) <= a and b;
    layer2_outputs(886) <= '0';
    layer2_outputs(887) <= b and not a;
    layer2_outputs(888) <= a;
    layer2_outputs(889) <= not b;
    layer2_outputs(890) <= a;
    layer2_outputs(891) <= b;
    layer2_outputs(892) <= a;
    layer2_outputs(893) <= not b or a;
    layer2_outputs(894) <= b;
    layer2_outputs(895) <= b;
    layer2_outputs(896) <= b and not a;
    layer2_outputs(897) <= not b or a;
    layer2_outputs(898) <= not (a or b);
    layer2_outputs(899) <= not (a and b);
    layer2_outputs(900) <= a or b;
    layer2_outputs(901) <= b;
    layer2_outputs(902) <= not (a or b);
    layer2_outputs(903) <= not a;
    layer2_outputs(904) <= a or b;
    layer2_outputs(905) <= not b;
    layer2_outputs(906) <= not a;
    layer2_outputs(907) <= b;
    layer2_outputs(908) <= not b;
    layer2_outputs(909) <= b;
    layer2_outputs(910) <= not a;
    layer2_outputs(911) <= not b or a;
    layer2_outputs(912) <= not a;
    layer2_outputs(913) <= a and not b;
    layer2_outputs(914) <= '1';
    layer2_outputs(915) <= not b;
    layer2_outputs(916) <= a and b;
    layer2_outputs(917) <= b;
    layer2_outputs(918) <= not (a and b);
    layer2_outputs(919) <= not a;
    layer2_outputs(920) <= a and not b;
    layer2_outputs(921) <= b;
    layer2_outputs(922) <= not b;
    layer2_outputs(923) <= not (a and b);
    layer2_outputs(924) <= not a or b;
    layer2_outputs(925) <= a and b;
    layer2_outputs(926) <= b and not a;
    layer2_outputs(927) <= '0';
    layer2_outputs(928) <= not a or b;
    layer2_outputs(929) <= b;
    layer2_outputs(930) <= a;
    layer2_outputs(931) <= not a;
    layer2_outputs(932) <= b;
    layer2_outputs(933) <= not a;
    layer2_outputs(934) <= a;
    layer2_outputs(935) <= b;
    layer2_outputs(936) <= not (a and b);
    layer2_outputs(937) <= not b;
    layer2_outputs(938) <= b;
    layer2_outputs(939) <= not (a or b);
    layer2_outputs(940) <= not b or a;
    layer2_outputs(941) <= not (a or b);
    layer2_outputs(942) <= not a or b;
    layer2_outputs(943) <= a and b;
    layer2_outputs(944) <= not a;
    layer2_outputs(945) <= not (a or b);
    layer2_outputs(946) <= not a;
    layer2_outputs(947) <= a or b;
    layer2_outputs(948) <= a;
    layer2_outputs(949) <= a xor b;
    layer2_outputs(950) <= a or b;
    layer2_outputs(951) <= b and not a;
    layer2_outputs(952) <= not a;
    layer2_outputs(953) <= not a;
    layer2_outputs(954) <= a or b;
    layer2_outputs(955) <= b;
    layer2_outputs(956) <= not a;
    layer2_outputs(957) <= not a or b;
    layer2_outputs(958) <= not b;
    layer2_outputs(959) <= not (a or b);
    layer2_outputs(960) <= a and not b;
    layer2_outputs(961) <= b and not a;
    layer2_outputs(962) <= not a;
    layer2_outputs(963) <= a;
    layer2_outputs(964) <= a xor b;
    layer2_outputs(965) <= a;
    layer2_outputs(966) <= a or b;
    layer2_outputs(967) <= not a;
    layer2_outputs(968) <= a xor b;
    layer2_outputs(969) <= a;
    layer2_outputs(970) <= a;
    layer2_outputs(971) <= a and b;
    layer2_outputs(972) <= a and not b;
    layer2_outputs(973) <= a and not b;
    layer2_outputs(974) <= a;
    layer2_outputs(975) <= not (a or b);
    layer2_outputs(976) <= a;
    layer2_outputs(977) <= b and not a;
    layer2_outputs(978) <= b;
    layer2_outputs(979) <= a;
    layer2_outputs(980) <= not b;
    layer2_outputs(981) <= not a or b;
    layer2_outputs(982) <= a or b;
    layer2_outputs(983) <= not (a and b);
    layer2_outputs(984) <= not b;
    layer2_outputs(985) <= b and not a;
    layer2_outputs(986) <= not b;
    layer2_outputs(987) <= a;
    layer2_outputs(988) <= a xor b;
    layer2_outputs(989) <= a;
    layer2_outputs(990) <= a and not b;
    layer2_outputs(991) <= a xor b;
    layer2_outputs(992) <= b and not a;
    layer2_outputs(993) <= not b;
    layer2_outputs(994) <= not b;
    layer2_outputs(995) <= a;
    layer2_outputs(996) <= a and b;
    layer2_outputs(997) <= a;
    layer2_outputs(998) <= '0';
    layer2_outputs(999) <= a;
    layer2_outputs(1000) <= not (a or b);
    layer2_outputs(1001) <= a or b;
    layer2_outputs(1002) <= a and b;
    layer2_outputs(1003) <= b;
    layer2_outputs(1004) <= a or b;
    layer2_outputs(1005) <= a and b;
    layer2_outputs(1006) <= a or b;
    layer2_outputs(1007) <= not (a or b);
    layer2_outputs(1008) <= a;
    layer2_outputs(1009) <= a or b;
    layer2_outputs(1010) <= not a or b;
    layer2_outputs(1011) <= '1';
    layer2_outputs(1012) <= a or b;
    layer2_outputs(1013) <= a or b;
    layer2_outputs(1014) <= b;
    layer2_outputs(1015) <= not a;
    layer2_outputs(1016) <= not a or b;
    layer2_outputs(1017) <= b;
    layer2_outputs(1018) <= a;
    layer2_outputs(1019) <= a or b;
    layer2_outputs(1020) <= a;
    layer2_outputs(1021) <= '1';
    layer2_outputs(1022) <= not b or a;
    layer2_outputs(1023) <= a xor b;
    layer2_outputs(1024) <= not b;
    layer2_outputs(1025) <= a or b;
    layer2_outputs(1026) <= not a or b;
    layer2_outputs(1027) <= a and b;
    layer2_outputs(1028) <= not (a or b);
    layer2_outputs(1029) <= not b;
    layer2_outputs(1030) <= not a;
    layer2_outputs(1031) <= not (a and b);
    layer2_outputs(1032) <= not a;
    layer2_outputs(1033) <= not (a or b);
    layer2_outputs(1034) <= not (a and b);
    layer2_outputs(1035) <= a and b;
    layer2_outputs(1036) <= not (a or b);
    layer2_outputs(1037) <= not (a or b);
    layer2_outputs(1038) <= '1';
    layer2_outputs(1039) <= a and b;
    layer2_outputs(1040) <= a;
    layer2_outputs(1041) <= '1';
    layer2_outputs(1042) <= a or b;
    layer2_outputs(1043) <= not (a or b);
    layer2_outputs(1044) <= not b;
    layer2_outputs(1045) <= not b;
    layer2_outputs(1046) <= b;
    layer2_outputs(1047) <= '1';
    layer2_outputs(1048) <= not b or a;
    layer2_outputs(1049) <= a and not b;
    layer2_outputs(1050) <= not a;
    layer2_outputs(1051) <= '0';
    layer2_outputs(1052) <= b;
    layer2_outputs(1053) <= not (a or b);
    layer2_outputs(1054) <= a or b;
    layer2_outputs(1055) <= a;
    layer2_outputs(1056) <= b and not a;
    layer2_outputs(1057) <= not (a and b);
    layer2_outputs(1058) <= '0';
    layer2_outputs(1059) <= not (a xor b);
    layer2_outputs(1060) <= a xor b;
    layer2_outputs(1061) <= b;
    layer2_outputs(1062) <= '1';
    layer2_outputs(1063) <= a and not b;
    layer2_outputs(1064) <= b and not a;
    layer2_outputs(1065) <= b;
    layer2_outputs(1066) <= not a;
    layer2_outputs(1067) <= not a or b;
    layer2_outputs(1068) <= not a;
    layer2_outputs(1069) <= a;
    layer2_outputs(1070) <= b and not a;
    layer2_outputs(1071) <= not b;
    layer2_outputs(1072) <= a;
    layer2_outputs(1073) <= a;
    layer2_outputs(1074) <= not a;
    layer2_outputs(1075) <= not a or b;
    layer2_outputs(1076) <= not a;
    layer2_outputs(1077) <= not b or a;
    layer2_outputs(1078) <= b and not a;
    layer2_outputs(1079) <= not b;
    layer2_outputs(1080) <= '0';
    layer2_outputs(1081) <= a and not b;
    layer2_outputs(1082) <= not a;
    layer2_outputs(1083) <= not a;
    layer2_outputs(1084) <= not a or b;
    layer2_outputs(1085) <= not (a or b);
    layer2_outputs(1086) <= a or b;
    layer2_outputs(1087) <= a and b;
    layer2_outputs(1088) <= a and b;
    layer2_outputs(1089) <= b;
    layer2_outputs(1090) <= not a;
    layer2_outputs(1091) <= not b or a;
    layer2_outputs(1092) <= not a;
    layer2_outputs(1093) <= not a;
    layer2_outputs(1094) <= not a;
    layer2_outputs(1095) <= b;
    layer2_outputs(1096) <= b;
    layer2_outputs(1097) <= b;
    layer2_outputs(1098) <= a or b;
    layer2_outputs(1099) <= not b or a;
    layer2_outputs(1100) <= not (a or b);
    layer2_outputs(1101) <= not a;
    layer2_outputs(1102) <= not a or b;
    layer2_outputs(1103) <= not b or a;
    layer2_outputs(1104) <= not a;
    layer2_outputs(1105) <= b and not a;
    layer2_outputs(1106) <= b and not a;
    layer2_outputs(1107) <= not (a and b);
    layer2_outputs(1108) <= not b or a;
    layer2_outputs(1109) <= a;
    layer2_outputs(1110) <= not a or b;
    layer2_outputs(1111) <= not (a and b);
    layer2_outputs(1112) <= not b;
    layer2_outputs(1113) <= not (a and b);
    layer2_outputs(1114) <= not a;
    layer2_outputs(1115) <= b;
    layer2_outputs(1116) <= a and b;
    layer2_outputs(1117) <= b and not a;
    layer2_outputs(1118) <= not a or b;
    layer2_outputs(1119) <= a and not b;
    layer2_outputs(1120) <= not (a xor b);
    layer2_outputs(1121) <= not b;
    layer2_outputs(1122) <= b and not a;
    layer2_outputs(1123) <= a or b;
    layer2_outputs(1124) <= a;
    layer2_outputs(1125) <= b;
    layer2_outputs(1126) <= a and b;
    layer2_outputs(1127) <= a;
    layer2_outputs(1128) <= a and not b;
    layer2_outputs(1129) <= not a;
    layer2_outputs(1130) <= not b or a;
    layer2_outputs(1131) <= a and not b;
    layer2_outputs(1132) <= b;
    layer2_outputs(1133) <= not b;
    layer2_outputs(1134) <= a;
    layer2_outputs(1135) <= not b;
    layer2_outputs(1136) <= not b;
    layer2_outputs(1137) <= not (a and b);
    layer2_outputs(1138) <= not a;
    layer2_outputs(1139) <= b and not a;
    layer2_outputs(1140) <= a and not b;
    layer2_outputs(1141) <= not (a xor b);
    layer2_outputs(1142) <= not a;
    layer2_outputs(1143) <= not (a and b);
    layer2_outputs(1144) <= a and b;
    layer2_outputs(1145) <= '1';
    layer2_outputs(1146) <= a xor b;
    layer2_outputs(1147) <= b and not a;
    layer2_outputs(1148) <= b and not a;
    layer2_outputs(1149) <= not (a or b);
    layer2_outputs(1150) <= not b or a;
    layer2_outputs(1151) <= a;
    layer2_outputs(1152) <= a or b;
    layer2_outputs(1153) <= '0';
    layer2_outputs(1154) <= not (a and b);
    layer2_outputs(1155) <= a;
    layer2_outputs(1156) <= '0';
    layer2_outputs(1157) <= a;
    layer2_outputs(1158) <= b;
    layer2_outputs(1159) <= not b;
    layer2_outputs(1160) <= not b;
    layer2_outputs(1161) <= b and not a;
    layer2_outputs(1162) <= b and not a;
    layer2_outputs(1163) <= a or b;
    layer2_outputs(1164) <= not a;
    layer2_outputs(1165) <= a;
    layer2_outputs(1166) <= b and not a;
    layer2_outputs(1167) <= not a;
    layer2_outputs(1168) <= not a;
    layer2_outputs(1169) <= a and not b;
    layer2_outputs(1170) <= a or b;
    layer2_outputs(1171) <= not (a or b);
    layer2_outputs(1172) <= not (a or b);
    layer2_outputs(1173) <= b;
    layer2_outputs(1174) <= a;
    layer2_outputs(1175) <= a;
    layer2_outputs(1176) <= a or b;
    layer2_outputs(1177) <= not (a or b);
    layer2_outputs(1178) <= not b or a;
    layer2_outputs(1179) <= a and b;
    layer2_outputs(1180) <= b and not a;
    layer2_outputs(1181) <= not (a or b);
    layer2_outputs(1182) <= not b;
    layer2_outputs(1183) <= not b or a;
    layer2_outputs(1184) <= b;
    layer2_outputs(1185) <= a xor b;
    layer2_outputs(1186) <= not b;
    layer2_outputs(1187) <= not b;
    layer2_outputs(1188) <= b;
    layer2_outputs(1189) <= not (a and b);
    layer2_outputs(1190) <= b;
    layer2_outputs(1191) <= b and not a;
    layer2_outputs(1192) <= a and b;
    layer2_outputs(1193) <= a or b;
    layer2_outputs(1194) <= not (a or b);
    layer2_outputs(1195) <= a and b;
    layer2_outputs(1196) <= not a or b;
    layer2_outputs(1197) <= not b;
    layer2_outputs(1198) <= not (a xor b);
    layer2_outputs(1199) <= b;
    layer2_outputs(1200) <= a;
    layer2_outputs(1201) <= not (a or b);
    layer2_outputs(1202) <= not b;
    layer2_outputs(1203) <= not a or b;
    layer2_outputs(1204) <= a and b;
    layer2_outputs(1205) <= a;
    layer2_outputs(1206) <= a and b;
    layer2_outputs(1207) <= not a or b;
    layer2_outputs(1208) <= a or b;
    layer2_outputs(1209) <= a or b;
    layer2_outputs(1210) <= b;
    layer2_outputs(1211) <= not a;
    layer2_outputs(1212) <= '0';
    layer2_outputs(1213) <= a or b;
    layer2_outputs(1214) <= not (a and b);
    layer2_outputs(1215) <= not b or a;
    layer2_outputs(1216) <= a;
    layer2_outputs(1217) <= a and not b;
    layer2_outputs(1218) <= a;
    layer2_outputs(1219) <= not b;
    layer2_outputs(1220) <= not b;
    layer2_outputs(1221) <= not a;
    layer2_outputs(1222) <= '0';
    layer2_outputs(1223) <= not a;
    layer2_outputs(1224) <= not b;
    layer2_outputs(1225) <= not (a and b);
    layer2_outputs(1226) <= not (a and b);
    layer2_outputs(1227) <= b and not a;
    layer2_outputs(1228) <= a;
    layer2_outputs(1229) <= b and not a;
    layer2_outputs(1230) <= b;
    layer2_outputs(1231) <= a;
    layer2_outputs(1232) <= a and b;
    layer2_outputs(1233) <= not (a or b);
    layer2_outputs(1234) <= a;
    layer2_outputs(1235) <= not b or a;
    layer2_outputs(1236) <= not b;
    layer2_outputs(1237) <= not b or a;
    layer2_outputs(1238) <= a and not b;
    layer2_outputs(1239) <= not b;
    layer2_outputs(1240) <= a or b;
    layer2_outputs(1241) <= not b or a;
    layer2_outputs(1242) <= not b;
    layer2_outputs(1243) <= not b or a;
    layer2_outputs(1244) <= b;
    layer2_outputs(1245) <= b;
    layer2_outputs(1246) <= a;
    layer2_outputs(1247) <= a xor b;
    layer2_outputs(1248) <= b and not a;
    layer2_outputs(1249) <= a or b;
    layer2_outputs(1250) <= b;
    layer2_outputs(1251) <= a and b;
    layer2_outputs(1252) <= a xor b;
    layer2_outputs(1253) <= not a or b;
    layer2_outputs(1254) <= not b;
    layer2_outputs(1255) <= b;
    layer2_outputs(1256) <= b;
    layer2_outputs(1257) <= '1';
    layer2_outputs(1258) <= not a;
    layer2_outputs(1259) <= b;
    layer2_outputs(1260) <= a and b;
    layer2_outputs(1261) <= not (a or b);
    layer2_outputs(1262) <= a and b;
    layer2_outputs(1263) <= not b or a;
    layer2_outputs(1264) <= not b;
    layer2_outputs(1265) <= b and not a;
    layer2_outputs(1266) <= '0';
    layer2_outputs(1267) <= not a;
    layer2_outputs(1268) <= b;
    layer2_outputs(1269) <= not (a xor b);
    layer2_outputs(1270) <= not (a or b);
    layer2_outputs(1271) <= not (a and b);
    layer2_outputs(1272) <= a;
    layer2_outputs(1273) <= a xor b;
    layer2_outputs(1274) <= b;
    layer2_outputs(1275) <= a and not b;
    layer2_outputs(1276) <= not a;
    layer2_outputs(1277) <= not (a and b);
    layer2_outputs(1278) <= b and not a;
    layer2_outputs(1279) <= a and b;
    layer2_outputs(1280) <= not (a and b);
    layer2_outputs(1281) <= not b;
    layer2_outputs(1282) <= not a or b;
    layer2_outputs(1283) <= a and b;
    layer2_outputs(1284) <= a;
    layer2_outputs(1285) <= not (a xor b);
    layer2_outputs(1286) <= a;
    layer2_outputs(1287) <= a and not b;
    layer2_outputs(1288) <= not a or b;
    layer2_outputs(1289) <= a;
    layer2_outputs(1290) <= a or b;
    layer2_outputs(1291) <= not b;
    layer2_outputs(1292) <= '1';
    layer2_outputs(1293) <= a and b;
    layer2_outputs(1294) <= '0';
    layer2_outputs(1295) <= not b;
    layer2_outputs(1296) <= not a or b;
    layer2_outputs(1297) <= not a or b;
    layer2_outputs(1298) <= not b or a;
    layer2_outputs(1299) <= not a or b;
    layer2_outputs(1300) <= not b;
    layer2_outputs(1301) <= a and b;
    layer2_outputs(1302) <= not a;
    layer2_outputs(1303) <= not (a and b);
    layer2_outputs(1304) <= b;
    layer2_outputs(1305) <= b;
    layer2_outputs(1306) <= a xor b;
    layer2_outputs(1307) <= not b;
    layer2_outputs(1308) <= not (a and b);
    layer2_outputs(1309) <= a;
    layer2_outputs(1310) <= '1';
    layer2_outputs(1311) <= b;
    layer2_outputs(1312) <= b and not a;
    layer2_outputs(1313) <= b;
    layer2_outputs(1314) <= not (a and b);
    layer2_outputs(1315) <= a or b;
    layer2_outputs(1316) <= b;
    layer2_outputs(1317) <= not b;
    layer2_outputs(1318) <= a;
    layer2_outputs(1319) <= not (a xor b);
    layer2_outputs(1320) <= a and not b;
    layer2_outputs(1321) <= not b;
    layer2_outputs(1322) <= a;
    layer2_outputs(1323) <= not (a and b);
    layer2_outputs(1324) <= not b;
    layer2_outputs(1325) <= not a or b;
    layer2_outputs(1326) <= '1';
    layer2_outputs(1327) <= a or b;
    layer2_outputs(1328) <= not (a and b);
    layer2_outputs(1329) <= '1';
    layer2_outputs(1330) <= not b or a;
    layer2_outputs(1331) <= a and b;
    layer2_outputs(1332) <= not a;
    layer2_outputs(1333) <= not a or b;
    layer2_outputs(1334) <= b and not a;
    layer2_outputs(1335) <= a and not b;
    layer2_outputs(1336) <= not (a and b);
    layer2_outputs(1337) <= '1';
    layer2_outputs(1338) <= a and not b;
    layer2_outputs(1339) <= b;
    layer2_outputs(1340) <= '1';
    layer2_outputs(1341) <= '0';
    layer2_outputs(1342) <= not a;
    layer2_outputs(1343) <= a or b;
    layer2_outputs(1344) <= b;
    layer2_outputs(1345) <= not (a or b);
    layer2_outputs(1346) <= not b;
    layer2_outputs(1347) <= not b or a;
    layer2_outputs(1348) <= b;
    layer2_outputs(1349) <= b;
    layer2_outputs(1350) <= not b;
    layer2_outputs(1351) <= a and not b;
    layer2_outputs(1352) <= a;
    layer2_outputs(1353) <= not a;
    layer2_outputs(1354) <= not a;
    layer2_outputs(1355) <= not a;
    layer2_outputs(1356) <= a and not b;
    layer2_outputs(1357) <= not a;
    layer2_outputs(1358) <= not b or a;
    layer2_outputs(1359) <= a and b;
    layer2_outputs(1360) <= not a;
    layer2_outputs(1361) <= a;
    layer2_outputs(1362) <= b;
    layer2_outputs(1363) <= not b;
    layer2_outputs(1364) <= not a;
    layer2_outputs(1365) <= not a;
    layer2_outputs(1366) <= not a or b;
    layer2_outputs(1367) <= not b;
    layer2_outputs(1368) <= not b or a;
    layer2_outputs(1369) <= '0';
    layer2_outputs(1370) <= a or b;
    layer2_outputs(1371) <= b;
    layer2_outputs(1372) <= a and b;
    layer2_outputs(1373) <= a;
    layer2_outputs(1374) <= a or b;
    layer2_outputs(1375) <= a and b;
    layer2_outputs(1376) <= not (a or b);
    layer2_outputs(1377) <= a xor b;
    layer2_outputs(1378) <= a and b;
    layer2_outputs(1379) <= '1';
    layer2_outputs(1380) <= a and not b;
    layer2_outputs(1381) <= b and not a;
    layer2_outputs(1382) <= not a or b;
    layer2_outputs(1383) <= not a;
    layer2_outputs(1384) <= not (a and b);
    layer2_outputs(1385) <= a;
    layer2_outputs(1386) <= not (a and b);
    layer2_outputs(1387) <= b and not a;
    layer2_outputs(1388) <= a;
    layer2_outputs(1389) <= b;
    layer2_outputs(1390) <= a xor b;
    layer2_outputs(1391) <= b;
    layer2_outputs(1392) <= not a;
    layer2_outputs(1393) <= a or b;
    layer2_outputs(1394) <= a xor b;
    layer2_outputs(1395) <= a and b;
    layer2_outputs(1396) <= not a;
    layer2_outputs(1397) <= a and b;
    layer2_outputs(1398) <= not (a and b);
    layer2_outputs(1399) <= a and b;
    layer2_outputs(1400) <= not a;
    layer2_outputs(1401) <= not b or a;
    layer2_outputs(1402) <= a;
    layer2_outputs(1403) <= '1';
    layer2_outputs(1404) <= a or b;
    layer2_outputs(1405) <= not a or b;
    layer2_outputs(1406) <= not (a and b);
    layer2_outputs(1407) <= a or b;
    layer2_outputs(1408) <= not (a or b);
    layer2_outputs(1409) <= a;
    layer2_outputs(1410) <= a and not b;
    layer2_outputs(1411) <= not (a and b);
    layer2_outputs(1412) <= a and not b;
    layer2_outputs(1413) <= not b;
    layer2_outputs(1414) <= not (a and b);
    layer2_outputs(1415) <= not b;
    layer2_outputs(1416) <= '1';
    layer2_outputs(1417) <= b;
    layer2_outputs(1418) <= b;
    layer2_outputs(1419) <= b;
    layer2_outputs(1420) <= a;
    layer2_outputs(1421) <= b;
    layer2_outputs(1422) <= b and not a;
    layer2_outputs(1423) <= not a;
    layer2_outputs(1424) <= '1';
    layer2_outputs(1425) <= a and b;
    layer2_outputs(1426) <= a xor b;
    layer2_outputs(1427) <= not a;
    layer2_outputs(1428) <= not (a or b);
    layer2_outputs(1429) <= not a;
    layer2_outputs(1430) <= a xor b;
    layer2_outputs(1431) <= not b or a;
    layer2_outputs(1432) <= a and not b;
    layer2_outputs(1433) <= not (a or b);
    layer2_outputs(1434) <= not b;
    layer2_outputs(1435) <= a and b;
    layer2_outputs(1436) <= not a;
    layer2_outputs(1437) <= not a;
    layer2_outputs(1438) <= b and not a;
    layer2_outputs(1439) <= not a or b;
    layer2_outputs(1440) <= a and not b;
    layer2_outputs(1441) <= a or b;
    layer2_outputs(1442) <= not a or b;
    layer2_outputs(1443) <= a;
    layer2_outputs(1444) <= a;
    layer2_outputs(1445) <= a and not b;
    layer2_outputs(1446) <= not (a xor b);
    layer2_outputs(1447) <= not b or a;
    layer2_outputs(1448) <= not a;
    layer2_outputs(1449) <= a and not b;
    layer2_outputs(1450) <= a;
    layer2_outputs(1451) <= a;
    layer2_outputs(1452) <= not (a xor b);
    layer2_outputs(1453) <= '0';
    layer2_outputs(1454) <= a and b;
    layer2_outputs(1455) <= not b or a;
    layer2_outputs(1456) <= b;
    layer2_outputs(1457) <= not b or a;
    layer2_outputs(1458) <= a;
    layer2_outputs(1459) <= a;
    layer2_outputs(1460) <= not a or b;
    layer2_outputs(1461) <= not b;
    layer2_outputs(1462) <= b;
    layer2_outputs(1463) <= not (a and b);
    layer2_outputs(1464) <= not a or b;
    layer2_outputs(1465) <= not a;
    layer2_outputs(1466) <= not a or b;
    layer2_outputs(1467) <= not b;
    layer2_outputs(1468) <= a and not b;
    layer2_outputs(1469) <= a and not b;
    layer2_outputs(1470) <= a and b;
    layer2_outputs(1471) <= b;
    layer2_outputs(1472) <= a and b;
    layer2_outputs(1473) <= not a or b;
    layer2_outputs(1474) <= not a;
    layer2_outputs(1475) <= b and not a;
    layer2_outputs(1476) <= a and not b;
    layer2_outputs(1477) <= not a;
    layer2_outputs(1478) <= a xor b;
    layer2_outputs(1479) <= not a or b;
    layer2_outputs(1480) <= b;
    layer2_outputs(1481) <= a xor b;
    layer2_outputs(1482) <= a;
    layer2_outputs(1483) <= not b;
    layer2_outputs(1484) <= not b;
    layer2_outputs(1485) <= a or b;
    layer2_outputs(1486) <= not b;
    layer2_outputs(1487) <= not b;
    layer2_outputs(1488) <= b;
    layer2_outputs(1489) <= not a;
    layer2_outputs(1490) <= not b;
    layer2_outputs(1491) <= b;
    layer2_outputs(1492) <= not a;
    layer2_outputs(1493) <= not b;
    layer2_outputs(1494) <= b and not a;
    layer2_outputs(1495) <= not a;
    layer2_outputs(1496) <= not (a and b);
    layer2_outputs(1497) <= a;
    layer2_outputs(1498) <= not a;
    layer2_outputs(1499) <= not (a xor b);
    layer2_outputs(1500) <= a and not b;
    layer2_outputs(1501) <= b and not a;
    layer2_outputs(1502) <= not (a xor b);
    layer2_outputs(1503) <= not a;
    layer2_outputs(1504) <= a and b;
    layer2_outputs(1505) <= not b or a;
    layer2_outputs(1506) <= a or b;
    layer2_outputs(1507) <= b;
    layer2_outputs(1508) <= b and not a;
    layer2_outputs(1509) <= a xor b;
    layer2_outputs(1510) <= not (a or b);
    layer2_outputs(1511) <= not (a or b);
    layer2_outputs(1512) <= b and not a;
    layer2_outputs(1513) <= a and b;
    layer2_outputs(1514) <= not a or b;
    layer2_outputs(1515) <= not (a and b);
    layer2_outputs(1516) <= b and not a;
    layer2_outputs(1517) <= not (a xor b);
    layer2_outputs(1518) <= not a;
    layer2_outputs(1519) <= not (a or b);
    layer2_outputs(1520) <= not a or b;
    layer2_outputs(1521) <= a and b;
    layer2_outputs(1522) <= a;
    layer2_outputs(1523) <= b;
    layer2_outputs(1524) <= not b or a;
    layer2_outputs(1525) <= not (a and b);
    layer2_outputs(1526) <= a;
    layer2_outputs(1527) <= not b;
    layer2_outputs(1528) <= not a or b;
    layer2_outputs(1529) <= not a or b;
    layer2_outputs(1530) <= a or b;
    layer2_outputs(1531) <= b and not a;
    layer2_outputs(1532) <= not (a or b);
    layer2_outputs(1533) <= not a or b;
    layer2_outputs(1534) <= '0';
    layer2_outputs(1535) <= a and not b;
    layer2_outputs(1536) <= '1';
    layer2_outputs(1537) <= b and not a;
    layer2_outputs(1538) <= '0';
    layer2_outputs(1539) <= a;
    layer2_outputs(1540) <= not (a or b);
    layer2_outputs(1541) <= a;
    layer2_outputs(1542) <= b;
    layer2_outputs(1543) <= b;
    layer2_outputs(1544) <= '0';
    layer2_outputs(1545) <= not b or a;
    layer2_outputs(1546) <= '1';
    layer2_outputs(1547) <= a and b;
    layer2_outputs(1548) <= b;
    layer2_outputs(1549) <= not (a xor b);
    layer2_outputs(1550) <= a or b;
    layer2_outputs(1551) <= not a;
    layer2_outputs(1552) <= b;
    layer2_outputs(1553) <= b and not a;
    layer2_outputs(1554) <= not b or a;
    layer2_outputs(1555) <= not b or a;
    layer2_outputs(1556) <= not b or a;
    layer2_outputs(1557) <= not b;
    layer2_outputs(1558) <= not (a and b);
    layer2_outputs(1559) <= not (a and b);
    layer2_outputs(1560) <= a;
    layer2_outputs(1561) <= a or b;
    layer2_outputs(1562) <= a or b;
    layer2_outputs(1563) <= not b;
    layer2_outputs(1564) <= a and not b;
    layer2_outputs(1565) <= a and b;
    layer2_outputs(1566) <= a and not b;
    layer2_outputs(1567) <= not b;
    layer2_outputs(1568) <= a;
    layer2_outputs(1569) <= b and not a;
    layer2_outputs(1570) <= not (a or b);
    layer2_outputs(1571) <= '1';
    layer2_outputs(1572) <= not (a and b);
    layer2_outputs(1573) <= b;
    layer2_outputs(1574) <= a and not b;
    layer2_outputs(1575) <= a and not b;
    layer2_outputs(1576) <= b and not a;
    layer2_outputs(1577) <= not (a and b);
    layer2_outputs(1578) <= not a;
    layer2_outputs(1579) <= not a;
    layer2_outputs(1580) <= a;
    layer2_outputs(1581) <= not (a or b);
    layer2_outputs(1582) <= not b;
    layer2_outputs(1583) <= not b or a;
    layer2_outputs(1584) <= not b or a;
    layer2_outputs(1585) <= not a;
    layer2_outputs(1586) <= '0';
    layer2_outputs(1587) <= not (a xor b);
    layer2_outputs(1588) <= a and not b;
    layer2_outputs(1589) <= not a;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= a xor b;
    layer2_outputs(1592) <= b and not a;
    layer2_outputs(1593) <= not (a xor b);
    layer2_outputs(1594) <= not b;
    layer2_outputs(1595) <= not a;
    layer2_outputs(1596) <= not a;
    layer2_outputs(1597) <= b;
    layer2_outputs(1598) <= not (a or b);
    layer2_outputs(1599) <= not (a and b);
    layer2_outputs(1600) <= not b;
    layer2_outputs(1601) <= not a;
    layer2_outputs(1602) <= a xor b;
    layer2_outputs(1603) <= not b;
    layer2_outputs(1604) <= b;
    layer2_outputs(1605) <= not (a and b);
    layer2_outputs(1606) <= b;
    layer2_outputs(1607) <= not (a xor b);
    layer2_outputs(1608) <= a xor b;
    layer2_outputs(1609) <= not a;
    layer2_outputs(1610) <= a;
    layer2_outputs(1611) <= not b or a;
    layer2_outputs(1612) <= a and not b;
    layer2_outputs(1613) <= b;
    layer2_outputs(1614) <= not b or a;
    layer2_outputs(1615) <= not a or b;
    layer2_outputs(1616) <= a or b;
    layer2_outputs(1617) <= '1';
    layer2_outputs(1618) <= a and not b;
    layer2_outputs(1619) <= not a or b;
    layer2_outputs(1620) <= not (a and b);
    layer2_outputs(1621) <= not a;
    layer2_outputs(1622) <= not (a and b);
    layer2_outputs(1623) <= not b or a;
    layer2_outputs(1624) <= a xor b;
    layer2_outputs(1625) <= not b or a;
    layer2_outputs(1626) <= not (a and b);
    layer2_outputs(1627) <= a and b;
    layer2_outputs(1628) <= not a or b;
    layer2_outputs(1629) <= not (a or b);
    layer2_outputs(1630) <= a xor b;
    layer2_outputs(1631) <= not b;
    layer2_outputs(1632) <= b;
    layer2_outputs(1633) <= a or b;
    layer2_outputs(1634) <= a and not b;
    layer2_outputs(1635) <= b and not a;
    layer2_outputs(1636) <= not a or b;
    layer2_outputs(1637) <= a xor b;
    layer2_outputs(1638) <= a and b;
    layer2_outputs(1639) <= b and not a;
    layer2_outputs(1640) <= not (a and b);
    layer2_outputs(1641) <= not b or a;
    layer2_outputs(1642) <= a;
    layer2_outputs(1643) <= not (a and b);
    layer2_outputs(1644) <= not a;
    layer2_outputs(1645) <= not b;
    layer2_outputs(1646) <= not b or a;
    layer2_outputs(1647) <= b;
    layer2_outputs(1648) <= a;
    layer2_outputs(1649) <= not (a or b);
    layer2_outputs(1650) <= a and not b;
    layer2_outputs(1651) <= not (a or b);
    layer2_outputs(1652) <= not a;
    layer2_outputs(1653) <= not b;
    layer2_outputs(1654) <= '1';
    layer2_outputs(1655) <= not a or b;
    layer2_outputs(1656) <= not b;
    layer2_outputs(1657) <= not b or a;
    layer2_outputs(1658) <= b;
    layer2_outputs(1659) <= not b;
    layer2_outputs(1660) <= a and b;
    layer2_outputs(1661) <= not a;
    layer2_outputs(1662) <= a;
    layer2_outputs(1663) <= b and not a;
    layer2_outputs(1664) <= a and b;
    layer2_outputs(1665) <= not b;
    layer2_outputs(1666) <= not b;
    layer2_outputs(1667) <= b;
    layer2_outputs(1668) <= a or b;
    layer2_outputs(1669) <= not b or a;
    layer2_outputs(1670) <= not b;
    layer2_outputs(1671) <= not a;
    layer2_outputs(1672) <= a and not b;
    layer2_outputs(1673) <= a;
    layer2_outputs(1674) <= '1';
    layer2_outputs(1675) <= not b;
    layer2_outputs(1676) <= not (a and b);
    layer2_outputs(1677) <= not b;
    layer2_outputs(1678) <= b;
    layer2_outputs(1679) <= not a;
    layer2_outputs(1680) <= a or b;
    layer2_outputs(1681) <= b;
    layer2_outputs(1682) <= not (a and b);
    layer2_outputs(1683) <= not a or b;
    layer2_outputs(1684) <= not b or a;
    layer2_outputs(1685) <= b and not a;
    layer2_outputs(1686) <= '1';
    layer2_outputs(1687) <= a or b;
    layer2_outputs(1688) <= b and not a;
    layer2_outputs(1689) <= not a;
    layer2_outputs(1690) <= not a or b;
    layer2_outputs(1691) <= not b or a;
    layer2_outputs(1692) <= b;
    layer2_outputs(1693) <= a;
    layer2_outputs(1694) <= not b;
    layer2_outputs(1695) <= not b or a;
    layer2_outputs(1696) <= b;
    layer2_outputs(1697) <= not b or a;
    layer2_outputs(1698) <= not a;
    layer2_outputs(1699) <= a and b;
    layer2_outputs(1700) <= '1';
    layer2_outputs(1701) <= not a;
    layer2_outputs(1702) <= not (a or b);
    layer2_outputs(1703) <= '1';
    layer2_outputs(1704) <= not (a and b);
    layer2_outputs(1705) <= a;
    layer2_outputs(1706) <= a or b;
    layer2_outputs(1707) <= not b;
    layer2_outputs(1708) <= a xor b;
    layer2_outputs(1709) <= not b;
    layer2_outputs(1710) <= a or b;
    layer2_outputs(1711) <= not a or b;
    layer2_outputs(1712) <= b;
    layer2_outputs(1713) <= not b;
    layer2_outputs(1714) <= not a or b;
    layer2_outputs(1715) <= a and not b;
    layer2_outputs(1716) <= a or b;
    layer2_outputs(1717) <= a and b;
    layer2_outputs(1718) <= a and b;
    layer2_outputs(1719) <= a and b;
    layer2_outputs(1720) <= b and not a;
    layer2_outputs(1721) <= b;
    layer2_outputs(1722) <= b;
    layer2_outputs(1723) <= not a or b;
    layer2_outputs(1724) <= b and not a;
    layer2_outputs(1725) <= a xor b;
    layer2_outputs(1726) <= not a;
    layer2_outputs(1727) <= a;
    layer2_outputs(1728) <= a and b;
    layer2_outputs(1729) <= not a;
    layer2_outputs(1730) <= a and not b;
    layer2_outputs(1731) <= not (a and b);
    layer2_outputs(1732) <= not a;
    layer2_outputs(1733) <= not b;
    layer2_outputs(1734) <= a xor b;
    layer2_outputs(1735) <= a;
    layer2_outputs(1736) <= not a or b;
    layer2_outputs(1737) <= '1';
    layer2_outputs(1738) <= a;
    layer2_outputs(1739) <= a and not b;
    layer2_outputs(1740) <= b;
    layer2_outputs(1741) <= b and not a;
    layer2_outputs(1742) <= not a;
    layer2_outputs(1743) <= not (a or b);
    layer2_outputs(1744) <= a;
    layer2_outputs(1745) <= a and not b;
    layer2_outputs(1746) <= not (a and b);
    layer2_outputs(1747) <= not a or b;
    layer2_outputs(1748) <= not b or a;
    layer2_outputs(1749) <= a;
    layer2_outputs(1750) <= a;
    layer2_outputs(1751) <= b;
    layer2_outputs(1752) <= '0';
    layer2_outputs(1753) <= not (a and b);
    layer2_outputs(1754) <= b;
    layer2_outputs(1755) <= b;
    layer2_outputs(1756) <= not b;
    layer2_outputs(1757) <= a or b;
    layer2_outputs(1758) <= not (a and b);
    layer2_outputs(1759) <= b;
    layer2_outputs(1760) <= a and b;
    layer2_outputs(1761) <= a;
    layer2_outputs(1762) <= a or b;
    layer2_outputs(1763) <= not a;
    layer2_outputs(1764) <= not (a xor b);
    layer2_outputs(1765) <= a and b;
    layer2_outputs(1766) <= a and not b;
    layer2_outputs(1767) <= not b;
    layer2_outputs(1768) <= a or b;
    layer2_outputs(1769) <= a and not b;
    layer2_outputs(1770) <= not a or b;
    layer2_outputs(1771) <= '0';
    layer2_outputs(1772) <= b;
    layer2_outputs(1773) <= a;
    layer2_outputs(1774) <= not a;
    layer2_outputs(1775) <= b;
    layer2_outputs(1776) <= not (a or b);
    layer2_outputs(1777) <= not a;
    layer2_outputs(1778) <= a and b;
    layer2_outputs(1779) <= a and not b;
    layer2_outputs(1780) <= a and b;
    layer2_outputs(1781) <= not b or a;
    layer2_outputs(1782) <= not a;
    layer2_outputs(1783) <= a;
    layer2_outputs(1784) <= a xor b;
    layer2_outputs(1785) <= a and b;
    layer2_outputs(1786) <= not b;
    layer2_outputs(1787) <= a xor b;
    layer2_outputs(1788) <= b;
    layer2_outputs(1789) <= not (a or b);
    layer2_outputs(1790) <= a and not b;
    layer2_outputs(1791) <= a and not b;
    layer2_outputs(1792) <= not b;
    layer2_outputs(1793) <= b;
    layer2_outputs(1794) <= not b;
    layer2_outputs(1795) <= a;
    layer2_outputs(1796) <= a;
    layer2_outputs(1797) <= b and not a;
    layer2_outputs(1798) <= '1';
    layer2_outputs(1799) <= a or b;
    layer2_outputs(1800) <= '0';
    layer2_outputs(1801) <= not (a or b);
    layer2_outputs(1802) <= not (a xor b);
    layer2_outputs(1803) <= not b;
    layer2_outputs(1804) <= a;
    layer2_outputs(1805) <= b and not a;
    layer2_outputs(1806) <= not a or b;
    layer2_outputs(1807) <= a and not b;
    layer2_outputs(1808) <= '1';
    layer2_outputs(1809) <= a;
    layer2_outputs(1810) <= a and b;
    layer2_outputs(1811) <= a or b;
    layer2_outputs(1812) <= a;
    layer2_outputs(1813) <= not b;
    layer2_outputs(1814) <= a xor b;
    layer2_outputs(1815) <= not a or b;
    layer2_outputs(1816) <= a or b;
    layer2_outputs(1817) <= not (a or b);
    layer2_outputs(1818) <= not b;
    layer2_outputs(1819) <= not a;
    layer2_outputs(1820) <= not b;
    layer2_outputs(1821) <= a xor b;
    layer2_outputs(1822) <= not (a or b);
    layer2_outputs(1823) <= not (a or b);
    layer2_outputs(1824) <= not a;
    layer2_outputs(1825) <= a and b;
    layer2_outputs(1826) <= a xor b;
    layer2_outputs(1827) <= not (a and b);
    layer2_outputs(1828) <= a xor b;
    layer2_outputs(1829) <= not b;
    layer2_outputs(1830) <= not b or a;
    layer2_outputs(1831) <= a;
    layer2_outputs(1832) <= a and not b;
    layer2_outputs(1833) <= b;
    layer2_outputs(1834) <= not b;
    layer2_outputs(1835) <= not (a xor b);
    layer2_outputs(1836) <= not b or a;
    layer2_outputs(1837) <= not (a xor b);
    layer2_outputs(1838) <= not a;
    layer2_outputs(1839) <= a and not b;
    layer2_outputs(1840) <= not b;
    layer2_outputs(1841) <= '0';
    layer2_outputs(1842) <= not a or b;
    layer2_outputs(1843) <= a or b;
    layer2_outputs(1844) <= a and b;
    layer2_outputs(1845) <= a and not b;
    layer2_outputs(1846) <= a and b;
    layer2_outputs(1847) <= not (a and b);
    layer2_outputs(1848) <= a;
    layer2_outputs(1849) <= not b;
    layer2_outputs(1850) <= not b;
    layer2_outputs(1851) <= not (a and b);
    layer2_outputs(1852) <= not b or a;
    layer2_outputs(1853) <= a and not b;
    layer2_outputs(1854) <= not (a or b);
    layer2_outputs(1855) <= not b or a;
    layer2_outputs(1856) <= not b or a;
    layer2_outputs(1857) <= b;
    layer2_outputs(1858) <= a and b;
    layer2_outputs(1859) <= not b;
    layer2_outputs(1860) <= not a or b;
    layer2_outputs(1861) <= b;
    layer2_outputs(1862) <= b and not a;
    layer2_outputs(1863) <= b and not a;
    layer2_outputs(1864) <= a;
    layer2_outputs(1865) <= not a;
    layer2_outputs(1866) <= not (a xor b);
    layer2_outputs(1867) <= not (a and b);
    layer2_outputs(1868) <= not a;
    layer2_outputs(1869) <= b and not a;
    layer2_outputs(1870) <= '0';
    layer2_outputs(1871) <= not (a xor b);
    layer2_outputs(1872) <= a and not b;
    layer2_outputs(1873) <= b;
    layer2_outputs(1874) <= a and not b;
    layer2_outputs(1875) <= '0';
    layer2_outputs(1876) <= a and not b;
    layer2_outputs(1877) <= b and not a;
    layer2_outputs(1878) <= not b;
    layer2_outputs(1879) <= a;
    layer2_outputs(1880) <= not (a and b);
    layer2_outputs(1881) <= '1';
    layer2_outputs(1882) <= b and not a;
    layer2_outputs(1883) <= a and b;
    layer2_outputs(1884) <= b;
    layer2_outputs(1885) <= not b;
    layer2_outputs(1886) <= a;
    layer2_outputs(1887) <= a or b;
    layer2_outputs(1888) <= b;
    layer2_outputs(1889) <= '1';
    layer2_outputs(1890) <= a;
    layer2_outputs(1891) <= not (a or b);
    layer2_outputs(1892) <= b;
    layer2_outputs(1893) <= a xor b;
    layer2_outputs(1894) <= '0';
    layer2_outputs(1895) <= b;
    layer2_outputs(1896) <= not b;
    layer2_outputs(1897) <= a and b;
    layer2_outputs(1898) <= a;
    layer2_outputs(1899) <= not a;
    layer2_outputs(1900) <= a xor b;
    layer2_outputs(1901) <= a;
    layer2_outputs(1902) <= not a;
    layer2_outputs(1903) <= b;
    layer2_outputs(1904) <= a;
    layer2_outputs(1905) <= '0';
    layer2_outputs(1906) <= not (a and b);
    layer2_outputs(1907) <= not a or b;
    layer2_outputs(1908) <= not a or b;
    layer2_outputs(1909) <= a and not b;
    layer2_outputs(1910) <= not a;
    layer2_outputs(1911) <= not (a or b);
    layer2_outputs(1912) <= a;
    layer2_outputs(1913) <= not a;
    layer2_outputs(1914) <= b and not a;
    layer2_outputs(1915) <= not b;
    layer2_outputs(1916) <= '1';
    layer2_outputs(1917) <= not a;
    layer2_outputs(1918) <= b and not a;
    layer2_outputs(1919) <= not (a xor b);
    layer2_outputs(1920) <= not a;
    layer2_outputs(1921) <= a xor b;
    layer2_outputs(1922) <= b;
    layer2_outputs(1923) <= a;
    layer2_outputs(1924) <= not (a or b);
    layer2_outputs(1925) <= a;
    layer2_outputs(1926) <= b;
    layer2_outputs(1927) <= a or b;
    layer2_outputs(1928) <= '0';
    layer2_outputs(1929) <= b;
    layer2_outputs(1930) <= a and b;
    layer2_outputs(1931) <= not b;
    layer2_outputs(1932) <= a and b;
    layer2_outputs(1933) <= not (a and b);
    layer2_outputs(1934) <= a or b;
    layer2_outputs(1935) <= b and not a;
    layer2_outputs(1936) <= not b;
    layer2_outputs(1937) <= not b;
    layer2_outputs(1938) <= a;
    layer2_outputs(1939) <= a and b;
    layer2_outputs(1940) <= not b or a;
    layer2_outputs(1941) <= b;
    layer2_outputs(1942) <= a or b;
    layer2_outputs(1943) <= not (a and b);
    layer2_outputs(1944) <= a;
    layer2_outputs(1945) <= '0';
    layer2_outputs(1946) <= not (a xor b);
    layer2_outputs(1947) <= a;
    layer2_outputs(1948) <= b;
    layer2_outputs(1949) <= a and b;
    layer2_outputs(1950) <= not b or a;
    layer2_outputs(1951) <= a and b;
    layer2_outputs(1952) <= not a;
    layer2_outputs(1953) <= '1';
    layer2_outputs(1954) <= not b or a;
    layer2_outputs(1955) <= not (a xor b);
    layer2_outputs(1956) <= not b;
    layer2_outputs(1957) <= b and not a;
    layer2_outputs(1958) <= '0';
    layer2_outputs(1959) <= a;
    layer2_outputs(1960) <= a and b;
    layer2_outputs(1961) <= a and b;
    layer2_outputs(1962) <= not b;
    layer2_outputs(1963) <= not a;
    layer2_outputs(1964) <= not (a or b);
    layer2_outputs(1965) <= not a;
    layer2_outputs(1966) <= a;
    layer2_outputs(1967) <= b and not a;
    layer2_outputs(1968) <= a and b;
    layer2_outputs(1969) <= not a;
    layer2_outputs(1970) <= b and not a;
    layer2_outputs(1971) <= not b;
    layer2_outputs(1972) <= not b;
    layer2_outputs(1973) <= not (a and b);
    layer2_outputs(1974) <= '0';
    layer2_outputs(1975) <= a and b;
    layer2_outputs(1976) <= a and not b;
    layer2_outputs(1977) <= not (a or b);
    layer2_outputs(1978) <= not b or a;
    layer2_outputs(1979) <= not a or b;
    layer2_outputs(1980) <= not (a and b);
    layer2_outputs(1981) <= b and not a;
    layer2_outputs(1982) <= not a or b;
    layer2_outputs(1983) <= not b;
    layer2_outputs(1984) <= b;
    layer2_outputs(1985) <= a and b;
    layer2_outputs(1986) <= a or b;
    layer2_outputs(1987) <= not b or a;
    layer2_outputs(1988) <= b;
    layer2_outputs(1989) <= not b or a;
    layer2_outputs(1990) <= not (a and b);
    layer2_outputs(1991) <= not (a and b);
    layer2_outputs(1992) <= not a;
    layer2_outputs(1993) <= not b;
    layer2_outputs(1994) <= not b;
    layer2_outputs(1995) <= not a;
    layer2_outputs(1996) <= not b or a;
    layer2_outputs(1997) <= a and b;
    layer2_outputs(1998) <= b;
    layer2_outputs(1999) <= a and b;
    layer2_outputs(2000) <= a xor b;
    layer2_outputs(2001) <= a or b;
    layer2_outputs(2002) <= b;
    layer2_outputs(2003) <= '1';
    layer2_outputs(2004) <= a and b;
    layer2_outputs(2005) <= '1';
    layer2_outputs(2006) <= b and not a;
    layer2_outputs(2007) <= a and b;
    layer2_outputs(2008) <= a;
    layer2_outputs(2009) <= not (a or b);
    layer2_outputs(2010) <= not b or a;
    layer2_outputs(2011) <= a xor b;
    layer2_outputs(2012) <= not b or a;
    layer2_outputs(2013) <= not a or b;
    layer2_outputs(2014) <= a and not b;
    layer2_outputs(2015) <= a or b;
    layer2_outputs(2016) <= b;
    layer2_outputs(2017) <= b;
    layer2_outputs(2018) <= not (a and b);
    layer2_outputs(2019) <= not a;
    layer2_outputs(2020) <= not a;
    layer2_outputs(2021) <= b and not a;
    layer2_outputs(2022) <= a and not b;
    layer2_outputs(2023) <= a or b;
    layer2_outputs(2024) <= not b;
    layer2_outputs(2025) <= a xor b;
    layer2_outputs(2026) <= a or b;
    layer2_outputs(2027) <= not (a or b);
    layer2_outputs(2028) <= b;
    layer2_outputs(2029) <= a and not b;
    layer2_outputs(2030) <= b;
    layer2_outputs(2031) <= '0';
    layer2_outputs(2032) <= a xor b;
    layer2_outputs(2033) <= a and not b;
    layer2_outputs(2034) <= not b;
    layer2_outputs(2035) <= not b;
    layer2_outputs(2036) <= not b;
    layer2_outputs(2037) <= b;
    layer2_outputs(2038) <= b;
    layer2_outputs(2039) <= not b;
    layer2_outputs(2040) <= not a or b;
    layer2_outputs(2041) <= not b or a;
    layer2_outputs(2042) <= not a;
    layer2_outputs(2043) <= not a or b;
    layer2_outputs(2044) <= a;
    layer2_outputs(2045) <= not a;
    layer2_outputs(2046) <= not b or a;
    layer2_outputs(2047) <= a and b;
    layer2_outputs(2048) <= not (a or b);
    layer2_outputs(2049) <= not b or a;
    layer2_outputs(2050) <= b;
    layer2_outputs(2051) <= b;
    layer2_outputs(2052) <= a or b;
    layer2_outputs(2053) <= a xor b;
    layer2_outputs(2054) <= a or b;
    layer2_outputs(2055) <= '0';
    layer2_outputs(2056) <= '1';
    layer2_outputs(2057) <= not b;
    layer2_outputs(2058) <= not b or a;
    layer2_outputs(2059) <= not a or b;
    layer2_outputs(2060) <= not b;
    layer2_outputs(2061) <= not b or a;
    layer2_outputs(2062) <= b;
    layer2_outputs(2063) <= not a;
    layer2_outputs(2064) <= a xor b;
    layer2_outputs(2065) <= not b;
    layer2_outputs(2066) <= a;
    layer2_outputs(2067) <= a and b;
    layer2_outputs(2068) <= a or b;
    layer2_outputs(2069) <= b;
    layer2_outputs(2070) <= a and b;
    layer2_outputs(2071) <= not (a or b);
    layer2_outputs(2072) <= not (a or b);
    layer2_outputs(2073) <= a xor b;
    layer2_outputs(2074) <= not (a or b);
    layer2_outputs(2075) <= not a or b;
    layer2_outputs(2076) <= b and not a;
    layer2_outputs(2077) <= not b or a;
    layer2_outputs(2078) <= not a;
    layer2_outputs(2079) <= b and not a;
    layer2_outputs(2080) <= a or b;
    layer2_outputs(2081) <= a;
    layer2_outputs(2082) <= b and not a;
    layer2_outputs(2083) <= not b or a;
    layer2_outputs(2084) <= not a;
    layer2_outputs(2085) <= a and b;
    layer2_outputs(2086) <= '1';
    layer2_outputs(2087) <= a or b;
    layer2_outputs(2088) <= a and not b;
    layer2_outputs(2089) <= a or b;
    layer2_outputs(2090) <= not a;
    layer2_outputs(2091) <= not b;
    layer2_outputs(2092) <= a;
    layer2_outputs(2093) <= a and b;
    layer2_outputs(2094) <= a;
    layer2_outputs(2095) <= not a;
    layer2_outputs(2096) <= not (a and b);
    layer2_outputs(2097) <= a and not b;
    layer2_outputs(2098) <= not a;
    layer2_outputs(2099) <= b and not a;
    layer2_outputs(2100) <= '1';
    layer2_outputs(2101) <= not a;
    layer2_outputs(2102) <= a;
    layer2_outputs(2103) <= b;
    layer2_outputs(2104) <= a xor b;
    layer2_outputs(2105) <= a or b;
    layer2_outputs(2106) <= a;
    layer2_outputs(2107) <= a and not b;
    layer2_outputs(2108) <= not b;
    layer2_outputs(2109) <= not a;
    layer2_outputs(2110) <= not a;
    layer2_outputs(2111) <= b;
    layer2_outputs(2112) <= a;
    layer2_outputs(2113) <= not b or a;
    layer2_outputs(2114) <= not (a xor b);
    layer2_outputs(2115) <= a xor b;
    layer2_outputs(2116) <= b;
    layer2_outputs(2117) <= a or b;
    layer2_outputs(2118) <= a and not b;
    layer2_outputs(2119) <= not a;
    layer2_outputs(2120) <= not (a or b);
    layer2_outputs(2121) <= a or b;
    layer2_outputs(2122) <= not b;
    layer2_outputs(2123) <= not b or a;
    layer2_outputs(2124) <= not a or b;
    layer2_outputs(2125) <= a or b;
    layer2_outputs(2126) <= not b;
    layer2_outputs(2127) <= b;
    layer2_outputs(2128) <= a;
    layer2_outputs(2129) <= a and b;
    layer2_outputs(2130) <= a xor b;
    layer2_outputs(2131) <= a and not b;
    layer2_outputs(2132) <= '1';
    layer2_outputs(2133) <= a;
    layer2_outputs(2134) <= '0';
    layer2_outputs(2135) <= not a or b;
    layer2_outputs(2136) <= a and b;
    layer2_outputs(2137) <= not (a or b);
    layer2_outputs(2138) <= not b or a;
    layer2_outputs(2139) <= not b;
    layer2_outputs(2140) <= not b or a;
    layer2_outputs(2141) <= not b or a;
    layer2_outputs(2142) <= a xor b;
    layer2_outputs(2143) <= a or b;
    layer2_outputs(2144) <= b;
    layer2_outputs(2145) <= a;
    layer2_outputs(2146) <= b;
    layer2_outputs(2147) <= not b or a;
    layer2_outputs(2148) <= b and not a;
    layer2_outputs(2149) <= not (a and b);
    layer2_outputs(2150) <= not (a or b);
    layer2_outputs(2151) <= not b;
    layer2_outputs(2152) <= not (a and b);
    layer2_outputs(2153) <= a xor b;
    layer2_outputs(2154) <= a or b;
    layer2_outputs(2155) <= not b or a;
    layer2_outputs(2156) <= b;
    layer2_outputs(2157) <= not b;
    layer2_outputs(2158) <= a;
    layer2_outputs(2159) <= not (a and b);
    layer2_outputs(2160) <= not (a and b);
    layer2_outputs(2161) <= not (a or b);
    layer2_outputs(2162) <= not (a xor b);
    layer2_outputs(2163) <= b;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= a;
    layer2_outputs(2166) <= b;
    layer2_outputs(2167) <= not b;
    layer2_outputs(2168) <= b;
    layer2_outputs(2169) <= a;
    layer2_outputs(2170) <= not (a xor b);
    layer2_outputs(2171) <= a or b;
    layer2_outputs(2172) <= b;
    layer2_outputs(2173) <= not (a and b);
    layer2_outputs(2174) <= not (a and b);
    layer2_outputs(2175) <= not (a xor b);
    layer2_outputs(2176) <= a;
    layer2_outputs(2177) <= b;
    layer2_outputs(2178) <= a;
    layer2_outputs(2179) <= a and not b;
    layer2_outputs(2180) <= a or b;
    layer2_outputs(2181) <= not (a xor b);
    layer2_outputs(2182) <= not (a and b);
    layer2_outputs(2183) <= not b;
    layer2_outputs(2184) <= not b;
    layer2_outputs(2185) <= not b;
    layer2_outputs(2186) <= not (a or b);
    layer2_outputs(2187) <= a and not b;
    layer2_outputs(2188) <= not (a or b);
    layer2_outputs(2189) <= not (a and b);
    layer2_outputs(2190) <= not a or b;
    layer2_outputs(2191) <= a;
    layer2_outputs(2192) <= a or b;
    layer2_outputs(2193) <= not b;
    layer2_outputs(2194) <= not a or b;
    layer2_outputs(2195) <= a and b;
    layer2_outputs(2196) <= not b;
    layer2_outputs(2197) <= b and not a;
    layer2_outputs(2198) <= a xor b;
    layer2_outputs(2199) <= not a;
    layer2_outputs(2200) <= a and not b;
    layer2_outputs(2201) <= a or b;
    layer2_outputs(2202) <= a;
    layer2_outputs(2203) <= not b;
    layer2_outputs(2204) <= not b;
    layer2_outputs(2205) <= a;
    layer2_outputs(2206) <= not a;
    layer2_outputs(2207) <= not b or a;
    layer2_outputs(2208) <= not (a xor b);
    layer2_outputs(2209) <= not (a or b);
    layer2_outputs(2210) <= not a or b;
    layer2_outputs(2211) <= a and not b;
    layer2_outputs(2212) <= not (a or b);
    layer2_outputs(2213) <= not b;
    layer2_outputs(2214) <= not (a and b);
    layer2_outputs(2215) <= a or b;
    layer2_outputs(2216) <= not (a and b);
    layer2_outputs(2217) <= a and not b;
    layer2_outputs(2218) <= a and not b;
    layer2_outputs(2219) <= a or b;
    layer2_outputs(2220) <= a and not b;
    layer2_outputs(2221) <= '1';
    layer2_outputs(2222) <= a and not b;
    layer2_outputs(2223) <= not a or b;
    layer2_outputs(2224) <= not (a and b);
    layer2_outputs(2225) <= not b;
    layer2_outputs(2226) <= not b;
    layer2_outputs(2227) <= not a;
    layer2_outputs(2228) <= not b or a;
    layer2_outputs(2229) <= not (a or b);
    layer2_outputs(2230) <= not a or b;
    layer2_outputs(2231) <= not a;
    layer2_outputs(2232) <= b;
    layer2_outputs(2233) <= a or b;
    layer2_outputs(2234) <= not (a and b);
    layer2_outputs(2235) <= '0';
    layer2_outputs(2236) <= not a or b;
    layer2_outputs(2237) <= a and b;
    layer2_outputs(2238) <= not b;
    layer2_outputs(2239) <= a and b;
    layer2_outputs(2240) <= a;
    layer2_outputs(2241) <= not a;
    layer2_outputs(2242) <= not (a and b);
    layer2_outputs(2243) <= '0';
    layer2_outputs(2244) <= not a;
    layer2_outputs(2245) <= not (a xor b);
    layer2_outputs(2246) <= not b or a;
    layer2_outputs(2247) <= not (a and b);
    layer2_outputs(2248) <= not b or a;
    layer2_outputs(2249) <= not a;
    layer2_outputs(2250) <= not b;
    layer2_outputs(2251) <= not (a and b);
    layer2_outputs(2252) <= a;
    layer2_outputs(2253) <= a;
    layer2_outputs(2254) <= not a;
    layer2_outputs(2255) <= '1';
    layer2_outputs(2256) <= not b or a;
    layer2_outputs(2257) <= a and b;
    layer2_outputs(2258) <= a and not b;
    layer2_outputs(2259) <= not (a xor b);
    layer2_outputs(2260) <= not a or b;
    layer2_outputs(2261) <= not (a and b);
    layer2_outputs(2262) <= '1';
    layer2_outputs(2263) <= a and not b;
    layer2_outputs(2264) <= a and not b;
    layer2_outputs(2265) <= b and not a;
    layer2_outputs(2266) <= not a or b;
    layer2_outputs(2267) <= a and not b;
    layer2_outputs(2268) <= b;
    layer2_outputs(2269) <= a;
    layer2_outputs(2270) <= not (a or b);
    layer2_outputs(2271) <= not (a and b);
    layer2_outputs(2272) <= a and not b;
    layer2_outputs(2273) <= a or b;
    layer2_outputs(2274) <= a and not b;
    layer2_outputs(2275) <= not a;
    layer2_outputs(2276) <= a;
    layer2_outputs(2277) <= not a;
    layer2_outputs(2278) <= not a or b;
    layer2_outputs(2279) <= not a;
    layer2_outputs(2280) <= not b or a;
    layer2_outputs(2281) <= not (a and b);
    layer2_outputs(2282) <= not a;
    layer2_outputs(2283) <= not a or b;
    layer2_outputs(2284) <= b;
    layer2_outputs(2285) <= not (a xor b);
    layer2_outputs(2286) <= '0';
    layer2_outputs(2287) <= not b or a;
    layer2_outputs(2288) <= a;
    layer2_outputs(2289) <= a;
    layer2_outputs(2290) <= a and b;
    layer2_outputs(2291) <= b;
    layer2_outputs(2292) <= a;
    layer2_outputs(2293) <= not (a and b);
    layer2_outputs(2294) <= '1';
    layer2_outputs(2295) <= not a or b;
    layer2_outputs(2296) <= not (a and b);
    layer2_outputs(2297) <= not (a and b);
    layer2_outputs(2298) <= b;
    layer2_outputs(2299) <= b and not a;
    layer2_outputs(2300) <= not a or b;
    layer2_outputs(2301) <= not a;
    layer2_outputs(2302) <= a and b;
    layer2_outputs(2303) <= not a;
    layer2_outputs(2304) <= '1';
    layer2_outputs(2305) <= b;
    layer2_outputs(2306) <= not a;
    layer2_outputs(2307) <= a and b;
    layer2_outputs(2308) <= not (a and b);
    layer2_outputs(2309) <= not b;
    layer2_outputs(2310) <= not a or b;
    layer2_outputs(2311) <= not b;
    layer2_outputs(2312) <= a and b;
    layer2_outputs(2313) <= b and not a;
    layer2_outputs(2314) <= a xor b;
    layer2_outputs(2315) <= '1';
    layer2_outputs(2316) <= a and b;
    layer2_outputs(2317) <= not (a xor b);
    layer2_outputs(2318) <= a;
    layer2_outputs(2319) <= not a or b;
    layer2_outputs(2320) <= b;
    layer2_outputs(2321) <= '0';
    layer2_outputs(2322) <= not (a xor b);
    layer2_outputs(2323) <= '1';
    layer2_outputs(2324) <= a and not b;
    layer2_outputs(2325) <= not (a or b);
    layer2_outputs(2326) <= not (a xor b);
    layer2_outputs(2327) <= not a;
    layer2_outputs(2328) <= a xor b;
    layer2_outputs(2329) <= a or b;
    layer2_outputs(2330) <= a or b;
    layer2_outputs(2331) <= not b;
    layer2_outputs(2332) <= b and not a;
    layer2_outputs(2333) <= not (a and b);
    layer2_outputs(2334) <= b and not a;
    layer2_outputs(2335) <= b and not a;
    layer2_outputs(2336) <= not a;
    layer2_outputs(2337) <= a or b;
    layer2_outputs(2338) <= not (a or b);
    layer2_outputs(2339) <= not a or b;
    layer2_outputs(2340) <= not a;
    layer2_outputs(2341) <= not (a or b);
    layer2_outputs(2342) <= a or b;
    layer2_outputs(2343) <= a and b;
    layer2_outputs(2344) <= not (a and b);
    layer2_outputs(2345) <= b and not a;
    layer2_outputs(2346) <= '1';
    layer2_outputs(2347) <= not b or a;
    layer2_outputs(2348) <= not (a and b);
    layer2_outputs(2349) <= not a;
    layer2_outputs(2350) <= not (a xor b);
    layer2_outputs(2351) <= a and not b;
    layer2_outputs(2352) <= a and b;
    layer2_outputs(2353) <= '1';
    layer2_outputs(2354) <= not b or a;
    layer2_outputs(2355) <= a;
    layer2_outputs(2356) <= not b or a;
    layer2_outputs(2357) <= not a or b;
    layer2_outputs(2358) <= b and not a;
    layer2_outputs(2359) <= not a;
    layer2_outputs(2360) <= not a or b;
    layer2_outputs(2361) <= not b or a;
    layer2_outputs(2362) <= b and not a;
    layer2_outputs(2363) <= b and not a;
    layer2_outputs(2364) <= a or b;
    layer2_outputs(2365) <= not (a or b);
    layer2_outputs(2366) <= a;
    layer2_outputs(2367) <= not a or b;
    layer2_outputs(2368) <= b and not a;
    layer2_outputs(2369) <= a;
    layer2_outputs(2370) <= not b or a;
    layer2_outputs(2371) <= b and not a;
    layer2_outputs(2372) <= '1';
    layer2_outputs(2373) <= '0';
    layer2_outputs(2374) <= not (a and b);
    layer2_outputs(2375) <= not b;
    layer2_outputs(2376) <= a and b;
    layer2_outputs(2377) <= b and not a;
    layer2_outputs(2378) <= a;
    layer2_outputs(2379) <= a and b;
    layer2_outputs(2380) <= a and not b;
    layer2_outputs(2381) <= not b;
    layer2_outputs(2382) <= a and not b;
    layer2_outputs(2383) <= not (a and b);
    layer2_outputs(2384) <= not a or b;
    layer2_outputs(2385) <= '1';
    layer2_outputs(2386) <= b and not a;
    layer2_outputs(2387) <= a or b;
    layer2_outputs(2388) <= a or b;
    layer2_outputs(2389) <= a xor b;
    layer2_outputs(2390) <= b and not a;
    layer2_outputs(2391) <= not (a or b);
    layer2_outputs(2392) <= not (a or b);
    layer2_outputs(2393) <= not a;
    layer2_outputs(2394) <= a;
    layer2_outputs(2395) <= not (a or b);
    layer2_outputs(2396) <= not (a and b);
    layer2_outputs(2397) <= a and not b;
    layer2_outputs(2398) <= not (a xor b);
    layer2_outputs(2399) <= a;
    layer2_outputs(2400) <= a xor b;
    layer2_outputs(2401) <= not b;
    layer2_outputs(2402) <= a and b;
    layer2_outputs(2403) <= not a or b;
    layer2_outputs(2404) <= a and not b;
    layer2_outputs(2405) <= a and b;
    layer2_outputs(2406) <= b and not a;
    layer2_outputs(2407) <= not (a or b);
    layer2_outputs(2408) <= b and not a;
    layer2_outputs(2409) <= b and not a;
    layer2_outputs(2410) <= a or b;
    layer2_outputs(2411) <= not (a or b);
    layer2_outputs(2412) <= b;
    layer2_outputs(2413) <= a;
    layer2_outputs(2414) <= not a;
    layer2_outputs(2415) <= a or b;
    layer2_outputs(2416) <= not a or b;
    layer2_outputs(2417) <= not b;
    layer2_outputs(2418) <= not b;
    layer2_outputs(2419) <= not a;
    layer2_outputs(2420) <= '1';
    layer2_outputs(2421) <= a;
    layer2_outputs(2422) <= not (a xor b);
    layer2_outputs(2423) <= not a;
    layer2_outputs(2424) <= a and not b;
    layer2_outputs(2425) <= b and not a;
    layer2_outputs(2426) <= not b or a;
    layer2_outputs(2427) <= '1';
    layer2_outputs(2428) <= a xor b;
    layer2_outputs(2429) <= not a or b;
    layer2_outputs(2430) <= '1';
    layer2_outputs(2431) <= b;
    layer2_outputs(2432) <= a and b;
    layer2_outputs(2433) <= not (a and b);
    layer2_outputs(2434) <= not a;
    layer2_outputs(2435) <= not b;
    layer2_outputs(2436) <= not b or a;
    layer2_outputs(2437) <= '1';
    layer2_outputs(2438) <= b;
    layer2_outputs(2439) <= not (a or b);
    layer2_outputs(2440) <= not b;
    layer2_outputs(2441) <= not a;
    layer2_outputs(2442) <= a;
    layer2_outputs(2443) <= a;
    layer2_outputs(2444) <= not b;
    layer2_outputs(2445) <= a and b;
    layer2_outputs(2446) <= a;
    layer2_outputs(2447) <= not a;
    layer2_outputs(2448) <= a or b;
    layer2_outputs(2449) <= a;
    layer2_outputs(2450) <= a and not b;
    layer2_outputs(2451) <= not b or a;
    layer2_outputs(2452) <= a and b;
    layer2_outputs(2453) <= not (a and b);
    layer2_outputs(2454) <= a and b;
    layer2_outputs(2455) <= b;
    layer2_outputs(2456) <= not b or a;
    layer2_outputs(2457) <= not (a and b);
    layer2_outputs(2458) <= not a;
    layer2_outputs(2459) <= not (a xor b);
    layer2_outputs(2460) <= a;
    layer2_outputs(2461) <= not (a and b);
    layer2_outputs(2462) <= not b;
    layer2_outputs(2463) <= not (a or b);
    layer2_outputs(2464) <= not (a or b);
    layer2_outputs(2465) <= not (a or b);
    layer2_outputs(2466) <= not b or a;
    layer2_outputs(2467) <= '0';
    layer2_outputs(2468) <= a and not b;
    layer2_outputs(2469) <= a or b;
    layer2_outputs(2470) <= b;
    layer2_outputs(2471) <= not a or b;
    layer2_outputs(2472) <= a xor b;
    layer2_outputs(2473) <= a;
    layer2_outputs(2474) <= a;
    layer2_outputs(2475) <= not b;
    layer2_outputs(2476) <= not a or b;
    layer2_outputs(2477) <= '0';
    layer2_outputs(2478) <= not (a and b);
    layer2_outputs(2479) <= not a;
    layer2_outputs(2480) <= a and not b;
    layer2_outputs(2481) <= b;
    layer2_outputs(2482) <= a;
    layer2_outputs(2483) <= a;
    layer2_outputs(2484) <= not b;
    layer2_outputs(2485) <= not (a xor b);
    layer2_outputs(2486) <= not (a or b);
    layer2_outputs(2487) <= a xor b;
    layer2_outputs(2488) <= not b;
    layer2_outputs(2489) <= not (a or b);
    layer2_outputs(2490) <= a or b;
    layer2_outputs(2491) <= '0';
    layer2_outputs(2492) <= a;
    layer2_outputs(2493) <= a and not b;
    layer2_outputs(2494) <= not (a or b);
    layer2_outputs(2495) <= a;
    layer2_outputs(2496) <= not b;
    layer2_outputs(2497) <= b and not a;
    layer2_outputs(2498) <= not a;
    layer2_outputs(2499) <= a;
    layer2_outputs(2500) <= b;
    layer2_outputs(2501) <= a and not b;
    layer2_outputs(2502) <= not b or a;
    layer2_outputs(2503) <= not (a and b);
    layer2_outputs(2504) <= not (a xor b);
    layer2_outputs(2505) <= not b or a;
    layer2_outputs(2506) <= a and not b;
    layer2_outputs(2507) <= not b or a;
    layer2_outputs(2508) <= not (a or b);
    layer2_outputs(2509) <= not a;
    layer2_outputs(2510) <= '1';
    layer2_outputs(2511) <= not a;
    layer2_outputs(2512) <= not a or b;
    layer2_outputs(2513) <= a;
    layer2_outputs(2514) <= not a or b;
    layer2_outputs(2515) <= not a;
    layer2_outputs(2516) <= b;
    layer2_outputs(2517) <= not b or a;
    layer2_outputs(2518) <= not (a and b);
    layer2_outputs(2519) <= not a;
    layer2_outputs(2520) <= b and not a;
    layer2_outputs(2521) <= not b;
    layer2_outputs(2522) <= not (a and b);
    layer2_outputs(2523) <= a;
    layer2_outputs(2524) <= not b or a;
    layer2_outputs(2525) <= a and b;
    layer2_outputs(2526) <= '1';
    layer2_outputs(2527) <= not a;
    layer2_outputs(2528) <= a;
    layer2_outputs(2529) <= a and not b;
    layer2_outputs(2530) <= not (a xor b);
    layer2_outputs(2531) <= not b;
    layer2_outputs(2532) <= not b or a;
    layer2_outputs(2533) <= not (a or b);
    layer2_outputs(2534) <= not (a or b);
    layer2_outputs(2535) <= not a or b;
    layer2_outputs(2536) <= not b or a;
    layer2_outputs(2537) <= a or b;
    layer2_outputs(2538) <= not (a xor b);
    layer2_outputs(2539) <= a;
    layer2_outputs(2540) <= not (a and b);
    layer2_outputs(2541) <= not b or a;
    layer2_outputs(2542) <= a;
    layer2_outputs(2543) <= not b;
    layer2_outputs(2544) <= not b;
    layer2_outputs(2545) <= not (a and b);
    layer2_outputs(2546) <= not a or b;
    layer2_outputs(2547) <= not b or a;
    layer2_outputs(2548) <= not a;
    layer2_outputs(2549) <= a;
    layer2_outputs(2550) <= not a;
    layer2_outputs(2551) <= a or b;
    layer2_outputs(2552) <= a and b;
    layer2_outputs(2553) <= a xor b;
    layer2_outputs(2554) <= not (a or b);
    layer2_outputs(2555) <= not b;
    layer2_outputs(2556) <= a or b;
    layer2_outputs(2557) <= not (a or b);
    layer2_outputs(2558) <= not (a or b);
    layer2_outputs(2559) <= a;
    layer2_outputs(2560) <= not a;
    layer2_outputs(2561) <= b and not a;
    layer2_outputs(2562) <= not a;
    layer2_outputs(2563) <= not a;
    layer2_outputs(2564) <= not a;
    layer2_outputs(2565) <= b;
    layer2_outputs(2566) <= not (a or b);
    layer2_outputs(2567) <= '0';
    layer2_outputs(2568) <= a or b;
    layer2_outputs(2569) <= not b;
    layer2_outputs(2570) <= b;
    layer2_outputs(2571) <= not b;
    layer2_outputs(2572) <= a;
    layer2_outputs(2573) <= a or b;
    layer2_outputs(2574) <= a and b;
    layer2_outputs(2575) <= '0';
    layer2_outputs(2576) <= not a;
    layer2_outputs(2577) <= b;
    layer2_outputs(2578) <= b and not a;
    layer2_outputs(2579) <= not b;
    layer2_outputs(2580) <= a;
    layer2_outputs(2581) <= a and not b;
    layer2_outputs(2582) <= a;
    layer2_outputs(2583) <= b;
    layer2_outputs(2584) <= not (a and b);
    layer2_outputs(2585) <= not b;
    layer2_outputs(2586) <= b;
    layer2_outputs(2587) <= a xor b;
    layer2_outputs(2588) <= a xor b;
    layer2_outputs(2589) <= not (a xor b);
    layer2_outputs(2590) <= a;
    layer2_outputs(2591) <= a;
    layer2_outputs(2592) <= b;
    layer2_outputs(2593) <= not b;
    layer2_outputs(2594) <= a or b;
    layer2_outputs(2595) <= not b or a;
    layer2_outputs(2596) <= not (a xor b);
    layer2_outputs(2597) <= not a or b;
    layer2_outputs(2598) <= a and not b;
    layer2_outputs(2599) <= a and b;
    layer2_outputs(2600) <= b and not a;
    layer2_outputs(2601) <= b;
    layer2_outputs(2602) <= '1';
    layer2_outputs(2603) <= b and not a;
    layer2_outputs(2604) <= a;
    layer2_outputs(2605) <= a and not b;
    layer2_outputs(2606) <= not (a or b);
    layer2_outputs(2607) <= a or b;
    layer2_outputs(2608) <= '1';
    layer2_outputs(2609) <= b;
    layer2_outputs(2610) <= not (a and b);
    layer2_outputs(2611) <= not b or a;
    layer2_outputs(2612) <= not a or b;
    layer2_outputs(2613) <= a and not b;
    layer2_outputs(2614) <= a;
    layer2_outputs(2615) <= not (a or b);
    layer2_outputs(2616) <= not a or b;
    layer2_outputs(2617) <= a and b;
    layer2_outputs(2618) <= not a;
    layer2_outputs(2619) <= b;
    layer2_outputs(2620) <= not (a and b);
    layer2_outputs(2621) <= not a;
    layer2_outputs(2622) <= not (a or b);
    layer2_outputs(2623) <= a and b;
    layer2_outputs(2624) <= b and not a;
    layer2_outputs(2625) <= not a;
    layer2_outputs(2626) <= b and not a;
    layer2_outputs(2627) <= not b or a;
    layer2_outputs(2628) <= not a or b;
    layer2_outputs(2629) <= not (a or b);
    layer2_outputs(2630) <= '0';
    layer2_outputs(2631) <= a or b;
    layer2_outputs(2632) <= a;
    layer2_outputs(2633) <= b and not a;
    layer2_outputs(2634) <= not a;
    layer2_outputs(2635) <= a xor b;
    layer2_outputs(2636) <= a or b;
    layer2_outputs(2637) <= a and not b;
    layer2_outputs(2638) <= a;
    layer2_outputs(2639) <= a;
    layer2_outputs(2640) <= a or b;
    layer2_outputs(2641) <= not a or b;
    layer2_outputs(2642) <= not a;
    layer2_outputs(2643) <= '1';
    layer2_outputs(2644) <= a;
    layer2_outputs(2645) <= a and not b;
    layer2_outputs(2646) <= not a or b;
    layer2_outputs(2647) <= not (a or b);
    layer2_outputs(2648) <= not (a and b);
    layer2_outputs(2649) <= not a;
    layer2_outputs(2650) <= b;
    layer2_outputs(2651) <= '0';
    layer2_outputs(2652) <= not a or b;
    layer2_outputs(2653) <= a or b;
    layer2_outputs(2654) <= '0';
    layer2_outputs(2655) <= b;
    layer2_outputs(2656) <= a and not b;
    layer2_outputs(2657) <= not b;
    layer2_outputs(2658) <= a;
    layer2_outputs(2659) <= b and not a;
    layer2_outputs(2660) <= not b;
    layer2_outputs(2661) <= not (a and b);
    layer2_outputs(2662) <= not (a xor b);
    layer2_outputs(2663) <= not a;
    layer2_outputs(2664) <= not a or b;
    layer2_outputs(2665) <= a xor b;
    layer2_outputs(2666) <= a;
    layer2_outputs(2667) <= a and not b;
    layer2_outputs(2668) <= not a or b;
    layer2_outputs(2669) <= not a;
    layer2_outputs(2670) <= not b;
    layer2_outputs(2671) <= not a or b;
    layer2_outputs(2672) <= not b;
    layer2_outputs(2673) <= a and not b;
    layer2_outputs(2674) <= a or b;
    layer2_outputs(2675) <= a and not b;
    layer2_outputs(2676) <= a and not b;
    layer2_outputs(2677) <= not (a or b);
    layer2_outputs(2678) <= not b;
    layer2_outputs(2679) <= a or b;
    layer2_outputs(2680) <= '0';
    layer2_outputs(2681) <= a and not b;
    layer2_outputs(2682) <= a xor b;
    layer2_outputs(2683) <= not (a or b);
    layer2_outputs(2684) <= not b;
    layer2_outputs(2685) <= a and not b;
    layer2_outputs(2686) <= not (a or b);
    layer2_outputs(2687) <= '1';
    layer2_outputs(2688) <= a and not b;
    layer2_outputs(2689) <= a;
    layer2_outputs(2690) <= a or b;
    layer2_outputs(2691) <= '0';
    layer2_outputs(2692) <= not a;
    layer2_outputs(2693) <= a xor b;
    layer2_outputs(2694) <= not b;
    layer2_outputs(2695) <= not (a and b);
    layer2_outputs(2696) <= a;
    layer2_outputs(2697) <= not (a xor b);
    layer2_outputs(2698) <= not b or a;
    layer2_outputs(2699) <= b;
    layer2_outputs(2700) <= '0';
    layer2_outputs(2701) <= a or b;
    layer2_outputs(2702) <= not b or a;
    layer2_outputs(2703) <= a;
    layer2_outputs(2704) <= '0';
    layer2_outputs(2705) <= a and b;
    layer2_outputs(2706) <= not (a or b);
    layer2_outputs(2707) <= not (a and b);
    layer2_outputs(2708) <= not (a or b);
    layer2_outputs(2709) <= b;
    layer2_outputs(2710) <= not b;
    layer2_outputs(2711) <= a xor b;
    layer2_outputs(2712) <= not a or b;
    layer2_outputs(2713) <= not a or b;
    layer2_outputs(2714) <= not (a or b);
    layer2_outputs(2715) <= not b;
    layer2_outputs(2716) <= not a;
    layer2_outputs(2717) <= not (a xor b);
    layer2_outputs(2718) <= a and not b;
    layer2_outputs(2719) <= b and not a;
    layer2_outputs(2720) <= not a or b;
    layer2_outputs(2721) <= a and b;
    layer2_outputs(2722) <= not a or b;
    layer2_outputs(2723) <= not (a xor b);
    layer2_outputs(2724) <= b and not a;
    layer2_outputs(2725) <= a and not b;
    layer2_outputs(2726) <= not (a or b);
    layer2_outputs(2727) <= not b;
    layer2_outputs(2728) <= a;
    layer2_outputs(2729) <= a;
    layer2_outputs(2730) <= b and not a;
    layer2_outputs(2731) <= b and not a;
    layer2_outputs(2732) <= not (a or b);
    layer2_outputs(2733) <= b and not a;
    layer2_outputs(2734) <= not b;
    layer2_outputs(2735) <= not b;
    layer2_outputs(2736) <= a and not b;
    layer2_outputs(2737) <= b;
    layer2_outputs(2738) <= not b or a;
    layer2_outputs(2739) <= a and not b;
    layer2_outputs(2740) <= not (a or b);
    layer2_outputs(2741) <= not b or a;
    layer2_outputs(2742) <= '0';
    layer2_outputs(2743) <= b;
    layer2_outputs(2744) <= not (a or b);
    layer2_outputs(2745) <= a;
    layer2_outputs(2746) <= not (a or b);
    layer2_outputs(2747) <= a or b;
    layer2_outputs(2748) <= '1';
    layer2_outputs(2749) <= a and not b;
    layer2_outputs(2750) <= not (a xor b);
    layer2_outputs(2751) <= not (a and b);
    layer2_outputs(2752) <= not b;
    layer2_outputs(2753) <= a xor b;
    layer2_outputs(2754) <= not b;
    layer2_outputs(2755) <= not b or a;
    layer2_outputs(2756) <= '0';
    layer2_outputs(2757) <= a;
    layer2_outputs(2758) <= not a;
    layer2_outputs(2759) <= b and not a;
    layer2_outputs(2760) <= not (a or b);
    layer2_outputs(2761) <= not a or b;
    layer2_outputs(2762) <= not a;
    layer2_outputs(2763) <= not a;
    layer2_outputs(2764) <= b;
    layer2_outputs(2765) <= not a;
    layer2_outputs(2766) <= a or b;
    layer2_outputs(2767) <= not (a or b);
    layer2_outputs(2768) <= a xor b;
    layer2_outputs(2769) <= not a;
    layer2_outputs(2770) <= not (a and b);
    layer2_outputs(2771) <= not (a and b);
    layer2_outputs(2772) <= b;
    layer2_outputs(2773) <= a and b;
    layer2_outputs(2774) <= not b or a;
    layer2_outputs(2775) <= a xor b;
    layer2_outputs(2776) <= not (a xor b);
    layer2_outputs(2777) <= not a or b;
    layer2_outputs(2778) <= '1';
    layer2_outputs(2779) <= not a;
    layer2_outputs(2780) <= not (a xor b);
    layer2_outputs(2781) <= b;
    layer2_outputs(2782) <= a and not b;
    layer2_outputs(2783) <= not b or a;
    layer2_outputs(2784) <= not a or b;
    layer2_outputs(2785) <= not (a or b);
    layer2_outputs(2786) <= not b;
    layer2_outputs(2787) <= '0';
    layer2_outputs(2788) <= not (a or b);
    layer2_outputs(2789) <= a and not b;
    layer2_outputs(2790) <= not a;
    layer2_outputs(2791) <= not b;
    layer2_outputs(2792) <= a xor b;
    layer2_outputs(2793) <= not b;
    layer2_outputs(2794) <= '0';
    layer2_outputs(2795) <= not (a or b);
    layer2_outputs(2796) <= b;
    layer2_outputs(2797) <= a;
    layer2_outputs(2798) <= a and b;
    layer2_outputs(2799) <= b;
    layer2_outputs(2800) <= not a or b;
    layer2_outputs(2801) <= not b;
    layer2_outputs(2802) <= not a or b;
    layer2_outputs(2803) <= not b or a;
    layer2_outputs(2804) <= not (a and b);
    layer2_outputs(2805) <= not (a or b);
    layer2_outputs(2806) <= a and not b;
    layer2_outputs(2807) <= '1';
    layer2_outputs(2808) <= a and b;
    layer2_outputs(2809) <= not a;
    layer2_outputs(2810) <= not (a and b);
    layer2_outputs(2811) <= not a or b;
    layer2_outputs(2812) <= a and not b;
    layer2_outputs(2813) <= not a;
    layer2_outputs(2814) <= a;
    layer2_outputs(2815) <= not a;
    layer2_outputs(2816) <= '1';
    layer2_outputs(2817) <= not (a or b);
    layer2_outputs(2818) <= a or b;
    layer2_outputs(2819) <= a;
    layer2_outputs(2820) <= a xor b;
    layer2_outputs(2821) <= a;
    layer2_outputs(2822) <= a;
    layer2_outputs(2823) <= not b or a;
    layer2_outputs(2824) <= not (a or b);
    layer2_outputs(2825) <= a;
    layer2_outputs(2826) <= b and not a;
    layer2_outputs(2827) <= not b or a;
    layer2_outputs(2828) <= not (a or b);
    layer2_outputs(2829) <= a and b;
    layer2_outputs(2830) <= a and b;
    layer2_outputs(2831) <= not a or b;
    layer2_outputs(2832) <= a and not b;
    layer2_outputs(2833) <= not (a or b);
    layer2_outputs(2834) <= not (a and b);
    layer2_outputs(2835) <= not b or a;
    layer2_outputs(2836) <= b and not a;
    layer2_outputs(2837) <= not b;
    layer2_outputs(2838) <= b and not a;
    layer2_outputs(2839) <= not b or a;
    layer2_outputs(2840) <= a or b;
    layer2_outputs(2841) <= not (a or b);
    layer2_outputs(2842) <= not b or a;
    layer2_outputs(2843) <= a and not b;
    layer2_outputs(2844) <= b;
    layer2_outputs(2845) <= a or b;
    layer2_outputs(2846) <= not (a and b);
    layer2_outputs(2847) <= a or b;
    layer2_outputs(2848) <= a or b;
    layer2_outputs(2849) <= a or b;
    layer2_outputs(2850) <= a or b;
    layer2_outputs(2851) <= not b;
    layer2_outputs(2852) <= not a;
    layer2_outputs(2853) <= not b;
    layer2_outputs(2854) <= '0';
    layer2_outputs(2855) <= a and b;
    layer2_outputs(2856) <= a or b;
    layer2_outputs(2857) <= not a;
    layer2_outputs(2858) <= not (a or b);
    layer2_outputs(2859) <= a;
    layer2_outputs(2860) <= b;
    layer2_outputs(2861) <= not b or a;
    layer2_outputs(2862) <= a and not b;
    layer2_outputs(2863) <= a xor b;
    layer2_outputs(2864) <= not b or a;
    layer2_outputs(2865) <= b;
    layer2_outputs(2866) <= not a or b;
    layer2_outputs(2867) <= b;
    layer2_outputs(2868) <= not b;
    layer2_outputs(2869) <= a and b;
    layer2_outputs(2870) <= not a;
    layer2_outputs(2871) <= not (a or b);
    layer2_outputs(2872) <= a and b;
    layer2_outputs(2873) <= not (a or b);
    layer2_outputs(2874) <= not a or b;
    layer2_outputs(2875) <= '1';
    layer2_outputs(2876) <= a and b;
    layer2_outputs(2877) <= '1';
    layer2_outputs(2878) <= not a;
    layer2_outputs(2879) <= b;
    layer2_outputs(2880) <= not (a xor b);
    layer2_outputs(2881) <= not a or b;
    layer2_outputs(2882) <= a and not b;
    layer2_outputs(2883) <= b;
    layer2_outputs(2884) <= b and not a;
    layer2_outputs(2885) <= b and not a;
    layer2_outputs(2886) <= b;
    layer2_outputs(2887) <= not b;
    layer2_outputs(2888) <= not b or a;
    layer2_outputs(2889) <= a;
    layer2_outputs(2890) <= a and not b;
    layer2_outputs(2891) <= a or b;
    layer2_outputs(2892) <= '1';
    layer2_outputs(2893) <= not b or a;
    layer2_outputs(2894) <= b and not a;
    layer2_outputs(2895) <= b;
    layer2_outputs(2896) <= a and b;
    layer2_outputs(2897) <= not a;
    layer2_outputs(2898) <= not a;
    layer2_outputs(2899) <= a and b;
    layer2_outputs(2900) <= not a or b;
    layer2_outputs(2901) <= not a;
    layer2_outputs(2902) <= not a or b;
    layer2_outputs(2903) <= a;
    layer2_outputs(2904) <= a;
    layer2_outputs(2905) <= b;
    layer2_outputs(2906) <= '1';
    layer2_outputs(2907) <= a;
    layer2_outputs(2908) <= a or b;
    layer2_outputs(2909) <= a;
    layer2_outputs(2910) <= '0';
    layer2_outputs(2911) <= not (a xor b);
    layer2_outputs(2912) <= not b;
    layer2_outputs(2913) <= b and not a;
    layer2_outputs(2914) <= not b;
    layer2_outputs(2915) <= b;
    layer2_outputs(2916) <= not (a and b);
    layer2_outputs(2917) <= not (a and b);
    layer2_outputs(2918) <= not (a xor b);
    layer2_outputs(2919) <= '0';
    layer2_outputs(2920) <= not (a or b);
    layer2_outputs(2921) <= not b or a;
    layer2_outputs(2922) <= not a;
    layer2_outputs(2923) <= not a or b;
    layer2_outputs(2924) <= b;
    layer2_outputs(2925) <= not a or b;
    layer2_outputs(2926) <= not (a or b);
    layer2_outputs(2927) <= not a;
    layer2_outputs(2928) <= b;
    layer2_outputs(2929) <= '1';
    layer2_outputs(2930) <= b;
    layer2_outputs(2931) <= b;
    layer2_outputs(2932) <= b;
    layer2_outputs(2933) <= not b or a;
    layer2_outputs(2934) <= not b;
    layer2_outputs(2935) <= a and not b;
    layer2_outputs(2936) <= a;
    layer2_outputs(2937) <= not b or a;
    layer2_outputs(2938) <= not a;
    layer2_outputs(2939) <= not (a or b);
    layer2_outputs(2940) <= a and not b;
    layer2_outputs(2941) <= a or b;
    layer2_outputs(2942) <= a and not b;
    layer2_outputs(2943) <= not b;
    layer2_outputs(2944) <= '0';
    layer2_outputs(2945) <= a;
    layer2_outputs(2946) <= not b or a;
    layer2_outputs(2947) <= a and b;
    layer2_outputs(2948) <= a xor b;
    layer2_outputs(2949) <= a xor b;
    layer2_outputs(2950) <= a;
    layer2_outputs(2951) <= b and not a;
    layer2_outputs(2952) <= not (a and b);
    layer2_outputs(2953) <= not a;
    layer2_outputs(2954) <= a and b;
    layer2_outputs(2955) <= b;
    layer2_outputs(2956) <= not (a and b);
    layer2_outputs(2957) <= not (a xor b);
    layer2_outputs(2958) <= not b;
    layer2_outputs(2959) <= b;
    layer2_outputs(2960) <= b and not a;
    layer2_outputs(2961) <= not a;
    layer2_outputs(2962) <= a and b;
    layer2_outputs(2963) <= b;
    layer2_outputs(2964) <= a or b;
    layer2_outputs(2965) <= not (a and b);
    layer2_outputs(2966) <= not (a or b);
    layer2_outputs(2967) <= not a;
    layer2_outputs(2968) <= '1';
    layer2_outputs(2969) <= a or b;
    layer2_outputs(2970) <= a and b;
    layer2_outputs(2971) <= not b or a;
    layer2_outputs(2972) <= not a or b;
    layer2_outputs(2973) <= not (a or b);
    layer2_outputs(2974) <= not (a xor b);
    layer2_outputs(2975) <= not b or a;
    layer2_outputs(2976) <= b;
    layer2_outputs(2977) <= b;
    layer2_outputs(2978) <= a and b;
    layer2_outputs(2979) <= b and not a;
    layer2_outputs(2980) <= not b or a;
    layer2_outputs(2981) <= a and not b;
    layer2_outputs(2982) <= b;
    layer2_outputs(2983) <= not (a or b);
    layer2_outputs(2984) <= a and b;
    layer2_outputs(2985) <= not (a and b);
    layer2_outputs(2986) <= not (a or b);
    layer2_outputs(2987) <= not b;
    layer2_outputs(2988) <= not (a and b);
    layer2_outputs(2989) <= not b;
    layer2_outputs(2990) <= not a or b;
    layer2_outputs(2991) <= not a or b;
    layer2_outputs(2992) <= b and not a;
    layer2_outputs(2993) <= not (a and b);
    layer2_outputs(2994) <= not (a and b);
    layer2_outputs(2995) <= a and not b;
    layer2_outputs(2996) <= a and not b;
    layer2_outputs(2997) <= a and not b;
    layer2_outputs(2998) <= a and not b;
    layer2_outputs(2999) <= b;
    layer2_outputs(3000) <= not b or a;
    layer2_outputs(3001) <= not (a or b);
    layer2_outputs(3002) <= not (a xor b);
    layer2_outputs(3003) <= '1';
    layer2_outputs(3004) <= a and not b;
    layer2_outputs(3005) <= '1';
    layer2_outputs(3006) <= not b;
    layer2_outputs(3007) <= a;
    layer2_outputs(3008) <= not (a or b);
    layer2_outputs(3009) <= not (a or b);
    layer2_outputs(3010) <= a;
    layer2_outputs(3011) <= a;
    layer2_outputs(3012) <= a and not b;
    layer2_outputs(3013) <= b;
    layer2_outputs(3014) <= a or b;
    layer2_outputs(3015) <= not (a and b);
    layer2_outputs(3016) <= a;
    layer2_outputs(3017) <= not a or b;
    layer2_outputs(3018) <= not a or b;
    layer2_outputs(3019) <= not (a or b);
    layer2_outputs(3020) <= a and not b;
    layer2_outputs(3021) <= not (a and b);
    layer2_outputs(3022) <= not a or b;
    layer2_outputs(3023) <= a and not b;
    layer2_outputs(3024) <= a and b;
    layer2_outputs(3025) <= a;
    layer2_outputs(3026) <= '1';
    layer2_outputs(3027) <= not (a xor b);
    layer2_outputs(3028) <= a and not b;
    layer2_outputs(3029) <= not (a xor b);
    layer2_outputs(3030) <= not (a and b);
    layer2_outputs(3031) <= b;
    layer2_outputs(3032) <= '1';
    layer2_outputs(3033) <= not (a and b);
    layer2_outputs(3034) <= a xor b;
    layer2_outputs(3035) <= not (a or b);
    layer2_outputs(3036) <= not a or b;
    layer2_outputs(3037) <= not b;
    layer2_outputs(3038) <= a;
    layer2_outputs(3039) <= not (a and b);
    layer2_outputs(3040) <= not a;
    layer2_outputs(3041) <= '0';
    layer2_outputs(3042) <= a and not b;
    layer2_outputs(3043) <= b and not a;
    layer2_outputs(3044) <= a and not b;
    layer2_outputs(3045) <= not (a and b);
    layer2_outputs(3046) <= a or b;
    layer2_outputs(3047) <= not (a or b);
    layer2_outputs(3048) <= not a or b;
    layer2_outputs(3049) <= not (a and b);
    layer2_outputs(3050) <= not a or b;
    layer2_outputs(3051) <= not b;
    layer2_outputs(3052) <= not a or b;
    layer2_outputs(3053) <= a;
    layer2_outputs(3054) <= not b;
    layer2_outputs(3055) <= b;
    layer2_outputs(3056) <= not b;
    layer2_outputs(3057) <= a and not b;
    layer2_outputs(3058) <= not b;
    layer2_outputs(3059) <= not b or a;
    layer2_outputs(3060) <= not (a or b);
    layer2_outputs(3061) <= not (a and b);
    layer2_outputs(3062) <= not a;
    layer2_outputs(3063) <= a or b;
    layer2_outputs(3064) <= a or b;
    layer2_outputs(3065) <= not (a and b);
    layer2_outputs(3066) <= a;
    layer2_outputs(3067) <= a;
    layer2_outputs(3068) <= not a;
    layer2_outputs(3069) <= a or b;
    layer2_outputs(3070) <= not a;
    layer2_outputs(3071) <= b and not a;
    layer2_outputs(3072) <= not (a xor b);
    layer2_outputs(3073) <= not (a or b);
    layer2_outputs(3074) <= a;
    layer2_outputs(3075) <= b;
    layer2_outputs(3076) <= not b or a;
    layer2_outputs(3077) <= a and b;
    layer2_outputs(3078) <= a and not b;
    layer2_outputs(3079) <= not a or b;
    layer2_outputs(3080) <= b and not a;
    layer2_outputs(3081) <= not a or b;
    layer2_outputs(3082) <= a and b;
    layer2_outputs(3083) <= a or b;
    layer2_outputs(3084) <= a and not b;
    layer2_outputs(3085) <= a and not b;
    layer2_outputs(3086) <= not (a xor b);
    layer2_outputs(3087) <= b and not a;
    layer2_outputs(3088) <= not a;
    layer2_outputs(3089) <= b;
    layer2_outputs(3090) <= not (a or b);
    layer2_outputs(3091) <= b;
    layer2_outputs(3092) <= b and not a;
    layer2_outputs(3093) <= not (a or b);
    layer2_outputs(3094) <= b;
    layer2_outputs(3095) <= '1';
    layer2_outputs(3096) <= b and not a;
    layer2_outputs(3097) <= not b;
    layer2_outputs(3098) <= a;
    layer2_outputs(3099) <= '0';
    layer2_outputs(3100) <= not (a or b);
    layer2_outputs(3101) <= a and not b;
    layer2_outputs(3102) <= not a or b;
    layer2_outputs(3103) <= a;
    layer2_outputs(3104) <= b and not a;
    layer2_outputs(3105) <= a xor b;
    layer2_outputs(3106) <= not (a or b);
    layer2_outputs(3107) <= a;
    layer2_outputs(3108) <= not (a and b);
    layer2_outputs(3109) <= not (a and b);
    layer2_outputs(3110) <= not (a and b);
    layer2_outputs(3111) <= not (a or b);
    layer2_outputs(3112) <= not b;
    layer2_outputs(3113) <= not b or a;
    layer2_outputs(3114) <= not a or b;
    layer2_outputs(3115) <= not b or a;
    layer2_outputs(3116) <= a and not b;
    layer2_outputs(3117) <= a;
    layer2_outputs(3118) <= not (a or b);
    layer2_outputs(3119) <= not a;
    layer2_outputs(3120) <= not a or b;
    layer2_outputs(3121) <= b;
    layer2_outputs(3122) <= a;
    layer2_outputs(3123) <= a and not b;
    layer2_outputs(3124) <= '1';
    layer2_outputs(3125) <= b;
    layer2_outputs(3126) <= a and not b;
    layer2_outputs(3127) <= not b or a;
    layer2_outputs(3128) <= not b;
    layer2_outputs(3129) <= not (a or b);
    layer2_outputs(3130) <= not b;
    layer2_outputs(3131) <= b;
    layer2_outputs(3132) <= not b;
    layer2_outputs(3133) <= a and b;
    layer2_outputs(3134) <= a or b;
    layer2_outputs(3135) <= a and b;
    layer2_outputs(3136) <= not a;
    layer2_outputs(3137) <= not (a and b);
    layer2_outputs(3138) <= a and not b;
    layer2_outputs(3139) <= not (a or b);
    layer2_outputs(3140) <= a or b;
    layer2_outputs(3141) <= a xor b;
    layer2_outputs(3142) <= b;
    layer2_outputs(3143) <= a or b;
    layer2_outputs(3144) <= not b;
    layer2_outputs(3145) <= '1';
    layer2_outputs(3146) <= not (a and b);
    layer2_outputs(3147) <= not (a xor b);
    layer2_outputs(3148) <= not (a or b);
    layer2_outputs(3149) <= not a or b;
    layer2_outputs(3150) <= not (a or b);
    layer2_outputs(3151) <= b;
    layer2_outputs(3152) <= not a;
    layer2_outputs(3153) <= not (a xor b);
    layer2_outputs(3154) <= not b;
    layer2_outputs(3155) <= a and not b;
    layer2_outputs(3156) <= not b;
    layer2_outputs(3157) <= not (a xor b);
    layer2_outputs(3158) <= a and not b;
    layer2_outputs(3159) <= a;
    layer2_outputs(3160) <= a and not b;
    layer2_outputs(3161) <= not (a or b);
    layer2_outputs(3162) <= a xor b;
    layer2_outputs(3163) <= not b;
    layer2_outputs(3164) <= a xor b;
    layer2_outputs(3165) <= b;
    layer2_outputs(3166) <= not b;
    layer2_outputs(3167) <= b;
    layer2_outputs(3168) <= a and b;
    layer2_outputs(3169) <= a;
    layer2_outputs(3170) <= a or b;
    layer2_outputs(3171) <= not a or b;
    layer2_outputs(3172) <= not b or a;
    layer2_outputs(3173) <= a and b;
    layer2_outputs(3174) <= not b;
    layer2_outputs(3175) <= not b or a;
    layer2_outputs(3176) <= not (a and b);
    layer2_outputs(3177) <= a;
    layer2_outputs(3178) <= not b or a;
    layer2_outputs(3179) <= not b or a;
    layer2_outputs(3180) <= not (a and b);
    layer2_outputs(3181) <= b;
    layer2_outputs(3182) <= not b or a;
    layer2_outputs(3183) <= a;
    layer2_outputs(3184) <= a and b;
    layer2_outputs(3185) <= a and b;
    layer2_outputs(3186) <= not a;
    layer2_outputs(3187) <= not a;
    layer2_outputs(3188) <= not b;
    layer2_outputs(3189) <= a and b;
    layer2_outputs(3190) <= a or b;
    layer2_outputs(3191) <= not (a and b);
    layer2_outputs(3192) <= not (a and b);
    layer2_outputs(3193) <= not b or a;
    layer2_outputs(3194) <= a and b;
    layer2_outputs(3195) <= not (a or b);
    layer2_outputs(3196) <= '0';
    layer2_outputs(3197) <= not b;
    layer2_outputs(3198) <= not b;
    layer2_outputs(3199) <= not a or b;
    layer2_outputs(3200) <= not a;
    layer2_outputs(3201) <= not b;
    layer2_outputs(3202) <= a;
    layer2_outputs(3203) <= b;
    layer2_outputs(3204) <= not a or b;
    layer2_outputs(3205) <= not a or b;
    layer2_outputs(3206) <= b and not a;
    layer2_outputs(3207) <= not (a and b);
    layer2_outputs(3208) <= not (a or b);
    layer2_outputs(3209) <= not (a and b);
    layer2_outputs(3210) <= not a;
    layer2_outputs(3211) <= a and b;
    layer2_outputs(3212) <= b;
    layer2_outputs(3213) <= not b;
    layer2_outputs(3214) <= b and not a;
    layer2_outputs(3215) <= a or b;
    layer2_outputs(3216) <= a or b;
    layer2_outputs(3217) <= a and not b;
    layer2_outputs(3218) <= not b;
    layer2_outputs(3219) <= '1';
    layer2_outputs(3220) <= '0';
    layer2_outputs(3221) <= a;
    layer2_outputs(3222) <= a;
    layer2_outputs(3223) <= b and not a;
    layer2_outputs(3224) <= not a;
    layer2_outputs(3225) <= not b;
    layer2_outputs(3226) <= '1';
    layer2_outputs(3227) <= b and not a;
    layer2_outputs(3228) <= not (a or b);
    layer2_outputs(3229) <= not b;
    layer2_outputs(3230) <= b;
    layer2_outputs(3231) <= not (a or b);
    layer2_outputs(3232) <= a;
    layer2_outputs(3233) <= '0';
    layer2_outputs(3234) <= not a;
    layer2_outputs(3235) <= not a;
    layer2_outputs(3236) <= not b;
    layer2_outputs(3237) <= b and not a;
    layer2_outputs(3238) <= not a;
    layer2_outputs(3239) <= a and b;
    layer2_outputs(3240) <= b and not a;
    layer2_outputs(3241) <= a;
    layer2_outputs(3242) <= not (a and b);
    layer2_outputs(3243) <= not a;
    layer2_outputs(3244) <= a or b;
    layer2_outputs(3245) <= a and b;
    layer2_outputs(3246) <= a or b;
    layer2_outputs(3247) <= b;
    layer2_outputs(3248) <= a and b;
    layer2_outputs(3249) <= not (a and b);
    layer2_outputs(3250) <= b and not a;
    layer2_outputs(3251) <= not b;
    layer2_outputs(3252) <= not a;
    layer2_outputs(3253) <= a and not b;
    layer2_outputs(3254) <= not a;
    layer2_outputs(3255) <= a and b;
    layer2_outputs(3256) <= a;
    layer2_outputs(3257) <= b and not a;
    layer2_outputs(3258) <= a xor b;
    layer2_outputs(3259) <= not a;
    layer2_outputs(3260) <= a or b;
    layer2_outputs(3261) <= a and not b;
    layer2_outputs(3262) <= not b or a;
    layer2_outputs(3263) <= a and b;
    layer2_outputs(3264) <= a;
    layer2_outputs(3265) <= b and not a;
    layer2_outputs(3266) <= b and not a;
    layer2_outputs(3267) <= a and b;
    layer2_outputs(3268) <= a;
    layer2_outputs(3269) <= a and b;
    layer2_outputs(3270) <= not a;
    layer2_outputs(3271) <= a and not b;
    layer2_outputs(3272) <= a;
    layer2_outputs(3273) <= not b or a;
    layer2_outputs(3274) <= b;
    layer2_outputs(3275) <= a and not b;
    layer2_outputs(3276) <= '1';
    layer2_outputs(3277) <= not b;
    layer2_outputs(3278) <= a;
    layer2_outputs(3279) <= '0';
    layer2_outputs(3280) <= a;
    layer2_outputs(3281) <= not b or a;
    layer2_outputs(3282) <= a;
    layer2_outputs(3283) <= not (a xor b);
    layer2_outputs(3284) <= not a or b;
    layer2_outputs(3285) <= not b or a;
    layer2_outputs(3286) <= b;
    layer2_outputs(3287) <= b and not a;
    layer2_outputs(3288) <= a or b;
    layer2_outputs(3289) <= not (a or b);
    layer2_outputs(3290) <= a and b;
    layer2_outputs(3291) <= a and not b;
    layer2_outputs(3292) <= not b;
    layer2_outputs(3293) <= a or b;
    layer2_outputs(3294) <= a and b;
    layer2_outputs(3295) <= not a or b;
    layer2_outputs(3296) <= not a;
    layer2_outputs(3297) <= not b or a;
    layer2_outputs(3298) <= not (a and b);
    layer2_outputs(3299) <= a and b;
    layer2_outputs(3300) <= not b;
    layer2_outputs(3301) <= not a;
    layer2_outputs(3302) <= not b;
    layer2_outputs(3303) <= not (a or b);
    layer2_outputs(3304) <= a;
    layer2_outputs(3305) <= a and b;
    layer2_outputs(3306) <= a or b;
    layer2_outputs(3307) <= '0';
    layer2_outputs(3308) <= not a or b;
    layer2_outputs(3309) <= b;
    layer2_outputs(3310) <= a;
    layer2_outputs(3311) <= a and not b;
    layer2_outputs(3312) <= a and b;
    layer2_outputs(3313) <= a xor b;
    layer2_outputs(3314) <= not a;
    layer2_outputs(3315) <= not b;
    layer2_outputs(3316) <= a and b;
    layer2_outputs(3317) <= not a or b;
    layer2_outputs(3318) <= a and not b;
    layer2_outputs(3319) <= not a or b;
    layer2_outputs(3320) <= a or b;
    layer2_outputs(3321) <= not a or b;
    layer2_outputs(3322) <= a;
    layer2_outputs(3323) <= not a;
    layer2_outputs(3324) <= b and not a;
    layer2_outputs(3325) <= not b or a;
    layer2_outputs(3326) <= b and not a;
    layer2_outputs(3327) <= a;
    layer2_outputs(3328) <= a and not b;
    layer2_outputs(3329) <= not b;
    layer2_outputs(3330) <= b;
    layer2_outputs(3331) <= not (a and b);
    layer2_outputs(3332) <= a and b;
    layer2_outputs(3333) <= not b or a;
    layer2_outputs(3334) <= a xor b;
    layer2_outputs(3335) <= not (a and b);
    layer2_outputs(3336) <= a;
    layer2_outputs(3337) <= not b;
    layer2_outputs(3338) <= not a or b;
    layer2_outputs(3339) <= not (a and b);
    layer2_outputs(3340) <= b and not a;
    layer2_outputs(3341) <= b;
    layer2_outputs(3342) <= b;
    layer2_outputs(3343) <= a and not b;
    layer2_outputs(3344) <= a;
    layer2_outputs(3345) <= b;
    layer2_outputs(3346) <= not a or b;
    layer2_outputs(3347) <= not a;
    layer2_outputs(3348) <= not b or a;
    layer2_outputs(3349) <= a;
    layer2_outputs(3350) <= not (a and b);
    layer2_outputs(3351) <= b and not a;
    layer2_outputs(3352) <= '1';
    layer2_outputs(3353) <= not b or a;
    layer2_outputs(3354) <= a or b;
    layer2_outputs(3355) <= not a or b;
    layer2_outputs(3356) <= b;
    layer2_outputs(3357) <= not a or b;
    layer2_outputs(3358) <= not b;
    layer2_outputs(3359) <= a and b;
    layer2_outputs(3360) <= a;
    layer2_outputs(3361) <= a and b;
    layer2_outputs(3362) <= not a or b;
    layer2_outputs(3363) <= a and b;
    layer2_outputs(3364) <= a and not b;
    layer2_outputs(3365) <= a;
    layer2_outputs(3366) <= a and not b;
    layer2_outputs(3367) <= not a;
    layer2_outputs(3368) <= a;
    layer2_outputs(3369) <= not (a or b);
    layer2_outputs(3370) <= not b;
    layer2_outputs(3371) <= a and not b;
    layer2_outputs(3372) <= a and b;
    layer2_outputs(3373) <= a and not b;
    layer2_outputs(3374) <= b;
    layer2_outputs(3375) <= not a;
    layer2_outputs(3376) <= not (a xor b);
    layer2_outputs(3377) <= a or b;
    layer2_outputs(3378) <= a and b;
    layer2_outputs(3379) <= a and b;
    layer2_outputs(3380) <= not b;
    layer2_outputs(3381) <= a;
    layer2_outputs(3382) <= a or b;
    layer2_outputs(3383) <= not a or b;
    layer2_outputs(3384) <= not b or a;
    layer2_outputs(3385) <= a and b;
    layer2_outputs(3386) <= a xor b;
    layer2_outputs(3387) <= not a;
    layer2_outputs(3388) <= not (a and b);
    layer2_outputs(3389) <= not a;
    layer2_outputs(3390) <= not b;
    layer2_outputs(3391) <= a;
    layer2_outputs(3392) <= not (a and b);
    layer2_outputs(3393) <= a and not b;
    layer2_outputs(3394) <= not (a and b);
    layer2_outputs(3395) <= not b;
    layer2_outputs(3396) <= not (a and b);
    layer2_outputs(3397) <= not a or b;
    layer2_outputs(3398) <= '0';
    layer2_outputs(3399) <= '0';
    layer2_outputs(3400) <= not a or b;
    layer2_outputs(3401) <= '0';
    layer2_outputs(3402) <= '1';
    layer2_outputs(3403) <= '1';
    layer2_outputs(3404) <= not b;
    layer2_outputs(3405) <= '0';
    layer2_outputs(3406) <= a xor b;
    layer2_outputs(3407) <= not b or a;
    layer2_outputs(3408) <= a or b;
    layer2_outputs(3409) <= not a;
    layer2_outputs(3410) <= not a;
    layer2_outputs(3411) <= not a;
    layer2_outputs(3412) <= a;
    layer2_outputs(3413) <= not a or b;
    layer2_outputs(3414) <= a;
    layer2_outputs(3415) <= not b;
    layer2_outputs(3416) <= a and not b;
    layer2_outputs(3417) <= not b;
    layer2_outputs(3418) <= not a or b;
    layer2_outputs(3419) <= a and not b;
    layer2_outputs(3420) <= '0';
    layer2_outputs(3421) <= a or b;
    layer2_outputs(3422) <= a and b;
    layer2_outputs(3423) <= not (a or b);
    layer2_outputs(3424) <= not (a and b);
    layer2_outputs(3425) <= b;
    layer2_outputs(3426) <= b and not a;
    layer2_outputs(3427) <= a;
    layer2_outputs(3428) <= not b;
    layer2_outputs(3429) <= a;
    layer2_outputs(3430) <= b and not a;
    layer2_outputs(3431) <= a and not b;
    layer2_outputs(3432) <= a xor b;
    layer2_outputs(3433) <= not (a and b);
    layer2_outputs(3434) <= a;
    layer2_outputs(3435) <= not b or a;
    layer2_outputs(3436) <= not (a or b);
    layer2_outputs(3437) <= not b;
    layer2_outputs(3438) <= b;
    layer2_outputs(3439) <= a and not b;
    layer2_outputs(3440) <= a;
    layer2_outputs(3441) <= a xor b;
    layer2_outputs(3442) <= not a;
    layer2_outputs(3443) <= not (a and b);
    layer2_outputs(3444) <= '1';
    layer2_outputs(3445) <= a and b;
    layer2_outputs(3446) <= a and b;
    layer2_outputs(3447) <= not a or b;
    layer2_outputs(3448) <= a xor b;
    layer2_outputs(3449) <= a or b;
    layer2_outputs(3450) <= not b or a;
    layer2_outputs(3451) <= b and not a;
    layer2_outputs(3452) <= a;
    layer2_outputs(3453) <= not (a xor b);
    layer2_outputs(3454) <= '0';
    layer2_outputs(3455) <= not (a or b);
    layer2_outputs(3456) <= not a;
    layer2_outputs(3457) <= a;
    layer2_outputs(3458) <= not a;
    layer2_outputs(3459) <= not b;
    layer2_outputs(3460) <= not b or a;
    layer2_outputs(3461) <= b;
    layer2_outputs(3462) <= a or b;
    layer2_outputs(3463) <= not b;
    layer2_outputs(3464) <= not a;
    layer2_outputs(3465) <= a or b;
    layer2_outputs(3466) <= a or b;
    layer2_outputs(3467) <= not b;
    layer2_outputs(3468) <= not a or b;
    layer2_outputs(3469) <= a and not b;
    layer2_outputs(3470) <= not b;
    layer2_outputs(3471) <= b and not a;
    layer2_outputs(3472) <= not b or a;
    layer2_outputs(3473) <= not b;
    layer2_outputs(3474) <= b;
    layer2_outputs(3475) <= b and not a;
    layer2_outputs(3476) <= b and not a;
    layer2_outputs(3477) <= b;
    layer2_outputs(3478) <= b;
    layer2_outputs(3479) <= not a;
    layer2_outputs(3480) <= b and not a;
    layer2_outputs(3481) <= b and not a;
    layer2_outputs(3482) <= not b or a;
    layer2_outputs(3483) <= not a or b;
    layer2_outputs(3484) <= not b or a;
    layer2_outputs(3485) <= a;
    layer2_outputs(3486) <= a and b;
    layer2_outputs(3487) <= a and b;
    layer2_outputs(3488) <= not a;
    layer2_outputs(3489) <= not b;
    layer2_outputs(3490) <= a and b;
    layer2_outputs(3491) <= a;
    layer2_outputs(3492) <= a xor b;
    layer2_outputs(3493) <= not a;
    layer2_outputs(3494) <= not (a or b);
    layer2_outputs(3495) <= not b;
    layer2_outputs(3496) <= a;
    layer2_outputs(3497) <= a and not b;
    layer2_outputs(3498) <= a and b;
    layer2_outputs(3499) <= a;
    layer2_outputs(3500) <= not b or a;
    layer2_outputs(3501) <= b;
    layer2_outputs(3502) <= not (a or b);
    layer2_outputs(3503) <= not a;
    layer2_outputs(3504) <= b;
    layer2_outputs(3505) <= not a or b;
    layer2_outputs(3506) <= a or b;
    layer2_outputs(3507) <= '1';
    layer2_outputs(3508) <= a;
    layer2_outputs(3509) <= a;
    layer2_outputs(3510) <= not b;
    layer2_outputs(3511) <= b and not a;
    layer2_outputs(3512) <= not a or b;
    layer2_outputs(3513) <= a or b;
    layer2_outputs(3514) <= not b;
    layer2_outputs(3515) <= not (a or b);
    layer2_outputs(3516) <= a;
    layer2_outputs(3517) <= a or b;
    layer2_outputs(3518) <= a and b;
    layer2_outputs(3519) <= not b or a;
    layer2_outputs(3520) <= a and b;
    layer2_outputs(3521) <= a;
    layer2_outputs(3522) <= b;
    layer2_outputs(3523) <= b and not a;
    layer2_outputs(3524) <= not (a xor b);
    layer2_outputs(3525) <= a;
    layer2_outputs(3526) <= '1';
    layer2_outputs(3527) <= not (a and b);
    layer2_outputs(3528) <= not b or a;
    layer2_outputs(3529) <= not b or a;
    layer2_outputs(3530) <= not b or a;
    layer2_outputs(3531) <= not (a or b);
    layer2_outputs(3532) <= '0';
    layer2_outputs(3533) <= a or b;
    layer2_outputs(3534) <= '0';
    layer2_outputs(3535) <= not (a xor b);
    layer2_outputs(3536) <= a;
    layer2_outputs(3537) <= not a;
    layer2_outputs(3538) <= a and b;
    layer2_outputs(3539) <= not (a or b);
    layer2_outputs(3540) <= not (a and b);
    layer2_outputs(3541) <= b;
    layer2_outputs(3542) <= not (a and b);
    layer2_outputs(3543) <= not a;
    layer2_outputs(3544) <= b and not a;
    layer2_outputs(3545) <= not b or a;
    layer2_outputs(3546) <= not b or a;
    layer2_outputs(3547) <= a and b;
    layer2_outputs(3548) <= b;
    layer2_outputs(3549) <= not a;
    layer2_outputs(3550) <= not (a and b);
    layer2_outputs(3551) <= not b or a;
    layer2_outputs(3552) <= not (a and b);
    layer2_outputs(3553) <= a;
    layer2_outputs(3554) <= a or b;
    layer2_outputs(3555) <= b and not a;
    layer2_outputs(3556) <= '1';
    layer2_outputs(3557) <= a and b;
    layer2_outputs(3558) <= '1';
    layer2_outputs(3559) <= not b;
    layer2_outputs(3560) <= a and not b;
    layer2_outputs(3561) <= not (a or b);
    layer2_outputs(3562) <= not a;
    layer2_outputs(3563) <= '1';
    layer2_outputs(3564) <= a xor b;
    layer2_outputs(3565) <= not b or a;
    layer2_outputs(3566) <= not a;
    layer2_outputs(3567) <= a;
    layer2_outputs(3568) <= not b;
    layer2_outputs(3569) <= not b;
    layer2_outputs(3570) <= '1';
    layer2_outputs(3571) <= not a;
    layer2_outputs(3572) <= not a;
    layer2_outputs(3573) <= not b;
    layer2_outputs(3574) <= a;
    layer2_outputs(3575) <= not (a or b);
    layer2_outputs(3576) <= not a or b;
    layer2_outputs(3577) <= not (a and b);
    layer2_outputs(3578) <= not a;
    layer2_outputs(3579) <= not b;
    layer2_outputs(3580) <= not (a xor b);
    layer2_outputs(3581) <= not b;
    layer2_outputs(3582) <= a and not b;
    layer2_outputs(3583) <= a and b;
    layer2_outputs(3584) <= a and b;
    layer2_outputs(3585) <= b;
    layer2_outputs(3586) <= a xor b;
    layer2_outputs(3587) <= not b or a;
    layer2_outputs(3588) <= not b;
    layer2_outputs(3589) <= a;
    layer2_outputs(3590) <= not a;
    layer2_outputs(3591) <= not a;
    layer2_outputs(3592) <= a or b;
    layer2_outputs(3593) <= not a or b;
    layer2_outputs(3594) <= not b or a;
    layer2_outputs(3595) <= not b;
    layer2_outputs(3596) <= not a;
    layer2_outputs(3597) <= not b;
    layer2_outputs(3598) <= a or b;
    layer2_outputs(3599) <= not a;
    layer2_outputs(3600) <= b;
    layer2_outputs(3601) <= not a or b;
    layer2_outputs(3602) <= a and b;
    layer2_outputs(3603) <= b and not a;
    layer2_outputs(3604) <= b;
    layer2_outputs(3605) <= '0';
    layer2_outputs(3606) <= not a or b;
    layer2_outputs(3607) <= a;
    layer2_outputs(3608) <= a and b;
    layer2_outputs(3609) <= not (a xor b);
    layer2_outputs(3610) <= a or b;
    layer2_outputs(3611) <= b;
    layer2_outputs(3612) <= a and not b;
    layer2_outputs(3613) <= a and b;
    layer2_outputs(3614) <= not (a or b);
    layer2_outputs(3615) <= not a or b;
    layer2_outputs(3616) <= b;
    layer2_outputs(3617) <= not a;
    layer2_outputs(3618) <= a xor b;
    layer2_outputs(3619) <= b;
    layer2_outputs(3620) <= b;
    layer2_outputs(3621) <= not a;
    layer2_outputs(3622) <= not b or a;
    layer2_outputs(3623) <= '1';
    layer2_outputs(3624) <= a xor b;
    layer2_outputs(3625) <= not b;
    layer2_outputs(3626) <= not (a or b);
    layer2_outputs(3627) <= not a or b;
    layer2_outputs(3628) <= b;
    layer2_outputs(3629) <= '1';
    layer2_outputs(3630) <= a and b;
    layer2_outputs(3631) <= a or b;
    layer2_outputs(3632) <= a and b;
    layer2_outputs(3633) <= a xor b;
    layer2_outputs(3634) <= a and b;
    layer2_outputs(3635) <= a;
    layer2_outputs(3636) <= b;
    layer2_outputs(3637) <= b;
    layer2_outputs(3638) <= not a or b;
    layer2_outputs(3639) <= not (a and b);
    layer2_outputs(3640) <= a and not b;
    layer2_outputs(3641) <= a;
    layer2_outputs(3642) <= not a or b;
    layer2_outputs(3643) <= not b;
    layer2_outputs(3644) <= not b;
    layer2_outputs(3645) <= a xor b;
    layer2_outputs(3646) <= not b or a;
    layer2_outputs(3647) <= a;
    layer2_outputs(3648) <= not b or a;
    layer2_outputs(3649) <= b and not a;
    layer2_outputs(3650) <= not b;
    layer2_outputs(3651) <= not b or a;
    layer2_outputs(3652) <= not (a or b);
    layer2_outputs(3653) <= b;
    layer2_outputs(3654) <= not a or b;
    layer2_outputs(3655) <= a;
    layer2_outputs(3656) <= '0';
    layer2_outputs(3657) <= a or b;
    layer2_outputs(3658) <= not (a xor b);
    layer2_outputs(3659) <= not a or b;
    layer2_outputs(3660) <= not (a xor b);
    layer2_outputs(3661) <= not a or b;
    layer2_outputs(3662) <= a and b;
    layer2_outputs(3663) <= not (a xor b);
    layer2_outputs(3664) <= not a or b;
    layer2_outputs(3665) <= not (a or b);
    layer2_outputs(3666) <= not b or a;
    layer2_outputs(3667) <= not (a or b);
    layer2_outputs(3668) <= a;
    layer2_outputs(3669) <= a;
    layer2_outputs(3670) <= not b or a;
    layer2_outputs(3671) <= a and b;
    layer2_outputs(3672) <= not (a or b);
    layer2_outputs(3673) <= a;
    layer2_outputs(3674) <= a;
    layer2_outputs(3675) <= not (a or b);
    layer2_outputs(3676) <= not a or b;
    layer2_outputs(3677) <= not (a or b);
    layer2_outputs(3678) <= a;
    layer2_outputs(3679) <= b and not a;
    layer2_outputs(3680) <= not b;
    layer2_outputs(3681) <= not (a or b);
    layer2_outputs(3682) <= '1';
    layer2_outputs(3683) <= a;
    layer2_outputs(3684) <= not b or a;
    layer2_outputs(3685) <= b;
    layer2_outputs(3686) <= b and not a;
    layer2_outputs(3687) <= b;
    layer2_outputs(3688) <= not b;
    layer2_outputs(3689) <= b;
    layer2_outputs(3690) <= a and not b;
    layer2_outputs(3691) <= not a or b;
    layer2_outputs(3692) <= not b or a;
    layer2_outputs(3693) <= not (a and b);
    layer2_outputs(3694) <= a or b;
    layer2_outputs(3695) <= '1';
    layer2_outputs(3696) <= not b or a;
    layer2_outputs(3697) <= a;
    layer2_outputs(3698) <= not b;
    layer2_outputs(3699) <= b and not a;
    layer2_outputs(3700) <= a;
    layer2_outputs(3701) <= not b or a;
    layer2_outputs(3702) <= not (a or b);
    layer2_outputs(3703) <= not a or b;
    layer2_outputs(3704) <= a and not b;
    layer2_outputs(3705) <= not b;
    layer2_outputs(3706) <= not b;
    layer2_outputs(3707) <= not b;
    layer2_outputs(3708) <= not b;
    layer2_outputs(3709) <= not a;
    layer2_outputs(3710) <= a;
    layer2_outputs(3711) <= not b;
    layer2_outputs(3712) <= b;
    layer2_outputs(3713) <= not b;
    layer2_outputs(3714) <= not (a and b);
    layer2_outputs(3715) <= not b or a;
    layer2_outputs(3716) <= a or b;
    layer2_outputs(3717) <= not b or a;
    layer2_outputs(3718) <= not b;
    layer2_outputs(3719) <= a or b;
    layer2_outputs(3720) <= not b;
    layer2_outputs(3721) <= not a or b;
    layer2_outputs(3722) <= not (a and b);
    layer2_outputs(3723) <= a or b;
    layer2_outputs(3724) <= not a or b;
    layer2_outputs(3725) <= not (a xor b);
    layer2_outputs(3726) <= not b;
    layer2_outputs(3727) <= a;
    layer2_outputs(3728) <= not a or b;
    layer2_outputs(3729) <= a xor b;
    layer2_outputs(3730) <= '1';
    layer2_outputs(3731) <= not a;
    layer2_outputs(3732) <= b and not a;
    layer2_outputs(3733) <= '0';
    layer2_outputs(3734) <= not a or b;
    layer2_outputs(3735) <= not (a xor b);
    layer2_outputs(3736) <= '0';
    layer2_outputs(3737) <= not b;
    layer2_outputs(3738) <= not (a xor b);
    layer2_outputs(3739) <= a;
    layer2_outputs(3740) <= b and not a;
    layer2_outputs(3741) <= not a;
    layer2_outputs(3742) <= not a;
    layer2_outputs(3743) <= a or b;
    layer2_outputs(3744) <= a or b;
    layer2_outputs(3745) <= '1';
    layer2_outputs(3746) <= not b or a;
    layer2_outputs(3747) <= not b;
    layer2_outputs(3748) <= not a or b;
    layer2_outputs(3749) <= b;
    layer2_outputs(3750) <= a and b;
    layer2_outputs(3751) <= a;
    layer2_outputs(3752) <= not b;
    layer2_outputs(3753) <= a or b;
    layer2_outputs(3754) <= a and not b;
    layer2_outputs(3755) <= a and b;
    layer2_outputs(3756) <= not a;
    layer2_outputs(3757) <= b and not a;
    layer2_outputs(3758) <= a xor b;
    layer2_outputs(3759) <= b;
    layer2_outputs(3760) <= a and b;
    layer2_outputs(3761) <= a xor b;
    layer2_outputs(3762) <= a and b;
    layer2_outputs(3763) <= b;
    layer2_outputs(3764) <= a or b;
    layer2_outputs(3765) <= a;
    layer2_outputs(3766) <= a;
    layer2_outputs(3767) <= not b or a;
    layer2_outputs(3768) <= not a or b;
    layer2_outputs(3769) <= not b or a;
    layer2_outputs(3770) <= not (a or b);
    layer2_outputs(3771) <= not b;
    layer2_outputs(3772) <= a and not b;
    layer2_outputs(3773) <= not b or a;
    layer2_outputs(3774) <= not (a and b);
    layer2_outputs(3775) <= b and not a;
    layer2_outputs(3776) <= not a or b;
    layer2_outputs(3777) <= a;
    layer2_outputs(3778) <= not b;
    layer2_outputs(3779) <= b;
    layer2_outputs(3780) <= not b;
    layer2_outputs(3781) <= not a;
    layer2_outputs(3782) <= not a;
    layer2_outputs(3783) <= b;
    layer2_outputs(3784) <= a or b;
    layer2_outputs(3785) <= not (a and b);
    layer2_outputs(3786) <= a or b;
    layer2_outputs(3787) <= a and b;
    layer2_outputs(3788) <= a and b;
    layer2_outputs(3789) <= a;
    layer2_outputs(3790) <= a;
    layer2_outputs(3791) <= b;
    layer2_outputs(3792) <= a;
    layer2_outputs(3793) <= b and not a;
    layer2_outputs(3794) <= b and not a;
    layer2_outputs(3795) <= not a;
    layer2_outputs(3796) <= not a;
    layer2_outputs(3797) <= not b or a;
    layer2_outputs(3798) <= a or b;
    layer2_outputs(3799) <= b;
    layer2_outputs(3800) <= not a;
    layer2_outputs(3801) <= b;
    layer2_outputs(3802) <= not (a and b);
    layer2_outputs(3803) <= not (a or b);
    layer2_outputs(3804) <= b;
    layer2_outputs(3805) <= a or b;
    layer2_outputs(3806) <= not b;
    layer2_outputs(3807) <= b and not a;
    layer2_outputs(3808) <= not a or b;
    layer2_outputs(3809) <= not (a or b);
    layer2_outputs(3810) <= not a or b;
    layer2_outputs(3811) <= not (a xor b);
    layer2_outputs(3812) <= not (a or b);
    layer2_outputs(3813) <= not (a and b);
    layer2_outputs(3814) <= b;
    layer2_outputs(3815) <= a and not b;
    layer2_outputs(3816) <= '0';
    layer2_outputs(3817) <= not b;
    layer2_outputs(3818) <= a and b;
    layer2_outputs(3819) <= not (a or b);
    layer2_outputs(3820) <= b;
    layer2_outputs(3821) <= not b;
    layer2_outputs(3822) <= a;
    layer2_outputs(3823) <= not b or a;
    layer2_outputs(3824) <= '0';
    layer2_outputs(3825) <= b;
    layer2_outputs(3826) <= a and not b;
    layer2_outputs(3827) <= not a or b;
    layer2_outputs(3828) <= not a or b;
    layer2_outputs(3829) <= b and not a;
    layer2_outputs(3830) <= not b;
    layer2_outputs(3831) <= not b or a;
    layer2_outputs(3832) <= '1';
    layer2_outputs(3833) <= a;
    layer2_outputs(3834) <= a;
    layer2_outputs(3835) <= a and b;
    layer2_outputs(3836) <= '0';
    layer2_outputs(3837) <= b and not a;
    layer2_outputs(3838) <= not (a xor b);
    layer2_outputs(3839) <= a and b;
    layer2_outputs(3840) <= not a;
    layer2_outputs(3841) <= b and not a;
    layer2_outputs(3842) <= a;
    layer2_outputs(3843) <= not (a and b);
    layer2_outputs(3844) <= a and b;
    layer2_outputs(3845) <= not a or b;
    layer2_outputs(3846) <= not b;
    layer2_outputs(3847) <= a;
    layer2_outputs(3848) <= a;
    layer2_outputs(3849) <= b;
    layer2_outputs(3850) <= not b or a;
    layer2_outputs(3851) <= a and not b;
    layer2_outputs(3852) <= '1';
    layer2_outputs(3853) <= not a or b;
    layer2_outputs(3854) <= a and b;
    layer2_outputs(3855) <= not (a or b);
    layer2_outputs(3856) <= a xor b;
    layer2_outputs(3857) <= b;
    layer2_outputs(3858) <= b;
    layer2_outputs(3859) <= a and b;
    layer2_outputs(3860) <= a;
    layer2_outputs(3861) <= not (a xor b);
    layer2_outputs(3862) <= b and not a;
    layer2_outputs(3863) <= not a or b;
    layer2_outputs(3864) <= a and not b;
    layer2_outputs(3865) <= b and not a;
    layer2_outputs(3866) <= not a;
    layer2_outputs(3867) <= '1';
    layer2_outputs(3868) <= not (a or b);
    layer2_outputs(3869) <= b;
    layer2_outputs(3870) <= not a;
    layer2_outputs(3871) <= not b;
    layer2_outputs(3872) <= a;
    layer2_outputs(3873) <= a and not b;
    layer2_outputs(3874) <= not (a and b);
    layer2_outputs(3875) <= a;
    layer2_outputs(3876) <= not (a or b);
    layer2_outputs(3877) <= a;
    layer2_outputs(3878) <= a or b;
    layer2_outputs(3879) <= a and b;
    layer2_outputs(3880) <= not a;
    layer2_outputs(3881) <= not b;
    layer2_outputs(3882) <= b;
    layer2_outputs(3883) <= b and not a;
    layer2_outputs(3884) <= not a;
    layer2_outputs(3885) <= a and b;
    layer2_outputs(3886) <= not a or b;
    layer2_outputs(3887) <= not b or a;
    layer2_outputs(3888) <= a;
    layer2_outputs(3889) <= not a or b;
    layer2_outputs(3890) <= a;
    layer2_outputs(3891) <= b;
    layer2_outputs(3892) <= b and not a;
    layer2_outputs(3893) <= not b;
    layer2_outputs(3894) <= not a;
    layer2_outputs(3895) <= '0';
    layer2_outputs(3896) <= a;
    layer2_outputs(3897) <= a;
    layer2_outputs(3898) <= a;
    layer2_outputs(3899) <= a and not b;
    layer2_outputs(3900) <= not a;
    layer2_outputs(3901) <= a;
    layer2_outputs(3902) <= not a;
    layer2_outputs(3903) <= not (a or b);
    layer2_outputs(3904) <= a and b;
    layer2_outputs(3905) <= a and b;
    layer2_outputs(3906) <= not (a and b);
    layer2_outputs(3907) <= not b or a;
    layer2_outputs(3908) <= not b;
    layer2_outputs(3909) <= not (a or b);
    layer2_outputs(3910) <= a;
    layer2_outputs(3911) <= a or b;
    layer2_outputs(3912) <= not (a and b);
    layer2_outputs(3913) <= '1';
    layer2_outputs(3914) <= a;
    layer2_outputs(3915) <= b and not a;
    layer2_outputs(3916) <= not a or b;
    layer2_outputs(3917) <= a and b;
    layer2_outputs(3918) <= b and not a;
    layer2_outputs(3919) <= not b;
    layer2_outputs(3920) <= not b;
    layer2_outputs(3921) <= a;
    layer2_outputs(3922) <= '0';
    layer2_outputs(3923) <= a and b;
    layer2_outputs(3924) <= not (a and b);
    layer2_outputs(3925) <= not a or b;
    layer2_outputs(3926) <= b and not a;
    layer2_outputs(3927) <= not a or b;
    layer2_outputs(3928) <= a and b;
    layer2_outputs(3929) <= not (a or b);
    layer2_outputs(3930) <= not (a and b);
    layer2_outputs(3931) <= not (a or b);
    layer2_outputs(3932) <= b and not a;
    layer2_outputs(3933) <= '1';
    layer2_outputs(3934) <= b;
    layer2_outputs(3935) <= '0';
    layer2_outputs(3936) <= not a;
    layer2_outputs(3937) <= a;
    layer2_outputs(3938) <= not b or a;
    layer2_outputs(3939) <= a and not b;
    layer2_outputs(3940) <= not b;
    layer2_outputs(3941) <= not a or b;
    layer2_outputs(3942) <= not b;
    layer2_outputs(3943) <= not a;
    layer2_outputs(3944) <= not b;
    layer2_outputs(3945) <= a xor b;
    layer2_outputs(3946) <= a or b;
    layer2_outputs(3947) <= b;
    layer2_outputs(3948) <= a;
    layer2_outputs(3949) <= not b or a;
    layer2_outputs(3950) <= not a or b;
    layer2_outputs(3951) <= not a;
    layer2_outputs(3952) <= not b;
    layer2_outputs(3953) <= not (a or b);
    layer2_outputs(3954) <= not b;
    layer2_outputs(3955) <= b;
    layer2_outputs(3956) <= not b;
    layer2_outputs(3957) <= a;
    layer2_outputs(3958) <= '1';
    layer2_outputs(3959) <= a and not b;
    layer2_outputs(3960) <= not b or a;
    layer2_outputs(3961) <= not (a or b);
    layer2_outputs(3962) <= not (a xor b);
    layer2_outputs(3963) <= not a or b;
    layer2_outputs(3964) <= a and b;
    layer2_outputs(3965) <= a and not b;
    layer2_outputs(3966) <= a xor b;
    layer2_outputs(3967) <= '1';
    layer2_outputs(3968) <= b;
    layer2_outputs(3969) <= a and b;
    layer2_outputs(3970) <= a;
    layer2_outputs(3971) <= not (a and b);
    layer2_outputs(3972) <= b;
    layer2_outputs(3973) <= not a;
    layer2_outputs(3974) <= b and not a;
    layer2_outputs(3975) <= '1';
    layer2_outputs(3976) <= b;
    layer2_outputs(3977) <= b and not a;
    layer2_outputs(3978) <= b and not a;
    layer2_outputs(3979) <= not a;
    layer2_outputs(3980) <= a;
    layer2_outputs(3981) <= not b or a;
    layer2_outputs(3982) <= b;
    layer2_outputs(3983) <= not a or b;
    layer2_outputs(3984) <= '1';
    layer2_outputs(3985) <= a;
    layer2_outputs(3986) <= a or b;
    layer2_outputs(3987) <= a or b;
    layer2_outputs(3988) <= b and not a;
    layer2_outputs(3989) <= not (a and b);
    layer2_outputs(3990) <= '1';
    layer2_outputs(3991) <= a;
    layer2_outputs(3992) <= not b or a;
    layer2_outputs(3993) <= a and b;
    layer2_outputs(3994) <= not (a or b);
    layer2_outputs(3995) <= a xor b;
    layer2_outputs(3996) <= a and b;
    layer2_outputs(3997) <= b and not a;
    layer2_outputs(3998) <= a or b;
    layer2_outputs(3999) <= a and not b;
    layer2_outputs(4000) <= b;
    layer2_outputs(4001) <= a or b;
    layer2_outputs(4002) <= a;
    layer2_outputs(4003) <= not (a and b);
    layer2_outputs(4004) <= '0';
    layer2_outputs(4005) <= not b;
    layer2_outputs(4006) <= b;
    layer2_outputs(4007) <= not (a xor b);
    layer2_outputs(4008) <= a and b;
    layer2_outputs(4009) <= a xor b;
    layer2_outputs(4010) <= not b or a;
    layer2_outputs(4011) <= a or b;
    layer2_outputs(4012) <= a and b;
    layer2_outputs(4013) <= a;
    layer2_outputs(4014) <= a;
    layer2_outputs(4015) <= not b;
    layer2_outputs(4016) <= not (a and b);
    layer2_outputs(4017) <= a and b;
    layer2_outputs(4018) <= a;
    layer2_outputs(4019) <= not a;
    layer2_outputs(4020) <= not b;
    layer2_outputs(4021) <= a and b;
    layer2_outputs(4022) <= '0';
    layer2_outputs(4023) <= b;
    layer2_outputs(4024) <= a;
    layer2_outputs(4025) <= a;
    layer2_outputs(4026) <= not (a or b);
    layer2_outputs(4027) <= a and not b;
    layer2_outputs(4028) <= a and not b;
    layer2_outputs(4029) <= a;
    layer2_outputs(4030) <= '1';
    layer2_outputs(4031) <= b;
    layer2_outputs(4032) <= not b;
    layer2_outputs(4033) <= b;
    layer2_outputs(4034) <= '0';
    layer2_outputs(4035) <= a xor b;
    layer2_outputs(4036) <= a;
    layer2_outputs(4037) <= a xor b;
    layer2_outputs(4038) <= a or b;
    layer2_outputs(4039) <= not a or b;
    layer2_outputs(4040) <= not (a and b);
    layer2_outputs(4041) <= not b;
    layer2_outputs(4042) <= a;
    layer2_outputs(4043) <= a;
    layer2_outputs(4044) <= a and b;
    layer2_outputs(4045) <= not a or b;
    layer2_outputs(4046) <= b;
    layer2_outputs(4047) <= b;
    layer2_outputs(4048) <= not b;
    layer2_outputs(4049) <= not (a xor b);
    layer2_outputs(4050) <= not b or a;
    layer2_outputs(4051) <= a and not b;
    layer2_outputs(4052) <= not b;
    layer2_outputs(4053) <= a or b;
    layer2_outputs(4054) <= a and b;
    layer2_outputs(4055) <= not (a or b);
    layer2_outputs(4056) <= not b;
    layer2_outputs(4057) <= not a;
    layer2_outputs(4058) <= not a;
    layer2_outputs(4059) <= a and not b;
    layer2_outputs(4060) <= b;
    layer2_outputs(4061) <= not (a xor b);
    layer2_outputs(4062) <= not (a xor b);
    layer2_outputs(4063) <= '1';
    layer2_outputs(4064) <= a xor b;
    layer2_outputs(4065) <= not b;
    layer2_outputs(4066) <= not (a or b);
    layer2_outputs(4067) <= a;
    layer2_outputs(4068) <= b;
    layer2_outputs(4069) <= a xor b;
    layer2_outputs(4070) <= a;
    layer2_outputs(4071) <= not a or b;
    layer2_outputs(4072) <= not a;
    layer2_outputs(4073) <= not a;
    layer2_outputs(4074) <= b and not a;
    layer2_outputs(4075) <= not b or a;
    layer2_outputs(4076) <= '1';
    layer2_outputs(4077) <= a or b;
    layer2_outputs(4078) <= not a or b;
    layer2_outputs(4079) <= a and not b;
    layer2_outputs(4080) <= not b;
    layer2_outputs(4081) <= a;
    layer2_outputs(4082) <= not (a and b);
    layer2_outputs(4083) <= '1';
    layer2_outputs(4084) <= a or b;
    layer2_outputs(4085) <= a;
    layer2_outputs(4086) <= not b or a;
    layer2_outputs(4087) <= not a or b;
    layer2_outputs(4088) <= b;
    layer2_outputs(4089) <= not a;
    layer2_outputs(4090) <= b and not a;
    layer2_outputs(4091) <= not b or a;
    layer2_outputs(4092) <= a or b;
    layer2_outputs(4093) <= a;
    layer2_outputs(4094) <= not (a xor b);
    layer2_outputs(4095) <= a and b;
    layer2_outputs(4096) <= b;
    layer2_outputs(4097) <= not b or a;
    layer2_outputs(4098) <= a or b;
    layer2_outputs(4099) <= a;
    layer2_outputs(4100) <= not a or b;
    layer2_outputs(4101) <= b;
    layer2_outputs(4102) <= not (a or b);
    layer2_outputs(4103) <= not (a or b);
    layer2_outputs(4104) <= not (a and b);
    layer2_outputs(4105) <= a;
    layer2_outputs(4106) <= not b;
    layer2_outputs(4107) <= b;
    layer2_outputs(4108) <= a;
    layer2_outputs(4109) <= not a or b;
    layer2_outputs(4110) <= b;
    layer2_outputs(4111) <= not b;
    layer2_outputs(4112) <= not (a xor b);
    layer2_outputs(4113) <= a and not b;
    layer2_outputs(4114) <= not (a xor b);
    layer2_outputs(4115) <= not a;
    layer2_outputs(4116) <= a;
    layer2_outputs(4117) <= a and not b;
    layer2_outputs(4118) <= b;
    layer2_outputs(4119) <= not (a or b);
    layer2_outputs(4120) <= not b;
    layer2_outputs(4121) <= not a;
    layer2_outputs(4122) <= '1';
    layer2_outputs(4123) <= not a or b;
    layer2_outputs(4124) <= b;
    layer2_outputs(4125) <= not (a and b);
    layer2_outputs(4126) <= not a;
    layer2_outputs(4127) <= a and not b;
    layer2_outputs(4128) <= not (a and b);
    layer2_outputs(4129) <= a and not b;
    layer2_outputs(4130) <= b;
    layer2_outputs(4131) <= not b;
    layer2_outputs(4132) <= a and not b;
    layer2_outputs(4133) <= not b;
    layer2_outputs(4134) <= not a;
    layer2_outputs(4135) <= not a or b;
    layer2_outputs(4136) <= a and not b;
    layer2_outputs(4137) <= a and b;
    layer2_outputs(4138) <= not (a xor b);
    layer2_outputs(4139) <= a or b;
    layer2_outputs(4140) <= not a;
    layer2_outputs(4141) <= '1';
    layer2_outputs(4142) <= not b;
    layer2_outputs(4143) <= a;
    layer2_outputs(4144) <= b;
    layer2_outputs(4145) <= a;
    layer2_outputs(4146) <= b;
    layer2_outputs(4147) <= not (a or b);
    layer2_outputs(4148) <= b;
    layer2_outputs(4149) <= a;
    layer2_outputs(4150) <= a and b;
    layer2_outputs(4151) <= not (a xor b);
    layer2_outputs(4152) <= b;
    layer2_outputs(4153) <= not (a or b);
    layer2_outputs(4154) <= not b;
    layer2_outputs(4155) <= a and b;
    layer2_outputs(4156) <= a;
    layer2_outputs(4157) <= not a;
    layer2_outputs(4158) <= a and not b;
    layer2_outputs(4159) <= a and b;
    layer2_outputs(4160) <= b;
    layer2_outputs(4161) <= b and not a;
    layer2_outputs(4162) <= not (a or b);
    layer2_outputs(4163) <= a and b;
    layer2_outputs(4164) <= a;
    layer2_outputs(4165) <= not b or a;
    layer2_outputs(4166) <= a and not b;
    layer2_outputs(4167) <= b;
    layer2_outputs(4168) <= a xor b;
    layer2_outputs(4169) <= '1';
    layer2_outputs(4170) <= not (a and b);
    layer2_outputs(4171) <= '1';
    layer2_outputs(4172) <= a or b;
    layer2_outputs(4173) <= '0';
    layer2_outputs(4174) <= not a or b;
    layer2_outputs(4175) <= not (a and b);
    layer2_outputs(4176) <= not (a and b);
    layer2_outputs(4177) <= not (a xor b);
    layer2_outputs(4178) <= not (a and b);
    layer2_outputs(4179) <= b;
    layer2_outputs(4180) <= not b;
    layer2_outputs(4181) <= b;
    layer2_outputs(4182) <= not a or b;
    layer2_outputs(4183) <= b and not a;
    layer2_outputs(4184) <= not a;
    layer2_outputs(4185) <= b and not a;
    layer2_outputs(4186) <= b;
    layer2_outputs(4187) <= b;
    layer2_outputs(4188) <= not (a xor b);
    layer2_outputs(4189) <= '1';
    layer2_outputs(4190) <= not b;
    layer2_outputs(4191) <= not a or b;
    layer2_outputs(4192) <= a and not b;
    layer2_outputs(4193) <= not (a or b);
    layer2_outputs(4194) <= b and not a;
    layer2_outputs(4195) <= not b or a;
    layer2_outputs(4196) <= a and not b;
    layer2_outputs(4197) <= a;
    layer2_outputs(4198) <= not a or b;
    layer2_outputs(4199) <= a;
    layer2_outputs(4200) <= not (a and b);
    layer2_outputs(4201) <= a xor b;
    layer2_outputs(4202) <= not (a or b);
    layer2_outputs(4203) <= not b or a;
    layer2_outputs(4204) <= not a;
    layer2_outputs(4205) <= a and b;
    layer2_outputs(4206) <= not a;
    layer2_outputs(4207) <= b and not a;
    layer2_outputs(4208) <= not a;
    layer2_outputs(4209) <= not (a xor b);
    layer2_outputs(4210) <= not (a or b);
    layer2_outputs(4211) <= '1';
    layer2_outputs(4212) <= not a or b;
    layer2_outputs(4213) <= a or b;
    layer2_outputs(4214) <= b and not a;
    layer2_outputs(4215) <= a xor b;
    layer2_outputs(4216) <= not a;
    layer2_outputs(4217) <= not a or b;
    layer2_outputs(4218) <= '0';
    layer2_outputs(4219) <= not b;
    layer2_outputs(4220) <= a and not b;
    layer2_outputs(4221) <= not (a or b);
    layer2_outputs(4222) <= a and not b;
    layer2_outputs(4223) <= not a;
    layer2_outputs(4224) <= '1';
    layer2_outputs(4225) <= not b;
    layer2_outputs(4226) <= not b or a;
    layer2_outputs(4227) <= not b;
    layer2_outputs(4228) <= b;
    layer2_outputs(4229) <= b;
    layer2_outputs(4230) <= a and b;
    layer2_outputs(4231) <= b and not a;
    layer2_outputs(4232) <= a;
    layer2_outputs(4233) <= not b;
    layer2_outputs(4234) <= a and b;
    layer2_outputs(4235) <= '0';
    layer2_outputs(4236) <= not (a xor b);
    layer2_outputs(4237) <= not (a xor b);
    layer2_outputs(4238) <= not (a and b);
    layer2_outputs(4239) <= not (a xor b);
    layer2_outputs(4240) <= not b or a;
    layer2_outputs(4241) <= not b or a;
    layer2_outputs(4242) <= not b;
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= a or b;
    layer2_outputs(4245) <= not b;
    layer2_outputs(4246) <= a;
    layer2_outputs(4247) <= not a;
    layer2_outputs(4248) <= b;
    layer2_outputs(4249) <= b;
    layer2_outputs(4250) <= a and b;
    layer2_outputs(4251) <= a;
    layer2_outputs(4252) <= not b or a;
    layer2_outputs(4253) <= not a;
    layer2_outputs(4254) <= not b or a;
    layer2_outputs(4255) <= b and not a;
    layer2_outputs(4256) <= a;
    layer2_outputs(4257) <= not (a and b);
    layer2_outputs(4258) <= a;
    layer2_outputs(4259) <= not a;
    layer2_outputs(4260) <= b and not a;
    layer2_outputs(4261) <= not (a and b);
    layer2_outputs(4262) <= not (a or b);
    layer2_outputs(4263) <= a and b;
    layer2_outputs(4264) <= b and not a;
    layer2_outputs(4265) <= a and not b;
    layer2_outputs(4266) <= not (a or b);
    layer2_outputs(4267) <= b;
    layer2_outputs(4268) <= not (a or b);
    layer2_outputs(4269) <= b and not a;
    layer2_outputs(4270) <= b;
    layer2_outputs(4271) <= a and b;
    layer2_outputs(4272) <= '1';
    layer2_outputs(4273) <= '1';
    layer2_outputs(4274) <= not b;
    layer2_outputs(4275) <= not b or a;
    layer2_outputs(4276) <= b;
    layer2_outputs(4277) <= a or b;
    layer2_outputs(4278) <= not b;
    layer2_outputs(4279) <= not a;
    layer2_outputs(4280) <= not (a or b);
    layer2_outputs(4281) <= not b;
    layer2_outputs(4282) <= a;
    layer2_outputs(4283) <= not (a and b);
    layer2_outputs(4284) <= a or b;
    layer2_outputs(4285) <= a;
    layer2_outputs(4286) <= '0';
    layer2_outputs(4287) <= not b;
    layer2_outputs(4288) <= b and not a;
    layer2_outputs(4289) <= not (a xor b);
    layer2_outputs(4290) <= a and not b;
    layer2_outputs(4291) <= not (a or b);
    layer2_outputs(4292) <= b and not a;
    layer2_outputs(4293) <= not b or a;
    layer2_outputs(4294) <= not a;
    layer2_outputs(4295) <= not a or b;
    layer2_outputs(4296) <= not (a or b);
    layer2_outputs(4297) <= a;
    layer2_outputs(4298) <= not a;
    layer2_outputs(4299) <= b and not a;
    layer2_outputs(4300) <= a and b;
    layer2_outputs(4301) <= '1';
    layer2_outputs(4302) <= not a or b;
    layer2_outputs(4303) <= not b;
    layer2_outputs(4304) <= b and not a;
    layer2_outputs(4305) <= b;
    layer2_outputs(4306) <= a and b;
    layer2_outputs(4307) <= not b;
    layer2_outputs(4308) <= not (a and b);
    layer2_outputs(4309) <= not b;
    layer2_outputs(4310) <= not (a or b);
    layer2_outputs(4311) <= b;
    layer2_outputs(4312) <= not a or b;
    layer2_outputs(4313) <= a or b;
    layer2_outputs(4314) <= not b;
    layer2_outputs(4315) <= not b;
    layer2_outputs(4316) <= not (a and b);
    layer2_outputs(4317) <= a;
    layer2_outputs(4318) <= a or b;
    layer2_outputs(4319) <= not b or a;
    layer2_outputs(4320) <= not a or b;
    layer2_outputs(4321) <= not a;
    layer2_outputs(4322) <= a and b;
    layer2_outputs(4323) <= '0';
    layer2_outputs(4324) <= not a or b;
    layer2_outputs(4325) <= not a or b;
    layer2_outputs(4326) <= not a;
    layer2_outputs(4327) <= not (a xor b);
    layer2_outputs(4328) <= b;
    layer2_outputs(4329) <= b;
    layer2_outputs(4330) <= '1';
    layer2_outputs(4331) <= not (a xor b);
    layer2_outputs(4332) <= not b or a;
    layer2_outputs(4333) <= not b;
    layer2_outputs(4334) <= b and not a;
    layer2_outputs(4335) <= a xor b;
    layer2_outputs(4336) <= a;
    layer2_outputs(4337) <= a xor b;
    layer2_outputs(4338) <= not b;
    layer2_outputs(4339) <= not b or a;
    layer2_outputs(4340) <= not b;
    layer2_outputs(4341) <= not b;
    layer2_outputs(4342) <= not a;
    layer2_outputs(4343) <= '0';
    layer2_outputs(4344) <= a and not b;
    layer2_outputs(4345) <= a or b;
    layer2_outputs(4346) <= not (a or b);
    layer2_outputs(4347) <= not a or b;
    layer2_outputs(4348) <= a and not b;
    layer2_outputs(4349) <= a;
    layer2_outputs(4350) <= not a;
    layer2_outputs(4351) <= a xor b;
    layer2_outputs(4352) <= b and not a;
    layer2_outputs(4353) <= a;
    layer2_outputs(4354) <= b;
    layer2_outputs(4355) <= a;
    layer2_outputs(4356) <= not b;
    layer2_outputs(4357) <= not b;
    layer2_outputs(4358) <= not a;
    layer2_outputs(4359) <= not (a or b);
    layer2_outputs(4360) <= '0';
    layer2_outputs(4361) <= not (a xor b);
    layer2_outputs(4362) <= a and b;
    layer2_outputs(4363) <= a and not b;
    layer2_outputs(4364) <= not (a or b);
    layer2_outputs(4365) <= not (a or b);
    layer2_outputs(4366) <= b and not a;
    layer2_outputs(4367) <= a and not b;
    layer2_outputs(4368) <= not a;
    layer2_outputs(4369) <= b;
    layer2_outputs(4370) <= not a;
    layer2_outputs(4371) <= a;
    layer2_outputs(4372) <= not a or b;
    layer2_outputs(4373) <= not b or a;
    layer2_outputs(4374) <= not b;
    layer2_outputs(4375) <= not b;
    layer2_outputs(4376) <= not b or a;
    layer2_outputs(4377) <= b;
    layer2_outputs(4378) <= not b;
    layer2_outputs(4379) <= a or b;
    layer2_outputs(4380) <= not a or b;
    layer2_outputs(4381) <= '0';
    layer2_outputs(4382) <= not b or a;
    layer2_outputs(4383) <= not a or b;
    layer2_outputs(4384) <= b and not a;
    layer2_outputs(4385) <= not b;
    layer2_outputs(4386) <= not b;
    layer2_outputs(4387) <= not (a or b);
    layer2_outputs(4388) <= b;
    layer2_outputs(4389) <= not (a or b);
    layer2_outputs(4390) <= a;
    layer2_outputs(4391) <= not b;
    layer2_outputs(4392) <= not a;
    layer2_outputs(4393) <= a;
    layer2_outputs(4394) <= not (a or b);
    layer2_outputs(4395) <= a and b;
    layer2_outputs(4396) <= not b;
    layer2_outputs(4397) <= not (a or b);
    layer2_outputs(4398) <= a and b;
    layer2_outputs(4399) <= a and not b;
    layer2_outputs(4400) <= b;
    layer2_outputs(4401) <= a and not b;
    layer2_outputs(4402) <= '0';
    layer2_outputs(4403) <= b and not a;
    layer2_outputs(4404) <= not a;
    layer2_outputs(4405) <= not b;
    layer2_outputs(4406) <= b and not a;
    layer2_outputs(4407) <= a xor b;
    layer2_outputs(4408) <= b;
    layer2_outputs(4409) <= not b or a;
    layer2_outputs(4410) <= not a;
    layer2_outputs(4411) <= a and b;
    layer2_outputs(4412) <= not (a xor b);
    layer2_outputs(4413) <= a;
    layer2_outputs(4414) <= a and not b;
    layer2_outputs(4415) <= not (a or b);
    layer2_outputs(4416) <= not (a and b);
    layer2_outputs(4417) <= not (a and b);
    layer2_outputs(4418) <= b;
    layer2_outputs(4419) <= a or b;
    layer2_outputs(4420) <= '0';
    layer2_outputs(4421) <= not (a or b);
    layer2_outputs(4422) <= not b or a;
    layer2_outputs(4423) <= a;
    layer2_outputs(4424) <= not b;
    layer2_outputs(4425) <= not a or b;
    layer2_outputs(4426) <= a or b;
    layer2_outputs(4427) <= not a or b;
    layer2_outputs(4428) <= b;
    layer2_outputs(4429) <= b and not a;
    layer2_outputs(4430) <= not a;
    layer2_outputs(4431) <= not a;
    layer2_outputs(4432) <= not (a and b);
    layer2_outputs(4433) <= a or b;
    layer2_outputs(4434) <= a;
    layer2_outputs(4435) <= not (a or b);
    layer2_outputs(4436) <= b and not a;
    layer2_outputs(4437) <= a and b;
    layer2_outputs(4438) <= b;
    layer2_outputs(4439) <= b;
    layer2_outputs(4440) <= not b;
    layer2_outputs(4441) <= not a or b;
    layer2_outputs(4442) <= a;
    layer2_outputs(4443) <= not (a and b);
    layer2_outputs(4444) <= not b or a;
    layer2_outputs(4445) <= a xor b;
    layer2_outputs(4446) <= a or b;
    layer2_outputs(4447) <= not a or b;
    layer2_outputs(4448) <= a or b;
    layer2_outputs(4449) <= a;
    layer2_outputs(4450) <= b and not a;
    layer2_outputs(4451) <= not (a xor b);
    layer2_outputs(4452) <= b and not a;
    layer2_outputs(4453) <= a xor b;
    layer2_outputs(4454) <= a and b;
    layer2_outputs(4455) <= not (a or b);
    layer2_outputs(4456) <= not a or b;
    layer2_outputs(4457) <= a or b;
    layer2_outputs(4458) <= not b;
    layer2_outputs(4459) <= not (a or b);
    layer2_outputs(4460) <= b;
    layer2_outputs(4461) <= b and not a;
    layer2_outputs(4462) <= not b or a;
    layer2_outputs(4463) <= a and b;
    layer2_outputs(4464) <= not (a and b);
    layer2_outputs(4465) <= not b;
    layer2_outputs(4466) <= b;
    layer2_outputs(4467) <= b and not a;
    layer2_outputs(4468) <= '0';
    layer2_outputs(4469) <= not a or b;
    layer2_outputs(4470) <= a;
    layer2_outputs(4471) <= not b;
    layer2_outputs(4472) <= b;
    layer2_outputs(4473) <= not (a or b);
    layer2_outputs(4474) <= not a;
    layer2_outputs(4475) <= a or b;
    layer2_outputs(4476) <= a and not b;
    layer2_outputs(4477) <= not a;
    layer2_outputs(4478) <= a;
    layer2_outputs(4479) <= a;
    layer2_outputs(4480) <= a and not b;
    layer2_outputs(4481) <= b;
    layer2_outputs(4482) <= not (a xor b);
    layer2_outputs(4483) <= not (a or b);
    layer2_outputs(4484) <= not (a or b);
    layer2_outputs(4485) <= a and b;
    layer2_outputs(4486) <= b;
    layer2_outputs(4487) <= not b;
    layer2_outputs(4488) <= not b or a;
    layer2_outputs(4489) <= not a or b;
    layer2_outputs(4490) <= not b or a;
    layer2_outputs(4491) <= not b;
    layer2_outputs(4492) <= not a;
    layer2_outputs(4493) <= not a;
    layer2_outputs(4494) <= a;
    layer2_outputs(4495) <= '1';
    layer2_outputs(4496) <= a xor b;
    layer2_outputs(4497) <= not a or b;
    layer2_outputs(4498) <= not (a and b);
    layer2_outputs(4499) <= not b;
    layer2_outputs(4500) <= a;
    layer2_outputs(4501) <= b and not a;
    layer2_outputs(4502) <= not b;
    layer2_outputs(4503) <= not b or a;
    layer2_outputs(4504) <= not b;
    layer2_outputs(4505) <= not b or a;
    layer2_outputs(4506) <= a and b;
    layer2_outputs(4507) <= not (a xor b);
    layer2_outputs(4508) <= '1';
    layer2_outputs(4509) <= not a or b;
    layer2_outputs(4510) <= a or b;
    layer2_outputs(4511) <= a and b;
    layer2_outputs(4512) <= not b or a;
    layer2_outputs(4513) <= b;
    layer2_outputs(4514) <= not b;
    layer2_outputs(4515) <= a and not b;
    layer2_outputs(4516) <= b;
    layer2_outputs(4517) <= a or b;
    layer2_outputs(4518) <= not a;
    layer2_outputs(4519) <= not a or b;
    layer2_outputs(4520) <= not a or b;
    layer2_outputs(4521) <= a;
    layer2_outputs(4522) <= not b;
    layer2_outputs(4523) <= not b;
    layer2_outputs(4524) <= not a;
    layer2_outputs(4525) <= not b or a;
    layer2_outputs(4526) <= not b;
    layer2_outputs(4527) <= a and not b;
    layer2_outputs(4528) <= not b or a;
    layer2_outputs(4529) <= '0';
    layer2_outputs(4530) <= not a or b;
    layer2_outputs(4531) <= not b or a;
    layer2_outputs(4532) <= b;
    layer2_outputs(4533) <= not a;
    layer2_outputs(4534) <= b;
    layer2_outputs(4535) <= a;
    layer2_outputs(4536) <= a and not b;
    layer2_outputs(4537) <= not b or a;
    layer2_outputs(4538) <= not (a or b);
    layer2_outputs(4539) <= not a or b;
    layer2_outputs(4540) <= not a;
    layer2_outputs(4541) <= a and not b;
    layer2_outputs(4542) <= a and not b;
    layer2_outputs(4543) <= not (a xor b);
    layer2_outputs(4544) <= not (a or b);
    layer2_outputs(4545) <= not a or b;
    layer2_outputs(4546) <= not a or b;
    layer2_outputs(4547) <= a;
    layer2_outputs(4548) <= not (a and b);
    layer2_outputs(4549) <= a;
    layer2_outputs(4550) <= not (a or b);
    layer2_outputs(4551) <= not (a or b);
    layer2_outputs(4552) <= not (a or b);
    layer2_outputs(4553) <= not a;
    layer2_outputs(4554) <= b;
    layer2_outputs(4555) <= '1';
    layer2_outputs(4556) <= a;
    layer2_outputs(4557) <= '0';
    layer2_outputs(4558) <= not (a xor b);
    layer2_outputs(4559) <= not (a and b);
    layer2_outputs(4560) <= not (a and b);
    layer2_outputs(4561) <= b and not a;
    layer2_outputs(4562) <= not b;
    layer2_outputs(4563) <= a;
    layer2_outputs(4564) <= not b or a;
    layer2_outputs(4565) <= b;
    layer2_outputs(4566) <= not a or b;
    layer2_outputs(4567) <= b;
    layer2_outputs(4568) <= not a;
    layer2_outputs(4569) <= not a;
    layer2_outputs(4570) <= a;
    layer2_outputs(4571) <= not (a and b);
    layer2_outputs(4572) <= a xor b;
    layer2_outputs(4573) <= a;
    layer2_outputs(4574) <= not a or b;
    layer2_outputs(4575) <= '1';
    layer2_outputs(4576) <= '1';
    layer2_outputs(4577) <= a and not b;
    layer2_outputs(4578) <= b;
    layer2_outputs(4579) <= not a or b;
    layer2_outputs(4580) <= not (a and b);
    layer2_outputs(4581) <= not b;
    layer2_outputs(4582) <= not (a or b);
    layer2_outputs(4583) <= b;
    layer2_outputs(4584) <= not a;
    layer2_outputs(4585) <= b and not a;
    layer2_outputs(4586) <= '1';
    layer2_outputs(4587) <= a and b;
    layer2_outputs(4588) <= not b or a;
    layer2_outputs(4589) <= not (a or b);
    layer2_outputs(4590) <= not a;
    layer2_outputs(4591) <= '0';
    layer2_outputs(4592) <= b;
    layer2_outputs(4593) <= not (a xor b);
    layer2_outputs(4594) <= b;
    layer2_outputs(4595) <= '1';
    layer2_outputs(4596) <= a;
    layer2_outputs(4597) <= a;
    layer2_outputs(4598) <= not (a or b);
    layer2_outputs(4599) <= b and not a;
    layer2_outputs(4600) <= '1';
    layer2_outputs(4601) <= a and not b;
    layer2_outputs(4602) <= not b;
    layer2_outputs(4603) <= not (a and b);
    layer2_outputs(4604) <= a and b;
    layer2_outputs(4605) <= not (a and b);
    layer2_outputs(4606) <= a xor b;
    layer2_outputs(4607) <= not a;
    layer2_outputs(4608) <= a;
    layer2_outputs(4609) <= b;
    layer2_outputs(4610) <= '1';
    layer2_outputs(4611) <= not b;
    layer2_outputs(4612) <= a or b;
    layer2_outputs(4613) <= b;
    layer2_outputs(4614) <= a and not b;
    layer2_outputs(4615) <= b and not a;
    layer2_outputs(4616) <= '1';
    layer2_outputs(4617) <= a or b;
    layer2_outputs(4618) <= not a or b;
    layer2_outputs(4619) <= not b;
    layer2_outputs(4620) <= b;
    layer2_outputs(4621) <= a;
    layer2_outputs(4622) <= a xor b;
    layer2_outputs(4623) <= not b or a;
    layer2_outputs(4624) <= not (a and b);
    layer2_outputs(4625) <= not (a or b);
    layer2_outputs(4626) <= b and not a;
    layer2_outputs(4627) <= not a or b;
    layer2_outputs(4628) <= not b or a;
    layer2_outputs(4629) <= not a;
    layer2_outputs(4630) <= not a or b;
    layer2_outputs(4631) <= a and b;
    layer2_outputs(4632) <= a;
    layer2_outputs(4633) <= not b;
    layer2_outputs(4634) <= '1';
    layer2_outputs(4635) <= a;
    layer2_outputs(4636) <= a xor b;
    layer2_outputs(4637) <= not a;
    layer2_outputs(4638) <= a xor b;
    layer2_outputs(4639) <= b and not a;
    layer2_outputs(4640) <= '1';
    layer2_outputs(4641) <= b;
    layer2_outputs(4642) <= a xor b;
    layer2_outputs(4643) <= '0';
    layer2_outputs(4644) <= not (a and b);
    layer2_outputs(4645) <= not b;
    layer2_outputs(4646) <= a and not b;
    layer2_outputs(4647) <= not (a or b);
    layer2_outputs(4648) <= not b or a;
    layer2_outputs(4649) <= b and not a;
    layer2_outputs(4650) <= not a;
    layer2_outputs(4651) <= not b;
    layer2_outputs(4652) <= a or b;
    layer2_outputs(4653) <= not (a or b);
    layer2_outputs(4654) <= not a;
    layer2_outputs(4655) <= not b or a;
    layer2_outputs(4656) <= a or b;
    layer2_outputs(4657) <= not b;
    layer2_outputs(4658) <= not a;
    layer2_outputs(4659) <= b;
    layer2_outputs(4660) <= not (a or b);
    layer2_outputs(4661) <= not a;
    layer2_outputs(4662) <= a;
    layer2_outputs(4663) <= not (a xor b);
    layer2_outputs(4664) <= not (a and b);
    layer2_outputs(4665) <= a;
    layer2_outputs(4666) <= not a or b;
    layer2_outputs(4667) <= not a;
    layer2_outputs(4668) <= b and not a;
    layer2_outputs(4669) <= not b or a;
    layer2_outputs(4670) <= '1';
    layer2_outputs(4671) <= not b;
    layer2_outputs(4672) <= b;
    layer2_outputs(4673) <= b and not a;
    layer2_outputs(4674) <= a;
    layer2_outputs(4675) <= not b;
    layer2_outputs(4676) <= not (a and b);
    layer2_outputs(4677) <= not b;
    layer2_outputs(4678) <= not a;
    layer2_outputs(4679) <= not b or a;
    layer2_outputs(4680) <= '0';
    layer2_outputs(4681) <= not b;
    layer2_outputs(4682) <= b and not a;
    layer2_outputs(4683) <= '1';
    layer2_outputs(4684) <= not a;
    layer2_outputs(4685) <= a and b;
    layer2_outputs(4686) <= a or b;
    layer2_outputs(4687) <= not a or b;
    layer2_outputs(4688) <= a and not b;
    layer2_outputs(4689) <= not (a xor b);
    layer2_outputs(4690) <= not (a xor b);
    layer2_outputs(4691) <= b and not a;
    layer2_outputs(4692) <= b;
    layer2_outputs(4693) <= not b;
    layer2_outputs(4694) <= not (a xor b);
    layer2_outputs(4695) <= not b;
    layer2_outputs(4696) <= not b;
    layer2_outputs(4697) <= not (a or b);
    layer2_outputs(4698) <= b;
    layer2_outputs(4699) <= a;
    layer2_outputs(4700) <= a;
    layer2_outputs(4701) <= not (a xor b);
    layer2_outputs(4702) <= a or b;
    layer2_outputs(4703) <= not (a or b);
    layer2_outputs(4704) <= not (a and b);
    layer2_outputs(4705) <= not (a or b);
    layer2_outputs(4706) <= a xor b;
    layer2_outputs(4707) <= a;
    layer2_outputs(4708) <= b;
    layer2_outputs(4709) <= not b or a;
    layer2_outputs(4710) <= not (a xor b);
    layer2_outputs(4711) <= b and not a;
    layer2_outputs(4712) <= b;
    layer2_outputs(4713) <= a or b;
    layer2_outputs(4714) <= not a or b;
    layer2_outputs(4715) <= not b;
    layer2_outputs(4716) <= not b;
    layer2_outputs(4717) <= not a;
    layer2_outputs(4718) <= not (a or b);
    layer2_outputs(4719) <= not a;
    layer2_outputs(4720) <= a and not b;
    layer2_outputs(4721) <= not a;
    layer2_outputs(4722) <= a xor b;
    layer2_outputs(4723) <= not b;
    layer2_outputs(4724) <= not (a or b);
    layer2_outputs(4725) <= not (a or b);
    layer2_outputs(4726) <= b;
    layer2_outputs(4727) <= a xor b;
    layer2_outputs(4728) <= a;
    layer2_outputs(4729) <= b;
    layer2_outputs(4730) <= not (a or b);
    layer2_outputs(4731) <= not a;
    layer2_outputs(4732) <= not b;
    layer2_outputs(4733) <= not a;
    layer2_outputs(4734) <= b and not a;
    layer2_outputs(4735) <= not b or a;
    layer2_outputs(4736) <= not (a and b);
    layer2_outputs(4737) <= b;
    layer2_outputs(4738) <= a;
    layer2_outputs(4739) <= not (a xor b);
    layer2_outputs(4740) <= not b or a;
    layer2_outputs(4741) <= a or b;
    layer2_outputs(4742) <= not (a or b);
    layer2_outputs(4743) <= not (a and b);
    layer2_outputs(4744) <= not a or b;
    layer2_outputs(4745) <= b;
    layer2_outputs(4746) <= not (a or b);
    layer2_outputs(4747) <= not (a xor b);
    layer2_outputs(4748) <= not a;
    layer2_outputs(4749) <= not a or b;
    layer2_outputs(4750) <= not a or b;
    layer2_outputs(4751) <= a or b;
    layer2_outputs(4752) <= not (a or b);
    layer2_outputs(4753) <= not a;
    layer2_outputs(4754) <= b;
    layer2_outputs(4755) <= not a;
    layer2_outputs(4756) <= not b;
    layer2_outputs(4757) <= not (a and b);
    layer2_outputs(4758) <= '1';
    layer2_outputs(4759) <= not a or b;
    layer2_outputs(4760) <= not a or b;
    layer2_outputs(4761) <= '1';
    layer2_outputs(4762) <= not (a and b);
    layer2_outputs(4763) <= a;
    layer2_outputs(4764) <= not b;
    layer2_outputs(4765) <= a and b;
    layer2_outputs(4766) <= not a;
    layer2_outputs(4767) <= a and not b;
    layer2_outputs(4768) <= '1';
    layer2_outputs(4769) <= not (a xor b);
    layer2_outputs(4770) <= a;
    layer2_outputs(4771) <= not b or a;
    layer2_outputs(4772) <= not b;
    layer2_outputs(4773) <= '1';
    layer2_outputs(4774) <= not a or b;
    layer2_outputs(4775) <= a and not b;
    layer2_outputs(4776) <= a;
    layer2_outputs(4777) <= not b;
    layer2_outputs(4778) <= '0';
    layer2_outputs(4779) <= a and not b;
    layer2_outputs(4780) <= not (a or b);
    layer2_outputs(4781) <= not b;
    layer2_outputs(4782) <= not (a xor b);
    layer2_outputs(4783) <= not a;
    layer2_outputs(4784) <= '1';
    layer2_outputs(4785) <= a;
    layer2_outputs(4786) <= not b or a;
    layer2_outputs(4787) <= not b;
    layer2_outputs(4788) <= b and not a;
    layer2_outputs(4789) <= not (a or b);
    layer2_outputs(4790) <= not a;
    layer2_outputs(4791) <= '0';
    layer2_outputs(4792) <= b;
    layer2_outputs(4793) <= not (a or b);
    layer2_outputs(4794) <= a or b;
    layer2_outputs(4795) <= a;
    layer2_outputs(4796) <= '1';
    layer2_outputs(4797) <= not (a xor b);
    layer2_outputs(4798) <= a and not b;
    layer2_outputs(4799) <= a;
    layer2_outputs(4800) <= not (a xor b);
    layer2_outputs(4801) <= not (a xor b);
    layer2_outputs(4802) <= b and not a;
    layer2_outputs(4803) <= a and b;
    layer2_outputs(4804) <= b;
    layer2_outputs(4805) <= not b or a;
    layer2_outputs(4806) <= b;
    layer2_outputs(4807) <= not a or b;
    layer2_outputs(4808) <= a or b;
    layer2_outputs(4809) <= not (a or b);
    layer2_outputs(4810) <= not a or b;
    layer2_outputs(4811) <= a;
    layer2_outputs(4812) <= '0';
    layer2_outputs(4813) <= not (a and b);
    layer2_outputs(4814) <= a;
    layer2_outputs(4815) <= not b or a;
    layer2_outputs(4816) <= b;
    layer2_outputs(4817) <= not b;
    layer2_outputs(4818) <= not b;
    layer2_outputs(4819) <= a and b;
    layer2_outputs(4820) <= not a or b;
    layer2_outputs(4821) <= b and not a;
    layer2_outputs(4822) <= a and b;
    layer2_outputs(4823) <= b and not a;
    layer2_outputs(4824) <= a xor b;
    layer2_outputs(4825) <= a and not b;
    layer2_outputs(4826) <= a;
    layer2_outputs(4827) <= a or b;
    layer2_outputs(4828) <= a;
    layer2_outputs(4829) <= not (a xor b);
    layer2_outputs(4830) <= b and not a;
    layer2_outputs(4831) <= not (a or b);
    layer2_outputs(4832) <= a and b;
    layer2_outputs(4833) <= a or b;
    layer2_outputs(4834) <= not b or a;
    layer2_outputs(4835) <= a and not b;
    layer2_outputs(4836) <= not b;
    layer2_outputs(4837) <= not b or a;
    layer2_outputs(4838) <= b;
    layer2_outputs(4839) <= '1';
    layer2_outputs(4840) <= not b or a;
    layer2_outputs(4841) <= a;
    layer2_outputs(4842) <= not a;
    layer2_outputs(4843) <= not a;
    layer2_outputs(4844) <= not b or a;
    layer2_outputs(4845) <= not (a or b);
    layer2_outputs(4846) <= not a or b;
    layer2_outputs(4847) <= a and b;
    layer2_outputs(4848) <= not (a xor b);
    layer2_outputs(4849) <= b;
    layer2_outputs(4850) <= a;
    layer2_outputs(4851) <= not (a or b);
    layer2_outputs(4852) <= not b or a;
    layer2_outputs(4853) <= a and b;
    layer2_outputs(4854) <= not a;
    layer2_outputs(4855) <= not b;
    layer2_outputs(4856) <= a and not b;
    layer2_outputs(4857) <= a and not b;
    layer2_outputs(4858) <= a;
    layer2_outputs(4859) <= not b or a;
    layer2_outputs(4860) <= not (a and b);
    layer2_outputs(4861) <= a and b;
    layer2_outputs(4862) <= a and b;
    layer2_outputs(4863) <= b and not a;
    layer2_outputs(4864) <= not (a or b);
    layer2_outputs(4865) <= a xor b;
    layer2_outputs(4866) <= not a or b;
    layer2_outputs(4867) <= a and b;
    layer2_outputs(4868) <= b;
    layer2_outputs(4869) <= b;
    layer2_outputs(4870) <= not (a xor b);
    layer2_outputs(4871) <= a or b;
    layer2_outputs(4872) <= not a or b;
    layer2_outputs(4873) <= not a;
    layer2_outputs(4874) <= not a;
    layer2_outputs(4875) <= a;
    layer2_outputs(4876) <= b;
    layer2_outputs(4877) <= not b;
    layer2_outputs(4878) <= not b or a;
    layer2_outputs(4879) <= b;
    layer2_outputs(4880) <= a and b;
    layer2_outputs(4881) <= not (a and b);
    layer2_outputs(4882) <= not (a or b);
    layer2_outputs(4883) <= not b;
    layer2_outputs(4884) <= not a or b;
    layer2_outputs(4885) <= not (a and b);
    layer2_outputs(4886) <= a and b;
    layer2_outputs(4887) <= not a;
    layer2_outputs(4888) <= '0';
    layer2_outputs(4889) <= not (a or b);
    layer2_outputs(4890) <= not b or a;
    layer2_outputs(4891) <= b;
    layer2_outputs(4892) <= not (a xor b);
    layer2_outputs(4893) <= a and b;
    layer2_outputs(4894) <= not (a or b);
    layer2_outputs(4895) <= b and not a;
    layer2_outputs(4896) <= b;
    layer2_outputs(4897) <= not b;
    layer2_outputs(4898) <= not (a and b);
    layer2_outputs(4899) <= a;
    layer2_outputs(4900) <= b and not a;
    layer2_outputs(4901) <= not b or a;
    layer2_outputs(4902) <= b;
    layer2_outputs(4903) <= not a or b;
    layer2_outputs(4904) <= not (a and b);
    layer2_outputs(4905) <= a or b;
    layer2_outputs(4906) <= not a or b;
    layer2_outputs(4907) <= not b;
    layer2_outputs(4908) <= not (a or b);
    layer2_outputs(4909) <= a;
    layer2_outputs(4910) <= a and not b;
    layer2_outputs(4911) <= not b;
    layer2_outputs(4912) <= not a;
    layer2_outputs(4913) <= not a or b;
    layer2_outputs(4914) <= b;
    layer2_outputs(4915) <= not (a or b);
    layer2_outputs(4916) <= a xor b;
    layer2_outputs(4917) <= not a or b;
    layer2_outputs(4918) <= a and not b;
    layer2_outputs(4919) <= '0';
    layer2_outputs(4920) <= a and not b;
    layer2_outputs(4921) <= not a;
    layer2_outputs(4922) <= not b;
    layer2_outputs(4923) <= a and not b;
    layer2_outputs(4924) <= b and not a;
    layer2_outputs(4925) <= b and not a;
    layer2_outputs(4926) <= not (a xor b);
    layer2_outputs(4927) <= a or b;
    layer2_outputs(4928) <= '1';
    layer2_outputs(4929) <= not (a and b);
    layer2_outputs(4930) <= not (a and b);
    layer2_outputs(4931) <= not (a or b);
    layer2_outputs(4932) <= a and b;
    layer2_outputs(4933) <= not a;
    layer2_outputs(4934) <= not (a or b);
    layer2_outputs(4935) <= not b;
    layer2_outputs(4936) <= b and not a;
    layer2_outputs(4937) <= a;
    layer2_outputs(4938) <= not (a or b);
    layer2_outputs(4939) <= '0';
    layer2_outputs(4940) <= b;
    layer2_outputs(4941) <= not a;
    layer2_outputs(4942) <= not b or a;
    layer2_outputs(4943) <= not a;
    layer2_outputs(4944) <= a;
    layer2_outputs(4945) <= not a;
    layer2_outputs(4946) <= not a or b;
    layer2_outputs(4947) <= not (a xor b);
    layer2_outputs(4948) <= b;
    layer2_outputs(4949) <= a and not b;
    layer2_outputs(4950) <= not b or a;
    layer2_outputs(4951) <= not a or b;
    layer2_outputs(4952) <= b;
    layer2_outputs(4953) <= a or b;
    layer2_outputs(4954) <= a and not b;
    layer2_outputs(4955) <= a;
    layer2_outputs(4956) <= a and b;
    layer2_outputs(4957) <= a or b;
    layer2_outputs(4958) <= not (a or b);
    layer2_outputs(4959) <= b;
    layer2_outputs(4960) <= a and b;
    layer2_outputs(4961) <= '1';
    layer2_outputs(4962) <= b and not a;
    layer2_outputs(4963) <= a or b;
    layer2_outputs(4964) <= not a or b;
    layer2_outputs(4965) <= b and not a;
    layer2_outputs(4966) <= not a or b;
    layer2_outputs(4967) <= not (a xor b);
    layer2_outputs(4968) <= b;
    layer2_outputs(4969) <= b;
    layer2_outputs(4970) <= a;
    layer2_outputs(4971) <= a;
    layer2_outputs(4972) <= a and not b;
    layer2_outputs(4973) <= a or b;
    layer2_outputs(4974) <= a;
    layer2_outputs(4975) <= not a;
    layer2_outputs(4976) <= not b;
    layer2_outputs(4977) <= not (a and b);
    layer2_outputs(4978) <= not b or a;
    layer2_outputs(4979) <= not (a or b);
    layer2_outputs(4980) <= a and not b;
    layer2_outputs(4981) <= a and not b;
    layer2_outputs(4982) <= not (a or b);
    layer2_outputs(4983) <= not a;
    layer2_outputs(4984) <= a and b;
    layer2_outputs(4985) <= not b;
    layer2_outputs(4986) <= a or b;
    layer2_outputs(4987) <= a xor b;
    layer2_outputs(4988) <= a;
    layer2_outputs(4989) <= b and not a;
    layer2_outputs(4990) <= b and not a;
    layer2_outputs(4991) <= not a;
    layer2_outputs(4992) <= b;
    layer2_outputs(4993) <= a and not b;
    layer2_outputs(4994) <= a or b;
    layer2_outputs(4995) <= not b or a;
    layer2_outputs(4996) <= b and not a;
    layer2_outputs(4997) <= b;
    layer2_outputs(4998) <= b and not a;
    layer2_outputs(4999) <= b and not a;
    layer2_outputs(5000) <= not a or b;
    layer2_outputs(5001) <= not (a and b);
    layer2_outputs(5002) <= not a or b;
    layer2_outputs(5003) <= b;
    layer2_outputs(5004) <= not (a and b);
    layer2_outputs(5005) <= not (a and b);
    layer2_outputs(5006) <= a and b;
    layer2_outputs(5007) <= not (a and b);
    layer2_outputs(5008) <= not (a or b);
    layer2_outputs(5009) <= not b;
    layer2_outputs(5010) <= not a;
    layer2_outputs(5011) <= a xor b;
    layer2_outputs(5012) <= not a;
    layer2_outputs(5013) <= a and not b;
    layer2_outputs(5014) <= not b;
    layer2_outputs(5015) <= b;
    layer2_outputs(5016) <= not b;
    layer2_outputs(5017) <= not a;
    layer2_outputs(5018) <= not a or b;
    layer2_outputs(5019) <= not (a and b);
    layer2_outputs(5020) <= '1';
    layer2_outputs(5021) <= not b;
    layer2_outputs(5022) <= b;
    layer2_outputs(5023) <= not (a and b);
    layer2_outputs(5024) <= a;
    layer2_outputs(5025) <= not (a or b);
    layer2_outputs(5026) <= '1';
    layer2_outputs(5027) <= a and b;
    layer2_outputs(5028) <= a and not b;
    layer2_outputs(5029) <= '0';
    layer2_outputs(5030) <= b;
    layer2_outputs(5031) <= a and b;
    layer2_outputs(5032) <= not (a and b);
    layer2_outputs(5033) <= a;
    layer2_outputs(5034) <= not (a and b);
    layer2_outputs(5035) <= a xor b;
    layer2_outputs(5036) <= b and not a;
    layer2_outputs(5037) <= a;
    layer2_outputs(5038) <= b and not a;
    layer2_outputs(5039) <= a;
    layer2_outputs(5040) <= a or b;
    layer2_outputs(5041) <= not (a or b);
    layer2_outputs(5042) <= a;
    layer2_outputs(5043) <= a xor b;
    layer2_outputs(5044) <= not a;
    layer2_outputs(5045) <= not (a xor b);
    layer2_outputs(5046) <= not (a and b);
    layer2_outputs(5047) <= b;
    layer2_outputs(5048) <= not b;
    layer2_outputs(5049) <= a and not b;
    layer2_outputs(5050) <= not b or a;
    layer2_outputs(5051) <= a and b;
    layer2_outputs(5052) <= a or b;
    layer2_outputs(5053) <= not (a and b);
    layer2_outputs(5054) <= '0';
    layer2_outputs(5055) <= not b;
    layer2_outputs(5056) <= a and b;
    layer2_outputs(5057) <= b and not a;
    layer2_outputs(5058) <= a and not b;
    layer2_outputs(5059) <= not a;
    layer2_outputs(5060) <= a and b;
    layer2_outputs(5061) <= a and not b;
    layer2_outputs(5062) <= not a;
    layer2_outputs(5063) <= a and not b;
    layer2_outputs(5064) <= not (a or b);
    layer2_outputs(5065) <= not (a and b);
    layer2_outputs(5066) <= a and b;
    layer2_outputs(5067) <= not a;
    layer2_outputs(5068) <= not (a and b);
    layer2_outputs(5069) <= b;
    layer2_outputs(5070) <= a xor b;
    layer2_outputs(5071) <= not a;
    layer2_outputs(5072) <= not b;
    layer2_outputs(5073) <= not a;
    layer2_outputs(5074) <= not b or a;
    layer2_outputs(5075) <= not a;
    layer2_outputs(5076) <= not a;
    layer2_outputs(5077) <= not a or b;
    layer2_outputs(5078) <= a and b;
    layer2_outputs(5079) <= not a or b;
    layer2_outputs(5080) <= not a;
    layer2_outputs(5081) <= a;
    layer2_outputs(5082) <= a and not b;
    layer2_outputs(5083) <= a xor b;
    layer2_outputs(5084) <= not b;
    layer2_outputs(5085) <= a;
    layer2_outputs(5086) <= not a;
    layer2_outputs(5087) <= not (a and b);
    layer2_outputs(5088) <= not (a or b);
    layer2_outputs(5089) <= not (a or b);
    layer2_outputs(5090) <= not (a and b);
    layer2_outputs(5091) <= b;
    layer2_outputs(5092) <= b;
    layer2_outputs(5093) <= a;
    layer2_outputs(5094) <= '0';
    layer2_outputs(5095) <= b;
    layer2_outputs(5096) <= not a or b;
    layer2_outputs(5097) <= a;
    layer2_outputs(5098) <= a;
    layer2_outputs(5099) <= not b;
    layer2_outputs(5100) <= not b or a;
    layer2_outputs(5101) <= a;
    layer2_outputs(5102) <= not a;
    layer2_outputs(5103) <= a or b;
    layer2_outputs(5104) <= not a;
    layer2_outputs(5105) <= b;
    layer2_outputs(5106) <= b;
    layer2_outputs(5107) <= not a;
    layer2_outputs(5108) <= a;
    layer2_outputs(5109) <= b and not a;
    layer2_outputs(5110) <= not b;
    layer2_outputs(5111) <= '1';
    layer2_outputs(5112) <= b and not a;
    layer2_outputs(5113) <= not (a or b);
    layer2_outputs(5114) <= a and b;
    layer2_outputs(5115) <= not a;
    layer2_outputs(5116) <= not (a and b);
    layer2_outputs(5117) <= '0';
    layer2_outputs(5118) <= not (a and b);
    layer2_outputs(5119) <= '0';
    layer3_outputs(0) <= not (a and b);
    layer3_outputs(1) <= not a;
    layer3_outputs(2) <= not a;
    layer3_outputs(3) <= not b;
    layer3_outputs(4) <= not a or b;
    layer3_outputs(5) <= not a;
    layer3_outputs(6) <= a and not b;
    layer3_outputs(7) <= a;
    layer3_outputs(8) <= not a;
    layer3_outputs(9) <= not (a and b);
    layer3_outputs(10) <= b;
    layer3_outputs(11) <= not (a and b);
    layer3_outputs(12) <= a;
    layer3_outputs(13) <= b;
    layer3_outputs(14) <= a;
    layer3_outputs(15) <= a and b;
    layer3_outputs(16) <= not (a and b);
    layer3_outputs(17) <= b and not a;
    layer3_outputs(18) <= b;
    layer3_outputs(19) <= not b or a;
    layer3_outputs(20) <= a or b;
    layer3_outputs(21) <= not (a xor b);
    layer3_outputs(22) <= '0';
    layer3_outputs(23) <= b;
    layer3_outputs(24) <= not a;
    layer3_outputs(25) <= a;
    layer3_outputs(26) <= not a;
    layer3_outputs(27) <= a and not b;
    layer3_outputs(28) <= a and not b;
    layer3_outputs(29) <= not a;
    layer3_outputs(30) <= a and b;
    layer3_outputs(31) <= not b;
    layer3_outputs(32) <= not (a and b);
    layer3_outputs(33) <= not a;
    layer3_outputs(34) <= a;
    layer3_outputs(35) <= not b;
    layer3_outputs(36) <= b and not a;
    layer3_outputs(37) <= a and b;
    layer3_outputs(38) <= '1';
    layer3_outputs(39) <= not b or a;
    layer3_outputs(40) <= a and not b;
    layer3_outputs(41) <= not (a xor b);
    layer3_outputs(42) <= a and b;
    layer3_outputs(43) <= not b;
    layer3_outputs(44) <= a or b;
    layer3_outputs(45) <= a;
    layer3_outputs(46) <= b and not a;
    layer3_outputs(47) <= not a;
    layer3_outputs(48) <= a and b;
    layer3_outputs(49) <= not a;
    layer3_outputs(50) <= not b;
    layer3_outputs(51) <= not a or b;
    layer3_outputs(52) <= not (a or b);
    layer3_outputs(53) <= b;
    layer3_outputs(54) <= not a;
    layer3_outputs(55) <= not b;
    layer3_outputs(56) <= not (a or b);
    layer3_outputs(57) <= b and not a;
    layer3_outputs(58) <= not a;
    layer3_outputs(59) <= not (a and b);
    layer3_outputs(60) <= a and b;
    layer3_outputs(61) <= not b or a;
    layer3_outputs(62) <= a and b;
    layer3_outputs(63) <= not (a or b);
    layer3_outputs(64) <= b;
    layer3_outputs(65) <= not a;
    layer3_outputs(66) <= a and b;
    layer3_outputs(67) <= not (a and b);
    layer3_outputs(68) <= not b or a;
    layer3_outputs(69) <= a or b;
    layer3_outputs(70) <= not b;
    layer3_outputs(71) <= a xor b;
    layer3_outputs(72) <= not a;
    layer3_outputs(73) <= b;
    layer3_outputs(74) <= a or b;
    layer3_outputs(75) <= not (a or b);
    layer3_outputs(76) <= b and not a;
    layer3_outputs(77) <= a;
    layer3_outputs(78) <= not b;
    layer3_outputs(79) <= not b or a;
    layer3_outputs(80) <= b and not a;
    layer3_outputs(81) <= not a or b;
    layer3_outputs(82) <= a;
    layer3_outputs(83) <= b;
    layer3_outputs(84) <= a;
    layer3_outputs(85) <= not b;
    layer3_outputs(86) <= not a;
    layer3_outputs(87) <= b and not a;
    layer3_outputs(88) <= a xor b;
    layer3_outputs(89) <= not (a and b);
    layer3_outputs(90) <= a;
    layer3_outputs(91) <= not b;
    layer3_outputs(92) <= a xor b;
    layer3_outputs(93) <= a;
    layer3_outputs(94) <= a and b;
    layer3_outputs(95) <= not a;
    layer3_outputs(96) <= '1';
    layer3_outputs(97) <= not b;
    layer3_outputs(98) <= not b or a;
    layer3_outputs(99) <= '0';
    layer3_outputs(100) <= not b;
    layer3_outputs(101) <= not a;
    layer3_outputs(102) <= b and not a;
    layer3_outputs(103) <= a and b;
    layer3_outputs(104) <= a;
    layer3_outputs(105) <= not b or a;
    layer3_outputs(106) <= a;
    layer3_outputs(107) <= a and b;
    layer3_outputs(108) <= a and b;
    layer3_outputs(109) <= not (a xor b);
    layer3_outputs(110) <= a or b;
    layer3_outputs(111) <= '0';
    layer3_outputs(112) <= a and not b;
    layer3_outputs(113) <= b and not a;
    layer3_outputs(114) <= b;
    layer3_outputs(115) <= b;
    layer3_outputs(116) <= not (a or b);
    layer3_outputs(117) <= not a;
    layer3_outputs(118) <= a;
    layer3_outputs(119) <= '0';
    layer3_outputs(120) <= b;
    layer3_outputs(121) <= a and not b;
    layer3_outputs(122) <= b;
    layer3_outputs(123) <= b and not a;
    layer3_outputs(124) <= not b;
    layer3_outputs(125) <= not b;
    layer3_outputs(126) <= a xor b;
    layer3_outputs(127) <= a;
    layer3_outputs(128) <= not (a or b);
    layer3_outputs(129) <= b and not a;
    layer3_outputs(130) <= not (a and b);
    layer3_outputs(131) <= not b;
    layer3_outputs(132) <= not a or b;
    layer3_outputs(133) <= not b;
    layer3_outputs(134) <= a;
    layer3_outputs(135) <= a;
    layer3_outputs(136) <= not b;
    layer3_outputs(137) <= not b;
    layer3_outputs(138) <= not (a or b);
    layer3_outputs(139) <= a and b;
    layer3_outputs(140) <= a xor b;
    layer3_outputs(141) <= not a;
    layer3_outputs(142) <= b and not a;
    layer3_outputs(143) <= not (a and b);
    layer3_outputs(144) <= not b or a;
    layer3_outputs(145) <= not (a or b);
    layer3_outputs(146) <= not b or a;
    layer3_outputs(147) <= not b;
    layer3_outputs(148) <= not b;
    layer3_outputs(149) <= a;
    layer3_outputs(150) <= not a;
    layer3_outputs(151) <= not a;
    layer3_outputs(152) <= not b;
    layer3_outputs(153) <= not (a xor b);
    layer3_outputs(154) <= b and not a;
    layer3_outputs(155) <= '0';
    layer3_outputs(156) <= '0';
    layer3_outputs(157) <= not b or a;
    layer3_outputs(158) <= a and not b;
    layer3_outputs(159) <= b;
    layer3_outputs(160) <= a xor b;
    layer3_outputs(161) <= '1';
    layer3_outputs(162) <= not (a and b);
    layer3_outputs(163) <= not a;
    layer3_outputs(164) <= not b;
    layer3_outputs(165) <= not a;
    layer3_outputs(166) <= not a;
    layer3_outputs(167) <= b and not a;
    layer3_outputs(168) <= a xor b;
    layer3_outputs(169) <= a;
    layer3_outputs(170) <= not (a and b);
    layer3_outputs(171) <= not a;
    layer3_outputs(172) <= not b or a;
    layer3_outputs(173) <= not a or b;
    layer3_outputs(174) <= not (a or b);
    layer3_outputs(175) <= not b or a;
    layer3_outputs(176) <= a and b;
    layer3_outputs(177) <= a and not b;
    layer3_outputs(178) <= not a;
    layer3_outputs(179) <= a;
    layer3_outputs(180) <= not (a or b);
    layer3_outputs(181) <= b;
    layer3_outputs(182) <= not b or a;
    layer3_outputs(183) <= b and not a;
    layer3_outputs(184) <= a;
    layer3_outputs(185) <= not b or a;
    layer3_outputs(186) <= not (a and b);
    layer3_outputs(187) <= a;
    layer3_outputs(188) <= '1';
    layer3_outputs(189) <= b;
    layer3_outputs(190) <= not b or a;
    layer3_outputs(191) <= a and b;
    layer3_outputs(192) <= not a or b;
    layer3_outputs(193) <= not a or b;
    layer3_outputs(194) <= not (a or b);
    layer3_outputs(195) <= a or b;
    layer3_outputs(196) <= not a;
    layer3_outputs(197) <= not (a and b);
    layer3_outputs(198) <= not (a and b);
    layer3_outputs(199) <= not (a or b);
    layer3_outputs(200) <= b;
    layer3_outputs(201) <= not (a xor b);
    layer3_outputs(202) <= not a;
    layer3_outputs(203) <= not b;
    layer3_outputs(204) <= a xor b;
    layer3_outputs(205) <= b;
    layer3_outputs(206) <= a;
    layer3_outputs(207) <= a and not b;
    layer3_outputs(208) <= b and not a;
    layer3_outputs(209) <= b and not a;
    layer3_outputs(210) <= not (a or b);
    layer3_outputs(211) <= not b;
    layer3_outputs(212) <= not b;
    layer3_outputs(213) <= '1';
    layer3_outputs(214) <= b;
    layer3_outputs(215) <= not b or a;
    layer3_outputs(216) <= a;
    layer3_outputs(217) <= not a;
    layer3_outputs(218) <= '1';
    layer3_outputs(219) <= a;
    layer3_outputs(220) <= a or b;
    layer3_outputs(221) <= not (a and b);
    layer3_outputs(222) <= not a;
    layer3_outputs(223) <= not (a xor b);
    layer3_outputs(224) <= not (a and b);
    layer3_outputs(225) <= a or b;
    layer3_outputs(226) <= not a;
    layer3_outputs(227) <= a;
    layer3_outputs(228) <= b and not a;
    layer3_outputs(229) <= not (a or b);
    layer3_outputs(230) <= a;
    layer3_outputs(231) <= not a;
    layer3_outputs(232) <= not (a and b);
    layer3_outputs(233) <= not (a xor b);
    layer3_outputs(234) <= a or b;
    layer3_outputs(235) <= a or b;
    layer3_outputs(236) <= b;
    layer3_outputs(237) <= not a or b;
    layer3_outputs(238) <= a and not b;
    layer3_outputs(239) <= '1';
    layer3_outputs(240) <= not (a and b);
    layer3_outputs(241) <= not b;
    layer3_outputs(242) <= not (a or b);
    layer3_outputs(243) <= '1';
    layer3_outputs(244) <= not (a or b);
    layer3_outputs(245) <= not a or b;
    layer3_outputs(246) <= not b or a;
    layer3_outputs(247) <= a or b;
    layer3_outputs(248) <= a;
    layer3_outputs(249) <= a xor b;
    layer3_outputs(250) <= not (a or b);
    layer3_outputs(251) <= not b;
    layer3_outputs(252) <= b and not a;
    layer3_outputs(253) <= a or b;
    layer3_outputs(254) <= not b;
    layer3_outputs(255) <= not a or b;
    layer3_outputs(256) <= a and not b;
    layer3_outputs(257) <= not a;
    layer3_outputs(258) <= b;
    layer3_outputs(259) <= a;
    layer3_outputs(260) <= not (a or b);
    layer3_outputs(261) <= '0';
    layer3_outputs(262) <= not (a or b);
    layer3_outputs(263) <= not b or a;
    layer3_outputs(264) <= not b or a;
    layer3_outputs(265) <= not (a or b);
    layer3_outputs(266) <= not a or b;
    layer3_outputs(267) <= not b or a;
    layer3_outputs(268) <= a and not b;
    layer3_outputs(269) <= b and not a;
    layer3_outputs(270) <= not b;
    layer3_outputs(271) <= not (a and b);
    layer3_outputs(272) <= not b;
    layer3_outputs(273) <= b;
    layer3_outputs(274) <= not a;
    layer3_outputs(275) <= not b;
    layer3_outputs(276) <= b;
    layer3_outputs(277) <= not (a or b);
    layer3_outputs(278) <= b;
    layer3_outputs(279) <= not a or b;
    layer3_outputs(280) <= not (a or b);
    layer3_outputs(281) <= a and not b;
    layer3_outputs(282) <= not b;
    layer3_outputs(283) <= b;
    layer3_outputs(284) <= not a;
    layer3_outputs(285) <= a or b;
    layer3_outputs(286) <= not a;
    layer3_outputs(287) <= b and not a;
    layer3_outputs(288) <= a and not b;
    layer3_outputs(289) <= b and not a;
    layer3_outputs(290) <= not b;
    layer3_outputs(291) <= a;
    layer3_outputs(292) <= b;
    layer3_outputs(293) <= b and not a;
    layer3_outputs(294) <= not b;
    layer3_outputs(295) <= a and b;
    layer3_outputs(296) <= not (a and b);
    layer3_outputs(297) <= not a or b;
    layer3_outputs(298) <= not a;
    layer3_outputs(299) <= not (a xor b);
    layer3_outputs(300) <= not a or b;
    layer3_outputs(301) <= b;
    layer3_outputs(302) <= not (a and b);
    layer3_outputs(303) <= not (a and b);
    layer3_outputs(304) <= not b;
    layer3_outputs(305) <= not (a and b);
    layer3_outputs(306) <= b and not a;
    layer3_outputs(307) <= b;
    layer3_outputs(308) <= b;
    layer3_outputs(309) <= a and b;
    layer3_outputs(310) <= not a;
    layer3_outputs(311) <= a or b;
    layer3_outputs(312) <= not b;
    layer3_outputs(313) <= not (a and b);
    layer3_outputs(314) <= not (a and b);
    layer3_outputs(315) <= b and not a;
    layer3_outputs(316) <= a xor b;
    layer3_outputs(317) <= a xor b;
    layer3_outputs(318) <= not b;
    layer3_outputs(319) <= not (a and b);
    layer3_outputs(320) <= b;
    layer3_outputs(321) <= not b;
    layer3_outputs(322) <= b;
    layer3_outputs(323) <= '0';
    layer3_outputs(324) <= b and not a;
    layer3_outputs(325) <= not (a xor b);
    layer3_outputs(326) <= not b;
    layer3_outputs(327) <= not a;
    layer3_outputs(328) <= not a;
    layer3_outputs(329) <= a;
    layer3_outputs(330) <= not a or b;
    layer3_outputs(331) <= a and not b;
    layer3_outputs(332) <= a;
    layer3_outputs(333) <= a and not b;
    layer3_outputs(334) <= a or b;
    layer3_outputs(335) <= not (a xor b);
    layer3_outputs(336) <= a;
    layer3_outputs(337) <= not a;
    layer3_outputs(338) <= '1';
    layer3_outputs(339) <= not b;
    layer3_outputs(340) <= not b;
    layer3_outputs(341) <= not a;
    layer3_outputs(342) <= not (a xor b);
    layer3_outputs(343) <= a or b;
    layer3_outputs(344) <= not b;
    layer3_outputs(345) <= not a or b;
    layer3_outputs(346) <= b and not a;
    layer3_outputs(347) <= a and b;
    layer3_outputs(348) <= a and b;
    layer3_outputs(349) <= b;
    layer3_outputs(350) <= not a;
    layer3_outputs(351) <= a;
    layer3_outputs(352) <= a and not b;
    layer3_outputs(353) <= a and b;
    layer3_outputs(354) <= not (a and b);
    layer3_outputs(355) <= a and not b;
    layer3_outputs(356) <= a and not b;
    layer3_outputs(357) <= not (a or b);
    layer3_outputs(358) <= a and b;
    layer3_outputs(359) <= b;
    layer3_outputs(360) <= a or b;
    layer3_outputs(361) <= b and not a;
    layer3_outputs(362) <= a or b;
    layer3_outputs(363) <= a and b;
    layer3_outputs(364) <= b and not a;
    layer3_outputs(365) <= a;
    layer3_outputs(366) <= not (a and b);
    layer3_outputs(367) <= not b;
    layer3_outputs(368) <= b;
    layer3_outputs(369) <= a xor b;
    layer3_outputs(370) <= b;
    layer3_outputs(371) <= a and b;
    layer3_outputs(372) <= not b or a;
    layer3_outputs(373) <= not a;
    layer3_outputs(374) <= not (a or b);
    layer3_outputs(375) <= a or b;
    layer3_outputs(376) <= a and not b;
    layer3_outputs(377) <= not b or a;
    layer3_outputs(378) <= not a;
    layer3_outputs(379) <= not b;
    layer3_outputs(380) <= not (a and b);
    layer3_outputs(381) <= not b;
    layer3_outputs(382) <= not a or b;
    layer3_outputs(383) <= b;
    layer3_outputs(384) <= not (a or b);
    layer3_outputs(385) <= b and not a;
    layer3_outputs(386) <= not b;
    layer3_outputs(387) <= b and not a;
    layer3_outputs(388) <= a or b;
    layer3_outputs(389) <= a or b;
    layer3_outputs(390) <= '0';
    layer3_outputs(391) <= not (a xor b);
    layer3_outputs(392) <= a and not b;
    layer3_outputs(393) <= not b or a;
    layer3_outputs(394) <= b and not a;
    layer3_outputs(395) <= a and not b;
    layer3_outputs(396) <= a;
    layer3_outputs(397) <= a xor b;
    layer3_outputs(398) <= a or b;
    layer3_outputs(399) <= b and not a;
    layer3_outputs(400) <= b;
    layer3_outputs(401) <= a and not b;
    layer3_outputs(402) <= b;
    layer3_outputs(403) <= not (a or b);
    layer3_outputs(404) <= b;
    layer3_outputs(405) <= a;
    layer3_outputs(406) <= not (a xor b);
    layer3_outputs(407) <= not a or b;
    layer3_outputs(408) <= a and not b;
    layer3_outputs(409) <= not (a and b);
    layer3_outputs(410) <= a or b;
    layer3_outputs(411) <= a;
    layer3_outputs(412) <= not (a or b);
    layer3_outputs(413) <= a;
    layer3_outputs(414) <= a;
    layer3_outputs(415) <= b and not a;
    layer3_outputs(416) <= b and not a;
    layer3_outputs(417) <= '1';
    layer3_outputs(418) <= '0';
    layer3_outputs(419) <= not (a and b);
    layer3_outputs(420) <= not a;
    layer3_outputs(421) <= not b or a;
    layer3_outputs(422) <= not a;
    layer3_outputs(423) <= not (a and b);
    layer3_outputs(424) <= not b;
    layer3_outputs(425) <= b and not a;
    layer3_outputs(426) <= b;
    layer3_outputs(427) <= not a;
    layer3_outputs(428) <= b;
    layer3_outputs(429) <= not b;
    layer3_outputs(430) <= not b;
    layer3_outputs(431) <= a;
    layer3_outputs(432) <= not b;
    layer3_outputs(433) <= a and not b;
    layer3_outputs(434) <= not b;
    layer3_outputs(435) <= b;
    layer3_outputs(436) <= a xor b;
    layer3_outputs(437) <= a and b;
    layer3_outputs(438) <= b;
    layer3_outputs(439) <= b;
    layer3_outputs(440) <= not a;
    layer3_outputs(441) <= b;
    layer3_outputs(442) <= b;
    layer3_outputs(443) <= not (a xor b);
    layer3_outputs(444) <= not b or a;
    layer3_outputs(445) <= not a;
    layer3_outputs(446) <= '0';
    layer3_outputs(447) <= not (a or b);
    layer3_outputs(448) <= not (a or b);
    layer3_outputs(449) <= not b;
    layer3_outputs(450) <= not (a xor b);
    layer3_outputs(451) <= not b;
    layer3_outputs(452) <= b;
    layer3_outputs(453) <= not a or b;
    layer3_outputs(454) <= '0';
    layer3_outputs(455) <= not a or b;
    layer3_outputs(456) <= not b;
    layer3_outputs(457) <= not (a and b);
    layer3_outputs(458) <= a or b;
    layer3_outputs(459) <= not (a or b);
    layer3_outputs(460) <= b and not a;
    layer3_outputs(461) <= not a;
    layer3_outputs(462) <= not (a and b);
    layer3_outputs(463) <= not a;
    layer3_outputs(464) <= a xor b;
    layer3_outputs(465) <= not (a or b);
    layer3_outputs(466) <= not (a or b);
    layer3_outputs(467) <= not b or a;
    layer3_outputs(468) <= b;
    layer3_outputs(469) <= not b;
    layer3_outputs(470) <= b;
    layer3_outputs(471) <= not a;
    layer3_outputs(472) <= a and b;
    layer3_outputs(473) <= not a;
    layer3_outputs(474) <= a;
    layer3_outputs(475) <= not (a xor b);
    layer3_outputs(476) <= not (a xor b);
    layer3_outputs(477) <= a and not b;
    layer3_outputs(478) <= a or b;
    layer3_outputs(479) <= not (a xor b);
    layer3_outputs(480) <= a and not b;
    layer3_outputs(481) <= a;
    layer3_outputs(482) <= not a or b;
    layer3_outputs(483) <= not a or b;
    layer3_outputs(484) <= a;
    layer3_outputs(485) <= not a;
    layer3_outputs(486) <= a;
    layer3_outputs(487) <= not (a and b);
    layer3_outputs(488) <= b and not a;
    layer3_outputs(489) <= not b;
    layer3_outputs(490) <= a or b;
    layer3_outputs(491) <= a and b;
    layer3_outputs(492) <= not a or b;
    layer3_outputs(493) <= a and not b;
    layer3_outputs(494) <= not (a or b);
    layer3_outputs(495) <= b;
    layer3_outputs(496) <= not b;
    layer3_outputs(497) <= b;
    layer3_outputs(498) <= not a;
    layer3_outputs(499) <= not (a and b);
    layer3_outputs(500) <= '1';
    layer3_outputs(501) <= a;
    layer3_outputs(502) <= a or b;
    layer3_outputs(503) <= b;
    layer3_outputs(504) <= a;
    layer3_outputs(505) <= a and not b;
    layer3_outputs(506) <= a xor b;
    layer3_outputs(507) <= not (a xor b);
    layer3_outputs(508) <= not a or b;
    layer3_outputs(509) <= not b;
    layer3_outputs(510) <= b and not a;
    layer3_outputs(511) <= a or b;
    layer3_outputs(512) <= a and b;
    layer3_outputs(513) <= a;
    layer3_outputs(514) <= b;
    layer3_outputs(515) <= b and not a;
    layer3_outputs(516) <= b and not a;
    layer3_outputs(517) <= not a;
    layer3_outputs(518) <= not (a xor b);
    layer3_outputs(519) <= a and not b;
    layer3_outputs(520) <= a and not b;
    layer3_outputs(521) <= not b;
    layer3_outputs(522) <= not b or a;
    layer3_outputs(523) <= not (a or b);
    layer3_outputs(524) <= a;
    layer3_outputs(525) <= not b;
    layer3_outputs(526) <= not b;
    layer3_outputs(527) <= not a;
    layer3_outputs(528) <= a or b;
    layer3_outputs(529) <= '0';
    layer3_outputs(530) <= not a or b;
    layer3_outputs(531) <= not a;
    layer3_outputs(532) <= b;
    layer3_outputs(533) <= a and b;
    layer3_outputs(534) <= b;
    layer3_outputs(535) <= a;
    layer3_outputs(536) <= a or b;
    layer3_outputs(537) <= not a or b;
    layer3_outputs(538) <= a or b;
    layer3_outputs(539) <= not (a and b);
    layer3_outputs(540) <= not b or a;
    layer3_outputs(541) <= b;
    layer3_outputs(542) <= '0';
    layer3_outputs(543) <= not (a xor b);
    layer3_outputs(544) <= not b or a;
    layer3_outputs(545) <= b;
    layer3_outputs(546) <= not (a or b);
    layer3_outputs(547) <= not (a xor b);
    layer3_outputs(548) <= not (a or b);
    layer3_outputs(549) <= a xor b;
    layer3_outputs(550) <= b;
    layer3_outputs(551) <= not a;
    layer3_outputs(552) <= not b;
    layer3_outputs(553) <= a;
    layer3_outputs(554) <= a or b;
    layer3_outputs(555) <= not b or a;
    layer3_outputs(556) <= a;
    layer3_outputs(557) <= a or b;
    layer3_outputs(558) <= b;
    layer3_outputs(559) <= not (a xor b);
    layer3_outputs(560) <= not b or a;
    layer3_outputs(561) <= not (a or b);
    layer3_outputs(562) <= a;
    layer3_outputs(563) <= not a or b;
    layer3_outputs(564) <= a;
    layer3_outputs(565) <= not (a xor b);
    layer3_outputs(566) <= a;
    layer3_outputs(567) <= a xor b;
    layer3_outputs(568) <= not (a or b);
    layer3_outputs(569) <= a;
    layer3_outputs(570) <= a or b;
    layer3_outputs(571) <= '1';
    layer3_outputs(572) <= not a or b;
    layer3_outputs(573) <= not (a or b);
    layer3_outputs(574) <= not a or b;
    layer3_outputs(575) <= a and not b;
    layer3_outputs(576) <= not a or b;
    layer3_outputs(577) <= b;
    layer3_outputs(578) <= b;
    layer3_outputs(579) <= a and not b;
    layer3_outputs(580) <= a and not b;
    layer3_outputs(581) <= a or b;
    layer3_outputs(582) <= a;
    layer3_outputs(583) <= b and not a;
    layer3_outputs(584) <= not (a and b);
    layer3_outputs(585) <= a;
    layer3_outputs(586) <= not a;
    layer3_outputs(587) <= not (a or b);
    layer3_outputs(588) <= a or b;
    layer3_outputs(589) <= not (a or b);
    layer3_outputs(590) <= not b;
    layer3_outputs(591) <= not a or b;
    layer3_outputs(592) <= a xor b;
    layer3_outputs(593) <= a and not b;
    layer3_outputs(594) <= a and b;
    layer3_outputs(595) <= b;
    layer3_outputs(596) <= not (a and b);
    layer3_outputs(597) <= not b or a;
    layer3_outputs(598) <= not (a or b);
    layer3_outputs(599) <= not b or a;
    layer3_outputs(600) <= a;
    layer3_outputs(601) <= not (a or b);
    layer3_outputs(602) <= not a or b;
    layer3_outputs(603) <= not b;
    layer3_outputs(604) <= b and not a;
    layer3_outputs(605) <= not a;
    layer3_outputs(606) <= b and not a;
    layer3_outputs(607) <= not a;
    layer3_outputs(608) <= a;
    layer3_outputs(609) <= not b;
    layer3_outputs(610) <= not (a or b);
    layer3_outputs(611) <= not b or a;
    layer3_outputs(612) <= not (a or b);
    layer3_outputs(613) <= b;
    layer3_outputs(614) <= a and b;
    layer3_outputs(615) <= a and b;
    layer3_outputs(616) <= a and b;
    layer3_outputs(617) <= b;
    layer3_outputs(618) <= not (a xor b);
    layer3_outputs(619) <= '0';
    layer3_outputs(620) <= b;
    layer3_outputs(621) <= b;
    layer3_outputs(622) <= b;
    layer3_outputs(623) <= b;
    layer3_outputs(624) <= not b or a;
    layer3_outputs(625) <= a and b;
    layer3_outputs(626) <= not (a xor b);
    layer3_outputs(627) <= not (a and b);
    layer3_outputs(628) <= not a;
    layer3_outputs(629) <= not b;
    layer3_outputs(630) <= not (a and b);
    layer3_outputs(631) <= a;
    layer3_outputs(632) <= b;
    layer3_outputs(633) <= b;
    layer3_outputs(634) <= not a;
    layer3_outputs(635) <= not a;
    layer3_outputs(636) <= not b;
    layer3_outputs(637) <= b;
    layer3_outputs(638) <= b;
    layer3_outputs(639) <= b and not a;
    layer3_outputs(640) <= b and not a;
    layer3_outputs(641) <= not b or a;
    layer3_outputs(642) <= a or b;
    layer3_outputs(643) <= a or b;
    layer3_outputs(644) <= not a;
    layer3_outputs(645) <= b;
    layer3_outputs(646) <= not a or b;
    layer3_outputs(647) <= not (a and b);
    layer3_outputs(648) <= a;
    layer3_outputs(649) <= not b or a;
    layer3_outputs(650) <= not b;
    layer3_outputs(651) <= not (a or b);
    layer3_outputs(652) <= a xor b;
    layer3_outputs(653) <= a;
    layer3_outputs(654) <= '0';
    layer3_outputs(655) <= a or b;
    layer3_outputs(656) <= not a;
    layer3_outputs(657) <= a;
    layer3_outputs(658) <= a and not b;
    layer3_outputs(659) <= not b or a;
    layer3_outputs(660) <= not (a or b);
    layer3_outputs(661) <= not (a xor b);
    layer3_outputs(662) <= a xor b;
    layer3_outputs(663) <= a and b;
    layer3_outputs(664) <= a or b;
    layer3_outputs(665) <= b and not a;
    layer3_outputs(666) <= b;
    layer3_outputs(667) <= a;
    layer3_outputs(668) <= not b;
    layer3_outputs(669) <= not a;
    layer3_outputs(670) <= b;
    layer3_outputs(671) <= not a;
    layer3_outputs(672) <= not a;
    layer3_outputs(673) <= not (a and b);
    layer3_outputs(674) <= b;
    layer3_outputs(675) <= a and not b;
    layer3_outputs(676) <= not a or b;
    layer3_outputs(677) <= not (a and b);
    layer3_outputs(678) <= not b or a;
    layer3_outputs(679) <= a;
    layer3_outputs(680) <= not (a or b);
    layer3_outputs(681) <= not b;
    layer3_outputs(682) <= not (a xor b);
    layer3_outputs(683) <= not (a and b);
    layer3_outputs(684) <= not (a or b);
    layer3_outputs(685) <= a;
    layer3_outputs(686) <= not (a or b);
    layer3_outputs(687) <= a or b;
    layer3_outputs(688) <= not b or a;
    layer3_outputs(689) <= not (a or b);
    layer3_outputs(690) <= not a;
    layer3_outputs(691) <= not a;
    layer3_outputs(692) <= b;
    layer3_outputs(693) <= b and not a;
    layer3_outputs(694) <= not (a and b);
    layer3_outputs(695) <= not (a xor b);
    layer3_outputs(696) <= a and not b;
    layer3_outputs(697) <= not b;
    layer3_outputs(698) <= not a;
    layer3_outputs(699) <= a;
    layer3_outputs(700) <= not b or a;
    layer3_outputs(701) <= b;
    layer3_outputs(702) <= a or b;
    layer3_outputs(703) <= not a or b;
    layer3_outputs(704) <= b and not a;
    layer3_outputs(705) <= a or b;
    layer3_outputs(706) <= a or b;
    layer3_outputs(707) <= not a;
    layer3_outputs(708) <= b;
    layer3_outputs(709) <= not a or b;
    layer3_outputs(710) <= a and b;
    layer3_outputs(711) <= a and not b;
    layer3_outputs(712) <= not (a and b);
    layer3_outputs(713) <= b;
    layer3_outputs(714) <= a xor b;
    layer3_outputs(715) <= not (a xor b);
    layer3_outputs(716) <= b;
    layer3_outputs(717) <= not a;
    layer3_outputs(718) <= a;
    layer3_outputs(719) <= a;
    layer3_outputs(720) <= not a;
    layer3_outputs(721) <= a;
    layer3_outputs(722) <= not b;
    layer3_outputs(723) <= not b;
    layer3_outputs(724) <= a or b;
    layer3_outputs(725) <= not (a xor b);
    layer3_outputs(726) <= not a or b;
    layer3_outputs(727) <= not b;
    layer3_outputs(728) <= '1';
    layer3_outputs(729) <= not a or b;
    layer3_outputs(730) <= not (a and b);
    layer3_outputs(731) <= not a or b;
    layer3_outputs(732) <= '1';
    layer3_outputs(733) <= not (a and b);
    layer3_outputs(734) <= a;
    layer3_outputs(735) <= not b;
    layer3_outputs(736) <= b and not a;
    layer3_outputs(737) <= b;
    layer3_outputs(738) <= b and not a;
    layer3_outputs(739) <= not b;
    layer3_outputs(740) <= not b;
    layer3_outputs(741) <= b;
    layer3_outputs(742) <= not a or b;
    layer3_outputs(743) <= not b;
    layer3_outputs(744) <= a and not b;
    layer3_outputs(745) <= not a;
    layer3_outputs(746) <= a and b;
    layer3_outputs(747) <= not b or a;
    layer3_outputs(748) <= a xor b;
    layer3_outputs(749) <= not b or a;
    layer3_outputs(750) <= not b or a;
    layer3_outputs(751) <= not a or b;
    layer3_outputs(752) <= a;
    layer3_outputs(753) <= not a or b;
    layer3_outputs(754) <= a;
    layer3_outputs(755) <= b and not a;
    layer3_outputs(756) <= not (a or b);
    layer3_outputs(757) <= '0';
    layer3_outputs(758) <= b;
    layer3_outputs(759) <= a and b;
    layer3_outputs(760) <= not b or a;
    layer3_outputs(761) <= a;
    layer3_outputs(762) <= a xor b;
    layer3_outputs(763) <= not (a and b);
    layer3_outputs(764) <= not (a or b);
    layer3_outputs(765) <= not (a or b);
    layer3_outputs(766) <= b;
    layer3_outputs(767) <= not a or b;
    layer3_outputs(768) <= a;
    layer3_outputs(769) <= not (a xor b);
    layer3_outputs(770) <= not a;
    layer3_outputs(771) <= a;
    layer3_outputs(772) <= not a or b;
    layer3_outputs(773) <= b and not a;
    layer3_outputs(774) <= a or b;
    layer3_outputs(775) <= a xor b;
    layer3_outputs(776) <= not (a or b);
    layer3_outputs(777) <= not a or b;
    layer3_outputs(778) <= a and b;
    layer3_outputs(779) <= not a;
    layer3_outputs(780) <= not (a or b);
    layer3_outputs(781) <= not b;
    layer3_outputs(782) <= a or b;
    layer3_outputs(783) <= a;
    layer3_outputs(784) <= not b or a;
    layer3_outputs(785) <= b and not a;
    layer3_outputs(786) <= not b or a;
    layer3_outputs(787) <= not (a xor b);
    layer3_outputs(788) <= b and not a;
    layer3_outputs(789) <= not (a or b);
    layer3_outputs(790) <= not a;
    layer3_outputs(791) <= '0';
    layer3_outputs(792) <= not (a or b);
    layer3_outputs(793) <= a and not b;
    layer3_outputs(794) <= a or b;
    layer3_outputs(795) <= a and not b;
    layer3_outputs(796) <= a;
    layer3_outputs(797) <= not b;
    layer3_outputs(798) <= b;
    layer3_outputs(799) <= '1';
    layer3_outputs(800) <= b and not a;
    layer3_outputs(801) <= a or b;
    layer3_outputs(802) <= not a or b;
    layer3_outputs(803) <= not b or a;
    layer3_outputs(804) <= not b;
    layer3_outputs(805) <= not (a xor b);
    layer3_outputs(806) <= a xor b;
    layer3_outputs(807) <= a;
    layer3_outputs(808) <= a and b;
    layer3_outputs(809) <= a and not b;
    layer3_outputs(810) <= '1';
    layer3_outputs(811) <= b and not a;
    layer3_outputs(812) <= b;
    layer3_outputs(813) <= not b;
    layer3_outputs(814) <= not a;
    layer3_outputs(815) <= not b;
    layer3_outputs(816) <= not (a and b);
    layer3_outputs(817) <= b and not a;
    layer3_outputs(818) <= '1';
    layer3_outputs(819) <= not (a xor b);
    layer3_outputs(820) <= not (a or b);
    layer3_outputs(821) <= b and not a;
    layer3_outputs(822) <= not b or a;
    layer3_outputs(823) <= a xor b;
    layer3_outputs(824) <= not a;
    layer3_outputs(825) <= a xor b;
    layer3_outputs(826) <= a or b;
    layer3_outputs(827) <= a and b;
    layer3_outputs(828) <= a;
    layer3_outputs(829) <= b and not a;
    layer3_outputs(830) <= b;
    layer3_outputs(831) <= a and not b;
    layer3_outputs(832) <= b;
    layer3_outputs(833) <= b and not a;
    layer3_outputs(834) <= not a;
    layer3_outputs(835) <= not a or b;
    layer3_outputs(836) <= not a or b;
    layer3_outputs(837) <= not a;
    layer3_outputs(838) <= not (a or b);
    layer3_outputs(839) <= a and not b;
    layer3_outputs(840) <= a and b;
    layer3_outputs(841) <= not (a and b);
    layer3_outputs(842) <= a xor b;
    layer3_outputs(843) <= a and b;
    layer3_outputs(844) <= a;
    layer3_outputs(845) <= not b or a;
    layer3_outputs(846) <= a and b;
    layer3_outputs(847) <= not b;
    layer3_outputs(848) <= a xor b;
    layer3_outputs(849) <= b and not a;
    layer3_outputs(850) <= not a;
    layer3_outputs(851) <= not (a xor b);
    layer3_outputs(852) <= b;
    layer3_outputs(853) <= b and not a;
    layer3_outputs(854) <= a or b;
    layer3_outputs(855) <= not a or b;
    layer3_outputs(856) <= not (a and b);
    layer3_outputs(857) <= not a;
    layer3_outputs(858) <= '1';
    layer3_outputs(859) <= b and not a;
    layer3_outputs(860) <= not b;
    layer3_outputs(861) <= not b or a;
    layer3_outputs(862) <= not (a xor b);
    layer3_outputs(863) <= a xor b;
    layer3_outputs(864) <= a;
    layer3_outputs(865) <= not a or b;
    layer3_outputs(866) <= b;
    layer3_outputs(867) <= a;
    layer3_outputs(868) <= a and not b;
    layer3_outputs(869) <= a and not b;
    layer3_outputs(870) <= not a or b;
    layer3_outputs(871) <= a;
    layer3_outputs(872) <= a and b;
    layer3_outputs(873) <= not a or b;
    layer3_outputs(874) <= not b;
    layer3_outputs(875) <= not (a xor b);
    layer3_outputs(876) <= not (a xor b);
    layer3_outputs(877) <= not a or b;
    layer3_outputs(878) <= a or b;
    layer3_outputs(879) <= a or b;
    layer3_outputs(880) <= a;
    layer3_outputs(881) <= not (a and b);
    layer3_outputs(882) <= a;
    layer3_outputs(883) <= a;
    layer3_outputs(884) <= a;
    layer3_outputs(885) <= not b or a;
    layer3_outputs(886) <= a and b;
    layer3_outputs(887) <= a;
    layer3_outputs(888) <= not a;
    layer3_outputs(889) <= not b;
    layer3_outputs(890) <= a or b;
    layer3_outputs(891) <= a and b;
    layer3_outputs(892) <= not (a or b);
    layer3_outputs(893) <= a and b;
    layer3_outputs(894) <= b;
    layer3_outputs(895) <= not (a xor b);
    layer3_outputs(896) <= not a;
    layer3_outputs(897) <= a and not b;
    layer3_outputs(898) <= a;
    layer3_outputs(899) <= not b;
    layer3_outputs(900) <= a xor b;
    layer3_outputs(901) <= a xor b;
    layer3_outputs(902) <= not a;
    layer3_outputs(903) <= a xor b;
    layer3_outputs(904) <= not (a or b);
    layer3_outputs(905) <= not b or a;
    layer3_outputs(906) <= '0';
    layer3_outputs(907) <= b;
    layer3_outputs(908) <= not a;
    layer3_outputs(909) <= not b;
    layer3_outputs(910) <= not a or b;
    layer3_outputs(911) <= a and b;
    layer3_outputs(912) <= not b or a;
    layer3_outputs(913) <= not a;
    layer3_outputs(914) <= a;
    layer3_outputs(915) <= not (a and b);
    layer3_outputs(916) <= not a or b;
    layer3_outputs(917) <= a;
    layer3_outputs(918) <= b;
    layer3_outputs(919) <= a or b;
    layer3_outputs(920) <= not a;
    layer3_outputs(921) <= a xor b;
    layer3_outputs(922) <= a or b;
    layer3_outputs(923) <= not b;
    layer3_outputs(924) <= a;
    layer3_outputs(925) <= not b;
    layer3_outputs(926) <= a;
    layer3_outputs(927) <= b and not a;
    layer3_outputs(928) <= a and not b;
    layer3_outputs(929) <= b;
    layer3_outputs(930) <= b;
    layer3_outputs(931) <= a xor b;
    layer3_outputs(932) <= not b;
    layer3_outputs(933) <= a;
    layer3_outputs(934) <= not a;
    layer3_outputs(935) <= not a or b;
    layer3_outputs(936) <= a;
    layer3_outputs(937) <= not (a or b);
    layer3_outputs(938) <= not (a or b);
    layer3_outputs(939) <= a and b;
    layer3_outputs(940) <= a;
    layer3_outputs(941) <= a and not b;
    layer3_outputs(942) <= not a;
    layer3_outputs(943) <= b;
    layer3_outputs(944) <= a and not b;
    layer3_outputs(945) <= not (a or b);
    layer3_outputs(946) <= b;
    layer3_outputs(947) <= a or b;
    layer3_outputs(948) <= not a;
    layer3_outputs(949) <= not (a or b);
    layer3_outputs(950) <= a xor b;
    layer3_outputs(951) <= not b;
    layer3_outputs(952) <= a xor b;
    layer3_outputs(953) <= not a or b;
    layer3_outputs(954) <= not b;
    layer3_outputs(955) <= a and not b;
    layer3_outputs(956) <= a and b;
    layer3_outputs(957) <= not a;
    layer3_outputs(958) <= not a;
    layer3_outputs(959) <= not a or b;
    layer3_outputs(960) <= not b;
    layer3_outputs(961) <= not (a xor b);
    layer3_outputs(962) <= not b;
    layer3_outputs(963) <= not a;
    layer3_outputs(964) <= b and not a;
    layer3_outputs(965) <= not a;
    layer3_outputs(966) <= not a or b;
    layer3_outputs(967) <= not (a and b);
    layer3_outputs(968) <= b;
    layer3_outputs(969) <= a and not b;
    layer3_outputs(970) <= not b;
    layer3_outputs(971) <= a and b;
    layer3_outputs(972) <= b and not a;
    layer3_outputs(973) <= not b;
    layer3_outputs(974) <= a or b;
    layer3_outputs(975) <= not (a and b);
    layer3_outputs(976) <= not a;
    layer3_outputs(977) <= not b or a;
    layer3_outputs(978) <= not b or a;
    layer3_outputs(979) <= not b;
    layer3_outputs(980) <= not b;
    layer3_outputs(981) <= '0';
    layer3_outputs(982) <= not b;
    layer3_outputs(983) <= not (a or b);
    layer3_outputs(984) <= b;
    layer3_outputs(985) <= not (a and b);
    layer3_outputs(986) <= b and not a;
    layer3_outputs(987) <= a;
    layer3_outputs(988) <= a xor b;
    layer3_outputs(989) <= a;
    layer3_outputs(990) <= a xor b;
    layer3_outputs(991) <= a;
    layer3_outputs(992) <= b;
    layer3_outputs(993) <= b and not a;
    layer3_outputs(994) <= a xor b;
    layer3_outputs(995) <= a or b;
    layer3_outputs(996) <= a and b;
    layer3_outputs(997) <= a and not b;
    layer3_outputs(998) <= b and not a;
    layer3_outputs(999) <= not a or b;
    layer3_outputs(1000) <= b and not a;
    layer3_outputs(1001) <= a;
    layer3_outputs(1002) <= b;
    layer3_outputs(1003) <= a or b;
    layer3_outputs(1004) <= a xor b;
    layer3_outputs(1005) <= a or b;
    layer3_outputs(1006) <= not a;
    layer3_outputs(1007) <= b;
    layer3_outputs(1008) <= '1';
    layer3_outputs(1009) <= not (a and b);
    layer3_outputs(1010) <= a and b;
    layer3_outputs(1011) <= '1';
    layer3_outputs(1012) <= b and not a;
    layer3_outputs(1013) <= not b;
    layer3_outputs(1014) <= not a or b;
    layer3_outputs(1015) <= a and not b;
    layer3_outputs(1016) <= not a;
    layer3_outputs(1017) <= not a or b;
    layer3_outputs(1018) <= b and not a;
    layer3_outputs(1019) <= not (a and b);
    layer3_outputs(1020) <= a;
    layer3_outputs(1021) <= a or b;
    layer3_outputs(1022) <= a;
    layer3_outputs(1023) <= '1';
    layer3_outputs(1024) <= a;
    layer3_outputs(1025) <= not a;
    layer3_outputs(1026) <= not b;
    layer3_outputs(1027) <= b;
    layer3_outputs(1028) <= a;
    layer3_outputs(1029) <= not b;
    layer3_outputs(1030) <= b;
    layer3_outputs(1031) <= a;
    layer3_outputs(1032) <= b and not a;
    layer3_outputs(1033) <= a;
    layer3_outputs(1034) <= '0';
    layer3_outputs(1035) <= b;
    layer3_outputs(1036) <= b and not a;
    layer3_outputs(1037) <= not b;
    layer3_outputs(1038) <= not (a xor b);
    layer3_outputs(1039) <= not a;
    layer3_outputs(1040) <= not a or b;
    layer3_outputs(1041) <= not b or a;
    layer3_outputs(1042) <= not a;
    layer3_outputs(1043) <= not a or b;
    layer3_outputs(1044) <= not a;
    layer3_outputs(1045) <= not b or a;
    layer3_outputs(1046) <= a;
    layer3_outputs(1047) <= not a or b;
    layer3_outputs(1048) <= a xor b;
    layer3_outputs(1049) <= not b or a;
    layer3_outputs(1050) <= a or b;
    layer3_outputs(1051) <= not a or b;
    layer3_outputs(1052) <= a;
    layer3_outputs(1053) <= not a;
    layer3_outputs(1054) <= not a or b;
    layer3_outputs(1055) <= not a;
    layer3_outputs(1056) <= b and not a;
    layer3_outputs(1057) <= a and not b;
    layer3_outputs(1058) <= a;
    layer3_outputs(1059) <= a or b;
    layer3_outputs(1060) <= not a;
    layer3_outputs(1061) <= a;
    layer3_outputs(1062) <= not a;
    layer3_outputs(1063) <= a;
    layer3_outputs(1064) <= b;
    layer3_outputs(1065) <= not (a and b);
    layer3_outputs(1066) <= not (a and b);
    layer3_outputs(1067) <= a;
    layer3_outputs(1068) <= a or b;
    layer3_outputs(1069) <= b and not a;
    layer3_outputs(1070) <= not b;
    layer3_outputs(1071) <= '1';
    layer3_outputs(1072) <= a and not b;
    layer3_outputs(1073) <= not (a or b);
    layer3_outputs(1074) <= b;
    layer3_outputs(1075) <= not (a and b);
    layer3_outputs(1076) <= a and b;
    layer3_outputs(1077) <= a;
    layer3_outputs(1078) <= not (a and b);
    layer3_outputs(1079) <= not a;
    layer3_outputs(1080) <= a and b;
    layer3_outputs(1081) <= b and not a;
    layer3_outputs(1082) <= not a;
    layer3_outputs(1083) <= not b;
    layer3_outputs(1084) <= not (a and b);
    layer3_outputs(1085) <= b;
    layer3_outputs(1086) <= a;
    layer3_outputs(1087) <= a xor b;
    layer3_outputs(1088) <= not a or b;
    layer3_outputs(1089) <= a or b;
    layer3_outputs(1090) <= not a or b;
    layer3_outputs(1091) <= not a;
    layer3_outputs(1092) <= not a;
    layer3_outputs(1093) <= a and b;
    layer3_outputs(1094) <= a;
    layer3_outputs(1095) <= not (a or b);
    layer3_outputs(1096) <= a xor b;
    layer3_outputs(1097) <= not (a or b);
    layer3_outputs(1098) <= a or b;
    layer3_outputs(1099) <= a and not b;
    layer3_outputs(1100) <= not (a xor b);
    layer3_outputs(1101) <= not (a and b);
    layer3_outputs(1102) <= a or b;
    layer3_outputs(1103) <= not b;
    layer3_outputs(1104) <= not a or b;
    layer3_outputs(1105) <= not b;
    layer3_outputs(1106) <= a and not b;
    layer3_outputs(1107) <= not a;
    layer3_outputs(1108) <= a;
    layer3_outputs(1109) <= not (a or b);
    layer3_outputs(1110) <= not b;
    layer3_outputs(1111) <= b;
    layer3_outputs(1112) <= a and b;
    layer3_outputs(1113) <= b and not a;
    layer3_outputs(1114) <= not b;
    layer3_outputs(1115) <= a or b;
    layer3_outputs(1116) <= a and not b;
    layer3_outputs(1117) <= not b;
    layer3_outputs(1118) <= a;
    layer3_outputs(1119) <= not b;
    layer3_outputs(1120) <= not a or b;
    layer3_outputs(1121) <= not (a or b);
    layer3_outputs(1122) <= a xor b;
    layer3_outputs(1123) <= a or b;
    layer3_outputs(1124) <= not (a and b);
    layer3_outputs(1125) <= not b or a;
    layer3_outputs(1126) <= not b;
    layer3_outputs(1127) <= a or b;
    layer3_outputs(1128) <= a;
    layer3_outputs(1129) <= a or b;
    layer3_outputs(1130) <= not a or b;
    layer3_outputs(1131) <= not b;
    layer3_outputs(1132) <= not b;
    layer3_outputs(1133) <= not b;
    layer3_outputs(1134) <= not b or a;
    layer3_outputs(1135) <= b;
    layer3_outputs(1136) <= not (a xor b);
    layer3_outputs(1137) <= not a or b;
    layer3_outputs(1138) <= not (a or b);
    layer3_outputs(1139) <= a and not b;
    layer3_outputs(1140) <= not a;
    layer3_outputs(1141) <= not b or a;
    layer3_outputs(1142) <= b;
    layer3_outputs(1143) <= a;
    layer3_outputs(1144) <= not (a xor b);
    layer3_outputs(1145) <= a;
    layer3_outputs(1146) <= not b;
    layer3_outputs(1147) <= not a;
    layer3_outputs(1148) <= not (a and b);
    layer3_outputs(1149) <= not b or a;
    layer3_outputs(1150) <= b;
    layer3_outputs(1151) <= a and b;
    layer3_outputs(1152) <= not b or a;
    layer3_outputs(1153) <= not a;
    layer3_outputs(1154) <= not (a xor b);
    layer3_outputs(1155) <= a and b;
    layer3_outputs(1156) <= not a;
    layer3_outputs(1157) <= a or b;
    layer3_outputs(1158) <= b and not a;
    layer3_outputs(1159) <= not (a xor b);
    layer3_outputs(1160) <= a and b;
    layer3_outputs(1161) <= not (a or b);
    layer3_outputs(1162) <= a;
    layer3_outputs(1163) <= not b;
    layer3_outputs(1164) <= a;
    layer3_outputs(1165) <= not b;
    layer3_outputs(1166) <= b;
    layer3_outputs(1167) <= a and not b;
    layer3_outputs(1168) <= not b;
    layer3_outputs(1169) <= not a or b;
    layer3_outputs(1170) <= b;
    layer3_outputs(1171) <= not a or b;
    layer3_outputs(1172) <= b;
    layer3_outputs(1173) <= a or b;
    layer3_outputs(1174) <= a xor b;
    layer3_outputs(1175) <= not (a or b);
    layer3_outputs(1176) <= not b or a;
    layer3_outputs(1177) <= not (a and b);
    layer3_outputs(1178) <= not (a and b);
    layer3_outputs(1179) <= not (a and b);
    layer3_outputs(1180) <= not a or b;
    layer3_outputs(1181) <= a or b;
    layer3_outputs(1182) <= not b or a;
    layer3_outputs(1183) <= '0';
    layer3_outputs(1184) <= a or b;
    layer3_outputs(1185) <= not b or a;
    layer3_outputs(1186) <= not (a and b);
    layer3_outputs(1187) <= not b;
    layer3_outputs(1188) <= a xor b;
    layer3_outputs(1189) <= not (a and b);
    layer3_outputs(1190) <= not a;
    layer3_outputs(1191) <= not b;
    layer3_outputs(1192) <= not (a and b);
    layer3_outputs(1193) <= not b;
    layer3_outputs(1194) <= not b or a;
    layer3_outputs(1195) <= a and not b;
    layer3_outputs(1196) <= a and b;
    layer3_outputs(1197) <= '0';
    layer3_outputs(1198) <= a and b;
    layer3_outputs(1199) <= not b;
    layer3_outputs(1200) <= a xor b;
    layer3_outputs(1201) <= not (a xor b);
    layer3_outputs(1202) <= a;
    layer3_outputs(1203) <= a or b;
    layer3_outputs(1204) <= not a;
    layer3_outputs(1205) <= not a;
    layer3_outputs(1206) <= b;
    layer3_outputs(1207) <= a and not b;
    layer3_outputs(1208) <= not a or b;
    layer3_outputs(1209) <= not a or b;
    layer3_outputs(1210) <= not (a and b);
    layer3_outputs(1211) <= not a or b;
    layer3_outputs(1212) <= not (a and b);
    layer3_outputs(1213) <= not b or a;
    layer3_outputs(1214) <= not b;
    layer3_outputs(1215) <= not a;
    layer3_outputs(1216) <= a;
    layer3_outputs(1217) <= not b;
    layer3_outputs(1218) <= not (a xor b);
    layer3_outputs(1219) <= a xor b;
    layer3_outputs(1220) <= not (a or b);
    layer3_outputs(1221) <= a;
    layer3_outputs(1222) <= a and not b;
    layer3_outputs(1223) <= b and not a;
    layer3_outputs(1224) <= not (a xor b);
    layer3_outputs(1225) <= a;
    layer3_outputs(1226) <= not a;
    layer3_outputs(1227) <= b and not a;
    layer3_outputs(1228) <= a and b;
    layer3_outputs(1229) <= a;
    layer3_outputs(1230) <= b and not a;
    layer3_outputs(1231) <= not a;
    layer3_outputs(1232) <= a;
    layer3_outputs(1233) <= a and not b;
    layer3_outputs(1234) <= a or b;
    layer3_outputs(1235) <= not (a and b);
    layer3_outputs(1236) <= not (a or b);
    layer3_outputs(1237) <= a and b;
    layer3_outputs(1238) <= not a or b;
    layer3_outputs(1239) <= not a or b;
    layer3_outputs(1240) <= not b or a;
    layer3_outputs(1241) <= not a or b;
    layer3_outputs(1242) <= a xor b;
    layer3_outputs(1243) <= not b or a;
    layer3_outputs(1244) <= not b;
    layer3_outputs(1245) <= b;
    layer3_outputs(1246) <= not a;
    layer3_outputs(1247) <= not b;
    layer3_outputs(1248) <= a;
    layer3_outputs(1249) <= not (a xor b);
    layer3_outputs(1250) <= b and not a;
    layer3_outputs(1251) <= not a or b;
    layer3_outputs(1252) <= not (a xor b);
    layer3_outputs(1253) <= not (a or b);
    layer3_outputs(1254) <= b and not a;
    layer3_outputs(1255) <= a or b;
    layer3_outputs(1256) <= a and b;
    layer3_outputs(1257) <= a;
    layer3_outputs(1258) <= a;
    layer3_outputs(1259) <= b and not a;
    layer3_outputs(1260) <= b;
    layer3_outputs(1261) <= not b;
    layer3_outputs(1262) <= b and not a;
    layer3_outputs(1263) <= a xor b;
    layer3_outputs(1264) <= b;
    layer3_outputs(1265) <= a or b;
    layer3_outputs(1266) <= a;
    layer3_outputs(1267) <= not (a and b);
    layer3_outputs(1268) <= b;
    layer3_outputs(1269) <= not a;
    layer3_outputs(1270) <= a;
    layer3_outputs(1271) <= not b;
    layer3_outputs(1272) <= a;
    layer3_outputs(1273) <= a or b;
    layer3_outputs(1274) <= a xor b;
    layer3_outputs(1275) <= not (a or b);
    layer3_outputs(1276) <= not a;
    layer3_outputs(1277) <= not a;
    layer3_outputs(1278) <= '0';
    layer3_outputs(1279) <= not b or a;
    layer3_outputs(1280) <= a xor b;
    layer3_outputs(1281) <= not b;
    layer3_outputs(1282) <= '0';
    layer3_outputs(1283) <= not b or a;
    layer3_outputs(1284) <= not b or a;
    layer3_outputs(1285) <= not b;
    layer3_outputs(1286) <= not a;
    layer3_outputs(1287) <= a xor b;
    layer3_outputs(1288) <= a;
    layer3_outputs(1289) <= not (a or b);
    layer3_outputs(1290) <= a and b;
    layer3_outputs(1291) <= a;
    layer3_outputs(1292) <= b and not a;
    layer3_outputs(1293) <= not b;
    layer3_outputs(1294) <= a and b;
    layer3_outputs(1295) <= not b or a;
    layer3_outputs(1296) <= not b;
    layer3_outputs(1297) <= a;
    layer3_outputs(1298) <= not a;
    layer3_outputs(1299) <= b and not a;
    layer3_outputs(1300) <= not a;
    layer3_outputs(1301) <= not a;
    layer3_outputs(1302) <= not b or a;
    layer3_outputs(1303) <= not (a and b);
    layer3_outputs(1304) <= b;
    layer3_outputs(1305) <= not (a xor b);
    layer3_outputs(1306) <= a and not b;
    layer3_outputs(1307) <= a and not b;
    layer3_outputs(1308) <= not (a xor b);
    layer3_outputs(1309) <= b and not a;
    layer3_outputs(1310) <= a and b;
    layer3_outputs(1311) <= a or b;
    layer3_outputs(1312) <= not (a xor b);
    layer3_outputs(1313) <= not b or a;
    layer3_outputs(1314) <= not b;
    layer3_outputs(1315) <= a and not b;
    layer3_outputs(1316) <= not a;
    layer3_outputs(1317) <= a xor b;
    layer3_outputs(1318) <= not a;
    layer3_outputs(1319) <= b;
    layer3_outputs(1320) <= not a;
    layer3_outputs(1321) <= a;
    layer3_outputs(1322) <= a and b;
    layer3_outputs(1323) <= not (a and b);
    layer3_outputs(1324) <= not (a or b);
    layer3_outputs(1325) <= a or b;
    layer3_outputs(1326) <= not a or b;
    layer3_outputs(1327) <= not a;
    layer3_outputs(1328) <= '1';
    layer3_outputs(1329) <= a xor b;
    layer3_outputs(1330) <= not a;
    layer3_outputs(1331) <= not b or a;
    layer3_outputs(1332) <= a and b;
    layer3_outputs(1333) <= b and not a;
    layer3_outputs(1334) <= a or b;
    layer3_outputs(1335) <= a;
    layer3_outputs(1336) <= a;
    layer3_outputs(1337) <= b and not a;
    layer3_outputs(1338) <= not (a and b);
    layer3_outputs(1339) <= a and b;
    layer3_outputs(1340) <= not a or b;
    layer3_outputs(1341) <= b and not a;
    layer3_outputs(1342) <= not (a and b);
    layer3_outputs(1343) <= '1';
    layer3_outputs(1344) <= not (a and b);
    layer3_outputs(1345) <= a or b;
    layer3_outputs(1346) <= a and not b;
    layer3_outputs(1347) <= not a;
    layer3_outputs(1348) <= b and not a;
    layer3_outputs(1349) <= b;
    layer3_outputs(1350) <= a or b;
    layer3_outputs(1351) <= b;
    layer3_outputs(1352) <= a or b;
    layer3_outputs(1353) <= not (a or b);
    layer3_outputs(1354) <= a and not b;
    layer3_outputs(1355) <= not (a or b);
    layer3_outputs(1356) <= not b;
    layer3_outputs(1357) <= not (a xor b);
    layer3_outputs(1358) <= b;
    layer3_outputs(1359) <= a or b;
    layer3_outputs(1360) <= not (a and b);
    layer3_outputs(1361) <= not a;
    layer3_outputs(1362) <= a and b;
    layer3_outputs(1363) <= b and not a;
    layer3_outputs(1364) <= not (a and b);
    layer3_outputs(1365) <= not (a and b);
    layer3_outputs(1366) <= a;
    layer3_outputs(1367) <= not (a xor b);
    layer3_outputs(1368) <= not (a and b);
    layer3_outputs(1369) <= not a or b;
    layer3_outputs(1370) <= b;
    layer3_outputs(1371) <= a;
    layer3_outputs(1372) <= not a;
    layer3_outputs(1373) <= not b or a;
    layer3_outputs(1374) <= '0';
    layer3_outputs(1375) <= not (a and b);
    layer3_outputs(1376) <= a and not b;
    layer3_outputs(1377) <= b;
    layer3_outputs(1378) <= a;
    layer3_outputs(1379) <= not b or a;
    layer3_outputs(1380) <= not a;
    layer3_outputs(1381) <= not (a or b);
    layer3_outputs(1382) <= b;
    layer3_outputs(1383) <= not b;
    layer3_outputs(1384) <= not (a xor b);
    layer3_outputs(1385) <= not b;
    layer3_outputs(1386) <= not (a or b);
    layer3_outputs(1387) <= not (a and b);
    layer3_outputs(1388) <= b and not a;
    layer3_outputs(1389) <= not b;
    layer3_outputs(1390) <= a and b;
    layer3_outputs(1391) <= not (a and b);
    layer3_outputs(1392) <= not (a xor b);
    layer3_outputs(1393) <= a and not b;
    layer3_outputs(1394) <= not a;
    layer3_outputs(1395) <= a;
    layer3_outputs(1396) <= a;
    layer3_outputs(1397) <= b;
    layer3_outputs(1398) <= not b;
    layer3_outputs(1399) <= not (a or b);
    layer3_outputs(1400) <= a;
    layer3_outputs(1401) <= a;
    layer3_outputs(1402) <= not a;
    layer3_outputs(1403) <= b;
    layer3_outputs(1404) <= not a;
    layer3_outputs(1405) <= b and not a;
    layer3_outputs(1406) <= not a;
    layer3_outputs(1407) <= not (a and b);
    layer3_outputs(1408) <= not a or b;
    layer3_outputs(1409) <= not (a or b);
    layer3_outputs(1410) <= a;
    layer3_outputs(1411) <= not a;
    layer3_outputs(1412) <= not a or b;
    layer3_outputs(1413) <= a and b;
    layer3_outputs(1414) <= b;
    layer3_outputs(1415) <= a and not b;
    layer3_outputs(1416) <= '1';
    layer3_outputs(1417) <= not a or b;
    layer3_outputs(1418) <= a;
    layer3_outputs(1419) <= not b;
    layer3_outputs(1420) <= b;
    layer3_outputs(1421) <= not a;
    layer3_outputs(1422) <= not a;
    layer3_outputs(1423) <= not b;
    layer3_outputs(1424) <= not (a and b);
    layer3_outputs(1425) <= not a;
    layer3_outputs(1426) <= a;
    layer3_outputs(1427) <= b;
    layer3_outputs(1428) <= a and b;
    layer3_outputs(1429) <= a;
    layer3_outputs(1430) <= not (a xor b);
    layer3_outputs(1431) <= a and b;
    layer3_outputs(1432) <= not a or b;
    layer3_outputs(1433) <= a xor b;
    layer3_outputs(1434) <= b;
    layer3_outputs(1435) <= not (a xor b);
    layer3_outputs(1436) <= not a;
    layer3_outputs(1437) <= a;
    layer3_outputs(1438) <= not a;
    layer3_outputs(1439) <= b and not a;
    layer3_outputs(1440) <= b and not a;
    layer3_outputs(1441) <= b and not a;
    layer3_outputs(1442) <= not b or a;
    layer3_outputs(1443) <= '1';
    layer3_outputs(1444) <= not a;
    layer3_outputs(1445) <= a and not b;
    layer3_outputs(1446) <= not a or b;
    layer3_outputs(1447) <= a;
    layer3_outputs(1448) <= a and b;
    layer3_outputs(1449) <= not b;
    layer3_outputs(1450) <= not a;
    layer3_outputs(1451) <= not b;
    layer3_outputs(1452) <= not (a and b);
    layer3_outputs(1453) <= not (a and b);
    layer3_outputs(1454) <= not (a and b);
    layer3_outputs(1455) <= not b or a;
    layer3_outputs(1456) <= not (a or b);
    layer3_outputs(1457) <= not a or b;
    layer3_outputs(1458) <= not b or a;
    layer3_outputs(1459) <= a or b;
    layer3_outputs(1460) <= '0';
    layer3_outputs(1461) <= a and b;
    layer3_outputs(1462) <= not b or a;
    layer3_outputs(1463) <= not b;
    layer3_outputs(1464) <= '0';
    layer3_outputs(1465) <= a;
    layer3_outputs(1466) <= a and not b;
    layer3_outputs(1467) <= b and not a;
    layer3_outputs(1468) <= not b;
    layer3_outputs(1469) <= not b;
    layer3_outputs(1470) <= not (a or b);
    layer3_outputs(1471) <= b;
    layer3_outputs(1472) <= not (a and b);
    layer3_outputs(1473) <= b and not a;
    layer3_outputs(1474) <= not (a and b);
    layer3_outputs(1475) <= not a or b;
    layer3_outputs(1476) <= not b;
    layer3_outputs(1477) <= a or b;
    layer3_outputs(1478) <= not a;
    layer3_outputs(1479) <= a or b;
    layer3_outputs(1480) <= not a;
    layer3_outputs(1481) <= a;
    layer3_outputs(1482) <= not a;
    layer3_outputs(1483) <= a xor b;
    layer3_outputs(1484) <= a and b;
    layer3_outputs(1485) <= not a;
    layer3_outputs(1486) <= not b;
    layer3_outputs(1487) <= a xor b;
    layer3_outputs(1488) <= a and not b;
    layer3_outputs(1489) <= a;
    layer3_outputs(1490) <= not (a or b);
    layer3_outputs(1491) <= not b or a;
    layer3_outputs(1492) <= a and b;
    layer3_outputs(1493) <= b;
    layer3_outputs(1494) <= not b or a;
    layer3_outputs(1495) <= not a or b;
    layer3_outputs(1496) <= b;
    layer3_outputs(1497) <= a and b;
    layer3_outputs(1498) <= not (a or b);
    layer3_outputs(1499) <= not a or b;
    layer3_outputs(1500) <= b and not a;
    layer3_outputs(1501) <= b and not a;
    layer3_outputs(1502) <= b;
    layer3_outputs(1503) <= a;
    layer3_outputs(1504) <= not b;
    layer3_outputs(1505) <= not (a and b);
    layer3_outputs(1506) <= a;
    layer3_outputs(1507) <= not b;
    layer3_outputs(1508) <= a and b;
    layer3_outputs(1509) <= not b;
    layer3_outputs(1510) <= not (a and b);
    layer3_outputs(1511) <= b;
    layer3_outputs(1512) <= b and not a;
    layer3_outputs(1513) <= not (a or b);
    layer3_outputs(1514) <= a and not b;
    layer3_outputs(1515) <= not (a and b);
    layer3_outputs(1516) <= '0';
    layer3_outputs(1517) <= a and not b;
    layer3_outputs(1518) <= not b;
    layer3_outputs(1519) <= not (a xor b);
    layer3_outputs(1520) <= not (a or b);
    layer3_outputs(1521) <= not b or a;
    layer3_outputs(1522) <= not a;
    layer3_outputs(1523) <= not a or b;
    layer3_outputs(1524) <= b and not a;
    layer3_outputs(1525) <= not (a or b);
    layer3_outputs(1526) <= a;
    layer3_outputs(1527) <= not a or b;
    layer3_outputs(1528) <= b and not a;
    layer3_outputs(1529) <= a and b;
    layer3_outputs(1530) <= b and not a;
    layer3_outputs(1531) <= b;
    layer3_outputs(1532) <= b;
    layer3_outputs(1533) <= a xor b;
    layer3_outputs(1534) <= not a or b;
    layer3_outputs(1535) <= not (a xor b);
    layer3_outputs(1536) <= a and b;
    layer3_outputs(1537) <= not (a xor b);
    layer3_outputs(1538) <= not b or a;
    layer3_outputs(1539) <= not (a xor b);
    layer3_outputs(1540) <= a and b;
    layer3_outputs(1541) <= not (a or b);
    layer3_outputs(1542) <= not (a xor b);
    layer3_outputs(1543) <= a;
    layer3_outputs(1544) <= not a or b;
    layer3_outputs(1545) <= a and not b;
    layer3_outputs(1546) <= not a or b;
    layer3_outputs(1547) <= b;
    layer3_outputs(1548) <= not b;
    layer3_outputs(1549) <= a;
    layer3_outputs(1550) <= b and not a;
    layer3_outputs(1551) <= not b;
    layer3_outputs(1552) <= a;
    layer3_outputs(1553) <= b;
    layer3_outputs(1554) <= not b;
    layer3_outputs(1555) <= not (a xor b);
    layer3_outputs(1556) <= not a;
    layer3_outputs(1557) <= b;
    layer3_outputs(1558) <= a and b;
    layer3_outputs(1559) <= a;
    layer3_outputs(1560) <= not (a or b);
    layer3_outputs(1561) <= not (a xor b);
    layer3_outputs(1562) <= not b or a;
    layer3_outputs(1563) <= a or b;
    layer3_outputs(1564) <= not a;
    layer3_outputs(1565) <= not b;
    layer3_outputs(1566) <= not (a and b);
    layer3_outputs(1567) <= not a or b;
    layer3_outputs(1568) <= a;
    layer3_outputs(1569) <= b;
    layer3_outputs(1570) <= b;
    layer3_outputs(1571) <= not (a and b);
    layer3_outputs(1572) <= b and not a;
    layer3_outputs(1573) <= b;
    layer3_outputs(1574) <= a;
    layer3_outputs(1575) <= a or b;
    layer3_outputs(1576) <= a xor b;
    layer3_outputs(1577) <= not a or b;
    layer3_outputs(1578) <= a and b;
    layer3_outputs(1579) <= not b or a;
    layer3_outputs(1580) <= a and not b;
    layer3_outputs(1581) <= b;
    layer3_outputs(1582) <= a xor b;
    layer3_outputs(1583) <= not (a and b);
    layer3_outputs(1584) <= not b;
    layer3_outputs(1585) <= a;
    layer3_outputs(1586) <= a;
    layer3_outputs(1587) <= b;
    layer3_outputs(1588) <= not a or b;
    layer3_outputs(1589) <= b;
    layer3_outputs(1590) <= not (a or b);
    layer3_outputs(1591) <= a xor b;
    layer3_outputs(1592) <= not a;
    layer3_outputs(1593) <= not a or b;
    layer3_outputs(1594) <= '1';
    layer3_outputs(1595) <= b;
    layer3_outputs(1596) <= not a;
    layer3_outputs(1597) <= not a;
    layer3_outputs(1598) <= not (a xor b);
    layer3_outputs(1599) <= b;
    layer3_outputs(1600) <= not b;
    layer3_outputs(1601) <= not a or b;
    layer3_outputs(1602) <= a and not b;
    layer3_outputs(1603) <= a xor b;
    layer3_outputs(1604) <= a;
    layer3_outputs(1605) <= not a;
    layer3_outputs(1606) <= a and b;
    layer3_outputs(1607) <= not b or a;
    layer3_outputs(1608) <= a or b;
    layer3_outputs(1609) <= '1';
    layer3_outputs(1610) <= not (a or b);
    layer3_outputs(1611) <= not (a or b);
    layer3_outputs(1612) <= a or b;
    layer3_outputs(1613) <= not b;
    layer3_outputs(1614) <= b and not a;
    layer3_outputs(1615) <= not (a xor b);
    layer3_outputs(1616) <= a;
    layer3_outputs(1617) <= not (a or b);
    layer3_outputs(1618) <= not b;
    layer3_outputs(1619) <= not (a and b);
    layer3_outputs(1620) <= b;
    layer3_outputs(1621) <= b and not a;
    layer3_outputs(1622) <= b;
    layer3_outputs(1623) <= a and b;
    layer3_outputs(1624) <= a and b;
    layer3_outputs(1625) <= b and not a;
    layer3_outputs(1626) <= not b;
    layer3_outputs(1627) <= not b or a;
    layer3_outputs(1628) <= not (a and b);
    layer3_outputs(1629) <= a xor b;
    layer3_outputs(1630) <= b;
    layer3_outputs(1631) <= not a;
    layer3_outputs(1632) <= not b;
    layer3_outputs(1633) <= a and not b;
    layer3_outputs(1634) <= a;
    layer3_outputs(1635) <= not (a or b);
    layer3_outputs(1636) <= b;
    layer3_outputs(1637) <= not a;
    layer3_outputs(1638) <= a xor b;
    layer3_outputs(1639) <= not b;
    layer3_outputs(1640) <= b;
    layer3_outputs(1641) <= not (a xor b);
    layer3_outputs(1642) <= not b or a;
    layer3_outputs(1643) <= b;
    layer3_outputs(1644) <= not (a xor b);
    layer3_outputs(1645) <= a or b;
    layer3_outputs(1646) <= a xor b;
    layer3_outputs(1647) <= b and not a;
    layer3_outputs(1648) <= not (a or b);
    layer3_outputs(1649) <= b;
    layer3_outputs(1650) <= not a;
    layer3_outputs(1651) <= b and not a;
    layer3_outputs(1652) <= not a;
    layer3_outputs(1653) <= b;
    layer3_outputs(1654) <= not b;
    layer3_outputs(1655) <= a and b;
    layer3_outputs(1656) <= b;
    layer3_outputs(1657) <= a or b;
    layer3_outputs(1658) <= not (a or b);
    layer3_outputs(1659) <= not a;
    layer3_outputs(1660) <= not (a xor b);
    layer3_outputs(1661) <= not (a and b);
    layer3_outputs(1662) <= not b;
    layer3_outputs(1663) <= b;
    layer3_outputs(1664) <= not (a and b);
    layer3_outputs(1665) <= b and not a;
    layer3_outputs(1666) <= not a;
    layer3_outputs(1667) <= not (a and b);
    layer3_outputs(1668) <= not (a and b);
    layer3_outputs(1669) <= a or b;
    layer3_outputs(1670) <= not (a and b);
    layer3_outputs(1671) <= a and not b;
    layer3_outputs(1672) <= not b;
    layer3_outputs(1673) <= a xor b;
    layer3_outputs(1674) <= b;
    layer3_outputs(1675) <= '1';
    layer3_outputs(1676) <= a or b;
    layer3_outputs(1677) <= not (a or b);
    layer3_outputs(1678) <= a;
    layer3_outputs(1679) <= a or b;
    layer3_outputs(1680) <= not a;
    layer3_outputs(1681) <= a;
    layer3_outputs(1682) <= b;
    layer3_outputs(1683) <= not a or b;
    layer3_outputs(1684) <= b and not a;
    layer3_outputs(1685) <= a and b;
    layer3_outputs(1686) <= a and b;
    layer3_outputs(1687) <= not a;
    layer3_outputs(1688) <= a xor b;
    layer3_outputs(1689) <= b;
    layer3_outputs(1690) <= not (a or b);
    layer3_outputs(1691) <= b;
    layer3_outputs(1692) <= not (a and b);
    layer3_outputs(1693) <= not b or a;
    layer3_outputs(1694) <= a xor b;
    layer3_outputs(1695) <= not (a or b);
    layer3_outputs(1696) <= not a or b;
    layer3_outputs(1697) <= not b;
    layer3_outputs(1698) <= not (a and b);
    layer3_outputs(1699) <= a or b;
    layer3_outputs(1700) <= a;
    layer3_outputs(1701) <= not b;
    layer3_outputs(1702) <= not b;
    layer3_outputs(1703) <= not a;
    layer3_outputs(1704) <= not b;
    layer3_outputs(1705) <= not a;
    layer3_outputs(1706) <= not a;
    layer3_outputs(1707) <= not b or a;
    layer3_outputs(1708) <= not b;
    layer3_outputs(1709) <= a and b;
    layer3_outputs(1710) <= a xor b;
    layer3_outputs(1711) <= not a or b;
    layer3_outputs(1712) <= not (a and b);
    layer3_outputs(1713) <= not (a or b);
    layer3_outputs(1714) <= not a or b;
    layer3_outputs(1715) <= a or b;
    layer3_outputs(1716) <= b;
    layer3_outputs(1717) <= a;
    layer3_outputs(1718) <= not b or a;
    layer3_outputs(1719) <= b;
    layer3_outputs(1720) <= b;
    layer3_outputs(1721) <= a;
    layer3_outputs(1722) <= not b;
    layer3_outputs(1723) <= not a or b;
    layer3_outputs(1724) <= not (a and b);
    layer3_outputs(1725) <= b and not a;
    layer3_outputs(1726) <= '1';
    layer3_outputs(1727) <= b and not a;
    layer3_outputs(1728) <= a and not b;
    layer3_outputs(1729) <= not (a and b);
    layer3_outputs(1730) <= a and b;
    layer3_outputs(1731) <= not b or a;
    layer3_outputs(1732) <= not b or a;
    layer3_outputs(1733) <= a or b;
    layer3_outputs(1734) <= not a;
    layer3_outputs(1735) <= a;
    layer3_outputs(1736) <= b and not a;
    layer3_outputs(1737) <= b;
    layer3_outputs(1738) <= a or b;
    layer3_outputs(1739) <= not b or a;
    layer3_outputs(1740) <= not (a and b);
    layer3_outputs(1741) <= a xor b;
    layer3_outputs(1742) <= not a;
    layer3_outputs(1743) <= b;
    layer3_outputs(1744) <= a xor b;
    layer3_outputs(1745) <= b;
    layer3_outputs(1746) <= not b;
    layer3_outputs(1747) <= b;
    layer3_outputs(1748) <= a or b;
    layer3_outputs(1749) <= not (a or b);
    layer3_outputs(1750) <= a xor b;
    layer3_outputs(1751) <= b;
    layer3_outputs(1752) <= not (a xor b);
    layer3_outputs(1753) <= not a;
    layer3_outputs(1754) <= b and not a;
    layer3_outputs(1755) <= '0';
    layer3_outputs(1756) <= not (a or b);
    layer3_outputs(1757) <= not b;
    layer3_outputs(1758) <= a and not b;
    layer3_outputs(1759) <= a and not b;
    layer3_outputs(1760) <= a xor b;
    layer3_outputs(1761) <= a;
    layer3_outputs(1762) <= not a or b;
    layer3_outputs(1763) <= not a or b;
    layer3_outputs(1764) <= a or b;
    layer3_outputs(1765) <= a xor b;
    layer3_outputs(1766) <= a and not b;
    layer3_outputs(1767) <= a and b;
    layer3_outputs(1768) <= not b;
    layer3_outputs(1769) <= a;
    layer3_outputs(1770) <= b;
    layer3_outputs(1771) <= '1';
    layer3_outputs(1772) <= not a;
    layer3_outputs(1773) <= '1';
    layer3_outputs(1774) <= not a or b;
    layer3_outputs(1775) <= not a;
    layer3_outputs(1776) <= not a or b;
    layer3_outputs(1777) <= b;
    layer3_outputs(1778) <= b;
    layer3_outputs(1779) <= a and b;
    layer3_outputs(1780) <= not a;
    layer3_outputs(1781) <= b;
    layer3_outputs(1782) <= b and not a;
    layer3_outputs(1783) <= not (a or b);
    layer3_outputs(1784) <= a;
    layer3_outputs(1785) <= b;
    layer3_outputs(1786) <= not b or a;
    layer3_outputs(1787) <= not b;
    layer3_outputs(1788) <= not a;
    layer3_outputs(1789) <= a;
    layer3_outputs(1790) <= b and not a;
    layer3_outputs(1791) <= '1';
    layer3_outputs(1792) <= not (a or b);
    layer3_outputs(1793) <= not (a or b);
    layer3_outputs(1794) <= not (a or b);
    layer3_outputs(1795) <= not b;
    layer3_outputs(1796) <= a;
    layer3_outputs(1797) <= a xor b;
    layer3_outputs(1798) <= not a or b;
    layer3_outputs(1799) <= not a;
    layer3_outputs(1800) <= not (a or b);
    layer3_outputs(1801) <= b;
    layer3_outputs(1802) <= not (a xor b);
    layer3_outputs(1803) <= not (a or b);
    layer3_outputs(1804) <= not b;
    layer3_outputs(1805) <= a;
    layer3_outputs(1806) <= not b;
    layer3_outputs(1807) <= a or b;
    layer3_outputs(1808) <= not a;
    layer3_outputs(1809) <= not b or a;
    layer3_outputs(1810) <= '1';
    layer3_outputs(1811) <= not b or a;
    layer3_outputs(1812) <= not a;
    layer3_outputs(1813) <= not b;
    layer3_outputs(1814) <= b;
    layer3_outputs(1815) <= '0';
    layer3_outputs(1816) <= a xor b;
    layer3_outputs(1817) <= a and not b;
    layer3_outputs(1818) <= b;
    layer3_outputs(1819) <= b;
    layer3_outputs(1820) <= a;
    layer3_outputs(1821) <= b;
    layer3_outputs(1822) <= not b or a;
    layer3_outputs(1823) <= a or b;
    layer3_outputs(1824) <= a xor b;
    layer3_outputs(1825) <= b and not a;
    layer3_outputs(1826) <= b;
    layer3_outputs(1827) <= a;
    layer3_outputs(1828) <= '1';
    layer3_outputs(1829) <= not a;
    layer3_outputs(1830) <= a or b;
    layer3_outputs(1831) <= not (a or b);
    layer3_outputs(1832) <= a and b;
    layer3_outputs(1833) <= a;
    layer3_outputs(1834) <= not (a and b);
    layer3_outputs(1835) <= not a;
    layer3_outputs(1836) <= a and not b;
    layer3_outputs(1837) <= '0';
    layer3_outputs(1838) <= '0';
    layer3_outputs(1839) <= a;
    layer3_outputs(1840) <= not b or a;
    layer3_outputs(1841) <= a or b;
    layer3_outputs(1842) <= '1';
    layer3_outputs(1843) <= b and not a;
    layer3_outputs(1844) <= not (a and b);
    layer3_outputs(1845) <= a and not b;
    layer3_outputs(1846) <= a and not b;
    layer3_outputs(1847) <= not a or b;
    layer3_outputs(1848) <= not b or a;
    layer3_outputs(1849) <= a xor b;
    layer3_outputs(1850) <= a or b;
    layer3_outputs(1851) <= not a or b;
    layer3_outputs(1852) <= not (a xor b);
    layer3_outputs(1853) <= b;
    layer3_outputs(1854) <= not b or a;
    layer3_outputs(1855) <= not a;
    layer3_outputs(1856) <= not (a xor b);
    layer3_outputs(1857) <= a;
    layer3_outputs(1858) <= a;
    layer3_outputs(1859) <= a or b;
    layer3_outputs(1860) <= not b or a;
    layer3_outputs(1861) <= a;
    layer3_outputs(1862) <= a;
    layer3_outputs(1863) <= b;
    layer3_outputs(1864) <= not (a and b);
    layer3_outputs(1865) <= '1';
    layer3_outputs(1866) <= not b or a;
    layer3_outputs(1867) <= not a or b;
    layer3_outputs(1868) <= not (a and b);
    layer3_outputs(1869) <= '1';
    layer3_outputs(1870) <= not b or a;
    layer3_outputs(1871) <= not a or b;
    layer3_outputs(1872) <= b;
    layer3_outputs(1873) <= a or b;
    layer3_outputs(1874) <= a or b;
    layer3_outputs(1875) <= a and not b;
    layer3_outputs(1876) <= a and not b;
    layer3_outputs(1877) <= not a;
    layer3_outputs(1878) <= not a or b;
    layer3_outputs(1879) <= not b;
    layer3_outputs(1880) <= not a or b;
    layer3_outputs(1881) <= not (a xor b);
    layer3_outputs(1882) <= a and not b;
    layer3_outputs(1883) <= not (a and b);
    layer3_outputs(1884) <= a and not b;
    layer3_outputs(1885) <= a;
    layer3_outputs(1886) <= not a;
    layer3_outputs(1887) <= a;
    layer3_outputs(1888) <= a or b;
    layer3_outputs(1889) <= not b;
    layer3_outputs(1890) <= b;
    layer3_outputs(1891) <= not a or b;
    layer3_outputs(1892) <= a or b;
    layer3_outputs(1893) <= a;
    layer3_outputs(1894) <= not (a xor b);
    layer3_outputs(1895) <= not b;
    layer3_outputs(1896) <= not a or b;
    layer3_outputs(1897) <= not b or a;
    layer3_outputs(1898) <= b;
    layer3_outputs(1899) <= '0';
    layer3_outputs(1900) <= a;
    layer3_outputs(1901) <= a and b;
    layer3_outputs(1902) <= not b;
    layer3_outputs(1903) <= a;
    layer3_outputs(1904) <= not a or b;
    layer3_outputs(1905) <= not a;
    layer3_outputs(1906) <= a;
    layer3_outputs(1907) <= a and not b;
    layer3_outputs(1908) <= not a or b;
    layer3_outputs(1909) <= not (a xor b);
    layer3_outputs(1910) <= a and b;
    layer3_outputs(1911) <= a and not b;
    layer3_outputs(1912) <= a and b;
    layer3_outputs(1913) <= not a;
    layer3_outputs(1914) <= a;
    layer3_outputs(1915) <= a;
    layer3_outputs(1916) <= b and not a;
    layer3_outputs(1917) <= a and b;
    layer3_outputs(1918) <= b;
    layer3_outputs(1919) <= not a or b;
    layer3_outputs(1920) <= '1';
    layer3_outputs(1921) <= a and b;
    layer3_outputs(1922) <= not a or b;
    layer3_outputs(1923) <= not b;
    layer3_outputs(1924) <= not a;
    layer3_outputs(1925) <= not (a or b);
    layer3_outputs(1926) <= b and not a;
    layer3_outputs(1927) <= a or b;
    layer3_outputs(1928) <= a xor b;
    layer3_outputs(1929) <= not (a and b);
    layer3_outputs(1930) <= b;
    layer3_outputs(1931) <= not a;
    layer3_outputs(1932) <= not (a xor b);
    layer3_outputs(1933) <= not b;
    layer3_outputs(1934) <= a and b;
    layer3_outputs(1935) <= a;
    layer3_outputs(1936) <= a and b;
    layer3_outputs(1937) <= not (a xor b);
    layer3_outputs(1938) <= not a;
    layer3_outputs(1939) <= a and not b;
    layer3_outputs(1940) <= not b or a;
    layer3_outputs(1941) <= a xor b;
    layer3_outputs(1942) <= b;
    layer3_outputs(1943) <= not b;
    layer3_outputs(1944) <= a xor b;
    layer3_outputs(1945) <= a or b;
    layer3_outputs(1946) <= a and b;
    layer3_outputs(1947) <= not b or a;
    layer3_outputs(1948) <= not a;
    layer3_outputs(1949) <= a and b;
    layer3_outputs(1950) <= not b;
    layer3_outputs(1951) <= not (a xor b);
    layer3_outputs(1952) <= b;
    layer3_outputs(1953) <= not b or a;
    layer3_outputs(1954) <= not a;
    layer3_outputs(1955) <= a or b;
    layer3_outputs(1956) <= not a;
    layer3_outputs(1957) <= not b;
    layer3_outputs(1958) <= not (a or b);
    layer3_outputs(1959) <= a or b;
    layer3_outputs(1960) <= b and not a;
    layer3_outputs(1961) <= not a or b;
    layer3_outputs(1962) <= not a;
    layer3_outputs(1963) <= a or b;
    layer3_outputs(1964) <= not (a xor b);
    layer3_outputs(1965) <= not b or a;
    layer3_outputs(1966) <= not (a or b);
    layer3_outputs(1967) <= a or b;
    layer3_outputs(1968) <= a;
    layer3_outputs(1969) <= a or b;
    layer3_outputs(1970) <= not (a or b);
    layer3_outputs(1971) <= a;
    layer3_outputs(1972) <= a;
    layer3_outputs(1973) <= b and not a;
    layer3_outputs(1974) <= not a;
    layer3_outputs(1975) <= b;
    layer3_outputs(1976) <= not b or a;
    layer3_outputs(1977) <= not (a or b);
    layer3_outputs(1978) <= not a;
    layer3_outputs(1979) <= not a;
    layer3_outputs(1980) <= not a;
    layer3_outputs(1981) <= not (a or b);
    layer3_outputs(1982) <= b and not a;
    layer3_outputs(1983) <= not b or a;
    layer3_outputs(1984) <= b;
    layer3_outputs(1985) <= a or b;
    layer3_outputs(1986) <= not (a xor b);
    layer3_outputs(1987) <= a and not b;
    layer3_outputs(1988) <= not (a or b);
    layer3_outputs(1989) <= a and not b;
    layer3_outputs(1990) <= a and not b;
    layer3_outputs(1991) <= not b or a;
    layer3_outputs(1992) <= not b or a;
    layer3_outputs(1993) <= a xor b;
    layer3_outputs(1994) <= a;
    layer3_outputs(1995) <= a or b;
    layer3_outputs(1996) <= a or b;
    layer3_outputs(1997) <= not a or b;
    layer3_outputs(1998) <= a or b;
    layer3_outputs(1999) <= a;
    layer3_outputs(2000) <= a and not b;
    layer3_outputs(2001) <= not (a or b);
    layer3_outputs(2002) <= not b or a;
    layer3_outputs(2003) <= not b;
    layer3_outputs(2004) <= b;
    layer3_outputs(2005) <= a xor b;
    layer3_outputs(2006) <= b;
    layer3_outputs(2007) <= a;
    layer3_outputs(2008) <= not a;
    layer3_outputs(2009) <= b;
    layer3_outputs(2010) <= a xor b;
    layer3_outputs(2011) <= b and not a;
    layer3_outputs(2012) <= not a or b;
    layer3_outputs(2013) <= not (a and b);
    layer3_outputs(2014) <= not b;
    layer3_outputs(2015) <= not b or a;
    layer3_outputs(2016) <= a or b;
    layer3_outputs(2017) <= a;
    layer3_outputs(2018) <= b;
    layer3_outputs(2019) <= b and not a;
    layer3_outputs(2020) <= not a;
    layer3_outputs(2021) <= a;
    layer3_outputs(2022) <= not b;
    layer3_outputs(2023) <= a and b;
    layer3_outputs(2024) <= not (a and b);
    layer3_outputs(2025) <= not b;
    layer3_outputs(2026) <= not a or b;
    layer3_outputs(2027) <= a and not b;
    layer3_outputs(2028) <= b;
    layer3_outputs(2029) <= a or b;
    layer3_outputs(2030) <= not (a or b);
    layer3_outputs(2031) <= not a;
    layer3_outputs(2032) <= not (a or b);
    layer3_outputs(2033) <= not b;
    layer3_outputs(2034) <= not a or b;
    layer3_outputs(2035) <= a;
    layer3_outputs(2036) <= a or b;
    layer3_outputs(2037) <= not (a xor b);
    layer3_outputs(2038) <= not b;
    layer3_outputs(2039) <= not a or b;
    layer3_outputs(2040) <= not (a or b);
    layer3_outputs(2041) <= not b;
    layer3_outputs(2042) <= not b;
    layer3_outputs(2043) <= not a or b;
    layer3_outputs(2044) <= not b or a;
    layer3_outputs(2045) <= not a;
    layer3_outputs(2046) <= b;
    layer3_outputs(2047) <= b;
    layer3_outputs(2048) <= a;
    layer3_outputs(2049) <= not a;
    layer3_outputs(2050) <= not b or a;
    layer3_outputs(2051) <= not (a xor b);
    layer3_outputs(2052) <= not a;
    layer3_outputs(2053) <= not (a and b);
    layer3_outputs(2054) <= not (a xor b);
    layer3_outputs(2055) <= b;
    layer3_outputs(2056) <= b;
    layer3_outputs(2057) <= not b;
    layer3_outputs(2058) <= not b or a;
    layer3_outputs(2059) <= not a or b;
    layer3_outputs(2060) <= b and not a;
    layer3_outputs(2061) <= a;
    layer3_outputs(2062) <= b;
    layer3_outputs(2063) <= '0';
    layer3_outputs(2064) <= '1';
    layer3_outputs(2065) <= not (a or b);
    layer3_outputs(2066) <= a and b;
    layer3_outputs(2067) <= not (a or b);
    layer3_outputs(2068) <= a and not b;
    layer3_outputs(2069) <= b;
    layer3_outputs(2070) <= not b;
    layer3_outputs(2071) <= a and b;
    layer3_outputs(2072) <= not (a or b);
    layer3_outputs(2073) <= not (a or b);
    layer3_outputs(2074) <= not a;
    layer3_outputs(2075) <= not (a and b);
    layer3_outputs(2076) <= a and not b;
    layer3_outputs(2077) <= not b;
    layer3_outputs(2078) <= '0';
    layer3_outputs(2079) <= not (a and b);
    layer3_outputs(2080) <= b and not a;
    layer3_outputs(2081) <= not (a or b);
    layer3_outputs(2082) <= not b;
    layer3_outputs(2083) <= a and b;
    layer3_outputs(2084) <= b;
    layer3_outputs(2085) <= b;
    layer3_outputs(2086) <= a;
    layer3_outputs(2087) <= not (a xor b);
    layer3_outputs(2088) <= b and not a;
    layer3_outputs(2089) <= a;
    layer3_outputs(2090) <= not b;
    layer3_outputs(2091) <= not a;
    layer3_outputs(2092) <= a and b;
    layer3_outputs(2093) <= b;
    layer3_outputs(2094) <= b and not a;
    layer3_outputs(2095) <= not (a xor b);
    layer3_outputs(2096) <= not b;
    layer3_outputs(2097) <= b;
    layer3_outputs(2098) <= not b;
    layer3_outputs(2099) <= a xor b;
    layer3_outputs(2100) <= not b;
    layer3_outputs(2101) <= not (a and b);
    layer3_outputs(2102) <= b;
    layer3_outputs(2103) <= a xor b;
    layer3_outputs(2104) <= a xor b;
    layer3_outputs(2105) <= a;
    layer3_outputs(2106) <= not (a and b);
    layer3_outputs(2107) <= a and not b;
    layer3_outputs(2108) <= b;
    layer3_outputs(2109) <= b;
    layer3_outputs(2110) <= a or b;
    layer3_outputs(2111) <= not (a or b);
    layer3_outputs(2112) <= not a;
    layer3_outputs(2113) <= a;
    layer3_outputs(2114) <= not (a and b);
    layer3_outputs(2115) <= a xor b;
    layer3_outputs(2116) <= b and not a;
    layer3_outputs(2117) <= not b;
    layer3_outputs(2118) <= a xor b;
    layer3_outputs(2119) <= a and not b;
    layer3_outputs(2120) <= a or b;
    layer3_outputs(2121) <= b and not a;
    layer3_outputs(2122) <= not b;
    layer3_outputs(2123) <= not a or b;
    layer3_outputs(2124) <= a and not b;
    layer3_outputs(2125) <= not (a and b);
    layer3_outputs(2126) <= b;
    layer3_outputs(2127) <= not a or b;
    layer3_outputs(2128) <= not b or a;
    layer3_outputs(2129) <= not b;
    layer3_outputs(2130) <= '0';
    layer3_outputs(2131) <= not b;
    layer3_outputs(2132) <= not (a and b);
    layer3_outputs(2133) <= not a or b;
    layer3_outputs(2134) <= a xor b;
    layer3_outputs(2135) <= not a;
    layer3_outputs(2136) <= not a;
    layer3_outputs(2137) <= not b;
    layer3_outputs(2138) <= b;
    layer3_outputs(2139) <= not (a or b);
    layer3_outputs(2140) <= a;
    layer3_outputs(2141) <= b and not a;
    layer3_outputs(2142) <= a or b;
    layer3_outputs(2143) <= not b;
    layer3_outputs(2144) <= not (a or b);
    layer3_outputs(2145) <= not (a and b);
    layer3_outputs(2146) <= b;
    layer3_outputs(2147) <= a and b;
    layer3_outputs(2148) <= a and b;
    layer3_outputs(2149) <= not (a or b);
    layer3_outputs(2150) <= b;
    layer3_outputs(2151) <= not a;
    layer3_outputs(2152) <= b and not a;
    layer3_outputs(2153) <= b and not a;
    layer3_outputs(2154) <= not (a and b);
    layer3_outputs(2155) <= not a;
    layer3_outputs(2156) <= a;
    layer3_outputs(2157) <= not a;
    layer3_outputs(2158) <= a;
    layer3_outputs(2159) <= b;
    layer3_outputs(2160) <= not b;
    layer3_outputs(2161) <= not (a or b);
    layer3_outputs(2162) <= '1';
    layer3_outputs(2163) <= a and b;
    layer3_outputs(2164) <= not b or a;
    layer3_outputs(2165) <= not (a xor b);
    layer3_outputs(2166) <= not b;
    layer3_outputs(2167) <= b;
    layer3_outputs(2168) <= a and b;
    layer3_outputs(2169) <= not a;
    layer3_outputs(2170) <= not a or b;
    layer3_outputs(2171) <= a;
    layer3_outputs(2172) <= not b;
    layer3_outputs(2173) <= not a;
    layer3_outputs(2174) <= not b;
    layer3_outputs(2175) <= not (a and b);
    layer3_outputs(2176) <= a or b;
    layer3_outputs(2177) <= not (a and b);
    layer3_outputs(2178) <= not a;
    layer3_outputs(2179) <= b;
    layer3_outputs(2180) <= a;
    layer3_outputs(2181) <= a xor b;
    layer3_outputs(2182) <= a and not b;
    layer3_outputs(2183) <= not b;
    layer3_outputs(2184) <= not b or a;
    layer3_outputs(2185) <= not a or b;
    layer3_outputs(2186) <= a and not b;
    layer3_outputs(2187) <= not a;
    layer3_outputs(2188) <= not (a or b);
    layer3_outputs(2189) <= not b or a;
    layer3_outputs(2190) <= not b or a;
    layer3_outputs(2191) <= not b or a;
    layer3_outputs(2192) <= not (a and b);
    layer3_outputs(2193) <= not b;
    layer3_outputs(2194) <= not a;
    layer3_outputs(2195) <= a;
    layer3_outputs(2196) <= not (a xor b);
    layer3_outputs(2197) <= a and not b;
    layer3_outputs(2198) <= not b or a;
    layer3_outputs(2199) <= b and not a;
    layer3_outputs(2200) <= not (a or b);
    layer3_outputs(2201) <= a or b;
    layer3_outputs(2202) <= b and not a;
    layer3_outputs(2203) <= a and not b;
    layer3_outputs(2204) <= a;
    layer3_outputs(2205) <= not b;
    layer3_outputs(2206) <= b;
    layer3_outputs(2207) <= not a;
    layer3_outputs(2208) <= a;
    layer3_outputs(2209) <= b;
    layer3_outputs(2210) <= a or b;
    layer3_outputs(2211) <= not b or a;
    layer3_outputs(2212) <= not a;
    layer3_outputs(2213) <= a and b;
    layer3_outputs(2214) <= not b;
    layer3_outputs(2215) <= '1';
    layer3_outputs(2216) <= not a;
    layer3_outputs(2217) <= not a or b;
    layer3_outputs(2218) <= a or b;
    layer3_outputs(2219) <= a or b;
    layer3_outputs(2220) <= not b or a;
    layer3_outputs(2221) <= a and b;
    layer3_outputs(2222) <= not b;
    layer3_outputs(2223) <= a;
    layer3_outputs(2224) <= a;
    layer3_outputs(2225) <= a and b;
    layer3_outputs(2226) <= a or b;
    layer3_outputs(2227) <= not b;
    layer3_outputs(2228) <= not a;
    layer3_outputs(2229) <= not (a or b);
    layer3_outputs(2230) <= a and b;
    layer3_outputs(2231) <= a and not b;
    layer3_outputs(2232) <= not (a or b);
    layer3_outputs(2233) <= not b;
    layer3_outputs(2234) <= a and b;
    layer3_outputs(2235) <= not b;
    layer3_outputs(2236) <= a and not b;
    layer3_outputs(2237) <= not b or a;
    layer3_outputs(2238) <= a;
    layer3_outputs(2239) <= a xor b;
    layer3_outputs(2240) <= b and not a;
    layer3_outputs(2241) <= b;
    layer3_outputs(2242) <= b;
    layer3_outputs(2243) <= not b or a;
    layer3_outputs(2244) <= not a or b;
    layer3_outputs(2245) <= b and not a;
    layer3_outputs(2246) <= b;
    layer3_outputs(2247) <= a and not b;
    layer3_outputs(2248) <= '0';
    layer3_outputs(2249) <= a;
    layer3_outputs(2250) <= not (a or b);
    layer3_outputs(2251) <= not (a and b);
    layer3_outputs(2252) <= a and not b;
    layer3_outputs(2253) <= not b;
    layer3_outputs(2254) <= not a;
    layer3_outputs(2255) <= a and b;
    layer3_outputs(2256) <= not (a or b);
    layer3_outputs(2257) <= b;
    layer3_outputs(2258) <= not a or b;
    layer3_outputs(2259) <= a xor b;
    layer3_outputs(2260) <= not (a xor b);
    layer3_outputs(2261) <= not (a xor b);
    layer3_outputs(2262) <= a or b;
    layer3_outputs(2263) <= not b;
    layer3_outputs(2264) <= b;
    layer3_outputs(2265) <= b and not a;
    layer3_outputs(2266) <= a;
    layer3_outputs(2267) <= '0';
    layer3_outputs(2268) <= not (a or b);
    layer3_outputs(2269) <= a and not b;
    layer3_outputs(2270) <= a or b;
    layer3_outputs(2271) <= not a;
    layer3_outputs(2272) <= b and not a;
    layer3_outputs(2273) <= not (a or b);
    layer3_outputs(2274) <= b;
    layer3_outputs(2275) <= a;
    layer3_outputs(2276) <= a xor b;
    layer3_outputs(2277) <= not a;
    layer3_outputs(2278) <= not (a xor b);
    layer3_outputs(2279) <= '0';
    layer3_outputs(2280) <= not a or b;
    layer3_outputs(2281) <= not (a and b);
    layer3_outputs(2282) <= a and not b;
    layer3_outputs(2283) <= not (a or b);
    layer3_outputs(2284) <= a and not b;
    layer3_outputs(2285) <= a or b;
    layer3_outputs(2286) <= a xor b;
    layer3_outputs(2287) <= not a;
    layer3_outputs(2288) <= a or b;
    layer3_outputs(2289) <= a;
    layer3_outputs(2290) <= a and b;
    layer3_outputs(2291) <= not (a or b);
    layer3_outputs(2292) <= b;
    layer3_outputs(2293) <= not a;
    layer3_outputs(2294) <= a;
    layer3_outputs(2295) <= not b;
    layer3_outputs(2296) <= not (a or b);
    layer3_outputs(2297) <= a and b;
    layer3_outputs(2298) <= a or b;
    layer3_outputs(2299) <= a and b;
    layer3_outputs(2300) <= not (a and b);
    layer3_outputs(2301) <= not (a and b);
    layer3_outputs(2302) <= a;
    layer3_outputs(2303) <= a xor b;
    layer3_outputs(2304) <= not b;
    layer3_outputs(2305) <= a;
    layer3_outputs(2306) <= not (a or b);
    layer3_outputs(2307) <= not b;
    layer3_outputs(2308) <= b and not a;
    layer3_outputs(2309) <= a;
    layer3_outputs(2310) <= not a;
    layer3_outputs(2311) <= not (a and b);
    layer3_outputs(2312) <= not b;
    layer3_outputs(2313) <= a;
    layer3_outputs(2314) <= not b;
    layer3_outputs(2315) <= not (a or b);
    layer3_outputs(2316) <= not b or a;
    layer3_outputs(2317) <= not a;
    layer3_outputs(2318) <= a and not b;
    layer3_outputs(2319) <= b;
    layer3_outputs(2320) <= b and not a;
    layer3_outputs(2321) <= a and not b;
    layer3_outputs(2322) <= not b;
    layer3_outputs(2323) <= not (a and b);
    layer3_outputs(2324) <= a xor b;
    layer3_outputs(2325) <= a;
    layer3_outputs(2326) <= a xor b;
    layer3_outputs(2327) <= a and b;
    layer3_outputs(2328) <= b;
    layer3_outputs(2329) <= not (a or b);
    layer3_outputs(2330) <= a or b;
    layer3_outputs(2331) <= not (a or b);
    layer3_outputs(2332) <= a and not b;
    layer3_outputs(2333) <= not (a and b);
    layer3_outputs(2334) <= '1';
    layer3_outputs(2335) <= a;
    layer3_outputs(2336) <= a;
    layer3_outputs(2337) <= not (a xor b);
    layer3_outputs(2338) <= a xor b;
    layer3_outputs(2339) <= not b;
    layer3_outputs(2340) <= not a or b;
    layer3_outputs(2341) <= a or b;
    layer3_outputs(2342) <= a and b;
    layer3_outputs(2343) <= not (a xor b);
    layer3_outputs(2344) <= not b;
    layer3_outputs(2345) <= a;
    layer3_outputs(2346) <= '1';
    layer3_outputs(2347) <= b;
    layer3_outputs(2348) <= not b;
    layer3_outputs(2349) <= not (a xor b);
    layer3_outputs(2350) <= not a or b;
    layer3_outputs(2351) <= not b or a;
    layer3_outputs(2352) <= b and not a;
    layer3_outputs(2353) <= a xor b;
    layer3_outputs(2354) <= b;
    layer3_outputs(2355) <= b;
    layer3_outputs(2356) <= not a;
    layer3_outputs(2357) <= not a;
    layer3_outputs(2358) <= not b;
    layer3_outputs(2359) <= not (a or b);
    layer3_outputs(2360) <= a or b;
    layer3_outputs(2361) <= not a;
    layer3_outputs(2362) <= a;
    layer3_outputs(2363) <= not a;
    layer3_outputs(2364) <= a;
    layer3_outputs(2365) <= not (a xor b);
    layer3_outputs(2366) <= a;
    layer3_outputs(2367) <= a xor b;
    layer3_outputs(2368) <= not a;
    layer3_outputs(2369) <= a;
    layer3_outputs(2370) <= a or b;
    layer3_outputs(2371) <= a;
    layer3_outputs(2372) <= b;
    layer3_outputs(2373) <= a or b;
    layer3_outputs(2374) <= not b;
    layer3_outputs(2375) <= not b;
    layer3_outputs(2376) <= b;
    layer3_outputs(2377) <= a;
    layer3_outputs(2378) <= not a or b;
    layer3_outputs(2379) <= not b or a;
    layer3_outputs(2380) <= not a;
    layer3_outputs(2381) <= a and b;
    layer3_outputs(2382) <= a;
    layer3_outputs(2383) <= '0';
    layer3_outputs(2384) <= a and not b;
    layer3_outputs(2385) <= b;
    layer3_outputs(2386) <= a or b;
    layer3_outputs(2387) <= a and b;
    layer3_outputs(2388) <= not (a and b);
    layer3_outputs(2389) <= not b;
    layer3_outputs(2390) <= b;
    layer3_outputs(2391) <= '0';
    layer3_outputs(2392) <= a xor b;
    layer3_outputs(2393) <= a and b;
    layer3_outputs(2394) <= a and b;
    layer3_outputs(2395) <= a;
    layer3_outputs(2396) <= not (a xor b);
    layer3_outputs(2397) <= not (a xor b);
    layer3_outputs(2398) <= not (a or b);
    layer3_outputs(2399) <= a or b;
    layer3_outputs(2400) <= a;
    layer3_outputs(2401) <= not a;
    layer3_outputs(2402) <= a or b;
    layer3_outputs(2403) <= a and b;
    layer3_outputs(2404) <= a xor b;
    layer3_outputs(2405) <= not b;
    layer3_outputs(2406) <= b and not a;
    layer3_outputs(2407) <= not b;
    layer3_outputs(2408) <= a;
    layer3_outputs(2409) <= a;
    layer3_outputs(2410) <= not b or a;
    layer3_outputs(2411) <= a xor b;
    layer3_outputs(2412) <= a;
    layer3_outputs(2413) <= not (a or b);
    layer3_outputs(2414) <= not (a xor b);
    layer3_outputs(2415) <= not b or a;
    layer3_outputs(2416) <= a and not b;
    layer3_outputs(2417) <= not b;
    layer3_outputs(2418) <= a or b;
    layer3_outputs(2419) <= not a;
    layer3_outputs(2420) <= not a;
    layer3_outputs(2421) <= not (a or b);
    layer3_outputs(2422) <= a;
    layer3_outputs(2423) <= a or b;
    layer3_outputs(2424) <= not a;
    layer3_outputs(2425) <= not a;
    layer3_outputs(2426) <= a;
    layer3_outputs(2427) <= a;
    layer3_outputs(2428) <= a or b;
    layer3_outputs(2429) <= not b or a;
    layer3_outputs(2430) <= not b;
    layer3_outputs(2431) <= not (a xor b);
    layer3_outputs(2432) <= a and not b;
    layer3_outputs(2433) <= not (a and b);
    layer3_outputs(2434) <= a or b;
    layer3_outputs(2435) <= not b or a;
    layer3_outputs(2436) <= a or b;
    layer3_outputs(2437) <= '1';
    layer3_outputs(2438) <= '0';
    layer3_outputs(2439) <= b;
    layer3_outputs(2440) <= not b;
    layer3_outputs(2441) <= not b;
    layer3_outputs(2442) <= not b or a;
    layer3_outputs(2443) <= b and not a;
    layer3_outputs(2444) <= a;
    layer3_outputs(2445) <= a;
    layer3_outputs(2446) <= a xor b;
    layer3_outputs(2447) <= not a or b;
    layer3_outputs(2448) <= not b;
    layer3_outputs(2449) <= not (a or b);
    layer3_outputs(2450) <= b and not a;
    layer3_outputs(2451) <= a and not b;
    layer3_outputs(2452) <= a and b;
    layer3_outputs(2453) <= not (a or b);
    layer3_outputs(2454) <= b;
    layer3_outputs(2455) <= '1';
    layer3_outputs(2456) <= a xor b;
    layer3_outputs(2457) <= not b;
    layer3_outputs(2458) <= not a;
    layer3_outputs(2459) <= a or b;
    layer3_outputs(2460) <= a and not b;
    layer3_outputs(2461) <= not b;
    layer3_outputs(2462) <= a;
    layer3_outputs(2463) <= not (a xor b);
    layer3_outputs(2464) <= not a or b;
    layer3_outputs(2465) <= not (a and b);
    layer3_outputs(2466) <= a and b;
    layer3_outputs(2467) <= not b;
    layer3_outputs(2468) <= a;
    layer3_outputs(2469) <= a;
    layer3_outputs(2470) <= not a or b;
    layer3_outputs(2471) <= not (a xor b);
    layer3_outputs(2472) <= not b or a;
    layer3_outputs(2473) <= a;
    layer3_outputs(2474) <= a;
    layer3_outputs(2475) <= b;
    layer3_outputs(2476) <= b;
    layer3_outputs(2477) <= a;
    layer3_outputs(2478) <= not (a and b);
    layer3_outputs(2479) <= not a;
    layer3_outputs(2480) <= a xor b;
    layer3_outputs(2481) <= not a or b;
    layer3_outputs(2482) <= not (a or b);
    layer3_outputs(2483) <= a;
    layer3_outputs(2484) <= not a or b;
    layer3_outputs(2485) <= not (a or b);
    layer3_outputs(2486) <= not a;
    layer3_outputs(2487) <= not (a and b);
    layer3_outputs(2488) <= a xor b;
    layer3_outputs(2489) <= not b or a;
    layer3_outputs(2490) <= not (a xor b);
    layer3_outputs(2491) <= a and not b;
    layer3_outputs(2492) <= not b or a;
    layer3_outputs(2493) <= a;
    layer3_outputs(2494) <= b;
    layer3_outputs(2495) <= a and b;
    layer3_outputs(2496) <= a;
    layer3_outputs(2497) <= a or b;
    layer3_outputs(2498) <= a;
    layer3_outputs(2499) <= a or b;
    layer3_outputs(2500) <= not (a xor b);
    layer3_outputs(2501) <= not b or a;
    layer3_outputs(2502) <= a;
    layer3_outputs(2503) <= not b;
    layer3_outputs(2504) <= b;
    layer3_outputs(2505) <= a xor b;
    layer3_outputs(2506) <= not b or a;
    layer3_outputs(2507) <= not a;
    layer3_outputs(2508) <= not a;
    layer3_outputs(2509) <= not (a or b);
    layer3_outputs(2510) <= a;
    layer3_outputs(2511) <= '1';
    layer3_outputs(2512) <= not a;
    layer3_outputs(2513) <= a or b;
    layer3_outputs(2514) <= a or b;
    layer3_outputs(2515) <= not a;
    layer3_outputs(2516) <= a or b;
    layer3_outputs(2517) <= not a or b;
    layer3_outputs(2518) <= a;
    layer3_outputs(2519) <= '1';
    layer3_outputs(2520) <= not (a or b);
    layer3_outputs(2521) <= b;
    layer3_outputs(2522) <= not b or a;
    layer3_outputs(2523) <= not b;
    layer3_outputs(2524) <= a;
    layer3_outputs(2525) <= a or b;
    layer3_outputs(2526) <= not a;
    layer3_outputs(2527) <= a and b;
    layer3_outputs(2528) <= not (a xor b);
    layer3_outputs(2529) <= a or b;
    layer3_outputs(2530) <= not a;
    layer3_outputs(2531) <= a;
    layer3_outputs(2532) <= b;
    layer3_outputs(2533) <= not a;
    layer3_outputs(2534) <= not b;
    layer3_outputs(2535) <= a and not b;
    layer3_outputs(2536) <= not a;
    layer3_outputs(2537) <= a or b;
    layer3_outputs(2538) <= not (a or b);
    layer3_outputs(2539) <= not a or b;
    layer3_outputs(2540) <= a or b;
    layer3_outputs(2541) <= not b;
    layer3_outputs(2542) <= not b or a;
    layer3_outputs(2543) <= not b;
    layer3_outputs(2544) <= not b;
    layer3_outputs(2545) <= not (a or b);
    layer3_outputs(2546) <= not b;
    layer3_outputs(2547) <= not a;
    layer3_outputs(2548) <= b;
    layer3_outputs(2549) <= a or b;
    layer3_outputs(2550) <= a or b;
    layer3_outputs(2551) <= not b;
    layer3_outputs(2552) <= not (a or b);
    layer3_outputs(2553) <= b and not a;
    layer3_outputs(2554) <= not b or a;
    layer3_outputs(2555) <= not b;
    layer3_outputs(2556) <= not a;
    layer3_outputs(2557) <= not b or a;
    layer3_outputs(2558) <= a;
    layer3_outputs(2559) <= not b;
    layer3_outputs(2560) <= not b;
    layer3_outputs(2561) <= a xor b;
    layer3_outputs(2562) <= not b;
    layer3_outputs(2563) <= b;
    layer3_outputs(2564) <= not b;
    layer3_outputs(2565) <= a and not b;
    layer3_outputs(2566) <= a and b;
    layer3_outputs(2567) <= not a;
    layer3_outputs(2568) <= a or b;
    layer3_outputs(2569) <= not a or b;
    layer3_outputs(2570) <= b;
    layer3_outputs(2571) <= a or b;
    layer3_outputs(2572) <= a;
    layer3_outputs(2573) <= a and b;
    layer3_outputs(2574) <= not b or a;
    layer3_outputs(2575) <= a xor b;
    layer3_outputs(2576) <= not b;
    layer3_outputs(2577) <= not (a and b);
    layer3_outputs(2578) <= not b or a;
    layer3_outputs(2579) <= a;
    layer3_outputs(2580) <= a or b;
    layer3_outputs(2581) <= b and not a;
    layer3_outputs(2582) <= '1';
    layer3_outputs(2583) <= a and not b;
    layer3_outputs(2584) <= a and not b;
    layer3_outputs(2585) <= a xor b;
    layer3_outputs(2586) <= a and b;
    layer3_outputs(2587) <= b;
    layer3_outputs(2588) <= not a or b;
    layer3_outputs(2589) <= b;
    layer3_outputs(2590) <= not b or a;
    layer3_outputs(2591) <= not b;
    layer3_outputs(2592) <= not b;
    layer3_outputs(2593) <= not (a or b);
    layer3_outputs(2594) <= a xor b;
    layer3_outputs(2595) <= a;
    layer3_outputs(2596) <= not b;
    layer3_outputs(2597) <= not a;
    layer3_outputs(2598) <= not a;
    layer3_outputs(2599) <= not (a or b);
    layer3_outputs(2600) <= not (a and b);
    layer3_outputs(2601) <= a and not b;
    layer3_outputs(2602) <= not b;
    layer3_outputs(2603) <= a xor b;
    layer3_outputs(2604) <= a;
    layer3_outputs(2605) <= not b;
    layer3_outputs(2606) <= not b;
    layer3_outputs(2607) <= b;
    layer3_outputs(2608) <= not a or b;
    layer3_outputs(2609) <= a;
    layer3_outputs(2610) <= a and b;
    layer3_outputs(2611) <= not b or a;
    layer3_outputs(2612) <= b;
    layer3_outputs(2613) <= not (a or b);
    layer3_outputs(2614) <= not a or b;
    layer3_outputs(2615) <= not (a or b);
    layer3_outputs(2616) <= a and not b;
    layer3_outputs(2617) <= not b;
    layer3_outputs(2618) <= not b or a;
    layer3_outputs(2619) <= a and b;
    layer3_outputs(2620) <= not a;
    layer3_outputs(2621) <= not a;
    layer3_outputs(2622) <= not a or b;
    layer3_outputs(2623) <= not b or a;
    layer3_outputs(2624) <= not (a and b);
    layer3_outputs(2625) <= not b;
    layer3_outputs(2626) <= '1';
    layer3_outputs(2627) <= not (a or b);
    layer3_outputs(2628) <= not a;
    layer3_outputs(2629) <= a and not b;
    layer3_outputs(2630) <= not a or b;
    layer3_outputs(2631) <= a and b;
    layer3_outputs(2632) <= a;
    layer3_outputs(2633) <= not (a or b);
    layer3_outputs(2634) <= not a;
    layer3_outputs(2635) <= not b;
    layer3_outputs(2636) <= not b;
    layer3_outputs(2637) <= not (a and b);
    layer3_outputs(2638) <= not b;
    layer3_outputs(2639) <= not b;
    layer3_outputs(2640) <= b;
    layer3_outputs(2641) <= '0';
    layer3_outputs(2642) <= not a;
    layer3_outputs(2643) <= b;
    layer3_outputs(2644) <= a;
    layer3_outputs(2645) <= a and not b;
    layer3_outputs(2646) <= not b;
    layer3_outputs(2647) <= b and not a;
    layer3_outputs(2648) <= not (a and b);
    layer3_outputs(2649) <= not a;
    layer3_outputs(2650) <= not b;
    layer3_outputs(2651) <= b and not a;
    layer3_outputs(2652) <= '1';
    layer3_outputs(2653) <= not a or b;
    layer3_outputs(2654) <= a or b;
    layer3_outputs(2655) <= a and b;
    layer3_outputs(2656) <= not (a xor b);
    layer3_outputs(2657) <= '1';
    layer3_outputs(2658) <= not b;
    layer3_outputs(2659) <= b;
    layer3_outputs(2660) <= a;
    layer3_outputs(2661) <= a xor b;
    layer3_outputs(2662) <= not a;
    layer3_outputs(2663) <= b;
    layer3_outputs(2664) <= a and not b;
    layer3_outputs(2665) <= not (a xor b);
    layer3_outputs(2666) <= a or b;
    layer3_outputs(2667) <= not a or b;
    layer3_outputs(2668) <= not b;
    layer3_outputs(2669) <= a and not b;
    layer3_outputs(2670) <= b and not a;
    layer3_outputs(2671) <= a xor b;
    layer3_outputs(2672) <= a;
    layer3_outputs(2673) <= a and b;
    layer3_outputs(2674) <= a or b;
    layer3_outputs(2675) <= not a or b;
    layer3_outputs(2676) <= a;
    layer3_outputs(2677) <= a or b;
    layer3_outputs(2678) <= b;
    layer3_outputs(2679) <= not b;
    layer3_outputs(2680) <= b and not a;
    layer3_outputs(2681) <= not a;
    layer3_outputs(2682) <= b and not a;
    layer3_outputs(2683) <= not (a and b);
    layer3_outputs(2684) <= a;
    layer3_outputs(2685) <= not b;
    layer3_outputs(2686) <= not a or b;
    layer3_outputs(2687) <= not a;
    layer3_outputs(2688) <= not (a and b);
    layer3_outputs(2689) <= not (a and b);
    layer3_outputs(2690) <= not a;
    layer3_outputs(2691) <= a and not b;
    layer3_outputs(2692) <= not a;
    layer3_outputs(2693) <= a and b;
    layer3_outputs(2694) <= a and b;
    layer3_outputs(2695) <= b;
    layer3_outputs(2696) <= b and not a;
    layer3_outputs(2697) <= not b;
    layer3_outputs(2698) <= a;
    layer3_outputs(2699) <= a and b;
    layer3_outputs(2700) <= not (a and b);
    layer3_outputs(2701) <= not b;
    layer3_outputs(2702) <= not b;
    layer3_outputs(2703) <= not b;
    layer3_outputs(2704) <= not b;
    layer3_outputs(2705) <= a or b;
    layer3_outputs(2706) <= b;
    layer3_outputs(2707) <= b;
    layer3_outputs(2708) <= not (a or b);
    layer3_outputs(2709) <= not b;
    layer3_outputs(2710) <= a and b;
    layer3_outputs(2711) <= not a;
    layer3_outputs(2712) <= not b or a;
    layer3_outputs(2713) <= a or b;
    layer3_outputs(2714) <= a and not b;
    layer3_outputs(2715) <= not (a or b);
    layer3_outputs(2716) <= b and not a;
    layer3_outputs(2717) <= a or b;
    layer3_outputs(2718) <= a or b;
    layer3_outputs(2719) <= a and not b;
    layer3_outputs(2720) <= not a or b;
    layer3_outputs(2721) <= not (a or b);
    layer3_outputs(2722) <= not a;
    layer3_outputs(2723) <= not b;
    layer3_outputs(2724) <= not (a and b);
    layer3_outputs(2725) <= a or b;
    layer3_outputs(2726) <= a or b;
    layer3_outputs(2727) <= a and not b;
    layer3_outputs(2728) <= not b;
    layer3_outputs(2729) <= not (a or b);
    layer3_outputs(2730) <= a and b;
    layer3_outputs(2731) <= not (a xor b);
    layer3_outputs(2732) <= not a;
    layer3_outputs(2733) <= a and not b;
    layer3_outputs(2734) <= a and b;
    layer3_outputs(2735) <= not b or a;
    layer3_outputs(2736) <= a xor b;
    layer3_outputs(2737) <= '0';
    layer3_outputs(2738) <= not b;
    layer3_outputs(2739) <= b and not a;
    layer3_outputs(2740) <= a;
    layer3_outputs(2741) <= not a;
    layer3_outputs(2742) <= not a or b;
    layer3_outputs(2743) <= a or b;
    layer3_outputs(2744) <= a;
    layer3_outputs(2745) <= b;
    layer3_outputs(2746) <= a or b;
    layer3_outputs(2747) <= not b;
    layer3_outputs(2748) <= a and not b;
    layer3_outputs(2749) <= b;
    layer3_outputs(2750) <= not (a xor b);
    layer3_outputs(2751) <= a;
    layer3_outputs(2752) <= a xor b;
    layer3_outputs(2753) <= not a;
    layer3_outputs(2754) <= '1';
    layer3_outputs(2755) <= b;
    layer3_outputs(2756) <= not a;
    layer3_outputs(2757) <= a and b;
    layer3_outputs(2758) <= not b or a;
    layer3_outputs(2759) <= not (a or b);
    layer3_outputs(2760) <= not (a or b);
    layer3_outputs(2761) <= a or b;
    layer3_outputs(2762) <= not (a or b);
    layer3_outputs(2763) <= not (a or b);
    layer3_outputs(2764) <= not (a xor b);
    layer3_outputs(2765) <= not a;
    layer3_outputs(2766) <= a;
    layer3_outputs(2767) <= a and not b;
    layer3_outputs(2768) <= a and not b;
    layer3_outputs(2769) <= not (a xor b);
    layer3_outputs(2770) <= a and not b;
    layer3_outputs(2771) <= a and b;
    layer3_outputs(2772) <= a;
    layer3_outputs(2773) <= not a;
    layer3_outputs(2774) <= b;
    layer3_outputs(2775) <= not a;
    layer3_outputs(2776) <= not a or b;
    layer3_outputs(2777) <= not (a or b);
    layer3_outputs(2778) <= a and not b;
    layer3_outputs(2779) <= b;
    layer3_outputs(2780) <= b;
    layer3_outputs(2781) <= a and b;
    layer3_outputs(2782) <= a and b;
    layer3_outputs(2783) <= '0';
    layer3_outputs(2784) <= a and b;
    layer3_outputs(2785) <= not b or a;
    layer3_outputs(2786) <= not b;
    layer3_outputs(2787) <= a xor b;
    layer3_outputs(2788) <= a;
    layer3_outputs(2789) <= b;
    layer3_outputs(2790) <= a and not b;
    layer3_outputs(2791) <= a;
    layer3_outputs(2792) <= b;
    layer3_outputs(2793) <= b;
    layer3_outputs(2794) <= not b;
    layer3_outputs(2795) <= not b;
    layer3_outputs(2796) <= a xor b;
    layer3_outputs(2797) <= not b or a;
    layer3_outputs(2798) <= not a;
    layer3_outputs(2799) <= not (a xor b);
    layer3_outputs(2800) <= a xor b;
    layer3_outputs(2801) <= '1';
    layer3_outputs(2802) <= not a;
    layer3_outputs(2803) <= not (a xor b);
    layer3_outputs(2804) <= a;
    layer3_outputs(2805) <= not b;
    layer3_outputs(2806) <= not b;
    layer3_outputs(2807) <= b;
    layer3_outputs(2808) <= not (a and b);
    layer3_outputs(2809) <= a;
    layer3_outputs(2810) <= not a;
    layer3_outputs(2811) <= b and not a;
    layer3_outputs(2812) <= b;
    layer3_outputs(2813) <= not a or b;
    layer3_outputs(2814) <= '0';
    layer3_outputs(2815) <= '1';
    layer3_outputs(2816) <= a;
    layer3_outputs(2817) <= a and b;
    layer3_outputs(2818) <= a;
    layer3_outputs(2819) <= b;
    layer3_outputs(2820) <= not (a and b);
    layer3_outputs(2821) <= not a or b;
    layer3_outputs(2822) <= '0';
    layer3_outputs(2823) <= not a;
    layer3_outputs(2824) <= not (a or b);
    layer3_outputs(2825) <= not (a and b);
    layer3_outputs(2826) <= b;
    layer3_outputs(2827) <= not b;
    layer3_outputs(2828) <= not b or a;
    layer3_outputs(2829) <= b;
    layer3_outputs(2830) <= not b;
    layer3_outputs(2831) <= b and not a;
    layer3_outputs(2832) <= not b;
    layer3_outputs(2833) <= not b or a;
    layer3_outputs(2834) <= not a or b;
    layer3_outputs(2835) <= not b;
    layer3_outputs(2836) <= a and not b;
    layer3_outputs(2837) <= not (a or b);
    layer3_outputs(2838) <= b and not a;
    layer3_outputs(2839) <= not b;
    layer3_outputs(2840) <= not a;
    layer3_outputs(2841) <= a xor b;
    layer3_outputs(2842) <= '0';
    layer3_outputs(2843) <= b;
    layer3_outputs(2844) <= not (a or b);
    layer3_outputs(2845) <= '0';
    layer3_outputs(2846) <= a and not b;
    layer3_outputs(2847) <= a or b;
    layer3_outputs(2848) <= not b;
    layer3_outputs(2849) <= b;
    layer3_outputs(2850) <= a;
    layer3_outputs(2851) <= not a;
    layer3_outputs(2852) <= a or b;
    layer3_outputs(2853) <= b;
    layer3_outputs(2854) <= not (a xor b);
    layer3_outputs(2855) <= a and not b;
    layer3_outputs(2856) <= b;
    layer3_outputs(2857) <= not (a or b);
    layer3_outputs(2858) <= a or b;
    layer3_outputs(2859) <= a and b;
    layer3_outputs(2860) <= not (a and b);
    layer3_outputs(2861) <= a xor b;
    layer3_outputs(2862) <= a;
    layer3_outputs(2863) <= not b;
    layer3_outputs(2864) <= a and b;
    layer3_outputs(2865) <= a and not b;
    layer3_outputs(2866) <= a;
    layer3_outputs(2867) <= a;
    layer3_outputs(2868) <= a or b;
    layer3_outputs(2869) <= a and b;
    layer3_outputs(2870) <= not (a or b);
    layer3_outputs(2871) <= not (a or b);
    layer3_outputs(2872) <= a;
    layer3_outputs(2873) <= b and not a;
    layer3_outputs(2874) <= not a or b;
    layer3_outputs(2875) <= a and b;
    layer3_outputs(2876) <= b;
    layer3_outputs(2877) <= a and not b;
    layer3_outputs(2878) <= not b;
    layer3_outputs(2879) <= b and not a;
    layer3_outputs(2880) <= not (a and b);
    layer3_outputs(2881) <= not a or b;
    layer3_outputs(2882) <= not (a or b);
    layer3_outputs(2883) <= a and b;
    layer3_outputs(2884) <= a and b;
    layer3_outputs(2885) <= not a;
    layer3_outputs(2886) <= not a or b;
    layer3_outputs(2887) <= not b;
    layer3_outputs(2888) <= b;
    layer3_outputs(2889) <= '0';
    layer3_outputs(2890) <= not (a or b);
    layer3_outputs(2891) <= not a;
    layer3_outputs(2892) <= not (a xor b);
    layer3_outputs(2893) <= not a or b;
    layer3_outputs(2894) <= not b;
    layer3_outputs(2895) <= not (a xor b);
    layer3_outputs(2896) <= not a or b;
    layer3_outputs(2897) <= a xor b;
    layer3_outputs(2898) <= a and not b;
    layer3_outputs(2899) <= not a or b;
    layer3_outputs(2900) <= not a or b;
    layer3_outputs(2901) <= not b or a;
    layer3_outputs(2902) <= not (a or b);
    layer3_outputs(2903) <= b;
    layer3_outputs(2904) <= a and b;
    layer3_outputs(2905) <= not (a xor b);
    layer3_outputs(2906) <= not (a and b);
    layer3_outputs(2907) <= b and not a;
    layer3_outputs(2908) <= a;
    layer3_outputs(2909) <= not b or a;
    layer3_outputs(2910) <= not b;
    layer3_outputs(2911) <= not a or b;
    layer3_outputs(2912) <= a xor b;
    layer3_outputs(2913) <= a and not b;
    layer3_outputs(2914) <= a xor b;
    layer3_outputs(2915) <= b and not a;
    layer3_outputs(2916) <= not a or b;
    layer3_outputs(2917) <= b and not a;
    layer3_outputs(2918) <= a;
    layer3_outputs(2919) <= a or b;
    layer3_outputs(2920) <= not b;
    layer3_outputs(2921) <= not a or b;
    layer3_outputs(2922) <= not b;
    layer3_outputs(2923) <= a and not b;
    layer3_outputs(2924) <= a;
    layer3_outputs(2925) <= a xor b;
    layer3_outputs(2926) <= a;
    layer3_outputs(2927) <= b;
    layer3_outputs(2928) <= b and not a;
    layer3_outputs(2929) <= not a;
    layer3_outputs(2930) <= not a;
    layer3_outputs(2931) <= a;
    layer3_outputs(2932) <= not b or a;
    layer3_outputs(2933) <= '1';
    layer3_outputs(2934) <= a;
    layer3_outputs(2935) <= not a;
    layer3_outputs(2936) <= not b;
    layer3_outputs(2937) <= not b;
    layer3_outputs(2938) <= a and b;
    layer3_outputs(2939) <= not (a xor b);
    layer3_outputs(2940) <= not b or a;
    layer3_outputs(2941) <= not a;
    layer3_outputs(2942) <= not (a xor b);
    layer3_outputs(2943) <= not b;
    layer3_outputs(2944) <= not (a xor b);
    layer3_outputs(2945) <= a or b;
    layer3_outputs(2946) <= b;
    layer3_outputs(2947) <= not a or b;
    layer3_outputs(2948) <= not (a xor b);
    layer3_outputs(2949) <= a or b;
    layer3_outputs(2950) <= a;
    layer3_outputs(2951) <= not (a or b);
    layer3_outputs(2952) <= not a or b;
    layer3_outputs(2953) <= b;
    layer3_outputs(2954) <= not (a or b);
    layer3_outputs(2955) <= not b or a;
    layer3_outputs(2956) <= a and not b;
    layer3_outputs(2957) <= not b or a;
    layer3_outputs(2958) <= not b;
    layer3_outputs(2959) <= b and not a;
    layer3_outputs(2960) <= b;
    layer3_outputs(2961) <= b and not a;
    layer3_outputs(2962) <= not (a or b);
    layer3_outputs(2963) <= not (a xor b);
    layer3_outputs(2964) <= not b;
    layer3_outputs(2965) <= not (a or b);
    layer3_outputs(2966) <= not b;
    layer3_outputs(2967) <= not (a xor b);
    layer3_outputs(2968) <= a xor b;
    layer3_outputs(2969) <= b;
    layer3_outputs(2970) <= a and b;
    layer3_outputs(2971) <= not (a xor b);
    layer3_outputs(2972) <= a xor b;
    layer3_outputs(2973) <= '1';
    layer3_outputs(2974) <= not a;
    layer3_outputs(2975) <= b;
    layer3_outputs(2976) <= not (a xor b);
    layer3_outputs(2977) <= a and b;
    layer3_outputs(2978) <= b;
    layer3_outputs(2979) <= a and not b;
    layer3_outputs(2980) <= a or b;
    layer3_outputs(2981) <= a or b;
    layer3_outputs(2982) <= b;
    layer3_outputs(2983) <= b;
    layer3_outputs(2984) <= a or b;
    layer3_outputs(2985) <= a and b;
    layer3_outputs(2986) <= a and not b;
    layer3_outputs(2987) <= a or b;
    layer3_outputs(2988) <= a and b;
    layer3_outputs(2989) <= not b;
    layer3_outputs(2990) <= not b;
    layer3_outputs(2991) <= not (a or b);
    layer3_outputs(2992) <= not (a and b);
    layer3_outputs(2993) <= a;
    layer3_outputs(2994) <= not a or b;
    layer3_outputs(2995) <= a and b;
    layer3_outputs(2996) <= not b or a;
    layer3_outputs(2997) <= not (a or b);
    layer3_outputs(2998) <= a;
    layer3_outputs(2999) <= not (a xor b);
    layer3_outputs(3000) <= not a or b;
    layer3_outputs(3001) <= not b;
    layer3_outputs(3002) <= b and not a;
    layer3_outputs(3003) <= not a or b;
    layer3_outputs(3004) <= not a or b;
    layer3_outputs(3005) <= not b or a;
    layer3_outputs(3006) <= '1';
    layer3_outputs(3007) <= a and not b;
    layer3_outputs(3008) <= not a or b;
    layer3_outputs(3009) <= b;
    layer3_outputs(3010) <= a;
    layer3_outputs(3011) <= not (a and b);
    layer3_outputs(3012) <= not (a xor b);
    layer3_outputs(3013) <= a and not b;
    layer3_outputs(3014) <= a and b;
    layer3_outputs(3015) <= not a or b;
    layer3_outputs(3016) <= not b or a;
    layer3_outputs(3017) <= a and b;
    layer3_outputs(3018) <= not b;
    layer3_outputs(3019) <= not b or a;
    layer3_outputs(3020) <= not (a and b);
    layer3_outputs(3021) <= not (a and b);
    layer3_outputs(3022) <= b;
    layer3_outputs(3023) <= b;
    layer3_outputs(3024) <= not b;
    layer3_outputs(3025) <= b;
    layer3_outputs(3026) <= not (a and b);
    layer3_outputs(3027) <= a or b;
    layer3_outputs(3028) <= not (a xor b);
    layer3_outputs(3029) <= a;
    layer3_outputs(3030) <= not b or a;
    layer3_outputs(3031) <= not (a or b);
    layer3_outputs(3032) <= b and not a;
    layer3_outputs(3033) <= a and not b;
    layer3_outputs(3034) <= a;
    layer3_outputs(3035) <= not (a and b);
    layer3_outputs(3036) <= b;
    layer3_outputs(3037) <= a;
    layer3_outputs(3038) <= not b;
    layer3_outputs(3039) <= not (a or b);
    layer3_outputs(3040) <= a;
    layer3_outputs(3041) <= not b or a;
    layer3_outputs(3042) <= not (a or b);
    layer3_outputs(3043) <= not a;
    layer3_outputs(3044) <= not a;
    layer3_outputs(3045) <= b;
    layer3_outputs(3046) <= not b or a;
    layer3_outputs(3047) <= not a;
    layer3_outputs(3048) <= b and not a;
    layer3_outputs(3049) <= a and not b;
    layer3_outputs(3050) <= a;
    layer3_outputs(3051) <= not a or b;
    layer3_outputs(3052) <= a and not b;
    layer3_outputs(3053) <= not a or b;
    layer3_outputs(3054) <= not a or b;
    layer3_outputs(3055) <= not a;
    layer3_outputs(3056) <= '1';
    layer3_outputs(3057) <= not (a or b);
    layer3_outputs(3058) <= not a;
    layer3_outputs(3059) <= b and not a;
    layer3_outputs(3060) <= a or b;
    layer3_outputs(3061) <= a and not b;
    layer3_outputs(3062) <= not (a and b);
    layer3_outputs(3063) <= not (a or b);
    layer3_outputs(3064) <= not a or b;
    layer3_outputs(3065) <= not a;
    layer3_outputs(3066) <= not a or b;
    layer3_outputs(3067) <= not a;
    layer3_outputs(3068) <= a xor b;
    layer3_outputs(3069) <= not a or b;
    layer3_outputs(3070) <= a xor b;
    layer3_outputs(3071) <= a;
    layer3_outputs(3072) <= a and not b;
    layer3_outputs(3073) <= not b or a;
    layer3_outputs(3074) <= not a or b;
    layer3_outputs(3075) <= b and not a;
    layer3_outputs(3076) <= b and not a;
    layer3_outputs(3077) <= not b;
    layer3_outputs(3078) <= not a or b;
    layer3_outputs(3079) <= a xor b;
    layer3_outputs(3080) <= '1';
    layer3_outputs(3081) <= not (a or b);
    layer3_outputs(3082) <= not b;
    layer3_outputs(3083) <= a;
    layer3_outputs(3084) <= b;
    layer3_outputs(3085) <= a or b;
    layer3_outputs(3086) <= a;
    layer3_outputs(3087) <= not (a and b);
    layer3_outputs(3088) <= a and b;
    layer3_outputs(3089) <= a;
    layer3_outputs(3090) <= b;
    layer3_outputs(3091) <= a;
    layer3_outputs(3092) <= b and not a;
    layer3_outputs(3093) <= not a or b;
    layer3_outputs(3094) <= b;
    layer3_outputs(3095) <= a;
    layer3_outputs(3096) <= a;
    layer3_outputs(3097) <= a and b;
    layer3_outputs(3098) <= not (a and b);
    layer3_outputs(3099) <= a and b;
    layer3_outputs(3100) <= '1';
    layer3_outputs(3101) <= b and not a;
    layer3_outputs(3102) <= a;
    layer3_outputs(3103) <= a and b;
    layer3_outputs(3104) <= not (a xor b);
    layer3_outputs(3105) <= '1';
    layer3_outputs(3106) <= not b;
    layer3_outputs(3107) <= not b;
    layer3_outputs(3108) <= b;
    layer3_outputs(3109) <= not b or a;
    layer3_outputs(3110) <= a;
    layer3_outputs(3111) <= not a;
    layer3_outputs(3112) <= a or b;
    layer3_outputs(3113) <= b;
    layer3_outputs(3114) <= not a or b;
    layer3_outputs(3115) <= b and not a;
    layer3_outputs(3116) <= not a;
    layer3_outputs(3117) <= not b;
    layer3_outputs(3118) <= '1';
    layer3_outputs(3119) <= not b or a;
    layer3_outputs(3120) <= b;
    layer3_outputs(3121) <= not b;
    layer3_outputs(3122) <= b and not a;
    layer3_outputs(3123) <= not b;
    layer3_outputs(3124) <= a and b;
    layer3_outputs(3125) <= b and not a;
    layer3_outputs(3126) <= a and b;
    layer3_outputs(3127) <= not (a and b);
    layer3_outputs(3128) <= b and not a;
    layer3_outputs(3129) <= not a;
    layer3_outputs(3130) <= a or b;
    layer3_outputs(3131) <= not b;
    layer3_outputs(3132) <= not a;
    layer3_outputs(3133) <= not b or a;
    layer3_outputs(3134) <= b;
    layer3_outputs(3135) <= not (a xor b);
    layer3_outputs(3136) <= not a or b;
    layer3_outputs(3137) <= a xor b;
    layer3_outputs(3138) <= not (a or b);
    layer3_outputs(3139) <= not a or b;
    layer3_outputs(3140) <= not a or b;
    layer3_outputs(3141) <= not b;
    layer3_outputs(3142) <= b and not a;
    layer3_outputs(3143) <= a or b;
    layer3_outputs(3144) <= b and not a;
    layer3_outputs(3145) <= not b;
    layer3_outputs(3146) <= a;
    layer3_outputs(3147) <= b;
    layer3_outputs(3148) <= b;
    layer3_outputs(3149) <= not (a or b);
    layer3_outputs(3150) <= not b or a;
    layer3_outputs(3151) <= a and b;
    layer3_outputs(3152) <= a and not b;
    layer3_outputs(3153) <= a or b;
    layer3_outputs(3154) <= not a;
    layer3_outputs(3155) <= b;
    layer3_outputs(3156) <= not (a or b);
    layer3_outputs(3157) <= a and not b;
    layer3_outputs(3158) <= not a;
    layer3_outputs(3159) <= not (a and b);
    layer3_outputs(3160) <= not b;
    layer3_outputs(3161) <= not b or a;
    layer3_outputs(3162) <= b and not a;
    layer3_outputs(3163) <= b;
    layer3_outputs(3164) <= not a;
    layer3_outputs(3165) <= not (a and b);
    layer3_outputs(3166) <= not a;
    layer3_outputs(3167) <= '0';
    layer3_outputs(3168) <= b and not a;
    layer3_outputs(3169) <= a or b;
    layer3_outputs(3170) <= a;
    layer3_outputs(3171) <= '1';
    layer3_outputs(3172) <= a xor b;
    layer3_outputs(3173) <= not (a xor b);
    layer3_outputs(3174) <= a and b;
    layer3_outputs(3175) <= '0';
    layer3_outputs(3176) <= a;
    layer3_outputs(3177) <= a xor b;
    layer3_outputs(3178) <= a;
    layer3_outputs(3179) <= not a or b;
    layer3_outputs(3180) <= b and not a;
    layer3_outputs(3181) <= a or b;
    layer3_outputs(3182) <= not (a xor b);
    layer3_outputs(3183) <= b and not a;
    layer3_outputs(3184) <= not b or a;
    layer3_outputs(3185) <= not b or a;
    layer3_outputs(3186) <= not a;
    layer3_outputs(3187) <= a xor b;
    layer3_outputs(3188) <= a or b;
    layer3_outputs(3189) <= '1';
    layer3_outputs(3190) <= b and not a;
    layer3_outputs(3191) <= a and b;
    layer3_outputs(3192) <= not (a or b);
    layer3_outputs(3193) <= b;
    layer3_outputs(3194) <= a;
    layer3_outputs(3195) <= not a or b;
    layer3_outputs(3196) <= a and not b;
    layer3_outputs(3197) <= not a;
    layer3_outputs(3198) <= not (a xor b);
    layer3_outputs(3199) <= b and not a;
    layer3_outputs(3200) <= b;
    layer3_outputs(3201) <= not b;
    layer3_outputs(3202) <= a or b;
    layer3_outputs(3203) <= b and not a;
    layer3_outputs(3204) <= b;
    layer3_outputs(3205) <= not (a or b);
    layer3_outputs(3206) <= not a;
    layer3_outputs(3207) <= a and b;
    layer3_outputs(3208) <= b;
    layer3_outputs(3209) <= a and b;
    layer3_outputs(3210) <= a and not b;
    layer3_outputs(3211) <= a;
    layer3_outputs(3212) <= a and not b;
    layer3_outputs(3213) <= not a;
    layer3_outputs(3214) <= a and b;
    layer3_outputs(3215) <= not a;
    layer3_outputs(3216) <= a xor b;
    layer3_outputs(3217) <= b and not a;
    layer3_outputs(3218) <= not a;
    layer3_outputs(3219) <= not (a or b);
    layer3_outputs(3220) <= a;
    layer3_outputs(3221) <= not (a xor b);
    layer3_outputs(3222) <= b;
    layer3_outputs(3223) <= a or b;
    layer3_outputs(3224) <= a and not b;
    layer3_outputs(3225) <= not b or a;
    layer3_outputs(3226) <= not (a and b);
    layer3_outputs(3227) <= b;
    layer3_outputs(3228) <= not (a or b);
    layer3_outputs(3229) <= a and not b;
    layer3_outputs(3230) <= not (a or b);
    layer3_outputs(3231) <= a and not b;
    layer3_outputs(3232) <= a xor b;
    layer3_outputs(3233) <= a or b;
    layer3_outputs(3234) <= not (a and b);
    layer3_outputs(3235) <= not a;
    layer3_outputs(3236) <= a;
    layer3_outputs(3237) <= a;
    layer3_outputs(3238) <= not (a or b);
    layer3_outputs(3239) <= b;
    layer3_outputs(3240) <= not a;
    layer3_outputs(3241) <= b;
    layer3_outputs(3242) <= not (a and b);
    layer3_outputs(3243) <= a;
    layer3_outputs(3244) <= not b;
    layer3_outputs(3245) <= a and not b;
    layer3_outputs(3246) <= not a or b;
    layer3_outputs(3247) <= not b;
    layer3_outputs(3248) <= not a or b;
    layer3_outputs(3249) <= a;
    layer3_outputs(3250) <= a or b;
    layer3_outputs(3251) <= b and not a;
    layer3_outputs(3252) <= not (a and b);
    layer3_outputs(3253) <= not b or a;
    layer3_outputs(3254) <= not b or a;
    layer3_outputs(3255) <= not b or a;
    layer3_outputs(3256) <= not (a and b);
    layer3_outputs(3257) <= a;
    layer3_outputs(3258) <= b;
    layer3_outputs(3259) <= not (a and b);
    layer3_outputs(3260) <= a or b;
    layer3_outputs(3261) <= a;
    layer3_outputs(3262) <= not (a and b);
    layer3_outputs(3263) <= not a or b;
    layer3_outputs(3264) <= not a;
    layer3_outputs(3265) <= a or b;
    layer3_outputs(3266) <= not (a and b);
    layer3_outputs(3267) <= not (a xor b);
    layer3_outputs(3268) <= not (a and b);
    layer3_outputs(3269) <= a and b;
    layer3_outputs(3270) <= not a or b;
    layer3_outputs(3271) <= a;
    layer3_outputs(3272) <= a and b;
    layer3_outputs(3273) <= not a;
    layer3_outputs(3274) <= not a or b;
    layer3_outputs(3275) <= not b or a;
    layer3_outputs(3276) <= a and not b;
    layer3_outputs(3277) <= b and not a;
    layer3_outputs(3278) <= not a or b;
    layer3_outputs(3279) <= not b;
    layer3_outputs(3280) <= b and not a;
    layer3_outputs(3281) <= not a;
    layer3_outputs(3282) <= not (a and b);
    layer3_outputs(3283) <= not a;
    layer3_outputs(3284) <= not (a or b);
    layer3_outputs(3285) <= a and b;
    layer3_outputs(3286) <= not a;
    layer3_outputs(3287) <= b;
    layer3_outputs(3288) <= not (a or b);
    layer3_outputs(3289) <= not (a xor b);
    layer3_outputs(3290) <= not (a or b);
    layer3_outputs(3291) <= not b;
    layer3_outputs(3292) <= not b or a;
    layer3_outputs(3293) <= b;
    layer3_outputs(3294) <= not a;
    layer3_outputs(3295) <= b and not a;
    layer3_outputs(3296) <= not b or a;
    layer3_outputs(3297) <= a;
    layer3_outputs(3298) <= a or b;
    layer3_outputs(3299) <= not a or b;
    layer3_outputs(3300) <= b;
    layer3_outputs(3301) <= not (a xor b);
    layer3_outputs(3302) <= a;
    layer3_outputs(3303) <= not a;
    layer3_outputs(3304) <= not a;
    layer3_outputs(3305) <= b;
    layer3_outputs(3306) <= not a;
    layer3_outputs(3307) <= a;
    layer3_outputs(3308) <= a and not b;
    layer3_outputs(3309) <= not (a and b);
    layer3_outputs(3310) <= '0';
    layer3_outputs(3311) <= a;
    layer3_outputs(3312) <= not b;
    layer3_outputs(3313) <= a or b;
    layer3_outputs(3314) <= a;
    layer3_outputs(3315) <= not (a and b);
    layer3_outputs(3316) <= b;
    layer3_outputs(3317) <= not a or b;
    layer3_outputs(3318) <= not (a xor b);
    layer3_outputs(3319) <= not a or b;
    layer3_outputs(3320) <= b and not a;
    layer3_outputs(3321) <= b;
    layer3_outputs(3322) <= not a;
    layer3_outputs(3323) <= a and b;
    layer3_outputs(3324) <= b;
    layer3_outputs(3325) <= a;
    layer3_outputs(3326) <= b and not a;
    layer3_outputs(3327) <= a and not b;
    layer3_outputs(3328) <= '0';
    layer3_outputs(3329) <= a xor b;
    layer3_outputs(3330) <= b;
    layer3_outputs(3331) <= not a;
    layer3_outputs(3332) <= not b;
    layer3_outputs(3333) <= not (a xor b);
    layer3_outputs(3334) <= not a;
    layer3_outputs(3335) <= a;
    layer3_outputs(3336) <= a xor b;
    layer3_outputs(3337) <= b;
    layer3_outputs(3338) <= not b;
    layer3_outputs(3339) <= not b or a;
    layer3_outputs(3340) <= not b;
    layer3_outputs(3341) <= a or b;
    layer3_outputs(3342) <= not b or a;
    layer3_outputs(3343) <= not a or b;
    layer3_outputs(3344) <= a or b;
    layer3_outputs(3345) <= a and b;
    layer3_outputs(3346) <= not (a and b);
    layer3_outputs(3347) <= b;
    layer3_outputs(3348) <= a and not b;
    layer3_outputs(3349) <= '0';
    layer3_outputs(3350) <= not a;
    layer3_outputs(3351) <= a or b;
    layer3_outputs(3352) <= a and b;
    layer3_outputs(3353) <= not b;
    layer3_outputs(3354) <= not (a xor b);
    layer3_outputs(3355) <= a and b;
    layer3_outputs(3356) <= b;
    layer3_outputs(3357) <= b and not a;
    layer3_outputs(3358) <= not a;
    layer3_outputs(3359) <= a or b;
    layer3_outputs(3360) <= b;
    layer3_outputs(3361) <= not b or a;
    layer3_outputs(3362) <= b and not a;
    layer3_outputs(3363) <= a xor b;
    layer3_outputs(3364) <= not a or b;
    layer3_outputs(3365) <= not b;
    layer3_outputs(3366) <= a and b;
    layer3_outputs(3367) <= not (a or b);
    layer3_outputs(3368) <= not a or b;
    layer3_outputs(3369) <= b;
    layer3_outputs(3370) <= not b;
    layer3_outputs(3371) <= a and not b;
    layer3_outputs(3372) <= a or b;
    layer3_outputs(3373) <= not b;
    layer3_outputs(3374) <= not a or b;
    layer3_outputs(3375) <= a;
    layer3_outputs(3376) <= '0';
    layer3_outputs(3377) <= not (a and b);
    layer3_outputs(3378) <= a and not b;
    layer3_outputs(3379) <= a or b;
    layer3_outputs(3380) <= a or b;
    layer3_outputs(3381) <= not a or b;
    layer3_outputs(3382) <= a;
    layer3_outputs(3383) <= '0';
    layer3_outputs(3384) <= not b;
    layer3_outputs(3385) <= not (a and b);
    layer3_outputs(3386) <= not (a xor b);
    layer3_outputs(3387) <= not a or b;
    layer3_outputs(3388) <= not (a or b);
    layer3_outputs(3389) <= a xor b;
    layer3_outputs(3390) <= not b;
    layer3_outputs(3391) <= not (a and b);
    layer3_outputs(3392) <= a;
    layer3_outputs(3393) <= a;
    layer3_outputs(3394) <= b;
    layer3_outputs(3395) <= not b or a;
    layer3_outputs(3396) <= not a;
    layer3_outputs(3397) <= '0';
    layer3_outputs(3398) <= a xor b;
    layer3_outputs(3399) <= not b;
    layer3_outputs(3400) <= not (a xor b);
    layer3_outputs(3401) <= b;
    layer3_outputs(3402) <= a and b;
    layer3_outputs(3403) <= b;
    layer3_outputs(3404) <= b and not a;
    layer3_outputs(3405) <= a;
    layer3_outputs(3406) <= not a;
    layer3_outputs(3407) <= a;
    layer3_outputs(3408) <= not b;
    layer3_outputs(3409) <= a;
    layer3_outputs(3410) <= b;
    layer3_outputs(3411) <= b;
    layer3_outputs(3412) <= not a or b;
    layer3_outputs(3413) <= a or b;
    layer3_outputs(3414) <= a and not b;
    layer3_outputs(3415) <= a or b;
    layer3_outputs(3416) <= not b or a;
    layer3_outputs(3417) <= not b;
    layer3_outputs(3418) <= b;
    layer3_outputs(3419) <= a and not b;
    layer3_outputs(3420) <= not a;
    layer3_outputs(3421) <= not (a xor b);
    layer3_outputs(3422) <= a;
    layer3_outputs(3423) <= not b or a;
    layer3_outputs(3424) <= not b;
    layer3_outputs(3425) <= not a;
    layer3_outputs(3426) <= a;
    layer3_outputs(3427) <= not a;
    layer3_outputs(3428) <= not b;
    layer3_outputs(3429) <= b;
    layer3_outputs(3430) <= '0';
    layer3_outputs(3431) <= not b;
    layer3_outputs(3432) <= not (a xor b);
    layer3_outputs(3433) <= b;
    layer3_outputs(3434) <= not b;
    layer3_outputs(3435) <= not b or a;
    layer3_outputs(3436) <= not b;
    layer3_outputs(3437) <= not b or a;
    layer3_outputs(3438) <= not (a and b);
    layer3_outputs(3439) <= b;
    layer3_outputs(3440) <= not (a xor b);
    layer3_outputs(3441) <= a;
    layer3_outputs(3442) <= a xor b;
    layer3_outputs(3443) <= a;
    layer3_outputs(3444) <= b;
    layer3_outputs(3445) <= not b;
    layer3_outputs(3446) <= b and not a;
    layer3_outputs(3447) <= not (a and b);
    layer3_outputs(3448) <= not (a xor b);
    layer3_outputs(3449) <= not b or a;
    layer3_outputs(3450) <= not b;
    layer3_outputs(3451) <= not a or b;
    layer3_outputs(3452) <= a;
    layer3_outputs(3453) <= b and not a;
    layer3_outputs(3454) <= '0';
    layer3_outputs(3455) <= a and not b;
    layer3_outputs(3456) <= not b;
    layer3_outputs(3457) <= not (a or b);
    layer3_outputs(3458) <= not b or a;
    layer3_outputs(3459) <= b;
    layer3_outputs(3460) <= not (a xor b);
    layer3_outputs(3461) <= not (a or b);
    layer3_outputs(3462) <= b;
    layer3_outputs(3463) <= not (a xor b);
    layer3_outputs(3464) <= not a;
    layer3_outputs(3465) <= a and b;
    layer3_outputs(3466) <= not b;
    layer3_outputs(3467) <= not (a or b);
    layer3_outputs(3468) <= a and b;
    layer3_outputs(3469) <= b;
    layer3_outputs(3470) <= not (a xor b);
    layer3_outputs(3471) <= not b or a;
    layer3_outputs(3472) <= not a;
    layer3_outputs(3473) <= not (a xor b);
    layer3_outputs(3474) <= not a or b;
    layer3_outputs(3475) <= a;
    layer3_outputs(3476) <= not (a xor b);
    layer3_outputs(3477) <= a and b;
    layer3_outputs(3478) <= not (a xor b);
    layer3_outputs(3479) <= not b or a;
    layer3_outputs(3480) <= a and not b;
    layer3_outputs(3481) <= not a;
    layer3_outputs(3482) <= b;
    layer3_outputs(3483) <= b;
    layer3_outputs(3484) <= a;
    layer3_outputs(3485) <= b;
    layer3_outputs(3486) <= not (a or b);
    layer3_outputs(3487) <= a;
    layer3_outputs(3488) <= a or b;
    layer3_outputs(3489) <= a and b;
    layer3_outputs(3490) <= not b or a;
    layer3_outputs(3491) <= b and not a;
    layer3_outputs(3492) <= b;
    layer3_outputs(3493) <= not (a xor b);
    layer3_outputs(3494) <= not a;
    layer3_outputs(3495) <= not (a xor b);
    layer3_outputs(3496) <= not b or a;
    layer3_outputs(3497) <= a xor b;
    layer3_outputs(3498) <= not (a or b);
    layer3_outputs(3499) <= not b;
    layer3_outputs(3500) <= a xor b;
    layer3_outputs(3501) <= not a;
    layer3_outputs(3502) <= a and not b;
    layer3_outputs(3503) <= not b;
    layer3_outputs(3504) <= b;
    layer3_outputs(3505) <= b;
    layer3_outputs(3506) <= a xor b;
    layer3_outputs(3507) <= not a;
    layer3_outputs(3508) <= b;
    layer3_outputs(3509) <= a xor b;
    layer3_outputs(3510) <= not a;
    layer3_outputs(3511) <= not a;
    layer3_outputs(3512) <= not (a xor b);
    layer3_outputs(3513) <= b;
    layer3_outputs(3514) <= not b or a;
    layer3_outputs(3515) <= a and not b;
    layer3_outputs(3516) <= not b;
    layer3_outputs(3517) <= b;
    layer3_outputs(3518) <= a;
    layer3_outputs(3519) <= not (a xor b);
    layer3_outputs(3520) <= a;
    layer3_outputs(3521) <= b;
    layer3_outputs(3522) <= not b;
    layer3_outputs(3523) <= not b;
    layer3_outputs(3524) <= not a or b;
    layer3_outputs(3525) <= not a or b;
    layer3_outputs(3526) <= b and not a;
    layer3_outputs(3527) <= not b;
    layer3_outputs(3528) <= a;
    layer3_outputs(3529) <= not a;
    layer3_outputs(3530) <= b and not a;
    layer3_outputs(3531) <= b;
    layer3_outputs(3532) <= '0';
    layer3_outputs(3533) <= b;
    layer3_outputs(3534) <= b;
    layer3_outputs(3535) <= '0';
    layer3_outputs(3536) <= a;
    layer3_outputs(3537) <= b;
    layer3_outputs(3538) <= not (a xor b);
    layer3_outputs(3539) <= '1';
    layer3_outputs(3540) <= not (a xor b);
    layer3_outputs(3541) <= not (a and b);
    layer3_outputs(3542) <= a and not b;
    layer3_outputs(3543) <= b;
    layer3_outputs(3544) <= not a;
    layer3_outputs(3545) <= not a;
    layer3_outputs(3546) <= b and not a;
    layer3_outputs(3547) <= a and b;
    layer3_outputs(3548) <= a;
    layer3_outputs(3549) <= not b or a;
    layer3_outputs(3550) <= b;
    layer3_outputs(3551) <= not (a or b);
    layer3_outputs(3552) <= a and not b;
    layer3_outputs(3553) <= not (a and b);
    layer3_outputs(3554) <= not b;
    layer3_outputs(3555) <= a;
    layer3_outputs(3556) <= a xor b;
    layer3_outputs(3557) <= not a;
    layer3_outputs(3558) <= not b or a;
    layer3_outputs(3559) <= a xor b;
    layer3_outputs(3560) <= not a;
    layer3_outputs(3561) <= not a or b;
    layer3_outputs(3562) <= not b;
    layer3_outputs(3563) <= a and b;
    layer3_outputs(3564) <= b;
    layer3_outputs(3565) <= not a;
    layer3_outputs(3566) <= not (a xor b);
    layer3_outputs(3567) <= a and not b;
    layer3_outputs(3568) <= not a;
    layer3_outputs(3569) <= not a;
    layer3_outputs(3570) <= b;
    layer3_outputs(3571) <= b and not a;
    layer3_outputs(3572) <= b;
    layer3_outputs(3573) <= not b or a;
    layer3_outputs(3574) <= not a;
    layer3_outputs(3575) <= not b;
    layer3_outputs(3576) <= not a;
    layer3_outputs(3577) <= a;
    layer3_outputs(3578) <= a or b;
    layer3_outputs(3579) <= a;
    layer3_outputs(3580) <= not (a xor b);
    layer3_outputs(3581) <= a and b;
    layer3_outputs(3582) <= not a or b;
    layer3_outputs(3583) <= not b or a;
    layer3_outputs(3584) <= b and not a;
    layer3_outputs(3585) <= not a or b;
    layer3_outputs(3586) <= not a;
    layer3_outputs(3587) <= '0';
    layer3_outputs(3588) <= not (a or b);
    layer3_outputs(3589) <= not b;
    layer3_outputs(3590) <= a;
    layer3_outputs(3591) <= not a or b;
    layer3_outputs(3592) <= b;
    layer3_outputs(3593) <= not (a and b);
    layer3_outputs(3594) <= not a or b;
    layer3_outputs(3595) <= a and b;
    layer3_outputs(3596) <= not (a and b);
    layer3_outputs(3597) <= not b or a;
    layer3_outputs(3598) <= a xor b;
    layer3_outputs(3599) <= b;
    layer3_outputs(3600) <= a xor b;
    layer3_outputs(3601) <= a and not b;
    layer3_outputs(3602) <= not b or a;
    layer3_outputs(3603) <= not a;
    layer3_outputs(3604) <= a and b;
    layer3_outputs(3605) <= not b;
    layer3_outputs(3606) <= not b or a;
    layer3_outputs(3607) <= '0';
    layer3_outputs(3608) <= b and not a;
    layer3_outputs(3609) <= a or b;
    layer3_outputs(3610) <= not a or b;
    layer3_outputs(3611) <= not b or a;
    layer3_outputs(3612) <= b;
    layer3_outputs(3613) <= not b;
    layer3_outputs(3614) <= not (a and b);
    layer3_outputs(3615) <= b;
    layer3_outputs(3616) <= not a or b;
    layer3_outputs(3617) <= a;
    layer3_outputs(3618) <= a;
    layer3_outputs(3619) <= a or b;
    layer3_outputs(3620) <= a or b;
    layer3_outputs(3621) <= b;
    layer3_outputs(3622) <= not a or b;
    layer3_outputs(3623) <= a and not b;
    layer3_outputs(3624) <= a or b;
    layer3_outputs(3625) <= a and not b;
    layer3_outputs(3626) <= a and b;
    layer3_outputs(3627) <= not (a or b);
    layer3_outputs(3628) <= a;
    layer3_outputs(3629) <= not a or b;
    layer3_outputs(3630) <= not (a xor b);
    layer3_outputs(3631) <= b and not a;
    layer3_outputs(3632) <= b and not a;
    layer3_outputs(3633) <= b and not a;
    layer3_outputs(3634) <= not b;
    layer3_outputs(3635) <= a and b;
    layer3_outputs(3636) <= a;
    layer3_outputs(3637) <= a;
    layer3_outputs(3638) <= not a;
    layer3_outputs(3639) <= not b;
    layer3_outputs(3640) <= not a or b;
    layer3_outputs(3641) <= b;
    layer3_outputs(3642) <= a and not b;
    layer3_outputs(3643) <= not (a and b);
    layer3_outputs(3644) <= not a;
    layer3_outputs(3645) <= not b;
    layer3_outputs(3646) <= not a;
    layer3_outputs(3647) <= not b;
    layer3_outputs(3648) <= a;
    layer3_outputs(3649) <= not b;
    layer3_outputs(3650) <= not b or a;
    layer3_outputs(3651) <= a and not b;
    layer3_outputs(3652) <= a;
    layer3_outputs(3653) <= a xor b;
    layer3_outputs(3654) <= b and not a;
    layer3_outputs(3655) <= not (a and b);
    layer3_outputs(3656) <= b and not a;
    layer3_outputs(3657) <= a;
    layer3_outputs(3658) <= not a;
    layer3_outputs(3659) <= not b;
    layer3_outputs(3660) <= a and b;
    layer3_outputs(3661) <= b;
    layer3_outputs(3662) <= a or b;
    layer3_outputs(3663) <= b and not a;
    layer3_outputs(3664) <= not b;
    layer3_outputs(3665) <= not a;
    layer3_outputs(3666) <= not b;
    layer3_outputs(3667) <= not (a and b);
    layer3_outputs(3668) <= not (a or b);
    layer3_outputs(3669) <= b;
    layer3_outputs(3670) <= a;
    layer3_outputs(3671) <= a;
    layer3_outputs(3672) <= b;
    layer3_outputs(3673) <= a or b;
    layer3_outputs(3674) <= b and not a;
    layer3_outputs(3675) <= b and not a;
    layer3_outputs(3676) <= not a or b;
    layer3_outputs(3677) <= a;
    layer3_outputs(3678) <= not a;
    layer3_outputs(3679) <= not (a xor b);
    layer3_outputs(3680) <= '1';
    layer3_outputs(3681) <= not (a and b);
    layer3_outputs(3682) <= not b;
    layer3_outputs(3683) <= not (a and b);
    layer3_outputs(3684) <= not b;
    layer3_outputs(3685) <= not (a or b);
    layer3_outputs(3686) <= a and not b;
    layer3_outputs(3687) <= not a;
    layer3_outputs(3688) <= not a;
    layer3_outputs(3689) <= not a;
    layer3_outputs(3690) <= not b;
    layer3_outputs(3691) <= a and b;
    layer3_outputs(3692) <= a xor b;
    layer3_outputs(3693) <= not (a or b);
    layer3_outputs(3694) <= a;
    layer3_outputs(3695) <= b and not a;
    layer3_outputs(3696) <= '1';
    layer3_outputs(3697) <= a;
    layer3_outputs(3698) <= not b;
    layer3_outputs(3699) <= not a;
    layer3_outputs(3700) <= not b;
    layer3_outputs(3701) <= not a or b;
    layer3_outputs(3702) <= not a;
    layer3_outputs(3703) <= '1';
    layer3_outputs(3704) <= a or b;
    layer3_outputs(3705) <= not a or b;
    layer3_outputs(3706) <= not (a or b);
    layer3_outputs(3707) <= not b or a;
    layer3_outputs(3708) <= a and b;
    layer3_outputs(3709) <= not (a or b);
    layer3_outputs(3710) <= a or b;
    layer3_outputs(3711) <= a;
    layer3_outputs(3712) <= not (a and b);
    layer3_outputs(3713) <= not (a xor b);
    layer3_outputs(3714) <= a and b;
    layer3_outputs(3715) <= a;
    layer3_outputs(3716) <= b;
    layer3_outputs(3717) <= not b or a;
    layer3_outputs(3718) <= a;
    layer3_outputs(3719) <= b;
    layer3_outputs(3720) <= b;
    layer3_outputs(3721) <= a and b;
    layer3_outputs(3722) <= not a;
    layer3_outputs(3723) <= a and b;
    layer3_outputs(3724) <= not (a or b);
    layer3_outputs(3725) <= not (a xor b);
    layer3_outputs(3726) <= a or b;
    layer3_outputs(3727) <= a;
    layer3_outputs(3728) <= '1';
    layer3_outputs(3729) <= b;
    layer3_outputs(3730) <= b;
    layer3_outputs(3731) <= not a or b;
    layer3_outputs(3732) <= not b or a;
    layer3_outputs(3733) <= not (a or b);
    layer3_outputs(3734) <= b;
    layer3_outputs(3735) <= a and not b;
    layer3_outputs(3736) <= not a or b;
    layer3_outputs(3737) <= b and not a;
    layer3_outputs(3738) <= not a or b;
    layer3_outputs(3739) <= a or b;
    layer3_outputs(3740) <= not (a xor b);
    layer3_outputs(3741) <= a and not b;
    layer3_outputs(3742) <= a and b;
    layer3_outputs(3743) <= a;
    layer3_outputs(3744) <= not (a xor b);
    layer3_outputs(3745) <= not (a or b);
    layer3_outputs(3746) <= b;
    layer3_outputs(3747) <= not b or a;
    layer3_outputs(3748) <= not (a and b);
    layer3_outputs(3749) <= not (a and b);
    layer3_outputs(3750) <= not (a and b);
    layer3_outputs(3751) <= not b;
    layer3_outputs(3752) <= not a or b;
    layer3_outputs(3753) <= not a or b;
    layer3_outputs(3754) <= not (a xor b);
    layer3_outputs(3755) <= not b;
    layer3_outputs(3756) <= a and b;
    layer3_outputs(3757) <= a;
    layer3_outputs(3758) <= a and not b;
    layer3_outputs(3759) <= not (a or b);
    layer3_outputs(3760) <= a;
    layer3_outputs(3761) <= not (a xor b);
    layer3_outputs(3762) <= a xor b;
    layer3_outputs(3763) <= b and not a;
    layer3_outputs(3764) <= b;
    layer3_outputs(3765) <= a xor b;
    layer3_outputs(3766) <= not a;
    layer3_outputs(3767) <= b;
    layer3_outputs(3768) <= b and not a;
    layer3_outputs(3769) <= b;
    layer3_outputs(3770) <= a and not b;
    layer3_outputs(3771) <= not (a and b);
    layer3_outputs(3772) <= not (a xor b);
    layer3_outputs(3773) <= not a or b;
    layer3_outputs(3774) <= a or b;
    layer3_outputs(3775) <= not b;
    layer3_outputs(3776) <= not (a or b);
    layer3_outputs(3777) <= b and not a;
    layer3_outputs(3778) <= not a;
    layer3_outputs(3779) <= a or b;
    layer3_outputs(3780) <= a or b;
    layer3_outputs(3781) <= not a or b;
    layer3_outputs(3782) <= not b;
    layer3_outputs(3783) <= not (a xor b);
    layer3_outputs(3784) <= a;
    layer3_outputs(3785) <= a and b;
    layer3_outputs(3786) <= b;
    layer3_outputs(3787) <= not b;
    layer3_outputs(3788) <= not b or a;
    layer3_outputs(3789) <= b and not a;
    layer3_outputs(3790) <= a xor b;
    layer3_outputs(3791) <= a and not b;
    layer3_outputs(3792) <= not (a or b);
    layer3_outputs(3793) <= '1';
    layer3_outputs(3794) <= not a or b;
    layer3_outputs(3795) <= a xor b;
    layer3_outputs(3796) <= a and not b;
    layer3_outputs(3797) <= not (a or b);
    layer3_outputs(3798) <= not a;
    layer3_outputs(3799) <= not b or a;
    layer3_outputs(3800) <= b and not a;
    layer3_outputs(3801) <= a and b;
    layer3_outputs(3802) <= a and not b;
    layer3_outputs(3803) <= a;
    layer3_outputs(3804) <= not a;
    layer3_outputs(3805) <= a and b;
    layer3_outputs(3806) <= a;
    layer3_outputs(3807) <= not b;
    layer3_outputs(3808) <= a xor b;
    layer3_outputs(3809) <= b;
    layer3_outputs(3810) <= a or b;
    layer3_outputs(3811) <= a or b;
    layer3_outputs(3812) <= a;
    layer3_outputs(3813) <= not a or b;
    layer3_outputs(3814) <= not b or a;
    layer3_outputs(3815) <= a and b;
    layer3_outputs(3816) <= a and not b;
    layer3_outputs(3817) <= a;
    layer3_outputs(3818) <= b;
    layer3_outputs(3819) <= not b;
    layer3_outputs(3820) <= not b;
    layer3_outputs(3821) <= b;
    layer3_outputs(3822) <= not a;
    layer3_outputs(3823) <= b;
    layer3_outputs(3824) <= a or b;
    layer3_outputs(3825) <= not a;
    layer3_outputs(3826) <= a and not b;
    layer3_outputs(3827) <= a and b;
    layer3_outputs(3828) <= b and not a;
    layer3_outputs(3829) <= not (a and b);
    layer3_outputs(3830) <= not b;
    layer3_outputs(3831) <= not (a or b);
    layer3_outputs(3832) <= a and not b;
    layer3_outputs(3833) <= not a;
    layer3_outputs(3834) <= a;
    layer3_outputs(3835) <= a or b;
    layer3_outputs(3836) <= '1';
    layer3_outputs(3837) <= b and not a;
    layer3_outputs(3838) <= not b;
    layer3_outputs(3839) <= not (a or b);
    layer3_outputs(3840) <= a and not b;
    layer3_outputs(3841) <= a;
    layer3_outputs(3842) <= not (a and b);
    layer3_outputs(3843) <= not a;
    layer3_outputs(3844) <= not b or a;
    layer3_outputs(3845) <= a xor b;
    layer3_outputs(3846) <= b;
    layer3_outputs(3847) <= a;
    layer3_outputs(3848) <= not (a or b);
    layer3_outputs(3849) <= not b or a;
    layer3_outputs(3850) <= a;
    layer3_outputs(3851) <= not (a xor b);
    layer3_outputs(3852) <= a and not b;
    layer3_outputs(3853) <= b;
    layer3_outputs(3854) <= not a;
    layer3_outputs(3855) <= not b;
    layer3_outputs(3856) <= not (a and b);
    layer3_outputs(3857) <= not (a and b);
    layer3_outputs(3858) <= not (a and b);
    layer3_outputs(3859) <= not a or b;
    layer3_outputs(3860) <= not a;
    layer3_outputs(3861) <= not (a xor b);
    layer3_outputs(3862) <= not a;
    layer3_outputs(3863) <= not a;
    layer3_outputs(3864) <= a xor b;
    layer3_outputs(3865) <= a xor b;
    layer3_outputs(3866) <= not b or a;
    layer3_outputs(3867) <= not b;
    layer3_outputs(3868) <= not a or b;
    layer3_outputs(3869) <= a;
    layer3_outputs(3870) <= not b or a;
    layer3_outputs(3871) <= b;
    layer3_outputs(3872) <= a;
    layer3_outputs(3873) <= not b;
    layer3_outputs(3874) <= not b;
    layer3_outputs(3875) <= not b;
    layer3_outputs(3876) <= a;
    layer3_outputs(3877) <= not a or b;
    layer3_outputs(3878) <= a;
    layer3_outputs(3879) <= not b;
    layer3_outputs(3880) <= a or b;
    layer3_outputs(3881) <= a and b;
    layer3_outputs(3882) <= not (a and b);
    layer3_outputs(3883) <= a or b;
    layer3_outputs(3884) <= not a or b;
    layer3_outputs(3885) <= not b or a;
    layer3_outputs(3886) <= b and not a;
    layer3_outputs(3887) <= a xor b;
    layer3_outputs(3888) <= not (a and b);
    layer3_outputs(3889) <= not b or a;
    layer3_outputs(3890) <= not b;
    layer3_outputs(3891) <= b and not a;
    layer3_outputs(3892) <= a or b;
    layer3_outputs(3893) <= '1';
    layer3_outputs(3894) <= b;
    layer3_outputs(3895) <= not (a or b);
    layer3_outputs(3896) <= not b or a;
    layer3_outputs(3897) <= not b;
    layer3_outputs(3898) <= not b;
    layer3_outputs(3899) <= not a;
    layer3_outputs(3900) <= not b;
    layer3_outputs(3901) <= b;
    layer3_outputs(3902) <= a and not b;
    layer3_outputs(3903) <= not a;
    layer3_outputs(3904) <= not b or a;
    layer3_outputs(3905) <= not (a or b);
    layer3_outputs(3906) <= b;
    layer3_outputs(3907) <= b and not a;
    layer3_outputs(3908) <= a and b;
    layer3_outputs(3909) <= b;
    layer3_outputs(3910) <= not b;
    layer3_outputs(3911) <= not a;
    layer3_outputs(3912) <= not b;
    layer3_outputs(3913) <= a;
    layer3_outputs(3914) <= a;
    layer3_outputs(3915) <= not (a xor b);
    layer3_outputs(3916) <= b;
    layer3_outputs(3917) <= not b or a;
    layer3_outputs(3918) <= not b;
    layer3_outputs(3919) <= not (a or b);
    layer3_outputs(3920) <= a and b;
    layer3_outputs(3921) <= not b or a;
    layer3_outputs(3922) <= not (a or b);
    layer3_outputs(3923) <= not (a and b);
    layer3_outputs(3924) <= a;
    layer3_outputs(3925) <= a or b;
    layer3_outputs(3926) <= '0';
    layer3_outputs(3927) <= not (a and b);
    layer3_outputs(3928) <= not (a xor b);
    layer3_outputs(3929) <= not (a xor b);
    layer3_outputs(3930) <= a xor b;
    layer3_outputs(3931) <= a xor b;
    layer3_outputs(3932) <= a;
    layer3_outputs(3933) <= a xor b;
    layer3_outputs(3934) <= not a or b;
    layer3_outputs(3935) <= not (a and b);
    layer3_outputs(3936) <= b;
    layer3_outputs(3937) <= not a;
    layer3_outputs(3938) <= a or b;
    layer3_outputs(3939) <= not (a xor b);
    layer3_outputs(3940) <= not a;
    layer3_outputs(3941) <= not a or b;
    layer3_outputs(3942) <= a and not b;
    layer3_outputs(3943) <= not a;
    layer3_outputs(3944) <= a xor b;
    layer3_outputs(3945) <= not (a and b);
    layer3_outputs(3946) <= '1';
    layer3_outputs(3947) <= a or b;
    layer3_outputs(3948) <= '0';
    layer3_outputs(3949) <= not a;
    layer3_outputs(3950) <= not b;
    layer3_outputs(3951) <= not b or a;
    layer3_outputs(3952) <= a;
    layer3_outputs(3953) <= b;
    layer3_outputs(3954) <= not a or b;
    layer3_outputs(3955) <= not b or a;
    layer3_outputs(3956) <= b;
    layer3_outputs(3957) <= not (a xor b);
    layer3_outputs(3958) <= not a;
    layer3_outputs(3959) <= a and b;
    layer3_outputs(3960) <= not b or a;
    layer3_outputs(3961) <= a;
    layer3_outputs(3962) <= a;
    layer3_outputs(3963) <= not (a or b);
    layer3_outputs(3964) <= not (a or b);
    layer3_outputs(3965) <= b;
    layer3_outputs(3966) <= '0';
    layer3_outputs(3967) <= a;
    layer3_outputs(3968) <= not (a xor b);
    layer3_outputs(3969) <= a xor b;
    layer3_outputs(3970) <= not a or b;
    layer3_outputs(3971) <= not (a and b);
    layer3_outputs(3972) <= not b;
    layer3_outputs(3973) <= not (a or b);
    layer3_outputs(3974) <= b;
    layer3_outputs(3975) <= a and not b;
    layer3_outputs(3976) <= not a;
    layer3_outputs(3977) <= a;
    layer3_outputs(3978) <= not b or a;
    layer3_outputs(3979) <= a and not b;
    layer3_outputs(3980) <= '0';
    layer3_outputs(3981) <= not a or b;
    layer3_outputs(3982) <= a;
    layer3_outputs(3983) <= not a or b;
    layer3_outputs(3984) <= not a;
    layer3_outputs(3985) <= not b;
    layer3_outputs(3986) <= not a;
    layer3_outputs(3987) <= not (a and b);
    layer3_outputs(3988) <= not (a and b);
    layer3_outputs(3989) <= not (a and b);
    layer3_outputs(3990) <= '0';
    layer3_outputs(3991) <= b;
    layer3_outputs(3992) <= not b;
    layer3_outputs(3993) <= a or b;
    layer3_outputs(3994) <= not a;
    layer3_outputs(3995) <= b and not a;
    layer3_outputs(3996) <= a;
    layer3_outputs(3997) <= b;
    layer3_outputs(3998) <= not b;
    layer3_outputs(3999) <= not b or a;
    layer3_outputs(4000) <= not a;
    layer3_outputs(4001) <= not (a or b);
    layer3_outputs(4002) <= not (a and b);
    layer3_outputs(4003) <= a and not b;
    layer3_outputs(4004) <= not (a xor b);
    layer3_outputs(4005) <= a xor b;
    layer3_outputs(4006) <= not b or a;
    layer3_outputs(4007) <= a and b;
    layer3_outputs(4008) <= b;
    layer3_outputs(4009) <= not b;
    layer3_outputs(4010) <= not b;
    layer3_outputs(4011) <= '0';
    layer3_outputs(4012) <= a or b;
    layer3_outputs(4013) <= a or b;
    layer3_outputs(4014) <= not a;
    layer3_outputs(4015) <= a xor b;
    layer3_outputs(4016) <= b and not a;
    layer3_outputs(4017) <= not a;
    layer3_outputs(4018) <= not a or b;
    layer3_outputs(4019) <= not a;
    layer3_outputs(4020) <= not b or a;
    layer3_outputs(4021) <= not b or a;
    layer3_outputs(4022) <= not (a and b);
    layer3_outputs(4023) <= b;
    layer3_outputs(4024) <= not b;
    layer3_outputs(4025) <= not (a xor b);
    layer3_outputs(4026) <= not a or b;
    layer3_outputs(4027) <= not (a xor b);
    layer3_outputs(4028) <= a or b;
    layer3_outputs(4029) <= not b;
    layer3_outputs(4030) <= not b;
    layer3_outputs(4031) <= not a;
    layer3_outputs(4032) <= not b or a;
    layer3_outputs(4033) <= a xor b;
    layer3_outputs(4034) <= not a or b;
    layer3_outputs(4035) <= a and b;
    layer3_outputs(4036) <= not b;
    layer3_outputs(4037) <= b;
    layer3_outputs(4038) <= a;
    layer3_outputs(4039) <= not (a and b);
    layer3_outputs(4040) <= a;
    layer3_outputs(4041) <= '1';
    layer3_outputs(4042) <= b and not a;
    layer3_outputs(4043) <= not a;
    layer3_outputs(4044) <= a and b;
    layer3_outputs(4045) <= b;
    layer3_outputs(4046) <= a;
    layer3_outputs(4047) <= a and b;
    layer3_outputs(4048) <= a;
    layer3_outputs(4049) <= a;
    layer3_outputs(4050) <= not (a or b);
    layer3_outputs(4051) <= not a;
    layer3_outputs(4052) <= a and not b;
    layer3_outputs(4053) <= a xor b;
    layer3_outputs(4054) <= not a or b;
    layer3_outputs(4055) <= not a;
    layer3_outputs(4056) <= not a or b;
    layer3_outputs(4057) <= not (a and b);
    layer3_outputs(4058) <= not b or a;
    layer3_outputs(4059) <= not b;
    layer3_outputs(4060) <= '0';
    layer3_outputs(4061) <= not a;
    layer3_outputs(4062) <= a and not b;
    layer3_outputs(4063) <= '0';
    layer3_outputs(4064) <= not a or b;
    layer3_outputs(4065) <= a and not b;
    layer3_outputs(4066) <= a and not b;
    layer3_outputs(4067) <= not (a or b);
    layer3_outputs(4068) <= not b or a;
    layer3_outputs(4069) <= not b;
    layer3_outputs(4070) <= a and b;
    layer3_outputs(4071) <= not (a or b);
    layer3_outputs(4072) <= a or b;
    layer3_outputs(4073) <= a and not b;
    layer3_outputs(4074) <= not b or a;
    layer3_outputs(4075) <= b;
    layer3_outputs(4076) <= not (a xor b);
    layer3_outputs(4077) <= not a;
    layer3_outputs(4078) <= not b;
    layer3_outputs(4079) <= a and b;
    layer3_outputs(4080) <= not b;
    layer3_outputs(4081) <= not b or a;
    layer3_outputs(4082) <= a xor b;
    layer3_outputs(4083) <= not b or a;
    layer3_outputs(4084) <= not a or b;
    layer3_outputs(4085) <= b;
    layer3_outputs(4086) <= not a;
    layer3_outputs(4087) <= not a;
    layer3_outputs(4088) <= b;
    layer3_outputs(4089) <= a;
    layer3_outputs(4090) <= not (a and b);
    layer3_outputs(4091) <= b and not a;
    layer3_outputs(4092) <= not b;
    layer3_outputs(4093) <= a or b;
    layer3_outputs(4094) <= a;
    layer3_outputs(4095) <= not (a and b);
    layer3_outputs(4096) <= not b;
    layer3_outputs(4097) <= not a;
    layer3_outputs(4098) <= not a or b;
    layer3_outputs(4099) <= not b;
    layer3_outputs(4100) <= a xor b;
    layer3_outputs(4101) <= not a or b;
    layer3_outputs(4102) <= a or b;
    layer3_outputs(4103) <= a;
    layer3_outputs(4104) <= not (a or b);
    layer3_outputs(4105) <= not a;
    layer3_outputs(4106) <= not (a or b);
    layer3_outputs(4107) <= b and not a;
    layer3_outputs(4108) <= not b;
    layer3_outputs(4109) <= not a or b;
    layer3_outputs(4110) <= not b;
    layer3_outputs(4111) <= not b;
    layer3_outputs(4112) <= a xor b;
    layer3_outputs(4113) <= b;
    layer3_outputs(4114) <= not (a or b);
    layer3_outputs(4115) <= not b;
    layer3_outputs(4116) <= b;
    layer3_outputs(4117) <= not a or b;
    layer3_outputs(4118) <= not b;
    layer3_outputs(4119) <= not b;
    layer3_outputs(4120) <= a;
    layer3_outputs(4121) <= b and not a;
    layer3_outputs(4122) <= not b;
    layer3_outputs(4123) <= b and not a;
    layer3_outputs(4124) <= a and not b;
    layer3_outputs(4125) <= '1';
    layer3_outputs(4126) <= not a;
    layer3_outputs(4127) <= a and b;
    layer3_outputs(4128) <= not b or a;
    layer3_outputs(4129) <= a or b;
    layer3_outputs(4130) <= not b or a;
    layer3_outputs(4131) <= not a or b;
    layer3_outputs(4132) <= not b or a;
    layer3_outputs(4133) <= not (a or b);
    layer3_outputs(4134) <= a and b;
    layer3_outputs(4135) <= not b or a;
    layer3_outputs(4136) <= '1';
    layer3_outputs(4137) <= a xor b;
    layer3_outputs(4138) <= a;
    layer3_outputs(4139) <= b;
    layer3_outputs(4140) <= a or b;
    layer3_outputs(4141) <= not b;
    layer3_outputs(4142) <= a;
    layer3_outputs(4143) <= not a;
    layer3_outputs(4144) <= a or b;
    layer3_outputs(4145) <= not (a or b);
    layer3_outputs(4146) <= not (a and b);
    layer3_outputs(4147) <= not b or a;
    layer3_outputs(4148) <= not (a and b);
    layer3_outputs(4149) <= a and not b;
    layer3_outputs(4150) <= a or b;
    layer3_outputs(4151) <= '0';
    layer3_outputs(4152) <= not b;
    layer3_outputs(4153) <= b;
    layer3_outputs(4154) <= b and not a;
    layer3_outputs(4155) <= not a or b;
    layer3_outputs(4156) <= not a;
    layer3_outputs(4157) <= b;
    layer3_outputs(4158) <= a and not b;
    layer3_outputs(4159) <= a xor b;
    layer3_outputs(4160) <= not (a xor b);
    layer3_outputs(4161) <= a or b;
    layer3_outputs(4162) <= not (a xor b);
    layer3_outputs(4163) <= a and b;
    layer3_outputs(4164) <= not a;
    layer3_outputs(4165) <= not a or b;
    layer3_outputs(4166) <= not a;
    layer3_outputs(4167) <= not a;
    layer3_outputs(4168) <= not b;
    layer3_outputs(4169) <= a;
    layer3_outputs(4170) <= a;
    layer3_outputs(4171) <= a and b;
    layer3_outputs(4172) <= not a or b;
    layer3_outputs(4173) <= b;
    layer3_outputs(4174) <= not a or b;
    layer3_outputs(4175) <= not (a or b);
    layer3_outputs(4176) <= '1';
    layer3_outputs(4177) <= '0';
    layer3_outputs(4178) <= not a;
    layer3_outputs(4179) <= b and not a;
    layer3_outputs(4180) <= a and not b;
    layer3_outputs(4181) <= not a;
    layer3_outputs(4182) <= not (a xor b);
    layer3_outputs(4183) <= not a;
    layer3_outputs(4184) <= a or b;
    layer3_outputs(4185) <= a;
    layer3_outputs(4186) <= not b;
    layer3_outputs(4187) <= a and b;
    layer3_outputs(4188) <= not b or a;
    layer3_outputs(4189) <= not a or b;
    layer3_outputs(4190) <= not (a or b);
    layer3_outputs(4191) <= not (a or b);
    layer3_outputs(4192) <= a;
    layer3_outputs(4193) <= not b;
    layer3_outputs(4194) <= not (a xor b);
    layer3_outputs(4195) <= not (a or b);
    layer3_outputs(4196) <= not (a or b);
    layer3_outputs(4197) <= not a;
    layer3_outputs(4198) <= not (a and b);
    layer3_outputs(4199) <= not (a and b);
    layer3_outputs(4200) <= a xor b;
    layer3_outputs(4201) <= not b or a;
    layer3_outputs(4202) <= b and not a;
    layer3_outputs(4203) <= a xor b;
    layer3_outputs(4204) <= b;
    layer3_outputs(4205) <= b;
    layer3_outputs(4206) <= not (a xor b);
    layer3_outputs(4207) <= a or b;
    layer3_outputs(4208) <= a and not b;
    layer3_outputs(4209) <= b;
    layer3_outputs(4210) <= b;
    layer3_outputs(4211) <= not a or b;
    layer3_outputs(4212) <= a and b;
    layer3_outputs(4213) <= not (a and b);
    layer3_outputs(4214) <= b;
    layer3_outputs(4215) <= not (a and b);
    layer3_outputs(4216) <= a and b;
    layer3_outputs(4217) <= not (a xor b);
    layer3_outputs(4218) <= a;
    layer3_outputs(4219) <= b and not a;
    layer3_outputs(4220) <= not b;
    layer3_outputs(4221) <= a or b;
    layer3_outputs(4222) <= not (a and b);
    layer3_outputs(4223) <= b and not a;
    layer3_outputs(4224) <= a xor b;
    layer3_outputs(4225) <= not b;
    layer3_outputs(4226) <= b and not a;
    layer3_outputs(4227) <= not a;
    layer3_outputs(4228) <= not (a or b);
    layer3_outputs(4229) <= b and not a;
    layer3_outputs(4230) <= '0';
    layer3_outputs(4231) <= not b;
    layer3_outputs(4232) <= not b;
    layer3_outputs(4233) <= not b or a;
    layer3_outputs(4234) <= not (a xor b);
    layer3_outputs(4235) <= not a or b;
    layer3_outputs(4236) <= b;
    layer3_outputs(4237) <= not a or b;
    layer3_outputs(4238) <= not b;
    layer3_outputs(4239) <= a;
    layer3_outputs(4240) <= b and not a;
    layer3_outputs(4241) <= not a or b;
    layer3_outputs(4242) <= '1';
    layer3_outputs(4243) <= b and not a;
    layer3_outputs(4244) <= not a or b;
    layer3_outputs(4245) <= b;
    layer3_outputs(4246) <= not b or a;
    layer3_outputs(4247) <= not a or b;
    layer3_outputs(4248) <= not b or a;
    layer3_outputs(4249) <= a and not b;
    layer3_outputs(4250) <= not a or b;
    layer3_outputs(4251) <= a;
    layer3_outputs(4252) <= not a;
    layer3_outputs(4253) <= not (a xor b);
    layer3_outputs(4254) <= b and not a;
    layer3_outputs(4255) <= not (a or b);
    layer3_outputs(4256) <= a and b;
    layer3_outputs(4257) <= not b or a;
    layer3_outputs(4258) <= a and b;
    layer3_outputs(4259) <= a;
    layer3_outputs(4260) <= not (a and b);
    layer3_outputs(4261) <= not (a or b);
    layer3_outputs(4262) <= b;
    layer3_outputs(4263) <= a or b;
    layer3_outputs(4264) <= b;
    layer3_outputs(4265) <= a;
    layer3_outputs(4266) <= a;
    layer3_outputs(4267) <= not (a or b);
    layer3_outputs(4268) <= b;
    layer3_outputs(4269) <= not a or b;
    layer3_outputs(4270) <= a;
    layer3_outputs(4271) <= b and not a;
    layer3_outputs(4272) <= not a;
    layer3_outputs(4273) <= a and not b;
    layer3_outputs(4274) <= not a;
    layer3_outputs(4275) <= a and not b;
    layer3_outputs(4276) <= a or b;
    layer3_outputs(4277) <= not b or a;
    layer3_outputs(4278) <= b;
    layer3_outputs(4279) <= not a or b;
    layer3_outputs(4280) <= a or b;
    layer3_outputs(4281) <= not (a xor b);
    layer3_outputs(4282) <= not b or a;
    layer3_outputs(4283) <= not a;
    layer3_outputs(4284) <= a;
    layer3_outputs(4285) <= a xor b;
    layer3_outputs(4286) <= a;
    layer3_outputs(4287) <= b;
    layer3_outputs(4288) <= not a;
    layer3_outputs(4289) <= not b;
    layer3_outputs(4290) <= a;
    layer3_outputs(4291) <= not a;
    layer3_outputs(4292) <= not b;
    layer3_outputs(4293) <= b;
    layer3_outputs(4294) <= not a;
    layer3_outputs(4295) <= a xor b;
    layer3_outputs(4296) <= a and not b;
    layer3_outputs(4297) <= a xor b;
    layer3_outputs(4298) <= b;
    layer3_outputs(4299) <= b;
    layer3_outputs(4300) <= not b or a;
    layer3_outputs(4301) <= not (a xor b);
    layer3_outputs(4302) <= a or b;
    layer3_outputs(4303) <= not b or a;
    layer3_outputs(4304) <= not a or b;
    layer3_outputs(4305) <= b and not a;
    layer3_outputs(4306) <= not b or a;
    layer3_outputs(4307) <= a xor b;
    layer3_outputs(4308) <= not b;
    layer3_outputs(4309) <= a;
    layer3_outputs(4310) <= a and b;
    layer3_outputs(4311) <= not (a and b);
    layer3_outputs(4312) <= not (a or b);
    layer3_outputs(4313) <= a or b;
    layer3_outputs(4314) <= a and not b;
    layer3_outputs(4315) <= a and not b;
    layer3_outputs(4316) <= not b or a;
    layer3_outputs(4317) <= not a or b;
    layer3_outputs(4318) <= not a or b;
    layer3_outputs(4319) <= not b;
    layer3_outputs(4320) <= not a;
    layer3_outputs(4321) <= not b or a;
    layer3_outputs(4322) <= a;
    layer3_outputs(4323) <= a;
    layer3_outputs(4324) <= not (a xor b);
    layer3_outputs(4325) <= not b;
    layer3_outputs(4326) <= a and not b;
    layer3_outputs(4327) <= not a;
    layer3_outputs(4328) <= not (a xor b);
    layer3_outputs(4329) <= b;
    layer3_outputs(4330) <= not b;
    layer3_outputs(4331) <= not (a or b);
    layer3_outputs(4332) <= b;
    layer3_outputs(4333) <= a;
    layer3_outputs(4334) <= b;
    layer3_outputs(4335) <= b;
    layer3_outputs(4336) <= not (a or b);
    layer3_outputs(4337) <= b;
    layer3_outputs(4338) <= a and b;
    layer3_outputs(4339) <= not b;
    layer3_outputs(4340) <= b;
    layer3_outputs(4341) <= a;
    layer3_outputs(4342) <= not (a or b);
    layer3_outputs(4343) <= a xor b;
    layer3_outputs(4344) <= a;
    layer3_outputs(4345) <= not (a or b);
    layer3_outputs(4346) <= not b or a;
    layer3_outputs(4347) <= a;
    layer3_outputs(4348) <= a or b;
    layer3_outputs(4349) <= not b;
    layer3_outputs(4350) <= a xor b;
    layer3_outputs(4351) <= not (a or b);
    layer3_outputs(4352) <= not b;
    layer3_outputs(4353) <= not b;
    layer3_outputs(4354) <= not (a or b);
    layer3_outputs(4355) <= not (a and b);
    layer3_outputs(4356) <= not (a and b);
    layer3_outputs(4357) <= not a;
    layer3_outputs(4358) <= not b;
    layer3_outputs(4359) <= a or b;
    layer3_outputs(4360) <= b;
    layer3_outputs(4361) <= b and not a;
    layer3_outputs(4362) <= not (a and b);
    layer3_outputs(4363) <= b and not a;
    layer3_outputs(4364) <= b and not a;
    layer3_outputs(4365) <= a or b;
    layer3_outputs(4366) <= not (a and b);
    layer3_outputs(4367) <= a and not b;
    layer3_outputs(4368) <= not a;
    layer3_outputs(4369) <= not a;
    layer3_outputs(4370) <= not a or b;
    layer3_outputs(4371) <= b;
    layer3_outputs(4372) <= not (a and b);
    layer3_outputs(4373) <= b and not a;
    layer3_outputs(4374) <= not b or a;
    layer3_outputs(4375) <= not b or a;
    layer3_outputs(4376) <= a;
    layer3_outputs(4377) <= b;
    layer3_outputs(4378) <= not (a or b);
    layer3_outputs(4379) <= a;
    layer3_outputs(4380) <= a;
    layer3_outputs(4381) <= b;
    layer3_outputs(4382) <= '1';
    layer3_outputs(4383) <= not (a xor b);
    layer3_outputs(4384) <= not (a and b);
    layer3_outputs(4385) <= a and not b;
    layer3_outputs(4386) <= not a;
    layer3_outputs(4387) <= a;
    layer3_outputs(4388) <= not (a or b);
    layer3_outputs(4389) <= b and not a;
    layer3_outputs(4390) <= b;
    layer3_outputs(4391) <= not a;
    layer3_outputs(4392) <= '1';
    layer3_outputs(4393) <= not b;
    layer3_outputs(4394) <= b;
    layer3_outputs(4395) <= not a or b;
    layer3_outputs(4396) <= not b;
    layer3_outputs(4397) <= a and b;
    layer3_outputs(4398) <= b and not a;
    layer3_outputs(4399) <= b and not a;
    layer3_outputs(4400) <= not b;
    layer3_outputs(4401) <= not b;
    layer3_outputs(4402) <= not a;
    layer3_outputs(4403) <= not b;
    layer3_outputs(4404) <= b;
    layer3_outputs(4405) <= not b or a;
    layer3_outputs(4406) <= not a or b;
    layer3_outputs(4407) <= a or b;
    layer3_outputs(4408) <= not (a and b);
    layer3_outputs(4409) <= not (a xor b);
    layer3_outputs(4410) <= not b;
    layer3_outputs(4411) <= b and not a;
    layer3_outputs(4412) <= not (a or b);
    layer3_outputs(4413) <= a xor b;
    layer3_outputs(4414) <= not (a or b);
    layer3_outputs(4415) <= not a or b;
    layer3_outputs(4416) <= a;
    layer3_outputs(4417) <= a and b;
    layer3_outputs(4418) <= not b or a;
    layer3_outputs(4419) <= a and not b;
    layer3_outputs(4420) <= not (a and b);
    layer3_outputs(4421) <= a;
    layer3_outputs(4422) <= not a;
    layer3_outputs(4423) <= a and not b;
    layer3_outputs(4424) <= b;
    layer3_outputs(4425) <= not b;
    layer3_outputs(4426) <= not a or b;
    layer3_outputs(4427) <= a;
    layer3_outputs(4428) <= not (a xor b);
    layer3_outputs(4429) <= a xor b;
    layer3_outputs(4430) <= not b or a;
    layer3_outputs(4431) <= not (a xor b);
    layer3_outputs(4432) <= not b;
    layer3_outputs(4433) <= not b or a;
    layer3_outputs(4434) <= '0';
    layer3_outputs(4435) <= a;
    layer3_outputs(4436) <= a;
    layer3_outputs(4437) <= not a or b;
    layer3_outputs(4438) <= a and not b;
    layer3_outputs(4439) <= a xor b;
    layer3_outputs(4440) <= not (a or b);
    layer3_outputs(4441) <= not (a and b);
    layer3_outputs(4442) <= b;
    layer3_outputs(4443) <= not a or b;
    layer3_outputs(4444) <= not b or a;
    layer3_outputs(4445) <= not b;
    layer3_outputs(4446) <= a or b;
    layer3_outputs(4447) <= not a;
    layer3_outputs(4448) <= a and not b;
    layer3_outputs(4449) <= a and not b;
    layer3_outputs(4450) <= b and not a;
    layer3_outputs(4451) <= b and not a;
    layer3_outputs(4452) <= b and not a;
    layer3_outputs(4453) <= b;
    layer3_outputs(4454) <= not a;
    layer3_outputs(4455) <= a;
    layer3_outputs(4456) <= not (a or b);
    layer3_outputs(4457) <= not a;
    layer3_outputs(4458) <= b;
    layer3_outputs(4459) <= not a;
    layer3_outputs(4460) <= not (a and b);
    layer3_outputs(4461) <= not b;
    layer3_outputs(4462) <= not b or a;
    layer3_outputs(4463) <= a;
    layer3_outputs(4464) <= b;
    layer3_outputs(4465) <= not (a and b);
    layer3_outputs(4466) <= b and not a;
    layer3_outputs(4467) <= not b;
    layer3_outputs(4468) <= not b;
    layer3_outputs(4469) <= a and b;
    layer3_outputs(4470) <= not (a or b);
    layer3_outputs(4471) <= b and not a;
    layer3_outputs(4472) <= not (a or b);
    layer3_outputs(4473) <= not (a xor b);
    layer3_outputs(4474) <= not b or a;
    layer3_outputs(4475) <= not a;
    layer3_outputs(4476) <= b;
    layer3_outputs(4477) <= a;
    layer3_outputs(4478) <= not a;
    layer3_outputs(4479) <= a;
    layer3_outputs(4480) <= b;
    layer3_outputs(4481) <= a and not b;
    layer3_outputs(4482) <= a xor b;
    layer3_outputs(4483) <= not a;
    layer3_outputs(4484) <= not (a and b);
    layer3_outputs(4485) <= not a or b;
    layer3_outputs(4486) <= not a;
    layer3_outputs(4487) <= a xor b;
    layer3_outputs(4488) <= not a;
    layer3_outputs(4489) <= a and not b;
    layer3_outputs(4490) <= not a;
    layer3_outputs(4491) <= not a;
    layer3_outputs(4492) <= a and b;
    layer3_outputs(4493) <= not (a or b);
    layer3_outputs(4494) <= a and b;
    layer3_outputs(4495) <= not a or b;
    layer3_outputs(4496) <= a and b;
    layer3_outputs(4497) <= a or b;
    layer3_outputs(4498) <= a or b;
    layer3_outputs(4499) <= a xor b;
    layer3_outputs(4500) <= not a;
    layer3_outputs(4501) <= not b;
    layer3_outputs(4502) <= b;
    layer3_outputs(4503) <= not b;
    layer3_outputs(4504) <= b;
    layer3_outputs(4505) <= not b;
    layer3_outputs(4506) <= a;
    layer3_outputs(4507) <= not b or a;
    layer3_outputs(4508) <= '0';
    layer3_outputs(4509) <= not a or b;
    layer3_outputs(4510) <= not b or a;
    layer3_outputs(4511) <= a and not b;
    layer3_outputs(4512) <= not a;
    layer3_outputs(4513) <= not b;
    layer3_outputs(4514) <= b;
    layer3_outputs(4515) <= not a or b;
    layer3_outputs(4516) <= a;
    layer3_outputs(4517) <= not (a and b);
    layer3_outputs(4518) <= b;
    layer3_outputs(4519) <= not b;
    layer3_outputs(4520) <= b;
    layer3_outputs(4521) <= not (a or b);
    layer3_outputs(4522) <= a and not b;
    layer3_outputs(4523) <= '1';
    layer3_outputs(4524) <= not b;
    layer3_outputs(4525) <= not (a xor b);
    layer3_outputs(4526) <= not a;
    layer3_outputs(4527) <= not b;
    layer3_outputs(4528) <= a and b;
    layer3_outputs(4529) <= not a or b;
    layer3_outputs(4530) <= a or b;
    layer3_outputs(4531) <= not (a or b);
    layer3_outputs(4532) <= not a;
    layer3_outputs(4533) <= not (a or b);
    layer3_outputs(4534) <= a or b;
    layer3_outputs(4535) <= not a;
    layer3_outputs(4536) <= not b or a;
    layer3_outputs(4537) <= a;
    layer3_outputs(4538) <= a xor b;
    layer3_outputs(4539) <= a;
    layer3_outputs(4540) <= a xor b;
    layer3_outputs(4541) <= not a or b;
    layer3_outputs(4542) <= a or b;
    layer3_outputs(4543) <= not (a xor b);
    layer3_outputs(4544) <= not b;
    layer3_outputs(4545) <= a;
    layer3_outputs(4546) <= a xor b;
    layer3_outputs(4547) <= not a;
    layer3_outputs(4548) <= a;
    layer3_outputs(4549) <= b and not a;
    layer3_outputs(4550) <= b;
    layer3_outputs(4551) <= not (a and b);
    layer3_outputs(4552) <= not b or a;
    layer3_outputs(4553) <= not b;
    layer3_outputs(4554) <= a and b;
    layer3_outputs(4555) <= not (a and b);
    layer3_outputs(4556) <= not a;
    layer3_outputs(4557) <= a and not b;
    layer3_outputs(4558) <= b;
    layer3_outputs(4559) <= b;
    layer3_outputs(4560) <= b and not a;
    layer3_outputs(4561) <= not a;
    layer3_outputs(4562) <= not (a or b);
    layer3_outputs(4563) <= not b or a;
    layer3_outputs(4564) <= a and b;
    layer3_outputs(4565) <= not (a xor b);
    layer3_outputs(4566) <= not (a xor b);
    layer3_outputs(4567) <= '1';
    layer3_outputs(4568) <= not a or b;
    layer3_outputs(4569) <= not (a xor b);
    layer3_outputs(4570) <= not b or a;
    layer3_outputs(4571) <= a xor b;
    layer3_outputs(4572) <= a or b;
    layer3_outputs(4573) <= '1';
    layer3_outputs(4574) <= not a;
    layer3_outputs(4575) <= not b or a;
    layer3_outputs(4576) <= '1';
    layer3_outputs(4577) <= not b or a;
    layer3_outputs(4578) <= not (a and b);
    layer3_outputs(4579) <= a and not b;
    layer3_outputs(4580) <= b;
    layer3_outputs(4581) <= a and not b;
    layer3_outputs(4582) <= a;
    layer3_outputs(4583) <= not b or a;
    layer3_outputs(4584) <= b and not a;
    layer3_outputs(4585) <= a and b;
    layer3_outputs(4586) <= not (a or b);
    layer3_outputs(4587) <= a and not b;
    layer3_outputs(4588) <= not (a xor b);
    layer3_outputs(4589) <= '0';
    layer3_outputs(4590) <= a and b;
    layer3_outputs(4591) <= not b;
    layer3_outputs(4592) <= not a;
    layer3_outputs(4593) <= b;
    layer3_outputs(4594) <= a and b;
    layer3_outputs(4595) <= a and not b;
    layer3_outputs(4596) <= b;
    layer3_outputs(4597) <= not b or a;
    layer3_outputs(4598) <= a xor b;
    layer3_outputs(4599) <= not a;
    layer3_outputs(4600) <= not a or b;
    layer3_outputs(4601) <= not a or b;
    layer3_outputs(4602) <= b;
    layer3_outputs(4603) <= not b or a;
    layer3_outputs(4604) <= not a or b;
    layer3_outputs(4605) <= '0';
    layer3_outputs(4606) <= a;
    layer3_outputs(4607) <= a and not b;
    layer3_outputs(4608) <= not (a and b);
    layer3_outputs(4609) <= a or b;
    layer3_outputs(4610) <= a xor b;
    layer3_outputs(4611) <= not b;
    layer3_outputs(4612) <= not b;
    layer3_outputs(4613) <= b;
    layer3_outputs(4614) <= not (a or b);
    layer3_outputs(4615) <= a xor b;
    layer3_outputs(4616) <= not b;
    layer3_outputs(4617) <= '0';
    layer3_outputs(4618) <= not a;
    layer3_outputs(4619) <= a xor b;
    layer3_outputs(4620) <= a;
    layer3_outputs(4621) <= b and not a;
    layer3_outputs(4622) <= '0';
    layer3_outputs(4623) <= b;
    layer3_outputs(4624) <= not b or a;
    layer3_outputs(4625) <= not b or a;
    layer3_outputs(4626) <= a;
    layer3_outputs(4627) <= '0';
    layer3_outputs(4628) <= not a;
    layer3_outputs(4629) <= not a;
    layer3_outputs(4630) <= not (a or b);
    layer3_outputs(4631) <= a;
    layer3_outputs(4632) <= not a;
    layer3_outputs(4633) <= not b;
    layer3_outputs(4634) <= a and not b;
    layer3_outputs(4635) <= not b or a;
    layer3_outputs(4636) <= '0';
    layer3_outputs(4637) <= not (a xor b);
    layer3_outputs(4638) <= b and not a;
    layer3_outputs(4639) <= not b;
    layer3_outputs(4640) <= not (a or b);
    layer3_outputs(4641) <= a xor b;
    layer3_outputs(4642) <= a;
    layer3_outputs(4643) <= not b;
    layer3_outputs(4644) <= not a or b;
    layer3_outputs(4645) <= b and not a;
    layer3_outputs(4646) <= not b;
    layer3_outputs(4647) <= b;
    layer3_outputs(4648) <= a;
    layer3_outputs(4649) <= '1';
    layer3_outputs(4650) <= not (a xor b);
    layer3_outputs(4651) <= not a;
    layer3_outputs(4652) <= b;
    layer3_outputs(4653) <= a;
    layer3_outputs(4654) <= not a or b;
    layer3_outputs(4655) <= a xor b;
    layer3_outputs(4656) <= not a;
    layer3_outputs(4657) <= not a;
    layer3_outputs(4658) <= not b;
    layer3_outputs(4659) <= not b;
    layer3_outputs(4660) <= b;
    layer3_outputs(4661) <= a and not b;
    layer3_outputs(4662) <= not a;
    layer3_outputs(4663) <= b and not a;
    layer3_outputs(4664) <= not a;
    layer3_outputs(4665) <= a or b;
    layer3_outputs(4666) <= b;
    layer3_outputs(4667) <= a;
    layer3_outputs(4668) <= not (a or b);
    layer3_outputs(4669) <= a or b;
    layer3_outputs(4670) <= not a or b;
    layer3_outputs(4671) <= not (a and b);
    layer3_outputs(4672) <= a or b;
    layer3_outputs(4673) <= not b;
    layer3_outputs(4674) <= a;
    layer3_outputs(4675) <= not b or a;
    layer3_outputs(4676) <= not b;
    layer3_outputs(4677) <= not b;
    layer3_outputs(4678) <= not a;
    layer3_outputs(4679) <= a or b;
    layer3_outputs(4680) <= not a;
    layer3_outputs(4681) <= a xor b;
    layer3_outputs(4682) <= not b;
    layer3_outputs(4683) <= not b;
    layer3_outputs(4684) <= not a;
    layer3_outputs(4685) <= b and not a;
    layer3_outputs(4686) <= not (a xor b);
    layer3_outputs(4687) <= not b;
    layer3_outputs(4688) <= not b or a;
    layer3_outputs(4689) <= not a;
    layer3_outputs(4690) <= a xor b;
    layer3_outputs(4691) <= a;
    layer3_outputs(4692) <= not b;
    layer3_outputs(4693) <= not (a and b);
    layer3_outputs(4694) <= not b;
    layer3_outputs(4695) <= not b;
    layer3_outputs(4696) <= a xor b;
    layer3_outputs(4697) <= not (a xor b);
    layer3_outputs(4698) <= '1';
    layer3_outputs(4699) <= a;
    layer3_outputs(4700) <= '0';
    layer3_outputs(4701) <= a or b;
    layer3_outputs(4702) <= a and b;
    layer3_outputs(4703) <= not b;
    layer3_outputs(4704) <= b;
    layer3_outputs(4705) <= not b;
    layer3_outputs(4706) <= not (a and b);
    layer3_outputs(4707) <= a and b;
    layer3_outputs(4708) <= not (a and b);
    layer3_outputs(4709) <= not b;
    layer3_outputs(4710) <= not a;
    layer3_outputs(4711) <= b and not a;
    layer3_outputs(4712) <= not (a or b);
    layer3_outputs(4713) <= not b or a;
    layer3_outputs(4714) <= not b;
    layer3_outputs(4715) <= b;
    layer3_outputs(4716) <= a and b;
    layer3_outputs(4717) <= b and not a;
    layer3_outputs(4718) <= a or b;
    layer3_outputs(4719) <= b and not a;
    layer3_outputs(4720) <= b and not a;
    layer3_outputs(4721) <= a;
    layer3_outputs(4722) <= a;
    layer3_outputs(4723) <= not (a xor b);
    layer3_outputs(4724) <= not b or a;
    layer3_outputs(4725) <= not (a and b);
    layer3_outputs(4726) <= not a;
    layer3_outputs(4727) <= b;
    layer3_outputs(4728) <= a;
    layer3_outputs(4729) <= a and b;
    layer3_outputs(4730) <= b;
    layer3_outputs(4731) <= a or b;
    layer3_outputs(4732) <= b;
    layer3_outputs(4733) <= b;
    layer3_outputs(4734) <= a;
    layer3_outputs(4735) <= a xor b;
    layer3_outputs(4736) <= not (a and b);
    layer3_outputs(4737) <= a;
    layer3_outputs(4738) <= b;
    layer3_outputs(4739) <= b;
    layer3_outputs(4740) <= not (a and b);
    layer3_outputs(4741) <= not a;
    layer3_outputs(4742) <= a;
    layer3_outputs(4743) <= not b or a;
    layer3_outputs(4744) <= not b;
    layer3_outputs(4745) <= not (a or b);
    layer3_outputs(4746) <= not (a or b);
    layer3_outputs(4747) <= a;
    layer3_outputs(4748) <= not b;
    layer3_outputs(4749) <= not b;
    layer3_outputs(4750) <= not (a and b);
    layer3_outputs(4751) <= a or b;
    layer3_outputs(4752) <= a and not b;
    layer3_outputs(4753) <= not a;
    layer3_outputs(4754) <= not (a and b);
    layer3_outputs(4755) <= a or b;
    layer3_outputs(4756) <= a or b;
    layer3_outputs(4757) <= a and not b;
    layer3_outputs(4758) <= a;
    layer3_outputs(4759) <= b;
    layer3_outputs(4760) <= a;
    layer3_outputs(4761) <= a and b;
    layer3_outputs(4762) <= b and not a;
    layer3_outputs(4763) <= a xor b;
    layer3_outputs(4764) <= a and b;
    layer3_outputs(4765) <= b;
    layer3_outputs(4766) <= not (a xor b);
    layer3_outputs(4767) <= a;
    layer3_outputs(4768) <= b and not a;
    layer3_outputs(4769) <= not a;
    layer3_outputs(4770) <= not a;
    layer3_outputs(4771) <= a and not b;
    layer3_outputs(4772) <= not (a or b);
    layer3_outputs(4773) <= not (a or b);
    layer3_outputs(4774) <= not (a and b);
    layer3_outputs(4775) <= not (a or b);
    layer3_outputs(4776) <= b;
    layer3_outputs(4777) <= not b or a;
    layer3_outputs(4778) <= a and not b;
    layer3_outputs(4779) <= not b or a;
    layer3_outputs(4780) <= not b or a;
    layer3_outputs(4781) <= not b;
    layer3_outputs(4782) <= not (a and b);
    layer3_outputs(4783) <= a or b;
    layer3_outputs(4784) <= not (a xor b);
    layer3_outputs(4785) <= a;
    layer3_outputs(4786) <= not (a or b);
    layer3_outputs(4787) <= not a or b;
    layer3_outputs(4788) <= a and not b;
    layer3_outputs(4789) <= a or b;
    layer3_outputs(4790) <= a;
    layer3_outputs(4791) <= not a or b;
    layer3_outputs(4792) <= b;
    layer3_outputs(4793) <= a and not b;
    layer3_outputs(4794) <= not (a and b);
    layer3_outputs(4795) <= a xor b;
    layer3_outputs(4796) <= a or b;
    layer3_outputs(4797) <= b;
    layer3_outputs(4798) <= a and not b;
    layer3_outputs(4799) <= not a or b;
    layer3_outputs(4800) <= a and not b;
    layer3_outputs(4801) <= a;
    layer3_outputs(4802) <= not b;
    layer3_outputs(4803) <= b;
    layer3_outputs(4804) <= a or b;
    layer3_outputs(4805) <= not b;
    layer3_outputs(4806) <= a and b;
    layer3_outputs(4807) <= not a;
    layer3_outputs(4808) <= a and not b;
    layer3_outputs(4809) <= not b;
    layer3_outputs(4810) <= not a;
    layer3_outputs(4811) <= '0';
    layer3_outputs(4812) <= '1';
    layer3_outputs(4813) <= not b;
    layer3_outputs(4814) <= not (a and b);
    layer3_outputs(4815) <= b;
    layer3_outputs(4816) <= not (a xor b);
    layer3_outputs(4817) <= not a;
    layer3_outputs(4818) <= not a or b;
    layer3_outputs(4819) <= b and not a;
    layer3_outputs(4820) <= not a;
    layer3_outputs(4821) <= not b or a;
    layer3_outputs(4822) <= not a;
    layer3_outputs(4823) <= a xor b;
    layer3_outputs(4824) <= a or b;
    layer3_outputs(4825) <= '1';
    layer3_outputs(4826) <= a and b;
    layer3_outputs(4827) <= a;
    layer3_outputs(4828) <= not (a xor b);
    layer3_outputs(4829) <= not a;
    layer3_outputs(4830) <= a and b;
    layer3_outputs(4831) <= not (a xor b);
    layer3_outputs(4832) <= not b;
    layer3_outputs(4833) <= b and not a;
    layer3_outputs(4834) <= b;
    layer3_outputs(4835) <= a or b;
    layer3_outputs(4836) <= '0';
    layer3_outputs(4837) <= not a;
    layer3_outputs(4838) <= a;
    layer3_outputs(4839) <= b and not a;
    layer3_outputs(4840) <= not a;
    layer3_outputs(4841) <= not b;
    layer3_outputs(4842) <= a xor b;
    layer3_outputs(4843) <= not (a or b);
    layer3_outputs(4844) <= a;
    layer3_outputs(4845) <= not (a or b);
    layer3_outputs(4846) <= a and not b;
    layer3_outputs(4847) <= not (a xor b);
    layer3_outputs(4848) <= a;
    layer3_outputs(4849) <= a;
    layer3_outputs(4850) <= a;
    layer3_outputs(4851) <= not (a xor b);
    layer3_outputs(4852) <= not b;
    layer3_outputs(4853) <= not (a and b);
    layer3_outputs(4854) <= not a;
    layer3_outputs(4855) <= not a or b;
    layer3_outputs(4856) <= not b or a;
    layer3_outputs(4857) <= '0';
    layer3_outputs(4858) <= b;
    layer3_outputs(4859) <= b;
    layer3_outputs(4860) <= a and b;
    layer3_outputs(4861) <= a or b;
    layer3_outputs(4862) <= not (a and b);
    layer3_outputs(4863) <= a or b;
    layer3_outputs(4864) <= not a or b;
    layer3_outputs(4865) <= a or b;
    layer3_outputs(4866) <= not a;
    layer3_outputs(4867) <= not b;
    layer3_outputs(4868) <= b;
    layer3_outputs(4869) <= not (a or b);
    layer3_outputs(4870) <= a xor b;
    layer3_outputs(4871) <= not a or b;
    layer3_outputs(4872) <= not a or b;
    layer3_outputs(4873) <= not b;
    layer3_outputs(4874) <= not b;
    layer3_outputs(4875) <= not (a or b);
    layer3_outputs(4876) <= not (a and b);
    layer3_outputs(4877) <= not b;
    layer3_outputs(4878) <= b and not a;
    layer3_outputs(4879) <= a;
    layer3_outputs(4880) <= b;
    layer3_outputs(4881) <= b;
    layer3_outputs(4882) <= a;
    layer3_outputs(4883) <= not a;
    layer3_outputs(4884) <= '0';
    layer3_outputs(4885) <= b;
    layer3_outputs(4886) <= b;
    layer3_outputs(4887) <= '0';
    layer3_outputs(4888) <= not b;
    layer3_outputs(4889) <= not b or a;
    layer3_outputs(4890) <= not b;
    layer3_outputs(4891) <= not a;
    layer3_outputs(4892) <= '0';
    layer3_outputs(4893) <= b;
    layer3_outputs(4894) <= not a or b;
    layer3_outputs(4895) <= not a or b;
    layer3_outputs(4896) <= b and not a;
    layer3_outputs(4897) <= '1';
    layer3_outputs(4898) <= not (a and b);
    layer3_outputs(4899) <= '1';
    layer3_outputs(4900) <= not (a xor b);
    layer3_outputs(4901) <= a;
    layer3_outputs(4902) <= not a;
    layer3_outputs(4903) <= not b;
    layer3_outputs(4904) <= a;
    layer3_outputs(4905) <= not (a and b);
    layer3_outputs(4906) <= a;
    layer3_outputs(4907) <= b and not a;
    layer3_outputs(4908) <= a and b;
    layer3_outputs(4909) <= not b or a;
    layer3_outputs(4910) <= a xor b;
    layer3_outputs(4911) <= b;
    layer3_outputs(4912) <= a or b;
    layer3_outputs(4913) <= a or b;
    layer3_outputs(4914) <= a and b;
    layer3_outputs(4915) <= not (a xor b);
    layer3_outputs(4916) <= not a or b;
    layer3_outputs(4917) <= a;
    layer3_outputs(4918) <= b;
    layer3_outputs(4919) <= not (a or b);
    layer3_outputs(4920) <= a and not b;
    layer3_outputs(4921) <= a and b;
    layer3_outputs(4922) <= not b or a;
    layer3_outputs(4923) <= b;
    layer3_outputs(4924) <= not a;
    layer3_outputs(4925) <= not b or a;
    layer3_outputs(4926) <= not b or a;
    layer3_outputs(4927) <= not a or b;
    layer3_outputs(4928) <= a and not b;
    layer3_outputs(4929) <= not b;
    layer3_outputs(4930) <= not b;
    layer3_outputs(4931) <= not (a and b);
    layer3_outputs(4932) <= b;
    layer3_outputs(4933) <= not (a xor b);
    layer3_outputs(4934) <= not (a and b);
    layer3_outputs(4935) <= not b or a;
    layer3_outputs(4936) <= not a or b;
    layer3_outputs(4937) <= not (a xor b);
    layer3_outputs(4938) <= b;
    layer3_outputs(4939) <= a and not b;
    layer3_outputs(4940) <= a or b;
    layer3_outputs(4941) <= a;
    layer3_outputs(4942) <= a and b;
    layer3_outputs(4943) <= not b;
    layer3_outputs(4944) <= not b;
    layer3_outputs(4945) <= not b;
    layer3_outputs(4946) <= not b;
    layer3_outputs(4947) <= a;
    layer3_outputs(4948) <= a and not b;
    layer3_outputs(4949) <= a and not b;
    layer3_outputs(4950) <= not (a or b);
    layer3_outputs(4951) <= not b or a;
    layer3_outputs(4952) <= a;
    layer3_outputs(4953) <= not b or a;
    layer3_outputs(4954) <= not a or b;
    layer3_outputs(4955) <= a and b;
    layer3_outputs(4956) <= a;
    layer3_outputs(4957) <= b;
    layer3_outputs(4958) <= not (a and b);
    layer3_outputs(4959) <= not a;
    layer3_outputs(4960) <= not (a and b);
    layer3_outputs(4961) <= b;
    layer3_outputs(4962) <= a;
    layer3_outputs(4963) <= b;
    layer3_outputs(4964) <= not a;
    layer3_outputs(4965) <= not b;
    layer3_outputs(4966) <= not b;
    layer3_outputs(4967) <= not a;
    layer3_outputs(4968) <= b;
    layer3_outputs(4969) <= not (a and b);
    layer3_outputs(4970) <= not a;
    layer3_outputs(4971) <= not (a xor b);
    layer3_outputs(4972) <= a xor b;
    layer3_outputs(4973) <= a and b;
    layer3_outputs(4974) <= not a;
    layer3_outputs(4975) <= b;
    layer3_outputs(4976) <= not a or b;
    layer3_outputs(4977) <= b;
    layer3_outputs(4978) <= not a;
    layer3_outputs(4979) <= a or b;
    layer3_outputs(4980) <= not a or b;
    layer3_outputs(4981) <= not (a xor b);
    layer3_outputs(4982) <= a and b;
    layer3_outputs(4983) <= not b;
    layer3_outputs(4984) <= a and b;
    layer3_outputs(4985) <= not (a and b);
    layer3_outputs(4986) <= a xor b;
    layer3_outputs(4987) <= b;
    layer3_outputs(4988) <= '1';
    layer3_outputs(4989) <= '1';
    layer3_outputs(4990) <= '0';
    layer3_outputs(4991) <= not b or a;
    layer3_outputs(4992) <= not a or b;
    layer3_outputs(4993) <= a and b;
    layer3_outputs(4994) <= not b or a;
    layer3_outputs(4995) <= b;
    layer3_outputs(4996) <= not a;
    layer3_outputs(4997) <= a xor b;
    layer3_outputs(4998) <= not a;
    layer3_outputs(4999) <= a and b;
    layer3_outputs(5000) <= a and b;
    layer3_outputs(5001) <= b;
    layer3_outputs(5002) <= not (a or b);
    layer3_outputs(5003) <= a;
    layer3_outputs(5004) <= a;
    layer3_outputs(5005) <= a;
    layer3_outputs(5006) <= a and not b;
    layer3_outputs(5007) <= not b;
    layer3_outputs(5008) <= b;
    layer3_outputs(5009) <= b;
    layer3_outputs(5010) <= b and not a;
    layer3_outputs(5011) <= not a;
    layer3_outputs(5012) <= not a or b;
    layer3_outputs(5013) <= not (a or b);
    layer3_outputs(5014) <= not a;
    layer3_outputs(5015) <= not (a or b);
    layer3_outputs(5016) <= a or b;
    layer3_outputs(5017) <= a xor b;
    layer3_outputs(5018) <= not b;
    layer3_outputs(5019) <= not b;
    layer3_outputs(5020) <= b;
    layer3_outputs(5021) <= b;
    layer3_outputs(5022) <= b and not a;
    layer3_outputs(5023) <= not (a xor b);
    layer3_outputs(5024) <= not a;
    layer3_outputs(5025) <= not b;
    layer3_outputs(5026) <= a;
    layer3_outputs(5027) <= b;
    layer3_outputs(5028) <= not b or a;
    layer3_outputs(5029) <= not a;
    layer3_outputs(5030) <= not b or a;
    layer3_outputs(5031) <= a xor b;
    layer3_outputs(5032) <= b and not a;
    layer3_outputs(5033) <= a;
    layer3_outputs(5034) <= a xor b;
    layer3_outputs(5035) <= not (a xor b);
    layer3_outputs(5036) <= not b or a;
    layer3_outputs(5037) <= not (a xor b);
    layer3_outputs(5038) <= not (a or b);
    layer3_outputs(5039) <= not b;
    layer3_outputs(5040) <= a;
    layer3_outputs(5041) <= not b;
    layer3_outputs(5042) <= a or b;
    layer3_outputs(5043) <= a and b;
    layer3_outputs(5044) <= b;
    layer3_outputs(5045) <= not a or b;
    layer3_outputs(5046) <= a and not b;
    layer3_outputs(5047) <= not b or a;
    layer3_outputs(5048) <= not b or a;
    layer3_outputs(5049) <= not (a and b);
    layer3_outputs(5050) <= not b;
    layer3_outputs(5051) <= b;
    layer3_outputs(5052) <= not (a xor b);
    layer3_outputs(5053) <= not (a and b);
    layer3_outputs(5054) <= not a;
    layer3_outputs(5055) <= not b or a;
    layer3_outputs(5056) <= a and b;
    layer3_outputs(5057) <= a xor b;
    layer3_outputs(5058) <= not (a or b);
    layer3_outputs(5059) <= a;
    layer3_outputs(5060) <= a and b;
    layer3_outputs(5061) <= not (a or b);
    layer3_outputs(5062) <= not a;
    layer3_outputs(5063) <= b;
    layer3_outputs(5064) <= a and b;
    layer3_outputs(5065) <= a;
    layer3_outputs(5066) <= not (a or b);
    layer3_outputs(5067) <= not a;
    layer3_outputs(5068) <= '1';
    layer3_outputs(5069) <= not b;
    layer3_outputs(5070) <= b;
    layer3_outputs(5071) <= a and b;
    layer3_outputs(5072) <= b and not a;
    layer3_outputs(5073) <= b;
    layer3_outputs(5074) <= not (a xor b);
    layer3_outputs(5075) <= a xor b;
    layer3_outputs(5076) <= not (a xor b);
    layer3_outputs(5077) <= not a or b;
    layer3_outputs(5078) <= a;
    layer3_outputs(5079) <= b;
    layer3_outputs(5080) <= not a;
    layer3_outputs(5081) <= b;
    layer3_outputs(5082) <= not b or a;
    layer3_outputs(5083) <= a;
    layer3_outputs(5084) <= a;
    layer3_outputs(5085) <= not (a and b);
    layer3_outputs(5086) <= not a;
    layer3_outputs(5087) <= a or b;
    layer3_outputs(5088) <= a and b;
    layer3_outputs(5089) <= a or b;
    layer3_outputs(5090) <= not (a and b);
    layer3_outputs(5091) <= a;
    layer3_outputs(5092) <= not a;
    layer3_outputs(5093) <= not b;
    layer3_outputs(5094) <= a or b;
    layer3_outputs(5095) <= a xor b;
    layer3_outputs(5096) <= a or b;
    layer3_outputs(5097) <= not b or a;
    layer3_outputs(5098) <= not b or a;
    layer3_outputs(5099) <= a or b;
    layer3_outputs(5100) <= not (a and b);
    layer3_outputs(5101) <= not a;
    layer3_outputs(5102) <= not b;
    layer3_outputs(5103) <= not a;
    layer3_outputs(5104) <= a xor b;
    layer3_outputs(5105) <= a and not b;
    layer3_outputs(5106) <= not b;
    layer3_outputs(5107) <= a and not b;
    layer3_outputs(5108) <= not b or a;
    layer3_outputs(5109) <= not a;
    layer3_outputs(5110) <= b;
    layer3_outputs(5111) <= not a or b;
    layer3_outputs(5112) <= not a;
    layer3_outputs(5113) <= not b;
    layer3_outputs(5114) <= a;
    layer3_outputs(5115) <= a and b;
    layer3_outputs(5116) <= b;
    layer3_outputs(5117) <= not a;
    layer3_outputs(5118) <= not a;
    layer3_outputs(5119) <= b;
    layer4_outputs(0) <= a and not b;
    layer4_outputs(1) <= b;
    layer4_outputs(2) <= not (a or b);
    layer4_outputs(3) <= b;
    layer4_outputs(4) <= a or b;
    layer4_outputs(5) <= not (a or b);
    layer4_outputs(6) <= not (a xor b);
    layer4_outputs(7) <= not (a and b);
    layer4_outputs(8) <= b;
    layer4_outputs(9) <= a xor b;
    layer4_outputs(10) <= b;
    layer4_outputs(11) <= not (a and b);
    layer4_outputs(12) <= b and not a;
    layer4_outputs(13) <= a or b;
    layer4_outputs(14) <= b and not a;
    layer4_outputs(15) <= not b or a;
    layer4_outputs(16) <= not (a xor b);
    layer4_outputs(17) <= a and b;
    layer4_outputs(18) <= b;
    layer4_outputs(19) <= b and not a;
    layer4_outputs(20) <= a;
    layer4_outputs(21) <= not a or b;
    layer4_outputs(22) <= not b;
    layer4_outputs(23) <= not (a xor b);
    layer4_outputs(24) <= not b;
    layer4_outputs(25) <= not b;
    layer4_outputs(26) <= b and not a;
    layer4_outputs(27) <= a;
    layer4_outputs(28) <= not a;
    layer4_outputs(29) <= not (a or b);
    layer4_outputs(30) <= b and not a;
    layer4_outputs(31) <= a;
    layer4_outputs(32) <= not (a xor b);
    layer4_outputs(33) <= not b;
    layer4_outputs(34) <= a;
    layer4_outputs(35) <= a and b;
    layer4_outputs(36) <= not a;
    layer4_outputs(37) <= not b;
    layer4_outputs(38) <= a or b;
    layer4_outputs(39) <= not b;
    layer4_outputs(40) <= a;
    layer4_outputs(41) <= a;
    layer4_outputs(42) <= a xor b;
    layer4_outputs(43) <= a;
    layer4_outputs(44) <= not b;
    layer4_outputs(45) <= b;
    layer4_outputs(46) <= a or b;
    layer4_outputs(47) <= not a;
    layer4_outputs(48) <= not (a and b);
    layer4_outputs(49) <= b;
    layer4_outputs(50) <= b;
    layer4_outputs(51) <= not b;
    layer4_outputs(52) <= b and not a;
    layer4_outputs(53) <= not (a and b);
    layer4_outputs(54) <= not a;
    layer4_outputs(55) <= a and not b;
    layer4_outputs(56) <= not a;
    layer4_outputs(57) <= b;
    layer4_outputs(58) <= a;
    layer4_outputs(59) <= not a;
    layer4_outputs(60) <= b and not a;
    layer4_outputs(61) <= not a;
    layer4_outputs(62) <= not (a xor b);
    layer4_outputs(63) <= not a;
    layer4_outputs(64) <= a and b;
    layer4_outputs(65) <= b and not a;
    layer4_outputs(66) <= not a;
    layer4_outputs(67) <= a xor b;
    layer4_outputs(68) <= not (a xor b);
    layer4_outputs(69) <= a;
    layer4_outputs(70) <= a and b;
    layer4_outputs(71) <= '0';
    layer4_outputs(72) <= not a;
    layer4_outputs(73) <= b and not a;
    layer4_outputs(74) <= not b;
    layer4_outputs(75) <= not b or a;
    layer4_outputs(76) <= not a;
    layer4_outputs(77) <= not a;
    layer4_outputs(78) <= not (a and b);
    layer4_outputs(79) <= not a or b;
    layer4_outputs(80) <= not (a xor b);
    layer4_outputs(81) <= a and not b;
    layer4_outputs(82) <= not b or a;
    layer4_outputs(83) <= b;
    layer4_outputs(84) <= not (a and b);
    layer4_outputs(85) <= not a;
    layer4_outputs(86) <= not (a and b);
    layer4_outputs(87) <= a and b;
    layer4_outputs(88) <= b;
    layer4_outputs(89) <= not b;
    layer4_outputs(90) <= a xor b;
    layer4_outputs(91) <= b;
    layer4_outputs(92) <= not b;
    layer4_outputs(93) <= a or b;
    layer4_outputs(94) <= a or b;
    layer4_outputs(95) <= a and b;
    layer4_outputs(96) <= not b;
    layer4_outputs(97) <= a and b;
    layer4_outputs(98) <= not a;
    layer4_outputs(99) <= not (a xor b);
    layer4_outputs(100) <= a or b;
    layer4_outputs(101) <= b;
    layer4_outputs(102) <= b;
    layer4_outputs(103) <= not a;
    layer4_outputs(104) <= not b;
    layer4_outputs(105) <= not (a xor b);
    layer4_outputs(106) <= b;
    layer4_outputs(107) <= not a or b;
    layer4_outputs(108) <= not (a and b);
    layer4_outputs(109) <= not (a or b);
    layer4_outputs(110) <= not a;
    layer4_outputs(111) <= not b or a;
    layer4_outputs(112) <= not (a and b);
    layer4_outputs(113) <= a;
    layer4_outputs(114) <= not (a xor b);
    layer4_outputs(115) <= not (a and b);
    layer4_outputs(116) <= b and not a;
    layer4_outputs(117) <= a;
    layer4_outputs(118) <= not b;
    layer4_outputs(119) <= not b;
    layer4_outputs(120) <= not (a or b);
    layer4_outputs(121) <= not (a xor b);
    layer4_outputs(122) <= not a or b;
    layer4_outputs(123) <= not b;
    layer4_outputs(124) <= not a;
    layer4_outputs(125) <= a;
    layer4_outputs(126) <= not (a or b);
    layer4_outputs(127) <= not (a xor b);
    layer4_outputs(128) <= not a;
    layer4_outputs(129) <= not a;
    layer4_outputs(130) <= not b or a;
    layer4_outputs(131) <= not b or a;
    layer4_outputs(132) <= a;
    layer4_outputs(133) <= a and b;
    layer4_outputs(134) <= not (a or b);
    layer4_outputs(135) <= not (a or b);
    layer4_outputs(136) <= not a;
    layer4_outputs(137) <= a;
    layer4_outputs(138) <= b;
    layer4_outputs(139) <= b;
    layer4_outputs(140) <= not b;
    layer4_outputs(141) <= a;
    layer4_outputs(142) <= b and not a;
    layer4_outputs(143) <= not b;
    layer4_outputs(144) <= not b;
    layer4_outputs(145) <= not b;
    layer4_outputs(146) <= not b;
    layer4_outputs(147) <= not a;
    layer4_outputs(148) <= b and not a;
    layer4_outputs(149) <= a;
    layer4_outputs(150) <= not (a or b);
    layer4_outputs(151) <= a;
    layer4_outputs(152) <= a and b;
    layer4_outputs(153) <= not a;
    layer4_outputs(154) <= not a;
    layer4_outputs(155) <= a or b;
    layer4_outputs(156) <= not b or a;
    layer4_outputs(157) <= not (a or b);
    layer4_outputs(158) <= not a;
    layer4_outputs(159) <= a xor b;
    layer4_outputs(160) <= not b;
    layer4_outputs(161) <= not (a or b);
    layer4_outputs(162) <= not (a and b);
    layer4_outputs(163) <= a and not b;
    layer4_outputs(164) <= not b;
    layer4_outputs(165) <= not (a and b);
    layer4_outputs(166) <= not b;
    layer4_outputs(167) <= a and not b;
    layer4_outputs(168) <= not (a xor b);
    layer4_outputs(169) <= a;
    layer4_outputs(170) <= not b;
    layer4_outputs(171) <= b;
    layer4_outputs(172) <= a and not b;
    layer4_outputs(173) <= not b;
    layer4_outputs(174) <= not b;
    layer4_outputs(175) <= not a;
    layer4_outputs(176) <= not (a and b);
    layer4_outputs(177) <= not (a xor b);
    layer4_outputs(178) <= not b;
    layer4_outputs(179) <= not b;
    layer4_outputs(180) <= not a;
    layer4_outputs(181) <= a and not b;
    layer4_outputs(182) <= a;
    layer4_outputs(183) <= b and not a;
    layer4_outputs(184) <= not b;
    layer4_outputs(185) <= not a;
    layer4_outputs(186) <= not b;
    layer4_outputs(187) <= not (a or b);
    layer4_outputs(188) <= not (a and b);
    layer4_outputs(189) <= a;
    layer4_outputs(190) <= a;
    layer4_outputs(191) <= a;
    layer4_outputs(192) <= not (a or b);
    layer4_outputs(193) <= not (a or b);
    layer4_outputs(194) <= a xor b;
    layer4_outputs(195) <= a and not b;
    layer4_outputs(196) <= a or b;
    layer4_outputs(197) <= a or b;
    layer4_outputs(198) <= a;
    layer4_outputs(199) <= not b;
    layer4_outputs(200) <= not a;
    layer4_outputs(201) <= not b;
    layer4_outputs(202) <= not b or a;
    layer4_outputs(203) <= a and b;
    layer4_outputs(204) <= b;
    layer4_outputs(205) <= b and not a;
    layer4_outputs(206) <= not a or b;
    layer4_outputs(207) <= b;
    layer4_outputs(208) <= a xor b;
    layer4_outputs(209) <= a xor b;
    layer4_outputs(210) <= not a or b;
    layer4_outputs(211) <= a;
    layer4_outputs(212) <= not a;
    layer4_outputs(213) <= not b;
    layer4_outputs(214) <= b and not a;
    layer4_outputs(215) <= a xor b;
    layer4_outputs(216) <= a and b;
    layer4_outputs(217) <= not (a xor b);
    layer4_outputs(218) <= not b;
    layer4_outputs(219) <= not b;
    layer4_outputs(220) <= b;
    layer4_outputs(221) <= b;
    layer4_outputs(222) <= b;
    layer4_outputs(223) <= b;
    layer4_outputs(224) <= not (a and b);
    layer4_outputs(225) <= not (a and b);
    layer4_outputs(226) <= b and not a;
    layer4_outputs(227) <= not a;
    layer4_outputs(228) <= not a or b;
    layer4_outputs(229) <= a;
    layer4_outputs(230) <= a xor b;
    layer4_outputs(231) <= a or b;
    layer4_outputs(232) <= not b;
    layer4_outputs(233) <= not a;
    layer4_outputs(234) <= not b;
    layer4_outputs(235) <= not (a xor b);
    layer4_outputs(236) <= not b;
    layer4_outputs(237) <= a;
    layer4_outputs(238) <= b;
    layer4_outputs(239) <= not b;
    layer4_outputs(240) <= a;
    layer4_outputs(241) <= not (a xor b);
    layer4_outputs(242) <= not (a and b);
    layer4_outputs(243) <= not b or a;
    layer4_outputs(244) <= a xor b;
    layer4_outputs(245) <= not b or a;
    layer4_outputs(246) <= a;
    layer4_outputs(247) <= a;
    layer4_outputs(248) <= not a or b;
    layer4_outputs(249) <= not b or a;
    layer4_outputs(250) <= not a;
    layer4_outputs(251) <= a;
    layer4_outputs(252) <= not (a xor b);
    layer4_outputs(253) <= not a or b;
    layer4_outputs(254) <= '0';
    layer4_outputs(255) <= not b or a;
    layer4_outputs(256) <= b;
    layer4_outputs(257) <= not b;
    layer4_outputs(258) <= a;
    layer4_outputs(259) <= '1';
    layer4_outputs(260) <= a and b;
    layer4_outputs(261) <= a xor b;
    layer4_outputs(262) <= not (a or b);
    layer4_outputs(263) <= not a;
    layer4_outputs(264) <= not b or a;
    layer4_outputs(265) <= b and not a;
    layer4_outputs(266) <= not a;
    layer4_outputs(267) <= not a or b;
    layer4_outputs(268) <= not b or a;
    layer4_outputs(269) <= a and not b;
    layer4_outputs(270) <= not a;
    layer4_outputs(271) <= not b or a;
    layer4_outputs(272) <= a xor b;
    layer4_outputs(273) <= a or b;
    layer4_outputs(274) <= a or b;
    layer4_outputs(275) <= b;
    layer4_outputs(276) <= not (a and b);
    layer4_outputs(277) <= a and b;
    layer4_outputs(278) <= not a;
    layer4_outputs(279) <= not (a and b);
    layer4_outputs(280) <= a or b;
    layer4_outputs(281) <= b;
    layer4_outputs(282) <= a xor b;
    layer4_outputs(283) <= b;
    layer4_outputs(284) <= a;
    layer4_outputs(285) <= a;
    layer4_outputs(286) <= not (a xor b);
    layer4_outputs(287) <= not b;
    layer4_outputs(288) <= a or b;
    layer4_outputs(289) <= '1';
    layer4_outputs(290) <= a and not b;
    layer4_outputs(291) <= not b;
    layer4_outputs(292) <= not b or a;
    layer4_outputs(293) <= b;
    layer4_outputs(294) <= not a;
    layer4_outputs(295) <= not b;
    layer4_outputs(296) <= not (a or b);
    layer4_outputs(297) <= a;
    layer4_outputs(298) <= a or b;
    layer4_outputs(299) <= not (a or b);
    layer4_outputs(300) <= a and b;
    layer4_outputs(301) <= not (a and b);
    layer4_outputs(302) <= a;
    layer4_outputs(303) <= a and not b;
    layer4_outputs(304) <= b;
    layer4_outputs(305) <= a or b;
    layer4_outputs(306) <= not a;
    layer4_outputs(307) <= not b;
    layer4_outputs(308) <= b;
    layer4_outputs(309) <= a;
    layer4_outputs(310) <= not (a xor b);
    layer4_outputs(311) <= not (a xor b);
    layer4_outputs(312) <= not a or b;
    layer4_outputs(313) <= not a;
    layer4_outputs(314) <= a and not b;
    layer4_outputs(315) <= b;
    layer4_outputs(316) <= b and not a;
    layer4_outputs(317) <= b and not a;
    layer4_outputs(318) <= a;
    layer4_outputs(319) <= a;
    layer4_outputs(320) <= a and b;
    layer4_outputs(321) <= not a or b;
    layer4_outputs(322) <= a or b;
    layer4_outputs(323) <= not b;
    layer4_outputs(324) <= a;
    layer4_outputs(325) <= b;
    layer4_outputs(326) <= b;
    layer4_outputs(327) <= a xor b;
    layer4_outputs(328) <= not b;
    layer4_outputs(329) <= b;
    layer4_outputs(330) <= a and not b;
    layer4_outputs(331) <= b;
    layer4_outputs(332) <= b and not a;
    layer4_outputs(333) <= not b;
    layer4_outputs(334) <= not a;
    layer4_outputs(335) <= a xor b;
    layer4_outputs(336) <= not (a xor b);
    layer4_outputs(337) <= not (a or b);
    layer4_outputs(338) <= a;
    layer4_outputs(339) <= b;
    layer4_outputs(340) <= b;
    layer4_outputs(341) <= not b;
    layer4_outputs(342) <= a xor b;
    layer4_outputs(343) <= not a or b;
    layer4_outputs(344) <= a and b;
    layer4_outputs(345) <= '0';
    layer4_outputs(346) <= a and b;
    layer4_outputs(347) <= not (a xor b);
    layer4_outputs(348) <= not (a and b);
    layer4_outputs(349) <= not b;
    layer4_outputs(350) <= b;
    layer4_outputs(351) <= not (a or b);
    layer4_outputs(352) <= a and b;
    layer4_outputs(353) <= b;
    layer4_outputs(354) <= a;
    layer4_outputs(355) <= not (a xor b);
    layer4_outputs(356) <= a and b;
    layer4_outputs(357) <= not a;
    layer4_outputs(358) <= not (a and b);
    layer4_outputs(359) <= a and not b;
    layer4_outputs(360) <= a and not b;
    layer4_outputs(361) <= not a or b;
    layer4_outputs(362) <= a;
    layer4_outputs(363) <= not b;
    layer4_outputs(364) <= a and b;
    layer4_outputs(365) <= b;
    layer4_outputs(366) <= not a or b;
    layer4_outputs(367) <= not a;
    layer4_outputs(368) <= b;
    layer4_outputs(369) <= a;
    layer4_outputs(370) <= a or b;
    layer4_outputs(371) <= not b or a;
    layer4_outputs(372) <= b;
    layer4_outputs(373) <= not (a or b);
    layer4_outputs(374) <= a;
    layer4_outputs(375) <= a;
    layer4_outputs(376) <= a xor b;
    layer4_outputs(377) <= not a;
    layer4_outputs(378) <= not b or a;
    layer4_outputs(379) <= not (a and b);
    layer4_outputs(380) <= not a or b;
    layer4_outputs(381) <= a xor b;
    layer4_outputs(382) <= b and not a;
    layer4_outputs(383) <= not b;
    layer4_outputs(384) <= a and b;
    layer4_outputs(385) <= not b or a;
    layer4_outputs(386) <= b and not a;
    layer4_outputs(387) <= not (a and b);
    layer4_outputs(388) <= b;
    layer4_outputs(389) <= a;
    layer4_outputs(390) <= a and b;
    layer4_outputs(391) <= a or b;
    layer4_outputs(392) <= not b;
    layer4_outputs(393) <= not b;
    layer4_outputs(394) <= not a;
    layer4_outputs(395) <= b;
    layer4_outputs(396) <= b;
    layer4_outputs(397) <= a and b;
    layer4_outputs(398) <= b;
    layer4_outputs(399) <= a;
    layer4_outputs(400) <= a and not b;
    layer4_outputs(401) <= not a;
    layer4_outputs(402) <= not (a xor b);
    layer4_outputs(403) <= a xor b;
    layer4_outputs(404) <= not a or b;
    layer4_outputs(405) <= not (a xor b);
    layer4_outputs(406) <= a or b;
    layer4_outputs(407) <= b and not a;
    layer4_outputs(408) <= a and not b;
    layer4_outputs(409) <= a;
    layer4_outputs(410) <= not a;
    layer4_outputs(411) <= a and not b;
    layer4_outputs(412) <= a and not b;
    layer4_outputs(413) <= not (a and b);
    layer4_outputs(414) <= b;
    layer4_outputs(415) <= b;
    layer4_outputs(416) <= not (a xor b);
    layer4_outputs(417) <= not (a or b);
    layer4_outputs(418) <= not (a and b);
    layer4_outputs(419) <= not (a xor b);
    layer4_outputs(420) <= a and b;
    layer4_outputs(421) <= not (a xor b);
    layer4_outputs(422) <= a;
    layer4_outputs(423) <= a and not b;
    layer4_outputs(424) <= not a;
    layer4_outputs(425) <= not b;
    layer4_outputs(426) <= a and b;
    layer4_outputs(427) <= not (a or b);
    layer4_outputs(428) <= not a;
    layer4_outputs(429) <= not (a and b);
    layer4_outputs(430) <= b and not a;
    layer4_outputs(431) <= a;
    layer4_outputs(432) <= a;
    layer4_outputs(433) <= b;
    layer4_outputs(434) <= not (a or b);
    layer4_outputs(435) <= a xor b;
    layer4_outputs(436) <= a;
    layer4_outputs(437) <= not b or a;
    layer4_outputs(438) <= a and not b;
    layer4_outputs(439) <= a or b;
    layer4_outputs(440) <= not a;
    layer4_outputs(441) <= not (a xor b);
    layer4_outputs(442) <= not (a and b);
    layer4_outputs(443) <= not b or a;
    layer4_outputs(444) <= b;
    layer4_outputs(445) <= a;
    layer4_outputs(446) <= a and b;
    layer4_outputs(447) <= a and not b;
    layer4_outputs(448) <= not (a or b);
    layer4_outputs(449) <= not a;
    layer4_outputs(450) <= not a;
    layer4_outputs(451) <= not (a xor b);
    layer4_outputs(452) <= a xor b;
    layer4_outputs(453) <= a xor b;
    layer4_outputs(454) <= a;
    layer4_outputs(455) <= b;
    layer4_outputs(456) <= not (a and b);
    layer4_outputs(457) <= b and not a;
    layer4_outputs(458) <= a and not b;
    layer4_outputs(459) <= a xor b;
    layer4_outputs(460) <= not b;
    layer4_outputs(461) <= b;
    layer4_outputs(462) <= a xor b;
    layer4_outputs(463) <= a and not b;
    layer4_outputs(464) <= '0';
    layer4_outputs(465) <= a and not b;
    layer4_outputs(466) <= not (a or b);
    layer4_outputs(467) <= not b;
    layer4_outputs(468) <= a xor b;
    layer4_outputs(469) <= a xor b;
    layer4_outputs(470) <= not b;
    layer4_outputs(471) <= a;
    layer4_outputs(472) <= a;
    layer4_outputs(473) <= not (a xor b);
    layer4_outputs(474) <= a and b;
    layer4_outputs(475) <= not b;
    layer4_outputs(476) <= not (a xor b);
    layer4_outputs(477) <= not a;
    layer4_outputs(478) <= b and not a;
    layer4_outputs(479) <= a;
    layer4_outputs(480) <= not b or a;
    layer4_outputs(481) <= not b;
    layer4_outputs(482) <= a or b;
    layer4_outputs(483) <= b and not a;
    layer4_outputs(484) <= not (a xor b);
    layer4_outputs(485) <= not a;
    layer4_outputs(486) <= a or b;
    layer4_outputs(487) <= a;
    layer4_outputs(488) <= not a;
    layer4_outputs(489) <= not a;
    layer4_outputs(490) <= not a;
    layer4_outputs(491) <= not (a or b);
    layer4_outputs(492) <= a;
    layer4_outputs(493) <= not (a and b);
    layer4_outputs(494) <= a and not b;
    layer4_outputs(495) <= b;
    layer4_outputs(496) <= b;
    layer4_outputs(497) <= not (a or b);
    layer4_outputs(498) <= not b or a;
    layer4_outputs(499) <= not (a xor b);
    layer4_outputs(500) <= not b;
    layer4_outputs(501) <= a and not b;
    layer4_outputs(502) <= a;
    layer4_outputs(503) <= not a or b;
    layer4_outputs(504) <= not a;
    layer4_outputs(505) <= not a;
    layer4_outputs(506) <= not (a and b);
    layer4_outputs(507) <= b;
    layer4_outputs(508) <= a xor b;
    layer4_outputs(509) <= b;
    layer4_outputs(510) <= a or b;
    layer4_outputs(511) <= a;
    layer4_outputs(512) <= b;
    layer4_outputs(513) <= not b;
    layer4_outputs(514) <= a;
    layer4_outputs(515) <= not (a xor b);
    layer4_outputs(516) <= a and not b;
    layer4_outputs(517) <= not (a xor b);
    layer4_outputs(518) <= b and not a;
    layer4_outputs(519) <= b;
    layer4_outputs(520) <= not b;
    layer4_outputs(521) <= not a;
    layer4_outputs(522) <= not b or a;
    layer4_outputs(523) <= a and b;
    layer4_outputs(524) <= b and not a;
    layer4_outputs(525) <= a and b;
    layer4_outputs(526) <= not (a and b);
    layer4_outputs(527) <= not b;
    layer4_outputs(528) <= a xor b;
    layer4_outputs(529) <= a or b;
    layer4_outputs(530) <= b;
    layer4_outputs(531) <= a or b;
    layer4_outputs(532) <= not b or a;
    layer4_outputs(533) <= not (a or b);
    layer4_outputs(534) <= not (a xor b);
    layer4_outputs(535) <= a;
    layer4_outputs(536) <= not (a or b);
    layer4_outputs(537) <= b and not a;
    layer4_outputs(538) <= not (a or b);
    layer4_outputs(539) <= not b or a;
    layer4_outputs(540) <= not b;
    layer4_outputs(541) <= not (a and b);
    layer4_outputs(542) <= not a;
    layer4_outputs(543) <= a xor b;
    layer4_outputs(544) <= a or b;
    layer4_outputs(545) <= a;
    layer4_outputs(546) <= a xor b;
    layer4_outputs(547) <= not a;
    layer4_outputs(548) <= not b;
    layer4_outputs(549) <= not a or b;
    layer4_outputs(550) <= not a;
    layer4_outputs(551) <= a;
    layer4_outputs(552) <= not (a xor b);
    layer4_outputs(553) <= b and not a;
    layer4_outputs(554) <= a xor b;
    layer4_outputs(555) <= not b or a;
    layer4_outputs(556) <= a;
    layer4_outputs(557) <= a and b;
    layer4_outputs(558) <= not (a and b);
    layer4_outputs(559) <= not (a and b);
    layer4_outputs(560) <= not a or b;
    layer4_outputs(561) <= a and b;
    layer4_outputs(562) <= not (a or b);
    layer4_outputs(563) <= not a;
    layer4_outputs(564) <= a and b;
    layer4_outputs(565) <= a and not b;
    layer4_outputs(566) <= not (a xor b);
    layer4_outputs(567) <= not (a and b);
    layer4_outputs(568) <= not b;
    layer4_outputs(569) <= not a;
    layer4_outputs(570) <= not a or b;
    layer4_outputs(571) <= not a or b;
    layer4_outputs(572) <= not (a or b);
    layer4_outputs(573) <= b;
    layer4_outputs(574) <= b;
    layer4_outputs(575) <= a and not b;
    layer4_outputs(576) <= not a or b;
    layer4_outputs(577) <= '0';
    layer4_outputs(578) <= not b;
    layer4_outputs(579) <= a or b;
    layer4_outputs(580) <= a and not b;
    layer4_outputs(581) <= a or b;
    layer4_outputs(582) <= not b or a;
    layer4_outputs(583) <= b;
    layer4_outputs(584) <= not a;
    layer4_outputs(585) <= not (a or b);
    layer4_outputs(586) <= not (a and b);
    layer4_outputs(587) <= not a;
    layer4_outputs(588) <= b;
    layer4_outputs(589) <= not a or b;
    layer4_outputs(590) <= not a;
    layer4_outputs(591) <= not a;
    layer4_outputs(592) <= not b;
    layer4_outputs(593) <= not b;
    layer4_outputs(594) <= b and not a;
    layer4_outputs(595) <= a and not b;
    layer4_outputs(596) <= '0';
    layer4_outputs(597) <= not (a xor b);
    layer4_outputs(598) <= not a;
    layer4_outputs(599) <= not b;
    layer4_outputs(600) <= a and b;
    layer4_outputs(601) <= b and not a;
    layer4_outputs(602) <= not b or a;
    layer4_outputs(603) <= not b or a;
    layer4_outputs(604) <= a or b;
    layer4_outputs(605) <= not b or a;
    layer4_outputs(606) <= b;
    layer4_outputs(607) <= not (a or b);
    layer4_outputs(608) <= a and not b;
    layer4_outputs(609) <= b;
    layer4_outputs(610) <= not (a and b);
    layer4_outputs(611) <= b;
    layer4_outputs(612) <= not b or a;
    layer4_outputs(613) <= not (a xor b);
    layer4_outputs(614) <= not (a or b);
    layer4_outputs(615) <= a or b;
    layer4_outputs(616) <= not a or b;
    layer4_outputs(617) <= not b or a;
    layer4_outputs(618) <= not b;
    layer4_outputs(619) <= a;
    layer4_outputs(620) <= b;
    layer4_outputs(621) <= not b;
    layer4_outputs(622) <= not b;
    layer4_outputs(623) <= not (a and b);
    layer4_outputs(624) <= not b;
    layer4_outputs(625) <= not b;
    layer4_outputs(626) <= not (a or b);
    layer4_outputs(627) <= a;
    layer4_outputs(628) <= a xor b;
    layer4_outputs(629) <= not a;
    layer4_outputs(630) <= b;
    layer4_outputs(631) <= b;
    layer4_outputs(632) <= a and not b;
    layer4_outputs(633) <= a xor b;
    layer4_outputs(634) <= not a;
    layer4_outputs(635) <= a;
    layer4_outputs(636) <= a and b;
    layer4_outputs(637) <= not (a xor b);
    layer4_outputs(638) <= a xor b;
    layer4_outputs(639) <= not a or b;
    layer4_outputs(640) <= not b;
    layer4_outputs(641) <= not (a and b);
    layer4_outputs(642) <= a and not b;
    layer4_outputs(643) <= not a;
    layer4_outputs(644) <= a and not b;
    layer4_outputs(645) <= a and b;
    layer4_outputs(646) <= a and b;
    layer4_outputs(647) <= '1';
    layer4_outputs(648) <= a and b;
    layer4_outputs(649) <= not a;
    layer4_outputs(650) <= not a or b;
    layer4_outputs(651) <= not (a and b);
    layer4_outputs(652) <= not b or a;
    layer4_outputs(653) <= b and not a;
    layer4_outputs(654) <= not b;
    layer4_outputs(655) <= a and not b;
    layer4_outputs(656) <= b;
    layer4_outputs(657) <= not a;
    layer4_outputs(658) <= a xor b;
    layer4_outputs(659) <= b;
    layer4_outputs(660) <= not (a and b);
    layer4_outputs(661) <= not (a or b);
    layer4_outputs(662) <= b and not a;
    layer4_outputs(663) <= not b;
    layer4_outputs(664) <= not a or b;
    layer4_outputs(665) <= not a or b;
    layer4_outputs(666) <= not a;
    layer4_outputs(667) <= a and not b;
    layer4_outputs(668) <= b;
    layer4_outputs(669) <= not (a xor b);
    layer4_outputs(670) <= a;
    layer4_outputs(671) <= a and not b;
    layer4_outputs(672) <= a and b;
    layer4_outputs(673) <= b;
    layer4_outputs(674) <= a and not b;
    layer4_outputs(675) <= a xor b;
    layer4_outputs(676) <= not (a and b);
    layer4_outputs(677) <= '1';
    layer4_outputs(678) <= a;
    layer4_outputs(679) <= not (a or b);
    layer4_outputs(680) <= b;
    layer4_outputs(681) <= a;
    layer4_outputs(682) <= not b;
    layer4_outputs(683) <= not a or b;
    layer4_outputs(684) <= b;
    layer4_outputs(685) <= a and b;
    layer4_outputs(686) <= not a;
    layer4_outputs(687) <= a and not b;
    layer4_outputs(688) <= not (a or b);
    layer4_outputs(689) <= not (a xor b);
    layer4_outputs(690) <= a and not b;
    layer4_outputs(691) <= b;
    layer4_outputs(692) <= b;
    layer4_outputs(693) <= b and not a;
    layer4_outputs(694) <= not b;
    layer4_outputs(695) <= not b;
    layer4_outputs(696) <= not (a and b);
    layer4_outputs(697) <= not (a xor b);
    layer4_outputs(698) <= not (a and b);
    layer4_outputs(699) <= not b;
    layer4_outputs(700) <= a or b;
    layer4_outputs(701) <= b;
    layer4_outputs(702) <= '1';
    layer4_outputs(703) <= not a;
    layer4_outputs(704) <= a;
    layer4_outputs(705) <= not a or b;
    layer4_outputs(706) <= not b or a;
    layer4_outputs(707) <= b and not a;
    layer4_outputs(708) <= not (a or b);
    layer4_outputs(709) <= a or b;
    layer4_outputs(710) <= not a or b;
    layer4_outputs(711) <= a;
    layer4_outputs(712) <= not (a xor b);
    layer4_outputs(713) <= not (a and b);
    layer4_outputs(714) <= a or b;
    layer4_outputs(715) <= not a or b;
    layer4_outputs(716) <= a;
    layer4_outputs(717) <= a;
    layer4_outputs(718) <= a xor b;
    layer4_outputs(719) <= a and not b;
    layer4_outputs(720) <= not (a and b);
    layer4_outputs(721) <= b;
    layer4_outputs(722) <= not b;
    layer4_outputs(723) <= not (a xor b);
    layer4_outputs(724) <= b;
    layer4_outputs(725) <= a and not b;
    layer4_outputs(726) <= a;
    layer4_outputs(727) <= not a;
    layer4_outputs(728) <= not (a and b);
    layer4_outputs(729) <= a;
    layer4_outputs(730) <= not a;
    layer4_outputs(731) <= b and not a;
    layer4_outputs(732) <= not a or b;
    layer4_outputs(733) <= b;
    layer4_outputs(734) <= b;
    layer4_outputs(735) <= not a;
    layer4_outputs(736) <= not b;
    layer4_outputs(737) <= not (a and b);
    layer4_outputs(738) <= not b;
    layer4_outputs(739) <= not (a or b);
    layer4_outputs(740) <= not (a or b);
    layer4_outputs(741) <= b;
    layer4_outputs(742) <= b;
    layer4_outputs(743) <= a;
    layer4_outputs(744) <= not a;
    layer4_outputs(745) <= not a or b;
    layer4_outputs(746) <= not b;
    layer4_outputs(747) <= a;
    layer4_outputs(748) <= not b or a;
    layer4_outputs(749) <= a or b;
    layer4_outputs(750) <= b;
    layer4_outputs(751) <= not a;
    layer4_outputs(752) <= not (a xor b);
    layer4_outputs(753) <= a;
    layer4_outputs(754) <= a and b;
    layer4_outputs(755) <= a xor b;
    layer4_outputs(756) <= a or b;
    layer4_outputs(757) <= not (a and b);
    layer4_outputs(758) <= b and not a;
    layer4_outputs(759) <= b;
    layer4_outputs(760) <= not a or b;
    layer4_outputs(761) <= not b;
    layer4_outputs(762) <= not b;
    layer4_outputs(763) <= a or b;
    layer4_outputs(764) <= not (a and b);
    layer4_outputs(765) <= a;
    layer4_outputs(766) <= not a;
    layer4_outputs(767) <= a or b;
    layer4_outputs(768) <= not b;
    layer4_outputs(769) <= a or b;
    layer4_outputs(770) <= not b;
    layer4_outputs(771) <= not (a and b);
    layer4_outputs(772) <= a;
    layer4_outputs(773) <= a or b;
    layer4_outputs(774) <= a and b;
    layer4_outputs(775) <= not b or a;
    layer4_outputs(776) <= a xor b;
    layer4_outputs(777) <= not a or b;
    layer4_outputs(778) <= b and not a;
    layer4_outputs(779) <= not (a xor b);
    layer4_outputs(780) <= not a;
    layer4_outputs(781) <= not a;
    layer4_outputs(782) <= '0';
    layer4_outputs(783) <= not (a and b);
    layer4_outputs(784) <= a and b;
    layer4_outputs(785) <= '1';
    layer4_outputs(786) <= not (a or b);
    layer4_outputs(787) <= not (a xor b);
    layer4_outputs(788) <= not a or b;
    layer4_outputs(789) <= a;
    layer4_outputs(790) <= b;
    layer4_outputs(791) <= a xor b;
    layer4_outputs(792) <= not a;
    layer4_outputs(793) <= not b;
    layer4_outputs(794) <= a xor b;
    layer4_outputs(795) <= not a;
    layer4_outputs(796) <= a or b;
    layer4_outputs(797) <= b;
    layer4_outputs(798) <= a or b;
    layer4_outputs(799) <= b;
    layer4_outputs(800) <= a and b;
    layer4_outputs(801) <= not b;
    layer4_outputs(802) <= not (a or b);
    layer4_outputs(803) <= b;
    layer4_outputs(804) <= b;
    layer4_outputs(805) <= a;
    layer4_outputs(806) <= not (a and b);
    layer4_outputs(807) <= not a;
    layer4_outputs(808) <= a or b;
    layer4_outputs(809) <= not a or b;
    layer4_outputs(810) <= a;
    layer4_outputs(811) <= not (a or b);
    layer4_outputs(812) <= a;
    layer4_outputs(813) <= not (a or b);
    layer4_outputs(814) <= '1';
    layer4_outputs(815) <= b and not a;
    layer4_outputs(816) <= b;
    layer4_outputs(817) <= b;
    layer4_outputs(818) <= b;
    layer4_outputs(819) <= not b or a;
    layer4_outputs(820) <= not a;
    layer4_outputs(821) <= not b;
    layer4_outputs(822) <= not a;
    layer4_outputs(823) <= a;
    layer4_outputs(824) <= not b;
    layer4_outputs(825) <= not a;
    layer4_outputs(826) <= not a or b;
    layer4_outputs(827) <= a and not b;
    layer4_outputs(828) <= a;
    layer4_outputs(829) <= not b;
    layer4_outputs(830) <= b and not a;
    layer4_outputs(831) <= not b or a;
    layer4_outputs(832) <= not a;
    layer4_outputs(833) <= b and not a;
    layer4_outputs(834) <= b;
    layer4_outputs(835) <= b and not a;
    layer4_outputs(836) <= '0';
    layer4_outputs(837) <= not b;
    layer4_outputs(838) <= a;
    layer4_outputs(839) <= '1';
    layer4_outputs(840) <= not a;
    layer4_outputs(841) <= a or b;
    layer4_outputs(842) <= a and b;
    layer4_outputs(843) <= not (a and b);
    layer4_outputs(844) <= a xor b;
    layer4_outputs(845) <= b;
    layer4_outputs(846) <= b;
    layer4_outputs(847) <= a xor b;
    layer4_outputs(848) <= b;
    layer4_outputs(849) <= not (a xor b);
    layer4_outputs(850) <= not b or a;
    layer4_outputs(851) <= not a;
    layer4_outputs(852) <= not b or a;
    layer4_outputs(853) <= b and not a;
    layer4_outputs(854) <= not a or b;
    layer4_outputs(855) <= not (a xor b);
    layer4_outputs(856) <= a;
    layer4_outputs(857) <= a and not b;
    layer4_outputs(858) <= not b or a;
    layer4_outputs(859) <= not b;
    layer4_outputs(860) <= not b or a;
    layer4_outputs(861) <= not (a or b);
    layer4_outputs(862) <= not (a or b);
    layer4_outputs(863) <= a xor b;
    layer4_outputs(864) <= not b;
    layer4_outputs(865) <= b and not a;
    layer4_outputs(866) <= not b;
    layer4_outputs(867) <= not b or a;
    layer4_outputs(868) <= not (a or b);
    layer4_outputs(869) <= not b;
    layer4_outputs(870) <= a or b;
    layer4_outputs(871) <= not a or b;
    layer4_outputs(872) <= a xor b;
    layer4_outputs(873) <= a xor b;
    layer4_outputs(874) <= b and not a;
    layer4_outputs(875) <= a and b;
    layer4_outputs(876) <= not (a or b);
    layer4_outputs(877) <= not b;
    layer4_outputs(878) <= not (a or b);
    layer4_outputs(879) <= a and b;
    layer4_outputs(880) <= not (a xor b);
    layer4_outputs(881) <= a;
    layer4_outputs(882) <= b;
    layer4_outputs(883) <= b and not a;
    layer4_outputs(884) <= b and not a;
    layer4_outputs(885) <= a;
    layer4_outputs(886) <= a;
    layer4_outputs(887) <= a or b;
    layer4_outputs(888) <= b and not a;
    layer4_outputs(889) <= not b or a;
    layer4_outputs(890) <= a;
    layer4_outputs(891) <= '0';
    layer4_outputs(892) <= a and b;
    layer4_outputs(893) <= not b;
    layer4_outputs(894) <= a;
    layer4_outputs(895) <= a;
    layer4_outputs(896) <= not b;
    layer4_outputs(897) <= not a;
    layer4_outputs(898) <= '0';
    layer4_outputs(899) <= a xor b;
    layer4_outputs(900) <= a or b;
    layer4_outputs(901) <= b;
    layer4_outputs(902) <= a;
    layer4_outputs(903) <= b;
    layer4_outputs(904) <= b and not a;
    layer4_outputs(905) <= a and b;
    layer4_outputs(906) <= not a or b;
    layer4_outputs(907) <= not (a and b);
    layer4_outputs(908) <= not (a xor b);
    layer4_outputs(909) <= not a;
    layer4_outputs(910) <= not b;
    layer4_outputs(911) <= not b or a;
    layer4_outputs(912) <= not b;
    layer4_outputs(913) <= a;
    layer4_outputs(914) <= not (a xor b);
    layer4_outputs(915) <= not b;
    layer4_outputs(916) <= not (a or b);
    layer4_outputs(917) <= b and not a;
    layer4_outputs(918) <= not (a or b);
    layer4_outputs(919) <= a xor b;
    layer4_outputs(920) <= not (a or b);
    layer4_outputs(921) <= not b or a;
    layer4_outputs(922) <= a or b;
    layer4_outputs(923) <= b;
    layer4_outputs(924) <= not a;
    layer4_outputs(925) <= a;
    layer4_outputs(926) <= not (a and b);
    layer4_outputs(927) <= b and not a;
    layer4_outputs(928) <= b;
    layer4_outputs(929) <= a xor b;
    layer4_outputs(930) <= b;
    layer4_outputs(931) <= a;
    layer4_outputs(932) <= a or b;
    layer4_outputs(933) <= not (a and b);
    layer4_outputs(934) <= b and not a;
    layer4_outputs(935) <= a and not b;
    layer4_outputs(936) <= a and not b;
    layer4_outputs(937) <= not a;
    layer4_outputs(938) <= b;
    layer4_outputs(939) <= not b;
    layer4_outputs(940) <= not (a and b);
    layer4_outputs(941) <= a and not b;
    layer4_outputs(942) <= a xor b;
    layer4_outputs(943) <= a and b;
    layer4_outputs(944) <= not b;
    layer4_outputs(945) <= not b;
    layer4_outputs(946) <= a;
    layer4_outputs(947) <= b;
    layer4_outputs(948) <= not b or a;
    layer4_outputs(949) <= not (a and b);
    layer4_outputs(950) <= a and b;
    layer4_outputs(951) <= b and not a;
    layer4_outputs(952) <= a;
    layer4_outputs(953) <= a;
    layer4_outputs(954) <= not b;
    layer4_outputs(955) <= not a;
    layer4_outputs(956) <= a or b;
    layer4_outputs(957) <= not a;
    layer4_outputs(958) <= a;
    layer4_outputs(959) <= a or b;
    layer4_outputs(960) <= a and b;
    layer4_outputs(961) <= '1';
    layer4_outputs(962) <= not a;
    layer4_outputs(963) <= not a or b;
    layer4_outputs(964) <= not a or b;
    layer4_outputs(965) <= not b;
    layer4_outputs(966) <= a and not b;
    layer4_outputs(967) <= a and not b;
    layer4_outputs(968) <= a;
    layer4_outputs(969) <= not (a xor b);
    layer4_outputs(970) <= not (a and b);
    layer4_outputs(971) <= not a;
    layer4_outputs(972) <= not a;
    layer4_outputs(973) <= not b;
    layer4_outputs(974) <= a xor b;
    layer4_outputs(975) <= b and not a;
    layer4_outputs(976) <= not (a xor b);
    layer4_outputs(977) <= not b or a;
    layer4_outputs(978) <= b and not a;
    layer4_outputs(979) <= a or b;
    layer4_outputs(980) <= a;
    layer4_outputs(981) <= a and b;
    layer4_outputs(982) <= a and b;
    layer4_outputs(983) <= b and not a;
    layer4_outputs(984) <= a or b;
    layer4_outputs(985) <= not a;
    layer4_outputs(986) <= not a;
    layer4_outputs(987) <= a and not b;
    layer4_outputs(988) <= b and not a;
    layer4_outputs(989) <= a and b;
    layer4_outputs(990) <= a and not b;
    layer4_outputs(991) <= not (a xor b);
    layer4_outputs(992) <= not a;
    layer4_outputs(993) <= b;
    layer4_outputs(994) <= a;
    layer4_outputs(995) <= b;
    layer4_outputs(996) <= not a or b;
    layer4_outputs(997) <= a xor b;
    layer4_outputs(998) <= b;
    layer4_outputs(999) <= a or b;
    layer4_outputs(1000) <= a;
    layer4_outputs(1001) <= b;
    layer4_outputs(1002) <= b;
    layer4_outputs(1003) <= not b;
    layer4_outputs(1004) <= not (a xor b);
    layer4_outputs(1005) <= not (a and b);
    layer4_outputs(1006) <= not (a and b);
    layer4_outputs(1007) <= not a or b;
    layer4_outputs(1008) <= a;
    layer4_outputs(1009) <= a;
    layer4_outputs(1010) <= a and b;
    layer4_outputs(1011) <= b and not a;
    layer4_outputs(1012) <= a xor b;
    layer4_outputs(1013) <= not b;
    layer4_outputs(1014) <= b;
    layer4_outputs(1015) <= a and b;
    layer4_outputs(1016) <= b and not a;
    layer4_outputs(1017) <= not (a or b);
    layer4_outputs(1018) <= not a;
    layer4_outputs(1019) <= not (a or b);
    layer4_outputs(1020) <= a;
    layer4_outputs(1021) <= a or b;
    layer4_outputs(1022) <= a xor b;
    layer4_outputs(1023) <= not (a xor b);
    layer4_outputs(1024) <= a or b;
    layer4_outputs(1025) <= not (a xor b);
    layer4_outputs(1026) <= not a;
    layer4_outputs(1027) <= '0';
    layer4_outputs(1028) <= not b;
    layer4_outputs(1029) <= not (a and b);
    layer4_outputs(1030) <= a and not b;
    layer4_outputs(1031) <= not a;
    layer4_outputs(1032) <= b and not a;
    layer4_outputs(1033) <= not b;
    layer4_outputs(1034) <= b;
    layer4_outputs(1035) <= not b or a;
    layer4_outputs(1036) <= not a;
    layer4_outputs(1037) <= a;
    layer4_outputs(1038) <= b and not a;
    layer4_outputs(1039) <= b and not a;
    layer4_outputs(1040) <= a and b;
    layer4_outputs(1041) <= b;
    layer4_outputs(1042) <= not (a xor b);
    layer4_outputs(1043) <= a or b;
    layer4_outputs(1044) <= a;
    layer4_outputs(1045) <= not b;
    layer4_outputs(1046) <= not (a and b);
    layer4_outputs(1047) <= b;
    layer4_outputs(1048) <= a xor b;
    layer4_outputs(1049) <= not b or a;
    layer4_outputs(1050) <= not b or a;
    layer4_outputs(1051) <= not a;
    layer4_outputs(1052) <= not a or b;
    layer4_outputs(1053) <= not (a or b);
    layer4_outputs(1054) <= not a;
    layer4_outputs(1055) <= a;
    layer4_outputs(1056) <= a xor b;
    layer4_outputs(1057) <= a and b;
    layer4_outputs(1058) <= not (a or b);
    layer4_outputs(1059) <= a;
    layer4_outputs(1060) <= not a;
    layer4_outputs(1061) <= a and b;
    layer4_outputs(1062) <= a and not b;
    layer4_outputs(1063) <= not b or a;
    layer4_outputs(1064) <= not a or b;
    layer4_outputs(1065) <= not b or a;
    layer4_outputs(1066) <= not (a or b);
    layer4_outputs(1067) <= not b or a;
    layer4_outputs(1068) <= a and b;
    layer4_outputs(1069) <= a and b;
    layer4_outputs(1070) <= not (a or b);
    layer4_outputs(1071) <= not b or a;
    layer4_outputs(1072) <= not (a xor b);
    layer4_outputs(1073) <= not b;
    layer4_outputs(1074) <= a;
    layer4_outputs(1075) <= a xor b;
    layer4_outputs(1076) <= a;
    layer4_outputs(1077) <= b;
    layer4_outputs(1078) <= not a or b;
    layer4_outputs(1079) <= a and not b;
    layer4_outputs(1080) <= a and not b;
    layer4_outputs(1081) <= not b or a;
    layer4_outputs(1082) <= not a;
    layer4_outputs(1083) <= not b or a;
    layer4_outputs(1084) <= '1';
    layer4_outputs(1085) <= not a;
    layer4_outputs(1086) <= a xor b;
    layer4_outputs(1087) <= not a;
    layer4_outputs(1088) <= a xor b;
    layer4_outputs(1089) <= not (a and b);
    layer4_outputs(1090) <= b;
    layer4_outputs(1091) <= b and not a;
    layer4_outputs(1092) <= not a or b;
    layer4_outputs(1093) <= not a;
    layer4_outputs(1094) <= not (a xor b);
    layer4_outputs(1095) <= a;
    layer4_outputs(1096) <= b and not a;
    layer4_outputs(1097) <= a and not b;
    layer4_outputs(1098) <= not b;
    layer4_outputs(1099) <= not (a and b);
    layer4_outputs(1100) <= a xor b;
    layer4_outputs(1101) <= a or b;
    layer4_outputs(1102) <= not b;
    layer4_outputs(1103) <= not (a xor b);
    layer4_outputs(1104) <= not a or b;
    layer4_outputs(1105) <= a and not b;
    layer4_outputs(1106) <= not a;
    layer4_outputs(1107) <= '0';
    layer4_outputs(1108) <= b;
    layer4_outputs(1109) <= a and not b;
    layer4_outputs(1110) <= b and not a;
    layer4_outputs(1111) <= b and not a;
    layer4_outputs(1112) <= a and b;
    layer4_outputs(1113) <= not (a or b);
    layer4_outputs(1114) <= not b;
    layer4_outputs(1115) <= a or b;
    layer4_outputs(1116) <= not a;
    layer4_outputs(1117) <= not (a xor b);
    layer4_outputs(1118) <= a and b;
    layer4_outputs(1119) <= a and b;
    layer4_outputs(1120) <= not b or a;
    layer4_outputs(1121) <= b;
    layer4_outputs(1122) <= b and not a;
    layer4_outputs(1123) <= not a;
    layer4_outputs(1124) <= not b;
    layer4_outputs(1125) <= a;
    layer4_outputs(1126) <= b;
    layer4_outputs(1127) <= b and not a;
    layer4_outputs(1128) <= not a;
    layer4_outputs(1129) <= not a or b;
    layer4_outputs(1130) <= b and not a;
    layer4_outputs(1131) <= not (a or b);
    layer4_outputs(1132) <= not b or a;
    layer4_outputs(1133) <= not b;
    layer4_outputs(1134) <= a and b;
    layer4_outputs(1135) <= not (a or b);
    layer4_outputs(1136) <= a and not b;
    layer4_outputs(1137) <= b;
    layer4_outputs(1138) <= not b;
    layer4_outputs(1139) <= b;
    layer4_outputs(1140) <= b;
    layer4_outputs(1141) <= b;
    layer4_outputs(1142) <= a and not b;
    layer4_outputs(1143) <= a and not b;
    layer4_outputs(1144) <= a;
    layer4_outputs(1145) <= b and not a;
    layer4_outputs(1146) <= not (a and b);
    layer4_outputs(1147) <= a xor b;
    layer4_outputs(1148) <= not (a or b);
    layer4_outputs(1149) <= not b or a;
    layer4_outputs(1150) <= not (a and b);
    layer4_outputs(1151) <= not (a and b);
    layer4_outputs(1152) <= a or b;
    layer4_outputs(1153) <= b;
    layer4_outputs(1154) <= not a;
    layer4_outputs(1155) <= a or b;
    layer4_outputs(1156) <= not (a xor b);
    layer4_outputs(1157) <= a;
    layer4_outputs(1158) <= not b or a;
    layer4_outputs(1159) <= not (a and b);
    layer4_outputs(1160) <= not a;
    layer4_outputs(1161) <= not b;
    layer4_outputs(1162) <= b and not a;
    layer4_outputs(1163) <= a;
    layer4_outputs(1164) <= a xor b;
    layer4_outputs(1165) <= a and b;
    layer4_outputs(1166) <= not (a or b);
    layer4_outputs(1167) <= b;
    layer4_outputs(1168) <= not b or a;
    layer4_outputs(1169) <= a and not b;
    layer4_outputs(1170) <= not (a xor b);
    layer4_outputs(1171) <= not (a or b);
    layer4_outputs(1172) <= a and b;
    layer4_outputs(1173) <= not a;
    layer4_outputs(1174) <= not b;
    layer4_outputs(1175) <= not b;
    layer4_outputs(1176) <= not b or a;
    layer4_outputs(1177) <= not b;
    layer4_outputs(1178) <= a xor b;
    layer4_outputs(1179) <= a or b;
    layer4_outputs(1180) <= not b or a;
    layer4_outputs(1181) <= a or b;
    layer4_outputs(1182) <= not a;
    layer4_outputs(1183) <= a xor b;
    layer4_outputs(1184) <= not a;
    layer4_outputs(1185) <= a xor b;
    layer4_outputs(1186) <= b;
    layer4_outputs(1187) <= not a or b;
    layer4_outputs(1188) <= a and b;
    layer4_outputs(1189) <= not (a and b);
    layer4_outputs(1190) <= not a;
    layer4_outputs(1191) <= a xor b;
    layer4_outputs(1192) <= not a;
    layer4_outputs(1193) <= a xor b;
    layer4_outputs(1194) <= b;
    layer4_outputs(1195) <= b;
    layer4_outputs(1196) <= a and not b;
    layer4_outputs(1197) <= not a;
    layer4_outputs(1198) <= not b or a;
    layer4_outputs(1199) <= not a;
    layer4_outputs(1200) <= a and b;
    layer4_outputs(1201) <= b;
    layer4_outputs(1202) <= a and b;
    layer4_outputs(1203) <= a;
    layer4_outputs(1204) <= not b;
    layer4_outputs(1205) <= not b;
    layer4_outputs(1206) <= '1';
    layer4_outputs(1207) <= not a or b;
    layer4_outputs(1208) <= a;
    layer4_outputs(1209) <= a and not b;
    layer4_outputs(1210) <= a or b;
    layer4_outputs(1211) <= a and not b;
    layer4_outputs(1212) <= not (a and b);
    layer4_outputs(1213) <= a;
    layer4_outputs(1214) <= a or b;
    layer4_outputs(1215) <= not (a and b);
    layer4_outputs(1216) <= not b;
    layer4_outputs(1217) <= not b;
    layer4_outputs(1218) <= b;
    layer4_outputs(1219) <= not (a or b);
    layer4_outputs(1220) <= not a or b;
    layer4_outputs(1221) <= not b;
    layer4_outputs(1222) <= a xor b;
    layer4_outputs(1223) <= a xor b;
    layer4_outputs(1224) <= a;
    layer4_outputs(1225) <= b and not a;
    layer4_outputs(1226) <= not (a or b);
    layer4_outputs(1227) <= a and not b;
    layer4_outputs(1228) <= not a;
    layer4_outputs(1229) <= not (a xor b);
    layer4_outputs(1230) <= not a;
    layer4_outputs(1231) <= b;
    layer4_outputs(1232) <= a or b;
    layer4_outputs(1233) <= a xor b;
    layer4_outputs(1234) <= not b;
    layer4_outputs(1235) <= not a;
    layer4_outputs(1236) <= not a or b;
    layer4_outputs(1237) <= a xor b;
    layer4_outputs(1238) <= b;
    layer4_outputs(1239) <= not (a and b);
    layer4_outputs(1240) <= a xor b;
    layer4_outputs(1241) <= a and not b;
    layer4_outputs(1242) <= a;
    layer4_outputs(1243) <= a and not b;
    layer4_outputs(1244) <= not a;
    layer4_outputs(1245) <= a and b;
    layer4_outputs(1246) <= a xor b;
    layer4_outputs(1247) <= not a;
    layer4_outputs(1248) <= b;
    layer4_outputs(1249) <= not (a or b);
    layer4_outputs(1250) <= b;
    layer4_outputs(1251) <= a or b;
    layer4_outputs(1252) <= not b or a;
    layer4_outputs(1253) <= not b;
    layer4_outputs(1254) <= a;
    layer4_outputs(1255) <= b;
    layer4_outputs(1256) <= a;
    layer4_outputs(1257) <= not a;
    layer4_outputs(1258) <= not a;
    layer4_outputs(1259) <= not b;
    layer4_outputs(1260) <= a xor b;
    layer4_outputs(1261) <= b;
    layer4_outputs(1262) <= a xor b;
    layer4_outputs(1263) <= a or b;
    layer4_outputs(1264) <= a;
    layer4_outputs(1265) <= not b or a;
    layer4_outputs(1266) <= not b;
    layer4_outputs(1267) <= not (a and b);
    layer4_outputs(1268) <= not a;
    layer4_outputs(1269) <= a and b;
    layer4_outputs(1270) <= not b;
    layer4_outputs(1271) <= a;
    layer4_outputs(1272) <= not (a xor b);
    layer4_outputs(1273) <= a and b;
    layer4_outputs(1274) <= not b;
    layer4_outputs(1275) <= a;
    layer4_outputs(1276) <= b;
    layer4_outputs(1277) <= not b;
    layer4_outputs(1278) <= a;
    layer4_outputs(1279) <= not b;
    layer4_outputs(1280) <= b;
    layer4_outputs(1281) <= a xor b;
    layer4_outputs(1282) <= a xor b;
    layer4_outputs(1283) <= a and not b;
    layer4_outputs(1284) <= b and not a;
    layer4_outputs(1285) <= not b or a;
    layer4_outputs(1286) <= a;
    layer4_outputs(1287) <= b;
    layer4_outputs(1288) <= a;
    layer4_outputs(1289) <= not b;
    layer4_outputs(1290) <= b;
    layer4_outputs(1291) <= b and not a;
    layer4_outputs(1292) <= not b;
    layer4_outputs(1293) <= b;
    layer4_outputs(1294) <= not b;
    layer4_outputs(1295) <= not (a or b);
    layer4_outputs(1296) <= not a;
    layer4_outputs(1297) <= b;
    layer4_outputs(1298) <= b;
    layer4_outputs(1299) <= b;
    layer4_outputs(1300) <= not a;
    layer4_outputs(1301) <= a or b;
    layer4_outputs(1302) <= b and not a;
    layer4_outputs(1303) <= not a;
    layer4_outputs(1304) <= not (a and b);
    layer4_outputs(1305) <= b;
    layer4_outputs(1306) <= not a;
    layer4_outputs(1307) <= not (a or b);
    layer4_outputs(1308) <= not a;
    layer4_outputs(1309) <= not (a xor b);
    layer4_outputs(1310) <= not b;
    layer4_outputs(1311) <= b;
    layer4_outputs(1312) <= a;
    layer4_outputs(1313) <= a;
    layer4_outputs(1314) <= not (a xor b);
    layer4_outputs(1315) <= not (a xor b);
    layer4_outputs(1316) <= not b or a;
    layer4_outputs(1317) <= b and not a;
    layer4_outputs(1318) <= b and not a;
    layer4_outputs(1319) <= not (a or b);
    layer4_outputs(1320) <= a and not b;
    layer4_outputs(1321) <= b and not a;
    layer4_outputs(1322) <= not b or a;
    layer4_outputs(1323) <= not (a or b);
    layer4_outputs(1324) <= a or b;
    layer4_outputs(1325) <= not a or b;
    layer4_outputs(1326) <= a and b;
    layer4_outputs(1327) <= a;
    layer4_outputs(1328) <= b and not a;
    layer4_outputs(1329) <= b and not a;
    layer4_outputs(1330) <= not (a and b);
    layer4_outputs(1331) <= a xor b;
    layer4_outputs(1332) <= a and not b;
    layer4_outputs(1333) <= a or b;
    layer4_outputs(1334) <= b;
    layer4_outputs(1335) <= a;
    layer4_outputs(1336) <= b;
    layer4_outputs(1337) <= a;
    layer4_outputs(1338) <= a and not b;
    layer4_outputs(1339) <= not a;
    layer4_outputs(1340) <= b;
    layer4_outputs(1341) <= a;
    layer4_outputs(1342) <= b and not a;
    layer4_outputs(1343) <= a xor b;
    layer4_outputs(1344) <= a xor b;
    layer4_outputs(1345) <= not (a or b);
    layer4_outputs(1346) <= a xor b;
    layer4_outputs(1347) <= a or b;
    layer4_outputs(1348) <= a and not b;
    layer4_outputs(1349) <= not (a xor b);
    layer4_outputs(1350) <= b;
    layer4_outputs(1351) <= a and b;
    layer4_outputs(1352) <= a or b;
    layer4_outputs(1353) <= not (a xor b);
    layer4_outputs(1354) <= not b or a;
    layer4_outputs(1355) <= not (a or b);
    layer4_outputs(1356) <= b and not a;
    layer4_outputs(1357) <= not (a or b);
    layer4_outputs(1358) <= not b;
    layer4_outputs(1359) <= not (a or b);
    layer4_outputs(1360) <= a;
    layer4_outputs(1361) <= a and not b;
    layer4_outputs(1362) <= not (a or b);
    layer4_outputs(1363) <= b;
    layer4_outputs(1364) <= a or b;
    layer4_outputs(1365) <= not b or a;
    layer4_outputs(1366) <= not (a and b);
    layer4_outputs(1367) <= not a;
    layer4_outputs(1368) <= not (a and b);
    layer4_outputs(1369) <= a or b;
    layer4_outputs(1370) <= not (a or b);
    layer4_outputs(1371) <= not a or b;
    layer4_outputs(1372) <= a and b;
    layer4_outputs(1373) <= not a;
    layer4_outputs(1374) <= not (a xor b);
    layer4_outputs(1375) <= not a or b;
    layer4_outputs(1376) <= not b;
    layer4_outputs(1377) <= b and not a;
    layer4_outputs(1378) <= a and b;
    layer4_outputs(1379) <= a and not b;
    layer4_outputs(1380) <= not (a and b);
    layer4_outputs(1381) <= not b;
    layer4_outputs(1382) <= not (a and b);
    layer4_outputs(1383) <= not a;
    layer4_outputs(1384) <= a;
    layer4_outputs(1385) <= not b or a;
    layer4_outputs(1386) <= not b;
    layer4_outputs(1387) <= not b;
    layer4_outputs(1388) <= b and not a;
    layer4_outputs(1389) <= a xor b;
    layer4_outputs(1390) <= b;
    layer4_outputs(1391) <= not b;
    layer4_outputs(1392) <= b;
    layer4_outputs(1393) <= not a;
    layer4_outputs(1394) <= not (a and b);
    layer4_outputs(1395) <= not a or b;
    layer4_outputs(1396) <= not a or b;
    layer4_outputs(1397) <= a or b;
    layer4_outputs(1398) <= not a;
    layer4_outputs(1399) <= not (a xor b);
    layer4_outputs(1400) <= a;
    layer4_outputs(1401) <= a and not b;
    layer4_outputs(1402) <= not (a or b);
    layer4_outputs(1403) <= b;
    layer4_outputs(1404) <= a xor b;
    layer4_outputs(1405) <= a;
    layer4_outputs(1406) <= a and not b;
    layer4_outputs(1407) <= b and not a;
    layer4_outputs(1408) <= not (a or b);
    layer4_outputs(1409) <= b;
    layer4_outputs(1410) <= b;
    layer4_outputs(1411) <= a and b;
    layer4_outputs(1412) <= b;
    layer4_outputs(1413) <= a or b;
    layer4_outputs(1414) <= a or b;
    layer4_outputs(1415) <= not (a xor b);
    layer4_outputs(1416) <= b;
    layer4_outputs(1417) <= not (a or b);
    layer4_outputs(1418) <= a xor b;
    layer4_outputs(1419) <= not a;
    layer4_outputs(1420) <= a and not b;
    layer4_outputs(1421) <= not (a xor b);
    layer4_outputs(1422) <= a and b;
    layer4_outputs(1423) <= a or b;
    layer4_outputs(1424) <= '1';
    layer4_outputs(1425) <= not (a and b);
    layer4_outputs(1426) <= '1';
    layer4_outputs(1427) <= b and not a;
    layer4_outputs(1428) <= not b;
    layer4_outputs(1429) <= a and not b;
    layer4_outputs(1430) <= not (a or b);
    layer4_outputs(1431) <= '1';
    layer4_outputs(1432) <= not (a or b);
    layer4_outputs(1433) <= not (a or b);
    layer4_outputs(1434) <= not a;
    layer4_outputs(1435) <= not b;
    layer4_outputs(1436) <= a xor b;
    layer4_outputs(1437) <= not (a or b);
    layer4_outputs(1438) <= not b;
    layer4_outputs(1439) <= not (a and b);
    layer4_outputs(1440) <= a and b;
    layer4_outputs(1441) <= a and not b;
    layer4_outputs(1442) <= not (a or b);
    layer4_outputs(1443) <= not (a and b);
    layer4_outputs(1444) <= a or b;
    layer4_outputs(1445) <= a and not b;
    layer4_outputs(1446) <= not (a xor b);
    layer4_outputs(1447) <= b;
    layer4_outputs(1448) <= not a;
    layer4_outputs(1449) <= not b or a;
    layer4_outputs(1450) <= not b;
    layer4_outputs(1451) <= not (a xor b);
    layer4_outputs(1452) <= a and b;
    layer4_outputs(1453) <= b;
    layer4_outputs(1454) <= a xor b;
    layer4_outputs(1455) <= not b;
    layer4_outputs(1456) <= a;
    layer4_outputs(1457) <= not (a or b);
    layer4_outputs(1458) <= b;
    layer4_outputs(1459) <= not (a or b);
    layer4_outputs(1460) <= a and not b;
    layer4_outputs(1461) <= b;
    layer4_outputs(1462) <= not a;
    layer4_outputs(1463) <= a and not b;
    layer4_outputs(1464) <= not (a xor b);
    layer4_outputs(1465) <= not b;
    layer4_outputs(1466) <= not a;
    layer4_outputs(1467) <= a;
    layer4_outputs(1468) <= not b;
    layer4_outputs(1469) <= not (a and b);
    layer4_outputs(1470) <= not a;
    layer4_outputs(1471) <= a;
    layer4_outputs(1472) <= not a;
    layer4_outputs(1473) <= b and not a;
    layer4_outputs(1474) <= not b;
    layer4_outputs(1475) <= not (a xor b);
    layer4_outputs(1476) <= a;
    layer4_outputs(1477) <= a and b;
    layer4_outputs(1478) <= a and b;
    layer4_outputs(1479) <= not (a or b);
    layer4_outputs(1480) <= a;
    layer4_outputs(1481) <= not b or a;
    layer4_outputs(1482) <= not (a and b);
    layer4_outputs(1483) <= b and not a;
    layer4_outputs(1484) <= a or b;
    layer4_outputs(1485) <= a and b;
    layer4_outputs(1486) <= not (a or b);
    layer4_outputs(1487) <= b and not a;
    layer4_outputs(1488) <= b;
    layer4_outputs(1489) <= not (a xor b);
    layer4_outputs(1490) <= b and not a;
    layer4_outputs(1491) <= a and not b;
    layer4_outputs(1492) <= not a or b;
    layer4_outputs(1493) <= a;
    layer4_outputs(1494) <= not b;
    layer4_outputs(1495) <= not (a and b);
    layer4_outputs(1496) <= not b;
    layer4_outputs(1497) <= b;
    layer4_outputs(1498) <= b;
    layer4_outputs(1499) <= not b;
    layer4_outputs(1500) <= a;
    layer4_outputs(1501) <= b and not a;
    layer4_outputs(1502) <= a or b;
    layer4_outputs(1503) <= not b;
    layer4_outputs(1504) <= a or b;
    layer4_outputs(1505) <= not (a xor b);
    layer4_outputs(1506) <= not b;
    layer4_outputs(1507) <= not a or b;
    layer4_outputs(1508) <= b;
    layer4_outputs(1509) <= not b;
    layer4_outputs(1510) <= not b or a;
    layer4_outputs(1511) <= a or b;
    layer4_outputs(1512) <= not a;
    layer4_outputs(1513) <= a and not b;
    layer4_outputs(1514) <= a;
    layer4_outputs(1515) <= a and b;
    layer4_outputs(1516) <= b;
    layer4_outputs(1517) <= a xor b;
    layer4_outputs(1518) <= a;
    layer4_outputs(1519) <= a xor b;
    layer4_outputs(1520) <= a;
    layer4_outputs(1521) <= a;
    layer4_outputs(1522) <= not (a or b);
    layer4_outputs(1523) <= not (a and b);
    layer4_outputs(1524) <= b and not a;
    layer4_outputs(1525) <= not a or b;
    layer4_outputs(1526) <= a xor b;
    layer4_outputs(1527) <= b;
    layer4_outputs(1528) <= not a or b;
    layer4_outputs(1529) <= a;
    layer4_outputs(1530) <= a;
    layer4_outputs(1531) <= b;
    layer4_outputs(1532) <= a;
    layer4_outputs(1533) <= b;
    layer4_outputs(1534) <= a and b;
    layer4_outputs(1535) <= a and not b;
    layer4_outputs(1536) <= b;
    layer4_outputs(1537) <= a or b;
    layer4_outputs(1538) <= b and not a;
    layer4_outputs(1539) <= not (a and b);
    layer4_outputs(1540) <= not (a or b);
    layer4_outputs(1541) <= not b;
    layer4_outputs(1542) <= a xor b;
    layer4_outputs(1543) <= a;
    layer4_outputs(1544) <= a and b;
    layer4_outputs(1545) <= not (a and b);
    layer4_outputs(1546) <= not b or a;
    layer4_outputs(1547) <= a;
    layer4_outputs(1548) <= b;
    layer4_outputs(1549) <= not a or b;
    layer4_outputs(1550) <= not a;
    layer4_outputs(1551) <= not (a xor b);
    layer4_outputs(1552) <= not b;
    layer4_outputs(1553) <= not a or b;
    layer4_outputs(1554) <= b;
    layer4_outputs(1555) <= b;
    layer4_outputs(1556) <= a xor b;
    layer4_outputs(1557) <= '1';
    layer4_outputs(1558) <= a or b;
    layer4_outputs(1559) <= b;
    layer4_outputs(1560) <= not b or a;
    layer4_outputs(1561) <= a xor b;
    layer4_outputs(1562) <= b;
    layer4_outputs(1563) <= a or b;
    layer4_outputs(1564) <= not b;
    layer4_outputs(1565) <= not (a xor b);
    layer4_outputs(1566) <= not b;
    layer4_outputs(1567) <= a and b;
    layer4_outputs(1568) <= not b;
    layer4_outputs(1569) <= b;
    layer4_outputs(1570) <= not (a xor b);
    layer4_outputs(1571) <= a and not b;
    layer4_outputs(1572) <= not a;
    layer4_outputs(1573) <= not (a and b);
    layer4_outputs(1574) <= a and not b;
    layer4_outputs(1575) <= '1';
    layer4_outputs(1576) <= not a;
    layer4_outputs(1577) <= a and b;
    layer4_outputs(1578) <= not b;
    layer4_outputs(1579) <= not (a xor b);
    layer4_outputs(1580) <= a;
    layer4_outputs(1581) <= not (a xor b);
    layer4_outputs(1582) <= a;
    layer4_outputs(1583) <= a;
    layer4_outputs(1584) <= a and not b;
    layer4_outputs(1585) <= a and b;
    layer4_outputs(1586) <= a;
    layer4_outputs(1587) <= not (a xor b);
    layer4_outputs(1588) <= not a;
    layer4_outputs(1589) <= not b or a;
    layer4_outputs(1590) <= not a;
    layer4_outputs(1591) <= a and not b;
    layer4_outputs(1592) <= not a or b;
    layer4_outputs(1593) <= not (a and b);
    layer4_outputs(1594) <= b and not a;
    layer4_outputs(1595) <= a;
    layer4_outputs(1596) <= b;
    layer4_outputs(1597) <= a;
    layer4_outputs(1598) <= not a;
    layer4_outputs(1599) <= not a;
    layer4_outputs(1600) <= b;
    layer4_outputs(1601) <= not a or b;
    layer4_outputs(1602) <= a;
    layer4_outputs(1603) <= not a;
    layer4_outputs(1604) <= not (a and b);
    layer4_outputs(1605) <= not b or a;
    layer4_outputs(1606) <= a and not b;
    layer4_outputs(1607) <= not (a and b);
    layer4_outputs(1608) <= not b;
    layer4_outputs(1609) <= not b or a;
    layer4_outputs(1610) <= a and not b;
    layer4_outputs(1611) <= a;
    layer4_outputs(1612) <= not b or a;
    layer4_outputs(1613) <= not b;
    layer4_outputs(1614) <= not (a or b);
    layer4_outputs(1615) <= a;
    layer4_outputs(1616) <= '0';
    layer4_outputs(1617) <= not a or b;
    layer4_outputs(1618) <= not (a and b);
    layer4_outputs(1619) <= a or b;
    layer4_outputs(1620) <= a and b;
    layer4_outputs(1621) <= b;
    layer4_outputs(1622) <= not a;
    layer4_outputs(1623) <= not (a and b);
    layer4_outputs(1624) <= b;
    layer4_outputs(1625) <= a xor b;
    layer4_outputs(1626) <= a and b;
    layer4_outputs(1627) <= a;
    layer4_outputs(1628) <= not b;
    layer4_outputs(1629) <= b;
    layer4_outputs(1630) <= a and not b;
    layer4_outputs(1631) <= a;
    layer4_outputs(1632) <= not a;
    layer4_outputs(1633) <= b;
    layer4_outputs(1634) <= not a;
    layer4_outputs(1635) <= b and not a;
    layer4_outputs(1636) <= not a;
    layer4_outputs(1637) <= not (a or b);
    layer4_outputs(1638) <= b;
    layer4_outputs(1639) <= not (a or b);
    layer4_outputs(1640) <= a or b;
    layer4_outputs(1641) <= not b;
    layer4_outputs(1642) <= not (a and b);
    layer4_outputs(1643) <= a;
    layer4_outputs(1644) <= a and not b;
    layer4_outputs(1645) <= a xor b;
    layer4_outputs(1646) <= b and not a;
    layer4_outputs(1647) <= a and not b;
    layer4_outputs(1648) <= not b;
    layer4_outputs(1649) <= not b;
    layer4_outputs(1650) <= a or b;
    layer4_outputs(1651) <= a;
    layer4_outputs(1652) <= not a;
    layer4_outputs(1653) <= b;
    layer4_outputs(1654) <= not (a xor b);
    layer4_outputs(1655) <= b and not a;
    layer4_outputs(1656) <= not b;
    layer4_outputs(1657) <= a;
    layer4_outputs(1658) <= b;
    layer4_outputs(1659) <= not a;
    layer4_outputs(1660) <= a and b;
    layer4_outputs(1661) <= a;
    layer4_outputs(1662) <= a and not b;
    layer4_outputs(1663) <= not (a and b);
    layer4_outputs(1664) <= a xor b;
    layer4_outputs(1665) <= not a or b;
    layer4_outputs(1666) <= a xor b;
    layer4_outputs(1667) <= not a;
    layer4_outputs(1668) <= a and not b;
    layer4_outputs(1669) <= a and b;
    layer4_outputs(1670) <= a or b;
    layer4_outputs(1671) <= a and not b;
    layer4_outputs(1672) <= not a;
    layer4_outputs(1673) <= b and not a;
    layer4_outputs(1674) <= a;
    layer4_outputs(1675) <= a or b;
    layer4_outputs(1676) <= not (a or b);
    layer4_outputs(1677) <= a and not b;
    layer4_outputs(1678) <= a;
    layer4_outputs(1679) <= a and not b;
    layer4_outputs(1680) <= a;
    layer4_outputs(1681) <= a and b;
    layer4_outputs(1682) <= a or b;
    layer4_outputs(1683) <= not a or b;
    layer4_outputs(1684) <= not (a or b);
    layer4_outputs(1685) <= a;
    layer4_outputs(1686) <= b;
    layer4_outputs(1687) <= not (a and b);
    layer4_outputs(1688) <= not (a or b);
    layer4_outputs(1689) <= a;
    layer4_outputs(1690) <= b and not a;
    layer4_outputs(1691) <= b;
    layer4_outputs(1692) <= not b;
    layer4_outputs(1693) <= not b;
    layer4_outputs(1694) <= not b;
    layer4_outputs(1695) <= b;
    layer4_outputs(1696) <= not a or b;
    layer4_outputs(1697) <= not a;
    layer4_outputs(1698) <= '0';
    layer4_outputs(1699) <= a or b;
    layer4_outputs(1700) <= not (a xor b);
    layer4_outputs(1701) <= not (a and b);
    layer4_outputs(1702) <= not (a xor b);
    layer4_outputs(1703) <= a;
    layer4_outputs(1704) <= a and not b;
    layer4_outputs(1705) <= b and not a;
    layer4_outputs(1706) <= not a;
    layer4_outputs(1707) <= not a;
    layer4_outputs(1708) <= a xor b;
    layer4_outputs(1709) <= not (a and b);
    layer4_outputs(1710) <= a xor b;
    layer4_outputs(1711) <= not (a xor b);
    layer4_outputs(1712) <= a and not b;
    layer4_outputs(1713) <= a;
    layer4_outputs(1714) <= a and b;
    layer4_outputs(1715) <= not b or a;
    layer4_outputs(1716) <= b;
    layer4_outputs(1717) <= not (a xor b);
    layer4_outputs(1718) <= b;
    layer4_outputs(1719) <= a;
    layer4_outputs(1720) <= a and b;
    layer4_outputs(1721) <= not a;
    layer4_outputs(1722) <= b and not a;
    layer4_outputs(1723) <= not (a or b);
    layer4_outputs(1724) <= b;
    layer4_outputs(1725) <= not (a xor b);
    layer4_outputs(1726) <= b;
    layer4_outputs(1727) <= a xor b;
    layer4_outputs(1728) <= not b;
    layer4_outputs(1729) <= a and not b;
    layer4_outputs(1730) <= a;
    layer4_outputs(1731) <= a and not b;
    layer4_outputs(1732) <= a;
    layer4_outputs(1733) <= not (a or b);
    layer4_outputs(1734) <= not (a or b);
    layer4_outputs(1735) <= a;
    layer4_outputs(1736) <= not a or b;
    layer4_outputs(1737) <= a and not b;
    layer4_outputs(1738) <= b;
    layer4_outputs(1739) <= not a or b;
    layer4_outputs(1740) <= not a;
    layer4_outputs(1741) <= not a;
    layer4_outputs(1742) <= a;
    layer4_outputs(1743) <= a;
    layer4_outputs(1744) <= a;
    layer4_outputs(1745) <= a and b;
    layer4_outputs(1746) <= not a;
    layer4_outputs(1747) <= not a or b;
    layer4_outputs(1748) <= not a or b;
    layer4_outputs(1749) <= b;
    layer4_outputs(1750) <= not a;
    layer4_outputs(1751) <= not b or a;
    layer4_outputs(1752) <= a;
    layer4_outputs(1753) <= not a;
    layer4_outputs(1754) <= not (a and b);
    layer4_outputs(1755) <= b and not a;
    layer4_outputs(1756) <= b;
    layer4_outputs(1757) <= not (a or b);
    layer4_outputs(1758) <= not a or b;
    layer4_outputs(1759) <= '0';
    layer4_outputs(1760) <= a;
    layer4_outputs(1761) <= not (a xor b);
    layer4_outputs(1762) <= not b or a;
    layer4_outputs(1763) <= not (a or b);
    layer4_outputs(1764) <= a;
    layer4_outputs(1765) <= not b;
    layer4_outputs(1766) <= b;
    layer4_outputs(1767) <= b and not a;
    layer4_outputs(1768) <= not b;
    layer4_outputs(1769) <= b;
    layer4_outputs(1770) <= not a;
    layer4_outputs(1771) <= b;
    layer4_outputs(1772) <= a;
    layer4_outputs(1773) <= b;
    layer4_outputs(1774) <= not a;
    layer4_outputs(1775) <= not (a and b);
    layer4_outputs(1776) <= not a or b;
    layer4_outputs(1777) <= not a;
    layer4_outputs(1778) <= a and b;
    layer4_outputs(1779) <= not (a and b);
    layer4_outputs(1780) <= not a;
    layer4_outputs(1781) <= a or b;
    layer4_outputs(1782) <= not a;
    layer4_outputs(1783) <= not a or b;
    layer4_outputs(1784) <= not a;
    layer4_outputs(1785) <= not a;
    layer4_outputs(1786) <= not a;
    layer4_outputs(1787) <= a;
    layer4_outputs(1788) <= not a;
    layer4_outputs(1789) <= not b;
    layer4_outputs(1790) <= not (a xor b);
    layer4_outputs(1791) <= not b;
    layer4_outputs(1792) <= not (a xor b);
    layer4_outputs(1793) <= not b or a;
    layer4_outputs(1794) <= not b;
    layer4_outputs(1795) <= a and b;
    layer4_outputs(1796) <= a;
    layer4_outputs(1797) <= a;
    layer4_outputs(1798) <= b;
    layer4_outputs(1799) <= not (a xor b);
    layer4_outputs(1800) <= b and not a;
    layer4_outputs(1801) <= b and not a;
    layer4_outputs(1802) <= b;
    layer4_outputs(1803) <= a or b;
    layer4_outputs(1804) <= a xor b;
    layer4_outputs(1805) <= a and b;
    layer4_outputs(1806) <= b and not a;
    layer4_outputs(1807) <= a;
    layer4_outputs(1808) <= a and not b;
    layer4_outputs(1809) <= a or b;
    layer4_outputs(1810) <= not a;
    layer4_outputs(1811) <= not (a and b);
    layer4_outputs(1812) <= not b or a;
    layer4_outputs(1813) <= not a or b;
    layer4_outputs(1814) <= a and not b;
    layer4_outputs(1815) <= a and not b;
    layer4_outputs(1816) <= not (a xor b);
    layer4_outputs(1817) <= not (a and b);
    layer4_outputs(1818) <= a and b;
    layer4_outputs(1819) <= a and b;
    layer4_outputs(1820) <= not (a and b);
    layer4_outputs(1821) <= not (a or b);
    layer4_outputs(1822) <= a and not b;
    layer4_outputs(1823) <= not a;
    layer4_outputs(1824) <= b;
    layer4_outputs(1825) <= a;
    layer4_outputs(1826) <= b and not a;
    layer4_outputs(1827) <= b and not a;
    layer4_outputs(1828) <= not b or a;
    layer4_outputs(1829) <= not b or a;
    layer4_outputs(1830) <= a and not b;
    layer4_outputs(1831) <= a or b;
    layer4_outputs(1832) <= b;
    layer4_outputs(1833) <= not b or a;
    layer4_outputs(1834) <= a;
    layer4_outputs(1835) <= a;
    layer4_outputs(1836) <= not a or b;
    layer4_outputs(1837) <= not b;
    layer4_outputs(1838) <= not (a or b);
    layer4_outputs(1839) <= a and b;
    layer4_outputs(1840) <= not a;
    layer4_outputs(1841) <= not (a or b);
    layer4_outputs(1842) <= not (a and b);
    layer4_outputs(1843) <= a;
    layer4_outputs(1844) <= not (a xor b);
    layer4_outputs(1845) <= not (a or b);
    layer4_outputs(1846) <= b;
    layer4_outputs(1847) <= not b;
    layer4_outputs(1848) <= a;
    layer4_outputs(1849) <= a xor b;
    layer4_outputs(1850) <= a;
    layer4_outputs(1851) <= a and b;
    layer4_outputs(1852) <= not a or b;
    layer4_outputs(1853) <= not b;
    layer4_outputs(1854) <= a and b;
    layer4_outputs(1855) <= not (a or b);
    layer4_outputs(1856) <= not a;
    layer4_outputs(1857) <= not (a xor b);
    layer4_outputs(1858) <= not (a or b);
    layer4_outputs(1859) <= not a;
    layer4_outputs(1860) <= a xor b;
    layer4_outputs(1861) <= not (a xor b);
    layer4_outputs(1862) <= not a;
    layer4_outputs(1863) <= not a;
    layer4_outputs(1864) <= not b or a;
    layer4_outputs(1865) <= b and not a;
    layer4_outputs(1866) <= not a;
    layer4_outputs(1867) <= not (a or b);
    layer4_outputs(1868) <= not b or a;
    layer4_outputs(1869) <= a and not b;
    layer4_outputs(1870) <= a and not b;
    layer4_outputs(1871) <= b;
    layer4_outputs(1872) <= not a or b;
    layer4_outputs(1873) <= a xor b;
    layer4_outputs(1874) <= a;
    layer4_outputs(1875) <= not b;
    layer4_outputs(1876) <= not b or a;
    layer4_outputs(1877) <= a;
    layer4_outputs(1878) <= not (a xor b);
    layer4_outputs(1879) <= b;
    layer4_outputs(1880) <= not (a xor b);
    layer4_outputs(1881) <= a;
    layer4_outputs(1882) <= not (a and b);
    layer4_outputs(1883) <= a and b;
    layer4_outputs(1884) <= not b or a;
    layer4_outputs(1885) <= b;
    layer4_outputs(1886) <= a;
    layer4_outputs(1887) <= a and b;
    layer4_outputs(1888) <= not (a xor b);
    layer4_outputs(1889) <= a;
    layer4_outputs(1890) <= not a or b;
    layer4_outputs(1891) <= a;
    layer4_outputs(1892) <= b;
    layer4_outputs(1893) <= not a;
    layer4_outputs(1894) <= not (a xor b);
    layer4_outputs(1895) <= a and not b;
    layer4_outputs(1896) <= not a;
    layer4_outputs(1897) <= a;
    layer4_outputs(1898) <= not b;
    layer4_outputs(1899) <= not a or b;
    layer4_outputs(1900) <= not a;
    layer4_outputs(1901) <= b and not a;
    layer4_outputs(1902) <= not b;
    layer4_outputs(1903) <= not (a or b);
    layer4_outputs(1904) <= not a;
    layer4_outputs(1905) <= not (a and b);
    layer4_outputs(1906) <= b and not a;
    layer4_outputs(1907) <= a;
    layer4_outputs(1908) <= not a or b;
    layer4_outputs(1909) <= a;
    layer4_outputs(1910) <= not a or b;
    layer4_outputs(1911) <= not a;
    layer4_outputs(1912) <= b and not a;
    layer4_outputs(1913) <= not a;
    layer4_outputs(1914) <= not (a or b);
    layer4_outputs(1915) <= a or b;
    layer4_outputs(1916) <= not b;
    layer4_outputs(1917) <= a;
    layer4_outputs(1918) <= a;
    layer4_outputs(1919) <= a;
    layer4_outputs(1920) <= a and not b;
    layer4_outputs(1921) <= '0';
    layer4_outputs(1922) <= not a;
    layer4_outputs(1923) <= not a;
    layer4_outputs(1924) <= a;
    layer4_outputs(1925) <= b;
    layer4_outputs(1926) <= b;
    layer4_outputs(1927) <= not (a or b);
    layer4_outputs(1928) <= not a or b;
    layer4_outputs(1929) <= not a;
    layer4_outputs(1930) <= not (a or b);
    layer4_outputs(1931) <= a;
    layer4_outputs(1932) <= not (a and b);
    layer4_outputs(1933) <= b;
    layer4_outputs(1934) <= not b;
    layer4_outputs(1935) <= not (a xor b);
    layer4_outputs(1936) <= not a;
    layer4_outputs(1937) <= a and b;
    layer4_outputs(1938) <= a;
    layer4_outputs(1939) <= not a;
    layer4_outputs(1940) <= not a;
    layer4_outputs(1941) <= not a;
    layer4_outputs(1942) <= not b;
    layer4_outputs(1943) <= b and not a;
    layer4_outputs(1944) <= not b or a;
    layer4_outputs(1945) <= not (a or b);
    layer4_outputs(1946) <= not a;
    layer4_outputs(1947) <= not a or b;
    layer4_outputs(1948) <= not a or b;
    layer4_outputs(1949) <= a or b;
    layer4_outputs(1950) <= a and b;
    layer4_outputs(1951) <= not a;
    layer4_outputs(1952) <= not a;
    layer4_outputs(1953) <= a;
    layer4_outputs(1954) <= not a or b;
    layer4_outputs(1955) <= b;
    layer4_outputs(1956) <= a or b;
    layer4_outputs(1957) <= a and not b;
    layer4_outputs(1958) <= not a;
    layer4_outputs(1959) <= not (a or b);
    layer4_outputs(1960) <= b and not a;
    layer4_outputs(1961) <= not (a xor b);
    layer4_outputs(1962) <= not a or b;
    layer4_outputs(1963) <= not a;
    layer4_outputs(1964) <= not (a or b);
    layer4_outputs(1965) <= not a;
    layer4_outputs(1966) <= not (a and b);
    layer4_outputs(1967) <= a;
    layer4_outputs(1968) <= a xor b;
    layer4_outputs(1969) <= a and not b;
    layer4_outputs(1970) <= a and not b;
    layer4_outputs(1971) <= not a;
    layer4_outputs(1972) <= a and b;
    layer4_outputs(1973) <= not (a and b);
    layer4_outputs(1974) <= not (a xor b);
    layer4_outputs(1975) <= not b or a;
    layer4_outputs(1976) <= not b;
    layer4_outputs(1977) <= a;
    layer4_outputs(1978) <= a and b;
    layer4_outputs(1979) <= not b or a;
    layer4_outputs(1980) <= not b;
    layer4_outputs(1981) <= a or b;
    layer4_outputs(1982) <= not a;
    layer4_outputs(1983) <= a xor b;
    layer4_outputs(1984) <= not b;
    layer4_outputs(1985) <= a;
    layer4_outputs(1986) <= not b or a;
    layer4_outputs(1987) <= b;
    layer4_outputs(1988) <= not a or b;
    layer4_outputs(1989) <= a;
    layer4_outputs(1990) <= not b;
    layer4_outputs(1991) <= a;
    layer4_outputs(1992) <= a or b;
    layer4_outputs(1993) <= not a;
    layer4_outputs(1994) <= not b or a;
    layer4_outputs(1995) <= a;
    layer4_outputs(1996) <= not a;
    layer4_outputs(1997) <= not a or b;
    layer4_outputs(1998) <= not b;
    layer4_outputs(1999) <= not a;
    layer4_outputs(2000) <= b;
    layer4_outputs(2001) <= not a;
    layer4_outputs(2002) <= not b;
    layer4_outputs(2003) <= not (a and b);
    layer4_outputs(2004) <= not b;
    layer4_outputs(2005) <= a xor b;
    layer4_outputs(2006) <= not b;
    layer4_outputs(2007) <= not a;
    layer4_outputs(2008) <= a and not b;
    layer4_outputs(2009) <= not a or b;
    layer4_outputs(2010) <= b;
    layer4_outputs(2011) <= a and b;
    layer4_outputs(2012) <= not a;
    layer4_outputs(2013) <= not b or a;
    layer4_outputs(2014) <= not b;
    layer4_outputs(2015) <= a and b;
    layer4_outputs(2016) <= a;
    layer4_outputs(2017) <= not (a xor b);
    layer4_outputs(2018) <= a or b;
    layer4_outputs(2019) <= not a;
    layer4_outputs(2020) <= not b;
    layer4_outputs(2021) <= not a;
    layer4_outputs(2022) <= not (a or b);
    layer4_outputs(2023) <= b;
    layer4_outputs(2024) <= b and not a;
    layer4_outputs(2025) <= a xor b;
    layer4_outputs(2026) <= a xor b;
    layer4_outputs(2027) <= a xor b;
    layer4_outputs(2028) <= not (a or b);
    layer4_outputs(2029) <= not (a or b);
    layer4_outputs(2030) <= a;
    layer4_outputs(2031) <= b and not a;
    layer4_outputs(2032) <= a or b;
    layer4_outputs(2033) <= b and not a;
    layer4_outputs(2034) <= b;
    layer4_outputs(2035) <= not (a and b);
    layer4_outputs(2036) <= not b;
    layer4_outputs(2037) <= not b;
    layer4_outputs(2038) <= b and not a;
    layer4_outputs(2039) <= not a or b;
    layer4_outputs(2040) <= not b or a;
    layer4_outputs(2041) <= not (a and b);
    layer4_outputs(2042) <= b;
    layer4_outputs(2043) <= b;
    layer4_outputs(2044) <= a;
    layer4_outputs(2045) <= not (a xor b);
    layer4_outputs(2046) <= a;
    layer4_outputs(2047) <= not (a xor b);
    layer4_outputs(2048) <= not (a and b);
    layer4_outputs(2049) <= b and not a;
    layer4_outputs(2050) <= not a;
    layer4_outputs(2051) <= a or b;
    layer4_outputs(2052) <= b;
    layer4_outputs(2053) <= a xor b;
    layer4_outputs(2054) <= not (a and b);
    layer4_outputs(2055) <= '0';
    layer4_outputs(2056) <= not a or b;
    layer4_outputs(2057) <= not (a xor b);
    layer4_outputs(2058) <= a and b;
    layer4_outputs(2059) <= not b;
    layer4_outputs(2060) <= a xor b;
    layer4_outputs(2061) <= a and not b;
    layer4_outputs(2062) <= a xor b;
    layer4_outputs(2063) <= a or b;
    layer4_outputs(2064) <= not (a or b);
    layer4_outputs(2065) <= a or b;
    layer4_outputs(2066) <= not a;
    layer4_outputs(2067) <= not b;
    layer4_outputs(2068) <= not a;
    layer4_outputs(2069) <= b;
    layer4_outputs(2070) <= a or b;
    layer4_outputs(2071) <= a xor b;
    layer4_outputs(2072) <= not a;
    layer4_outputs(2073) <= a and b;
    layer4_outputs(2074) <= a and not b;
    layer4_outputs(2075) <= not a;
    layer4_outputs(2076) <= a;
    layer4_outputs(2077) <= a;
    layer4_outputs(2078) <= not (a or b);
    layer4_outputs(2079) <= not b;
    layer4_outputs(2080) <= not b or a;
    layer4_outputs(2081) <= b and not a;
    layer4_outputs(2082) <= not a;
    layer4_outputs(2083) <= not (a and b);
    layer4_outputs(2084) <= not (a or b);
    layer4_outputs(2085) <= not (a or b);
    layer4_outputs(2086) <= not (a and b);
    layer4_outputs(2087) <= not b;
    layer4_outputs(2088) <= not b;
    layer4_outputs(2089) <= not b;
    layer4_outputs(2090) <= b;
    layer4_outputs(2091) <= a xor b;
    layer4_outputs(2092) <= b;
    layer4_outputs(2093) <= a and b;
    layer4_outputs(2094) <= a and b;
    layer4_outputs(2095) <= not a or b;
    layer4_outputs(2096) <= a xor b;
    layer4_outputs(2097) <= not b;
    layer4_outputs(2098) <= b;
    layer4_outputs(2099) <= not b;
    layer4_outputs(2100) <= not b;
    layer4_outputs(2101) <= not b;
    layer4_outputs(2102) <= b and not a;
    layer4_outputs(2103) <= not (a and b);
    layer4_outputs(2104) <= not (a xor b);
    layer4_outputs(2105) <= '1';
    layer4_outputs(2106) <= not b or a;
    layer4_outputs(2107) <= a;
    layer4_outputs(2108) <= not a;
    layer4_outputs(2109) <= not b or a;
    layer4_outputs(2110) <= not b;
    layer4_outputs(2111) <= a xor b;
    layer4_outputs(2112) <= b;
    layer4_outputs(2113) <= a and b;
    layer4_outputs(2114) <= not (a and b);
    layer4_outputs(2115) <= not (a xor b);
    layer4_outputs(2116) <= a xor b;
    layer4_outputs(2117) <= a xor b;
    layer4_outputs(2118) <= a and not b;
    layer4_outputs(2119) <= not b;
    layer4_outputs(2120) <= a or b;
    layer4_outputs(2121) <= a and not b;
    layer4_outputs(2122) <= not a;
    layer4_outputs(2123) <= b;
    layer4_outputs(2124) <= not b;
    layer4_outputs(2125) <= not a;
    layer4_outputs(2126) <= not a or b;
    layer4_outputs(2127) <= b and not a;
    layer4_outputs(2128) <= a;
    layer4_outputs(2129) <= b;
    layer4_outputs(2130) <= a and not b;
    layer4_outputs(2131) <= not a;
    layer4_outputs(2132) <= a xor b;
    layer4_outputs(2133) <= not a or b;
    layer4_outputs(2134) <= a xor b;
    layer4_outputs(2135) <= b;
    layer4_outputs(2136) <= a;
    layer4_outputs(2137) <= a and not b;
    layer4_outputs(2138) <= not a or b;
    layer4_outputs(2139) <= not a or b;
    layer4_outputs(2140) <= not a or b;
    layer4_outputs(2141) <= a;
    layer4_outputs(2142) <= a;
    layer4_outputs(2143) <= b;
    layer4_outputs(2144) <= not (a and b);
    layer4_outputs(2145) <= a;
    layer4_outputs(2146) <= not a or b;
    layer4_outputs(2147) <= not b;
    layer4_outputs(2148) <= b and not a;
    layer4_outputs(2149) <= not b or a;
    layer4_outputs(2150) <= not (a or b);
    layer4_outputs(2151) <= not a or b;
    layer4_outputs(2152) <= not b;
    layer4_outputs(2153) <= a and not b;
    layer4_outputs(2154) <= not b;
    layer4_outputs(2155) <= not (a or b);
    layer4_outputs(2156) <= b and not a;
    layer4_outputs(2157) <= not b;
    layer4_outputs(2158) <= not (a or b);
    layer4_outputs(2159) <= not a;
    layer4_outputs(2160) <= not a;
    layer4_outputs(2161) <= b;
    layer4_outputs(2162) <= not a;
    layer4_outputs(2163) <= not a or b;
    layer4_outputs(2164) <= not a;
    layer4_outputs(2165) <= not a or b;
    layer4_outputs(2166) <= not (a and b);
    layer4_outputs(2167) <= not a or b;
    layer4_outputs(2168) <= a and b;
    layer4_outputs(2169) <= a and not b;
    layer4_outputs(2170) <= a or b;
    layer4_outputs(2171) <= not (a xor b);
    layer4_outputs(2172) <= b;
    layer4_outputs(2173) <= '0';
    layer4_outputs(2174) <= not (a and b);
    layer4_outputs(2175) <= not (a and b);
    layer4_outputs(2176) <= a or b;
    layer4_outputs(2177) <= not a;
    layer4_outputs(2178) <= not b or a;
    layer4_outputs(2179) <= not a or b;
    layer4_outputs(2180) <= a and not b;
    layer4_outputs(2181) <= not b;
    layer4_outputs(2182) <= not (a or b);
    layer4_outputs(2183) <= not a or b;
    layer4_outputs(2184) <= not (a and b);
    layer4_outputs(2185) <= b and not a;
    layer4_outputs(2186) <= not b;
    layer4_outputs(2187) <= a and not b;
    layer4_outputs(2188) <= a and b;
    layer4_outputs(2189) <= b;
    layer4_outputs(2190) <= not (a and b);
    layer4_outputs(2191) <= not (a xor b);
    layer4_outputs(2192) <= a;
    layer4_outputs(2193) <= a and not b;
    layer4_outputs(2194) <= not a or b;
    layer4_outputs(2195) <= not b;
    layer4_outputs(2196) <= a or b;
    layer4_outputs(2197) <= a or b;
    layer4_outputs(2198) <= a or b;
    layer4_outputs(2199) <= a and not b;
    layer4_outputs(2200) <= not a;
    layer4_outputs(2201) <= a and b;
    layer4_outputs(2202) <= b;
    layer4_outputs(2203) <= not b;
    layer4_outputs(2204) <= b;
    layer4_outputs(2205) <= a and not b;
    layer4_outputs(2206) <= '0';
    layer4_outputs(2207) <= a;
    layer4_outputs(2208) <= not (a and b);
    layer4_outputs(2209) <= b;
    layer4_outputs(2210) <= b;
    layer4_outputs(2211) <= not b;
    layer4_outputs(2212) <= a and b;
    layer4_outputs(2213) <= a;
    layer4_outputs(2214) <= not (a and b);
    layer4_outputs(2215) <= not a or b;
    layer4_outputs(2216) <= a;
    layer4_outputs(2217) <= a or b;
    layer4_outputs(2218) <= a or b;
    layer4_outputs(2219) <= not (a or b);
    layer4_outputs(2220) <= not b;
    layer4_outputs(2221) <= a and not b;
    layer4_outputs(2222) <= not a;
    layer4_outputs(2223) <= not (a and b);
    layer4_outputs(2224) <= not (a xor b);
    layer4_outputs(2225) <= b;
    layer4_outputs(2226) <= a xor b;
    layer4_outputs(2227) <= a;
    layer4_outputs(2228) <= not a or b;
    layer4_outputs(2229) <= not (a and b);
    layer4_outputs(2230) <= not a or b;
    layer4_outputs(2231) <= a xor b;
    layer4_outputs(2232) <= not a;
    layer4_outputs(2233) <= not b;
    layer4_outputs(2234) <= a and b;
    layer4_outputs(2235) <= a;
    layer4_outputs(2236) <= not (a xor b);
    layer4_outputs(2237) <= not (a xor b);
    layer4_outputs(2238) <= not (a and b);
    layer4_outputs(2239) <= not (a xor b);
    layer4_outputs(2240) <= a and b;
    layer4_outputs(2241) <= a and b;
    layer4_outputs(2242) <= a;
    layer4_outputs(2243) <= b;
    layer4_outputs(2244) <= not b;
    layer4_outputs(2245) <= a xor b;
    layer4_outputs(2246) <= a;
    layer4_outputs(2247) <= not b;
    layer4_outputs(2248) <= a and b;
    layer4_outputs(2249) <= not (a xor b);
    layer4_outputs(2250) <= b;
    layer4_outputs(2251) <= b;
    layer4_outputs(2252) <= not a;
    layer4_outputs(2253) <= a and b;
    layer4_outputs(2254) <= a xor b;
    layer4_outputs(2255) <= a and b;
    layer4_outputs(2256) <= not (a and b);
    layer4_outputs(2257) <= not (a and b);
    layer4_outputs(2258) <= b and not a;
    layer4_outputs(2259) <= b;
    layer4_outputs(2260) <= not b or a;
    layer4_outputs(2261) <= not b;
    layer4_outputs(2262) <= not b;
    layer4_outputs(2263) <= a;
    layer4_outputs(2264) <= not (a and b);
    layer4_outputs(2265) <= not b;
    layer4_outputs(2266) <= a and b;
    layer4_outputs(2267) <= not (a and b);
    layer4_outputs(2268) <= a and b;
    layer4_outputs(2269) <= not b;
    layer4_outputs(2270) <= not a or b;
    layer4_outputs(2271) <= not (a xor b);
    layer4_outputs(2272) <= '1';
    layer4_outputs(2273) <= not a;
    layer4_outputs(2274) <= a or b;
    layer4_outputs(2275) <= not b;
    layer4_outputs(2276) <= a and not b;
    layer4_outputs(2277) <= not b;
    layer4_outputs(2278) <= not b or a;
    layer4_outputs(2279) <= not b;
    layer4_outputs(2280) <= a or b;
    layer4_outputs(2281) <= not (a or b);
    layer4_outputs(2282) <= a xor b;
    layer4_outputs(2283) <= b;
    layer4_outputs(2284) <= a;
    layer4_outputs(2285) <= a;
    layer4_outputs(2286) <= b;
    layer4_outputs(2287) <= not a;
    layer4_outputs(2288) <= not (a or b);
    layer4_outputs(2289) <= not a;
    layer4_outputs(2290) <= not b;
    layer4_outputs(2291) <= b;
    layer4_outputs(2292) <= a or b;
    layer4_outputs(2293) <= not (a xor b);
    layer4_outputs(2294) <= not a;
    layer4_outputs(2295) <= not (a xor b);
    layer4_outputs(2296) <= not (a or b);
    layer4_outputs(2297) <= a and b;
    layer4_outputs(2298) <= b;
    layer4_outputs(2299) <= a and not b;
    layer4_outputs(2300) <= a or b;
    layer4_outputs(2301) <= not a;
    layer4_outputs(2302) <= a or b;
    layer4_outputs(2303) <= b and not a;
    layer4_outputs(2304) <= not a or b;
    layer4_outputs(2305) <= not b or a;
    layer4_outputs(2306) <= not b;
    layer4_outputs(2307) <= not b;
    layer4_outputs(2308) <= a;
    layer4_outputs(2309) <= not b or a;
    layer4_outputs(2310) <= b and not a;
    layer4_outputs(2311) <= not (a and b);
    layer4_outputs(2312) <= b and not a;
    layer4_outputs(2313) <= a;
    layer4_outputs(2314) <= a;
    layer4_outputs(2315) <= a or b;
    layer4_outputs(2316) <= a;
    layer4_outputs(2317) <= not (a xor b);
    layer4_outputs(2318) <= not a;
    layer4_outputs(2319) <= not b;
    layer4_outputs(2320) <= '1';
    layer4_outputs(2321) <= a;
    layer4_outputs(2322) <= a or b;
    layer4_outputs(2323) <= not b;
    layer4_outputs(2324) <= not (a xor b);
    layer4_outputs(2325) <= not a;
    layer4_outputs(2326) <= b and not a;
    layer4_outputs(2327) <= a;
    layer4_outputs(2328) <= a and not b;
    layer4_outputs(2329) <= not a;
    layer4_outputs(2330) <= not b or a;
    layer4_outputs(2331) <= a and b;
    layer4_outputs(2332) <= a and b;
    layer4_outputs(2333) <= not (a and b);
    layer4_outputs(2334) <= not a;
    layer4_outputs(2335) <= not a;
    layer4_outputs(2336) <= not b or a;
    layer4_outputs(2337) <= b and not a;
    layer4_outputs(2338) <= not a or b;
    layer4_outputs(2339) <= not a or b;
    layer4_outputs(2340) <= a or b;
    layer4_outputs(2341) <= not a or b;
    layer4_outputs(2342) <= not (a xor b);
    layer4_outputs(2343) <= a or b;
    layer4_outputs(2344) <= not (a xor b);
    layer4_outputs(2345) <= a;
    layer4_outputs(2346) <= not b;
    layer4_outputs(2347) <= a xor b;
    layer4_outputs(2348) <= not b;
    layer4_outputs(2349) <= not b;
    layer4_outputs(2350) <= a;
    layer4_outputs(2351) <= a;
    layer4_outputs(2352) <= not a or b;
    layer4_outputs(2353) <= not (a xor b);
    layer4_outputs(2354) <= not b;
    layer4_outputs(2355) <= a and b;
    layer4_outputs(2356) <= not (a xor b);
    layer4_outputs(2357) <= b;
    layer4_outputs(2358) <= b;
    layer4_outputs(2359) <= not (a xor b);
    layer4_outputs(2360) <= not (a xor b);
    layer4_outputs(2361) <= not b or a;
    layer4_outputs(2362) <= not b;
    layer4_outputs(2363) <= a;
    layer4_outputs(2364) <= a;
    layer4_outputs(2365) <= a;
    layer4_outputs(2366) <= not a;
    layer4_outputs(2367) <= not b;
    layer4_outputs(2368) <= b;
    layer4_outputs(2369) <= not b or a;
    layer4_outputs(2370) <= not b or a;
    layer4_outputs(2371) <= not b or a;
    layer4_outputs(2372) <= a;
    layer4_outputs(2373) <= a and not b;
    layer4_outputs(2374) <= b and not a;
    layer4_outputs(2375) <= not a;
    layer4_outputs(2376) <= not a;
    layer4_outputs(2377) <= not (a and b);
    layer4_outputs(2378) <= a and b;
    layer4_outputs(2379) <= not a;
    layer4_outputs(2380) <= a;
    layer4_outputs(2381) <= not a;
    layer4_outputs(2382) <= not a or b;
    layer4_outputs(2383) <= not a;
    layer4_outputs(2384) <= not b or a;
    layer4_outputs(2385) <= b;
    layer4_outputs(2386) <= a;
    layer4_outputs(2387) <= not (a or b);
    layer4_outputs(2388) <= b;
    layer4_outputs(2389) <= not a;
    layer4_outputs(2390) <= b;
    layer4_outputs(2391) <= '0';
    layer4_outputs(2392) <= not (a xor b);
    layer4_outputs(2393) <= b and not a;
    layer4_outputs(2394) <= not b;
    layer4_outputs(2395) <= not (a or b);
    layer4_outputs(2396) <= not a;
    layer4_outputs(2397) <= a and not b;
    layer4_outputs(2398) <= a xor b;
    layer4_outputs(2399) <= a xor b;
    layer4_outputs(2400) <= not b or a;
    layer4_outputs(2401) <= not b;
    layer4_outputs(2402) <= not a;
    layer4_outputs(2403) <= b and not a;
    layer4_outputs(2404) <= a xor b;
    layer4_outputs(2405) <= a and b;
    layer4_outputs(2406) <= not b;
    layer4_outputs(2407) <= b and not a;
    layer4_outputs(2408) <= a;
    layer4_outputs(2409) <= not a;
    layer4_outputs(2410) <= a;
    layer4_outputs(2411) <= not a;
    layer4_outputs(2412) <= not b;
    layer4_outputs(2413) <= not a or b;
    layer4_outputs(2414) <= b and not a;
    layer4_outputs(2415) <= not b;
    layer4_outputs(2416) <= b and not a;
    layer4_outputs(2417) <= b;
    layer4_outputs(2418) <= a and not b;
    layer4_outputs(2419) <= not (a xor b);
    layer4_outputs(2420) <= a and not b;
    layer4_outputs(2421) <= b;
    layer4_outputs(2422) <= b;
    layer4_outputs(2423) <= not a;
    layer4_outputs(2424) <= '1';
    layer4_outputs(2425) <= a;
    layer4_outputs(2426) <= a xor b;
    layer4_outputs(2427) <= not a;
    layer4_outputs(2428) <= not b;
    layer4_outputs(2429) <= not (a xor b);
    layer4_outputs(2430) <= b;
    layer4_outputs(2431) <= b and not a;
    layer4_outputs(2432) <= a or b;
    layer4_outputs(2433) <= not b;
    layer4_outputs(2434) <= not b;
    layer4_outputs(2435) <= b;
    layer4_outputs(2436) <= not (a or b);
    layer4_outputs(2437) <= a and b;
    layer4_outputs(2438) <= not (a xor b);
    layer4_outputs(2439) <= a;
    layer4_outputs(2440) <= not b or a;
    layer4_outputs(2441) <= a and not b;
    layer4_outputs(2442) <= a;
    layer4_outputs(2443) <= not b or a;
    layer4_outputs(2444) <= a;
    layer4_outputs(2445) <= not b;
    layer4_outputs(2446) <= a;
    layer4_outputs(2447) <= not (a xor b);
    layer4_outputs(2448) <= a and not b;
    layer4_outputs(2449) <= b and not a;
    layer4_outputs(2450) <= a;
    layer4_outputs(2451) <= not b;
    layer4_outputs(2452) <= b;
    layer4_outputs(2453) <= b;
    layer4_outputs(2454) <= not b;
    layer4_outputs(2455) <= b and not a;
    layer4_outputs(2456) <= '1';
    layer4_outputs(2457) <= a and b;
    layer4_outputs(2458) <= not a;
    layer4_outputs(2459) <= not (a xor b);
    layer4_outputs(2460) <= not a;
    layer4_outputs(2461) <= b and not a;
    layer4_outputs(2462) <= a and b;
    layer4_outputs(2463) <= not b;
    layer4_outputs(2464) <= a xor b;
    layer4_outputs(2465) <= not b;
    layer4_outputs(2466) <= b;
    layer4_outputs(2467) <= b;
    layer4_outputs(2468) <= not a;
    layer4_outputs(2469) <= not (a and b);
    layer4_outputs(2470) <= not b or a;
    layer4_outputs(2471) <= not b;
    layer4_outputs(2472) <= not b;
    layer4_outputs(2473) <= b;
    layer4_outputs(2474) <= not (a or b);
    layer4_outputs(2475) <= not a;
    layer4_outputs(2476) <= a or b;
    layer4_outputs(2477) <= not (a xor b);
    layer4_outputs(2478) <= a and b;
    layer4_outputs(2479) <= not a or b;
    layer4_outputs(2480) <= a;
    layer4_outputs(2481) <= a and b;
    layer4_outputs(2482) <= not (a or b);
    layer4_outputs(2483) <= not (a and b);
    layer4_outputs(2484) <= a and not b;
    layer4_outputs(2485) <= not b;
    layer4_outputs(2486) <= not a or b;
    layer4_outputs(2487) <= a or b;
    layer4_outputs(2488) <= not a;
    layer4_outputs(2489) <= not (a or b);
    layer4_outputs(2490) <= b;
    layer4_outputs(2491) <= not (a and b);
    layer4_outputs(2492) <= b and not a;
    layer4_outputs(2493) <= not a;
    layer4_outputs(2494) <= a xor b;
    layer4_outputs(2495) <= a or b;
    layer4_outputs(2496) <= a;
    layer4_outputs(2497) <= b;
    layer4_outputs(2498) <= b and not a;
    layer4_outputs(2499) <= b;
    layer4_outputs(2500) <= not b;
    layer4_outputs(2501) <= a xor b;
    layer4_outputs(2502) <= a or b;
    layer4_outputs(2503) <= b;
    layer4_outputs(2504) <= not (a or b);
    layer4_outputs(2505) <= b;
    layer4_outputs(2506) <= a xor b;
    layer4_outputs(2507) <= a or b;
    layer4_outputs(2508) <= b;
    layer4_outputs(2509) <= not a;
    layer4_outputs(2510) <= b and not a;
    layer4_outputs(2511) <= not a or b;
    layer4_outputs(2512) <= a or b;
    layer4_outputs(2513) <= not a;
    layer4_outputs(2514) <= '1';
    layer4_outputs(2515) <= a;
    layer4_outputs(2516) <= a xor b;
    layer4_outputs(2517) <= a and not b;
    layer4_outputs(2518) <= a and b;
    layer4_outputs(2519) <= a;
    layer4_outputs(2520) <= not b;
    layer4_outputs(2521) <= not (a and b);
    layer4_outputs(2522) <= not a;
    layer4_outputs(2523) <= not b;
    layer4_outputs(2524) <= not b or a;
    layer4_outputs(2525) <= a and not b;
    layer4_outputs(2526) <= not b or a;
    layer4_outputs(2527) <= not b or a;
    layer4_outputs(2528) <= a;
    layer4_outputs(2529) <= a or b;
    layer4_outputs(2530) <= b;
    layer4_outputs(2531) <= a and not b;
    layer4_outputs(2532) <= b;
    layer4_outputs(2533) <= a and not b;
    layer4_outputs(2534) <= not b;
    layer4_outputs(2535) <= not a;
    layer4_outputs(2536) <= '1';
    layer4_outputs(2537) <= not (a or b);
    layer4_outputs(2538) <= not a;
    layer4_outputs(2539) <= a and not b;
    layer4_outputs(2540) <= a;
    layer4_outputs(2541) <= not b;
    layer4_outputs(2542) <= a xor b;
    layer4_outputs(2543) <= a;
    layer4_outputs(2544) <= b;
    layer4_outputs(2545) <= not b;
    layer4_outputs(2546) <= a;
    layer4_outputs(2547) <= a;
    layer4_outputs(2548) <= b;
    layer4_outputs(2549) <= a or b;
    layer4_outputs(2550) <= a or b;
    layer4_outputs(2551) <= not b;
    layer4_outputs(2552) <= b;
    layer4_outputs(2553) <= a and b;
    layer4_outputs(2554) <= not b;
    layer4_outputs(2555) <= not b;
    layer4_outputs(2556) <= not (a or b);
    layer4_outputs(2557) <= a and b;
    layer4_outputs(2558) <= not (a xor b);
    layer4_outputs(2559) <= not (a and b);
    layer4_outputs(2560) <= not (a xor b);
    layer4_outputs(2561) <= '0';
    layer4_outputs(2562) <= b;
    layer4_outputs(2563) <= not a or b;
    layer4_outputs(2564) <= a xor b;
    layer4_outputs(2565) <= not a;
    layer4_outputs(2566) <= not b;
    layer4_outputs(2567) <= not b;
    layer4_outputs(2568) <= not (a and b);
    layer4_outputs(2569) <= not a or b;
    layer4_outputs(2570) <= not b or a;
    layer4_outputs(2571) <= not a;
    layer4_outputs(2572) <= b;
    layer4_outputs(2573) <= a and b;
    layer4_outputs(2574) <= not (a and b);
    layer4_outputs(2575) <= not (a and b);
    layer4_outputs(2576) <= not b or a;
    layer4_outputs(2577) <= not a;
    layer4_outputs(2578) <= b;
    layer4_outputs(2579) <= b and not a;
    layer4_outputs(2580) <= not (a xor b);
    layer4_outputs(2581) <= a;
    layer4_outputs(2582) <= not b;
    layer4_outputs(2583) <= a and b;
    layer4_outputs(2584) <= not (a and b);
    layer4_outputs(2585) <= a or b;
    layer4_outputs(2586) <= not (a or b);
    layer4_outputs(2587) <= b;
    layer4_outputs(2588) <= a;
    layer4_outputs(2589) <= not b;
    layer4_outputs(2590) <= not b or a;
    layer4_outputs(2591) <= not (a xor b);
    layer4_outputs(2592) <= b;
    layer4_outputs(2593) <= b;
    layer4_outputs(2594) <= not (a and b);
    layer4_outputs(2595) <= not (a and b);
    layer4_outputs(2596) <= a;
    layer4_outputs(2597) <= not a or b;
    layer4_outputs(2598) <= not b;
    layer4_outputs(2599) <= a;
    layer4_outputs(2600) <= not a or b;
    layer4_outputs(2601) <= b and not a;
    layer4_outputs(2602) <= not (a and b);
    layer4_outputs(2603) <= not (a xor b);
    layer4_outputs(2604) <= not (a xor b);
    layer4_outputs(2605) <= not a or b;
    layer4_outputs(2606) <= not a;
    layer4_outputs(2607) <= b;
    layer4_outputs(2608) <= not b;
    layer4_outputs(2609) <= a xor b;
    layer4_outputs(2610) <= a and not b;
    layer4_outputs(2611) <= a;
    layer4_outputs(2612) <= b;
    layer4_outputs(2613) <= not b;
    layer4_outputs(2614) <= a and not b;
    layer4_outputs(2615) <= not b;
    layer4_outputs(2616) <= not a or b;
    layer4_outputs(2617) <= a xor b;
    layer4_outputs(2618) <= a;
    layer4_outputs(2619) <= not a or b;
    layer4_outputs(2620) <= not (a or b);
    layer4_outputs(2621) <= a or b;
    layer4_outputs(2622) <= a;
    layer4_outputs(2623) <= a;
    layer4_outputs(2624) <= a xor b;
    layer4_outputs(2625) <= a;
    layer4_outputs(2626) <= a;
    layer4_outputs(2627) <= a;
    layer4_outputs(2628) <= not (a or b);
    layer4_outputs(2629) <= a;
    layer4_outputs(2630) <= a;
    layer4_outputs(2631) <= a;
    layer4_outputs(2632) <= not (a xor b);
    layer4_outputs(2633) <= not (a and b);
    layer4_outputs(2634) <= a;
    layer4_outputs(2635) <= not (a or b);
    layer4_outputs(2636) <= not (a or b);
    layer4_outputs(2637) <= not (a and b);
    layer4_outputs(2638) <= not a;
    layer4_outputs(2639) <= a and b;
    layer4_outputs(2640) <= a and not b;
    layer4_outputs(2641) <= b and not a;
    layer4_outputs(2642) <= b and not a;
    layer4_outputs(2643) <= not b;
    layer4_outputs(2644) <= a xor b;
    layer4_outputs(2645) <= a and not b;
    layer4_outputs(2646) <= not (a and b);
    layer4_outputs(2647) <= not a;
    layer4_outputs(2648) <= a xor b;
    layer4_outputs(2649) <= not a;
    layer4_outputs(2650) <= not b;
    layer4_outputs(2651) <= b;
    layer4_outputs(2652) <= a;
    layer4_outputs(2653) <= a;
    layer4_outputs(2654) <= a;
    layer4_outputs(2655) <= not (a and b);
    layer4_outputs(2656) <= not (a and b);
    layer4_outputs(2657) <= not (a and b);
    layer4_outputs(2658) <= not (a xor b);
    layer4_outputs(2659) <= a and b;
    layer4_outputs(2660) <= '0';
    layer4_outputs(2661) <= a xor b;
    layer4_outputs(2662) <= not a;
    layer4_outputs(2663) <= '0';
    layer4_outputs(2664) <= not (a or b);
    layer4_outputs(2665) <= a;
    layer4_outputs(2666) <= not (a and b);
    layer4_outputs(2667) <= not a;
    layer4_outputs(2668) <= b;
    layer4_outputs(2669) <= a and not b;
    layer4_outputs(2670) <= not a;
    layer4_outputs(2671) <= a and b;
    layer4_outputs(2672) <= a and not b;
    layer4_outputs(2673) <= a;
    layer4_outputs(2674) <= not (a and b);
    layer4_outputs(2675) <= not (a xor b);
    layer4_outputs(2676) <= b and not a;
    layer4_outputs(2677) <= not a;
    layer4_outputs(2678) <= b;
    layer4_outputs(2679) <= a xor b;
    layer4_outputs(2680) <= not (a xor b);
    layer4_outputs(2681) <= not b;
    layer4_outputs(2682) <= not b;
    layer4_outputs(2683) <= a and not b;
    layer4_outputs(2684) <= a xor b;
    layer4_outputs(2685) <= not a;
    layer4_outputs(2686) <= b and not a;
    layer4_outputs(2687) <= not a;
    layer4_outputs(2688) <= not a;
    layer4_outputs(2689) <= not a;
    layer4_outputs(2690) <= a xor b;
    layer4_outputs(2691) <= not (a or b);
    layer4_outputs(2692) <= b and not a;
    layer4_outputs(2693) <= a and not b;
    layer4_outputs(2694) <= b;
    layer4_outputs(2695) <= not b;
    layer4_outputs(2696) <= not a;
    layer4_outputs(2697) <= not b;
    layer4_outputs(2698) <= a or b;
    layer4_outputs(2699) <= b;
    layer4_outputs(2700) <= not a;
    layer4_outputs(2701) <= not (a and b);
    layer4_outputs(2702) <= a xor b;
    layer4_outputs(2703) <= not (a or b);
    layer4_outputs(2704) <= a or b;
    layer4_outputs(2705) <= not a;
    layer4_outputs(2706) <= b and not a;
    layer4_outputs(2707) <= b and not a;
    layer4_outputs(2708) <= not (a or b);
    layer4_outputs(2709) <= not b;
    layer4_outputs(2710) <= b;
    layer4_outputs(2711) <= not (a and b);
    layer4_outputs(2712) <= not a;
    layer4_outputs(2713) <= b;
    layer4_outputs(2714) <= a and b;
    layer4_outputs(2715) <= a;
    layer4_outputs(2716) <= not (a or b);
    layer4_outputs(2717) <= a and not b;
    layer4_outputs(2718) <= a;
    layer4_outputs(2719) <= not a;
    layer4_outputs(2720) <= not b;
    layer4_outputs(2721) <= b;
    layer4_outputs(2722) <= a;
    layer4_outputs(2723) <= not a or b;
    layer4_outputs(2724) <= not a;
    layer4_outputs(2725) <= not b;
    layer4_outputs(2726) <= not a;
    layer4_outputs(2727) <= a;
    layer4_outputs(2728) <= not a;
    layer4_outputs(2729) <= a and not b;
    layer4_outputs(2730) <= a;
    layer4_outputs(2731) <= a and b;
    layer4_outputs(2732) <= b;
    layer4_outputs(2733) <= not (a or b);
    layer4_outputs(2734) <= a and not b;
    layer4_outputs(2735) <= not a;
    layer4_outputs(2736) <= b and not a;
    layer4_outputs(2737) <= a xor b;
    layer4_outputs(2738) <= not a or b;
    layer4_outputs(2739) <= not (a or b);
    layer4_outputs(2740) <= not (a xor b);
    layer4_outputs(2741) <= b;
    layer4_outputs(2742) <= not b;
    layer4_outputs(2743) <= a;
    layer4_outputs(2744) <= a and b;
    layer4_outputs(2745) <= not a;
    layer4_outputs(2746) <= not b;
    layer4_outputs(2747) <= a and not b;
    layer4_outputs(2748) <= not (a and b);
    layer4_outputs(2749) <= a and b;
    layer4_outputs(2750) <= not b;
    layer4_outputs(2751) <= a and not b;
    layer4_outputs(2752) <= b;
    layer4_outputs(2753) <= '1';
    layer4_outputs(2754) <= not b;
    layer4_outputs(2755) <= a or b;
    layer4_outputs(2756) <= not (a and b);
    layer4_outputs(2757) <= not (a or b);
    layer4_outputs(2758) <= a;
    layer4_outputs(2759) <= a and b;
    layer4_outputs(2760) <= not b;
    layer4_outputs(2761) <= a and not b;
    layer4_outputs(2762) <= not (a and b);
    layer4_outputs(2763) <= a;
    layer4_outputs(2764) <= b and not a;
    layer4_outputs(2765) <= b;
    layer4_outputs(2766) <= a xor b;
    layer4_outputs(2767) <= not a or b;
    layer4_outputs(2768) <= a or b;
    layer4_outputs(2769) <= not (a xor b);
    layer4_outputs(2770) <= not (a and b);
    layer4_outputs(2771) <= a and b;
    layer4_outputs(2772) <= not b or a;
    layer4_outputs(2773) <= b;
    layer4_outputs(2774) <= not a or b;
    layer4_outputs(2775) <= a;
    layer4_outputs(2776) <= not (a xor b);
    layer4_outputs(2777) <= b and not a;
    layer4_outputs(2778) <= not (a and b);
    layer4_outputs(2779) <= a xor b;
    layer4_outputs(2780) <= b;
    layer4_outputs(2781) <= a;
    layer4_outputs(2782) <= b;
    layer4_outputs(2783) <= not b or a;
    layer4_outputs(2784) <= not (a or b);
    layer4_outputs(2785) <= a and b;
    layer4_outputs(2786) <= not b or a;
    layer4_outputs(2787) <= not (a and b);
    layer4_outputs(2788) <= not a;
    layer4_outputs(2789) <= not b;
    layer4_outputs(2790) <= a or b;
    layer4_outputs(2791) <= not a;
    layer4_outputs(2792) <= b and not a;
    layer4_outputs(2793) <= not b;
    layer4_outputs(2794) <= a and not b;
    layer4_outputs(2795) <= not a;
    layer4_outputs(2796) <= a and b;
    layer4_outputs(2797) <= b;
    layer4_outputs(2798) <= a and b;
    layer4_outputs(2799) <= not a;
    layer4_outputs(2800) <= a;
    layer4_outputs(2801) <= not (a xor b);
    layer4_outputs(2802) <= not b;
    layer4_outputs(2803) <= a xor b;
    layer4_outputs(2804) <= not a;
    layer4_outputs(2805) <= not b;
    layer4_outputs(2806) <= not (a xor b);
    layer4_outputs(2807) <= a;
    layer4_outputs(2808) <= a xor b;
    layer4_outputs(2809) <= not b;
    layer4_outputs(2810) <= not b or a;
    layer4_outputs(2811) <= not (a xor b);
    layer4_outputs(2812) <= a or b;
    layer4_outputs(2813) <= not b;
    layer4_outputs(2814) <= not a;
    layer4_outputs(2815) <= b;
    layer4_outputs(2816) <= a;
    layer4_outputs(2817) <= a and not b;
    layer4_outputs(2818) <= not a or b;
    layer4_outputs(2819) <= not b;
    layer4_outputs(2820) <= b;
    layer4_outputs(2821) <= b;
    layer4_outputs(2822) <= a and not b;
    layer4_outputs(2823) <= not b;
    layer4_outputs(2824) <= not (a and b);
    layer4_outputs(2825) <= not (a or b);
    layer4_outputs(2826) <= a or b;
    layer4_outputs(2827) <= not (a xor b);
    layer4_outputs(2828) <= not b;
    layer4_outputs(2829) <= not a;
    layer4_outputs(2830) <= not (a xor b);
    layer4_outputs(2831) <= not b;
    layer4_outputs(2832) <= a and not b;
    layer4_outputs(2833) <= not (a or b);
    layer4_outputs(2834) <= not (a xor b);
    layer4_outputs(2835) <= b;
    layer4_outputs(2836) <= a;
    layer4_outputs(2837) <= a;
    layer4_outputs(2838) <= not b;
    layer4_outputs(2839) <= b and not a;
    layer4_outputs(2840) <= a;
    layer4_outputs(2841) <= a;
    layer4_outputs(2842) <= not a;
    layer4_outputs(2843) <= b and not a;
    layer4_outputs(2844) <= not (a xor b);
    layer4_outputs(2845) <= a or b;
    layer4_outputs(2846) <= not b;
    layer4_outputs(2847) <= not a or b;
    layer4_outputs(2848) <= b and not a;
    layer4_outputs(2849) <= b and not a;
    layer4_outputs(2850) <= a and b;
    layer4_outputs(2851) <= a;
    layer4_outputs(2852) <= a;
    layer4_outputs(2853) <= b and not a;
    layer4_outputs(2854) <= a or b;
    layer4_outputs(2855) <= not b;
    layer4_outputs(2856) <= a and b;
    layer4_outputs(2857) <= not (a and b);
    layer4_outputs(2858) <= not a or b;
    layer4_outputs(2859) <= b;
    layer4_outputs(2860) <= a xor b;
    layer4_outputs(2861) <= not (a or b);
    layer4_outputs(2862) <= b;
    layer4_outputs(2863) <= b;
    layer4_outputs(2864) <= not (a xor b);
    layer4_outputs(2865) <= not (a or b);
    layer4_outputs(2866) <= a;
    layer4_outputs(2867) <= not b;
    layer4_outputs(2868) <= not a or b;
    layer4_outputs(2869) <= a;
    layer4_outputs(2870) <= not b;
    layer4_outputs(2871) <= not (a xor b);
    layer4_outputs(2872) <= not b;
    layer4_outputs(2873) <= a and b;
    layer4_outputs(2874) <= a;
    layer4_outputs(2875) <= b;
    layer4_outputs(2876) <= not (a or b);
    layer4_outputs(2877) <= not b or a;
    layer4_outputs(2878) <= '1';
    layer4_outputs(2879) <= a and b;
    layer4_outputs(2880) <= not b;
    layer4_outputs(2881) <= a;
    layer4_outputs(2882) <= a or b;
    layer4_outputs(2883) <= b;
    layer4_outputs(2884) <= a or b;
    layer4_outputs(2885) <= not a;
    layer4_outputs(2886) <= not b;
    layer4_outputs(2887) <= not a;
    layer4_outputs(2888) <= not a;
    layer4_outputs(2889) <= not (a and b);
    layer4_outputs(2890) <= b and not a;
    layer4_outputs(2891) <= a;
    layer4_outputs(2892) <= a xor b;
    layer4_outputs(2893) <= not (a and b);
    layer4_outputs(2894) <= not (a or b);
    layer4_outputs(2895) <= b and not a;
    layer4_outputs(2896) <= a;
    layer4_outputs(2897) <= b;
    layer4_outputs(2898) <= a;
    layer4_outputs(2899) <= not (a or b);
    layer4_outputs(2900) <= not (a and b);
    layer4_outputs(2901) <= not (a or b);
    layer4_outputs(2902) <= not (a or b);
    layer4_outputs(2903) <= not a or b;
    layer4_outputs(2904) <= b;
    layer4_outputs(2905) <= not a or b;
    layer4_outputs(2906) <= a and not b;
    layer4_outputs(2907) <= not (a or b);
    layer4_outputs(2908) <= a;
    layer4_outputs(2909) <= a;
    layer4_outputs(2910) <= a and b;
    layer4_outputs(2911) <= a or b;
    layer4_outputs(2912) <= not a or b;
    layer4_outputs(2913) <= '1';
    layer4_outputs(2914) <= b;
    layer4_outputs(2915) <= b;
    layer4_outputs(2916) <= b;
    layer4_outputs(2917) <= b and not a;
    layer4_outputs(2918) <= not (a or b);
    layer4_outputs(2919) <= not b;
    layer4_outputs(2920) <= a and b;
    layer4_outputs(2921) <= not (a xor b);
    layer4_outputs(2922) <= not a;
    layer4_outputs(2923) <= a;
    layer4_outputs(2924) <= a;
    layer4_outputs(2925) <= not (a xor b);
    layer4_outputs(2926) <= b;
    layer4_outputs(2927) <= not b;
    layer4_outputs(2928) <= b and not a;
    layer4_outputs(2929) <= a;
    layer4_outputs(2930) <= not a or b;
    layer4_outputs(2931) <= not b;
    layer4_outputs(2932) <= not b;
    layer4_outputs(2933) <= b and not a;
    layer4_outputs(2934) <= not (a xor b);
    layer4_outputs(2935) <= not (a xor b);
    layer4_outputs(2936) <= a;
    layer4_outputs(2937) <= not a;
    layer4_outputs(2938) <= not b;
    layer4_outputs(2939) <= not a or b;
    layer4_outputs(2940) <= b;
    layer4_outputs(2941) <= not a;
    layer4_outputs(2942) <= a and b;
    layer4_outputs(2943) <= not (a xor b);
    layer4_outputs(2944) <= b;
    layer4_outputs(2945) <= not b or a;
    layer4_outputs(2946) <= not a;
    layer4_outputs(2947) <= not (a and b);
    layer4_outputs(2948) <= not a;
    layer4_outputs(2949) <= a and b;
    layer4_outputs(2950) <= b and not a;
    layer4_outputs(2951) <= not (a or b);
    layer4_outputs(2952) <= not (a and b);
    layer4_outputs(2953) <= b;
    layer4_outputs(2954) <= a;
    layer4_outputs(2955) <= a;
    layer4_outputs(2956) <= not (a and b);
    layer4_outputs(2957) <= not (a or b);
    layer4_outputs(2958) <= b and not a;
    layer4_outputs(2959) <= not b or a;
    layer4_outputs(2960) <= not b;
    layer4_outputs(2961) <= not b or a;
    layer4_outputs(2962) <= not a;
    layer4_outputs(2963) <= a;
    layer4_outputs(2964) <= not a;
    layer4_outputs(2965) <= not b;
    layer4_outputs(2966) <= a;
    layer4_outputs(2967) <= not (a and b);
    layer4_outputs(2968) <= a and not b;
    layer4_outputs(2969) <= b;
    layer4_outputs(2970) <= b;
    layer4_outputs(2971) <= not (a xor b);
    layer4_outputs(2972) <= b;
    layer4_outputs(2973) <= a and b;
    layer4_outputs(2974) <= b and not a;
    layer4_outputs(2975) <= b;
    layer4_outputs(2976) <= not (a xor b);
    layer4_outputs(2977) <= a;
    layer4_outputs(2978) <= a or b;
    layer4_outputs(2979) <= not (a and b);
    layer4_outputs(2980) <= not a;
    layer4_outputs(2981) <= not (a xor b);
    layer4_outputs(2982) <= not a;
    layer4_outputs(2983) <= not (a and b);
    layer4_outputs(2984) <= a xor b;
    layer4_outputs(2985) <= a and b;
    layer4_outputs(2986) <= not (a xor b);
    layer4_outputs(2987) <= a xor b;
    layer4_outputs(2988) <= not a;
    layer4_outputs(2989) <= '0';
    layer4_outputs(2990) <= not (a and b);
    layer4_outputs(2991) <= not b;
    layer4_outputs(2992) <= a and b;
    layer4_outputs(2993) <= not (a and b);
    layer4_outputs(2994) <= not (a and b);
    layer4_outputs(2995) <= not b or a;
    layer4_outputs(2996) <= not a;
    layer4_outputs(2997) <= b;
    layer4_outputs(2998) <= not (a and b);
    layer4_outputs(2999) <= not (a and b);
    layer4_outputs(3000) <= not a or b;
    layer4_outputs(3001) <= a xor b;
    layer4_outputs(3002) <= not (a and b);
    layer4_outputs(3003) <= not (a xor b);
    layer4_outputs(3004) <= not (a xor b);
    layer4_outputs(3005) <= a or b;
    layer4_outputs(3006) <= a and b;
    layer4_outputs(3007) <= not b or a;
    layer4_outputs(3008) <= b;
    layer4_outputs(3009) <= a;
    layer4_outputs(3010) <= not b;
    layer4_outputs(3011) <= a xor b;
    layer4_outputs(3012) <= not b;
    layer4_outputs(3013) <= b;
    layer4_outputs(3014) <= not a;
    layer4_outputs(3015) <= a;
    layer4_outputs(3016) <= b;
    layer4_outputs(3017) <= not a or b;
    layer4_outputs(3018) <= not a;
    layer4_outputs(3019) <= not a;
    layer4_outputs(3020) <= b;
    layer4_outputs(3021) <= not (a xor b);
    layer4_outputs(3022) <= a xor b;
    layer4_outputs(3023) <= not a;
    layer4_outputs(3024) <= not a or b;
    layer4_outputs(3025) <= a;
    layer4_outputs(3026) <= not (a xor b);
    layer4_outputs(3027) <= a;
    layer4_outputs(3028) <= not a or b;
    layer4_outputs(3029) <= not a or b;
    layer4_outputs(3030) <= a;
    layer4_outputs(3031) <= not b or a;
    layer4_outputs(3032) <= a or b;
    layer4_outputs(3033) <= not (a xor b);
    layer4_outputs(3034) <= not (a xor b);
    layer4_outputs(3035) <= b;
    layer4_outputs(3036) <= a and b;
    layer4_outputs(3037) <= not a;
    layer4_outputs(3038) <= not a;
    layer4_outputs(3039) <= not b;
    layer4_outputs(3040) <= not a or b;
    layer4_outputs(3041) <= not b;
    layer4_outputs(3042) <= a or b;
    layer4_outputs(3043) <= b and not a;
    layer4_outputs(3044) <= not b or a;
    layer4_outputs(3045) <= a;
    layer4_outputs(3046) <= b and not a;
    layer4_outputs(3047) <= b;
    layer4_outputs(3048) <= not (a xor b);
    layer4_outputs(3049) <= not a;
    layer4_outputs(3050) <= a and b;
    layer4_outputs(3051) <= b and not a;
    layer4_outputs(3052) <= not b;
    layer4_outputs(3053) <= not (a xor b);
    layer4_outputs(3054) <= not a;
    layer4_outputs(3055) <= b;
    layer4_outputs(3056) <= a;
    layer4_outputs(3057) <= not a;
    layer4_outputs(3058) <= a xor b;
    layer4_outputs(3059) <= not b;
    layer4_outputs(3060) <= a and b;
    layer4_outputs(3061) <= not a;
    layer4_outputs(3062) <= a xor b;
    layer4_outputs(3063) <= b and not a;
    layer4_outputs(3064) <= not a;
    layer4_outputs(3065) <= not a;
    layer4_outputs(3066) <= a;
    layer4_outputs(3067) <= a and not b;
    layer4_outputs(3068) <= not a;
    layer4_outputs(3069) <= not (a xor b);
    layer4_outputs(3070) <= not a;
    layer4_outputs(3071) <= a and not b;
    layer4_outputs(3072) <= not b;
    layer4_outputs(3073) <= a and b;
    layer4_outputs(3074) <= not (a or b);
    layer4_outputs(3075) <= not (a xor b);
    layer4_outputs(3076) <= not b;
    layer4_outputs(3077) <= a;
    layer4_outputs(3078) <= not b;
    layer4_outputs(3079) <= '0';
    layer4_outputs(3080) <= a;
    layer4_outputs(3081) <= a or b;
    layer4_outputs(3082) <= not a or b;
    layer4_outputs(3083) <= a;
    layer4_outputs(3084) <= not (a and b);
    layer4_outputs(3085) <= a and not b;
    layer4_outputs(3086) <= a xor b;
    layer4_outputs(3087) <= a or b;
    layer4_outputs(3088) <= a;
    layer4_outputs(3089) <= not a;
    layer4_outputs(3090) <= b;
    layer4_outputs(3091) <= a and b;
    layer4_outputs(3092) <= not b;
    layer4_outputs(3093) <= b;
    layer4_outputs(3094) <= a and not b;
    layer4_outputs(3095) <= a and b;
    layer4_outputs(3096) <= b and not a;
    layer4_outputs(3097) <= not a;
    layer4_outputs(3098) <= not a;
    layer4_outputs(3099) <= b;
    layer4_outputs(3100) <= a and not b;
    layer4_outputs(3101) <= a xor b;
    layer4_outputs(3102) <= not (a or b);
    layer4_outputs(3103) <= not (a and b);
    layer4_outputs(3104) <= not b or a;
    layer4_outputs(3105) <= a or b;
    layer4_outputs(3106) <= not (a or b);
    layer4_outputs(3107) <= not (a or b);
    layer4_outputs(3108) <= a and b;
    layer4_outputs(3109) <= not b;
    layer4_outputs(3110) <= a and b;
    layer4_outputs(3111) <= b;
    layer4_outputs(3112) <= b;
    layer4_outputs(3113) <= '0';
    layer4_outputs(3114) <= not a or b;
    layer4_outputs(3115) <= a xor b;
    layer4_outputs(3116) <= a;
    layer4_outputs(3117) <= not b;
    layer4_outputs(3118) <= not b;
    layer4_outputs(3119) <= b;
    layer4_outputs(3120) <= not b;
    layer4_outputs(3121) <= not a;
    layer4_outputs(3122) <= b;
    layer4_outputs(3123) <= not b;
    layer4_outputs(3124) <= not b;
    layer4_outputs(3125) <= not (a xor b);
    layer4_outputs(3126) <= a;
    layer4_outputs(3127) <= a and b;
    layer4_outputs(3128) <= a and not b;
    layer4_outputs(3129) <= not (a xor b);
    layer4_outputs(3130) <= b;
    layer4_outputs(3131) <= a xor b;
    layer4_outputs(3132) <= not a;
    layer4_outputs(3133) <= not (a and b);
    layer4_outputs(3134) <= not a;
    layer4_outputs(3135) <= not a or b;
    layer4_outputs(3136) <= not b;
    layer4_outputs(3137) <= not a or b;
    layer4_outputs(3138) <= a;
    layer4_outputs(3139) <= a and not b;
    layer4_outputs(3140) <= not b or a;
    layer4_outputs(3141) <= '0';
    layer4_outputs(3142) <= a and b;
    layer4_outputs(3143) <= not b;
    layer4_outputs(3144) <= not b or a;
    layer4_outputs(3145) <= not (a xor b);
    layer4_outputs(3146) <= not (a and b);
    layer4_outputs(3147) <= not b;
    layer4_outputs(3148) <= a;
    layer4_outputs(3149) <= not a or b;
    layer4_outputs(3150) <= a;
    layer4_outputs(3151) <= a;
    layer4_outputs(3152) <= not a;
    layer4_outputs(3153) <= not a;
    layer4_outputs(3154) <= not a;
    layer4_outputs(3155) <= not b;
    layer4_outputs(3156) <= not a;
    layer4_outputs(3157) <= not a;
    layer4_outputs(3158) <= not b or a;
    layer4_outputs(3159) <= a and b;
    layer4_outputs(3160) <= not b;
    layer4_outputs(3161) <= b and not a;
    layer4_outputs(3162) <= a xor b;
    layer4_outputs(3163) <= a;
    layer4_outputs(3164) <= a or b;
    layer4_outputs(3165) <= not a;
    layer4_outputs(3166) <= a xor b;
    layer4_outputs(3167) <= a;
    layer4_outputs(3168) <= a and b;
    layer4_outputs(3169) <= a and b;
    layer4_outputs(3170) <= not (a and b);
    layer4_outputs(3171) <= b;
    layer4_outputs(3172) <= not b;
    layer4_outputs(3173) <= not (a xor b);
    layer4_outputs(3174) <= not b or a;
    layer4_outputs(3175) <= a and b;
    layer4_outputs(3176) <= not a;
    layer4_outputs(3177) <= not (a and b);
    layer4_outputs(3178) <= a and b;
    layer4_outputs(3179) <= a;
    layer4_outputs(3180) <= b;
    layer4_outputs(3181) <= not a or b;
    layer4_outputs(3182) <= not b;
    layer4_outputs(3183) <= a and b;
    layer4_outputs(3184) <= b;
    layer4_outputs(3185) <= not (a and b);
    layer4_outputs(3186) <= not b;
    layer4_outputs(3187) <= a xor b;
    layer4_outputs(3188) <= a or b;
    layer4_outputs(3189) <= not b or a;
    layer4_outputs(3190) <= a or b;
    layer4_outputs(3191) <= a;
    layer4_outputs(3192) <= a xor b;
    layer4_outputs(3193) <= b and not a;
    layer4_outputs(3194) <= a;
    layer4_outputs(3195) <= not (a xor b);
    layer4_outputs(3196) <= not (a xor b);
    layer4_outputs(3197) <= a and b;
    layer4_outputs(3198) <= b and not a;
    layer4_outputs(3199) <= a and not b;
    layer4_outputs(3200) <= a xor b;
    layer4_outputs(3201) <= b and not a;
    layer4_outputs(3202) <= b;
    layer4_outputs(3203) <= not (a xor b);
    layer4_outputs(3204) <= not b;
    layer4_outputs(3205) <= not (a or b);
    layer4_outputs(3206) <= a xor b;
    layer4_outputs(3207) <= not a;
    layer4_outputs(3208) <= a;
    layer4_outputs(3209) <= b;
    layer4_outputs(3210) <= not (a and b);
    layer4_outputs(3211) <= a;
    layer4_outputs(3212) <= not a;
    layer4_outputs(3213) <= a xor b;
    layer4_outputs(3214) <= not a or b;
    layer4_outputs(3215) <= b and not a;
    layer4_outputs(3216) <= not b;
    layer4_outputs(3217) <= not a;
    layer4_outputs(3218) <= not b;
    layer4_outputs(3219) <= a and not b;
    layer4_outputs(3220) <= a or b;
    layer4_outputs(3221) <= a;
    layer4_outputs(3222) <= not (a or b);
    layer4_outputs(3223) <= b;
    layer4_outputs(3224) <= not b;
    layer4_outputs(3225) <= a and not b;
    layer4_outputs(3226) <= a and not b;
    layer4_outputs(3227) <= not b;
    layer4_outputs(3228) <= not b;
    layer4_outputs(3229) <= not (a xor b);
    layer4_outputs(3230) <= b;
    layer4_outputs(3231) <= not a or b;
    layer4_outputs(3232) <= not b;
    layer4_outputs(3233) <= not a;
    layer4_outputs(3234) <= not b or a;
    layer4_outputs(3235) <= a;
    layer4_outputs(3236) <= not a;
    layer4_outputs(3237) <= not (a and b);
    layer4_outputs(3238) <= a;
    layer4_outputs(3239) <= not b;
    layer4_outputs(3240) <= a;
    layer4_outputs(3241) <= not b;
    layer4_outputs(3242) <= a;
    layer4_outputs(3243) <= a;
    layer4_outputs(3244) <= b and not a;
    layer4_outputs(3245) <= not a;
    layer4_outputs(3246) <= a;
    layer4_outputs(3247) <= a and b;
    layer4_outputs(3248) <= a or b;
    layer4_outputs(3249) <= not (a xor b);
    layer4_outputs(3250) <= not (a xor b);
    layer4_outputs(3251) <= a and b;
    layer4_outputs(3252) <= a;
    layer4_outputs(3253) <= a;
    layer4_outputs(3254) <= b and not a;
    layer4_outputs(3255) <= not a;
    layer4_outputs(3256) <= not (a or b);
    layer4_outputs(3257) <= b;
    layer4_outputs(3258) <= not (a xor b);
    layer4_outputs(3259) <= not (a xor b);
    layer4_outputs(3260) <= a or b;
    layer4_outputs(3261) <= a xor b;
    layer4_outputs(3262) <= a;
    layer4_outputs(3263) <= not b;
    layer4_outputs(3264) <= not b;
    layer4_outputs(3265) <= b and not a;
    layer4_outputs(3266) <= not (a xor b);
    layer4_outputs(3267) <= not (a xor b);
    layer4_outputs(3268) <= not (a xor b);
    layer4_outputs(3269) <= not a;
    layer4_outputs(3270) <= a and b;
    layer4_outputs(3271) <= a and b;
    layer4_outputs(3272) <= a and not b;
    layer4_outputs(3273) <= not b or a;
    layer4_outputs(3274) <= not (a xor b);
    layer4_outputs(3275) <= not a;
    layer4_outputs(3276) <= not b;
    layer4_outputs(3277) <= not (a and b);
    layer4_outputs(3278) <= not a;
    layer4_outputs(3279) <= not (a or b);
    layer4_outputs(3280) <= not (a and b);
    layer4_outputs(3281) <= a or b;
    layer4_outputs(3282) <= b;
    layer4_outputs(3283) <= not b;
    layer4_outputs(3284) <= a xor b;
    layer4_outputs(3285) <= a xor b;
    layer4_outputs(3286) <= not (a and b);
    layer4_outputs(3287) <= not (a or b);
    layer4_outputs(3288) <= a;
    layer4_outputs(3289) <= not (a or b);
    layer4_outputs(3290) <= a or b;
    layer4_outputs(3291) <= a xor b;
    layer4_outputs(3292) <= a;
    layer4_outputs(3293) <= not b or a;
    layer4_outputs(3294) <= not a or b;
    layer4_outputs(3295) <= not b or a;
    layer4_outputs(3296) <= a;
    layer4_outputs(3297) <= not b or a;
    layer4_outputs(3298) <= not a or b;
    layer4_outputs(3299) <= a;
    layer4_outputs(3300) <= a xor b;
    layer4_outputs(3301) <= a and b;
    layer4_outputs(3302) <= not b;
    layer4_outputs(3303) <= not a or b;
    layer4_outputs(3304) <= a and not b;
    layer4_outputs(3305) <= not (a and b);
    layer4_outputs(3306) <= not (a and b);
    layer4_outputs(3307) <= a and b;
    layer4_outputs(3308) <= not (a and b);
    layer4_outputs(3309) <= a;
    layer4_outputs(3310) <= '0';
    layer4_outputs(3311) <= b and not a;
    layer4_outputs(3312) <= not (a and b);
    layer4_outputs(3313) <= a xor b;
    layer4_outputs(3314) <= a or b;
    layer4_outputs(3315) <= not a;
    layer4_outputs(3316) <= not a;
    layer4_outputs(3317) <= not a or b;
    layer4_outputs(3318) <= not (a or b);
    layer4_outputs(3319) <= not a or b;
    layer4_outputs(3320) <= not b or a;
    layer4_outputs(3321) <= b;
    layer4_outputs(3322) <= a and not b;
    layer4_outputs(3323) <= not (a or b);
    layer4_outputs(3324) <= b;
    layer4_outputs(3325) <= a xor b;
    layer4_outputs(3326) <= not (a or b);
    layer4_outputs(3327) <= not a;
    layer4_outputs(3328) <= b;
    layer4_outputs(3329) <= a;
    layer4_outputs(3330) <= b;
    layer4_outputs(3331) <= b;
    layer4_outputs(3332) <= a;
    layer4_outputs(3333) <= not (a xor b);
    layer4_outputs(3334) <= not b;
    layer4_outputs(3335) <= a or b;
    layer4_outputs(3336) <= not b or a;
    layer4_outputs(3337) <= b;
    layer4_outputs(3338) <= b;
    layer4_outputs(3339) <= not b;
    layer4_outputs(3340) <= not a or b;
    layer4_outputs(3341) <= not b or a;
    layer4_outputs(3342) <= b;
    layer4_outputs(3343) <= a;
    layer4_outputs(3344) <= a xor b;
    layer4_outputs(3345) <= not a or b;
    layer4_outputs(3346) <= not a;
    layer4_outputs(3347) <= not (a and b);
    layer4_outputs(3348) <= b and not a;
    layer4_outputs(3349) <= a or b;
    layer4_outputs(3350) <= not a;
    layer4_outputs(3351) <= a or b;
    layer4_outputs(3352) <= a and not b;
    layer4_outputs(3353) <= not a;
    layer4_outputs(3354) <= not a or b;
    layer4_outputs(3355) <= not b or a;
    layer4_outputs(3356) <= not b;
    layer4_outputs(3357) <= not b;
    layer4_outputs(3358) <= a and b;
    layer4_outputs(3359) <= a;
    layer4_outputs(3360) <= not (a or b);
    layer4_outputs(3361) <= not b;
    layer4_outputs(3362) <= a;
    layer4_outputs(3363) <= b;
    layer4_outputs(3364) <= b;
    layer4_outputs(3365) <= b;
    layer4_outputs(3366) <= not b;
    layer4_outputs(3367) <= b and not a;
    layer4_outputs(3368) <= b and not a;
    layer4_outputs(3369) <= not a or b;
    layer4_outputs(3370) <= not (a and b);
    layer4_outputs(3371) <= a;
    layer4_outputs(3372) <= not a or b;
    layer4_outputs(3373) <= a and not b;
    layer4_outputs(3374) <= a xor b;
    layer4_outputs(3375) <= not (a and b);
    layer4_outputs(3376) <= b;
    layer4_outputs(3377) <= not b;
    layer4_outputs(3378) <= not b;
    layer4_outputs(3379) <= a xor b;
    layer4_outputs(3380) <= b;
    layer4_outputs(3381) <= b;
    layer4_outputs(3382) <= not (a and b);
    layer4_outputs(3383) <= a xor b;
    layer4_outputs(3384) <= not (a xor b);
    layer4_outputs(3385) <= a;
    layer4_outputs(3386) <= not a;
    layer4_outputs(3387) <= not b;
    layer4_outputs(3388) <= b;
    layer4_outputs(3389) <= not a;
    layer4_outputs(3390) <= not a or b;
    layer4_outputs(3391) <= b;
    layer4_outputs(3392) <= not (a or b);
    layer4_outputs(3393) <= not b or a;
    layer4_outputs(3394) <= not a;
    layer4_outputs(3395) <= not a;
    layer4_outputs(3396) <= not a or b;
    layer4_outputs(3397) <= a xor b;
    layer4_outputs(3398) <= a and not b;
    layer4_outputs(3399) <= b;
    layer4_outputs(3400) <= a or b;
    layer4_outputs(3401) <= a;
    layer4_outputs(3402) <= a and b;
    layer4_outputs(3403) <= b;
    layer4_outputs(3404) <= not a;
    layer4_outputs(3405) <= not b or a;
    layer4_outputs(3406) <= not (a xor b);
    layer4_outputs(3407) <= a xor b;
    layer4_outputs(3408) <= not b;
    layer4_outputs(3409) <= a and b;
    layer4_outputs(3410) <= not b or a;
    layer4_outputs(3411) <= a and not b;
    layer4_outputs(3412) <= a xor b;
    layer4_outputs(3413) <= not (a and b);
    layer4_outputs(3414) <= a;
    layer4_outputs(3415) <= not a;
    layer4_outputs(3416) <= not a or b;
    layer4_outputs(3417) <= not a;
    layer4_outputs(3418) <= not (a xor b);
    layer4_outputs(3419) <= not b;
    layer4_outputs(3420) <= not a or b;
    layer4_outputs(3421) <= not b;
    layer4_outputs(3422) <= a xor b;
    layer4_outputs(3423) <= not a;
    layer4_outputs(3424) <= not a;
    layer4_outputs(3425) <= a or b;
    layer4_outputs(3426) <= a and not b;
    layer4_outputs(3427) <= a and not b;
    layer4_outputs(3428) <= not b or a;
    layer4_outputs(3429) <= not (a xor b);
    layer4_outputs(3430) <= not a;
    layer4_outputs(3431) <= b;
    layer4_outputs(3432) <= not a or b;
    layer4_outputs(3433) <= a;
    layer4_outputs(3434) <= not a or b;
    layer4_outputs(3435) <= not a or b;
    layer4_outputs(3436) <= not a or b;
    layer4_outputs(3437) <= not a;
    layer4_outputs(3438) <= not a;
    layer4_outputs(3439) <= not a;
    layer4_outputs(3440) <= not (a or b);
    layer4_outputs(3441) <= a;
    layer4_outputs(3442) <= a xor b;
    layer4_outputs(3443) <= not (a or b);
    layer4_outputs(3444) <= a;
    layer4_outputs(3445) <= '1';
    layer4_outputs(3446) <= b and not a;
    layer4_outputs(3447) <= a and not b;
    layer4_outputs(3448) <= a xor b;
    layer4_outputs(3449) <= b and not a;
    layer4_outputs(3450) <= a xor b;
    layer4_outputs(3451) <= b;
    layer4_outputs(3452) <= not a or b;
    layer4_outputs(3453) <= a and b;
    layer4_outputs(3454) <= not (a xor b);
    layer4_outputs(3455) <= not (a or b);
    layer4_outputs(3456) <= not (a or b);
    layer4_outputs(3457) <= a;
    layer4_outputs(3458) <= a;
    layer4_outputs(3459) <= not (a or b);
    layer4_outputs(3460) <= not (a xor b);
    layer4_outputs(3461) <= not b or a;
    layer4_outputs(3462) <= not a;
    layer4_outputs(3463) <= not (a and b);
    layer4_outputs(3464) <= not (a and b);
    layer4_outputs(3465) <= a and not b;
    layer4_outputs(3466) <= not b;
    layer4_outputs(3467) <= a and not b;
    layer4_outputs(3468) <= a;
    layer4_outputs(3469) <= not b or a;
    layer4_outputs(3470) <= a and not b;
    layer4_outputs(3471) <= not (a and b);
    layer4_outputs(3472) <= not a or b;
    layer4_outputs(3473) <= not a;
    layer4_outputs(3474) <= not b;
    layer4_outputs(3475) <= b;
    layer4_outputs(3476) <= a;
    layer4_outputs(3477) <= a and b;
    layer4_outputs(3478) <= not b;
    layer4_outputs(3479) <= a;
    layer4_outputs(3480) <= not b;
    layer4_outputs(3481) <= not b;
    layer4_outputs(3482) <= not (a or b);
    layer4_outputs(3483) <= not a;
    layer4_outputs(3484) <= not b or a;
    layer4_outputs(3485) <= a xor b;
    layer4_outputs(3486) <= not (a or b);
    layer4_outputs(3487) <= not a or b;
    layer4_outputs(3488) <= a xor b;
    layer4_outputs(3489) <= not a;
    layer4_outputs(3490) <= a;
    layer4_outputs(3491) <= not a;
    layer4_outputs(3492) <= not a or b;
    layer4_outputs(3493) <= a and not b;
    layer4_outputs(3494) <= not b;
    layer4_outputs(3495) <= a;
    layer4_outputs(3496) <= b and not a;
    layer4_outputs(3497) <= not a;
    layer4_outputs(3498) <= b and not a;
    layer4_outputs(3499) <= not b or a;
    layer4_outputs(3500) <= a or b;
    layer4_outputs(3501) <= not a or b;
    layer4_outputs(3502) <= a;
    layer4_outputs(3503) <= not a;
    layer4_outputs(3504) <= not (a xor b);
    layer4_outputs(3505) <= a xor b;
    layer4_outputs(3506) <= a;
    layer4_outputs(3507) <= b and not a;
    layer4_outputs(3508) <= not b or a;
    layer4_outputs(3509) <= not a;
    layer4_outputs(3510) <= not a or b;
    layer4_outputs(3511) <= not (a and b);
    layer4_outputs(3512) <= a xor b;
    layer4_outputs(3513) <= b;
    layer4_outputs(3514) <= not b or a;
    layer4_outputs(3515) <= not (a or b);
    layer4_outputs(3516) <= not (a xor b);
    layer4_outputs(3517) <= a xor b;
    layer4_outputs(3518) <= a and not b;
    layer4_outputs(3519) <= a and b;
    layer4_outputs(3520) <= not a;
    layer4_outputs(3521) <= b;
    layer4_outputs(3522) <= a or b;
    layer4_outputs(3523) <= not b;
    layer4_outputs(3524) <= a or b;
    layer4_outputs(3525) <= a or b;
    layer4_outputs(3526) <= not (a xor b);
    layer4_outputs(3527) <= not (a or b);
    layer4_outputs(3528) <= not b;
    layer4_outputs(3529) <= not a;
    layer4_outputs(3530) <= a and b;
    layer4_outputs(3531) <= a and b;
    layer4_outputs(3532) <= b;
    layer4_outputs(3533) <= a and not b;
    layer4_outputs(3534) <= not (a xor b);
    layer4_outputs(3535) <= not (a or b);
    layer4_outputs(3536) <= a;
    layer4_outputs(3537) <= b;
    layer4_outputs(3538) <= a and b;
    layer4_outputs(3539) <= a and not b;
    layer4_outputs(3540) <= not b or a;
    layer4_outputs(3541) <= not (a or b);
    layer4_outputs(3542) <= b;
    layer4_outputs(3543) <= not a or b;
    layer4_outputs(3544) <= a and b;
    layer4_outputs(3545) <= not b;
    layer4_outputs(3546) <= not b;
    layer4_outputs(3547) <= not a;
    layer4_outputs(3548) <= a;
    layer4_outputs(3549) <= b and not a;
    layer4_outputs(3550) <= a and not b;
    layer4_outputs(3551) <= a or b;
    layer4_outputs(3552) <= a and b;
    layer4_outputs(3553) <= b;
    layer4_outputs(3554) <= not (a and b);
    layer4_outputs(3555) <= a;
    layer4_outputs(3556) <= b;
    layer4_outputs(3557) <= a and not b;
    layer4_outputs(3558) <= not b or a;
    layer4_outputs(3559) <= '0';
    layer4_outputs(3560) <= not b;
    layer4_outputs(3561) <= not a;
    layer4_outputs(3562) <= not (a or b);
    layer4_outputs(3563) <= a;
    layer4_outputs(3564) <= a xor b;
    layer4_outputs(3565) <= a or b;
    layer4_outputs(3566) <= not b;
    layer4_outputs(3567) <= not b;
    layer4_outputs(3568) <= a;
    layer4_outputs(3569) <= not a;
    layer4_outputs(3570) <= b;
    layer4_outputs(3571) <= not a;
    layer4_outputs(3572) <= not a or b;
    layer4_outputs(3573) <= not a or b;
    layer4_outputs(3574) <= a;
    layer4_outputs(3575) <= not b;
    layer4_outputs(3576) <= b and not a;
    layer4_outputs(3577) <= not b;
    layer4_outputs(3578) <= not (a xor b);
    layer4_outputs(3579) <= b;
    layer4_outputs(3580) <= not (a xor b);
    layer4_outputs(3581) <= b;
    layer4_outputs(3582) <= b and not a;
    layer4_outputs(3583) <= not a;
    layer4_outputs(3584) <= not a;
    layer4_outputs(3585) <= a or b;
    layer4_outputs(3586) <= not a;
    layer4_outputs(3587) <= a xor b;
    layer4_outputs(3588) <= b;
    layer4_outputs(3589) <= b and not a;
    layer4_outputs(3590) <= not a;
    layer4_outputs(3591) <= a;
    layer4_outputs(3592) <= b;
    layer4_outputs(3593) <= not a;
    layer4_outputs(3594) <= a or b;
    layer4_outputs(3595) <= not (a xor b);
    layer4_outputs(3596) <= not b;
    layer4_outputs(3597) <= a;
    layer4_outputs(3598) <= a or b;
    layer4_outputs(3599) <= a and b;
    layer4_outputs(3600) <= not a or b;
    layer4_outputs(3601) <= not b or a;
    layer4_outputs(3602) <= not (a xor b);
    layer4_outputs(3603) <= not (a or b);
    layer4_outputs(3604) <= not b;
    layer4_outputs(3605) <= a;
    layer4_outputs(3606) <= not (a xor b);
    layer4_outputs(3607) <= a;
    layer4_outputs(3608) <= a;
    layer4_outputs(3609) <= a;
    layer4_outputs(3610) <= not a or b;
    layer4_outputs(3611) <= a and not b;
    layer4_outputs(3612) <= not a;
    layer4_outputs(3613) <= b and not a;
    layer4_outputs(3614) <= a and b;
    layer4_outputs(3615) <= not (a or b);
    layer4_outputs(3616) <= not a or b;
    layer4_outputs(3617) <= not (a and b);
    layer4_outputs(3618) <= not a;
    layer4_outputs(3619) <= a;
    layer4_outputs(3620) <= b;
    layer4_outputs(3621) <= not b;
    layer4_outputs(3622) <= a or b;
    layer4_outputs(3623) <= not (a and b);
    layer4_outputs(3624) <= a;
    layer4_outputs(3625) <= not b;
    layer4_outputs(3626) <= not b;
    layer4_outputs(3627) <= not b or a;
    layer4_outputs(3628) <= b;
    layer4_outputs(3629) <= a or b;
    layer4_outputs(3630) <= a and b;
    layer4_outputs(3631) <= not (a or b);
    layer4_outputs(3632) <= not a or b;
    layer4_outputs(3633) <= not (a or b);
    layer4_outputs(3634) <= b;
    layer4_outputs(3635) <= not b or a;
    layer4_outputs(3636) <= not b or a;
    layer4_outputs(3637) <= not (a xor b);
    layer4_outputs(3638) <= not a;
    layer4_outputs(3639) <= not a;
    layer4_outputs(3640) <= not (a or b);
    layer4_outputs(3641) <= a;
    layer4_outputs(3642) <= not a;
    layer4_outputs(3643) <= b and not a;
    layer4_outputs(3644) <= a;
    layer4_outputs(3645) <= not a;
    layer4_outputs(3646) <= a xor b;
    layer4_outputs(3647) <= b and not a;
    layer4_outputs(3648) <= not (a and b);
    layer4_outputs(3649) <= not a or b;
    layer4_outputs(3650) <= not (a or b);
    layer4_outputs(3651) <= b;
    layer4_outputs(3652) <= b;
    layer4_outputs(3653) <= not (a xor b);
    layer4_outputs(3654) <= a xor b;
    layer4_outputs(3655) <= b;
    layer4_outputs(3656) <= not a or b;
    layer4_outputs(3657) <= b;
    layer4_outputs(3658) <= a;
    layer4_outputs(3659) <= b;
    layer4_outputs(3660) <= not (a and b);
    layer4_outputs(3661) <= not a;
    layer4_outputs(3662) <= a and not b;
    layer4_outputs(3663) <= b and not a;
    layer4_outputs(3664) <= a xor b;
    layer4_outputs(3665) <= a and not b;
    layer4_outputs(3666) <= a;
    layer4_outputs(3667) <= not b;
    layer4_outputs(3668) <= a xor b;
    layer4_outputs(3669) <= not a;
    layer4_outputs(3670) <= a;
    layer4_outputs(3671) <= a and b;
    layer4_outputs(3672) <= not (a or b);
    layer4_outputs(3673) <= b and not a;
    layer4_outputs(3674) <= a and not b;
    layer4_outputs(3675) <= not (a and b);
    layer4_outputs(3676) <= a;
    layer4_outputs(3677) <= b;
    layer4_outputs(3678) <= a xor b;
    layer4_outputs(3679) <= '1';
    layer4_outputs(3680) <= a;
    layer4_outputs(3681) <= not b;
    layer4_outputs(3682) <= not b;
    layer4_outputs(3683) <= not b;
    layer4_outputs(3684) <= not b;
    layer4_outputs(3685) <= not a;
    layer4_outputs(3686) <= not a or b;
    layer4_outputs(3687) <= not (a or b);
    layer4_outputs(3688) <= a xor b;
    layer4_outputs(3689) <= not a or b;
    layer4_outputs(3690) <= not a;
    layer4_outputs(3691) <= not (a xor b);
    layer4_outputs(3692) <= a xor b;
    layer4_outputs(3693) <= not b;
    layer4_outputs(3694) <= not (a and b);
    layer4_outputs(3695) <= not b;
    layer4_outputs(3696) <= b;
    layer4_outputs(3697) <= b;
    layer4_outputs(3698) <= not (a or b);
    layer4_outputs(3699) <= a;
    layer4_outputs(3700) <= not b or a;
    layer4_outputs(3701) <= not a;
    layer4_outputs(3702) <= not a or b;
    layer4_outputs(3703) <= not a;
    layer4_outputs(3704) <= not a or b;
    layer4_outputs(3705) <= a xor b;
    layer4_outputs(3706) <= not (a xor b);
    layer4_outputs(3707) <= a;
    layer4_outputs(3708) <= a;
    layer4_outputs(3709) <= not a or b;
    layer4_outputs(3710) <= a;
    layer4_outputs(3711) <= b;
    layer4_outputs(3712) <= not a or b;
    layer4_outputs(3713) <= a xor b;
    layer4_outputs(3714) <= b and not a;
    layer4_outputs(3715) <= not a or b;
    layer4_outputs(3716) <= not a;
    layer4_outputs(3717) <= a and b;
    layer4_outputs(3718) <= a or b;
    layer4_outputs(3719) <= not a or b;
    layer4_outputs(3720) <= '1';
    layer4_outputs(3721) <= a or b;
    layer4_outputs(3722) <= a xor b;
    layer4_outputs(3723) <= not a;
    layer4_outputs(3724) <= not a;
    layer4_outputs(3725) <= not (a and b);
    layer4_outputs(3726) <= a;
    layer4_outputs(3727) <= not a;
    layer4_outputs(3728) <= b and not a;
    layer4_outputs(3729) <= not (a and b);
    layer4_outputs(3730) <= a and b;
    layer4_outputs(3731) <= a and not b;
    layer4_outputs(3732) <= a and not b;
    layer4_outputs(3733) <= not b or a;
    layer4_outputs(3734) <= not b;
    layer4_outputs(3735) <= not a or b;
    layer4_outputs(3736) <= not (a xor b);
    layer4_outputs(3737) <= not (a or b);
    layer4_outputs(3738) <= b;
    layer4_outputs(3739) <= not (a and b);
    layer4_outputs(3740) <= not a or b;
    layer4_outputs(3741) <= b and not a;
    layer4_outputs(3742) <= not b or a;
    layer4_outputs(3743) <= a xor b;
    layer4_outputs(3744) <= not a;
    layer4_outputs(3745) <= not a;
    layer4_outputs(3746) <= a xor b;
    layer4_outputs(3747) <= not (a and b);
    layer4_outputs(3748) <= a xor b;
    layer4_outputs(3749) <= not b or a;
    layer4_outputs(3750) <= not (a and b);
    layer4_outputs(3751) <= not (a or b);
    layer4_outputs(3752) <= not (a and b);
    layer4_outputs(3753) <= not a;
    layer4_outputs(3754) <= a;
    layer4_outputs(3755) <= a and not b;
    layer4_outputs(3756) <= not (a or b);
    layer4_outputs(3757) <= not (a xor b);
    layer4_outputs(3758) <= a or b;
    layer4_outputs(3759) <= a xor b;
    layer4_outputs(3760) <= a and not b;
    layer4_outputs(3761) <= a;
    layer4_outputs(3762) <= not b or a;
    layer4_outputs(3763) <= not a;
    layer4_outputs(3764) <= not a;
    layer4_outputs(3765) <= a and b;
    layer4_outputs(3766) <= a;
    layer4_outputs(3767) <= a or b;
    layer4_outputs(3768) <= not b;
    layer4_outputs(3769) <= not a or b;
    layer4_outputs(3770) <= not (a or b);
    layer4_outputs(3771) <= a;
    layer4_outputs(3772) <= a;
    layer4_outputs(3773) <= not (a and b);
    layer4_outputs(3774) <= not b;
    layer4_outputs(3775) <= a and b;
    layer4_outputs(3776) <= b and not a;
    layer4_outputs(3777) <= a;
    layer4_outputs(3778) <= a and b;
    layer4_outputs(3779) <= b and not a;
    layer4_outputs(3780) <= a and b;
    layer4_outputs(3781) <= a;
    layer4_outputs(3782) <= b;
    layer4_outputs(3783) <= b and not a;
    layer4_outputs(3784) <= not b;
    layer4_outputs(3785) <= b;
    layer4_outputs(3786) <= a;
    layer4_outputs(3787) <= not a;
    layer4_outputs(3788) <= not (a xor b);
    layer4_outputs(3789) <= a and not b;
    layer4_outputs(3790) <= b;
    layer4_outputs(3791) <= not a or b;
    layer4_outputs(3792) <= not a or b;
    layer4_outputs(3793) <= a;
    layer4_outputs(3794) <= not a;
    layer4_outputs(3795) <= not (a xor b);
    layer4_outputs(3796) <= b;
    layer4_outputs(3797) <= not (a or b);
    layer4_outputs(3798) <= b;
    layer4_outputs(3799) <= not a;
    layer4_outputs(3800) <= not (a xor b);
    layer4_outputs(3801) <= not a;
    layer4_outputs(3802) <= not b;
    layer4_outputs(3803) <= not (a and b);
    layer4_outputs(3804) <= not (a or b);
    layer4_outputs(3805) <= a and b;
    layer4_outputs(3806) <= b;
    layer4_outputs(3807) <= not a;
    layer4_outputs(3808) <= b and not a;
    layer4_outputs(3809) <= a;
    layer4_outputs(3810) <= not a;
    layer4_outputs(3811) <= '1';
    layer4_outputs(3812) <= not a or b;
    layer4_outputs(3813) <= not (a xor b);
    layer4_outputs(3814) <= not a;
    layer4_outputs(3815) <= '0';
    layer4_outputs(3816) <= a and b;
    layer4_outputs(3817) <= a or b;
    layer4_outputs(3818) <= a or b;
    layer4_outputs(3819) <= a xor b;
    layer4_outputs(3820) <= not a or b;
    layer4_outputs(3821) <= not a;
    layer4_outputs(3822) <= a and b;
    layer4_outputs(3823) <= not a or b;
    layer4_outputs(3824) <= not a;
    layer4_outputs(3825) <= b;
    layer4_outputs(3826) <= b and not a;
    layer4_outputs(3827) <= not b;
    layer4_outputs(3828) <= b;
    layer4_outputs(3829) <= not a or b;
    layer4_outputs(3830) <= a or b;
    layer4_outputs(3831) <= not b or a;
    layer4_outputs(3832) <= not (a or b);
    layer4_outputs(3833) <= '0';
    layer4_outputs(3834) <= a xor b;
    layer4_outputs(3835) <= not b;
    layer4_outputs(3836) <= b;
    layer4_outputs(3837) <= not b or a;
    layer4_outputs(3838) <= a xor b;
    layer4_outputs(3839) <= '0';
    layer4_outputs(3840) <= a;
    layer4_outputs(3841) <= not (a or b);
    layer4_outputs(3842) <= a and not b;
    layer4_outputs(3843) <= a xor b;
    layer4_outputs(3844) <= b and not a;
    layer4_outputs(3845) <= not (a and b);
    layer4_outputs(3846) <= b;
    layer4_outputs(3847) <= b and not a;
    layer4_outputs(3848) <= not (a and b);
    layer4_outputs(3849) <= not a;
    layer4_outputs(3850) <= a or b;
    layer4_outputs(3851) <= b;
    layer4_outputs(3852) <= not a;
    layer4_outputs(3853) <= not (a xor b);
    layer4_outputs(3854) <= not (a or b);
    layer4_outputs(3855) <= a and b;
    layer4_outputs(3856) <= a or b;
    layer4_outputs(3857) <= a and b;
    layer4_outputs(3858) <= a and not b;
    layer4_outputs(3859) <= b and not a;
    layer4_outputs(3860) <= not a;
    layer4_outputs(3861) <= '1';
    layer4_outputs(3862) <= not b;
    layer4_outputs(3863) <= not (a or b);
    layer4_outputs(3864) <= a and not b;
    layer4_outputs(3865) <= a and not b;
    layer4_outputs(3866) <= a xor b;
    layer4_outputs(3867) <= not (a or b);
    layer4_outputs(3868) <= b and not a;
    layer4_outputs(3869) <= b and not a;
    layer4_outputs(3870) <= not (a xor b);
    layer4_outputs(3871) <= a xor b;
    layer4_outputs(3872) <= not b;
    layer4_outputs(3873) <= not a;
    layer4_outputs(3874) <= b;
    layer4_outputs(3875) <= not a;
    layer4_outputs(3876) <= not (a and b);
    layer4_outputs(3877) <= not a or b;
    layer4_outputs(3878) <= a or b;
    layer4_outputs(3879) <= not a or b;
    layer4_outputs(3880) <= not a or b;
    layer4_outputs(3881) <= a or b;
    layer4_outputs(3882) <= b;
    layer4_outputs(3883) <= not (a xor b);
    layer4_outputs(3884) <= not b;
    layer4_outputs(3885) <= not a;
    layer4_outputs(3886) <= not a;
    layer4_outputs(3887) <= not (a and b);
    layer4_outputs(3888) <= a;
    layer4_outputs(3889) <= not a or b;
    layer4_outputs(3890) <= a or b;
    layer4_outputs(3891) <= a;
    layer4_outputs(3892) <= not b or a;
    layer4_outputs(3893) <= not b or a;
    layer4_outputs(3894) <= a or b;
    layer4_outputs(3895) <= not b;
    layer4_outputs(3896) <= b and not a;
    layer4_outputs(3897) <= not a;
    layer4_outputs(3898) <= a and not b;
    layer4_outputs(3899) <= not (a or b);
    layer4_outputs(3900) <= a;
    layer4_outputs(3901) <= a and b;
    layer4_outputs(3902) <= a and b;
    layer4_outputs(3903) <= '0';
    layer4_outputs(3904) <= not a;
    layer4_outputs(3905) <= not (a or b);
    layer4_outputs(3906) <= b;
    layer4_outputs(3907) <= a or b;
    layer4_outputs(3908) <= b;
    layer4_outputs(3909) <= not b;
    layer4_outputs(3910) <= not b or a;
    layer4_outputs(3911) <= not b or a;
    layer4_outputs(3912) <= a;
    layer4_outputs(3913) <= '0';
    layer4_outputs(3914) <= not (a or b);
    layer4_outputs(3915) <= b and not a;
    layer4_outputs(3916) <= not a;
    layer4_outputs(3917) <= not a;
    layer4_outputs(3918) <= not (a and b);
    layer4_outputs(3919) <= not a or b;
    layer4_outputs(3920) <= not a;
    layer4_outputs(3921) <= a or b;
    layer4_outputs(3922) <= not (a or b);
    layer4_outputs(3923) <= a;
    layer4_outputs(3924) <= a;
    layer4_outputs(3925) <= b and not a;
    layer4_outputs(3926) <= not a or b;
    layer4_outputs(3927) <= a or b;
    layer4_outputs(3928) <= a and not b;
    layer4_outputs(3929) <= not b or a;
    layer4_outputs(3930) <= a xor b;
    layer4_outputs(3931) <= not a or b;
    layer4_outputs(3932) <= not b;
    layer4_outputs(3933) <= not (a xor b);
    layer4_outputs(3934) <= not (a or b);
    layer4_outputs(3935) <= b;
    layer4_outputs(3936) <= not b;
    layer4_outputs(3937) <= not (a xor b);
    layer4_outputs(3938) <= not b;
    layer4_outputs(3939) <= not a or b;
    layer4_outputs(3940) <= not (a and b);
    layer4_outputs(3941) <= not (a or b);
    layer4_outputs(3942) <= a xor b;
    layer4_outputs(3943) <= b;
    layer4_outputs(3944) <= not (a and b);
    layer4_outputs(3945) <= not b;
    layer4_outputs(3946) <= not (a and b);
    layer4_outputs(3947) <= not b or a;
    layer4_outputs(3948) <= not (a xor b);
    layer4_outputs(3949) <= not a;
    layer4_outputs(3950) <= a and not b;
    layer4_outputs(3951) <= b and not a;
    layer4_outputs(3952) <= a or b;
    layer4_outputs(3953) <= a;
    layer4_outputs(3954) <= not (a and b);
    layer4_outputs(3955) <= b and not a;
    layer4_outputs(3956) <= not a or b;
    layer4_outputs(3957) <= not (a xor b);
    layer4_outputs(3958) <= not (a or b);
    layer4_outputs(3959) <= a xor b;
    layer4_outputs(3960) <= not (a xor b);
    layer4_outputs(3961) <= a;
    layer4_outputs(3962) <= a and b;
    layer4_outputs(3963) <= a;
    layer4_outputs(3964) <= b;
    layer4_outputs(3965) <= not b;
    layer4_outputs(3966) <= not (a or b);
    layer4_outputs(3967) <= a and not b;
    layer4_outputs(3968) <= a and b;
    layer4_outputs(3969) <= not a or b;
    layer4_outputs(3970) <= a and not b;
    layer4_outputs(3971) <= not b;
    layer4_outputs(3972) <= not (a or b);
    layer4_outputs(3973) <= not b;
    layer4_outputs(3974) <= a or b;
    layer4_outputs(3975) <= b;
    layer4_outputs(3976) <= not a or b;
    layer4_outputs(3977) <= '0';
    layer4_outputs(3978) <= not (a or b);
    layer4_outputs(3979) <= a xor b;
    layer4_outputs(3980) <= not b or a;
    layer4_outputs(3981) <= not (a and b);
    layer4_outputs(3982) <= not a or b;
    layer4_outputs(3983) <= not b;
    layer4_outputs(3984) <= not b;
    layer4_outputs(3985) <= not a;
    layer4_outputs(3986) <= a;
    layer4_outputs(3987) <= a or b;
    layer4_outputs(3988) <= a xor b;
    layer4_outputs(3989) <= b;
    layer4_outputs(3990) <= a or b;
    layer4_outputs(3991) <= not (a xor b);
    layer4_outputs(3992) <= not a or b;
    layer4_outputs(3993) <= not a;
    layer4_outputs(3994) <= '1';
    layer4_outputs(3995) <= not b or a;
    layer4_outputs(3996) <= a or b;
    layer4_outputs(3997) <= not a;
    layer4_outputs(3998) <= a and b;
    layer4_outputs(3999) <= not (a and b);
    layer4_outputs(4000) <= not b or a;
    layer4_outputs(4001) <= not b;
    layer4_outputs(4002) <= not b;
    layer4_outputs(4003) <= a and not b;
    layer4_outputs(4004) <= not b or a;
    layer4_outputs(4005) <= not a;
    layer4_outputs(4006) <= a;
    layer4_outputs(4007) <= not a or b;
    layer4_outputs(4008) <= a;
    layer4_outputs(4009) <= '1';
    layer4_outputs(4010) <= a and not b;
    layer4_outputs(4011) <= b;
    layer4_outputs(4012) <= not (a or b);
    layer4_outputs(4013) <= not (a or b);
    layer4_outputs(4014) <= not b;
    layer4_outputs(4015) <= not a or b;
    layer4_outputs(4016) <= not b or a;
    layer4_outputs(4017) <= b;
    layer4_outputs(4018) <= b;
    layer4_outputs(4019) <= not a or b;
    layer4_outputs(4020) <= not a or b;
    layer4_outputs(4021) <= a xor b;
    layer4_outputs(4022) <= not b;
    layer4_outputs(4023) <= not a;
    layer4_outputs(4024) <= not (a xor b);
    layer4_outputs(4025) <= not a or b;
    layer4_outputs(4026) <= a and not b;
    layer4_outputs(4027) <= not (a and b);
    layer4_outputs(4028) <= '0';
    layer4_outputs(4029) <= a or b;
    layer4_outputs(4030) <= not a;
    layer4_outputs(4031) <= not (a xor b);
    layer4_outputs(4032) <= not (a xor b);
    layer4_outputs(4033) <= not a;
    layer4_outputs(4034) <= not a;
    layer4_outputs(4035) <= not b;
    layer4_outputs(4036) <= a and b;
    layer4_outputs(4037) <= b and not a;
    layer4_outputs(4038) <= not b or a;
    layer4_outputs(4039) <= a or b;
    layer4_outputs(4040) <= b;
    layer4_outputs(4041) <= a;
    layer4_outputs(4042) <= a;
    layer4_outputs(4043) <= not b or a;
    layer4_outputs(4044) <= not b;
    layer4_outputs(4045) <= a;
    layer4_outputs(4046) <= not a;
    layer4_outputs(4047) <= not a or b;
    layer4_outputs(4048) <= b and not a;
    layer4_outputs(4049) <= '1';
    layer4_outputs(4050) <= a and b;
    layer4_outputs(4051) <= not a;
    layer4_outputs(4052) <= not (a xor b);
    layer4_outputs(4053) <= not a;
    layer4_outputs(4054) <= not (a or b);
    layer4_outputs(4055) <= not (a and b);
    layer4_outputs(4056) <= not (a and b);
    layer4_outputs(4057) <= not b;
    layer4_outputs(4058) <= b;
    layer4_outputs(4059) <= not a;
    layer4_outputs(4060) <= a and b;
    layer4_outputs(4061) <= b;
    layer4_outputs(4062) <= b;
    layer4_outputs(4063) <= not (a or b);
    layer4_outputs(4064) <= a;
    layer4_outputs(4065) <= not (a xor b);
    layer4_outputs(4066) <= b;
    layer4_outputs(4067) <= b and not a;
    layer4_outputs(4068) <= not b or a;
    layer4_outputs(4069) <= b;
    layer4_outputs(4070) <= not b or a;
    layer4_outputs(4071) <= b;
    layer4_outputs(4072) <= not a;
    layer4_outputs(4073) <= b;
    layer4_outputs(4074) <= a and not b;
    layer4_outputs(4075) <= a xor b;
    layer4_outputs(4076) <= a xor b;
    layer4_outputs(4077) <= not (a or b);
    layer4_outputs(4078) <= b;
    layer4_outputs(4079) <= not (a and b);
    layer4_outputs(4080) <= b;
    layer4_outputs(4081) <= a or b;
    layer4_outputs(4082) <= not (a xor b);
    layer4_outputs(4083) <= b and not a;
    layer4_outputs(4084) <= a;
    layer4_outputs(4085) <= a;
    layer4_outputs(4086) <= not a;
    layer4_outputs(4087) <= not (a xor b);
    layer4_outputs(4088) <= not a or b;
    layer4_outputs(4089) <= not b;
    layer4_outputs(4090) <= b and not a;
    layer4_outputs(4091) <= a and b;
    layer4_outputs(4092) <= not (a xor b);
    layer4_outputs(4093) <= not a or b;
    layer4_outputs(4094) <= not b or a;
    layer4_outputs(4095) <= b;
    layer4_outputs(4096) <= a or b;
    layer4_outputs(4097) <= a and b;
    layer4_outputs(4098) <= not b or a;
    layer4_outputs(4099) <= not b or a;
    layer4_outputs(4100) <= not (a and b);
    layer4_outputs(4101) <= not a;
    layer4_outputs(4102) <= b;
    layer4_outputs(4103) <= b;
    layer4_outputs(4104) <= a and b;
    layer4_outputs(4105) <= a and not b;
    layer4_outputs(4106) <= not a;
    layer4_outputs(4107) <= b;
    layer4_outputs(4108) <= not (a xor b);
    layer4_outputs(4109) <= not (a xor b);
    layer4_outputs(4110) <= a and not b;
    layer4_outputs(4111) <= a xor b;
    layer4_outputs(4112) <= a xor b;
    layer4_outputs(4113) <= a and not b;
    layer4_outputs(4114) <= not b or a;
    layer4_outputs(4115) <= b;
    layer4_outputs(4116) <= not b;
    layer4_outputs(4117) <= not (a xor b);
    layer4_outputs(4118) <= not (a or b);
    layer4_outputs(4119) <= a and not b;
    layer4_outputs(4120) <= not b;
    layer4_outputs(4121) <= a and b;
    layer4_outputs(4122) <= a;
    layer4_outputs(4123) <= not b;
    layer4_outputs(4124) <= not a;
    layer4_outputs(4125) <= a;
    layer4_outputs(4126) <= not b;
    layer4_outputs(4127) <= not (a and b);
    layer4_outputs(4128) <= a and b;
    layer4_outputs(4129) <= a and b;
    layer4_outputs(4130) <= b;
    layer4_outputs(4131) <= not b or a;
    layer4_outputs(4132) <= not (a xor b);
    layer4_outputs(4133) <= a and b;
    layer4_outputs(4134) <= a xor b;
    layer4_outputs(4135) <= a;
    layer4_outputs(4136) <= not (a xor b);
    layer4_outputs(4137) <= a;
    layer4_outputs(4138) <= a;
    layer4_outputs(4139) <= not (a or b);
    layer4_outputs(4140) <= a and not b;
    layer4_outputs(4141) <= a;
    layer4_outputs(4142) <= a;
    layer4_outputs(4143) <= a or b;
    layer4_outputs(4144) <= b and not a;
    layer4_outputs(4145) <= not a;
    layer4_outputs(4146) <= a;
    layer4_outputs(4147) <= not b;
    layer4_outputs(4148) <= b;
    layer4_outputs(4149) <= not b;
    layer4_outputs(4150) <= not b;
    layer4_outputs(4151) <= b;
    layer4_outputs(4152) <= b and not a;
    layer4_outputs(4153) <= not b;
    layer4_outputs(4154) <= a;
    layer4_outputs(4155) <= a xor b;
    layer4_outputs(4156) <= b and not a;
    layer4_outputs(4157) <= not (a xor b);
    layer4_outputs(4158) <= not (a xor b);
    layer4_outputs(4159) <= not a;
    layer4_outputs(4160) <= a;
    layer4_outputs(4161) <= a;
    layer4_outputs(4162) <= not (a xor b);
    layer4_outputs(4163) <= b and not a;
    layer4_outputs(4164) <= not a or b;
    layer4_outputs(4165) <= b and not a;
    layer4_outputs(4166) <= a;
    layer4_outputs(4167) <= b;
    layer4_outputs(4168) <= a and not b;
    layer4_outputs(4169) <= not b;
    layer4_outputs(4170) <= a and b;
    layer4_outputs(4171) <= a or b;
    layer4_outputs(4172) <= a and not b;
    layer4_outputs(4173) <= not a or b;
    layer4_outputs(4174) <= not a;
    layer4_outputs(4175) <= b;
    layer4_outputs(4176) <= not (a xor b);
    layer4_outputs(4177) <= not b;
    layer4_outputs(4178) <= not b;
    layer4_outputs(4179) <= a;
    layer4_outputs(4180) <= b;
    layer4_outputs(4181) <= not a;
    layer4_outputs(4182) <= not b;
    layer4_outputs(4183) <= a;
    layer4_outputs(4184) <= b;
    layer4_outputs(4185) <= not b;
    layer4_outputs(4186) <= a;
    layer4_outputs(4187) <= not a;
    layer4_outputs(4188) <= not b;
    layer4_outputs(4189) <= not b;
    layer4_outputs(4190) <= not a or b;
    layer4_outputs(4191) <= not (a and b);
    layer4_outputs(4192) <= b and not a;
    layer4_outputs(4193) <= a xor b;
    layer4_outputs(4194) <= a;
    layer4_outputs(4195) <= b;
    layer4_outputs(4196) <= not a;
    layer4_outputs(4197) <= not b;
    layer4_outputs(4198) <= b and not a;
    layer4_outputs(4199) <= not a;
    layer4_outputs(4200) <= a and not b;
    layer4_outputs(4201) <= '1';
    layer4_outputs(4202) <= not (a xor b);
    layer4_outputs(4203) <= not a;
    layer4_outputs(4204) <= a or b;
    layer4_outputs(4205) <= not b;
    layer4_outputs(4206) <= a;
    layer4_outputs(4207) <= a;
    layer4_outputs(4208) <= not (a xor b);
    layer4_outputs(4209) <= a;
    layer4_outputs(4210) <= not a or b;
    layer4_outputs(4211) <= a or b;
    layer4_outputs(4212) <= b and not a;
    layer4_outputs(4213) <= not b;
    layer4_outputs(4214) <= not (a and b);
    layer4_outputs(4215) <= a;
    layer4_outputs(4216) <= not b or a;
    layer4_outputs(4217) <= not b or a;
    layer4_outputs(4218) <= a;
    layer4_outputs(4219) <= a and b;
    layer4_outputs(4220) <= b and not a;
    layer4_outputs(4221) <= not b;
    layer4_outputs(4222) <= a xor b;
    layer4_outputs(4223) <= a;
    layer4_outputs(4224) <= not (a and b);
    layer4_outputs(4225) <= a or b;
    layer4_outputs(4226) <= not a;
    layer4_outputs(4227) <= a and not b;
    layer4_outputs(4228) <= not (a or b);
    layer4_outputs(4229) <= b and not a;
    layer4_outputs(4230) <= a xor b;
    layer4_outputs(4231) <= b;
    layer4_outputs(4232) <= a xor b;
    layer4_outputs(4233) <= a and not b;
    layer4_outputs(4234) <= b;
    layer4_outputs(4235) <= a;
    layer4_outputs(4236) <= not b or a;
    layer4_outputs(4237) <= a;
    layer4_outputs(4238) <= a or b;
    layer4_outputs(4239) <= not b;
    layer4_outputs(4240) <= a;
    layer4_outputs(4241) <= b;
    layer4_outputs(4242) <= not (a and b);
    layer4_outputs(4243) <= b;
    layer4_outputs(4244) <= not b;
    layer4_outputs(4245) <= not a;
    layer4_outputs(4246) <= not a or b;
    layer4_outputs(4247) <= not b;
    layer4_outputs(4248) <= not (a and b);
    layer4_outputs(4249) <= b;
    layer4_outputs(4250) <= a;
    layer4_outputs(4251) <= a;
    layer4_outputs(4252) <= a xor b;
    layer4_outputs(4253) <= not a;
    layer4_outputs(4254) <= a xor b;
    layer4_outputs(4255) <= a or b;
    layer4_outputs(4256) <= not a;
    layer4_outputs(4257) <= not b;
    layer4_outputs(4258) <= not (a or b);
    layer4_outputs(4259) <= a and not b;
    layer4_outputs(4260) <= a or b;
    layer4_outputs(4261) <= not (a xor b);
    layer4_outputs(4262) <= a and b;
    layer4_outputs(4263) <= a;
    layer4_outputs(4264) <= b;
    layer4_outputs(4265) <= a or b;
    layer4_outputs(4266) <= b;
    layer4_outputs(4267) <= not a;
    layer4_outputs(4268) <= b and not a;
    layer4_outputs(4269) <= a xor b;
    layer4_outputs(4270) <= not a or b;
    layer4_outputs(4271) <= not (a or b);
    layer4_outputs(4272) <= a;
    layer4_outputs(4273) <= a xor b;
    layer4_outputs(4274) <= not b;
    layer4_outputs(4275) <= not b;
    layer4_outputs(4276) <= not a;
    layer4_outputs(4277) <= not (a and b);
    layer4_outputs(4278) <= a and not b;
    layer4_outputs(4279) <= a;
    layer4_outputs(4280) <= not (a or b);
    layer4_outputs(4281) <= not (a or b);
    layer4_outputs(4282) <= a;
    layer4_outputs(4283) <= not (a or b);
    layer4_outputs(4284) <= a;
    layer4_outputs(4285) <= not b or a;
    layer4_outputs(4286) <= not (a and b);
    layer4_outputs(4287) <= not a;
    layer4_outputs(4288) <= not (a xor b);
    layer4_outputs(4289) <= not a or b;
    layer4_outputs(4290) <= not a;
    layer4_outputs(4291) <= not a;
    layer4_outputs(4292) <= '1';
    layer4_outputs(4293) <= not (a and b);
    layer4_outputs(4294) <= not (a xor b);
    layer4_outputs(4295) <= a xor b;
    layer4_outputs(4296) <= '1';
    layer4_outputs(4297) <= a;
    layer4_outputs(4298) <= not a or b;
    layer4_outputs(4299) <= a;
    layer4_outputs(4300) <= not b;
    layer4_outputs(4301) <= not b or a;
    layer4_outputs(4302) <= b and not a;
    layer4_outputs(4303) <= not (a or b);
    layer4_outputs(4304) <= not (a and b);
    layer4_outputs(4305) <= not (a xor b);
    layer4_outputs(4306) <= a and not b;
    layer4_outputs(4307) <= not a or b;
    layer4_outputs(4308) <= not b or a;
    layer4_outputs(4309) <= b;
    layer4_outputs(4310) <= not b;
    layer4_outputs(4311) <= not b;
    layer4_outputs(4312) <= not b or a;
    layer4_outputs(4313) <= not b or a;
    layer4_outputs(4314) <= not a or b;
    layer4_outputs(4315) <= b and not a;
    layer4_outputs(4316) <= a or b;
    layer4_outputs(4317) <= not a or b;
    layer4_outputs(4318) <= a or b;
    layer4_outputs(4319) <= b;
    layer4_outputs(4320) <= not b;
    layer4_outputs(4321) <= a;
    layer4_outputs(4322) <= a;
    layer4_outputs(4323) <= not (a and b);
    layer4_outputs(4324) <= not (a and b);
    layer4_outputs(4325) <= a and not b;
    layer4_outputs(4326) <= a;
    layer4_outputs(4327) <= not (a and b);
    layer4_outputs(4328) <= a and not b;
    layer4_outputs(4329) <= b;
    layer4_outputs(4330) <= a or b;
    layer4_outputs(4331) <= a;
    layer4_outputs(4332) <= not b or a;
    layer4_outputs(4333) <= a or b;
    layer4_outputs(4334) <= a;
    layer4_outputs(4335) <= '0';
    layer4_outputs(4336) <= b;
    layer4_outputs(4337) <= a;
    layer4_outputs(4338) <= a xor b;
    layer4_outputs(4339) <= not (a and b);
    layer4_outputs(4340) <= not a;
    layer4_outputs(4341) <= a and b;
    layer4_outputs(4342) <= b;
    layer4_outputs(4343) <= not b;
    layer4_outputs(4344) <= not a;
    layer4_outputs(4345) <= not b;
    layer4_outputs(4346) <= a or b;
    layer4_outputs(4347) <= not (a and b);
    layer4_outputs(4348) <= not b;
    layer4_outputs(4349) <= a;
    layer4_outputs(4350) <= a;
    layer4_outputs(4351) <= not b;
    layer4_outputs(4352) <= not a;
    layer4_outputs(4353) <= not (a and b);
    layer4_outputs(4354) <= b;
    layer4_outputs(4355) <= b;
    layer4_outputs(4356) <= not (a or b);
    layer4_outputs(4357) <= a;
    layer4_outputs(4358) <= b;
    layer4_outputs(4359) <= not b or a;
    layer4_outputs(4360) <= not b;
    layer4_outputs(4361) <= a or b;
    layer4_outputs(4362) <= not (a xor b);
    layer4_outputs(4363) <= b and not a;
    layer4_outputs(4364) <= not a or b;
    layer4_outputs(4365) <= a;
    layer4_outputs(4366) <= b;
    layer4_outputs(4367) <= not a or b;
    layer4_outputs(4368) <= not (a xor b);
    layer4_outputs(4369) <= b and not a;
    layer4_outputs(4370) <= not b;
    layer4_outputs(4371) <= '0';
    layer4_outputs(4372) <= b;
    layer4_outputs(4373) <= not a;
    layer4_outputs(4374) <= not a;
    layer4_outputs(4375) <= a;
    layer4_outputs(4376) <= not b;
    layer4_outputs(4377) <= not a or b;
    layer4_outputs(4378) <= a;
    layer4_outputs(4379) <= not (a xor b);
    layer4_outputs(4380) <= a and not b;
    layer4_outputs(4381) <= not (a xor b);
    layer4_outputs(4382) <= not a;
    layer4_outputs(4383) <= a and b;
    layer4_outputs(4384) <= b;
    layer4_outputs(4385) <= a or b;
    layer4_outputs(4386) <= a and b;
    layer4_outputs(4387) <= b;
    layer4_outputs(4388) <= a;
    layer4_outputs(4389) <= not (a xor b);
    layer4_outputs(4390) <= not b;
    layer4_outputs(4391) <= a and not b;
    layer4_outputs(4392) <= a and not b;
    layer4_outputs(4393) <= a;
    layer4_outputs(4394) <= not a or b;
    layer4_outputs(4395) <= a;
    layer4_outputs(4396) <= a and not b;
    layer4_outputs(4397) <= not a;
    layer4_outputs(4398) <= not b;
    layer4_outputs(4399) <= not (a or b);
    layer4_outputs(4400) <= not (a and b);
    layer4_outputs(4401) <= not (a xor b);
    layer4_outputs(4402) <= not b;
    layer4_outputs(4403) <= not a;
    layer4_outputs(4404) <= not b;
    layer4_outputs(4405) <= b and not a;
    layer4_outputs(4406) <= not (a xor b);
    layer4_outputs(4407) <= not (a xor b);
    layer4_outputs(4408) <= not a;
    layer4_outputs(4409) <= b;
    layer4_outputs(4410) <= a xor b;
    layer4_outputs(4411) <= a and not b;
    layer4_outputs(4412) <= a or b;
    layer4_outputs(4413) <= not b or a;
    layer4_outputs(4414) <= not b or a;
    layer4_outputs(4415) <= not (a xor b);
    layer4_outputs(4416) <= a;
    layer4_outputs(4417) <= a;
    layer4_outputs(4418) <= b;
    layer4_outputs(4419) <= not (a and b);
    layer4_outputs(4420) <= a;
    layer4_outputs(4421) <= not (a and b);
    layer4_outputs(4422) <= '0';
    layer4_outputs(4423) <= b;
    layer4_outputs(4424) <= not (a xor b);
    layer4_outputs(4425) <= not a;
    layer4_outputs(4426) <= not a;
    layer4_outputs(4427) <= not a;
    layer4_outputs(4428) <= a xor b;
    layer4_outputs(4429) <= a or b;
    layer4_outputs(4430) <= a or b;
    layer4_outputs(4431) <= not b or a;
    layer4_outputs(4432) <= not (a or b);
    layer4_outputs(4433) <= b and not a;
    layer4_outputs(4434) <= not b;
    layer4_outputs(4435) <= not b;
    layer4_outputs(4436) <= a xor b;
    layer4_outputs(4437) <= a and not b;
    layer4_outputs(4438) <= a xor b;
    layer4_outputs(4439) <= not b;
    layer4_outputs(4440) <= not (a and b);
    layer4_outputs(4441) <= a xor b;
    layer4_outputs(4442) <= not a;
    layer4_outputs(4443) <= not (a xor b);
    layer4_outputs(4444) <= not a;
    layer4_outputs(4445) <= a and not b;
    layer4_outputs(4446) <= not b or a;
    layer4_outputs(4447) <= a xor b;
    layer4_outputs(4448) <= not b;
    layer4_outputs(4449) <= b and not a;
    layer4_outputs(4450) <= not a;
    layer4_outputs(4451) <= a;
    layer4_outputs(4452) <= b;
    layer4_outputs(4453) <= a and b;
    layer4_outputs(4454) <= not (a xor b);
    layer4_outputs(4455) <= not a or b;
    layer4_outputs(4456) <= not b or a;
    layer4_outputs(4457) <= b and not a;
    layer4_outputs(4458) <= not a;
    layer4_outputs(4459) <= a xor b;
    layer4_outputs(4460) <= a and b;
    layer4_outputs(4461) <= a and b;
    layer4_outputs(4462) <= b;
    layer4_outputs(4463) <= b;
    layer4_outputs(4464) <= a;
    layer4_outputs(4465) <= a;
    layer4_outputs(4466) <= not a;
    layer4_outputs(4467) <= a or b;
    layer4_outputs(4468) <= a or b;
    layer4_outputs(4469) <= a;
    layer4_outputs(4470) <= not (a and b);
    layer4_outputs(4471) <= a;
    layer4_outputs(4472) <= not a;
    layer4_outputs(4473) <= not b;
    layer4_outputs(4474) <= not b;
    layer4_outputs(4475) <= a xor b;
    layer4_outputs(4476) <= b and not a;
    layer4_outputs(4477) <= not (a and b);
    layer4_outputs(4478) <= b;
    layer4_outputs(4479) <= a;
    layer4_outputs(4480) <= not (a and b);
    layer4_outputs(4481) <= not (a and b);
    layer4_outputs(4482) <= b and not a;
    layer4_outputs(4483) <= a;
    layer4_outputs(4484) <= a and b;
    layer4_outputs(4485) <= '1';
    layer4_outputs(4486) <= not b;
    layer4_outputs(4487) <= a;
    layer4_outputs(4488) <= not b;
    layer4_outputs(4489) <= not a;
    layer4_outputs(4490) <= not b or a;
    layer4_outputs(4491) <= not (a xor b);
    layer4_outputs(4492) <= not b;
    layer4_outputs(4493) <= b and not a;
    layer4_outputs(4494) <= b;
    layer4_outputs(4495) <= not a;
    layer4_outputs(4496) <= b and not a;
    layer4_outputs(4497) <= not (a xor b);
    layer4_outputs(4498) <= a and b;
    layer4_outputs(4499) <= not b;
    layer4_outputs(4500) <= not (a or b);
    layer4_outputs(4501) <= a xor b;
    layer4_outputs(4502) <= not (a and b);
    layer4_outputs(4503) <= a;
    layer4_outputs(4504) <= a;
    layer4_outputs(4505) <= b and not a;
    layer4_outputs(4506) <= a;
    layer4_outputs(4507) <= a;
    layer4_outputs(4508) <= a and not b;
    layer4_outputs(4509) <= not (a xor b);
    layer4_outputs(4510) <= b and not a;
    layer4_outputs(4511) <= '0';
    layer4_outputs(4512) <= a or b;
    layer4_outputs(4513) <= a xor b;
    layer4_outputs(4514) <= b and not a;
    layer4_outputs(4515) <= not a;
    layer4_outputs(4516) <= not (a xor b);
    layer4_outputs(4517) <= not b;
    layer4_outputs(4518) <= a or b;
    layer4_outputs(4519) <= not a;
    layer4_outputs(4520) <= a and b;
    layer4_outputs(4521) <= not a or b;
    layer4_outputs(4522) <= not (a xor b);
    layer4_outputs(4523) <= b;
    layer4_outputs(4524) <= not (a or b);
    layer4_outputs(4525) <= a;
    layer4_outputs(4526) <= not b;
    layer4_outputs(4527) <= not (a or b);
    layer4_outputs(4528) <= not (a xor b);
    layer4_outputs(4529) <= not b;
    layer4_outputs(4530) <= a and not b;
    layer4_outputs(4531) <= not (a and b);
    layer4_outputs(4532) <= not a;
    layer4_outputs(4533) <= not a;
    layer4_outputs(4534) <= not a;
    layer4_outputs(4535) <= not (a and b);
    layer4_outputs(4536) <= b;
    layer4_outputs(4537) <= b and not a;
    layer4_outputs(4538) <= a and b;
    layer4_outputs(4539) <= b and not a;
    layer4_outputs(4540) <= a and b;
    layer4_outputs(4541) <= a;
    layer4_outputs(4542) <= b;
    layer4_outputs(4543) <= not b or a;
    layer4_outputs(4544) <= not b;
    layer4_outputs(4545) <= a;
    layer4_outputs(4546) <= a and not b;
    layer4_outputs(4547) <= b and not a;
    layer4_outputs(4548) <= not b;
    layer4_outputs(4549) <= not (a and b);
    layer4_outputs(4550) <= b and not a;
    layer4_outputs(4551) <= b;
    layer4_outputs(4552) <= b and not a;
    layer4_outputs(4553) <= not b;
    layer4_outputs(4554) <= b;
    layer4_outputs(4555) <= a;
    layer4_outputs(4556) <= not (a xor b);
    layer4_outputs(4557) <= a and not b;
    layer4_outputs(4558) <= a and not b;
    layer4_outputs(4559) <= not b;
    layer4_outputs(4560) <= b;
    layer4_outputs(4561) <= not (a xor b);
    layer4_outputs(4562) <= a;
    layer4_outputs(4563) <= not (a xor b);
    layer4_outputs(4564) <= b;
    layer4_outputs(4565) <= not a;
    layer4_outputs(4566) <= a or b;
    layer4_outputs(4567) <= b;
    layer4_outputs(4568) <= a;
    layer4_outputs(4569) <= a;
    layer4_outputs(4570) <= a xor b;
    layer4_outputs(4571) <= a;
    layer4_outputs(4572) <= b;
    layer4_outputs(4573) <= not (a or b);
    layer4_outputs(4574) <= not b;
    layer4_outputs(4575) <= b;
    layer4_outputs(4576) <= not a;
    layer4_outputs(4577) <= a;
    layer4_outputs(4578) <= not (a xor b);
    layer4_outputs(4579) <= a and b;
    layer4_outputs(4580) <= not (a and b);
    layer4_outputs(4581) <= b;
    layer4_outputs(4582) <= not a;
    layer4_outputs(4583) <= b and not a;
    layer4_outputs(4584) <= a and not b;
    layer4_outputs(4585) <= not a;
    layer4_outputs(4586) <= b;
    layer4_outputs(4587) <= not a or b;
    layer4_outputs(4588) <= a xor b;
    layer4_outputs(4589) <= a or b;
    layer4_outputs(4590) <= not b;
    layer4_outputs(4591) <= a;
    layer4_outputs(4592) <= a;
    layer4_outputs(4593) <= not b or a;
    layer4_outputs(4594) <= a and b;
    layer4_outputs(4595) <= not (a xor b);
    layer4_outputs(4596) <= b;
    layer4_outputs(4597) <= a;
    layer4_outputs(4598) <= not b or a;
    layer4_outputs(4599) <= not b;
    layer4_outputs(4600) <= not (a and b);
    layer4_outputs(4601) <= b;
    layer4_outputs(4602) <= a and not b;
    layer4_outputs(4603) <= a xor b;
    layer4_outputs(4604) <= not b;
    layer4_outputs(4605) <= not (a and b);
    layer4_outputs(4606) <= not b or a;
    layer4_outputs(4607) <= not a or b;
    layer4_outputs(4608) <= not b or a;
    layer4_outputs(4609) <= b and not a;
    layer4_outputs(4610) <= not a;
    layer4_outputs(4611) <= a;
    layer4_outputs(4612) <= a xor b;
    layer4_outputs(4613) <= a or b;
    layer4_outputs(4614) <= not a or b;
    layer4_outputs(4615) <= not a or b;
    layer4_outputs(4616) <= not b or a;
    layer4_outputs(4617) <= not a or b;
    layer4_outputs(4618) <= a and not b;
    layer4_outputs(4619) <= not a or b;
    layer4_outputs(4620) <= b and not a;
    layer4_outputs(4621) <= a and b;
    layer4_outputs(4622) <= b;
    layer4_outputs(4623) <= a;
    layer4_outputs(4624) <= b;
    layer4_outputs(4625) <= not a;
    layer4_outputs(4626) <= not (a xor b);
    layer4_outputs(4627) <= not (a xor b);
    layer4_outputs(4628) <= a and not b;
    layer4_outputs(4629) <= a and not b;
    layer4_outputs(4630) <= not b or a;
    layer4_outputs(4631) <= not b;
    layer4_outputs(4632) <= not (a and b);
    layer4_outputs(4633) <= a and b;
    layer4_outputs(4634) <= not b;
    layer4_outputs(4635) <= a or b;
    layer4_outputs(4636) <= b;
    layer4_outputs(4637) <= not (a or b);
    layer4_outputs(4638) <= not b or a;
    layer4_outputs(4639) <= not a;
    layer4_outputs(4640) <= a;
    layer4_outputs(4641) <= not b;
    layer4_outputs(4642) <= a or b;
    layer4_outputs(4643) <= b;
    layer4_outputs(4644) <= not (a or b);
    layer4_outputs(4645) <= a xor b;
    layer4_outputs(4646) <= not (a or b);
    layer4_outputs(4647) <= not a or b;
    layer4_outputs(4648) <= a;
    layer4_outputs(4649) <= a xor b;
    layer4_outputs(4650) <= a xor b;
    layer4_outputs(4651) <= not a;
    layer4_outputs(4652) <= not b;
    layer4_outputs(4653) <= a xor b;
    layer4_outputs(4654) <= not (a or b);
    layer4_outputs(4655) <= a;
    layer4_outputs(4656) <= not a or b;
    layer4_outputs(4657) <= a or b;
    layer4_outputs(4658) <= a;
    layer4_outputs(4659) <= not b or a;
    layer4_outputs(4660) <= b and not a;
    layer4_outputs(4661) <= b;
    layer4_outputs(4662) <= not a;
    layer4_outputs(4663) <= not (a xor b);
    layer4_outputs(4664) <= b;
    layer4_outputs(4665) <= b and not a;
    layer4_outputs(4666) <= a;
    layer4_outputs(4667) <= a and b;
    layer4_outputs(4668) <= not b or a;
    layer4_outputs(4669) <= a or b;
    layer4_outputs(4670) <= a and b;
    layer4_outputs(4671) <= a xor b;
    layer4_outputs(4672) <= not a or b;
    layer4_outputs(4673) <= not b;
    layer4_outputs(4674) <= a and not b;
    layer4_outputs(4675) <= not b;
    layer4_outputs(4676) <= b and not a;
    layer4_outputs(4677) <= b;
    layer4_outputs(4678) <= not a;
    layer4_outputs(4679) <= b;
    layer4_outputs(4680) <= not a;
    layer4_outputs(4681) <= not a;
    layer4_outputs(4682) <= not a;
    layer4_outputs(4683) <= not a or b;
    layer4_outputs(4684) <= a;
    layer4_outputs(4685) <= not a;
    layer4_outputs(4686) <= not (a and b);
    layer4_outputs(4687) <= not a or b;
    layer4_outputs(4688) <= not b or a;
    layer4_outputs(4689) <= a and b;
    layer4_outputs(4690) <= b and not a;
    layer4_outputs(4691) <= not b;
    layer4_outputs(4692) <= not (a or b);
    layer4_outputs(4693) <= a xor b;
    layer4_outputs(4694) <= a;
    layer4_outputs(4695) <= '0';
    layer4_outputs(4696) <= not a;
    layer4_outputs(4697) <= b and not a;
    layer4_outputs(4698) <= not a;
    layer4_outputs(4699) <= not b;
    layer4_outputs(4700) <= a xor b;
    layer4_outputs(4701) <= not (a and b);
    layer4_outputs(4702) <= b and not a;
    layer4_outputs(4703) <= not (a and b);
    layer4_outputs(4704) <= not b or a;
    layer4_outputs(4705) <= not (a xor b);
    layer4_outputs(4706) <= not (a xor b);
    layer4_outputs(4707) <= not b;
    layer4_outputs(4708) <= a xor b;
    layer4_outputs(4709) <= a xor b;
    layer4_outputs(4710) <= a or b;
    layer4_outputs(4711) <= a and b;
    layer4_outputs(4712) <= not (a or b);
    layer4_outputs(4713) <= a;
    layer4_outputs(4714) <= a and not b;
    layer4_outputs(4715) <= a;
    layer4_outputs(4716) <= a and not b;
    layer4_outputs(4717) <= not b or a;
    layer4_outputs(4718) <= not (a and b);
    layer4_outputs(4719) <= not a;
    layer4_outputs(4720) <= a;
    layer4_outputs(4721) <= a and b;
    layer4_outputs(4722) <= not b;
    layer4_outputs(4723) <= a xor b;
    layer4_outputs(4724) <= not a;
    layer4_outputs(4725) <= a and b;
    layer4_outputs(4726) <= not (a and b);
    layer4_outputs(4727) <= not b or a;
    layer4_outputs(4728) <= not b;
    layer4_outputs(4729) <= a;
    layer4_outputs(4730) <= b and not a;
    layer4_outputs(4731) <= a and not b;
    layer4_outputs(4732) <= not b;
    layer4_outputs(4733) <= b;
    layer4_outputs(4734) <= b and not a;
    layer4_outputs(4735) <= not a or b;
    layer4_outputs(4736) <= b;
    layer4_outputs(4737) <= not b or a;
    layer4_outputs(4738) <= b;
    layer4_outputs(4739) <= b and not a;
    layer4_outputs(4740) <= not (a and b);
    layer4_outputs(4741) <= not a or b;
    layer4_outputs(4742) <= b;
    layer4_outputs(4743) <= a or b;
    layer4_outputs(4744) <= a;
    layer4_outputs(4745) <= a;
    layer4_outputs(4746) <= not b or a;
    layer4_outputs(4747) <= not b;
    layer4_outputs(4748) <= not b;
    layer4_outputs(4749) <= not a;
    layer4_outputs(4750) <= b and not a;
    layer4_outputs(4751) <= not a or b;
    layer4_outputs(4752) <= b;
    layer4_outputs(4753) <= not a;
    layer4_outputs(4754) <= not a;
    layer4_outputs(4755) <= not a;
    layer4_outputs(4756) <= not b or a;
    layer4_outputs(4757) <= a or b;
    layer4_outputs(4758) <= not a;
    layer4_outputs(4759) <= not b;
    layer4_outputs(4760) <= not a or b;
    layer4_outputs(4761) <= not (a or b);
    layer4_outputs(4762) <= not (a xor b);
    layer4_outputs(4763) <= a or b;
    layer4_outputs(4764) <= not (a xor b);
    layer4_outputs(4765) <= not b;
    layer4_outputs(4766) <= not b;
    layer4_outputs(4767) <= not a or b;
    layer4_outputs(4768) <= b;
    layer4_outputs(4769) <= not b;
    layer4_outputs(4770) <= b and not a;
    layer4_outputs(4771) <= b;
    layer4_outputs(4772) <= '1';
    layer4_outputs(4773) <= b;
    layer4_outputs(4774) <= not a;
    layer4_outputs(4775) <= a and b;
    layer4_outputs(4776) <= b and not a;
    layer4_outputs(4777) <= not a;
    layer4_outputs(4778) <= b;
    layer4_outputs(4779) <= not (a and b);
    layer4_outputs(4780) <= not b;
    layer4_outputs(4781) <= a xor b;
    layer4_outputs(4782) <= b;
    layer4_outputs(4783) <= a and b;
    layer4_outputs(4784) <= not (a or b);
    layer4_outputs(4785) <= a;
    layer4_outputs(4786) <= a and b;
    layer4_outputs(4787) <= a or b;
    layer4_outputs(4788) <= a;
    layer4_outputs(4789) <= b;
    layer4_outputs(4790) <= a and b;
    layer4_outputs(4791) <= not b or a;
    layer4_outputs(4792) <= b;
    layer4_outputs(4793) <= a;
    layer4_outputs(4794) <= not (a xor b);
    layer4_outputs(4795) <= a xor b;
    layer4_outputs(4796) <= b and not a;
    layer4_outputs(4797) <= not b;
    layer4_outputs(4798) <= a xor b;
    layer4_outputs(4799) <= not b;
    layer4_outputs(4800) <= a;
    layer4_outputs(4801) <= not (a or b);
    layer4_outputs(4802) <= not a;
    layer4_outputs(4803) <= not b or a;
    layer4_outputs(4804) <= not a;
    layer4_outputs(4805) <= b;
    layer4_outputs(4806) <= a;
    layer4_outputs(4807) <= a;
    layer4_outputs(4808) <= a;
    layer4_outputs(4809) <= b and not a;
    layer4_outputs(4810) <= a and not b;
    layer4_outputs(4811) <= a and b;
    layer4_outputs(4812) <= a;
    layer4_outputs(4813) <= not b;
    layer4_outputs(4814) <= not a;
    layer4_outputs(4815) <= not (a or b);
    layer4_outputs(4816) <= not (a and b);
    layer4_outputs(4817) <= not a;
    layer4_outputs(4818) <= '1';
    layer4_outputs(4819) <= not (a or b);
    layer4_outputs(4820) <= not a or b;
    layer4_outputs(4821) <= not a;
    layer4_outputs(4822) <= a or b;
    layer4_outputs(4823) <= not (a xor b);
    layer4_outputs(4824) <= not b;
    layer4_outputs(4825) <= a and b;
    layer4_outputs(4826) <= not a or b;
    layer4_outputs(4827) <= a and not b;
    layer4_outputs(4828) <= not (a xor b);
    layer4_outputs(4829) <= not a;
    layer4_outputs(4830) <= not a;
    layer4_outputs(4831) <= not (a or b);
    layer4_outputs(4832) <= not a;
    layer4_outputs(4833) <= a xor b;
    layer4_outputs(4834) <= a;
    layer4_outputs(4835) <= not a;
    layer4_outputs(4836) <= not a;
    layer4_outputs(4837) <= a or b;
    layer4_outputs(4838) <= not a;
    layer4_outputs(4839) <= not a or b;
    layer4_outputs(4840) <= b;
    layer4_outputs(4841) <= not b or a;
    layer4_outputs(4842) <= b and not a;
    layer4_outputs(4843) <= a;
    layer4_outputs(4844) <= not b;
    layer4_outputs(4845) <= not a;
    layer4_outputs(4846) <= b and not a;
    layer4_outputs(4847) <= b;
    layer4_outputs(4848) <= b;
    layer4_outputs(4849) <= not (a or b);
    layer4_outputs(4850) <= a xor b;
    layer4_outputs(4851) <= not b;
    layer4_outputs(4852) <= not b or a;
    layer4_outputs(4853) <= a;
    layer4_outputs(4854) <= not b;
    layer4_outputs(4855) <= not (a or b);
    layer4_outputs(4856) <= a and b;
    layer4_outputs(4857) <= not a;
    layer4_outputs(4858) <= b;
    layer4_outputs(4859) <= not (a xor b);
    layer4_outputs(4860) <= a;
    layer4_outputs(4861) <= a or b;
    layer4_outputs(4862) <= a and not b;
    layer4_outputs(4863) <= a or b;
    layer4_outputs(4864) <= b;
    layer4_outputs(4865) <= not a or b;
    layer4_outputs(4866) <= not (a xor b);
    layer4_outputs(4867) <= a or b;
    layer4_outputs(4868) <= not a or b;
    layer4_outputs(4869) <= a;
    layer4_outputs(4870) <= a or b;
    layer4_outputs(4871) <= a;
    layer4_outputs(4872) <= not a or b;
    layer4_outputs(4873) <= not a;
    layer4_outputs(4874) <= not b or a;
    layer4_outputs(4875) <= not (a and b);
    layer4_outputs(4876) <= a;
    layer4_outputs(4877) <= a;
    layer4_outputs(4878) <= b and not a;
    layer4_outputs(4879) <= a and b;
    layer4_outputs(4880) <= not (a xor b);
    layer4_outputs(4881) <= b and not a;
    layer4_outputs(4882) <= b;
    layer4_outputs(4883) <= a xor b;
    layer4_outputs(4884) <= a and b;
    layer4_outputs(4885) <= a xor b;
    layer4_outputs(4886) <= not b or a;
    layer4_outputs(4887) <= a xor b;
    layer4_outputs(4888) <= b and not a;
    layer4_outputs(4889) <= not a;
    layer4_outputs(4890) <= not (a and b);
    layer4_outputs(4891) <= a and not b;
    layer4_outputs(4892) <= b;
    layer4_outputs(4893) <= not (a xor b);
    layer4_outputs(4894) <= not b or a;
    layer4_outputs(4895) <= b;
    layer4_outputs(4896) <= not (a or b);
    layer4_outputs(4897) <= not a;
    layer4_outputs(4898) <= a xor b;
    layer4_outputs(4899) <= not b;
    layer4_outputs(4900) <= b;
    layer4_outputs(4901) <= a;
    layer4_outputs(4902) <= not (a xor b);
    layer4_outputs(4903) <= a;
    layer4_outputs(4904) <= not (a and b);
    layer4_outputs(4905) <= not b;
    layer4_outputs(4906) <= not (a or b);
    layer4_outputs(4907) <= not a;
    layer4_outputs(4908) <= b;
    layer4_outputs(4909) <= b and not a;
    layer4_outputs(4910) <= a and b;
    layer4_outputs(4911) <= not a or b;
    layer4_outputs(4912) <= a or b;
    layer4_outputs(4913) <= a;
    layer4_outputs(4914) <= not b;
    layer4_outputs(4915) <= not b or a;
    layer4_outputs(4916) <= a xor b;
    layer4_outputs(4917) <= not b;
    layer4_outputs(4918) <= '0';
    layer4_outputs(4919) <= not a;
    layer4_outputs(4920) <= not b;
    layer4_outputs(4921) <= a xor b;
    layer4_outputs(4922) <= not (a and b);
    layer4_outputs(4923) <= not b;
    layer4_outputs(4924) <= not b;
    layer4_outputs(4925) <= a xor b;
    layer4_outputs(4926) <= a xor b;
    layer4_outputs(4927) <= not (a or b);
    layer4_outputs(4928) <= a;
    layer4_outputs(4929) <= b;
    layer4_outputs(4930) <= b;
    layer4_outputs(4931) <= a xor b;
    layer4_outputs(4932) <= not b or a;
    layer4_outputs(4933) <= not (a and b);
    layer4_outputs(4934) <= not a;
    layer4_outputs(4935) <= a and b;
    layer4_outputs(4936) <= b;
    layer4_outputs(4937) <= a and b;
    layer4_outputs(4938) <= a;
    layer4_outputs(4939) <= b and not a;
    layer4_outputs(4940) <= b;
    layer4_outputs(4941) <= a and b;
    layer4_outputs(4942) <= b and not a;
    layer4_outputs(4943) <= a xor b;
    layer4_outputs(4944) <= a;
    layer4_outputs(4945) <= not (a or b);
    layer4_outputs(4946) <= not b;
    layer4_outputs(4947) <= a and not b;
    layer4_outputs(4948) <= not (a xor b);
    layer4_outputs(4949) <= not b;
    layer4_outputs(4950) <= not a;
    layer4_outputs(4951) <= not a or b;
    layer4_outputs(4952) <= not a;
    layer4_outputs(4953) <= not a or b;
    layer4_outputs(4954) <= a and not b;
    layer4_outputs(4955) <= a or b;
    layer4_outputs(4956) <= not (a xor b);
    layer4_outputs(4957) <= not a or b;
    layer4_outputs(4958) <= not (a and b);
    layer4_outputs(4959) <= a;
    layer4_outputs(4960) <= not (a or b);
    layer4_outputs(4961) <= b;
    layer4_outputs(4962) <= a;
    layer4_outputs(4963) <= not a;
    layer4_outputs(4964) <= not a;
    layer4_outputs(4965) <= not b;
    layer4_outputs(4966) <= not a;
    layer4_outputs(4967) <= not b;
    layer4_outputs(4968) <= a and not b;
    layer4_outputs(4969) <= not b;
    layer4_outputs(4970) <= not b or a;
    layer4_outputs(4971) <= not b or a;
    layer4_outputs(4972) <= not a or b;
    layer4_outputs(4973) <= not (a xor b);
    layer4_outputs(4974) <= a and not b;
    layer4_outputs(4975) <= b;
    layer4_outputs(4976) <= not a;
    layer4_outputs(4977) <= not b;
    layer4_outputs(4978) <= a xor b;
    layer4_outputs(4979) <= a and b;
    layer4_outputs(4980) <= not (a and b);
    layer4_outputs(4981) <= not b or a;
    layer4_outputs(4982) <= b and not a;
    layer4_outputs(4983) <= a;
    layer4_outputs(4984) <= not b;
    layer4_outputs(4985) <= a or b;
    layer4_outputs(4986) <= not b;
    layer4_outputs(4987) <= b and not a;
    layer4_outputs(4988) <= a xor b;
    layer4_outputs(4989) <= b and not a;
    layer4_outputs(4990) <= not b;
    layer4_outputs(4991) <= not a;
    layer4_outputs(4992) <= b;
    layer4_outputs(4993) <= a and not b;
    layer4_outputs(4994) <= not b;
    layer4_outputs(4995) <= a;
    layer4_outputs(4996) <= a and not b;
    layer4_outputs(4997) <= a xor b;
    layer4_outputs(4998) <= not b;
    layer4_outputs(4999) <= a or b;
    layer4_outputs(5000) <= not (a and b);
    layer4_outputs(5001) <= a;
    layer4_outputs(5002) <= not (a and b);
    layer4_outputs(5003) <= a and b;
    layer4_outputs(5004) <= a xor b;
    layer4_outputs(5005) <= not a;
    layer4_outputs(5006) <= a;
    layer4_outputs(5007) <= not a or b;
    layer4_outputs(5008) <= a and not b;
    layer4_outputs(5009) <= b;
    layer4_outputs(5010) <= a and b;
    layer4_outputs(5011) <= a and not b;
    layer4_outputs(5012) <= b and not a;
    layer4_outputs(5013) <= not a or b;
    layer4_outputs(5014) <= b and not a;
    layer4_outputs(5015) <= not b;
    layer4_outputs(5016) <= a;
    layer4_outputs(5017) <= b and not a;
    layer4_outputs(5018) <= b;
    layer4_outputs(5019) <= not a;
    layer4_outputs(5020) <= not (a xor b);
    layer4_outputs(5021) <= not (a and b);
    layer4_outputs(5022) <= a;
    layer4_outputs(5023) <= a xor b;
    layer4_outputs(5024) <= not b;
    layer4_outputs(5025) <= a or b;
    layer4_outputs(5026) <= a;
    layer4_outputs(5027) <= b;
    layer4_outputs(5028) <= b;
    layer4_outputs(5029) <= a;
    layer4_outputs(5030) <= not a or b;
    layer4_outputs(5031) <= not (a and b);
    layer4_outputs(5032) <= not a or b;
    layer4_outputs(5033) <= a xor b;
    layer4_outputs(5034) <= b;
    layer4_outputs(5035) <= not (a or b);
    layer4_outputs(5036) <= a or b;
    layer4_outputs(5037) <= b;
    layer4_outputs(5038) <= not b;
    layer4_outputs(5039) <= a;
    layer4_outputs(5040) <= not a;
    layer4_outputs(5041) <= not b or a;
    layer4_outputs(5042) <= a;
    layer4_outputs(5043) <= b;
    layer4_outputs(5044) <= not a;
    layer4_outputs(5045) <= b;
    layer4_outputs(5046) <= not (a or b);
    layer4_outputs(5047) <= a and not b;
    layer4_outputs(5048) <= b and not a;
    layer4_outputs(5049) <= a xor b;
    layer4_outputs(5050) <= b;
    layer4_outputs(5051) <= not b or a;
    layer4_outputs(5052) <= b;
    layer4_outputs(5053) <= b;
    layer4_outputs(5054) <= not a or b;
    layer4_outputs(5055) <= not a or b;
    layer4_outputs(5056) <= not (a or b);
    layer4_outputs(5057) <= a and b;
    layer4_outputs(5058) <= a and b;
    layer4_outputs(5059) <= b;
    layer4_outputs(5060) <= b and not a;
    layer4_outputs(5061) <= a;
    layer4_outputs(5062) <= a;
    layer4_outputs(5063) <= a and not b;
    layer4_outputs(5064) <= b and not a;
    layer4_outputs(5065) <= not b or a;
    layer4_outputs(5066) <= not b;
    layer4_outputs(5067) <= not a or b;
    layer4_outputs(5068) <= a;
    layer4_outputs(5069) <= not a or b;
    layer4_outputs(5070) <= a;
    layer4_outputs(5071) <= not b;
    layer4_outputs(5072) <= not b;
    layer4_outputs(5073) <= not (a xor b);
    layer4_outputs(5074) <= not a;
    layer4_outputs(5075) <= a and not b;
    layer4_outputs(5076) <= a;
    layer4_outputs(5077) <= not (a xor b);
    layer4_outputs(5078) <= not b or a;
    layer4_outputs(5079) <= a and b;
    layer4_outputs(5080) <= not a;
    layer4_outputs(5081) <= a and b;
    layer4_outputs(5082) <= a xor b;
    layer4_outputs(5083) <= a or b;
    layer4_outputs(5084) <= b;
    layer4_outputs(5085) <= b;
    layer4_outputs(5086) <= not b;
    layer4_outputs(5087) <= not b or a;
    layer4_outputs(5088) <= a or b;
    layer4_outputs(5089) <= not (a or b);
    layer4_outputs(5090) <= not (a or b);
    layer4_outputs(5091) <= not b;
    layer4_outputs(5092) <= b and not a;
    layer4_outputs(5093) <= not a;
    layer4_outputs(5094) <= not b or a;
    layer4_outputs(5095) <= not a;
    layer4_outputs(5096) <= a and not b;
    layer4_outputs(5097) <= not b;
    layer4_outputs(5098) <= not a;
    layer4_outputs(5099) <= not (a or b);
    layer4_outputs(5100) <= not b;
    layer4_outputs(5101) <= a and not b;
    layer4_outputs(5102) <= b;
    layer4_outputs(5103) <= a;
    layer4_outputs(5104) <= not b or a;
    layer4_outputs(5105) <= a;
    layer4_outputs(5106) <= not a;
    layer4_outputs(5107) <= a;
    layer4_outputs(5108) <= b;
    layer4_outputs(5109) <= b;
    layer4_outputs(5110) <= a xor b;
    layer4_outputs(5111) <= not a;
    layer4_outputs(5112) <= not a;
    layer4_outputs(5113) <= a and not b;
    layer4_outputs(5114) <= a;
    layer4_outputs(5115) <= a;
    layer4_outputs(5116) <= b;
    layer4_outputs(5117) <= a and not b;
    layer4_outputs(5118) <= not (a and b);
    layer4_outputs(5119) <= not a or b;
    outputs(0) <= b;
    outputs(1) <= not a;
    outputs(2) <= a;
    outputs(3) <= not (a xor b);
    outputs(4) <= not b;
    outputs(5) <= not (a xor b);
    outputs(6) <= not a;
    outputs(7) <= a xor b;
    outputs(8) <= not b;
    outputs(9) <= not a;
    outputs(10) <= not b;
    outputs(11) <= not b;
    outputs(12) <= not a or b;
    outputs(13) <= not a;
    outputs(14) <= a and b;
    outputs(15) <= not (a xor b);
    outputs(16) <= a;
    outputs(17) <= a and b;
    outputs(18) <= a;
    outputs(19) <= a and not b;
    outputs(20) <= not (a and b);
    outputs(21) <= a and not b;
    outputs(22) <= not a;
    outputs(23) <= not b;
    outputs(24) <= a xor b;
    outputs(25) <= not a;
    outputs(26) <= a xor b;
    outputs(27) <= a;
    outputs(28) <= not (a or b);
    outputs(29) <= b;
    outputs(30) <= b;
    outputs(31) <= not b;
    outputs(32) <= not (a or b);
    outputs(33) <= a and not b;
    outputs(34) <= a xor b;
    outputs(35) <= not b;
    outputs(36) <= not (a and b);
    outputs(37) <= a;
    outputs(38) <= not a;
    outputs(39) <= a;
    outputs(40) <= a xor b;
    outputs(41) <= a;
    outputs(42) <= a;
    outputs(43) <= b;
    outputs(44) <= not b;
    outputs(45) <= not a;
    outputs(46) <= a or b;
    outputs(47) <= not b;
    outputs(48) <= not a;
    outputs(49) <= a and b;
    outputs(50) <= a and not b;
    outputs(51) <= not a;
    outputs(52) <= not (a xor b);
    outputs(53) <= a or b;
    outputs(54) <= not (a xor b);
    outputs(55) <= b;
    outputs(56) <= not b;
    outputs(57) <= a and not b;
    outputs(58) <= not (a and b);
    outputs(59) <= not (a xor b);
    outputs(60) <= not a;
    outputs(61) <= b and not a;
    outputs(62) <= a;
    outputs(63) <= not a;
    outputs(64) <= a xor b;
    outputs(65) <= not (a or b);
    outputs(66) <= not b;
    outputs(67) <= not b;
    outputs(68) <= not (a or b);
    outputs(69) <= a and b;
    outputs(70) <= a;
    outputs(71) <= b;
    outputs(72) <= a and not b;
    outputs(73) <= a and not b;
    outputs(74) <= not b;
    outputs(75) <= not (a xor b);
    outputs(76) <= not b;
    outputs(77) <= not (a or b);
    outputs(78) <= b and not a;
    outputs(79) <= a;
    outputs(80) <= not a;
    outputs(81) <= not (a xor b);
    outputs(82) <= not (a and b);
    outputs(83) <= b and not a;
    outputs(84) <= b;
    outputs(85) <= not (a or b);
    outputs(86) <= not b;
    outputs(87) <= not b;
    outputs(88) <= not a;
    outputs(89) <= not a;
    outputs(90) <= a;
    outputs(91) <= not (a xor b);
    outputs(92) <= a xor b;
    outputs(93) <= not (a or b);
    outputs(94) <= b;
    outputs(95) <= b and not a;
    outputs(96) <= a;
    outputs(97) <= a;
    outputs(98) <= b;
    outputs(99) <= not b;
    outputs(100) <= b;
    outputs(101) <= not a;
    outputs(102) <= not (a or b);
    outputs(103) <= not b;
    outputs(104) <= b;
    outputs(105) <= b;
    outputs(106) <= not (a or b);
    outputs(107) <= b;
    outputs(108) <= not b;
    outputs(109) <= a;
    outputs(110) <= b;
    outputs(111) <= not a;
    outputs(112) <= a;
    outputs(113) <= not b;
    outputs(114) <= not b;
    outputs(115) <= a xor b;
    outputs(116) <= not b;
    outputs(117) <= a xor b;
    outputs(118) <= a;
    outputs(119) <= not (a xor b);
    outputs(120) <= not a;
    outputs(121) <= not (a or b);
    outputs(122) <= b;
    outputs(123) <= a xor b;
    outputs(124) <= b and not a;
    outputs(125) <= a;
    outputs(126) <= a and b;
    outputs(127) <= b;
    outputs(128) <= a;
    outputs(129) <= a xor b;
    outputs(130) <= not a;
    outputs(131) <= not a or b;
    outputs(132) <= a;
    outputs(133) <= a;
    outputs(134) <= a or b;
    outputs(135) <= a;
    outputs(136) <= not a;
    outputs(137) <= a;
    outputs(138) <= not (a xor b);
    outputs(139) <= a;
    outputs(140) <= not b;
    outputs(141) <= not (a or b);
    outputs(142) <= not (a xor b);
    outputs(143) <= b;
    outputs(144) <= a and not b;
    outputs(145) <= not b;
    outputs(146) <= not b;
    outputs(147) <= a;
    outputs(148) <= a and not b;
    outputs(149) <= a;
    outputs(150) <= not a;
    outputs(151) <= not b;
    outputs(152) <= b;
    outputs(153) <= b and not a;
    outputs(154) <= not b;
    outputs(155) <= a and not b;
    outputs(156) <= a and not b;
    outputs(157) <= b;
    outputs(158) <= not b;
    outputs(159) <= a;
    outputs(160) <= a;
    outputs(161) <= not (a xor b);
    outputs(162) <= b;
    outputs(163) <= not b;
    outputs(164) <= not a;
    outputs(165) <= a and not b;
    outputs(166) <= not (a xor b);
    outputs(167) <= a and not b;
    outputs(168) <= not b;
    outputs(169) <= a and not b;
    outputs(170) <= not (a or b);
    outputs(171) <= a or b;
    outputs(172) <= a xor b;
    outputs(173) <= b and not a;
    outputs(174) <= a;
    outputs(175) <= not (a or b);
    outputs(176) <= not a or b;
    outputs(177) <= a;
    outputs(178) <= b;
    outputs(179) <= not b;
    outputs(180) <= not (a xor b);
    outputs(181) <= a;
    outputs(182) <= a xor b;
    outputs(183) <= not a or b;
    outputs(184) <= b;
    outputs(185) <= not b;
    outputs(186) <= not b;
    outputs(187) <= not b;
    outputs(188) <= a xor b;
    outputs(189) <= not (a xor b);
    outputs(190) <= a;
    outputs(191) <= a and b;
    outputs(192) <= not b;
    outputs(193) <= not (a or b);
    outputs(194) <= not b or a;
    outputs(195) <= not (a or b);
    outputs(196) <= not (a xor b);
    outputs(197) <= not a or b;
    outputs(198) <= not a;
    outputs(199) <= not a;
    outputs(200) <= b;
    outputs(201) <= not b;
    outputs(202) <= not b or a;
    outputs(203) <= not (a xor b);
    outputs(204) <= a;
    outputs(205) <= not (a xor b);
    outputs(206) <= b;
    outputs(207) <= b and not a;
    outputs(208) <= b;
    outputs(209) <= a and not b;
    outputs(210) <= a;
    outputs(211) <= b;
    outputs(212) <= not a;
    outputs(213) <= not (a xor b);
    outputs(214) <= not a;
    outputs(215) <= not (a xor b);
    outputs(216) <= not b;
    outputs(217) <= a;
    outputs(218) <= not b;
    outputs(219) <= b and not a;
    outputs(220) <= not (a xor b);
    outputs(221) <= not b;
    outputs(222) <= not b;
    outputs(223) <= not (a and b);
    outputs(224) <= b;
    outputs(225) <= not (a xor b);
    outputs(226) <= a xor b;
    outputs(227) <= not a;
    outputs(228) <= a;
    outputs(229) <= a xor b;
    outputs(230) <= a xor b;
    outputs(231) <= not a;
    outputs(232) <= a and b;
    outputs(233) <= b;
    outputs(234) <= a and not b;
    outputs(235) <= not (a or b);
    outputs(236) <= a;
    outputs(237) <= b and not a;
    outputs(238) <= not b;
    outputs(239) <= not a;
    outputs(240) <= not b;
    outputs(241) <= a xor b;
    outputs(242) <= a;
    outputs(243) <= a;
    outputs(244) <= not b;
    outputs(245) <= not b;
    outputs(246) <= not b;
    outputs(247) <= not a;
    outputs(248) <= b;
    outputs(249) <= not b;
    outputs(250) <= not b;
    outputs(251) <= a xor b;
    outputs(252) <= b;
    outputs(253) <= b;
    outputs(254) <= a and not b;
    outputs(255) <= b and not a;
    outputs(256) <= not b;
    outputs(257) <= a;
    outputs(258) <= not a;
    outputs(259) <= b and not a;
    outputs(260) <= not b or a;
    outputs(261) <= not (a xor b);
    outputs(262) <= not a;
    outputs(263) <= a and b;
    outputs(264) <= not a;
    outputs(265) <= not (a or b);
    outputs(266) <= not (a or b);
    outputs(267) <= not b;
    outputs(268) <= a and b;
    outputs(269) <= not b;
    outputs(270) <= b and not a;
    outputs(271) <= a or b;
    outputs(272) <= not a;
    outputs(273) <= not a;
    outputs(274) <= not (a and b);
    outputs(275) <= b;
    outputs(276) <= b;
    outputs(277) <= a and b;
    outputs(278) <= b and not a;
    outputs(279) <= not b;
    outputs(280) <= a and b;
    outputs(281) <= not (a xor b);
    outputs(282) <= a and not b;
    outputs(283) <= b;
    outputs(284) <= a and b;
    outputs(285) <= a or b;
    outputs(286) <= a and not b;
    outputs(287) <= not a;
    outputs(288) <= a;
    outputs(289) <= a xor b;
    outputs(290) <= not a;
    outputs(291) <= not a;
    outputs(292) <= b;
    outputs(293) <= a and not b;
    outputs(294) <= a;
    outputs(295) <= b;
    outputs(296) <= not (a xor b);
    outputs(297) <= not a;
    outputs(298) <= not b or a;
    outputs(299) <= not a;
    outputs(300) <= not a;
    outputs(301) <= a xor b;
    outputs(302) <= not a;
    outputs(303) <= a xor b;
    outputs(304) <= b;
    outputs(305) <= not a;
    outputs(306) <= a and b;
    outputs(307) <= not (a or b);
    outputs(308) <= a;
    outputs(309) <= not (a xor b);
    outputs(310) <= not b;
    outputs(311) <= not (a xor b);
    outputs(312) <= not (a and b);
    outputs(313) <= b;
    outputs(314) <= not b;
    outputs(315) <= a xor b;
    outputs(316) <= a and not b;
    outputs(317) <= not a;
    outputs(318) <= a xor b;
    outputs(319) <= not a;
    outputs(320) <= not b;
    outputs(321) <= a xor b;
    outputs(322) <= a;
    outputs(323) <= a;
    outputs(324) <= a xor b;
    outputs(325) <= a and b;
    outputs(326) <= not b;
    outputs(327) <= not a;
    outputs(328) <= not b;
    outputs(329) <= a or b;
    outputs(330) <= a;
    outputs(331) <= not a;
    outputs(332) <= b;
    outputs(333) <= not b;
    outputs(334) <= a;
    outputs(335) <= a and not b;
    outputs(336) <= a;
    outputs(337) <= not a;
    outputs(338) <= a;
    outputs(339) <= not a;
    outputs(340) <= not (a and b);
    outputs(341) <= not a or b;
    outputs(342) <= b and not a;
    outputs(343) <= b and not a;
    outputs(344) <= not (a and b);
    outputs(345) <= not (a xor b);
    outputs(346) <= b and not a;
    outputs(347) <= a;
    outputs(348) <= not b;
    outputs(349) <= a and b;
    outputs(350) <= a or b;
    outputs(351) <= a and not b;
    outputs(352) <= not b;
    outputs(353) <= not b;
    outputs(354) <= a;
    outputs(355) <= not (a xor b);
    outputs(356) <= b;
    outputs(357) <= a;
    outputs(358) <= not b;
    outputs(359) <= a and b;
    outputs(360) <= not b;
    outputs(361) <= a and not b;
    outputs(362) <= not (a xor b);
    outputs(363) <= b;
    outputs(364) <= not (a or b);
    outputs(365) <= b;
    outputs(366) <= a xor b;
    outputs(367) <= a;
    outputs(368) <= b;
    outputs(369) <= a and not b;
    outputs(370) <= a and not b;
    outputs(371) <= a and not b;
    outputs(372) <= not b;
    outputs(373) <= not a;
    outputs(374) <= b;
    outputs(375) <= not b;
    outputs(376) <= not a;
    outputs(377) <= a and b;
    outputs(378) <= a xor b;
    outputs(379) <= a and b;
    outputs(380) <= b and not a;
    outputs(381) <= a;
    outputs(382) <= b;
    outputs(383) <= not b;
    outputs(384) <= b and not a;
    outputs(385) <= not (a or b);
    outputs(386) <= not a;
    outputs(387) <= a;
    outputs(388) <= a or b;
    outputs(389) <= not a;
    outputs(390) <= a xor b;
    outputs(391) <= b and not a;
    outputs(392) <= a xor b;
    outputs(393) <= a xor b;
    outputs(394) <= b;
    outputs(395) <= a;
    outputs(396) <= a and not b;
    outputs(397) <= b and not a;
    outputs(398) <= a xor b;
    outputs(399) <= b and not a;
    outputs(400) <= not a;
    outputs(401) <= a;
    outputs(402) <= not (a xor b);
    outputs(403) <= not (a xor b);
    outputs(404) <= a xor b;
    outputs(405) <= not b;
    outputs(406) <= a;
    outputs(407) <= not b;
    outputs(408) <= not b;
    outputs(409) <= not b or a;
    outputs(410) <= a xor b;
    outputs(411) <= b;
    outputs(412) <= b and not a;
    outputs(413) <= not a;
    outputs(414) <= not (a xor b);
    outputs(415) <= a;
    outputs(416) <= not (a xor b);
    outputs(417) <= b and not a;
    outputs(418) <= a xor b;
    outputs(419) <= not (a or b);
    outputs(420) <= b and not a;
    outputs(421) <= b;
    outputs(422) <= not (a and b);
    outputs(423) <= a and not b;
    outputs(424) <= not (a or b);
    outputs(425) <= b;
    outputs(426) <= a and b;
    outputs(427) <= a xor b;
    outputs(428) <= not b;
    outputs(429) <= a and b;
    outputs(430) <= a;
    outputs(431) <= not a;
    outputs(432) <= not a;
    outputs(433) <= a;
    outputs(434) <= not a;
    outputs(435) <= not b;
    outputs(436) <= not b;
    outputs(437) <= not b;
    outputs(438) <= a;
    outputs(439) <= a and b;
    outputs(440) <= a;
    outputs(441) <= not a;
    outputs(442) <= not a;
    outputs(443) <= not (a xor b);
    outputs(444) <= not a;
    outputs(445) <= not b or a;
    outputs(446) <= a xor b;
    outputs(447) <= not (a and b);
    outputs(448) <= a xor b;
    outputs(449) <= not b;
    outputs(450) <= not (a xor b);
    outputs(451) <= not a;
    outputs(452) <= not b;
    outputs(453) <= not (a or b);
    outputs(454) <= not b;
    outputs(455) <= a and not b;
    outputs(456) <= a;
    outputs(457) <= not b;
    outputs(458) <= a xor b;
    outputs(459) <= not b;
    outputs(460) <= not b;
    outputs(461) <= not b;
    outputs(462) <= not (a xor b);
    outputs(463) <= b;
    outputs(464) <= a and b;
    outputs(465) <= not b;
    outputs(466) <= a;
    outputs(467) <= not a;
    outputs(468) <= not b;
    outputs(469) <= not b;
    outputs(470) <= not a;
    outputs(471) <= not b;
    outputs(472) <= a and not b;
    outputs(473) <= not (a and b);
    outputs(474) <= a xor b;
    outputs(475) <= b;
    outputs(476) <= not (a xor b);
    outputs(477) <= not (a or b);
    outputs(478) <= b;
    outputs(479) <= a;
    outputs(480) <= not a;
    outputs(481) <= not b or a;
    outputs(482) <= not a or b;
    outputs(483) <= a;
    outputs(484) <= not (a or b);
    outputs(485) <= b;
    outputs(486) <= not (a and b);
    outputs(487) <= b;
    outputs(488) <= not b or a;
    outputs(489) <= b and not a;
    outputs(490) <= not b;
    outputs(491) <= not b;
    outputs(492) <= not b;
    outputs(493) <= not (a xor b);
    outputs(494) <= not a;
    outputs(495) <= a;
    outputs(496) <= not b;
    outputs(497) <= a;
    outputs(498) <= not (a xor b);
    outputs(499) <= not a;
    outputs(500) <= a;
    outputs(501) <= not b;
    outputs(502) <= b;
    outputs(503) <= a;
    outputs(504) <= a and not b;
    outputs(505) <= not (a xor b);
    outputs(506) <= not (a and b);
    outputs(507) <= b and not a;
    outputs(508) <= not a;
    outputs(509) <= b;
    outputs(510) <= not a;
    outputs(511) <= not b;
    outputs(512) <= not a;
    outputs(513) <= a and not b;
    outputs(514) <= not b;
    outputs(515) <= a and b;
    outputs(516) <= a and b;
    outputs(517) <= a xor b;
    outputs(518) <= a and b;
    outputs(519) <= a and b;
    outputs(520) <= a xor b;
    outputs(521) <= not (a or b);
    outputs(522) <= b and not a;
    outputs(523) <= not a;
    outputs(524) <= b;
    outputs(525) <= a and b;
    outputs(526) <= not a or b;
    outputs(527) <= not (a xor b);
    outputs(528) <= a and not b;
    outputs(529) <= b and not a;
    outputs(530) <= a;
    outputs(531) <= not a;
    outputs(532) <= b and not a;
    outputs(533) <= b and not a;
    outputs(534) <= a xor b;
    outputs(535) <= a and b;
    outputs(536) <= not (a or b);
    outputs(537) <= a xor b;
    outputs(538) <= a xor b;
    outputs(539) <= a and b;
    outputs(540) <= b and not a;
    outputs(541) <= not (a or b);
    outputs(542) <= a and not b;
    outputs(543) <= a and not b;
    outputs(544) <= not b;
    outputs(545) <= a and not b;
    outputs(546) <= a and b;
    outputs(547) <= b and not a;
    outputs(548) <= a;
    outputs(549) <= a;
    outputs(550) <= a and not b;
    outputs(551) <= b and not a;
    outputs(552) <= a and not b;
    outputs(553) <= a and b;
    outputs(554) <= a and not b;
    outputs(555) <= a and b;
    outputs(556) <= a;
    outputs(557) <= a xor b;
    outputs(558) <= a;
    outputs(559) <= a and b;
    outputs(560) <= not a;
    outputs(561) <= not (a or b);
    outputs(562) <= a and b;
    outputs(563) <= b;
    outputs(564) <= a and not b;
    outputs(565) <= a and b;
    outputs(566) <= b and not a;
    outputs(567) <= not b;
    outputs(568) <= a and b;
    outputs(569) <= not a;
    outputs(570) <= a and not b;
    outputs(571) <= not (a or b);
    outputs(572) <= not (a xor b);
    outputs(573) <= not a or b;
    outputs(574) <= a;
    outputs(575) <= not (a xor b);
    outputs(576) <= b and not a;
    outputs(577) <= a;
    outputs(578) <= a or b;
    outputs(579) <= b;
    outputs(580) <= a and b;
    outputs(581) <= not (a or b);
    outputs(582) <= not (a or b);
    outputs(583) <= a and b;
    outputs(584) <= a and b;
    outputs(585) <= not (a or b);
    outputs(586) <= not b;
    outputs(587) <= b;
    outputs(588) <= not (a or b);
    outputs(589) <= not (a or b);
    outputs(590) <= not b;
    outputs(591) <= a;
    outputs(592) <= not b;
    outputs(593) <= not b;
    outputs(594) <= not (a and b);
    outputs(595) <= not b;
    outputs(596) <= not b;
    outputs(597) <= not (a or b);
    outputs(598) <= a;
    outputs(599) <= a and not b;
    outputs(600) <= not a;
    outputs(601) <= b;
    outputs(602) <= not a;
    outputs(603) <= a and not b;
    outputs(604) <= not b;
    outputs(605) <= b and not a;
    outputs(606) <= b and not a;
    outputs(607) <= not a;
    outputs(608) <= a and b;
    outputs(609) <= not (a or b);
    outputs(610) <= a xor b;
    outputs(611) <= not b;
    outputs(612) <= a;
    outputs(613) <= not (a or b);
    outputs(614) <= b and not a;
    outputs(615) <= a and not b;
    outputs(616) <= a xor b;
    outputs(617) <= b and not a;
    outputs(618) <= not (a xor b);
    outputs(619) <= not (a or b);
    outputs(620) <= a and not b;
    outputs(621) <= b and not a;
    outputs(622) <= not a;
    outputs(623) <= a and not b;
    outputs(624) <= a and b;
    outputs(625) <= b and not a;
    outputs(626) <= not b;
    outputs(627) <= not (a or b);
    outputs(628) <= not a;
    outputs(629) <= a and b;
    outputs(630) <= not (a or b);
    outputs(631) <= a and not b;
    outputs(632) <= b;
    outputs(633) <= a and not b;
    outputs(634) <= not (a or b);
    outputs(635) <= a xor b;
    outputs(636) <= a and b;
    outputs(637) <= b and not a;
    outputs(638) <= not (a or b);
    outputs(639) <= not (a or b);
    outputs(640) <= a and b;
    outputs(641) <= a and not b;
    outputs(642) <= b and not a;
    outputs(643) <= not (a or b);
    outputs(644) <= b and not a;
    outputs(645) <= a;
    outputs(646) <= not (a or b);
    outputs(647) <= b and not a;
    outputs(648) <= not (a or b);
    outputs(649) <= not a;
    outputs(650) <= not b;
    outputs(651) <= not b;
    outputs(652) <= a and not b;
    outputs(653) <= b;
    outputs(654) <= a and b;
    outputs(655) <= b and not a;
    outputs(656) <= a and b;
    outputs(657) <= a and not b;
    outputs(658) <= a and not b;
    outputs(659) <= b;
    outputs(660) <= not a or b;
    outputs(661) <= a and not b;
    outputs(662) <= not a;
    outputs(663) <= not a or b;
    outputs(664) <= not b;
    outputs(665) <= not b or a;
    outputs(666) <= not a;
    outputs(667) <= not (a xor b);
    outputs(668) <= not (a or b);
    outputs(669) <= not a;
    outputs(670) <= a and not b;
    outputs(671) <= a and b;
    outputs(672) <= b;
    outputs(673) <= not (a or b);
    outputs(674) <= a;
    outputs(675) <= a and not b;
    outputs(676) <= a xor b;
    outputs(677) <= not a;
    outputs(678) <= not (a or b);
    outputs(679) <= a;
    outputs(680) <= a and not b;
    outputs(681) <= a and b;
    outputs(682) <= not (a or b);
    outputs(683) <= not b;
    outputs(684) <= not (a xor b);
    outputs(685) <= a;
    outputs(686) <= not b;
    outputs(687) <= a and not b;
    outputs(688) <= a or b;
    outputs(689) <= a;
    outputs(690) <= a;
    outputs(691) <= a;
    outputs(692) <= a xor b;
    outputs(693) <= not (a or b);
    outputs(694) <= b and not a;
    outputs(695) <= not a;
    outputs(696) <= a and b;
    outputs(697) <= b and not a;
    outputs(698) <= a xor b;
    outputs(699) <= a;
    outputs(700) <= not (a or b);
    outputs(701) <= a and b;
    outputs(702) <= a and not b;
    outputs(703) <= a;
    outputs(704) <= a xor b;
    outputs(705) <= not b;
    outputs(706) <= a;
    outputs(707) <= a and not b;
    outputs(708) <= a xor b;
    outputs(709) <= a xor b;
    outputs(710) <= b and not a;
    outputs(711) <= b;
    outputs(712) <= a and b;
    outputs(713) <= a xor b;
    outputs(714) <= a and not b;
    outputs(715) <= a and b;
    outputs(716) <= a and not b;
    outputs(717) <= not a;
    outputs(718) <= not (a or b);
    outputs(719) <= not (a or b);
    outputs(720) <= not (a or b);
    outputs(721) <= b;
    outputs(722) <= b;
    outputs(723) <= a xor b;
    outputs(724) <= a and b;
    outputs(725) <= a xor b;
    outputs(726) <= a and b;
    outputs(727) <= b;
    outputs(728) <= b and not a;
    outputs(729) <= not a;
    outputs(730) <= not (a xor b);
    outputs(731) <= b and not a;
    outputs(732) <= a and b;
    outputs(733) <= not (a xor b);
    outputs(734) <= not a;
    outputs(735) <= not a;
    outputs(736) <= a and not b;
    outputs(737) <= not (a or b);
    outputs(738) <= a or b;
    outputs(739) <= a and not b;
    outputs(740) <= a and b;
    outputs(741) <= not a;
    outputs(742) <= not a;
    outputs(743) <= not (a or b);
    outputs(744) <= not b;
    outputs(745) <= a;
    outputs(746) <= a;
    outputs(747) <= b;
    outputs(748) <= not b;
    outputs(749) <= not b;
    outputs(750) <= b and not a;
    outputs(751) <= not b;
    outputs(752) <= not a;
    outputs(753) <= b and not a;
    outputs(754) <= b and not a;
    outputs(755) <= not (a or b);
    outputs(756) <= b;
    outputs(757) <= not (a or b);
    outputs(758) <= a;
    outputs(759) <= b and not a;
    outputs(760) <= b;
    outputs(761) <= not (a or b);
    outputs(762) <= not b;
    outputs(763) <= b;
    outputs(764) <= a and b;
    outputs(765) <= a and not b;
    outputs(766) <= a xor b;
    outputs(767) <= not a or b;
    outputs(768) <= b;
    outputs(769) <= not (a or b);
    outputs(770) <= b and not a;
    outputs(771) <= a and not b;
    outputs(772) <= a xor b;
    outputs(773) <= b and not a;
    outputs(774) <= not (a or b);
    outputs(775) <= a and b;
    outputs(776) <= not (a or b);
    outputs(777) <= a;
    outputs(778) <= a and not b;
    outputs(779) <= a xor b;
    outputs(780) <= not b;
    outputs(781) <= b and not a;
    outputs(782) <= b;
    outputs(783) <= a and b;
    outputs(784) <= a and not b;
    outputs(785) <= not a or b;
    outputs(786) <= a and not b;
    outputs(787) <= a and b;
    outputs(788) <= b and not a;
    outputs(789) <= not a;
    outputs(790) <= b and not a;
    outputs(791) <= not (a or b);
    outputs(792) <= a and not b;
    outputs(793) <= a and not b;
    outputs(794) <= a and not b;
    outputs(795) <= a and b;
    outputs(796) <= a and not b;
    outputs(797) <= a and not b;
    outputs(798) <= a and b;
    outputs(799) <= not a;
    outputs(800) <= not b;
    outputs(801) <= a and b;
    outputs(802) <= not b;
    outputs(803) <= not (a xor b);
    outputs(804) <= a and b;
    outputs(805) <= a;
    outputs(806) <= b and not a;
    outputs(807) <= not (a or b);
    outputs(808) <= a and not b;
    outputs(809) <= a;
    outputs(810) <= b;
    outputs(811) <= a and not b;
    outputs(812) <= not (a or b);
    outputs(813) <= a and b;
    outputs(814) <= b and not a;
    outputs(815) <= a and not b;
    outputs(816) <= not (a xor b);
    outputs(817) <= a and b;
    outputs(818) <= not a;
    outputs(819) <= a and b;
    outputs(820) <= a and not b;
    outputs(821) <= a and not b;
    outputs(822) <= not (a or b);
    outputs(823) <= b and not a;
    outputs(824) <= not (a xor b);
    outputs(825) <= a and b;
    outputs(826) <= not (a or b);
    outputs(827) <= a and b;
    outputs(828) <= a and not b;
    outputs(829) <= not (a or b);
    outputs(830) <= a and b;
    outputs(831) <= not (a or b);
    outputs(832) <= a and not b;
    outputs(833) <= b and not a;
    outputs(834) <= a and b;
    outputs(835) <= a and b;
    outputs(836) <= not (a xor b);
    outputs(837) <= not (a xor b);
    outputs(838) <= not (a xor b);
    outputs(839) <= a and b;
    outputs(840) <= not b;
    outputs(841) <= a xor b;
    outputs(842) <= a and not b;
    outputs(843) <= b;
    outputs(844) <= a xor b;
    outputs(845) <= not (a or b);
    outputs(846) <= a xor b;
    outputs(847) <= a and not b;
    outputs(848) <= not (a or b);
    outputs(849) <= not a;
    outputs(850) <= a and not b;
    outputs(851) <= b;
    outputs(852) <= not (a or b);
    outputs(853) <= not (a or b);
    outputs(854) <= not a or b;
    outputs(855) <= a and not b;
    outputs(856) <= a and b;
    outputs(857) <= not a;
    outputs(858) <= not a;
    outputs(859) <= a and b;
    outputs(860) <= a;
    outputs(861) <= a;
    outputs(862) <= not a or b;
    outputs(863) <= a and b;
    outputs(864) <= b and not a;
    outputs(865) <= a;
    outputs(866) <= a;
    outputs(867) <= not b;
    outputs(868) <= a and not b;
    outputs(869) <= not b;
    outputs(870) <= not a;
    outputs(871) <= a and not b;
    outputs(872) <= a xor b;
    outputs(873) <= a;
    outputs(874) <= b and not a;
    outputs(875) <= a and not b;
    outputs(876) <= not b;
    outputs(877) <= a xor b;
    outputs(878) <= b and not a;
    outputs(879) <= not (a or b);
    outputs(880) <= a and b;
    outputs(881) <= not (a or b);
    outputs(882) <= a and not b;
    outputs(883) <= a and not b;
    outputs(884) <= b;
    outputs(885) <= a;
    outputs(886) <= b;
    outputs(887) <= a xor b;
    outputs(888) <= b and not a;
    outputs(889) <= not (a and b);
    outputs(890) <= b and not a;
    outputs(891) <= not (a xor b);
    outputs(892) <= not a;
    outputs(893) <= a xor b;
    outputs(894) <= not (a or b);
    outputs(895) <= a xor b;
    outputs(896) <= not (a or b);
    outputs(897) <= b;
    outputs(898) <= b and not a;
    outputs(899) <= b and not a;
    outputs(900) <= not (a xor b);
    outputs(901) <= a;
    outputs(902) <= not a;
    outputs(903) <= not (a or b);
    outputs(904) <= not (a xor b);
    outputs(905) <= not a;
    outputs(906) <= b and not a;
    outputs(907) <= b;
    outputs(908) <= b and not a;
    outputs(909) <= not (a or b);
    outputs(910) <= b and not a;
    outputs(911) <= a xor b;
    outputs(912) <= not b;
    outputs(913) <= a xor b;
    outputs(914) <= a;
    outputs(915) <= not a;
    outputs(916) <= a xor b;
    outputs(917) <= not a;
    outputs(918) <= not (a or b);
    outputs(919) <= a;
    outputs(920) <= a and not b;
    outputs(921) <= b;
    outputs(922) <= not (a or b);
    outputs(923) <= a and not b;
    outputs(924) <= not (a or b);
    outputs(925) <= a and b;
    outputs(926) <= a and not b;
    outputs(927) <= b and not a;
    outputs(928) <= a xor b;
    outputs(929) <= b;
    outputs(930) <= not (a or b);
    outputs(931) <= not (a xor b);
    outputs(932) <= not (a xor b);
    outputs(933) <= a and not b;
    outputs(934) <= b and not a;
    outputs(935) <= not (a or b);
    outputs(936) <= a and not b;
    outputs(937) <= b;
    outputs(938) <= not b;
    outputs(939) <= a and b;
    outputs(940) <= not (a or b);
    outputs(941) <= not (a or b);
    outputs(942) <= not a;
    outputs(943) <= not a or b;
    outputs(944) <= a xor b;
    outputs(945) <= b;
    outputs(946) <= not b or a;
    outputs(947) <= b and not a;
    outputs(948) <= not b;
    outputs(949) <= b and not a;
    outputs(950) <= not b;
    outputs(951) <= not (a or b);
    outputs(952) <= a and b;
    outputs(953) <= a;
    outputs(954) <= a and not b;
    outputs(955) <= a and b;
    outputs(956) <= a and not b;
    outputs(957) <= a;
    outputs(958) <= a xor b;
    outputs(959) <= a and b;
    outputs(960) <= a or b;
    outputs(961) <= not a;
    outputs(962) <= a and not b;
    outputs(963) <= not (a or b);
    outputs(964) <= a and not b;
    outputs(965) <= a and not b;
    outputs(966) <= not (a or b);
    outputs(967) <= a and b;
    outputs(968) <= a and not b;
    outputs(969) <= b and not a;
    outputs(970) <= not (a or b);
    outputs(971) <= a and b;
    outputs(972) <= '0';
    outputs(973) <= a and b;
    outputs(974) <= not (a or b);
    outputs(975) <= a and not b;
    outputs(976) <= a xor b;
    outputs(977) <= a and not b;
    outputs(978) <= a and not b;
    outputs(979) <= not b;
    outputs(980) <= b;
    outputs(981) <= a and not b;
    outputs(982) <= a and not b;
    outputs(983) <= b;
    outputs(984) <= a and b;
    outputs(985) <= b and not a;
    outputs(986) <= not (a xor b);
    outputs(987) <= not (a or b);
    outputs(988) <= a;
    outputs(989) <= not a;
    outputs(990) <= not (a and b);
    outputs(991) <= b and not a;
    outputs(992) <= b;
    outputs(993) <= b and not a;
    outputs(994) <= not b;
    outputs(995) <= not a;
    outputs(996) <= b;
    outputs(997) <= not b or a;
    outputs(998) <= not (a or b);
    outputs(999) <= not a;
    outputs(1000) <= b;
    outputs(1001) <= not (a or b);
    outputs(1002) <= not (a or b);
    outputs(1003) <= b;
    outputs(1004) <= a;
    outputs(1005) <= not (a or b);
    outputs(1006) <= a and not b;
    outputs(1007) <= a xor b;
    outputs(1008) <= not a;
    outputs(1009) <= a and b;
    outputs(1010) <= a and b;
    outputs(1011) <= not (a or b);
    outputs(1012) <= a and not b;
    outputs(1013) <= a and b;
    outputs(1014) <= a and b;
    outputs(1015) <= not (a xor b);
    outputs(1016) <= a xor b;
    outputs(1017) <= not (a or b);
    outputs(1018) <= b and not a;
    outputs(1019) <= a and not b;
    outputs(1020) <= b and not a;
    outputs(1021) <= a;
    outputs(1022) <= a xor b;
    outputs(1023) <= not b;
    outputs(1024) <= not (a or b);
    outputs(1025) <= not (a or b);
    outputs(1026) <= not (a xor b);
    outputs(1027) <= a;
    outputs(1028) <= b;
    outputs(1029) <= not a;
    outputs(1030) <= not (a and b);
    outputs(1031) <= not (a xor b);
    outputs(1032) <= not b or a;
    outputs(1033) <= not (a xor b);
    outputs(1034) <= not b;
    outputs(1035) <= b and not a;
    outputs(1036) <= not (a xor b);
    outputs(1037) <= not (a xor b);
    outputs(1038) <= a xor b;
    outputs(1039) <= b;
    outputs(1040) <= not b or a;
    outputs(1041) <= not b or a;
    outputs(1042) <= a and not b;
    outputs(1043) <= not (a and b);
    outputs(1044) <= not a or b;
    outputs(1045) <= b;
    outputs(1046) <= a xor b;
    outputs(1047) <= not a;
    outputs(1048) <= b;
    outputs(1049) <= not b;
    outputs(1050) <= b and not a;
    outputs(1051) <= a xor b;
    outputs(1052) <= a;
    outputs(1053) <= not b;
    outputs(1054) <= not b;
    outputs(1055) <= not b;
    outputs(1056) <= a and not b;
    outputs(1057) <= not (a or b);
    outputs(1058) <= b;
    outputs(1059) <= b and not a;
    outputs(1060) <= a or b;
    outputs(1061) <= not b;
    outputs(1062) <= a xor b;
    outputs(1063) <= not a;
    outputs(1064) <= a and b;
    outputs(1065) <= not (a and b);
    outputs(1066) <= not a or b;
    outputs(1067) <= not b;
    outputs(1068) <= a;
    outputs(1069) <= not a;
    outputs(1070) <= not b;
    outputs(1071) <= a and b;
    outputs(1072) <= a xor b;
    outputs(1073) <= a or b;
    outputs(1074) <= b and not a;
    outputs(1075) <= a and not b;
    outputs(1076) <= not (a xor b);
    outputs(1077) <= not (a xor b);
    outputs(1078) <= not a;
    outputs(1079) <= a xor b;
    outputs(1080) <= not a;
    outputs(1081) <= not a or b;
    outputs(1082) <= a;
    outputs(1083) <= a or b;
    outputs(1084) <= not b;
    outputs(1085) <= a and not b;
    outputs(1086) <= a xor b;
    outputs(1087) <= not b;
    outputs(1088) <= a xor b;
    outputs(1089) <= a xor b;
    outputs(1090) <= not a;
    outputs(1091) <= a;
    outputs(1092) <= not a;
    outputs(1093) <= not a;
    outputs(1094) <= a;
    outputs(1095) <= a or b;
    outputs(1096) <= not b;
    outputs(1097) <= not a or b;
    outputs(1098) <= not a;
    outputs(1099) <= a xor b;
    outputs(1100) <= not (a or b);
    outputs(1101) <= a xor b;
    outputs(1102) <= b and not a;
    outputs(1103) <= not a;
    outputs(1104) <= not (a xor b);
    outputs(1105) <= b;
    outputs(1106) <= not a;
    outputs(1107) <= not a or b;
    outputs(1108) <= a;
    outputs(1109) <= a xor b;
    outputs(1110) <= not (a xor b);
    outputs(1111) <= b;
    outputs(1112) <= a xor b;
    outputs(1113) <= not a;
    outputs(1114) <= not b;
    outputs(1115) <= a;
    outputs(1116) <= not a;
    outputs(1117) <= not b;
    outputs(1118) <= not b or a;
    outputs(1119) <= b;
    outputs(1120) <= not b;
    outputs(1121) <= a;
    outputs(1122) <= a or b;
    outputs(1123) <= a;
    outputs(1124) <= a;
    outputs(1125) <= not (a and b);
    outputs(1126) <= not (a xor b);
    outputs(1127) <= a and b;
    outputs(1128) <= a or b;
    outputs(1129) <= a;
    outputs(1130) <= not b;
    outputs(1131) <= b;
    outputs(1132) <= b;
    outputs(1133) <= not (a xor b);
    outputs(1134) <= a;
    outputs(1135) <= a and b;
    outputs(1136) <= a and not b;
    outputs(1137) <= not (a or b);
    outputs(1138) <= not a;
    outputs(1139) <= a;
    outputs(1140) <= not b;
    outputs(1141) <= b;
    outputs(1142) <= a xor b;
    outputs(1143) <= not a;
    outputs(1144) <= b;
    outputs(1145) <= a;
    outputs(1146) <= not b;
    outputs(1147) <= a and not b;
    outputs(1148) <= b;
    outputs(1149) <= a xor b;
    outputs(1150) <= not a or b;
    outputs(1151) <= not b;
    outputs(1152) <= a and not b;
    outputs(1153) <= a and b;
    outputs(1154) <= a and not b;
    outputs(1155) <= not a;
    outputs(1156) <= not (a and b);
    outputs(1157) <= not (a and b);
    outputs(1158) <= a;
    outputs(1159) <= b;
    outputs(1160) <= b;
    outputs(1161) <= not (a or b);
    outputs(1162) <= b;
    outputs(1163) <= b;
    outputs(1164) <= b and not a;
    outputs(1165) <= a;
    outputs(1166) <= b;
    outputs(1167) <= not a;
    outputs(1168) <= not (a and b);
    outputs(1169) <= not a;
    outputs(1170) <= not (a xor b);
    outputs(1171) <= b;
    outputs(1172) <= not a or b;
    outputs(1173) <= a xor b;
    outputs(1174) <= not a;
    outputs(1175) <= not a;
    outputs(1176) <= not b or a;
    outputs(1177) <= b;
    outputs(1178) <= b and not a;
    outputs(1179) <= not (a xor b);
    outputs(1180) <= b and not a;
    outputs(1181) <= b;
    outputs(1182) <= b;
    outputs(1183) <= not b;
    outputs(1184) <= a;
    outputs(1185) <= a;
    outputs(1186) <= not a;
    outputs(1187) <= a or b;
    outputs(1188) <= not a or b;
    outputs(1189) <= not b;
    outputs(1190) <= not (a or b);
    outputs(1191) <= b;
    outputs(1192) <= not b;
    outputs(1193) <= not (a xor b);
    outputs(1194) <= a;
    outputs(1195) <= not (a and b);
    outputs(1196) <= a and not b;
    outputs(1197) <= not a;
    outputs(1198) <= a;
    outputs(1199) <= not (a or b);
    outputs(1200) <= not b;
    outputs(1201) <= not b;
    outputs(1202) <= a and not b;
    outputs(1203) <= not (a or b);
    outputs(1204) <= not b or a;
    outputs(1205) <= not b or a;
    outputs(1206) <= b;
    outputs(1207) <= a;
    outputs(1208) <= not (a xor b);
    outputs(1209) <= not a or b;
    outputs(1210) <= not (a or b);
    outputs(1211) <= not b;
    outputs(1212) <= a or b;
    outputs(1213) <= b;
    outputs(1214) <= a and not b;
    outputs(1215) <= not a or b;
    outputs(1216) <= not a;
    outputs(1217) <= not b;
    outputs(1218) <= b;
    outputs(1219) <= not (a xor b);
    outputs(1220) <= b and not a;
    outputs(1221) <= a and b;
    outputs(1222) <= not (a xor b);
    outputs(1223) <= a xor b;
    outputs(1224) <= a and not b;
    outputs(1225) <= b;
    outputs(1226) <= b;
    outputs(1227) <= a and not b;
    outputs(1228) <= not b or a;
    outputs(1229) <= a;
    outputs(1230) <= b;
    outputs(1231) <= b;
    outputs(1232) <= not (a or b);
    outputs(1233) <= not b;
    outputs(1234) <= not (a xor b);
    outputs(1235) <= a xor b;
    outputs(1236) <= b and not a;
    outputs(1237) <= b;
    outputs(1238) <= not a or b;
    outputs(1239) <= a and b;
    outputs(1240) <= not b;
    outputs(1241) <= a and not b;
    outputs(1242) <= a xor b;
    outputs(1243) <= a;
    outputs(1244) <= not a;
    outputs(1245) <= a xor b;
    outputs(1246) <= a;
    outputs(1247) <= b and not a;
    outputs(1248) <= not a;
    outputs(1249) <= not b;
    outputs(1250) <= not (a and b);
    outputs(1251) <= not (a or b);
    outputs(1252) <= a and b;
    outputs(1253) <= b;
    outputs(1254) <= not (a xor b);
    outputs(1255) <= not b or a;
    outputs(1256) <= a xor b;
    outputs(1257) <= not b;
    outputs(1258) <= not b;
    outputs(1259) <= not (a or b);
    outputs(1260) <= b and not a;
    outputs(1261) <= not (a xor b);
    outputs(1262) <= a and not b;
    outputs(1263) <= b;
    outputs(1264) <= not a;
    outputs(1265) <= not b;
    outputs(1266) <= not b;
    outputs(1267) <= a xor b;
    outputs(1268) <= b and not a;
    outputs(1269) <= a and b;
    outputs(1270) <= b and not a;
    outputs(1271) <= a and b;
    outputs(1272) <= not b or a;
    outputs(1273) <= a;
    outputs(1274) <= not b;
    outputs(1275) <= a and b;
    outputs(1276) <= a and b;
    outputs(1277) <= not b;
    outputs(1278) <= not (a and b);
    outputs(1279) <= a;
    outputs(1280) <= a xor b;
    outputs(1281) <= a or b;
    outputs(1282) <= a xor b;
    outputs(1283) <= a;
    outputs(1284) <= not (a xor b);
    outputs(1285) <= b and not a;
    outputs(1286) <= a xor b;
    outputs(1287) <= b;
    outputs(1288) <= not b;
    outputs(1289) <= not b;
    outputs(1290) <= not b;
    outputs(1291) <= b;
    outputs(1292) <= a;
    outputs(1293) <= not (a xor b);
    outputs(1294) <= not (a xor b);
    outputs(1295) <= b;
    outputs(1296) <= a and not b;
    outputs(1297) <= not b;
    outputs(1298) <= not a;
    outputs(1299) <= b;
    outputs(1300) <= not a;
    outputs(1301) <= not a;
    outputs(1302) <= a;
    outputs(1303) <= a;
    outputs(1304) <= a;
    outputs(1305) <= a and not b;
    outputs(1306) <= not (a xor b);
    outputs(1307) <= not b;
    outputs(1308) <= not b or a;
    outputs(1309) <= a;
    outputs(1310) <= a xor b;
    outputs(1311) <= not a;
    outputs(1312) <= a;
    outputs(1313) <= a or b;
    outputs(1314) <= not a;
    outputs(1315) <= b;
    outputs(1316) <= not b;
    outputs(1317) <= b;
    outputs(1318) <= not (a or b);
    outputs(1319) <= not a;
    outputs(1320) <= b and not a;
    outputs(1321) <= not b or a;
    outputs(1322) <= not b;
    outputs(1323) <= b;
    outputs(1324) <= not b;
    outputs(1325) <= a xor b;
    outputs(1326) <= b and not a;
    outputs(1327) <= not (a xor b);
    outputs(1328) <= not b or a;
    outputs(1329) <= not b;
    outputs(1330) <= b and not a;
    outputs(1331) <= not b or a;
    outputs(1332) <= not (a xor b);
    outputs(1333) <= a;
    outputs(1334) <= a and b;
    outputs(1335) <= a and b;
    outputs(1336) <= b;
    outputs(1337) <= a;
    outputs(1338) <= a;
    outputs(1339) <= a xor b;
    outputs(1340) <= not a or b;
    outputs(1341) <= a and b;
    outputs(1342) <= not a or b;
    outputs(1343) <= b and not a;
    outputs(1344) <= b;
    outputs(1345) <= b and not a;
    outputs(1346) <= not (a xor b);
    outputs(1347) <= b and not a;
    outputs(1348) <= not (a xor b);
    outputs(1349) <= a xor b;
    outputs(1350) <= not (a or b);
    outputs(1351) <= not a;
    outputs(1352) <= a and not b;
    outputs(1353) <= not a or b;
    outputs(1354) <= a or b;
    outputs(1355) <= a and not b;
    outputs(1356) <= a xor b;
    outputs(1357) <= not (a or b);
    outputs(1358) <= not (a or b);
    outputs(1359) <= not (a xor b);
    outputs(1360) <= a xor b;
    outputs(1361) <= not (a or b);
    outputs(1362) <= not b or a;
    outputs(1363) <= a;
    outputs(1364) <= not b;
    outputs(1365) <= a xor b;
    outputs(1366) <= not b;
    outputs(1367) <= b;
    outputs(1368) <= a;
    outputs(1369) <= not a or b;
    outputs(1370) <= not (a and b);
    outputs(1371) <= not a;
    outputs(1372) <= not (a and b);
    outputs(1373) <= not b;
    outputs(1374) <= not a;
    outputs(1375) <= not b;
    outputs(1376) <= not (a xor b);
    outputs(1377) <= not a;
    outputs(1378) <= a or b;
    outputs(1379) <= not b;
    outputs(1380) <= a or b;
    outputs(1381) <= a and b;
    outputs(1382) <= not b;
    outputs(1383) <= a;
    outputs(1384) <= b;
    outputs(1385) <= a xor b;
    outputs(1386) <= not b;
    outputs(1387) <= not b;
    outputs(1388) <= a xor b;
    outputs(1389) <= not b;
    outputs(1390) <= b and not a;
    outputs(1391) <= not (a or b);
    outputs(1392) <= a and not b;
    outputs(1393) <= b;
    outputs(1394) <= a and b;
    outputs(1395) <= not (a xor b);
    outputs(1396) <= not a;
    outputs(1397) <= not a or b;
    outputs(1398) <= a xor b;
    outputs(1399) <= not (a xor b);
    outputs(1400) <= not b;
    outputs(1401) <= b;
    outputs(1402) <= b;
    outputs(1403) <= a and b;
    outputs(1404) <= b;
    outputs(1405) <= b;
    outputs(1406) <= not a;
    outputs(1407) <= b;
    outputs(1408) <= not b or a;
    outputs(1409) <= a;
    outputs(1410) <= a xor b;
    outputs(1411) <= a;
    outputs(1412) <= a;
    outputs(1413) <= not (a xor b);
    outputs(1414) <= b and not a;
    outputs(1415) <= a and b;
    outputs(1416) <= b;
    outputs(1417) <= a and not b;
    outputs(1418) <= b and not a;
    outputs(1419) <= b;
    outputs(1420) <= a xor b;
    outputs(1421) <= a xor b;
    outputs(1422) <= not b;
    outputs(1423) <= not a;
    outputs(1424) <= a and not b;
    outputs(1425) <= a xor b;
    outputs(1426) <= not b;
    outputs(1427) <= not (a and b);
    outputs(1428) <= a or b;
    outputs(1429) <= not (a or b);
    outputs(1430) <= b;
    outputs(1431) <= b and not a;
    outputs(1432) <= not (a xor b);
    outputs(1433) <= not (a xor b);
    outputs(1434) <= b;
    outputs(1435) <= not a or b;
    outputs(1436) <= not a;
    outputs(1437) <= a;
    outputs(1438) <= a and not b;
    outputs(1439) <= not b;
    outputs(1440) <= b;
    outputs(1441) <= not b;
    outputs(1442) <= not (a xor b);
    outputs(1443) <= b and not a;
    outputs(1444) <= a xor b;
    outputs(1445) <= not a;
    outputs(1446) <= a;
    outputs(1447) <= not b or a;
    outputs(1448) <= a and b;
    outputs(1449) <= not (a xor b);
    outputs(1450) <= not (a or b);
    outputs(1451) <= not (a and b);
    outputs(1452) <= a xor b;
    outputs(1453) <= a and b;
    outputs(1454) <= a xor b;
    outputs(1455) <= a and not b;
    outputs(1456) <= a xor b;
    outputs(1457) <= not b;
    outputs(1458) <= not a;
    outputs(1459) <= a;
    outputs(1460) <= b;
    outputs(1461) <= b;
    outputs(1462) <= not b or a;
    outputs(1463) <= b;
    outputs(1464) <= not a or b;
    outputs(1465) <= a;
    outputs(1466) <= not a;
    outputs(1467) <= not b;
    outputs(1468) <= b;
    outputs(1469) <= not b;
    outputs(1470) <= not (a xor b);
    outputs(1471) <= not a or b;
    outputs(1472) <= b and not a;
    outputs(1473) <= a or b;
    outputs(1474) <= a and not b;
    outputs(1475) <= not a;
    outputs(1476) <= a or b;
    outputs(1477) <= not (a xor b);
    outputs(1478) <= not a;
    outputs(1479) <= b;
    outputs(1480) <= b;
    outputs(1481) <= b;
    outputs(1482) <= a;
    outputs(1483) <= not (a or b);
    outputs(1484) <= not (a and b);
    outputs(1485) <= a or b;
    outputs(1486) <= not (a xor b);
    outputs(1487) <= not (a xor b);
    outputs(1488) <= not b;
    outputs(1489) <= not b;
    outputs(1490) <= a;
    outputs(1491) <= not (a xor b);
    outputs(1492) <= not b;
    outputs(1493) <= b and not a;
    outputs(1494) <= a xor b;
    outputs(1495) <= a;
    outputs(1496) <= a;
    outputs(1497) <= not (a xor b);
    outputs(1498) <= not a;
    outputs(1499) <= not b;
    outputs(1500) <= not (a xor b);
    outputs(1501) <= a or b;
    outputs(1502) <= not b;
    outputs(1503) <= not b;
    outputs(1504) <= not b or a;
    outputs(1505) <= a or b;
    outputs(1506) <= not (a and b);
    outputs(1507) <= not b;
    outputs(1508) <= not (a or b);
    outputs(1509) <= a and not b;
    outputs(1510) <= b;
    outputs(1511) <= a xor b;
    outputs(1512) <= a;
    outputs(1513) <= b;
    outputs(1514) <= a xor b;
    outputs(1515) <= a;
    outputs(1516) <= a;
    outputs(1517) <= b;
    outputs(1518) <= not a;
    outputs(1519) <= not b or a;
    outputs(1520) <= a and not b;
    outputs(1521) <= a and not b;
    outputs(1522) <= not (a or b);
    outputs(1523) <= a and not b;
    outputs(1524) <= a xor b;
    outputs(1525) <= a;
    outputs(1526) <= not b;
    outputs(1527) <= a;
    outputs(1528) <= a xor b;
    outputs(1529) <= not (a xor b);
    outputs(1530) <= a and not b;
    outputs(1531) <= a and b;
    outputs(1532) <= a;
    outputs(1533) <= not a;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= a;
    outputs(1536) <= a xor b;
    outputs(1537) <= not (a xor b);
    outputs(1538) <= a and not b;
    outputs(1539) <= not a;
    outputs(1540) <= a;
    outputs(1541) <= a and b;
    outputs(1542) <= b;
    outputs(1543) <= a;
    outputs(1544) <= not b;
    outputs(1545) <= not (a or b);
    outputs(1546) <= not a;
    outputs(1547) <= not a or b;
    outputs(1548) <= not b;
    outputs(1549) <= not (a or b);
    outputs(1550) <= b and not a;
    outputs(1551) <= a and not b;
    outputs(1552) <= a and b;
    outputs(1553) <= a;
    outputs(1554) <= not b;
    outputs(1555) <= not a;
    outputs(1556) <= b;
    outputs(1557) <= not b;
    outputs(1558) <= not b;
    outputs(1559) <= a;
    outputs(1560) <= not (a xor b);
    outputs(1561) <= a;
    outputs(1562) <= not (a xor b);
    outputs(1563) <= a and not b;
    outputs(1564) <= not a;
    outputs(1565) <= a or b;
    outputs(1566) <= not a or b;
    outputs(1567) <= not b;
    outputs(1568) <= not (a xor b);
    outputs(1569) <= a xor b;
    outputs(1570) <= b;
    outputs(1571) <= not (a and b);
    outputs(1572) <= a or b;
    outputs(1573) <= a or b;
    outputs(1574) <= not a;
    outputs(1575) <= a;
    outputs(1576) <= not b;
    outputs(1577) <= a and not b;
    outputs(1578) <= a xor b;
    outputs(1579) <= a or b;
    outputs(1580) <= not a;
    outputs(1581) <= a xor b;
    outputs(1582) <= a and not b;
    outputs(1583) <= not (a or b);
    outputs(1584) <= not (a xor b);
    outputs(1585) <= not b or a;
    outputs(1586) <= a and not b;
    outputs(1587) <= b;
    outputs(1588) <= a and b;
    outputs(1589) <= a xor b;
    outputs(1590) <= b;
    outputs(1591) <= a;
    outputs(1592) <= a and not b;
    outputs(1593) <= a and not b;
    outputs(1594) <= b and not a;
    outputs(1595) <= a xor b;
    outputs(1596) <= not b;
    outputs(1597) <= not (a xor b);
    outputs(1598) <= not (a xor b);
    outputs(1599) <= a;
    outputs(1600) <= b;
    outputs(1601) <= not a;
    outputs(1602) <= a and not b;
    outputs(1603) <= b and not a;
    outputs(1604) <= not a;
    outputs(1605) <= b;
    outputs(1606) <= a;
    outputs(1607) <= a;
    outputs(1608) <= not b or a;
    outputs(1609) <= not (a and b);
    outputs(1610) <= not (a xor b);
    outputs(1611) <= a;
    outputs(1612) <= not a;
    outputs(1613) <= b;
    outputs(1614) <= not a;
    outputs(1615) <= not b;
    outputs(1616) <= not (a xor b);
    outputs(1617) <= not a;
    outputs(1618) <= b and not a;
    outputs(1619) <= a and b;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= b and not a;
    outputs(1622) <= not (a xor b);
    outputs(1623) <= not a;
    outputs(1624) <= a and b;
    outputs(1625) <= not (a xor b);
    outputs(1626) <= not a;
    outputs(1627) <= not (a or b);
    outputs(1628) <= not b;
    outputs(1629) <= not b;
    outputs(1630) <= not b or a;
    outputs(1631) <= b;
    outputs(1632) <= not b;
    outputs(1633) <= not b or a;
    outputs(1634) <= not b;
    outputs(1635) <= a and not b;
    outputs(1636) <= not (a or b);
    outputs(1637) <= a;
    outputs(1638) <= not b;
    outputs(1639) <= b and not a;
    outputs(1640) <= a xor b;
    outputs(1641) <= not b;
    outputs(1642) <= not (a xor b);
    outputs(1643) <= not (a or b);
    outputs(1644) <= a and b;
    outputs(1645) <= not (a or b);
    outputs(1646) <= b and not a;
    outputs(1647) <= b;
    outputs(1648) <= b;
    outputs(1649) <= a and b;
    outputs(1650) <= not (a xor b);
    outputs(1651) <= a;
    outputs(1652) <= a and not b;
    outputs(1653) <= a;
    outputs(1654) <= not b;
    outputs(1655) <= a and not b;
    outputs(1656) <= b;
    outputs(1657) <= a and b;
    outputs(1658) <= not a;
    outputs(1659) <= not (a and b);
    outputs(1660) <= a xor b;
    outputs(1661) <= a;
    outputs(1662) <= b;
    outputs(1663) <= a;
    outputs(1664) <= not a;
    outputs(1665) <= b and not a;
    outputs(1666) <= not a;
    outputs(1667) <= not a;
    outputs(1668) <= not b or a;
    outputs(1669) <= not b;
    outputs(1670) <= not b;
    outputs(1671) <= not (a xor b);
    outputs(1672) <= a xor b;
    outputs(1673) <= a;
    outputs(1674) <= not b or a;
    outputs(1675) <= not (a or b);
    outputs(1676) <= a;
    outputs(1677) <= not b or a;
    outputs(1678) <= not (a or b);
    outputs(1679) <= not (a xor b);
    outputs(1680) <= a;
    outputs(1681) <= not a;
    outputs(1682) <= a and not b;
    outputs(1683) <= not (a xor b);
    outputs(1684) <= a and not b;
    outputs(1685) <= a and not b;
    outputs(1686) <= b and not a;
    outputs(1687) <= not a;
    outputs(1688) <= a;
    outputs(1689) <= a;
    outputs(1690) <= not (a xor b);
    outputs(1691) <= a xor b;
    outputs(1692) <= not a;
    outputs(1693) <= not (a or b);
    outputs(1694) <= not a;
    outputs(1695) <= b;
    outputs(1696) <= not (a or b);
    outputs(1697) <= a xor b;
    outputs(1698) <= b;
    outputs(1699) <= a;
    outputs(1700) <= b;
    outputs(1701) <= a and b;
    outputs(1702) <= not a;
    outputs(1703) <= not a;
    outputs(1704) <= b;
    outputs(1705) <= a;
    outputs(1706) <= a and not b;
    outputs(1707) <= a or b;
    outputs(1708) <= not (a or b);
    outputs(1709) <= not b;
    outputs(1710) <= not a;
    outputs(1711) <= not b;
    outputs(1712) <= not b;
    outputs(1713) <= a xor b;
    outputs(1714) <= a and not b;
    outputs(1715) <= a;
    outputs(1716) <= not (a or b);
    outputs(1717) <= b;
    outputs(1718) <= a and not b;
    outputs(1719) <= a and not b;
    outputs(1720) <= not (a xor b);
    outputs(1721) <= not (a xor b);
    outputs(1722) <= not (a xor b);
    outputs(1723) <= not b;
    outputs(1724) <= not a;
    outputs(1725) <= not (a xor b);
    outputs(1726) <= not (a xor b);
    outputs(1727) <= not b or a;
    outputs(1728) <= not b;
    outputs(1729) <= not a;
    outputs(1730) <= b;
    outputs(1731) <= a and b;
    outputs(1732) <= not b;
    outputs(1733) <= a and b;
    outputs(1734) <= b;
    outputs(1735) <= a and not b;
    outputs(1736) <= a;
    outputs(1737) <= not a;
    outputs(1738) <= b;
    outputs(1739) <= not b;
    outputs(1740) <= a and not b;
    outputs(1741) <= a xor b;
    outputs(1742) <= not a;
    outputs(1743) <= a or b;
    outputs(1744) <= a and b;
    outputs(1745) <= not a;
    outputs(1746) <= a xor b;
    outputs(1747) <= b;
    outputs(1748) <= not b;
    outputs(1749) <= not a;
    outputs(1750) <= b and not a;
    outputs(1751) <= b;
    outputs(1752) <= not (a or b);
    outputs(1753) <= a and b;
    outputs(1754) <= not a;
    outputs(1755) <= not (a xor b);
    outputs(1756) <= not (a and b);
    outputs(1757) <= not b;
    outputs(1758) <= not a;
    outputs(1759) <= not a;
    outputs(1760) <= a;
    outputs(1761) <= not a;
    outputs(1762) <= b;
    outputs(1763) <= a;
    outputs(1764) <= not a;
    outputs(1765) <= not b;
    outputs(1766) <= a;
    outputs(1767) <= b;
    outputs(1768) <= b;
    outputs(1769) <= not (a and b);
    outputs(1770) <= a;
    outputs(1771) <= not b or a;
    outputs(1772) <= not (a or b);
    outputs(1773) <= a and b;
    outputs(1774) <= not b;
    outputs(1775) <= not (a xor b);
    outputs(1776) <= not (a and b);
    outputs(1777) <= a xor b;
    outputs(1778) <= a and b;
    outputs(1779) <= not (a xor b);
    outputs(1780) <= not b;
    outputs(1781) <= not a or b;
    outputs(1782) <= not b;
    outputs(1783) <= a;
    outputs(1784) <= b;
    outputs(1785) <= a;
    outputs(1786) <= a and not b;
    outputs(1787) <= a;
    outputs(1788) <= not a;
    outputs(1789) <= not a;
    outputs(1790) <= b and not a;
    outputs(1791) <= a xor b;
    outputs(1792) <= b;
    outputs(1793) <= b;
    outputs(1794) <= b and not a;
    outputs(1795) <= a and not b;
    outputs(1796) <= a and b;
    outputs(1797) <= not (a xor b);
    outputs(1798) <= not b;
    outputs(1799) <= a or b;
    outputs(1800) <= a;
    outputs(1801) <= not (a xor b);
    outputs(1802) <= a and b;
    outputs(1803) <= a;
    outputs(1804) <= a or b;
    outputs(1805) <= a or b;
    outputs(1806) <= not a;
    outputs(1807) <= not a;
    outputs(1808) <= not (a xor b);
    outputs(1809) <= b;
    outputs(1810) <= a and b;
    outputs(1811) <= a and b;
    outputs(1812) <= a;
    outputs(1813) <= not (a xor b);
    outputs(1814) <= not b;
    outputs(1815) <= a;
    outputs(1816) <= a and not b;
    outputs(1817) <= not b;
    outputs(1818) <= a;
    outputs(1819) <= not b;
    outputs(1820) <= not b;
    outputs(1821) <= not a;
    outputs(1822) <= a;
    outputs(1823) <= not (a or b);
    outputs(1824) <= a or b;
    outputs(1825) <= not b;
    outputs(1826) <= not b or a;
    outputs(1827) <= b;
    outputs(1828) <= not b;
    outputs(1829) <= not b or a;
    outputs(1830) <= b and not a;
    outputs(1831) <= a xor b;
    outputs(1832) <= b and not a;
    outputs(1833) <= not a;
    outputs(1834) <= a;
    outputs(1835) <= a and b;
    outputs(1836) <= a or b;
    outputs(1837) <= a and not b;
    outputs(1838) <= not (a and b);
    outputs(1839) <= a;
    outputs(1840) <= a and not b;
    outputs(1841) <= b and not a;
    outputs(1842) <= not b;
    outputs(1843) <= not a;
    outputs(1844) <= not (a xor b);
    outputs(1845) <= not a;
    outputs(1846) <= b;
    outputs(1847) <= a xor b;
    outputs(1848) <= b;
    outputs(1849) <= not b or a;
    outputs(1850) <= b and not a;
    outputs(1851) <= a and not b;
    outputs(1852) <= not b or a;
    outputs(1853) <= a or b;
    outputs(1854) <= not a or b;
    outputs(1855) <= not (a xor b);
    outputs(1856) <= not a;
    outputs(1857) <= not (a or b);
    outputs(1858) <= not (a or b);
    outputs(1859) <= a xor b;
    outputs(1860) <= a and b;
    outputs(1861) <= not a;
    outputs(1862) <= not b;
    outputs(1863) <= a;
    outputs(1864) <= b and not a;
    outputs(1865) <= not (a or b);
    outputs(1866) <= b and not a;
    outputs(1867) <= a;
    outputs(1868) <= b and not a;
    outputs(1869) <= a;
    outputs(1870) <= not a or b;
    outputs(1871) <= not (a xor b);
    outputs(1872) <= a or b;
    outputs(1873) <= a;
    outputs(1874) <= b;
    outputs(1875) <= not (a and b);
    outputs(1876) <= b;
    outputs(1877) <= not (a or b);
    outputs(1878) <= a xor b;
    outputs(1879) <= a and not b;
    outputs(1880) <= b;
    outputs(1881) <= not (a and b);
    outputs(1882) <= not (a xor b);
    outputs(1883) <= a and not b;
    outputs(1884) <= a;
    outputs(1885) <= a;
    outputs(1886) <= a or b;
    outputs(1887) <= a xor b;
    outputs(1888) <= b;
    outputs(1889) <= a;
    outputs(1890) <= not a;
    outputs(1891) <= a;
    outputs(1892) <= b;
    outputs(1893) <= not b;
    outputs(1894) <= b;
    outputs(1895) <= b;
    outputs(1896) <= a;
    outputs(1897) <= a and not b;
    outputs(1898) <= a;
    outputs(1899) <= a;
    outputs(1900) <= not (a xor b);
    outputs(1901) <= a and b;
    outputs(1902) <= a xor b;
    outputs(1903) <= a;
    outputs(1904) <= not (a xor b);
    outputs(1905) <= not b or a;
    outputs(1906) <= not a;
    outputs(1907) <= not a;
    outputs(1908) <= not b;
    outputs(1909) <= a xor b;
    outputs(1910) <= not (a xor b);
    outputs(1911) <= not (a or b);
    outputs(1912) <= a;
    outputs(1913) <= not b;
    outputs(1914) <= b;
    outputs(1915) <= a xor b;
    outputs(1916) <= b and not a;
    outputs(1917) <= not (a xor b);
    outputs(1918) <= a and not b;
    outputs(1919) <= not b;
    outputs(1920) <= not b;
    outputs(1921) <= not b;
    outputs(1922) <= not (a xor b);
    outputs(1923) <= a and not b;
    outputs(1924) <= b and not a;
    outputs(1925) <= not a;
    outputs(1926) <= b;
    outputs(1927) <= not a or b;
    outputs(1928) <= not b or a;
    outputs(1929) <= a and b;
    outputs(1930) <= b;
    outputs(1931) <= a or b;
    outputs(1932) <= not b;
    outputs(1933) <= a and not b;
    outputs(1934) <= a xor b;
    outputs(1935) <= b and not a;
    outputs(1936) <= not a;
    outputs(1937) <= not b;
    outputs(1938) <= a xor b;
    outputs(1939) <= not b or a;
    outputs(1940) <= a;
    outputs(1941) <= a xor b;
    outputs(1942) <= a xor b;
    outputs(1943) <= b;
    outputs(1944) <= not a;
    outputs(1945) <= not (a xor b);
    outputs(1946) <= not a;
    outputs(1947) <= not a;
    outputs(1948) <= a xor b;
    outputs(1949) <= b;
    outputs(1950) <= not (a xor b);
    outputs(1951) <= not b;
    outputs(1952) <= b;
    outputs(1953) <= not a;
    outputs(1954) <= not b;
    outputs(1955) <= a and b;
    outputs(1956) <= not a;
    outputs(1957) <= not (a and b);
    outputs(1958) <= a;
    outputs(1959) <= not (a xor b);
    outputs(1960) <= not (a xor b);
    outputs(1961) <= not (a xor b);
    outputs(1962) <= b;
    outputs(1963) <= b;
    outputs(1964) <= not (a xor b);
    outputs(1965) <= not b;
    outputs(1966) <= a;
    outputs(1967) <= not b or a;
    outputs(1968) <= not a;
    outputs(1969) <= not b;
    outputs(1970) <= b;
    outputs(1971) <= a and b;
    outputs(1972) <= not b;
    outputs(1973) <= not a;
    outputs(1974) <= a xor b;
    outputs(1975) <= b;
    outputs(1976) <= not (a and b);
    outputs(1977) <= a and not b;
    outputs(1978) <= b;
    outputs(1979) <= not (a xor b);
    outputs(1980) <= a;
    outputs(1981) <= not a or b;
    outputs(1982) <= b;
    outputs(1983) <= a xor b;
    outputs(1984) <= a;
    outputs(1985) <= not a;
    outputs(1986) <= not b;
    outputs(1987) <= b and not a;
    outputs(1988) <= b;
    outputs(1989) <= not a;
    outputs(1990) <= b;
    outputs(1991) <= a and b;
    outputs(1992) <= b;
    outputs(1993) <= a and b;
    outputs(1994) <= not a;
    outputs(1995) <= not (a xor b);
    outputs(1996) <= a xor b;
    outputs(1997) <= not (a and b);
    outputs(1998) <= a and b;
    outputs(1999) <= b;
    outputs(2000) <= a xor b;
    outputs(2001) <= a and not b;
    outputs(2002) <= not (a and b);
    outputs(2003) <= a xor b;
    outputs(2004) <= a;
    outputs(2005) <= not (a xor b);
    outputs(2006) <= not (a or b);
    outputs(2007) <= a and b;
    outputs(2008) <= not a;
    outputs(2009) <= a and not b;
    outputs(2010) <= a;
    outputs(2011) <= not a;
    outputs(2012) <= not a;
    outputs(2013) <= not a or b;
    outputs(2014) <= a;
    outputs(2015) <= not (a and b);
    outputs(2016) <= a and not b;
    outputs(2017) <= not a;
    outputs(2018) <= not a;
    outputs(2019) <= a or b;
    outputs(2020) <= not b;
    outputs(2021) <= a and b;
    outputs(2022) <= not b;
    outputs(2023) <= a xor b;
    outputs(2024) <= not b;
    outputs(2025) <= not a;
    outputs(2026) <= b;
    outputs(2027) <= a;
    outputs(2028) <= a or b;
    outputs(2029) <= b;
    outputs(2030) <= not a;
    outputs(2031) <= a and not b;
    outputs(2032) <= not b or a;
    outputs(2033) <= not a;
    outputs(2034) <= not (a or b);
    outputs(2035) <= not a;
    outputs(2036) <= a and not b;
    outputs(2037) <= b and not a;
    outputs(2038) <= a;
    outputs(2039) <= not (a xor b);
    outputs(2040) <= a and not b;
    outputs(2041) <= not (a or b);
    outputs(2042) <= not (a or b);
    outputs(2043) <= a xor b;
    outputs(2044) <= not b;
    outputs(2045) <= a or b;
    outputs(2046) <= a or b;
    outputs(2047) <= not a;
    outputs(2048) <= a;
    outputs(2049) <= a and b;
    outputs(2050) <= a;
    outputs(2051) <= b;
    outputs(2052) <= a xor b;
    outputs(2053) <= not b;
    outputs(2054) <= a and not b;
    outputs(2055) <= a and b;
    outputs(2056) <= a xor b;
    outputs(2057) <= a;
    outputs(2058) <= b;
    outputs(2059) <= b;
    outputs(2060) <= not a or b;
    outputs(2061) <= a xor b;
    outputs(2062) <= a;
    outputs(2063) <= a and not b;
    outputs(2064) <= b and not a;
    outputs(2065) <= not b;
    outputs(2066) <= b;
    outputs(2067) <= not b;
    outputs(2068) <= b and not a;
    outputs(2069) <= b;
    outputs(2070) <= b;
    outputs(2071) <= b;
    outputs(2072) <= not b;
    outputs(2073) <= not (a xor b);
    outputs(2074) <= not a;
    outputs(2075) <= not a;
    outputs(2076) <= b;
    outputs(2077) <= not b;
    outputs(2078) <= not b;
    outputs(2079) <= a and b;
    outputs(2080) <= a and not b;
    outputs(2081) <= b and not a;
    outputs(2082) <= a;
    outputs(2083) <= not (a xor b);
    outputs(2084) <= b;
    outputs(2085) <= b;
    outputs(2086) <= a xor b;
    outputs(2087) <= a;
    outputs(2088) <= not (a xor b);
    outputs(2089) <= not b;
    outputs(2090) <= not (a or b);
    outputs(2091) <= not a;
    outputs(2092) <= a;
    outputs(2093) <= a;
    outputs(2094) <= b;
    outputs(2095) <= a;
    outputs(2096) <= not (a xor b);
    outputs(2097) <= not a;
    outputs(2098) <= a;
    outputs(2099) <= b;
    outputs(2100) <= a xor b;
    outputs(2101) <= not (a xor b);
    outputs(2102) <= a;
    outputs(2103) <= b and not a;
    outputs(2104) <= a and not b;
    outputs(2105) <= not a;
    outputs(2106) <= a xor b;
    outputs(2107) <= b;
    outputs(2108) <= b and not a;
    outputs(2109) <= b;
    outputs(2110) <= not (a or b);
    outputs(2111) <= not b;
    outputs(2112) <= not a;
    outputs(2113) <= not (a xor b);
    outputs(2114) <= a xor b;
    outputs(2115) <= not b;
    outputs(2116) <= not b or a;
    outputs(2117) <= a;
    outputs(2118) <= not a;
    outputs(2119) <= b;
    outputs(2120) <= not (a and b);
    outputs(2121) <= b;
    outputs(2122) <= not a or b;
    outputs(2123) <= b;
    outputs(2124) <= a xor b;
    outputs(2125) <= not a;
    outputs(2126) <= not b;
    outputs(2127) <= a and b;
    outputs(2128) <= not (a or b);
    outputs(2129) <= a and not b;
    outputs(2130) <= b;
    outputs(2131) <= not a;
    outputs(2132) <= a;
    outputs(2133) <= b;
    outputs(2134) <= not a;
    outputs(2135) <= not a;
    outputs(2136) <= a xor b;
    outputs(2137) <= b;
    outputs(2138) <= a and b;
    outputs(2139) <= not (a or b);
    outputs(2140) <= not b or a;
    outputs(2141) <= a and not b;
    outputs(2142) <= b;
    outputs(2143) <= b and not a;
    outputs(2144) <= b and not a;
    outputs(2145) <= b and not a;
    outputs(2146) <= not b;
    outputs(2147) <= b;
    outputs(2148) <= not (a xor b);
    outputs(2149) <= a;
    outputs(2150) <= not b;
    outputs(2151) <= a;
    outputs(2152) <= not a;
    outputs(2153) <= not a or b;
    outputs(2154) <= not (a xor b);
    outputs(2155) <= not (a or b);
    outputs(2156) <= a or b;
    outputs(2157) <= not b;
    outputs(2158) <= a and b;
    outputs(2159) <= a and b;
    outputs(2160) <= not a;
    outputs(2161) <= not (a or b);
    outputs(2162) <= not b;
    outputs(2163) <= not (a or b);
    outputs(2164) <= not (a or b);
    outputs(2165) <= not (a xor b);
    outputs(2166) <= a xor b;
    outputs(2167) <= b;
    outputs(2168) <= b and not a;
    outputs(2169) <= not b;
    outputs(2170) <= not (a xor b);
    outputs(2171) <= b;
    outputs(2172) <= not (a or b);
    outputs(2173) <= b;
    outputs(2174) <= not b;
    outputs(2175) <= not b;
    outputs(2176) <= not b;
    outputs(2177) <= not b;
    outputs(2178) <= not b;
    outputs(2179) <= a and b;
    outputs(2180) <= a;
    outputs(2181) <= not b;
    outputs(2182) <= a;
    outputs(2183) <= a or b;
    outputs(2184) <= b;
    outputs(2185) <= a;
    outputs(2186) <= not a;
    outputs(2187) <= a;
    outputs(2188) <= not a;
    outputs(2189) <= a and b;
    outputs(2190) <= not b;
    outputs(2191) <= a and not b;
    outputs(2192) <= not b;
    outputs(2193) <= a and not b;
    outputs(2194) <= not (a or b);
    outputs(2195) <= not (a xor b);
    outputs(2196) <= b;
    outputs(2197) <= a and not b;
    outputs(2198) <= not a;
    outputs(2199) <= not (a and b);
    outputs(2200) <= a;
    outputs(2201) <= not a;
    outputs(2202) <= not (a xor b);
    outputs(2203) <= not b or a;
    outputs(2204) <= not a;
    outputs(2205) <= b;
    outputs(2206) <= b;
    outputs(2207) <= a and not b;
    outputs(2208) <= a xor b;
    outputs(2209) <= b;
    outputs(2210) <= not (a and b);
    outputs(2211) <= b and not a;
    outputs(2212) <= a xor b;
    outputs(2213) <= a or b;
    outputs(2214) <= not (a or b);
    outputs(2215) <= a and not b;
    outputs(2216) <= a and b;
    outputs(2217) <= not (a xor b);
    outputs(2218) <= not b;
    outputs(2219) <= not b or a;
    outputs(2220) <= not b;
    outputs(2221) <= a;
    outputs(2222) <= not b;
    outputs(2223) <= a or b;
    outputs(2224) <= a;
    outputs(2225) <= a or b;
    outputs(2226) <= not a;
    outputs(2227) <= a xor b;
    outputs(2228) <= not a;
    outputs(2229) <= not a;
    outputs(2230) <= not a;
    outputs(2231) <= not (a xor b);
    outputs(2232) <= a and b;
    outputs(2233) <= b and not a;
    outputs(2234) <= not (a xor b);
    outputs(2235) <= not a or b;
    outputs(2236) <= not b;
    outputs(2237) <= b;
    outputs(2238) <= a xor b;
    outputs(2239) <= b and not a;
    outputs(2240) <= b;
    outputs(2241) <= a xor b;
    outputs(2242) <= not b;
    outputs(2243) <= b;
    outputs(2244) <= not a;
    outputs(2245) <= a;
    outputs(2246) <= a;
    outputs(2247) <= not b or a;
    outputs(2248) <= not (a or b);
    outputs(2249) <= not (a xor b);
    outputs(2250) <= a and b;
    outputs(2251) <= not b;
    outputs(2252) <= not b;
    outputs(2253) <= b and not a;
    outputs(2254) <= a or b;
    outputs(2255) <= not (a or b);
    outputs(2256) <= not b;
    outputs(2257) <= a;
    outputs(2258) <= not b;
    outputs(2259) <= b and not a;
    outputs(2260) <= a xor b;
    outputs(2261) <= not b or a;
    outputs(2262) <= not (a xor b);
    outputs(2263) <= not a;
    outputs(2264) <= not (a xor b);
    outputs(2265) <= not a or b;
    outputs(2266) <= not (a xor b);
    outputs(2267) <= a;
    outputs(2268) <= a;
    outputs(2269) <= not (a xor b);
    outputs(2270) <= not a;
    outputs(2271) <= not a;
    outputs(2272) <= a and not b;
    outputs(2273) <= b;
    outputs(2274) <= a xor b;
    outputs(2275) <= b;
    outputs(2276) <= b;
    outputs(2277) <= b and not a;
    outputs(2278) <= a;
    outputs(2279) <= a and not b;
    outputs(2280) <= a and not b;
    outputs(2281) <= not a or b;
    outputs(2282) <= not a;
    outputs(2283) <= a and not b;
    outputs(2284) <= a xor b;
    outputs(2285) <= a;
    outputs(2286) <= not (a and b);
    outputs(2287) <= a;
    outputs(2288) <= not a;
    outputs(2289) <= not a;
    outputs(2290) <= not (a xor b);
    outputs(2291) <= a and not b;
    outputs(2292) <= not (a or b);
    outputs(2293) <= a or b;
    outputs(2294) <= a and b;
    outputs(2295) <= not a;
    outputs(2296) <= not (a xor b);
    outputs(2297) <= a;
    outputs(2298) <= b;
    outputs(2299) <= not (a or b);
    outputs(2300) <= not a;
    outputs(2301) <= not a or b;
    outputs(2302) <= a;
    outputs(2303) <= b;
    outputs(2304) <= a;
    outputs(2305) <= a or b;
    outputs(2306) <= not a;
    outputs(2307) <= not a;
    outputs(2308) <= not (a and b);
    outputs(2309) <= a and b;
    outputs(2310) <= a or b;
    outputs(2311) <= a;
    outputs(2312) <= not b;
    outputs(2313) <= not (a xor b);
    outputs(2314) <= a and not b;
    outputs(2315) <= a and b;
    outputs(2316) <= not (a xor b);
    outputs(2317) <= a and not b;
    outputs(2318) <= b;
    outputs(2319) <= not b;
    outputs(2320) <= not a;
    outputs(2321) <= not a;
    outputs(2322) <= b;
    outputs(2323) <= a xor b;
    outputs(2324) <= not a;
    outputs(2325) <= a xor b;
    outputs(2326) <= b;
    outputs(2327) <= b and not a;
    outputs(2328) <= not a;
    outputs(2329) <= a and b;
    outputs(2330) <= a and not b;
    outputs(2331) <= not a or b;
    outputs(2332) <= b;
    outputs(2333) <= not (a xor b);
    outputs(2334) <= not b or a;
    outputs(2335) <= a;
    outputs(2336) <= b;
    outputs(2337) <= not b;
    outputs(2338) <= b and not a;
    outputs(2339) <= not (a xor b);
    outputs(2340) <= b;
    outputs(2341) <= not a;
    outputs(2342) <= not (a xor b);
    outputs(2343) <= b and not a;
    outputs(2344) <= not a;
    outputs(2345) <= not (a or b);
    outputs(2346) <= a and b;
    outputs(2347) <= a or b;
    outputs(2348) <= not (a xor b);
    outputs(2349) <= not b;
    outputs(2350) <= not b;
    outputs(2351) <= b;
    outputs(2352) <= a and b;
    outputs(2353) <= not a;
    outputs(2354) <= not b;
    outputs(2355) <= not (a or b);
    outputs(2356) <= a;
    outputs(2357) <= b and not a;
    outputs(2358) <= a and b;
    outputs(2359) <= not b;
    outputs(2360) <= not b;
    outputs(2361) <= b;
    outputs(2362) <= a and b;
    outputs(2363) <= not (a xor b);
    outputs(2364) <= not (a or b);
    outputs(2365) <= b;
    outputs(2366) <= not (a or b);
    outputs(2367) <= not a;
    outputs(2368) <= a xor b;
    outputs(2369) <= a and not b;
    outputs(2370) <= a;
    outputs(2371) <= not a;
    outputs(2372) <= not a;
    outputs(2373) <= a and not b;
    outputs(2374) <= a and not b;
    outputs(2375) <= not (a or b);
    outputs(2376) <= not a or b;
    outputs(2377) <= not b or a;
    outputs(2378) <= not (a xor b);
    outputs(2379) <= a and b;
    outputs(2380) <= not a;
    outputs(2381) <= a;
    outputs(2382) <= not a;
    outputs(2383) <= not a;
    outputs(2384) <= not b;
    outputs(2385) <= a and b;
    outputs(2386) <= not a;
    outputs(2387) <= a;
    outputs(2388) <= not a;
    outputs(2389) <= a and not b;
    outputs(2390) <= not b or a;
    outputs(2391) <= a;
    outputs(2392) <= a and not b;
    outputs(2393) <= not a;
    outputs(2394) <= b;
    outputs(2395) <= a and b;
    outputs(2396) <= not a;
    outputs(2397) <= b and not a;
    outputs(2398) <= not b;
    outputs(2399) <= a;
    outputs(2400) <= not a or b;
    outputs(2401) <= a or b;
    outputs(2402) <= a;
    outputs(2403) <= not (a or b);
    outputs(2404) <= not (a and b);
    outputs(2405) <= a;
    outputs(2406) <= b;
    outputs(2407) <= a and not b;
    outputs(2408) <= a;
    outputs(2409) <= not (a or b);
    outputs(2410) <= not a;
    outputs(2411) <= a and b;
    outputs(2412) <= not b;
    outputs(2413) <= not (a xor b);
    outputs(2414) <= not (a xor b);
    outputs(2415) <= not (a or b);
    outputs(2416) <= b and not a;
    outputs(2417) <= not b;
    outputs(2418) <= a;
    outputs(2419) <= not a or b;
    outputs(2420) <= a;
    outputs(2421) <= not a;
    outputs(2422) <= a and b;
    outputs(2423) <= a;
    outputs(2424) <= not b;
    outputs(2425) <= a and b;
    outputs(2426) <= a and b;
    outputs(2427) <= not (a or b);
    outputs(2428) <= a and b;
    outputs(2429) <= a;
    outputs(2430) <= a;
    outputs(2431) <= a;
    outputs(2432) <= not a;
    outputs(2433) <= not a;
    outputs(2434) <= a or b;
    outputs(2435) <= a and not b;
    outputs(2436) <= not (a or b);
    outputs(2437) <= not a;
    outputs(2438) <= not a;
    outputs(2439) <= a;
    outputs(2440) <= not b;
    outputs(2441) <= b and not a;
    outputs(2442) <= a and b;
    outputs(2443) <= not (a xor b);
    outputs(2444) <= not a;
    outputs(2445) <= a and not b;
    outputs(2446) <= a;
    outputs(2447) <= a and not b;
    outputs(2448) <= b and not a;
    outputs(2449) <= b and not a;
    outputs(2450) <= a and not b;
    outputs(2451) <= b and not a;
    outputs(2452) <= a and not b;
    outputs(2453) <= not (a or b);
    outputs(2454) <= a;
    outputs(2455) <= b and not a;
    outputs(2456) <= a and b;
    outputs(2457) <= not a;
    outputs(2458) <= a and not b;
    outputs(2459) <= b and not a;
    outputs(2460) <= not (a xor b);
    outputs(2461) <= not b;
    outputs(2462) <= a and not b;
    outputs(2463) <= not (a or b);
    outputs(2464) <= not a;
    outputs(2465) <= a;
    outputs(2466) <= not b;
    outputs(2467) <= not b;
    outputs(2468) <= not b or a;
    outputs(2469) <= not a;
    outputs(2470) <= a;
    outputs(2471) <= not a;
    outputs(2472) <= b;
    outputs(2473) <= not a;
    outputs(2474) <= not a;
    outputs(2475) <= a xor b;
    outputs(2476) <= not b;
    outputs(2477) <= not b;
    outputs(2478) <= b;
    outputs(2479) <= a xor b;
    outputs(2480) <= a;
    outputs(2481) <= a;
    outputs(2482) <= b;
    outputs(2483) <= b;
    outputs(2484) <= a and not b;
    outputs(2485) <= not (a or b);
    outputs(2486) <= a and not b;
    outputs(2487) <= not b;
    outputs(2488) <= not a;
    outputs(2489) <= a or b;
    outputs(2490) <= b;
    outputs(2491) <= b;
    outputs(2492) <= a and not b;
    outputs(2493) <= not b;
    outputs(2494) <= a and b;
    outputs(2495) <= a and b;
    outputs(2496) <= not (a or b);
    outputs(2497) <= b;
    outputs(2498) <= b;
    outputs(2499) <= not b;
    outputs(2500) <= not b;
    outputs(2501) <= not b;
    outputs(2502) <= a;
    outputs(2503) <= a;
    outputs(2504) <= b and not a;
    outputs(2505) <= not a;
    outputs(2506) <= not a or b;
    outputs(2507) <= not (a or b);
    outputs(2508) <= a;
    outputs(2509) <= a;
    outputs(2510) <= not a;
    outputs(2511) <= b and not a;
    outputs(2512) <= a;
    outputs(2513) <= not a;
    outputs(2514) <= a;
    outputs(2515) <= a;
    outputs(2516) <= b;
    outputs(2517) <= a;
    outputs(2518) <= not (a and b);
    outputs(2519) <= a and not b;
    outputs(2520) <= not a;
    outputs(2521) <= not a or b;
    outputs(2522) <= not a or b;
    outputs(2523) <= a xor b;
    outputs(2524) <= b;
    outputs(2525) <= not a;
    outputs(2526) <= a;
    outputs(2527) <= not b;
    outputs(2528) <= a and not b;
    outputs(2529) <= a and not b;
    outputs(2530) <= not (a and b);
    outputs(2531) <= not a;
    outputs(2532) <= b;
    outputs(2533) <= a and b;
    outputs(2534) <= not a;
    outputs(2535) <= not b;
    outputs(2536) <= a;
    outputs(2537) <= not (a xor b);
    outputs(2538) <= not a;
    outputs(2539) <= not (a or b);
    outputs(2540) <= a and b;
    outputs(2541) <= a xor b;
    outputs(2542) <= a;
    outputs(2543) <= not (a or b);
    outputs(2544) <= a or b;
    outputs(2545) <= a and not b;
    outputs(2546) <= b;
    outputs(2547) <= b;
    outputs(2548) <= not b;
    outputs(2549) <= not (a or b);
    outputs(2550) <= a;
    outputs(2551) <= a and not b;
    outputs(2552) <= a and not b;
    outputs(2553) <= a;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= b;
    outputs(2556) <= not b;
    outputs(2557) <= not (a xor b);
    outputs(2558) <= b;
    outputs(2559) <= a and not b;
    outputs(2560) <= not b;
    outputs(2561) <= a;
    outputs(2562) <= not a;
    outputs(2563) <= a;
    outputs(2564) <= not b;
    outputs(2565) <= a;
    outputs(2566) <= not (a xor b);
    outputs(2567) <= not a;
    outputs(2568) <= not b or a;
    outputs(2569) <= a and b;
    outputs(2570) <= a;
    outputs(2571) <= b;
    outputs(2572) <= not (a xor b);
    outputs(2573) <= not b;
    outputs(2574) <= not a;
    outputs(2575) <= not a;
    outputs(2576) <= not (a xor b);
    outputs(2577) <= not a;
    outputs(2578) <= not a;
    outputs(2579) <= a and not b;
    outputs(2580) <= not (a or b);
    outputs(2581) <= b;
    outputs(2582) <= b;
    outputs(2583) <= not a;
    outputs(2584) <= not b;
    outputs(2585) <= a and b;
    outputs(2586) <= a and not b;
    outputs(2587) <= a;
    outputs(2588) <= a;
    outputs(2589) <= not (a xor b);
    outputs(2590) <= a xor b;
    outputs(2591) <= not (a xor b);
    outputs(2592) <= not a;
    outputs(2593) <= not (a xor b);
    outputs(2594) <= not a;
    outputs(2595) <= a xor b;
    outputs(2596) <= not a;
    outputs(2597) <= not (a xor b);
    outputs(2598) <= a xor b;
    outputs(2599) <= not (a xor b);
    outputs(2600) <= not (a xor b);
    outputs(2601) <= a xor b;
    outputs(2602) <= a and not b;
    outputs(2603) <= a;
    outputs(2604) <= not (a or b);
    outputs(2605) <= a;
    outputs(2606) <= not b;
    outputs(2607) <= not a;
    outputs(2608) <= not (a xor b);
    outputs(2609) <= b and not a;
    outputs(2610) <= a or b;
    outputs(2611) <= a;
    outputs(2612) <= a and b;
    outputs(2613) <= a;
    outputs(2614) <= not b;
    outputs(2615) <= a and not b;
    outputs(2616) <= b;
    outputs(2617) <= not b;
    outputs(2618) <= b;
    outputs(2619) <= a;
    outputs(2620) <= not b or a;
    outputs(2621) <= a;
    outputs(2622) <= a;
    outputs(2623) <= a xor b;
    outputs(2624) <= a and b;
    outputs(2625) <= not (a xor b);
    outputs(2626) <= a and not b;
    outputs(2627) <= not b;
    outputs(2628) <= a xor b;
    outputs(2629) <= a;
    outputs(2630) <= not a;
    outputs(2631) <= not b or a;
    outputs(2632) <= a;
    outputs(2633) <= a;
    outputs(2634) <= a xor b;
    outputs(2635) <= not (a xor b);
    outputs(2636) <= b;
    outputs(2637) <= b;
    outputs(2638) <= a and not b;
    outputs(2639) <= not (a xor b);
    outputs(2640) <= not a;
    outputs(2641) <= a or b;
    outputs(2642) <= a;
    outputs(2643) <= not (a and b);
    outputs(2644) <= a or b;
    outputs(2645) <= not b;
    outputs(2646) <= b and not a;
    outputs(2647) <= b;
    outputs(2648) <= a;
    outputs(2649) <= a or b;
    outputs(2650) <= a xor b;
    outputs(2651) <= not (a xor b);
    outputs(2652) <= not a;
    outputs(2653) <= not b or a;
    outputs(2654) <= not a;
    outputs(2655) <= not (a xor b);
    outputs(2656) <= a or b;
    outputs(2657) <= b;
    outputs(2658) <= a or b;
    outputs(2659) <= not (a xor b);
    outputs(2660) <= a xor b;
    outputs(2661) <= not a or b;
    outputs(2662) <= not (a or b);
    outputs(2663) <= not a;
    outputs(2664) <= a and not b;
    outputs(2665) <= not b;
    outputs(2666) <= not a;
    outputs(2667) <= not b;
    outputs(2668) <= a xor b;
    outputs(2669) <= not a;
    outputs(2670) <= a xor b;
    outputs(2671) <= a and not b;
    outputs(2672) <= a xor b;
    outputs(2673) <= a xor b;
    outputs(2674) <= a xor b;
    outputs(2675) <= not b;
    outputs(2676) <= not b;
    outputs(2677) <= a and not b;
    outputs(2678) <= not b or a;
    outputs(2679) <= not b;
    outputs(2680) <= not (a xor b);
    outputs(2681) <= not a;
    outputs(2682) <= not b;
    outputs(2683) <= not (a or b);
    outputs(2684) <= not (a xor b);
    outputs(2685) <= b and not a;
    outputs(2686) <= not a;
    outputs(2687) <= a xor b;
    outputs(2688) <= a xor b;
    outputs(2689) <= a or b;
    outputs(2690) <= not (a xor b);
    outputs(2691) <= a xor b;
    outputs(2692) <= a xor b;
    outputs(2693) <= a;
    outputs(2694) <= not (a or b);
    outputs(2695) <= a and b;
    outputs(2696) <= a and b;
    outputs(2697) <= b;
    outputs(2698) <= a xor b;
    outputs(2699) <= a;
    outputs(2700) <= not (a or b);
    outputs(2701) <= not a;
    outputs(2702) <= a;
    outputs(2703) <= b and not a;
    outputs(2704) <= b;
    outputs(2705) <= a;
    outputs(2706) <= not (a xor b);
    outputs(2707) <= not (a or b);
    outputs(2708) <= a xor b;
    outputs(2709) <= not b or a;
    outputs(2710) <= a xor b;
    outputs(2711) <= not a;
    outputs(2712) <= not a;
    outputs(2713) <= not a;
    outputs(2714) <= a;
    outputs(2715) <= a or b;
    outputs(2716) <= a and b;
    outputs(2717) <= not (a xor b);
    outputs(2718) <= not a or b;
    outputs(2719) <= a xor b;
    outputs(2720) <= not (a and b);
    outputs(2721) <= a and b;
    outputs(2722) <= not (a xor b);
    outputs(2723) <= not b;
    outputs(2724) <= not (a xor b);
    outputs(2725) <= b;
    outputs(2726) <= a;
    outputs(2727) <= b;
    outputs(2728) <= a or b;
    outputs(2729) <= a xor b;
    outputs(2730) <= b;
    outputs(2731) <= a xor b;
    outputs(2732) <= not (a and b);
    outputs(2733) <= b and not a;
    outputs(2734) <= a;
    outputs(2735) <= a xor b;
    outputs(2736) <= b;
    outputs(2737) <= not (a or b);
    outputs(2738) <= not (a xor b);
    outputs(2739) <= not a;
    outputs(2740) <= not b;
    outputs(2741) <= not a;
    outputs(2742) <= a and b;
    outputs(2743) <= not (a xor b);
    outputs(2744) <= not b;
    outputs(2745) <= not a;
    outputs(2746) <= not a;
    outputs(2747) <= not a or b;
    outputs(2748) <= a;
    outputs(2749) <= not a or b;
    outputs(2750) <= not b;
    outputs(2751) <= not b;
    outputs(2752) <= not (a xor b);
    outputs(2753) <= not b or a;
    outputs(2754) <= a and not b;
    outputs(2755) <= not b;
    outputs(2756) <= a and b;
    outputs(2757) <= a;
    outputs(2758) <= not a;
    outputs(2759) <= not b;
    outputs(2760) <= b and not a;
    outputs(2761) <= a;
    outputs(2762) <= a;
    outputs(2763) <= not b;
    outputs(2764) <= a xor b;
    outputs(2765) <= not (a xor b);
    outputs(2766) <= b;
    outputs(2767) <= a xor b;
    outputs(2768) <= not a;
    outputs(2769) <= not a;
    outputs(2770) <= b;
    outputs(2771) <= not (a and b);
    outputs(2772) <= not a;
    outputs(2773) <= not (a or b);
    outputs(2774) <= b;
    outputs(2775) <= b and not a;
    outputs(2776) <= not a;
    outputs(2777) <= a xor b;
    outputs(2778) <= b;
    outputs(2779) <= not a;
    outputs(2780) <= a xor b;
    outputs(2781) <= b;
    outputs(2782) <= not b;
    outputs(2783) <= not b;
    outputs(2784) <= not (a xor b);
    outputs(2785) <= a and b;
    outputs(2786) <= b and not a;
    outputs(2787) <= b;
    outputs(2788) <= not a;
    outputs(2789) <= a and not b;
    outputs(2790) <= a and not b;
    outputs(2791) <= not (a and b);
    outputs(2792) <= not b;
    outputs(2793) <= a xor b;
    outputs(2794) <= a and b;
    outputs(2795) <= not (a xor b);
    outputs(2796) <= not b;
    outputs(2797) <= not b;
    outputs(2798) <= a;
    outputs(2799) <= not b or a;
    outputs(2800) <= not (a xor b);
    outputs(2801) <= not (a xor b);
    outputs(2802) <= not (a and b);
    outputs(2803) <= a xor b;
    outputs(2804) <= not (a or b);
    outputs(2805) <= not (a xor b);
    outputs(2806) <= not b;
    outputs(2807) <= a and not b;
    outputs(2808) <= a or b;
    outputs(2809) <= b;
    outputs(2810) <= not b;
    outputs(2811) <= b;
    outputs(2812) <= not (a xor b);
    outputs(2813) <= not b;
    outputs(2814) <= a xor b;
    outputs(2815) <= not a;
    outputs(2816) <= a;
    outputs(2817) <= not (a or b);
    outputs(2818) <= not (a and b);
    outputs(2819) <= b;
    outputs(2820) <= a and not b;
    outputs(2821) <= not b or a;
    outputs(2822) <= a and not b;
    outputs(2823) <= b;
    outputs(2824) <= a;
    outputs(2825) <= not (a xor b);
    outputs(2826) <= b;
    outputs(2827) <= not (a or b);
    outputs(2828) <= not (a or b);
    outputs(2829) <= not (a or b);
    outputs(2830) <= a xor b;
    outputs(2831) <= not b or a;
    outputs(2832) <= a and b;
    outputs(2833) <= not (a or b);
    outputs(2834) <= not a;
    outputs(2835) <= not b;
    outputs(2836) <= not a;
    outputs(2837) <= not a;
    outputs(2838) <= not a or b;
    outputs(2839) <= b;
    outputs(2840) <= b and not a;
    outputs(2841) <= b and not a;
    outputs(2842) <= not a;
    outputs(2843) <= b and not a;
    outputs(2844) <= a and b;
    outputs(2845) <= not (a xor b);
    outputs(2846) <= a and b;
    outputs(2847) <= b;
    outputs(2848) <= a xor b;
    outputs(2849) <= not (a and b);
    outputs(2850) <= a or b;
    outputs(2851) <= not (a xor b);
    outputs(2852) <= not b;
    outputs(2853) <= a and not b;
    outputs(2854) <= b and not a;
    outputs(2855) <= not (a xor b);
    outputs(2856) <= a and b;
    outputs(2857) <= a and b;
    outputs(2858) <= b;
    outputs(2859) <= a;
    outputs(2860) <= not b;
    outputs(2861) <= not a;
    outputs(2862) <= a and not b;
    outputs(2863) <= a or b;
    outputs(2864) <= not a or b;
    outputs(2865) <= not (a or b);
    outputs(2866) <= a;
    outputs(2867) <= b;
    outputs(2868) <= b and not a;
    outputs(2869) <= a xor b;
    outputs(2870) <= a;
    outputs(2871) <= a xor b;
    outputs(2872) <= b;
    outputs(2873) <= not (a and b);
    outputs(2874) <= a xor b;
    outputs(2875) <= a xor b;
    outputs(2876) <= b;
    outputs(2877) <= a and not b;
    outputs(2878) <= a;
    outputs(2879) <= b;
    outputs(2880) <= not a;
    outputs(2881) <= b;
    outputs(2882) <= b and not a;
    outputs(2883) <= not a;
    outputs(2884) <= not b;
    outputs(2885) <= not a or b;
    outputs(2886) <= b;
    outputs(2887) <= b;
    outputs(2888) <= b;
    outputs(2889) <= a xor b;
    outputs(2890) <= not (a and b);
    outputs(2891) <= not (a and b);
    outputs(2892) <= not (a xor b);
    outputs(2893) <= a xor b;
    outputs(2894) <= not (a xor b);
    outputs(2895) <= b and not a;
    outputs(2896) <= not a;
    outputs(2897) <= a xor b;
    outputs(2898) <= a;
    outputs(2899) <= not b or a;
    outputs(2900) <= a xor b;
    outputs(2901) <= not (a xor b);
    outputs(2902) <= b and not a;
    outputs(2903) <= not a;
    outputs(2904) <= not a or b;
    outputs(2905) <= not b;
    outputs(2906) <= b;
    outputs(2907) <= a;
    outputs(2908) <= a;
    outputs(2909) <= not a;
    outputs(2910) <= b;
    outputs(2911) <= a;
    outputs(2912) <= not (a xor b);
    outputs(2913) <= not (a xor b);
    outputs(2914) <= not (a xor b);
    outputs(2915) <= not (a and b);
    outputs(2916) <= a xor b;
    outputs(2917) <= a xor b;
    outputs(2918) <= not a;
    outputs(2919) <= a xor b;
    outputs(2920) <= a xor b;
    outputs(2921) <= not b or a;
    outputs(2922) <= not (a xor b);
    outputs(2923) <= b;
    outputs(2924) <= not (a xor b);
    outputs(2925) <= a and b;
    outputs(2926) <= a and b;
    outputs(2927) <= not (a xor b);
    outputs(2928) <= not a;
    outputs(2929) <= not b;
    outputs(2930) <= a;
    outputs(2931) <= b;
    outputs(2932) <= b and not a;
    outputs(2933) <= not (a or b);
    outputs(2934) <= a and b;
    outputs(2935) <= a xor b;
    outputs(2936) <= not a;
    outputs(2937) <= b and not a;
    outputs(2938) <= not (a xor b);
    outputs(2939) <= not a;
    outputs(2940) <= b;
    outputs(2941) <= b and not a;
    outputs(2942) <= not (a xor b);
    outputs(2943) <= not a;
    outputs(2944) <= not (a xor b);
    outputs(2945) <= a;
    outputs(2946) <= a;
    outputs(2947) <= a xor b;
    outputs(2948) <= not (a or b);
    outputs(2949) <= not (a xor b);
    outputs(2950) <= a xor b;
    outputs(2951) <= not (a xor b);
    outputs(2952) <= b;
    outputs(2953) <= not a;
    outputs(2954) <= not a;
    outputs(2955) <= a xor b;
    outputs(2956) <= not b;
    outputs(2957) <= not (a or b);
    outputs(2958) <= b;
    outputs(2959) <= not a or b;
    outputs(2960) <= not (a xor b);
    outputs(2961) <= b and not a;
    outputs(2962) <= not b;
    outputs(2963) <= not b;
    outputs(2964) <= not a;
    outputs(2965) <= not a;
    outputs(2966) <= not b;
    outputs(2967) <= not a or b;
    outputs(2968) <= a xor b;
    outputs(2969) <= a xor b;
    outputs(2970) <= not (a xor b);
    outputs(2971) <= a;
    outputs(2972) <= not (a xor b);
    outputs(2973) <= not b;
    outputs(2974) <= a or b;
    outputs(2975) <= not a;
    outputs(2976) <= not a;
    outputs(2977) <= not b;
    outputs(2978) <= a and b;
    outputs(2979) <= b;
    outputs(2980) <= b;
    outputs(2981) <= a;
    outputs(2982) <= b;
    outputs(2983) <= not (a xor b);
    outputs(2984) <= a xor b;
    outputs(2985) <= a;
    outputs(2986) <= not (a or b);
    outputs(2987) <= a xor b;
    outputs(2988) <= a and b;
    outputs(2989) <= not (a xor b);
    outputs(2990) <= not (a xor b);
    outputs(2991) <= a and b;
    outputs(2992) <= not (a or b);
    outputs(2993) <= not (a xor b);
    outputs(2994) <= not b or a;
    outputs(2995) <= b and not a;
    outputs(2996) <= a xor b;
    outputs(2997) <= not (a xor b);
    outputs(2998) <= not a or b;
    outputs(2999) <= not (a xor b);
    outputs(3000) <= not a;
    outputs(3001) <= not a;
    outputs(3002) <= not b or a;
    outputs(3003) <= not b;
    outputs(3004) <= not (a or b);
    outputs(3005) <= not b or a;
    outputs(3006) <= a and b;
    outputs(3007) <= a xor b;
    outputs(3008) <= not a;
    outputs(3009) <= b and not a;
    outputs(3010) <= not (a xor b);
    outputs(3011) <= a xor b;
    outputs(3012) <= a and not b;
    outputs(3013) <= a xor b;
    outputs(3014) <= not a or b;
    outputs(3015) <= not b;
    outputs(3016) <= not a;
    outputs(3017) <= a;
    outputs(3018) <= not b or a;
    outputs(3019) <= not (a and b);
    outputs(3020) <= not a or b;
    outputs(3021) <= b;
    outputs(3022) <= not b;
    outputs(3023) <= a xor b;
    outputs(3024) <= not a or b;
    outputs(3025) <= not (a xor b);
    outputs(3026) <= b;
    outputs(3027) <= a xor b;
    outputs(3028) <= a or b;
    outputs(3029) <= not a;
    outputs(3030) <= not a or b;
    outputs(3031) <= not (a or b);
    outputs(3032) <= a xor b;
    outputs(3033) <= b;
    outputs(3034) <= a xor b;
    outputs(3035) <= not b;
    outputs(3036) <= a or b;
    outputs(3037) <= not (a or b);
    outputs(3038) <= not (a xor b);
    outputs(3039) <= not (a or b);
    outputs(3040) <= a xor b;
    outputs(3041) <= b and not a;
    outputs(3042) <= a and not b;
    outputs(3043) <= not a;
    outputs(3044) <= not a;
    outputs(3045) <= a;
    outputs(3046) <= a or b;
    outputs(3047) <= a and not b;
    outputs(3048) <= not b;
    outputs(3049) <= not a;
    outputs(3050) <= not (a xor b);
    outputs(3051) <= not a;
    outputs(3052) <= b;
    outputs(3053) <= not a;
    outputs(3054) <= a xor b;
    outputs(3055) <= a xor b;
    outputs(3056) <= not b;
    outputs(3057) <= not b or a;
    outputs(3058) <= b and not a;
    outputs(3059) <= b and not a;
    outputs(3060) <= not (a xor b);
    outputs(3061) <= not a;
    outputs(3062) <= b;
    outputs(3063) <= not b;
    outputs(3064) <= not a;
    outputs(3065) <= b;
    outputs(3066) <= not a;
    outputs(3067) <= not (a xor b);
    outputs(3068) <= a xor b;
    outputs(3069) <= a and b;
    outputs(3070) <= b;
    outputs(3071) <= not (a or b);
    outputs(3072) <= not b;
    outputs(3073) <= not a;
    outputs(3074) <= b;
    outputs(3075) <= not b;
    outputs(3076) <= a xor b;
    outputs(3077) <= not (a or b);
    outputs(3078) <= not b;
    outputs(3079) <= not a;
    outputs(3080) <= not a;
    outputs(3081) <= not (a or b);
    outputs(3082) <= a and b;
    outputs(3083) <= not (a xor b);
    outputs(3084) <= b;
    outputs(3085) <= b;
    outputs(3086) <= a;
    outputs(3087) <= a and not b;
    outputs(3088) <= not (a xor b);
    outputs(3089) <= not b;
    outputs(3090) <= a;
    outputs(3091) <= not b or a;
    outputs(3092) <= not (a xor b);
    outputs(3093) <= a;
    outputs(3094) <= a xor b;
    outputs(3095) <= not (a xor b);
    outputs(3096) <= b;
    outputs(3097) <= a xor b;
    outputs(3098) <= not b;
    outputs(3099) <= a xor b;
    outputs(3100) <= not (a xor b);
    outputs(3101) <= not a;
    outputs(3102) <= not (a and b);
    outputs(3103) <= a and b;
    outputs(3104) <= a and not b;
    outputs(3105) <= not b or a;
    outputs(3106) <= not b;
    outputs(3107) <= a;
    outputs(3108) <= a;
    outputs(3109) <= a xor b;
    outputs(3110) <= b;
    outputs(3111) <= not b;
    outputs(3112) <= not b;
    outputs(3113) <= a xor b;
    outputs(3114) <= a;
    outputs(3115) <= not (a xor b);
    outputs(3116) <= a;
    outputs(3117) <= a;
    outputs(3118) <= a;
    outputs(3119) <= b;
    outputs(3120) <= not b;
    outputs(3121) <= b and not a;
    outputs(3122) <= not b;
    outputs(3123) <= a;
    outputs(3124) <= a and not b;
    outputs(3125) <= b;
    outputs(3126) <= a xor b;
    outputs(3127) <= a;
    outputs(3128) <= not (a xor b);
    outputs(3129) <= a and not b;
    outputs(3130) <= not b;
    outputs(3131) <= a xor b;
    outputs(3132) <= a;
    outputs(3133) <= b;
    outputs(3134) <= not a;
    outputs(3135) <= b and not a;
    outputs(3136) <= b and not a;
    outputs(3137) <= not b;
    outputs(3138) <= not (a xor b);
    outputs(3139) <= not (a xor b);
    outputs(3140) <= not b;
    outputs(3141) <= not a or b;
    outputs(3142) <= not (a or b);
    outputs(3143) <= a xor b;
    outputs(3144) <= a;
    outputs(3145) <= a xor b;
    outputs(3146) <= not b;
    outputs(3147) <= b and not a;
    outputs(3148) <= not b;
    outputs(3149) <= not a;
    outputs(3150) <= b;
    outputs(3151) <= not b;
    outputs(3152) <= b and not a;
    outputs(3153) <= not (a or b);
    outputs(3154) <= b and not a;
    outputs(3155) <= a and not b;
    outputs(3156) <= a and not b;
    outputs(3157) <= a;
    outputs(3158) <= not (a xor b);
    outputs(3159) <= a xor b;
    outputs(3160) <= not a or b;
    outputs(3161) <= a xor b;
    outputs(3162) <= a;
    outputs(3163) <= b;
    outputs(3164) <= a and b;
    outputs(3165) <= not (a or b);
    outputs(3166) <= not b;
    outputs(3167) <= a or b;
    outputs(3168) <= b;
    outputs(3169) <= b;
    outputs(3170) <= not (a or b);
    outputs(3171) <= not (a and b);
    outputs(3172) <= not (a and b);
    outputs(3173) <= a and b;
    outputs(3174) <= not (a xor b);
    outputs(3175) <= not a;
    outputs(3176) <= not (a or b);
    outputs(3177) <= not b;
    outputs(3178) <= not b;
    outputs(3179) <= a and b;
    outputs(3180) <= not a;
    outputs(3181) <= a or b;
    outputs(3182) <= not a;
    outputs(3183) <= b;
    outputs(3184) <= not a;
    outputs(3185) <= not a;
    outputs(3186) <= not b;
    outputs(3187) <= not b;
    outputs(3188) <= a;
    outputs(3189) <= not (a or b);
    outputs(3190) <= not b;
    outputs(3191) <= a and not b;
    outputs(3192) <= a;
    outputs(3193) <= b and not a;
    outputs(3194) <= not (a xor b);
    outputs(3195) <= not a;
    outputs(3196) <= a;
    outputs(3197) <= a xor b;
    outputs(3198) <= not (a and b);
    outputs(3199) <= not (a xor b);
    outputs(3200) <= not b;
    outputs(3201) <= not (a and b);
    outputs(3202) <= b and not a;
    outputs(3203) <= a;
    outputs(3204) <= b;
    outputs(3205) <= b;
    outputs(3206) <= b and not a;
    outputs(3207) <= not (a xor b);
    outputs(3208) <= not a;
    outputs(3209) <= a xor b;
    outputs(3210) <= b;
    outputs(3211) <= not (a or b);
    outputs(3212) <= a;
    outputs(3213) <= not a;
    outputs(3214) <= a;
    outputs(3215) <= b;
    outputs(3216) <= a and not b;
    outputs(3217) <= b;
    outputs(3218) <= not a;
    outputs(3219) <= a;
    outputs(3220) <= a;
    outputs(3221) <= not a;
    outputs(3222) <= not (a xor b);
    outputs(3223) <= a and not b;
    outputs(3224) <= not a;
    outputs(3225) <= a;
    outputs(3226) <= not (a xor b);
    outputs(3227) <= not a;
    outputs(3228) <= not a or b;
    outputs(3229) <= a;
    outputs(3230) <= not b or a;
    outputs(3231) <= a;
    outputs(3232) <= a and not b;
    outputs(3233) <= a;
    outputs(3234) <= not (a and b);
    outputs(3235) <= not a;
    outputs(3236) <= b;
    outputs(3237) <= not (a or b);
    outputs(3238) <= not (a or b);
    outputs(3239) <= not a;
    outputs(3240) <= not b or a;
    outputs(3241) <= a and not b;
    outputs(3242) <= not b;
    outputs(3243) <= not b;
    outputs(3244) <= not b;
    outputs(3245) <= not a or b;
    outputs(3246) <= a xor b;
    outputs(3247) <= a xor b;
    outputs(3248) <= a;
    outputs(3249) <= a xor b;
    outputs(3250) <= b;
    outputs(3251) <= b and not a;
    outputs(3252) <= not a;
    outputs(3253) <= b;
    outputs(3254) <= b;
    outputs(3255) <= not b;
    outputs(3256) <= not b or a;
    outputs(3257) <= a and b;
    outputs(3258) <= b;
    outputs(3259) <= not a;
    outputs(3260) <= not a or b;
    outputs(3261) <= a;
    outputs(3262) <= not b or a;
    outputs(3263) <= b;
    outputs(3264) <= b and not a;
    outputs(3265) <= b;
    outputs(3266) <= a xor b;
    outputs(3267) <= b and not a;
    outputs(3268) <= not b;
    outputs(3269) <= a;
    outputs(3270) <= b;
    outputs(3271) <= not (a or b);
    outputs(3272) <= not b;
    outputs(3273) <= a;
    outputs(3274) <= not a or b;
    outputs(3275) <= b;
    outputs(3276) <= a;
    outputs(3277) <= a xor b;
    outputs(3278) <= a xor b;
    outputs(3279) <= a xor b;
    outputs(3280) <= not b;
    outputs(3281) <= not a;
    outputs(3282) <= a and b;
    outputs(3283) <= a;
    outputs(3284) <= b and not a;
    outputs(3285) <= a or b;
    outputs(3286) <= a xor b;
    outputs(3287) <= b and not a;
    outputs(3288) <= not (a or b);
    outputs(3289) <= b;
    outputs(3290) <= a;
    outputs(3291) <= b;
    outputs(3292) <= a and not b;
    outputs(3293) <= not (a xor b);
    outputs(3294) <= a xor b;
    outputs(3295) <= b and not a;
    outputs(3296) <= b;
    outputs(3297) <= not a;
    outputs(3298) <= a and b;
    outputs(3299) <= b;
    outputs(3300) <= not b;
    outputs(3301) <= a or b;
    outputs(3302) <= not (a xor b);
    outputs(3303) <= a;
    outputs(3304) <= not b;
    outputs(3305) <= b;
    outputs(3306) <= not (a or b);
    outputs(3307) <= a xor b;
    outputs(3308) <= not (a xor b);
    outputs(3309) <= not a;
    outputs(3310) <= b;
    outputs(3311) <= a and b;
    outputs(3312) <= not a;
    outputs(3313) <= not (a and b);
    outputs(3314) <= not b;
    outputs(3315) <= a;
    outputs(3316) <= not (a and b);
    outputs(3317) <= b;
    outputs(3318) <= not a;
    outputs(3319) <= not b;
    outputs(3320) <= a;
    outputs(3321) <= a and not b;
    outputs(3322) <= a xor b;
    outputs(3323) <= a;
    outputs(3324) <= b and not a;
    outputs(3325) <= a xor b;
    outputs(3326) <= not (a or b);
    outputs(3327) <= not (a or b);
    outputs(3328) <= a xor b;
    outputs(3329) <= a and b;
    outputs(3330) <= not a;
    outputs(3331) <= not b or a;
    outputs(3332) <= a;
    outputs(3333) <= a and not b;
    outputs(3334) <= a;
    outputs(3335) <= a and b;
    outputs(3336) <= not (a or b);
    outputs(3337) <= not (a and b);
    outputs(3338) <= not b;
    outputs(3339) <= b;
    outputs(3340) <= b;
    outputs(3341) <= not a;
    outputs(3342) <= b;
    outputs(3343) <= b and not a;
    outputs(3344) <= not (a or b);
    outputs(3345) <= not a;
    outputs(3346) <= b;
    outputs(3347) <= not a;
    outputs(3348) <= not b;
    outputs(3349) <= a or b;
    outputs(3350) <= a xor b;
    outputs(3351) <= not b;
    outputs(3352) <= a;
    outputs(3353) <= b;
    outputs(3354) <= a and not b;
    outputs(3355) <= not (a xor b);
    outputs(3356) <= a xor b;
    outputs(3357) <= not a;
    outputs(3358) <= not a;
    outputs(3359) <= not b;
    outputs(3360) <= not (a or b);
    outputs(3361) <= a;
    outputs(3362) <= a;
    outputs(3363) <= not a or b;
    outputs(3364) <= a;
    outputs(3365) <= not b;
    outputs(3366) <= b;
    outputs(3367) <= not a;
    outputs(3368) <= a or b;
    outputs(3369) <= not a;
    outputs(3370) <= a and b;
    outputs(3371) <= b;
    outputs(3372) <= not a;
    outputs(3373) <= b;
    outputs(3374) <= not b;
    outputs(3375) <= b;
    outputs(3376) <= not b;
    outputs(3377) <= not a or b;
    outputs(3378) <= a and not b;
    outputs(3379) <= a and b;
    outputs(3380) <= not (a or b);
    outputs(3381) <= b;
    outputs(3382) <= a and not b;
    outputs(3383) <= a;
    outputs(3384) <= not b;
    outputs(3385) <= a and b;
    outputs(3386) <= not a;
    outputs(3387) <= not b or a;
    outputs(3388) <= a xor b;
    outputs(3389) <= not (a xor b);
    outputs(3390) <= a;
    outputs(3391) <= not b;
    outputs(3392) <= a and not b;
    outputs(3393) <= not b;
    outputs(3394) <= b and not a;
    outputs(3395) <= not (a xor b);
    outputs(3396) <= a xor b;
    outputs(3397) <= not (a and b);
    outputs(3398) <= not a;
    outputs(3399) <= b;
    outputs(3400) <= not b;
    outputs(3401) <= not a;
    outputs(3402) <= not b or a;
    outputs(3403) <= not a;
    outputs(3404) <= not (a or b);
    outputs(3405) <= not a;
    outputs(3406) <= a;
    outputs(3407) <= not (a xor b);
    outputs(3408) <= b;
    outputs(3409) <= a and not b;
    outputs(3410) <= not b or a;
    outputs(3411) <= a;
    outputs(3412) <= a or b;
    outputs(3413) <= a;
    outputs(3414) <= a and not b;
    outputs(3415) <= a xor b;
    outputs(3416) <= not (a xor b);
    outputs(3417) <= b and not a;
    outputs(3418) <= a;
    outputs(3419) <= not (a xor b);
    outputs(3420) <= a xor b;
    outputs(3421) <= a and b;
    outputs(3422) <= a xor b;
    outputs(3423) <= not a or b;
    outputs(3424) <= not b;
    outputs(3425) <= a and not b;
    outputs(3426) <= b;
    outputs(3427) <= b;
    outputs(3428) <= b;
    outputs(3429) <= a and not b;
    outputs(3430) <= not (a or b);
    outputs(3431) <= a;
    outputs(3432) <= a and b;
    outputs(3433) <= not b or a;
    outputs(3434) <= a;
    outputs(3435) <= a xor b;
    outputs(3436) <= not b;
    outputs(3437) <= b;
    outputs(3438) <= not a;
    outputs(3439) <= not (a or b);
    outputs(3440) <= not (a xor b);
    outputs(3441) <= not a;
    outputs(3442) <= a;
    outputs(3443) <= a;
    outputs(3444) <= a xor b;
    outputs(3445) <= not (a xor b);
    outputs(3446) <= a xor b;
    outputs(3447) <= not b;
    outputs(3448) <= not (a or b);
    outputs(3449) <= not (a or b);
    outputs(3450) <= not a;
    outputs(3451) <= a xor b;
    outputs(3452) <= not (a or b);
    outputs(3453) <= not a;
    outputs(3454) <= a and b;
    outputs(3455) <= not b;
    outputs(3456) <= not b;
    outputs(3457) <= not (a or b);
    outputs(3458) <= a xor b;
    outputs(3459) <= a and not b;
    outputs(3460) <= b and not a;
    outputs(3461) <= not (a xor b);
    outputs(3462) <= not (a xor b);
    outputs(3463) <= a;
    outputs(3464) <= b;
    outputs(3465) <= not (a and b);
    outputs(3466) <= not (a or b);
    outputs(3467) <= not b;
    outputs(3468) <= b;
    outputs(3469) <= not a or b;
    outputs(3470) <= not (a xor b);
    outputs(3471) <= not (a xor b);
    outputs(3472) <= a;
    outputs(3473) <= b;
    outputs(3474) <= not b or a;
    outputs(3475) <= not (a xor b);
    outputs(3476) <= a xor b;
    outputs(3477) <= a;
    outputs(3478) <= not a or b;
    outputs(3479) <= not (a xor b);
    outputs(3480) <= a xor b;
    outputs(3481) <= not b;
    outputs(3482) <= not (a xor b);
    outputs(3483) <= not b;
    outputs(3484) <= not b;
    outputs(3485) <= not a;
    outputs(3486) <= b;
    outputs(3487) <= a;
    outputs(3488) <= not a;
    outputs(3489) <= not (a xor b);
    outputs(3490) <= a;
    outputs(3491) <= not b;
    outputs(3492) <= not (a or b);
    outputs(3493) <= not a;
    outputs(3494) <= a;
    outputs(3495) <= b;
    outputs(3496) <= a and b;
    outputs(3497) <= not (a and b);
    outputs(3498) <= not a;
    outputs(3499) <= a;
    outputs(3500) <= not (a or b);
    outputs(3501) <= not b;
    outputs(3502) <= not b;
    outputs(3503) <= not b;
    outputs(3504) <= a xor b;
    outputs(3505) <= b;
    outputs(3506) <= a xor b;
    outputs(3507) <= not (a or b);
    outputs(3508) <= b;
    outputs(3509) <= a and not b;
    outputs(3510) <= a;
    outputs(3511) <= b;
    outputs(3512) <= a xor b;
    outputs(3513) <= not (a xor b);
    outputs(3514) <= b and not a;
    outputs(3515) <= b;
    outputs(3516) <= a xor b;
    outputs(3517) <= not a;
    outputs(3518) <= a xor b;
    outputs(3519) <= a;
    outputs(3520) <= b;
    outputs(3521) <= not b;
    outputs(3522) <= b;
    outputs(3523) <= a and b;
    outputs(3524) <= b;
    outputs(3525) <= not a;
    outputs(3526) <= a xor b;
    outputs(3527) <= a;
    outputs(3528) <= a;
    outputs(3529) <= not a;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= not (a xor b);
    outputs(3532) <= not b;
    outputs(3533) <= a;
    outputs(3534) <= not a;
    outputs(3535) <= not (a xor b);
    outputs(3536) <= not b or a;
    outputs(3537) <= not (a or b);
    outputs(3538) <= a xor b;
    outputs(3539) <= not b;
    outputs(3540) <= b;
    outputs(3541) <= b;
    outputs(3542) <= a and not b;
    outputs(3543) <= not b;
    outputs(3544) <= not b;
    outputs(3545) <= b;
    outputs(3546) <= a;
    outputs(3547) <= not (a or b);
    outputs(3548) <= b;
    outputs(3549) <= not a or b;
    outputs(3550) <= a xor b;
    outputs(3551) <= not b;
    outputs(3552) <= a xor b;
    outputs(3553) <= b;
    outputs(3554) <= a xor b;
    outputs(3555) <= not (a xor b);
    outputs(3556) <= a and b;
    outputs(3557) <= a;
    outputs(3558) <= b;
    outputs(3559) <= not b;
    outputs(3560) <= a;
    outputs(3561) <= b and not a;
    outputs(3562) <= a and b;
    outputs(3563) <= not a or b;
    outputs(3564) <= b and not a;
    outputs(3565) <= a and not b;
    outputs(3566) <= a xor b;
    outputs(3567) <= not b;
    outputs(3568) <= b;
    outputs(3569) <= not b;
    outputs(3570) <= a and not b;
    outputs(3571) <= a;
    outputs(3572) <= not b;
    outputs(3573) <= b;
    outputs(3574) <= a xor b;
    outputs(3575) <= a;
    outputs(3576) <= not (a xor b);
    outputs(3577) <= not a;
    outputs(3578) <= b;
    outputs(3579) <= not a;
    outputs(3580) <= a and not b;
    outputs(3581) <= b and not a;
    outputs(3582) <= b and not a;
    outputs(3583) <= not (a or b);
    outputs(3584) <= b;
    outputs(3585) <= a and b;
    outputs(3586) <= a and b;
    outputs(3587) <= not (a and b);
    outputs(3588) <= a;
    outputs(3589) <= not (a or b);
    outputs(3590) <= b and not a;
    outputs(3591) <= b;
    outputs(3592) <= not b;
    outputs(3593) <= not a;
    outputs(3594) <= not (a or b);
    outputs(3595) <= a and not b;
    outputs(3596) <= not a;
    outputs(3597) <= not (a or b);
    outputs(3598) <= a;
    outputs(3599) <= not (a or b);
    outputs(3600) <= not b;
    outputs(3601) <= b;
    outputs(3602) <= not (a or b);
    outputs(3603) <= a;
    outputs(3604) <= not b;
    outputs(3605) <= not a or b;
    outputs(3606) <= b and not a;
    outputs(3607) <= a and b;
    outputs(3608) <= not b;
    outputs(3609) <= not a or b;
    outputs(3610) <= not (a xor b);
    outputs(3611) <= not (a and b);
    outputs(3612) <= a and b;
    outputs(3613) <= not b;
    outputs(3614) <= b;
    outputs(3615) <= a and not b;
    outputs(3616) <= not (a or b);
    outputs(3617) <= a and b;
    outputs(3618) <= not a;
    outputs(3619) <= not a;
    outputs(3620) <= not a;
    outputs(3621) <= b;
    outputs(3622) <= a and b;
    outputs(3623) <= b;
    outputs(3624) <= a and not b;
    outputs(3625) <= not b;
    outputs(3626) <= a and b;
    outputs(3627) <= b;
    outputs(3628) <= not a or b;
    outputs(3629) <= a xor b;
    outputs(3630) <= a and not b;
    outputs(3631) <= b;
    outputs(3632) <= a and not b;
    outputs(3633) <= b;
    outputs(3634) <= b and not a;
    outputs(3635) <= b and not a;
    outputs(3636) <= a and b;
    outputs(3637) <= a xor b;
    outputs(3638) <= not a;
    outputs(3639) <= b and not a;
    outputs(3640) <= not b or a;
    outputs(3641) <= not (a or b);
    outputs(3642) <= not b;
    outputs(3643) <= a;
    outputs(3644) <= a and not b;
    outputs(3645) <= a and b;
    outputs(3646) <= a xor b;
    outputs(3647) <= not a;
    outputs(3648) <= not b;
    outputs(3649) <= not b or a;
    outputs(3650) <= not b;
    outputs(3651) <= a;
    outputs(3652) <= a;
    outputs(3653) <= a and b;
    outputs(3654) <= a xor b;
    outputs(3655) <= b;
    outputs(3656) <= not b;
    outputs(3657) <= b;
    outputs(3658) <= not a;
    outputs(3659) <= not (a or b);
    outputs(3660) <= a;
    outputs(3661) <= not (a or b);
    outputs(3662) <= a;
    outputs(3663) <= not a;
    outputs(3664) <= not a;
    outputs(3665) <= not (a or b);
    outputs(3666) <= not (a xor b);
    outputs(3667) <= b and not a;
    outputs(3668) <= not b;
    outputs(3669) <= not b;
    outputs(3670) <= a;
    outputs(3671) <= not a;
    outputs(3672) <= a;
    outputs(3673) <= a and not b;
    outputs(3674) <= b;
    outputs(3675) <= a and b;
    outputs(3676) <= not (a and b);
    outputs(3677) <= not a;
    outputs(3678) <= a and not b;
    outputs(3679) <= a;
    outputs(3680) <= a xor b;
    outputs(3681) <= a;
    outputs(3682) <= a;
    outputs(3683) <= a;
    outputs(3684) <= not b;
    outputs(3685) <= a;
    outputs(3686) <= a and b;
    outputs(3687) <= a;
    outputs(3688) <= not a;
    outputs(3689) <= a and b;
    outputs(3690) <= a;
    outputs(3691) <= a;
    outputs(3692) <= not b;
    outputs(3693) <= not (a xor b);
    outputs(3694) <= a;
    outputs(3695) <= a and b;
    outputs(3696) <= not (a or b);
    outputs(3697) <= a;
    outputs(3698) <= b and not a;
    outputs(3699) <= not b;
    outputs(3700) <= not (a or b);
    outputs(3701) <= b and not a;
    outputs(3702) <= a;
    outputs(3703) <= b and not a;
    outputs(3704) <= a and not b;
    outputs(3705) <= not (a xor b);
    outputs(3706) <= b;
    outputs(3707) <= a;
    outputs(3708) <= a xor b;
    outputs(3709) <= not b or a;
    outputs(3710) <= a and b;
    outputs(3711) <= not (a xor b);
    outputs(3712) <= not (a xor b);
    outputs(3713) <= not a;
    outputs(3714) <= a and b;
    outputs(3715) <= a or b;
    outputs(3716) <= b;
    outputs(3717) <= b;
    outputs(3718) <= a;
    outputs(3719) <= a and b;
    outputs(3720) <= b;
    outputs(3721) <= a;
    outputs(3722) <= b and not a;
    outputs(3723) <= a and b;
    outputs(3724) <= not (a or b);
    outputs(3725) <= b;
    outputs(3726) <= not b;
    outputs(3727) <= not (a or b);
    outputs(3728) <= a xor b;
    outputs(3729) <= a;
    outputs(3730) <= b and not a;
    outputs(3731) <= not (a and b);
    outputs(3732) <= b and not a;
    outputs(3733) <= not (a or b);
    outputs(3734) <= not a;
    outputs(3735) <= not b;
    outputs(3736) <= a and not b;
    outputs(3737) <= not (a or b);
    outputs(3738) <= not a or b;
    outputs(3739) <= b;
    outputs(3740) <= a;
    outputs(3741) <= b and not a;
    outputs(3742) <= not a;
    outputs(3743) <= not b;
    outputs(3744) <= not b;
    outputs(3745) <= not (a xor b);
    outputs(3746) <= not a or b;
    outputs(3747) <= not a;
    outputs(3748) <= not b;
    outputs(3749) <= b and not a;
    outputs(3750) <= a and b;
    outputs(3751) <= not (a or b);
    outputs(3752) <= not a;
    outputs(3753) <= b and not a;
    outputs(3754) <= b and not a;
    outputs(3755) <= a;
    outputs(3756) <= b;
    outputs(3757) <= not b;
    outputs(3758) <= not a;
    outputs(3759) <= not (a xor b);
    outputs(3760) <= not a;
    outputs(3761) <= b;
    outputs(3762) <= b;
    outputs(3763) <= not (a or b);
    outputs(3764) <= not (a or b);
    outputs(3765) <= not b;
    outputs(3766) <= not (a and b);
    outputs(3767) <= b and not a;
    outputs(3768) <= b;
    outputs(3769) <= not (a or b);
    outputs(3770) <= not (a and b);
    outputs(3771) <= a;
    outputs(3772) <= not a;
    outputs(3773) <= a and b;
    outputs(3774) <= not (a and b);
    outputs(3775) <= a and not b;
    outputs(3776) <= not a or b;
    outputs(3777) <= not b;
    outputs(3778) <= a xor b;
    outputs(3779) <= a and b;
    outputs(3780) <= not (a or b);
    outputs(3781) <= not a;
    outputs(3782) <= not (a or b);
    outputs(3783) <= b and not a;
    outputs(3784) <= not a;
    outputs(3785) <= not b;
    outputs(3786) <= not a or b;
    outputs(3787) <= not a;
    outputs(3788) <= a xor b;
    outputs(3789) <= not b;
    outputs(3790) <= a;
    outputs(3791) <= not a;
    outputs(3792) <= a;
    outputs(3793) <= not b or a;
    outputs(3794) <= b and not a;
    outputs(3795) <= not (a and b);
    outputs(3796) <= b;
    outputs(3797) <= not b;
    outputs(3798) <= a xor b;
    outputs(3799) <= not a;
    outputs(3800) <= a and not b;
    outputs(3801) <= not (a or b);
    outputs(3802) <= not (a xor b);
    outputs(3803) <= not b;
    outputs(3804) <= not (a xor b);
    outputs(3805) <= not (a and b);
    outputs(3806) <= not (a and b);
    outputs(3807) <= not b;
    outputs(3808) <= not (a and b);
    outputs(3809) <= a xor b;
    outputs(3810) <= not (a or b);
    outputs(3811) <= not b;
    outputs(3812) <= b and not a;
    outputs(3813) <= b;
    outputs(3814) <= a;
    outputs(3815) <= not a;
    outputs(3816) <= a and not b;
    outputs(3817) <= a and not b;
    outputs(3818) <= not a;
    outputs(3819) <= not (a xor b);
    outputs(3820) <= a and b;
    outputs(3821) <= not b;
    outputs(3822) <= a;
    outputs(3823) <= not b;
    outputs(3824) <= a xor b;
    outputs(3825) <= a and not b;
    outputs(3826) <= b;
    outputs(3827) <= not a;
    outputs(3828) <= a and b;
    outputs(3829) <= b;
    outputs(3830) <= b and not a;
    outputs(3831) <= not a;
    outputs(3832) <= a;
    outputs(3833) <= not b;
    outputs(3834) <= not (a or b);
    outputs(3835) <= b;
    outputs(3836) <= a and b;
    outputs(3837) <= a;
    outputs(3838) <= not a or b;
    outputs(3839) <= a and not b;
    outputs(3840) <= not b;
    outputs(3841) <= a or b;
    outputs(3842) <= not a;
    outputs(3843) <= b;
    outputs(3844) <= a;
    outputs(3845) <= a and b;
    outputs(3846) <= b;
    outputs(3847) <= a and not b;
    outputs(3848) <= b;
    outputs(3849) <= b and not a;
    outputs(3850) <= a;
    outputs(3851) <= not b or a;
    outputs(3852) <= not a;
    outputs(3853) <= a and b;
    outputs(3854) <= not a;
    outputs(3855) <= a and not b;
    outputs(3856) <= a and not b;
    outputs(3857) <= a and not b;
    outputs(3858) <= a and not b;
    outputs(3859) <= b and not a;
    outputs(3860) <= a and b;
    outputs(3861) <= not b;
    outputs(3862) <= a and b;
    outputs(3863) <= not (a xor b);
    outputs(3864) <= not a;
    outputs(3865) <= a xor b;
    outputs(3866) <= not a;
    outputs(3867) <= not (a xor b);
    outputs(3868) <= a and not b;
    outputs(3869) <= not b;
    outputs(3870) <= not a;
    outputs(3871) <= a and b;
    outputs(3872) <= b;
    outputs(3873) <= not (a or b);
    outputs(3874) <= not (a and b);
    outputs(3875) <= not b;
    outputs(3876) <= a and b;
    outputs(3877) <= a and b;
    outputs(3878) <= not a;
    outputs(3879) <= a and b;
    outputs(3880) <= not a;
    outputs(3881) <= not (a or b);
    outputs(3882) <= a;
    outputs(3883) <= a and not b;
    outputs(3884) <= a xor b;
    outputs(3885) <= not a;
    outputs(3886) <= not (a xor b);
    outputs(3887) <= not a;
    outputs(3888) <= b and not a;
    outputs(3889) <= a and not b;
    outputs(3890) <= not b;
    outputs(3891) <= not a;
    outputs(3892) <= a xor b;
    outputs(3893) <= a or b;
    outputs(3894) <= b and not a;
    outputs(3895) <= a xor b;
    outputs(3896) <= b and not a;
    outputs(3897) <= a xor b;
    outputs(3898) <= a xor b;
    outputs(3899) <= a and b;
    outputs(3900) <= not (a or b);
    outputs(3901) <= not a;
    outputs(3902) <= a and not b;
    outputs(3903) <= b;
    outputs(3904) <= not a;
    outputs(3905) <= b;
    outputs(3906) <= b and not a;
    outputs(3907) <= a and not b;
    outputs(3908) <= not (a xor b);
    outputs(3909) <= a or b;
    outputs(3910) <= a;
    outputs(3911) <= a;
    outputs(3912) <= a and not b;
    outputs(3913) <= not a or b;
    outputs(3914) <= a and not b;
    outputs(3915) <= not b;
    outputs(3916) <= a xor b;
    outputs(3917) <= not b;
    outputs(3918) <= a;
    outputs(3919) <= not (a or b);
    outputs(3920) <= not b or a;
    outputs(3921) <= not (a xor b);
    outputs(3922) <= not b;
    outputs(3923) <= not b;
    outputs(3924) <= a;
    outputs(3925) <= not (a xor b);
    outputs(3926) <= not (a xor b);
    outputs(3927) <= b;
    outputs(3928) <= not b;
    outputs(3929) <= a and not b;
    outputs(3930) <= a;
    outputs(3931) <= a and b;
    outputs(3932) <= not b;
    outputs(3933) <= a and b;
    outputs(3934) <= not a;
    outputs(3935) <= not b;
    outputs(3936) <= not a or b;
    outputs(3937) <= b;
    outputs(3938) <= not b;
    outputs(3939) <= a and not b;
    outputs(3940) <= a and b;
    outputs(3941) <= b and not a;
    outputs(3942) <= not b;
    outputs(3943) <= a;
    outputs(3944) <= a or b;
    outputs(3945) <= not a;
    outputs(3946) <= b;
    outputs(3947) <= not a;
    outputs(3948) <= a;
    outputs(3949) <= b;
    outputs(3950) <= a xor b;
    outputs(3951) <= b and not a;
    outputs(3952) <= not (a and b);
    outputs(3953) <= b and not a;
    outputs(3954) <= b;
    outputs(3955) <= b;
    outputs(3956) <= a or b;
    outputs(3957) <= not a or b;
    outputs(3958) <= b and not a;
    outputs(3959) <= a and not b;
    outputs(3960) <= b and not a;
    outputs(3961) <= a or b;
    outputs(3962) <= b;
    outputs(3963) <= a and b;
    outputs(3964) <= not b;
    outputs(3965) <= not (a xor b);
    outputs(3966) <= a and b;
    outputs(3967) <= b;
    outputs(3968) <= a and not b;
    outputs(3969) <= a xor b;
    outputs(3970) <= not a;
    outputs(3971) <= b and not a;
    outputs(3972) <= a;
    outputs(3973) <= a and b;
    outputs(3974) <= b;
    outputs(3975) <= a and not b;
    outputs(3976) <= a and not b;
    outputs(3977) <= b and not a;
    outputs(3978) <= a and b;
    outputs(3979) <= a and not b;
    outputs(3980) <= a;
    outputs(3981) <= a xor b;
    outputs(3982) <= a and not b;
    outputs(3983) <= not a;
    outputs(3984) <= not a;
    outputs(3985) <= a and b;
    outputs(3986) <= not (a or b);
    outputs(3987) <= a and b;
    outputs(3988) <= b and not a;
    outputs(3989) <= a and b;
    outputs(3990) <= not a;
    outputs(3991) <= a and b;
    outputs(3992) <= b;
    outputs(3993) <= a;
    outputs(3994) <= not (a xor b);
    outputs(3995) <= a or b;
    outputs(3996) <= not b;
    outputs(3997) <= not (a or b);
    outputs(3998) <= b;
    outputs(3999) <= not b or a;
    outputs(4000) <= a;
    outputs(4001) <= a and b;
    outputs(4002) <= not (a or b);
    outputs(4003) <= not (a xor b);
    outputs(4004) <= not (a or b);
    outputs(4005) <= b and not a;
    outputs(4006) <= a and not b;
    outputs(4007) <= a and not b;
    outputs(4008) <= not b;
    outputs(4009) <= not (a or b);
    outputs(4010) <= b and not a;
    outputs(4011) <= a and not b;
    outputs(4012) <= b and not a;
    outputs(4013) <= not a;
    outputs(4014) <= a and b;
    outputs(4015) <= not (a xor b);
    outputs(4016) <= not b;
    outputs(4017) <= a and b;
    outputs(4018) <= a or b;
    outputs(4019) <= a or b;
    outputs(4020) <= a;
    outputs(4021) <= not (a xor b);
    outputs(4022) <= a and b;
    outputs(4023) <= a;
    outputs(4024) <= not a;
    outputs(4025) <= a and not b;
    outputs(4026) <= a and not b;
    outputs(4027) <= a and not b;
    outputs(4028) <= not a;
    outputs(4029) <= not b;
    outputs(4030) <= a and b;
    outputs(4031) <= a and not b;
    outputs(4032) <= not b;
    outputs(4033) <= not b;
    outputs(4034) <= a;
    outputs(4035) <= a and b;
    outputs(4036) <= a;
    outputs(4037) <= a;
    outputs(4038) <= a or b;
    outputs(4039) <= a;
    outputs(4040) <= b and not a;
    outputs(4041) <= b;
    outputs(4042) <= not a;
    outputs(4043) <= b and not a;
    outputs(4044) <= not b;
    outputs(4045) <= a;
    outputs(4046) <= not b or a;
    outputs(4047) <= a;
    outputs(4048) <= not (a xor b);
    outputs(4049) <= a;
    outputs(4050) <= not (a or b);
    outputs(4051) <= not (a or b);
    outputs(4052) <= a;
    outputs(4053) <= not a;
    outputs(4054) <= b;
    outputs(4055) <= a;
    outputs(4056) <= not a;
    outputs(4057) <= not (a xor b);
    outputs(4058) <= b;
    outputs(4059) <= a xor b;
    outputs(4060) <= not b;
    outputs(4061) <= b;
    outputs(4062) <= b and not a;
    outputs(4063) <= b and not a;
    outputs(4064) <= not a;
    outputs(4065) <= not b;
    outputs(4066) <= a;
    outputs(4067) <= a or b;
    outputs(4068) <= not a;
    outputs(4069) <= a;
    outputs(4070) <= not a;
    outputs(4071) <= b;
    outputs(4072) <= b and not a;
    outputs(4073) <= not (a xor b);
    outputs(4074) <= not (a or b);
    outputs(4075) <= not (a or b);
    outputs(4076) <= not (a and b);
    outputs(4077) <= b and not a;
    outputs(4078) <= b and not a;
    outputs(4079) <= b and not a;
    outputs(4080) <= not a;
    outputs(4081) <= not (a or b);
    outputs(4082) <= a and not b;
    outputs(4083) <= a xor b;
    outputs(4084) <= not a or b;
    outputs(4085) <= not (a or b);
    outputs(4086) <= a and b;
    outputs(4087) <= a and b;
    outputs(4088) <= not b;
    outputs(4089) <= b and not a;
    outputs(4090) <= not a;
    outputs(4091) <= b and not a;
    outputs(4092) <= not b;
    outputs(4093) <= not (a and b);
    outputs(4094) <= a xor b;
    outputs(4095) <= a xor b;
    outputs(4096) <= a;
    outputs(4097) <= a;
    outputs(4098) <= not a;
    outputs(4099) <= not b;
    outputs(4100) <= not (a xor b);
    outputs(4101) <= a and not b;
    outputs(4102) <= not a;
    outputs(4103) <= not b;
    outputs(4104) <= not a;
    outputs(4105) <= not a;
    outputs(4106) <= a;
    outputs(4107) <= a;
    outputs(4108) <= not a;
    outputs(4109) <= not b;
    outputs(4110) <= not a;
    outputs(4111) <= not a;
    outputs(4112) <= b;
    outputs(4113) <= not a;
    outputs(4114) <= not b;
    outputs(4115) <= not (a xor b);
    outputs(4116) <= a;
    outputs(4117) <= a or b;
    outputs(4118) <= not b or a;
    outputs(4119) <= a;
    outputs(4120) <= not a or b;
    outputs(4121) <= a;
    outputs(4122) <= b and not a;
    outputs(4123) <= a or b;
    outputs(4124) <= not b;
    outputs(4125) <= not b or a;
    outputs(4126) <= not b;
    outputs(4127) <= not b;
    outputs(4128) <= not (a xor b);
    outputs(4129) <= b;
    outputs(4130) <= b;
    outputs(4131) <= a;
    outputs(4132) <= a;
    outputs(4133) <= a xor b;
    outputs(4134) <= not b;
    outputs(4135) <= not (a xor b);
    outputs(4136) <= not a or b;
    outputs(4137) <= a;
    outputs(4138) <= a xor b;
    outputs(4139) <= b and not a;
    outputs(4140) <= not (a or b);
    outputs(4141) <= not a or b;
    outputs(4142) <= a;
    outputs(4143) <= b;
    outputs(4144) <= b and not a;
    outputs(4145) <= a and b;
    outputs(4146) <= not b;
    outputs(4147) <= a xor b;
    outputs(4148) <= a or b;
    outputs(4149) <= not a;
    outputs(4150) <= a or b;
    outputs(4151) <= a and b;
    outputs(4152) <= b;
    outputs(4153) <= not b;
    outputs(4154) <= not b;
    outputs(4155) <= not b;
    outputs(4156) <= b and not a;
    outputs(4157) <= b;
    outputs(4158) <= not b;
    outputs(4159) <= not a or b;
    outputs(4160) <= not b;
    outputs(4161) <= not a;
    outputs(4162) <= a and b;
    outputs(4163) <= a xor b;
    outputs(4164) <= a xor b;
    outputs(4165) <= not a;
    outputs(4166) <= b;
    outputs(4167) <= not (a or b);
    outputs(4168) <= not a;
    outputs(4169) <= a;
    outputs(4170) <= a xor b;
    outputs(4171) <= a and not b;
    outputs(4172) <= not a;
    outputs(4173) <= b and not a;
    outputs(4174) <= b;
    outputs(4175) <= not b;
    outputs(4176) <= not (a xor b);
    outputs(4177) <= not b;
    outputs(4178) <= not b;
    outputs(4179) <= not b;
    outputs(4180) <= not b;
    outputs(4181) <= a xor b;
    outputs(4182) <= a and not b;
    outputs(4183) <= a and b;
    outputs(4184) <= not a or b;
    outputs(4185) <= not (a xor b);
    outputs(4186) <= b and not a;
    outputs(4187) <= a or b;
    outputs(4188) <= not b;
    outputs(4189) <= b;
    outputs(4190) <= a xor b;
    outputs(4191) <= a;
    outputs(4192) <= not (a xor b);
    outputs(4193) <= not (a xor b);
    outputs(4194) <= b;
    outputs(4195) <= b and not a;
    outputs(4196) <= not (a or b);
    outputs(4197) <= a;
    outputs(4198) <= a xor b;
    outputs(4199) <= not b or a;
    outputs(4200) <= not b;
    outputs(4201) <= not b;
    outputs(4202) <= a;
    outputs(4203) <= a or b;
    outputs(4204) <= not a;
    outputs(4205) <= not a;
    outputs(4206) <= b and not a;
    outputs(4207) <= not a or b;
    outputs(4208) <= a;
    outputs(4209) <= b and not a;
    outputs(4210) <= a;
    outputs(4211) <= a and b;
    outputs(4212) <= a or b;
    outputs(4213) <= a xor b;
    outputs(4214) <= not a or b;
    outputs(4215) <= b;
    outputs(4216) <= not (a xor b);
    outputs(4217) <= not a;
    outputs(4218) <= a;
    outputs(4219) <= a or b;
    outputs(4220) <= not a;
    outputs(4221) <= b;
    outputs(4222) <= b and not a;
    outputs(4223) <= b;
    outputs(4224) <= not a;
    outputs(4225) <= not b;
    outputs(4226) <= a xor b;
    outputs(4227) <= not b;
    outputs(4228) <= a or b;
    outputs(4229) <= not a;
    outputs(4230) <= a and not b;
    outputs(4231) <= a and b;
    outputs(4232) <= not a;
    outputs(4233) <= a xor b;
    outputs(4234) <= a xor b;
    outputs(4235) <= not b;
    outputs(4236) <= a xor b;
    outputs(4237) <= not a;
    outputs(4238) <= b;
    outputs(4239) <= not a or b;
    outputs(4240) <= not b;
    outputs(4241) <= a and not b;
    outputs(4242) <= not (a xor b);
    outputs(4243) <= b and not a;
    outputs(4244) <= a;
    outputs(4245) <= not b;
    outputs(4246) <= not b or a;
    outputs(4247) <= not a;
    outputs(4248) <= b;
    outputs(4249) <= a and b;
    outputs(4250) <= a and b;
    outputs(4251) <= not (a xor b);
    outputs(4252) <= a;
    outputs(4253) <= not a;
    outputs(4254) <= b;
    outputs(4255) <= b;
    outputs(4256) <= not b or a;
    outputs(4257) <= a xor b;
    outputs(4258) <= not (a xor b);
    outputs(4259) <= not (a xor b);
    outputs(4260) <= not b;
    outputs(4261) <= not a;
    outputs(4262) <= not b or a;
    outputs(4263) <= not b;
    outputs(4264) <= a;
    outputs(4265) <= b and not a;
    outputs(4266) <= not a;
    outputs(4267) <= a xor b;
    outputs(4268) <= b;
    outputs(4269) <= a xor b;
    outputs(4270) <= b;
    outputs(4271) <= b;
    outputs(4272) <= a xor b;
    outputs(4273) <= not (a and b);
    outputs(4274) <= not a;
    outputs(4275) <= not a;
    outputs(4276) <= a;
    outputs(4277) <= not b;
    outputs(4278) <= a;
    outputs(4279) <= not b;
    outputs(4280) <= b;
    outputs(4281) <= a xor b;
    outputs(4282) <= not a;
    outputs(4283) <= not b;
    outputs(4284) <= not b;
    outputs(4285) <= not b;
    outputs(4286) <= b and not a;
    outputs(4287) <= a and b;
    outputs(4288) <= a;
    outputs(4289) <= not (a and b);
    outputs(4290) <= not a;
    outputs(4291) <= b;
    outputs(4292) <= not (a xor b);
    outputs(4293) <= a and b;
    outputs(4294) <= b and not a;
    outputs(4295) <= b and not a;
    outputs(4296) <= not (a and b);
    outputs(4297) <= a xor b;
    outputs(4298) <= not (a xor b);
    outputs(4299) <= b;
    outputs(4300) <= a;
    outputs(4301) <= b;
    outputs(4302) <= not a or b;
    outputs(4303) <= a and not b;
    outputs(4304) <= not (a xor b);
    outputs(4305) <= not a;
    outputs(4306) <= b;
    outputs(4307) <= a;
    outputs(4308) <= not (a xor b);
    outputs(4309) <= not (a or b);
    outputs(4310) <= b;
    outputs(4311) <= a xor b;
    outputs(4312) <= a;
    outputs(4313) <= not (a xor b);
    outputs(4314) <= b;
    outputs(4315) <= b;
    outputs(4316) <= not (a xor b);
    outputs(4317) <= not (a xor b);
    outputs(4318) <= a and not b;
    outputs(4319) <= b and not a;
    outputs(4320) <= not a;
    outputs(4321) <= not a or b;
    outputs(4322) <= b;
    outputs(4323) <= b;
    outputs(4324) <= not (a or b);
    outputs(4325) <= not a or b;
    outputs(4326) <= not b;
    outputs(4327) <= not (a xor b);
    outputs(4328) <= not (a and b);
    outputs(4329) <= a;
    outputs(4330) <= a xor b;
    outputs(4331) <= not b;
    outputs(4332) <= a;
    outputs(4333) <= not (a xor b);
    outputs(4334) <= a xor b;
    outputs(4335) <= not a;
    outputs(4336) <= b;
    outputs(4337) <= a and b;
    outputs(4338) <= not (a xor b);
    outputs(4339) <= not a or b;
    outputs(4340) <= a xor b;
    outputs(4341) <= a;
    outputs(4342) <= a xor b;
    outputs(4343) <= not a;
    outputs(4344) <= a xor b;
    outputs(4345) <= not (a xor b);
    outputs(4346) <= a and not b;
    outputs(4347) <= not a;
    outputs(4348) <= not a;
    outputs(4349) <= not (a or b);
    outputs(4350) <= not b or a;
    outputs(4351) <= a and b;
    outputs(4352) <= not b;
    outputs(4353) <= not a;
    outputs(4354) <= not a;
    outputs(4355) <= a;
    outputs(4356) <= not a;
    outputs(4357) <= not b;
    outputs(4358) <= a and b;
    outputs(4359) <= not (a or b);
    outputs(4360) <= a xor b;
    outputs(4361) <= not b;
    outputs(4362) <= a;
    outputs(4363) <= a xor b;
    outputs(4364) <= not b or a;
    outputs(4365) <= a or b;
    outputs(4366) <= b;
    outputs(4367) <= not a;
    outputs(4368) <= b and not a;
    outputs(4369) <= b;
    outputs(4370) <= not a;
    outputs(4371) <= not b or a;
    outputs(4372) <= not a;
    outputs(4373) <= a and not b;
    outputs(4374) <= b;
    outputs(4375) <= not (a xor b);
    outputs(4376) <= a xor b;
    outputs(4377) <= a xor b;
    outputs(4378) <= not (a xor b);
    outputs(4379) <= not a;
    outputs(4380) <= not b or a;
    outputs(4381) <= not b;
    outputs(4382) <= not b;
    outputs(4383) <= not b;
    outputs(4384) <= not b;
    outputs(4385) <= a or b;
    outputs(4386) <= a;
    outputs(4387) <= not b or a;
    outputs(4388) <= a;
    outputs(4389) <= not (a xor b);
    outputs(4390) <= a or b;
    outputs(4391) <= a;
    outputs(4392) <= a;
    outputs(4393) <= a and b;
    outputs(4394) <= a xor b;
    outputs(4395) <= b and not a;
    outputs(4396) <= b and not a;
    outputs(4397) <= b and not a;
    outputs(4398) <= not (a xor b);
    outputs(4399) <= not b;
    outputs(4400) <= a xor b;
    outputs(4401) <= a and b;
    outputs(4402) <= b;
    outputs(4403) <= not b or a;
    outputs(4404) <= not (a or b);
    outputs(4405) <= a xor b;
    outputs(4406) <= not a;
    outputs(4407) <= a;
    outputs(4408) <= b;
    outputs(4409) <= not b or a;
    outputs(4410) <= not a;
    outputs(4411) <= not (a xor b);
    outputs(4412) <= not a;
    outputs(4413) <= a and not b;
    outputs(4414) <= not (a or b);
    outputs(4415) <= not (a and b);
    outputs(4416) <= a or b;
    outputs(4417) <= not a;
    outputs(4418) <= not (a xor b);
    outputs(4419) <= not b;
    outputs(4420) <= not (a xor b);
    outputs(4421) <= not b or a;
    outputs(4422) <= not b;
    outputs(4423) <= not b;
    outputs(4424) <= a and not b;
    outputs(4425) <= not b;
    outputs(4426) <= not b;
    outputs(4427) <= not (a xor b);
    outputs(4428) <= not (a xor b);
    outputs(4429) <= not (a or b);
    outputs(4430) <= a and not b;
    outputs(4431) <= a and not b;
    outputs(4432) <= a and not b;
    outputs(4433) <= b;
    outputs(4434) <= not a;
    outputs(4435) <= not b or a;
    outputs(4436) <= a xor b;
    outputs(4437) <= a;
    outputs(4438) <= not b or a;
    outputs(4439) <= b;
    outputs(4440) <= a xor b;
    outputs(4441) <= b;
    outputs(4442) <= b;
    outputs(4443) <= a;
    outputs(4444) <= a and not b;
    outputs(4445) <= not a;
    outputs(4446) <= a;
    outputs(4447) <= b and not a;
    outputs(4448) <= not a;
    outputs(4449) <= b;
    outputs(4450) <= a or b;
    outputs(4451) <= not (a or b);
    outputs(4452) <= not a;
    outputs(4453) <= a and not b;
    outputs(4454) <= not b;
    outputs(4455) <= b;
    outputs(4456) <= a xor b;
    outputs(4457) <= not b;
    outputs(4458) <= b;
    outputs(4459) <= a;
    outputs(4460) <= not b;
    outputs(4461) <= b;
    outputs(4462) <= b and not a;
    outputs(4463) <= a;
    outputs(4464) <= not (a xor b);
    outputs(4465) <= not a;
    outputs(4466) <= a;
    outputs(4467) <= b;
    outputs(4468) <= not (a or b);
    outputs(4469) <= a xor b;
    outputs(4470) <= not b;
    outputs(4471) <= not a;
    outputs(4472) <= not a;
    outputs(4473) <= a xor b;
    outputs(4474) <= a xor b;
    outputs(4475) <= a xor b;
    outputs(4476) <= not (a xor b);
    outputs(4477) <= not a;
    outputs(4478) <= b;
    outputs(4479) <= a xor b;
    outputs(4480) <= not b;
    outputs(4481) <= not b;
    outputs(4482) <= b;
    outputs(4483) <= not (a xor b);
    outputs(4484) <= not b;
    outputs(4485) <= not b;
    outputs(4486) <= b;
    outputs(4487) <= not a;
    outputs(4488) <= not (a xor b);
    outputs(4489) <= b and not a;
    outputs(4490) <= a or b;
    outputs(4491) <= a or b;
    outputs(4492) <= a or b;
    outputs(4493) <= a;
    outputs(4494) <= not a;
    outputs(4495) <= a xor b;
    outputs(4496) <= not (a or b);
    outputs(4497) <= b;
    outputs(4498) <= not b;
    outputs(4499) <= not a or b;
    outputs(4500) <= not b;
    outputs(4501) <= b and not a;
    outputs(4502) <= a;
    outputs(4503) <= a and not b;
    outputs(4504) <= not a;
    outputs(4505) <= a and not b;
    outputs(4506) <= not a or b;
    outputs(4507) <= b;
    outputs(4508) <= b;
    outputs(4509) <= not a;
    outputs(4510) <= a xor b;
    outputs(4511) <= a and b;
    outputs(4512) <= not (a xor b);
    outputs(4513) <= b;
    outputs(4514) <= a;
    outputs(4515) <= a xor b;
    outputs(4516) <= not (a xor b);
    outputs(4517) <= not a;
    outputs(4518) <= not b;
    outputs(4519) <= a or b;
    outputs(4520) <= not b;
    outputs(4521) <= a and not b;
    outputs(4522) <= b and not a;
    outputs(4523) <= b;
    outputs(4524) <= not (a xor b);
    outputs(4525) <= b and not a;
    outputs(4526) <= not a or b;
    outputs(4527) <= not a or b;
    outputs(4528) <= a and not b;
    outputs(4529) <= not (a xor b);
    outputs(4530) <= a xor b;
    outputs(4531) <= b;
    outputs(4532) <= b and not a;
    outputs(4533) <= b;
    outputs(4534) <= not a;
    outputs(4535) <= not b or a;
    outputs(4536) <= a xor b;
    outputs(4537) <= b;
    outputs(4538) <= a or b;
    outputs(4539) <= a and not b;
    outputs(4540) <= not b;
    outputs(4541) <= not b or a;
    outputs(4542) <= a xor b;
    outputs(4543) <= a and b;
    outputs(4544) <= not a;
    outputs(4545) <= a;
    outputs(4546) <= not (a xor b);
    outputs(4547) <= not b;
    outputs(4548) <= b;
    outputs(4549) <= a;
    outputs(4550) <= a and not b;
    outputs(4551) <= a;
    outputs(4552) <= not (a xor b);
    outputs(4553) <= a xor b;
    outputs(4554) <= not (a xor b);
    outputs(4555) <= not b;
    outputs(4556) <= not a;
    outputs(4557) <= a;
    outputs(4558) <= not (a and b);
    outputs(4559) <= not (a and b);
    outputs(4560) <= b;
    outputs(4561) <= not (a and b);
    outputs(4562) <= not a;
    outputs(4563) <= b;
    outputs(4564) <= not (a xor b);
    outputs(4565) <= not a;
    outputs(4566) <= a;
    outputs(4567) <= b;
    outputs(4568) <= not (a xor b);
    outputs(4569) <= a xor b;
    outputs(4570) <= a xor b;
    outputs(4571) <= a;
    outputs(4572) <= not (a xor b);
    outputs(4573) <= not (a xor b);
    outputs(4574) <= not b or a;
    outputs(4575) <= not (a xor b);
    outputs(4576) <= a or b;
    outputs(4577) <= a;
    outputs(4578) <= not a;
    outputs(4579) <= b;
    outputs(4580) <= not b;
    outputs(4581) <= not (a and b);
    outputs(4582) <= not a;
    outputs(4583) <= a;
    outputs(4584) <= not a;
    outputs(4585) <= not b;
    outputs(4586) <= not a;
    outputs(4587) <= a and not b;
    outputs(4588) <= not (a xor b);
    outputs(4589) <= a xor b;
    outputs(4590) <= not a;
    outputs(4591) <= not a;
    outputs(4592) <= b;
    outputs(4593) <= not a;
    outputs(4594) <= b;
    outputs(4595) <= not b;
    outputs(4596) <= a xor b;
    outputs(4597) <= a or b;
    outputs(4598) <= not b;
    outputs(4599) <= not a;
    outputs(4600) <= b;
    outputs(4601) <= a xor b;
    outputs(4602) <= not (a xor b);
    outputs(4603) <= a or b;
    outputs(4604) <= not a;
    outputs(4605) <= a and b;
    outputs(4606) <= a xor b;
    outputs(4607) <= not a;
    outputs(4608) <= not b;
    outputs(4609) <= a and not b;
    outputs(4610) <= not a or b;
    outputs(4611) <= not b or a;
    outputs(4612) <= not (a xor b);
    outputs(4613) <= not a;
    outputs(4614) <= not (a or b);
    outputs(4615) <= a xor b;
    outputs(4616) <= not a;
    outputs(4617) <= not (a or b);
    outputs(4618) <= b and not a;
    outputs(4619) <= not b;
    outputs(4620) <= not (a xor b);
    outputs(4621) <= a and b;
    outputs(4622) <= a;
    outputs(4623) <= a xor b;
    outputs(4624) <= a;
    outputs(4625) <= not b;
    outputs(4626) <= a xor b;
    outputs(4627) <= a;
    outputs(4628) <= b and not a;
    outputs(4629) <= a;
    outputs(4630) <= not (a xor b);
    outputs(4631) <= a or b;
    outputs(4632) <= b and not a;
    outputs(4633) <= a;
    outputs(4634) <= a and not b;
    outputs(4635) <= not b;
    outputs(4636) <= a xor b;
    outputs(4637) <= b and not a;
    outputs(4638) <= not b;
    outputs(4639) <= a xor b;
    outputs(4640) <= not (a or b);
    outputs(4641) <= b;
    outputs(4642) <= not b or a;
    outputs(4643) <= not a;
    outputs(4644) <= not (a xor b);
    outputs(4645) <= a;
    outputs(4646) <= not b or a;
    outputs(4647) <= a and not b;
    outputs(4648) <= not b;
    outputs(4649) <= b;
    outputs(4650) <= b;
    outputs(4651) <= not (a xor b);
    outputs(4652) <= not a or b;
    outputs(4653) <= not (a xor b);
    outputs(4654) <= a or b;
    outputs(4655) <= a and not b;
    outputs(4656) <= not a;
    outputs(4657) <= a and b;
    outputs(4658) <= a and b;
    outputs(4659) <= not a;
    outputs(4660) <= b;
    outputs(4661) <= a;
    outputs(4662) <= a xor b;
    outputs(4663) <= b;
    outputs(4664) <= not b;
    outputs(4665) <= not a;
    outputs(4666) <= not a or b;
    outputs(4667) <= b;
    outputs(4668) <= a and b;
    outputs(4669) <= not b;
    outputs(4670) <= a and not b;
    outputs(4671) <= a;
    outputs(4672) <= a xor b;
    outputs(4673) <= a and b;
    outputs(4674) <= not a;
    outputs(4675) <= a and b;
    outputs(4676) <= not b or a;
    outputs(4677) <= not b;
    outputs(4678) <= not (a or b);
    outputs(4679) <= not b;
    outputs(4680) <= a xor b;
    outputs(4681) <= not b or a;
    outputs(4682) <= a xor b;
    outputs(4683) <= not b;
    outputs(4684) <= not b;
    outputs(4685) <= b and not a;
    outputs(4686) <= a or b;
    outputs(4687) <= not a or b;
    outputs(4688) <= not a or b;
    outputs(4689) <= not b or a;
    outputs(4690) <= a xor b;
    outputs(4691) <= not a;
    outputs(4692) <= not a;
    outputs(4693) <= b and not a;
    outputs(4694) <= not b;
    outputs(4695) <= a xor b;
    outputs(4696) <= not a;
    outputs(4697) <= not a;
    outputs(4698) <= b;
    outputs(4699) <= a xor b;
    outputs(4700) <= a xor b;
    outputs(4701) <= not (a or b);
    outputs(4702) <= a and b;
    outputs(4703) <= a;
    outputs(4704) <= not (a xor b);
    outputs(4705) <= not (a xor b);
    outputs(4706) <= not a or b;
    outputs(4707) <= a and not b;
    outputs(4708) <= b;
    outputs(4709) <= not a or b;
    outputs(4710) <= not (a or b);
    outputs(4711) <= not a;
    outputs(4712) <= not (a or b);
    outputs(4713) <= b;
    outputs(4714) <= b;
    outputs(4715) <= not b or a;
    outputs(4716) <= b;
    outputs(4717) <= a xor b;
    outputs(4718) <= a;
    outputs(4719) <= a and b;
    outputs(4720) <= a;
    outputs(4721) <= a and not b;
    outputs(4722) <= a;
    outputs(4723) <= b;
    outputs(4724) <= a;
    outputs(4725) <= not b;
    outputs(4726) <= b and not a;
    outputs(4727) <= b;
    outputs(4728) <= not b;
    outputs(4729) <= not b;
    outputs(4730) <= a;
    outputs(4731) <= a;
    outputs(4732) <= a;
    outputs(4733) <= a;
    outputs(4734) <= b;
    outputs(4735) <= not b;
    outputs(4736) <= a xor b;
    outputs(4737) <= b and not a;
    outputs(4738) <= a;
    outputs(4739) <= not b or a;
    outputs(4740) <= a and b;
    outputs(4741) <= not a;
    outputs(4742) <= a and b;
    outputs(4743) <= a xor b;
    outputs(4744) <= b and not a;
    outputs(4745) <= not b;
    outputs(4746) <= a;
    outputs(4747) <= a;
    outputs(4748) <= b;
    outputs(4749) <= not (a and b);
    outputs(4750) <= not (a xor b);
    outputs(4751) <= not (a xor b);
    outputs(4752) <= a and b;
    outputs(4753) <= b;
    outputs(4754) <= a and b;
    outputs(4755) <= not b;
    outputs(4756) <= not (a xor b);
    outputs(4757) <= a;
    outputs(4758) <= b;
    outputs(4759) <= not a;
    outputs(4760) <= not (a or b);
    outputs(4761) <= b;
    outputs(4762) <= a;
    outputs(4763) <= not b;
    outputs(4764) <= not b;
    outputs(4765) <= a xor b;
    outputs(4766) <= b;
    outputs(4767) <= not (a xor b);
    outputs(4768) <= not a;
    outputs(4769) <= not a;
    outputs(4770) <= b;
    outputs(4771) <= b and not a;
    outputs(4772) <= not b;
    outputs(4773) <= b;
    outputs(4774) <= a;
    outputs(4775) <= a;
    outputs(4776) <= a or b;
    outputs(4777) <= a xor b;
    outputs(4778) <= b;
    outputs(4779) <= not (a xor b);
    outputs(4780) <= not b;
    outputs(4781) <= a xor b;
    outputs(4782) <= a xor b;
    outputs(4783) <= not b;
    outputs(4784) <= not a;
    outputs(4785) <= a and b;
    outputs(4786) <= not b;
    outputs(4787) <= not a;
    outputs(4788) <= a;
    outputs(4789) <= not (a xor b);
    outputs(4790) <= not (a or b);
    outputs(4791) <= a and not b;
    outputs(4792) <= not a;
    outputs(4793) <= a xor b;
    outputs(4794) <= not b;
    outputs(4795) <= a and b;
    outputs(4796) <= not a;
    outputs(4797) <= b;
    outputs(4798) <= a or b;
    outputs(4799) <= b;
    outputs(4800) <= not (a xor b);
    outputs(4801) <= a;
    outputs(4802) <= not (a or b);
    outputs(4803) <= not b or a;
    outputs(4804) <= not (a xor b);
    outputs(4805) <= not b;
    outputs(4806) <= not a or b;
    outputs(4807) <= a xor b;
    outputs(4808) <= a xor b;
    outputs(4809) <= b and not a;
    outputs(4810) <= not b;
    outputs(4811) <= not b;
    outputs(4812) <= a;
    outputs(4813) <= a and not b;
    outputs(4814) <= not a;
    outputs(4815) <= not a;
    outputs(4816) <= not b;
    outputs(4817) <= b;
    outputs(4818) <= a and b;
    outputs(4819) <= a;
    outputs(4820) <= not a;
    outputs(4821) <= not a;
    outputs(4822) <= not a or b;
    outputs(4823) <= a;
    outputs(4824) <= b;
    outputs(4825) <= a;
    outputs(4826) <= a;
    outputs(4827) <= a;
    outputs(4828) <= b and not a;
    outputs(4829) <= not (a or b);
    outputs(4830) <= not a;
    outputs(4831) <= not b;
    outputs(4832) <= a xor b;
    outputs(4833) <= not (a or b);
    outputs(4834) <= a;
    outputs(4835) <= a and b;
    outputs(4836) <= a;
    outputs(4837) <= not b;
    outputs(4838) <= a;
    outputs(4839) <= not a or b;
    outputs(4840) <= a and b;
    outputs(4841) <= a;
    outputs(4842) <= not (a xor b);
    outputs(4843) <= a;
    outputs(4844) <= not a;
    outputs(4845) <= not a;
    outputs(4846) <= a xor b;
    outputs(4847) <= b and not a;
    outputs(4848) <= b;
    outputs(4849) <= a and not b;
    outputs(4850) <= not a;
    outputs(4851) <= a and b;
    outputs(4852) <= a and b;
    outputs(4853) <= a and not b;
    outputs(4854) <= not b;
    outputs(4855) <= not a;
    outputs(4856) <= not b;
    outputs(4857) <= not (a xor b);
    outputs(4858) <= b and not a;
    outputs(4859) <= a or b;
    outputs(4860) <= a;
    outputs(4861) <= not (a and b);
    outputs(4862) <= not (a or b);
    outputs(4863) <= not b;
    outputs(4864) <= a;
    outputs(4865) <= b and not a;
    outputs(4866) <= not (a or b);
    outputs(4867) <= not b or a;
    outputs(4868) <= not b or a;
    outputs(4869) <= a and not b;
    outputs(4870) <= not a;
    outputs(4871) <= not b;
    outputs(4872) <= not b;
    outputs(4873) <= b;
    outputs(4874) <= b;
    outputs(4875) <= a and b;
    outputs(4876) <= not (a xor b);
    outputs(4877) <= b and not a;
    outputs(4878) <= not (a xor b);
    outputs(4879) <= b and not a;
    outputs(4880) <= a and b;
    outputs(4881) <= b;
    outputs(4882) <= not (a xor b);
    outputs(4883) <= not (a xor b);
    outputs(4884) <= not (a or b);
    outputs(4885) <= b and not a;
    outputs(4886) <= b and not a;
    outputs(4887) <= a;
    outputs(4888) <= not b;
    outputs(4889) <= not b;
    outputs(4890) <= b and not a;
    outputs(4891) <= not b or a;
    outputs(4892) <= a and not b;
    outputs(4893) <= b;
    outputs(4894) <= not b;
    outputs(4895) <= not a;
    outputs(4896) <= not b;
    outputs(4897) <= a and b;
    outputs(4898) <= a;
    outputs(4899) <= a xor b;
    outputs(4900) <= a;
    outputs(4901) <= b;
    outputs(4902) <= not a;
    outputs(4903) <= a and b;
    outputs(4904) <= b and not a;
    outputs(4905) <= not b;
    outputs(4906) <= a;
    outputs(4907) <= b and not a;
    outputs(4908) <= a xor b;
    outputs(4909) <= b;
    outputs(4910) <= a and b;
    outputs(4911) <= a or b;
    outputs(4912) <= a;
    outputs(4913) <= a;
    outputs(4914) <= a and b;
    outputs(4915) <= b and not a;
    outputs(4916) <= a xor b;
    outputs(4917) <= a;
    outputs(4918) <= not (a or b);
    outputs(4919) <= a;
    outputs(4920) <= a;
    outputs(4921) <= a and b;
    outputs(4922) <= not (a xor b);
    outputs(4923) <= not a;
    outputs(4924) <= a;
    outputs(4925) <= b;
    outputs(4926) <= not (a xor b);
    outputs(4927) <= not a;
    outputs(4928) <= not a;
    outputs(4929) <= b;
    outputs(4930) <= a;
    outputs(4931) <= a or b;
    outputs(4932) <= a;
    outputs(4933) <= b;
    outputs(4934) <= not b;
    outputs(4935) <= not a;
    outputs(4936) <= not b;
    outputs(4937) <= b and not a;
    outputs(4938) <= b and not a;
    outputs(4939) <= b;
    outputs(4940) <= b and not a;
    outputs(4941) <= a;
    outputs(4942) <= a and b;
    outputs(4943) <= not a;
    outputs(4944) <= b;
    outputs(4945) <= b and not a;
    outputs(4946) <= not b;
    outputs(4947) <= a xor b;
    outputs(4948) <= b;
    outputs(4949) <= not (a xor b);
    outputs(4950) <= not b;
    outputs(4951) <= a and not b;
    outputs(4952) <= a and not b;
    outputs(4953) <= not (a xor b);
    outputs(4954) <= a xor b;
    outputs(4955) <= a xor b;
    outputs(4956) <= not a;
    outputs(4957) <= a and not b;
    outputs(4958) <= not (a xor b);
    outputs(4959) <= not a;
    outputs(4960) <= b;
    outputs(4961) <= not b;
    outputs(4962) <= a;
    outputs(4963) <= a;
    outputs(4964) <= not a or b;
    outputs(4965) <= a;
    outputs(4966) <= not a;
    outputs(4967) <= a and b;
    outputs(4968) <= not (a xor b);
    outputs(4969) <= b;
    outputs(4970) <= not a;
    outputs(4971) <= not b;
    outputs(4972) <= a and b;
    outputs(4973) <= not (a or b);
    outputs(4974) <= a xor b;
    outputs(4975) <= not (a and b);
    outputs(4976) <= b;
    outputs(4977) <= not (a or b);
    outputs(4978) <= a and b;
    outputs(4979) <= a and b;
    outputs(4980) <= b;
    outputs(4981) <= not (a and b);
    outputs(4982) <= not a or b;
    outputs(4983) <= a and b;
    outputs(4984) <= not (a xor b);
    outputs(4985) <= a;
    outputs(4986) <= not b;
    outputs(4987) <= a and b;
    outputs(4988) <= b;
    outputs(4989) <= a or b;
    outputs(4990) <= not a;
    outputs(4991) <= b;
    outputs(4992) <= b;
    outputs(4993) <= a and b;
    outputs(4994) <= not a or b;
    outputs(4995) <= a xor b;
    outputs(4996) <= not b;
    outputs(4997) <= not (a or b);
    outputs(4998) <= a or b;
    outputs(4999) <= not b;
    outputs(5000) <= not b;
    outputs(5001) <= b;
    outputs(5002) <= not a;
    outputs(5003) <= not (a xor b);
    outputs(5004) <= a xor b;
    outputs(5005) <= a and b;
    outputs(5006) <= b and not a;
    outputs(5007) <= a and not b;
    outputs(5008) <= not a;
    outputs(5009) <= not a;
    outputs(5010) <= not (a xor b);
    outputs(5011) <= b and not a;
    outputs(5012) <= a and not b;
    outputs(5013) <= b and not a;
    outputs(5014) <= not (a xor b);
    outputs(5015) <= not a;
    outputs(5016) <= not a;
    outputs(5017) <= not b;
    outputs(5018) <= not a;
    outputs(5019) <= not (a or b);
    outputs(5020) <= not b;
    outputs(5021) <= a;
    outputs(5022) <= b and not a;
    outputs(5023) <= a;
    outputs(5024) <= a and not b;
    outputs(5025) <= a xor b;
    outputs(5026) <= a and b;
    outputs(5027) <= not (a or b);
    outputs(5028) <= not b;
    outputs(5029) <= a and not b;
    outputs(5030) <= a;
    outputs(5031) <= not (a xor b);
    outputs(5032) <= not (a xor b);
    outputs(5033) <= not a;
    outputs(5034) <= not (a xor b);
    outputs(5035) <= a and not b;
    outputs(5036) <= b and not a;
    outputs(5037) <= a;
    outputs(5038) <= b;
    outputs(5039) <= a or b;
    outputs(5040) <= not b;
    outputs(5041) <= a;
    outputs(5042) <= not (a xor b);
    outputs(5043) <= a and not b;
    outputs(5044) <= a and b;
    outputs(5045) <= a xor b;
    outputs(5046) <= a xor b;
    outputs(5047) <= not a;
    outputs(5048) <= a;
    outputs(5049) <= not (a xor b);
    outputs(5050) <= a xor b;
    outputs(5051) <= not (a or b);
    outputs(5052) <= a;
    outputs(5053) <= not b;
    outputs(5054) <= b;
    outputs(5055) <= a and b;
    outputs(5056) <= a and b;
    outputs(5057) <= not b;
    outputs(5058) <= not (a xor b);
    outputs(5059) <= b;
    outputs(5060) <= a and b;
    outputs(5061) <= not a;
    outputs(5062) <= not (a xor b);
    outputs(5063) <= a and not b;
    outputs(5064) <= b;
    outputs(5065) <= not b;
    outputs(5066) <= b and not a;
    outputs(5067) <= a and not b;
    outputs(5068) <= not b;
    outputs(5069) <= not (a xor b);
    outputs(5070) <= not a;
    outputs(5071) <= a and b;
    outputs(5072) <= not (a xor b);
    outputs(5073) <= a and not b;
    outputs(5074) <= not a or b;
    outputs(5075) <= not a or b;
    outputs(5076) <= not b or a;
    outputs(5077) <= b and not a;
    outputs(5078) <= not a;
    outputs(5079) <= a;
    outputs(5080) <= a and b;
    outputs(5081) <= a xor b;
    outputs(5082) <= b and not a;
    outputs(5083) <= a and not b;
    outputs(5084) <= a or b;
    outputs(5085) <= not (a xor b);
    outputs(5086) <= a and b;
    outputs(5087) <= a;
    outputs(5088) <= not (a or b);
    outputs(5089) <= a;
    outputs(5090) <= not b;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= not b;
    outputs(5093) <= not a or b;
    outputs(5094) <= a or b;
    outputs(5095) <= not b;
    outputs(5096) <= a xor b;
    outputs(5097) <= a or b;
    outputs(5098) <= not b;
    outputs(5099) <= b;
    outputs(5100) <= b;
    outputs(5101) <= not a or b;
    outputs(5102) <= b;
    outputs(5103) <= not (a and b);
    outputs(5104) <= b;
    outputs(5105) <= b;
    outputs(5106) <= not a;
    outputs(5107) <= b;
    outputs(5108) <= not b;
    outputs(5109) <= a;
    outputs(5110) <= a xor b;
    outputs(5111) <= not (a xor b);
    outputs(5112) <= not b;
    outputs(5113) <= a or b;
    outputs(5114) <= not (a or b);
    outputs(5115) <= b;
    outputs(5116) <= a;
    outputs(5117) <= a or b;
    outputs(5118) <= not a;
    outputs(5119) <= a and b;
end Behavioral;
