library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(7679 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(7679 downto 0);

begin

    layer0_outputs(0) <= (inputs(22)) and not (inputs(142));
    layer0_outputs(1) <= (inputs(66)) and (inputs(235));
    layer0_outputs(2) <= (inputs(151)) or (inputs(224));
    layer0_outputs(3) <= (inputs(41)) or (inputs(8));
    layer0_outputs(4) <= (inputs(52)) and (inputs(29));
    layer0_outputs(5) <= not(inputs(121));
    layer0_outputs(6) <= not(inputs(29));
    layer0_outputs(7) <= not((inputs(138)) or (inputs(217)));
    layer0_outputs(8) <= not((inputs(11)) and (inputs(186)));
    layer0_outputs(9) <= inputs(136);
    layer0_outputs(10) <= inputs(33);
    layer0_outputs(11) <= not(inputs(33)) or (inputs(105));
    layer0_outputs(12) <= not((inputs(20)) or (inputs(195)));
    layer0_outputs(13) <= not(inputs(252));
    layer0_outputs(14) <= (inputs(178)) xor (inputs(189));
    layer0_outputs(15) <= not(inputs(138)) or (inputs(26));
    layer0_outputs(16) <= not(inputs(155)) or (inputs(18));
    layer0_outputs(17) <= not(inputs(133)) or (inputs(132));
    layer0_outputs(18) <= not(inputs(26));
    layer0_outputs(19) <= not(inputs(40));
    layer0_outputs(20) <= not(inputs(69));
    layer0_outputs(21) <= not(inputs(254));
    layer0_outputs(22) <= not((inputs(153)) and (inputs(151)));
    layer0_outputs(23) <= not(inputs(231));
    layer0_outputs(24) <= not((inputs(233)) or (inputs(64)));
    layer0_outputs(25) <= (inputs(125)) and not (inputs(80));
    layer0_outputs(26) <= not((inputs(202)) xor (inputs(130)));
    layer0_outputs(27) <= not((inputs(176)) or (inputs(30)));
    layer0_outputs(28) <= not(inputs(23)) or (inputs(208));
    layer0_outputs(29) <= not((inputs(164)) xor (inputs(61)));
    layer0_outputs(30) <= (inputs(252)) or (inputs(123));
    layer0_outputs(31) <= not((inputs(133)) or (inputs(175)));
    layer0_outputs(32) <= (inputs(224)) xor (inputs(237));
    layer0_outputs(33) <= not((inputs(40)) and (inputs(165)));
    layer0_outputs(34) <= not(inputs(202)) or (inputs(109));
    layer0_outputs(35) <= not(inputs(173)) or (inputs(139));
    layer0_outputs(36) <= not(inputs(93)) or (inputs(183));
    layer0_outputs(37) <= not(inputs(187));
    layer0_outputs(38) <= inputs(210);
    layer0_outputs(39) <= inputs(246);
    layer0_outputs(40) <= not(inputs(89)) or (inputs(22));
    layer0_outputs(41) <= inputs(2);
    layer0_outputs(42) <= not((inputs(80)) or (inputs(29)));
    layer0_outputs(43) <= (inputs(28)) xor (inputs(164));
    layer0_outputs(44) <= not((inputs(132)) xor (inputs(196)));
    layer0_outputs(45) <= not(inputs(80)) or (inputs(95));
    layer0_outputs(46) <= not(inputs(6));
    layer0_outputs(47) <= not(inputs(249));
    layer0_outputs(48) <= not((inputs(109)) xor (inputs(111)));
    layer0_outputs(49) <= not((inputs(21)) or (inputs(145)));
    layer0_outputs(50) <= not(inputs(130));
    layer0_outputs(51) <= (inputs(166)) and not (inputs(139));
    layer0_outputs(52) <= not((inputs(126)) xor (inputs(18)));
    layer0_outputs(53) <= (inputs(228)) and not (inputs(208));
    layer0_outputs(54) <= (inputs(220)) xor (inputs(139));
    layer0_outputs(55) <= (inputs(209)) or (inputs(28));
    layer0_outputs(56) <= (inputs(209)) xor (inputs(158));
    layer0_outputs(57) <= not(inputs(30));
    layer0_outputs(58) <= not(inputs(24));
    layer0_outputs(59) <= not((inputs(253)) xor (inputs(171)));
    layer0_outputs(60) <= (inputs(247)) and not (inputs(6));
    layer0_outputs(61) <= (inputs(104)) or (inputs(177));
    layer0_outputs(62) <= (inputs(109)) or (inputs(150));
    layer0_outputs(63) <= not(inputs(194)) or (inputs(130));
    layer0_outputs(64) <= not((inputs(56)) or (inputs(112)));
    layer0_outputs(65) <= not(inputs(241)) or (inputs(175));
    layer0_outputs(66) <= not(inputs(212)) or (inputs(31));
    layer0_outputs(67) <= not(inputs(187));
    layer0_outputs(68) <= not(inputs(223));
    layer0_outputs(69) <= '1';
    layer0_outputs(70) <= (inputs(23)) and not (inputs(178));
    layer0_outputs(71) <= (inputs(113)) or (inputs(58));
    layer0_outputs(72) <= not(inputs(228));
    layer0_outputs(73) <= inputs(35);
    layer0_outputs(74) <= (inputs(124)) and not (inputs(162));
    layer0_outputs(75) <= not((inputs(133)) xor (inputs(102)));
    layer0_outputs(76) <= not(inputs(231)) or (inputs(240));
    layer0_outputs(77) <= (inputs(7)) or (inputs(111));
    layer0_outputs(78) <= (inputs(126)) xor (inputs(57));
    layer0_outputs(79) <= not(inputs(214)) or (inputs(49));
    layer0_outputs(80) <= not((inputs(217)) xor (inputs(248)));
    layer0_outputs(81) <= (inputs(240)) or (inputs(242));
    layer0_outputs(82) <= not(inputs(41)) or (inputs(114));
    layer0_outputs(83) <= (inputs(91)) or (inputs(245));
    layer0_outputs(84) <= (inputs(26)) or (inputs(64));
    layer0_outputs(85) <= not(inputs(137));
    layer0_outputs(86) <= inputs(72);
    layer0_outputs(87) <= not(inputs(26)) or (inputs(143));
    layer0_outputs(88) <= (inputs(172)) and not (inputs(178));
    layer0_outputs(89) <= (inputs(22)) or (inputs(96));
    layer0_outputs(90) <= not((inputs(53)) or (inputs(13)));
    layer0_outputs(91) <= (inputs(250)) xor (inputs(108));
    layer0_outputs(92) <= not(inputs(30)) or (inputs(87));
    layer0_outputs(93) <= not((inputs(187)) xor (inputs(98)));
    layer0_outputs(94) <= (inputs(188)) or (inputs(161));
    layer0_outputs(95) <= not(inputs(115)) or (inputs(192));
    layer0_outputs(96) <= not(inputs(94));
    layer0_outputs(97) <= inputs(193);
    layer0_outputs(98) <= (inputs(22)) or (inputs(192));
    layer0_outputs(99) <= not((inputs(255)) and (inputs(150)));
    layer0_outputs(100) <= not(inputs(203));
    layer0_outputs(101) <= (inputs(108)) or (inputs(64));
    layer0_outputs(102) <= (inputs(189)) xor (inputs(156));
    layer0_outputs(103) <= (inputs(109)) and not (inputs(208));
    layer0_outputs(104) <= not(inputs(25));
    layer0_outputs(105) <= (inputs(224)) and (inputs(239));
    layer0_outputs(106) <= not((inputs(250)) or (inputs(104)));
    layer0_outputs(107) <= (inputs(95)) or (inputs(170));
    layer0_outputs(108) <= not((inputs(189)) or (inputs(78)));
    layer0_outputs(109) <= (inputs(18)) and (inputs(175));
    layer0_outputs(110) <= (inputs(222)) or (inputs(239));
    layer0_outputs(111) <= (inputs(195)) and not (inputs(79));
    layer0_outputs(112) <= not(inputs(232));
    layer0_outputs(113) <= (inputs(196)) or (inputs(56));
    layer0_outputs(114) <= inputs(165);
    layer0_outputs(115) <= not(inputs(4)) or (inputs(130));
    layer0_outputs(116) <= (inputs(154)) xor (inputs(218));
    layer0_outputs(117) <= (inputs(125)) and not (inputs(237));
    layer0_outputs(118) <= (inputs(27)) or (inputs(197));
    layer0_outputs(119) <= (inputs(84)) or (inputs(94));
    layer0_outputs(120) <= not((inputs(85)) or (inputs(249)));
    layer0_outputs(121) <= (inputs(13)) or (inputs(127));
    layer0_outputs(122) <= not(inputs(175));
    layer0_outputs(123) <= (inputs(245)) xor (inputs(112));
    layer0_outputs(124) <= not(inputs(44));
    layer0_outputs(125) <= not((inputs(173)) or (inputs(83)));
    layer0_outputs(126) <= (inputs(73)) and not (inputs(155));
    layer0_outputs(127) <= (inputs(191)) and not (inputs(216));
    layer0_outputs(128) <= inputs(85);
    layer0_outputs(129) <= not(inputs(81));
    layer0_outputs(130) <= not(inputs(19));
    layer0_outputs(131) <= (inputs(102)) and not (inputs(65));
    layer0_outputs(132) <= inputs(136);
    layer0_outputs(133) <= not(inputs(44));
    layer0_outputs(134) <= not(inputs(83));
    layer0_outputs(135) <= (inputs(233)) or (inputs(41));
    layer0_outputs(136) <= (inputs(54)) or (inputs(81));
    layer0_outputs(137) <= not(inputs(24));
    layer0_outputs(138) <= not((inputs(87)) xor (inputs(50)));
    layer0_outputs(139) <= not((inputs(63)) or (inputs(160)));
    layer0_outputs(140) <= (inputs(187)) or (inputs(99));
    layer0_outputs(141) <= (inputs(168)) and not (inputs(49));
    layer0_outputs(142) <= (inputs(51)) xor (inputs(11));
    layer0_outputs(143) <= (inputs(14)) or (inputs(247));
    layer0_outputs(144) <= (inputs(142)) or (inputs(135));
    layer0_outputs(145) <= '1';
    layer0_outputs(146) <= inputs(212);
    layer0_outputs(147) <= not(inputs(85));
    layer0_outputs(148) <= (inputs(179)) xor (inputs(174));
    layer0_outputs(149) <= not(inputs(97));
    layer0_outputs(150) <= (inputs(1)) and (inputs(19));
    layer0_outputs(151) <= inputs(117);
    layer0_outputs(152) <= inputs(75);
    layer0_outputs(153) <= not(inputs(166)) or (inputs(12));
    layer0_outputs(154) <= (inputs(156)) or (inputs(206));
    layer0_outputs(155) <= not(inputs(146)) or (inputs(87));
    layer0_outputs(156) <= not((inputs(21)) or (inputs(193)));
    layer0_outputs(157) <= not(inputs(5)) or (inputs(173));
    layer0_outputs(158) <= '1';
    layer0_outputs(159) <= not((inputs(206)) xor (inputs(95)));
    layer0_outputs(160) <= not((inputs(55)) and (inputs(242)));
    layer0_outputs(161) <= (inputs(243)) or (inputs(104));
    layer0_outputs(162) <= not((inputs(125)) or (inputs(187)));
    layer0_outputs(163) <= (inputs(35)) or (inputs(210));
    layer0_outputs(164) <= not((inputs(241)) or (inputs(151)));
    layer0_outputs(165) <= (inputs(161)) xor (inputs(103));
    layer0_outputs(166) <= not(inputs(98));
    layer0_outputs(167) <= (inputs(176)) xor (inputs(147));
    layer0_outputs(168) <= (inputs(221)) xor (inputs(56));
    layer0_outputs(169) <= (inputs(198)) or (inputs(192));
    layer0_outputs(170) <= (inputs(61)) and not (inputs(219));
    layer0_outputs(171) <= (inputs(105)) and not (inputs(172));
    layer0_outputs(172) <= (inputs(20)) and (inputs(188));
    layer0_outputs(173) <= (inputs(166)) or (inputs(110));
    layer0_outputs(174) <= (inputs(211)) xor (inputs(200));
    layer0_outputs(175) <= (inputs(8)) and not (inputs(97));
    layer0_outputs(176) <= not(inputs(83)) or (inputs(240));
    layer0_outputs(177) <= inputs(131);
    layer0_outputs(178) <= not(inputs(218));
    layer0_outputs(179) <= (inputs(229)) xor (inputs(161));
    layer0_outputs(180) <= (inputs(92)) xor (inputs(150));
    layer0_outputs(181) <= not(inputs(188)) or (inputs(14));
    layer0_outputs(182) <= not((inputs(183)) and (inputs(190)));
    layer0_outputs(183) <= not((inputs(108)) and (inputs(139)));
    layer0_outputs(184) <= not(inputs(234));
    layer0_outputs(185) <= (inputs(162)) xor (inputs(168));
    layer0_outputs(186) <= (inputs(68)) or (inputs(24));
    layer0_outputs(187) <= (inputs(5)) xor (inputs(238));
    layer0_outputs(188) <= not(inputs(156));
    layer0_outputs(189) <= (inputs(188)) or (inputs(210));
    layer0_outputs(190) <= (inputs(111)) and not (inputs(235));
    layer0_outputs(191) <= (inputs(103)) or (inputs(137));
    layer0_outputs(192) <= not((inputs(41)) xor (inputs(117)));
    layer0_outputs(193) <= not((inputs(26)) or (inputs(63)));
    layer0_outputs(194) <= (inputs(172)) or (inputs(71));
    layer0_outputs(195) <= not(inputs(125));
    layer0_outputs(196) <= (inputs(178)) xor (inputs(142));
    layer0_outputs(197) <= (inputs(156)) xor (inputs(39));
    layer0_outputs(198) <= not((inputs(65)) or (inputs(240)));
    layer0_outputs(199) <= not(inputs(228));
    layer0_outputs(200) <= not((inputs(217)) xor (inputs(4)));
    layer0_outputs(201) <= not(inputs(91));
    layer0_outputs(202) <= inputs(231);
    layer0_outputs(203) <= not((inputs(237)) or (inputs(7)));
    layer0_outputs(204) <= (inputs(88)) and (inputs(68));
    layer0_outputs(205) <= not((inputs(187)) and (inputs(155)));
    layer0_outputs(206) <= not((inputs(143)) or (inputs(58)));
    layer0_outputs(207) <= inputs(169);
    layer0_outputs(208) <= not(inputs(104));
    layer0_outputs(209) <= (inputs(252)) or (inputs(121));
    layer0_outputs(210) <= (inputs(108)) and not (inputs(3));
    layer0_outputs(211) <= not(inputs(163));
    layer0_outputs(212) <= (inputs(15)) or (inputs(141));
    layer0_outputs(213) <= (inputs(113)) and (inputs(97));
    layer0_outputs(214) <= (inputs(33)) or (inputs(153));
    layer0_outputs(215) <= inputs(36);
    layer0_outputs(216) <= inputs(10);
    layer0_outputs(217) <= (inputs(37)) or (inputs(93));
    layer0_outputs(218) <= inputs(158);
    layer0_outputs(219) <= not((inputs(20)) xor (inputs(123)));
    layer0_outputs(220) <= not((inputs(217)) and (inputs(230)));
    layer0_outputs(221) <= not(inputs(139)) or (inputs(160));
    layer0_outputs(222) <= inputs(59);
    layer0_outputs(223) <= not(inputs(229));
    layer0_outputs(224) <= inputs(170);
    layer0_outputs(225) <= not((inputs(104)) or (inputs(92)));
    layer0_outputs(226) <= inputs(37);
    layer0_outputs(227) <= not((inputs(189)) or (inputs(0)));
    layer0_outputs(228) <= not((inputs(39)) and (inputs(53)));
    layer0_outputs(229) <= not((inputs(73)) xor (inputs(250)));
    layer0_outputs(230) <= (inputs(196)) and not (inputs(108));
    layer0_outputs(231) <= (inputs(85)) or (inputs(178));
    layer0_outputs(232) <= (inputs(18)) or (inputs(110));
    layer0_outputs(233) <= not(inputs(231)) or (inputs(147));
    layer0_outputs(234) <= inputs(98);
    layer0_outputs(235) <= not((inputs(132)) or (inputs(52)));
    layer0_outputs(236) <= (inputs(14)) or (inputs(215));
    layer0_outputs(237) <= '1';
    layer0_outputs(238) <= not(inputs(172));
    layer0_outputs(239) <= not(inputs(26));
    layer0_outputs(240) <= (inputs(148)) and not (inputs(1));
    layer0_outputs(241) <= inputs(169);
    layer0_outputs(242) <= inputs(135);
    layer0_outputs(243) <= not(inputs(126)) or (inputs(177));
    layer0_outputs(244) <= inputs(86);
    layer0_outputs(245) <= inputs(98);
    layer0_outputs(246) <= (inputs(234)) and not (inputs(99));
    layer0_outputs(247) <= (inputs(73)) or (inputs(83));
    layer0_outputs(248) <= not(inputs(212));
    layer0_outputs(249) <= (inputs(246)) and not (inputs(244));
    layer0_outputs(250) <= (inputs(205)) and not (inputs(132));
    layer0_outputs(251) <= (inputs(69)) xor (inputs(176));
    layer0_outputs(252) <= not(inputs(46)) or (inputs(208));
    layer0_outputs(253) <= inputs(108);
    layer0_outputs(254) <= (inputs(9)) or (inputs(50));
    layer0_outputs(255) <= inputs(246);
    layer0_outputs(256) <= inputs(180);
    layer0_outputs(257) <= inputs(94);
    layer0_outputs(258) <= (inputs(213)) or (inputs(79));
    layer0_outputs(259) <= inputs(222);
    layer0_outputs(260) <= (inputs(48)) xor (inputs(98));
    layer0_outputs(261) <= (inputs(114)) xor (inputs(144));
    layer0_outputs(262) <= (inputs(2)) xor (inputs(29));
    layer0_outputs(263) <= not(inputs(80));
    layer0_outputs(264) <= (inputs(216)) xor (inputs(184));
    layer0_outputs(265) <= (inputs(188)) and not (inputs(127));
    layer0_outputs(266) <= not((inputs(195)) or (inputs(53)));
    layer0_outputs(267) <= (inputs(141)) or (inputs(181));
    layer0_outputs(268) <= inputs(6);
    layer0_outputs(269) <= (inputs(247)) xor (inputs(213));
    layer0_outputs(270) <= not(inputs(122));
    layer0_outputs(271) <= inputs(232);
    layer0_outputs(272) <= not(inputs(23)) or (inputs(30));
    layer0_outputs(273) <= (inputs(72)) and not (inputs(27));
    layer0_outputs(274) <= not((inputs(35)) xor (inputs(224)));
    layer0_outputs(275) <= (inputs(129)) and not (inputs(145));
    layer0_outputs(276) <= not(inputs(182));
    layer0_outputs(277) <= (inputs(120)) and not (inputs(99));
    layer0_outputs(278) <= not((inputs(0)) xor (inputs(253)));
    layer0_outputs(279) <= inputs(243);
    layer0_outputs(280) <= not((inputs(163)) xor (inputs(145)));
    layer0_outputs(281) <= not((inputs(175)) xor (inputs(202)));
    layer0_outputs(282) <= not(inputs(60));
    layer0_outputs(283) <= not(inputs(128));
    layer0_outputs(284) <= (inputs(142)) or (inputs(235));
    layer0_outputs(285) <= (inputs(160)) or (inputs(170));
    layer0_outputs(286) <= inputs(23);
    layer0_outputs(287) <= inputs(231);
    layer0_outputs(288) <= (inputs(156)) and not (inputs(50));
    layer0_outputs(289) <= (inputs(118)) and not (inputs(241));
    layer0_outputs(290) <= inputs(231);
    layer0_outputs(291) <= not(inputs(212));
    layer0_outputs(292) <= not(inputs(113));
    layer0_outputs(293) <= not((inputs(61)) or (inputs(9)));
    layer0_outputs(294) <= not(inputs(5));
    layer0_outputs(295) <= not((inputs(73)) xor (inputs(150)));
    layer0_outputs(296) <= not((inputs(180)) xor (inputs(110)));
    layer0_outputs(297) <= inputs(196);
    layer0_outputs(298) <= not((inputs(154)) or (inputs(37)));
    layer0_outputs(299) <= not(inputs(155)) or (inputs(199));
    layer0_outputs(300) <= not(inputs(12));
    layer0_outputs(301) <= (inputs(27)) and not (inputs(153));
    layer0_outputs(302) <= not((inputs(160)) or (inputs(182)));
    layer0_outputs(303) <= (inputs(108)) or (inputs(191));
    layer0_outputs(304) <= not(inputs(120));
    layer0_outputs(305) <= not(inputs(147));
    layer0_outputs(306) <= (inputs(173)) and not (inputs(122));
    layer0_outputs(307) <= not(inputs(195)) or (inputs(110));
    layer0_outputs(308) <= inputs(85);
    layer0_outputs(309) <= not(inputs(22));
    layer0_outputs(310) <= not((inputs(214)) or (inputs(112)));
    layer0_outputs(311) <= not((inputs(169)) or (inputs(100)));
    layer0_outputs(312) <= '1';
    layer0_outputs(313) <= (inputs(71)) xor (inputs(200));
    layer0_outputs(314) <= inputs(158);
    layer0_outputs(315) <= not(inputs(137)) or (inputs(55));
    layer0_outputs(316) <= (inputs(18)) and not (inputs(81));
    layer0_outputs(317) <= inputs(216);
    layer0_outputs(318) <= not(inputs(44));
    layer0_outputs(319) <= not((inputs(104)) xor (inputs(169)));
    layer0_outputs(320) <= inputs(144);
    layer0_outputs(321) <= (inputs(210)) or (inputs(80));
    layer0_outputs(322) <= not(inputs(179));
    layer0_outputs(323) <= not(inputs(82));
    layer0_outputs(324) <= not(inputs(160));
    layer0_outputs(325) <= (inputs(0)) or (inputs(155));
    layer0_outputs(326) <= (inputs(161)) or (inputs(230));
    layer0_outputs(327) <= (inputs(245)) or (inputs(177));
    layer0_outputs(328) <= (inputs(126)) or (inputs(166));
    layer0_outputs(329) <= not((inputs(36)) and (inputs(28)));
    layer0_outputs(330) <= not((inputs(227)) and (inputs(184)));
    layer0_outputs(331) <= (inputs(60)) and not (inputs(145));
    layer0_outputs(332) <= not((inputs(223)) xor (inputs(54)));
    layer0_outputs(333) <= (inputs(241)) xor (inputs(37));
    layer0_outputs(334) <= not(inputs(52));
    layer0_outputs(335) <= not(inputs(185)) or (inputs(87));
    layer0_outputs(336) <= (inputs(127)) or (inputs(5));
    layer0_outputs(337) <= inputs(194);
    layer0_outputs(338) <= not((inputs(102)) xor (inputs(189)));
    layer0_outputs(339) <= not((inputs(71)) or (inputs(234)));
    layer0_outputs(340) <= (inputs(106)) or (inputs(131));
    layer0_outputs(341) <= not(inputs(58)) or (inputs(63));
    layer0_outputs(342) <= not((inputs(61)) xor (inputs(240)));
    layer0_outputs(343) <= (inputs(230)) and (inputs(6));
    layer0_outputs(344) <= not(inputs(61)) or (inputs(225));
    layer0_outputs(345) <= inputs(150);
    layer0_outputs(346) <= inputs(192);
    layer0_outputs(347) <= not((inputs(226)) xor (inputs(12)));
    layer0_outputs(348) <= inputs(178);
    layer0_outputs(349) <= not((inputs(178)) or (inputs(127)));
    layer0_outputs(350) <= not((inputs(38)) or (inputs(155)));
    layer0_outputs(351) <= (inputs(6)) or (inputs(19));
    layer0_outputs(352) <= not((inputs(137)) or (inputs(117)));
    layer0_outputs(353) <= inputs(36);
    layer0_outputs(354) <= not((inputs(100)) xor (inputs(113)));
    layer0_outputs(355) <= not(inputs(176));
    layer0_outputs(356) <= (inputs(61)) or (inputs(125));
    layer0_outputs(357) <= inputs(141);
    layer0_outputs(358) <= inputs(182);
    layer0_outputs(359) <= (inputs(28)) or (inputs(113));
    layer0_outputs(360) <= (inputs(211)) or (inputs(114));
    layer0_outputs(361) <= '0';
    layer0_outputs(362) <= (inputs(192)) or (inputs(17));
    layer0_outputs(363) <= inputs(82);
    layer0_outputs(364) <= inputs(130);
    layer0_outputs(365) <= not(inputs(216)) or (inputs(107));
    layer0_outputs(366) <= (inputs(179)) or (inputs(252));
    layer0_outputs(367) <= (inputs(2)) and (inputs(58));
    layer0_outputs(368) <= (inputs(12)) and not (inputs(76));
    layer0_outputs(369) <= not((inputs(126)) or (inputs(27)));
    layer0_outputs(370) <= (inputs(141)) and not (inputs(253));
    layer0_outputs(371) <= not(inputs(33));
    layer0_outputs(372) <= not((inputs(32)) xor (inputs(66)));
    layer0_outputs(373) <= not((inputs(88)) xor (inputs(141)));
    layer0_outputs(374) <= (inputs(113)) and not (inputs(79));
    layer0_outputs(375) <= not((inputs(10)) or (inputs(155)));
    layer0_outputs(376) <= not(inputs(1)) or (inputs(18));
    layer0_outputs(377) <= (inputs(127)) or (inputs(98));
    layer0_outputs(378) <= not((inputs(230)) and (inputs(26)));
    layer0_outputs(379) <= inputs(140);
    layer0_outputs(380) <= inputs(237);
    layer0_outputs(381) <= (inputs(172)) and not (inputs(46));
    layer0_outputs(382) <= not(inputs(220));
    layer0_outputs(383) <= inputs(198);
    layer0_outputs(384) <= inputs(62);
    layer0_outputs(385) <= not(inputs(218)) or (inputs(54));
    layer0_outputs(386) <= inputs(141);
    layer0_outputs(387) <= not((inputs(60)) xor (inputs(255)));
    layer0_outputs(388) <= '1';
    layer0_outputs(389) <= inputs(101);
    layer0_outputs(390) <= not(inputs(93)) or (inputs(238));
    layer0_outputs(391) <= inputs(213);
    layer0_outputs(392) <= (inputs(158)) or (inputs(103));
    layer0_outputs(393) <= (inputs(117)) and not (inputs(188));
    layer0_outputs(394) <= '1';
    layer0_outputs(395) <= (inputs(235)) and not (inputs(128));
    layer0_outputs(396) <= (inputs(122)) xor (inputs(91));
    layer0_outputs(397) <= (inputs(23)) and not (inputs(236));
    layer0_outputs(398) <= (inputs(74)) xor (inputs(72));
    layer0_outputs(399) <= (inputs(82)) or (inputs(116));
    layer0_outputs(400) <= (inputs(54)) or (inputs(108));
    layer0_outputs(401) <= not(inputs(22));
    layer0_outputs(402) <= (inputs(183)) and not (inputs(99));
    layer0_outputs(403) <= not((inputs(23)) xor (inputs(142)));
    layer0_outputs(404) <= inputs(53);
    layer0_outputs(405) <= inputs(231);
    layer0_outputs(406) <= (inputs(216)) xor (inputs(139));
    layer0_outputs(407) <= not(inputs(78));
    layer0_outputs(408) <= not(inputs(150)) or (inputs(80));
    layer0_outputs(409) <= (inputs(186)) and not (inputs(194));
    layer0_outputs(410) <= not(inputs(3));
    layer0_outputs(411) <= inputs(203);
    layer0_outputs(412) <= not((inputs(163)) or (inputs(165)));
    layer0_outputs(413) <= (inputs(148)) or (inputs(13));
    layer0_outputs(414) <= (inputs(210)) or (inputs(230));
    layer0_outputs(415) <= '1';
    layer0_outputs(416) <= (inputs(148)) and not (inputs(94));
    layer0_outputs(417) <= (inputs(7)) and not (inputs(3));
    layer0_outputs(418) <= not((inputs(95)) or (inputs(253)));
    layer0_outputs(419) <= (inputs(204)) or (inputs(152));
    layer0_outputs(420) <= (inputs(42)) and not (inputs(203));
    layer0_outputs(421) <= not(inputs(78));
    layer0_outputs(422) <= not(inputs(226)) or (inputs(243));
    layer0_outputs(423) <= not(inputs(235));
    layer0_outputs(424) <= (inputs(102)) and not (inputs(189));
    layer0_outputs(425) <= '0';
    layer0_outputs(426) <= (inputs(186)) and not (inputs(1));
    layer0_outputs(427) <= not((inputs(21)) or (inputs(120)));
    layer0_outputs(428) <= not(inputs(109));
    layer0_outputs(429) <= not((inputs(8)) xor (inputs(59)));
    layer0_outputs(430) <= not(inputs(21));
    layer0_outputs(431) <= (inputs(105)) xor (inputs(223));
    layer0_outputs(432) <= not(inputs(234));
    layer0_outputs(433) <= not((inputs(78)) or (inputs(226)));
    layer0_outputs(434) <= (inputs(121)) and not (inputs(39));
    layer0_outputs(435) <= not(inputs(150));
    layer0_outputs(436) <= not(inputs(134));
    layer0_outputs(437) <= not(inputs(19));
    layer0_outputs(438) <= inputs(78);
    layer0_outputs(439) <= inputs(198);
    layer0_outputs(440) <= (inputs(194)) and (inputs(58));
    layer0_outputs(441) <= inputs(102);
    layer0_outputs(442) <= inputs(119);
    layer0_outputs(443) <= not(inputs(177));
    layer0_outputs(444) <= not(inputs(246));
    layer0_outputs(445) <= not((inputs(12)) and (inputs(26)));
    layer0_outputs(446) <= inputs(100);
    layer0_outputs(447) <= not(inputs(255));
    layer0_outputs(448) <= (inputs(27)) and not (inputs(220));
    layer0_outputs(449) <= not(inputs(249)) or (inputs(123));
    layer0_outputs(450) <= inputs(211);
    layer0_outputs(451) <= not(inputs(233)) or (inputs(22));
    layer0_outputs(452) <= not(inputs(59)) or (inputs(191));
    layer0_outputs(453) <= not((inputs(89)) and (inputs(73)));
    layer0_outputs(454) <= not(inputs(79));
    layer0_outputs(455) <= (inputs(196)) or (inputs(208));
    layer0_outputs(456) <= (inputs(97)) and not (inputs(218));
    layer0_outputs(457) <= (inputs(26)) xor (inputs(63));
    layer0_outputs(458) <= (inputs(40)) and not (inputs(135));
    layer0_outputs(459) <= not((inputs(85)) xor (inputs(21)));
    layer0_outputs(460) <= inputs(137);
    layer0_outputs(461) <= (inputs(171)) xor (inputs(96));
    layer0_outputs(462) <= inputs(205);
    layer0_outputs(463) <= (inputs(9)) and (inputs(174));
    layer0_outputs(464) <= not(inputs(120)) or (inputs(179));
    layer0_outputs(465) <= not(inputs(198)) or (inputs(226));
    layer0_outputs(466) <= (inputs(182)) and (inputs(192));
    layer0_outputs(467) <= (inputs(162)) or (inputs(129));
    layer0_outputs(468) <= not(inputs(186)) or (inputs(53));
    layer0_outputs(469) <= (inputs(211)) and not (inputs(48));
    layer0_outputs(470) <= not((inputs(124)) xor (inputs(128)));
    layer0_outputs(471) <= inputs(148);
    layer0_outputs(472) <= not((inputs(97)) xor (inputs(208)));
    layer0_outputs(473) <= not(inputs(93)) or (inputs(223));
    layer0_outputs(474) <= not((inputs(168)) or (inputs(139)));
    layer0_outputs(475) <= not(inputs(72)) or (inputs(124));
    layer0_outputs(476) <= (inputs(58)) xor (inputs(224));
    layer0_outputs(477) <= not(inputs(197));
    layer0_outputs(478) <= (inputs(58)) or (inputs(77));
    layer0_outputs(479) <= (inputs(135)) and not (inputs(49));
    layer0_outputs(480) <= not(inputs(30));
    layer0_outputs(481) <= (inputs(234)) or (inputs(192));
    layer0_outputs(482) <= inputs(197);
    layer0_outputs(483) <= (inputs(66)) xor (inputs(186));
    layer0_outputs(484) <= (inputs(56)) or (inputs(33));
    layer0_outputs(485) <= inputs(98);
    layer0_outputs(486) <= not(inputs(116));
    layer0_outputs(487) <= inputs(32);
    layer0_outputs(488) <= not(inputs(134)) or (inputs(188));
    layer0_outputs(489) <= not(inputs(242)) or (inputs(17));
    layer0_outputs(490) <= inputs(110);
    layer0_outputs(491) <= not((inputs(124)) or (inputs(82)));
    layer0_outputs(492) <= not(inputs(179));
    layer0_outputs(493) <= (inputs(10)) and (inputs(44));
    layer0_outputs(494) <= not((inputs(219)) or (inputs(158)));
    layer0_outputs(495) <= not(inputs(82));
    layer0_outputs(496) <= (inputs(42)) xor (inputs(32));
    layer0_outputs(497) <= (inputs(172)) or (inputs(88));
    layer0_outputs(498) <= not(inputs(51));
    layer0_outputs(499) <= (inputs(170)) and not (inputs(49));
    layer0_outputs(500) <= not(inputs(4));
    layer0_outputs(501) <= inputs(70);
    layer0_outputs(502) <= not((inputs(126)) or (inputs(59)));
    layer0_outputs(503) <= inputs(118);
    layer0_outputs(504) <= (inputs(62)) and not (inputs(254));
    layer0_outputs(505) <= not(inputs(130));
    layer0_outputs(506) <= not((inputs(181)) or (inputs(190)));
    layer0_outputs(507) <= inputs(229);
    layer0_outputs(508) <= not(inputs(110)) or (inputs(239));
    layer0_outputs(509) <= not(inputs(245)) or (inputs(254));
    layer0_outputs(510) <= not((inputs(153)) xor (inputs(63)));
    layer0_outputs(511) <= not(inputs(86)) or (inputs(174));
    layer0_outputs(512) <= not(inputs(204)) or (inputs(41));
    layer0_outputs(513) <= inputs(100);
    layer0_outputs(514) <= (inputs(227)) xor (inputs(15));
    layer0_outputs(515) <= not(inputs(195)) or (inputs(46));
    layer0_outputs(516) <= '1';
    layer0_outputs(517) <= not(inputs(108));
    layer0_outputs(518) <= not((inputs(180)) and (inputs(140)));
    layer0_outputs(519) <= (inputs(137)) or (inputs(126));
    layer0_outputs(520) <= not(inputs(137)) or (inputs(38));
    layer0_outputs(521) <= not(inputs(126));
    layer0_outputs(522) <= not(inputs(152)) or (inputs(154));
    layer0_outputs(523) <= not(inputs(132)) or (inputs(207));
    layer0_outputs(524) <= (inputs(240)) or (inputs(44));
    layer0_outputs(525) <= inputs(82);
    layer0_outputs(526) <= not(inputs(28));
    layer0_outputs(527) <= (inputs(53)) and not (inputs(170));
    layer0_outputs(528) <= inputs(183);
    layer0_outputs(529) <= inputs(25);
    layer0_outputs(530) <= inputs(104);
    layer0_outputs(531) <= (inputs(250)) xor (inputs(159));
    layer0_outputs(532) <= (inputs(67)) and not (inputs(221));
    layer0_outputs(533) <= (inputs(203)) and not (inputs(1));
    layer0_outputs(534) <= not(inputs(244));
    layer0_outputs(535) <= not((inputs(101)) or (inputs(50)));
    layer0_outputs(536) <= not((inputs(148)) xor (inputs(190)));
    layer0_outputs(537) <= not(inputs(244));
    layer0_outputs(538) <= (inputs(29)) and (inputs(27));
    layer0_outputs(539) <= not((inputs(255)) xor (inputs(168)));
    layer0_outputs(540) <= not((inputs(163)) or (inputs(121)));
    layer0_outputs(541) <= (inputs(146)) or (inputs(248));
    layer0_outputs(542) <= (inputs(216)) and (inputs(216));
    layer0_outputs(543) <= (inputs(137)) xor (inputs(244));
    layer0_outputs(544) <= (inputs(46)) xor (inputs(218));
    layer0_outputs(545) <= not(inputs(2));
    layer0_outputs(546) <= not((inputs(173)) and (inputs(10)));
    layer0_outputs(547) <= inputs(233);
    layer0_outputs(548) <= inputs(145);
    layer0_outputs(549) <= (inputs(254)) xor (inputs(211));
    layer0_outputs(550) <= inputs(234);
    layer0_outputs(551) <= inputs(36);
    layer0_outputs(552) <= inputs(163);
    layer0_outputs(553) <= not(inputs(113));
    layer0_outputs(554) <= (inputs(13)) or (inputs(237));
    layer0_outputs(555) <= not(inputs(197));
    layer0_outputs(556) <= not(inputs(24)) or (inputs(81));
    layer0_outputs(557) <= inputs(126);
    layer0_outputs(558) <= (inputs(167)) and not (inputs(79));
    layer0_outputs(559) <= inputs(171);
    layer0_outputs(560) <= inputs(85);
    layer0_outputs(561) <= (inputs(234)) and (inputs(162));
    layer0_outputs(562) <= (inputs(149)) or (inputs(50));
    layer0_outputs(563) <= not(inputs(21));
    layer0_outputs(564) <= (inputs(67)) and not (inputs(143));
    layer0_outputs(565) <= (inputs(202)) or (inputs(206));
    layer0_outputs(566) <= '1';
    layer0_outputs(567) <= not(inputs(14)) or (inputs(127));
    layer0_outputs(568) <= (inputs(46)) and not (inputs(213));
    layer0_outputs(569) <= (inputs(139)) or (inputs(116));
    layer0_outputs(570) <= not(inputs(94));
    layer0_outputs(571) <= inputs(213);
    layer0_outputs(572) <= (inputs(23)) and not (inputs(178));
    layer0_outputs(573) <= inputs(249);
    layer0_outputs(574) <= not(inputs(140));
    layer0_outputs(575) <= not((inputs(4)) or (inputs(222)));
    layer0_outputs(576) <= (inputs(49)) or (inputs(67));
    layer0_outputs(577) <= not(inputs(157)) or (inputs(12));
    layer0_outputs(578) <= not((inputs(175)) or (inputs(244)));
    layer0_outputs(579) <= inputs(236);
    layer0_outputs(580) <= (inputs(248)) or (inputs(217));
    layer0_outputs(581) <= not((inputs(221)) xor (inputs(13)));
    layer0_outputs(582) <= inputs(120);
    layer0_outputs(583) <= (inputs(140)) or (inputs(223));
    layer0_outputs(584) <= not((inputs(239)) xor (inputs(139)));
    layer0_outputs(585) <= (inputs(177)) and not (inputs(128));
    layer0_outputs(586) <= (inputs(146)) or (inputs(251));
    layer0_outputs(587) <= not(inputs(166));
    layer0_outputs(588) <= inputs(205);
    layer0_outputs(589) <= (inputs(76)) or (inputs(195));
    layer0_outputs(590) <= not(inputs(226)) or (inputs(118));
    layer0_outputs(591) <= not(inputs(119));
    layer0_outputs(592) <= not(inputs(166)) or (inputs(114));
    layer0_outputs(593) <= not(inputs(58));
    layer0_outputs(594) <= (inputs(179)) or (inputs(91));
    layer0_outputs(595) <= not((inputs(110)) or (inputs(181)));
    layer0_outputs(596) <= (inputs(160)) or (inputs(109));
    layer0_outputs(597) <= (inputs(205)) or (inputs(89));
    layer0_outputs(598) <= not((inputs(113)) or (inputs(252)));
    layer0_outputs(599) <= inputs(227);
    layer0_outputs(600) <= inputs(216);
    layer0_outputs(601) <= not(inputs(129));
    layer0_outputs(602) <= (inputs(40)) and not (inputs(101));
    layer0_outputs(603) <= (inputs(246)) xor (inputs(96));
    layer0_outputs(604) <= not((inputs(31)) xor (inputs(245)));
    layer0_outputs(605) <= '0';
    layer0_outputs(606) <= (inputs(142)) xor (inputs(95));
    layer0_outputs(607) <= (inputs(245)) xor (inputs(218));
    layer0_outputs(608) <= inputs(160);
    layer0_outputs(609) <= inputs(237);
    layer0_outputs(610) <= not(inputs(94)) or (inputs(224));
    layer0_outputs(611) <= not((inputs(176)) and (inputs(131)));
    layer0_outputs(612) <= (inputs(34)) xor (inputs(129));
    layer0_outputs(613) <= inputs(109);
    layer0_outputs(614) <= not(inputs(219));
    layer0_outputs(615) <= (inputs(137)) or (inputs(241));
    layer0_outputs(616) <= not(inputs(137)) or (inputs(34));
    layer0_outputs(617) <= (inputs(239)) xor (inputs(3));
    layer0_outputs(618) <= not((inputs(7)) xor (inputs(208)));
    layer0_outputs(619) <= (inputs(111)) or (inputs(245));
    layer0_outputs(620) <= not(inputs(40));
    layer0_outputs(621) <= not(inputs(233));
    layer0_outputs(622) <= (inputs(36)) xor (inputs(186));
    layer0_outputs(623) <= not((inputs(14)) or (inputs(197)));
    layer0_outputs(624) <= not((inputs(174)) or (inputs(136)));
    layer0_outputs(625) <= not((inputs(43)) or (inputs(63)));
    layer0_outputs(626) <= (inputs(255)) or (inputs(119));
    layer0_outputs(627) <= not((inputs(236)) or (inputs(254)));
    layer0_outputs(628) <= not(inputs(59)) or (inputs(236));
    layer0_outputs(629) <= inputs(248);
    layer0_outputs(630) <= (inputs(110)) or (inputs(234));
    layer0_outputs(631) <= not(inputs(93)) or (inputs(120));
    layer0_outputs(632) <= not(inputs(128));
    layer0_outputs(633) <= inputs(41);
    layer0_outputs(634) <= (inputs(7)) xor (inputs(64));
    layer0_outputs(635) <= not(inputs(90));
    layer0_outputs(636) <= not(inputs(172)) or (inputs(108));
    layer0_outputs(637) <= not(inputs(146));
    layer0_outputs(638) <= not((inputs(240)) xor (inputs(12)));
    layer0_outputs(639) <= (inputs(208)) or (inputs(212));
    layer0_outputs(640) <= not(inputs(79)) or (inputs(29));
    layer0_outputs(641) <= (inputs(62)) and not (inputs(31));
    layer0_outputs(642) <= (inputs(60)) and not (inputs(219));
    layer0_outputs(643) <= inputs(23);
    layer0_outputs(644) <= inputs(148);
    layer0_outputs(645) <= not(inputs(83));
    layer0_outputs(646) <= not(inputs(1));
    layer0_outputs(647) <= inputs(92);
    layer0_outputs(648) <= not((inputs(53)) or (inputs(79)));
    layer0_outputs(649) <= (inputs(230)) and not (inputs(60));
    layer0_outputs(650) <= not(inputs(210));
    layer0_outputs(651) <= not(inputs(75)) or (inputs(237));
    layer0_outputs(652) <= (inputs(148)) and not (inputs(215));
    layer0_outputs(653) <= not((inputs(242)) or (inputs(78)));
    layer0_outputs(654) <= not(inputs(85)) or (inputs(108));
    layer0_outputs(655) <= not(inputs(231));
    layer0_outputs(656) <= not((inputs(164)) or (inputs(129)));
    layer0_outputs(657) <= not(inputs(79));
    layer0_outputs(658) <= (inputs(29)) or (inputs(233));
    layer0_outputs(659) <= '0';
    layer0_outputs(660) <= (inputs(86)) xor (inputs(114));
    layer0_outputs(661) <= not(inputs(180));
    layer0_outputs(662) <= (inputs(4)) or (inputs(94));
    layer0_outputs(663) <= (inputs(89)) and not (inputs(50));
    layer0_outputs(664) <= not((inputs(145)) or (inputs(115)));
    layer0_outputs(665) <= inputs(98);
    layer0_outputs(666) <= not((inputs(4)) or (inputs(91)));
    layer0_outputs(667) <= not(inputs(1)) or (inputs(237));
    layer0_outputs(668) <= (inputs(223)) or (inputs(85));
    layer0_outputs(669) <= inputs(85);
    layer0_outputs(670) <= inputs(39);
    layer0_outputs(671) <= not(inputs(38)) or (inputs(147));
    layer0_outputs(672) <= (inputs(166)) or (inputs(222));
    layer0_outputs(673) <= '1';
    layer0_outputs(674) <= (inputs(37)) and (inputs(89));
    layer0_outputs(675) <= not(inputs(99)) or (inputs(15));
    layer0_outputs(676) <= (inputs(2)) or (inputs(36));
    layer0_outputs(677) <= inputs(84);
    layer0_outputs(678) <= not(inputs(246)) or (inputs(0));
    layer0_outputs(679) <= not(inputs(54));
    layer0_outputs(680) <= inputs(247);
    layer0_outputs(681) <= not(inputs(85)) or (inputs(48));
    layer0_outputs(682) <= not(inputs(204));
    layer0_outputs(683) <= not(inputs(237)) or (inputs(143));
    layer0_outputs(684) <= not(inputs(24));
    layer0_outputs(685) <= inputs(8);
    layer0_outputs(686) <= (inputs(26)) and not (inputs(187));
    layer0_outputs(687) <= inputs(227);
    layer0_outputs(688) <= (inputs(107)) and not (inputs(126));
    layer0_outputs(689) <= (inputs(200)) or (inputs(133));
    layer0_outputs(690) <= (inputs(51)) or (inputs(96));
    layer0_outputs(691) <= not((inputs(119)) or (inputs(249)));
    layer0_outputs(692) <= not((inputs(192)) xor (inputs(42)));
    layer0_outputs(693) <= not((inputs(115)) or (inputs(142)));
    layer0_outputs(694) <= '1';
    layer0_outputs(695) <= not(inputs(223));
    layer0_outputs(696) <= not((inputs(180)) xor (inputs(88)));
    layer0_outputs(697) <= inputs(221);
    layer0_outputs(698) <= not(inputs(94));
    layer0_outputs(699) <= inputs(175);
    layer0_outputs(700) <= not(inputs(163));
    layer0_outputs(701) <= inputs(20);
    layer0_outputs(702) <= (inputs(178)) or (inputs(246));
    layer0_outputs(703) <= '1';
    layer0_outputs(704) <= not((inputs(33)) xor (inputs(91)));
    layer0_outputs(705) <= (inputs(126)) xor (inputs(107));
    layer0_outputs(706) <= not((inputs(249)) or (inputs(45)));
    layer0_outputs(707) <= not((inputs(182)) or (inputs(19)));
    layer0_outputs(708) <= (inputs(39)) or (inputs(230));
    layer0_outputs(709) <= not(inputs(231));
    layer0_outputs(710) <= (inputs(48)) or (inputs(94));
    layer0_outputs(711) <= (inputs(248)) or (inputs(27));
    layer0_outputs(712) <= (inputs(21)) and not (inputs(99));
    layer0_outputs(713) <= not(inputs(106)) or (inputs(49));
    layer0_outputs(714) <= not(inputs(38)) or (inputs(112));
    layer0_outputs(715) <= not(inputs(41)) or (inputs(168));
    layer0_outputs(716) <= inputs(107);
    layer0_outputs(717) <= (inputs(63)) or (inputs(215));
    layer0_outputs(718) <= not((inputs(119)) xor (inputs(241)));
    layer0_outputs(719) <= inputs(120);
    layer0_outputs(720) <= (inputs(124)) or (inputs(20));
    layer0_outputs(721) <= not((inputs(46)) and (inputs(42)));
    layer0_outputs(722) <= not(inputs(68)) or (inputs(192));
    layer0_outputs(723) <= inputs(88);
    layer0_outputs(724) <= not((inputs(3)) or (inputs(42)));
    layer0_outputs(725) <= not(inputs(68)) or (inputs(78));
    layer0_outputs(726) <= (inputs(70)) or (inputs(249));
    layer0_outputs(727) <= not(inputs(30)) or (inputs(57));
    layer0_outputs(728) <= inputs(186);
    layer0_outputs(729) <= (inputs(162)) and not (inputs(153));
    layer0_outputs(730) <= (inputs(244)) xor (inputs(4));
    layer0_outputs(731) <= (inputs(213)) or (inputs(140));
    layer0_outputs(732) <= inputs(9);
    layer0_outputs(733) <= not((inputs(130)) or (inputs(176)));
    layer0_outputs(734) <= (inputs(161)) xor (inputs(19));
    layer0_outputs(735) <= inputs(253);
    layer0_outputs(736) <= '1';
    layer0_outputs(737) <= (inputs(128)) or (inputs(177));
    layer0_outputs(738) <= not((inputs(80)) xor (inputs(105)));
    layer0_outputs(739) <= '1';
    layer0_outputs(740) <= not((inputs(173)) or (inputs(179)));
    layer0_outputs(741) <= not(inputs(130)) or (inputs(238));
    layer0_outputs(742) <= not(inputs(229));
    layer0_outputs(743) <= (inputs(86)) and (inputs(225));
    layer0_outputs(744) <= not(inputs(100)) or (inputs(225));
    layer0_outputs(745) <= not(inputs(79));
    layer0_outputs(746) <= not(inputs(116));
    layer0_outputs(747) <= (inputs(141)) or (inputs(108));
    layer0_outputs(748) <= not(inputs(75));
    layer0_outputs(749) <= not(inputs(86)) or (inputs(183));
    layer0_outputs(750) <= not(inputs(125));
    layer0_outputs(751) <= inputs(110);
    layer0_outputs(752) <= (inputs(129)) or (inputs(149));
    layer0_outputs(753) <= not(inputs(120));
    layer0_outputs(754) <= (inputs(2)) or (inputs(203));
    layer0_outputs(755) <= not((inputs(138)) or (inputs(49)));
    layer0_outputs(756) <= (inputs(35)) or (inputs(122));
    layer0_outputs(757) <= (inputs(158)) xor (inputs(26));
    layer0_outputs(758) <= (inputs(189)) or (inputs(169));
    layer0_outputs(759) <= not(inputs(72));
    layer0_outputs(760) <= inputs(120);
    layer0_outputs(761) <= not(inputs(165)) or (inputs(125));
    layer0_outputs(762) <= not((inputs(181)) xor (inputs(226)));
    layer0_outputs(763) <= not(inputs(181));
    layer0_outputs(764) <= not(inputs(89)) or (inputs(144));
    layer0_outputs(765) <= not(inputs(167));
    layer0_outputs(766) <= not((inputs(231)) or (inputs(65)));
    layer0_outputs(767) <= not((inputs(41)) or (inputs(1)));
    layer0_outputs(768) <= (inputs(255)) and not (inputs(36));
    layer0_outputs(769) <= not((inputs(223)) xor (inputs(85)));
    layer0_outputs(770) <= not((inputs(26)) and (inputs(25)));
    layer0_outputs(771) <= not(inputs(25)) or (inputs(1));
    layer0_outputs(772) <= (inputs(69)) and not (inputs(154));
    layer0_outputs(773) <= not(inputs(194)) or (inputs(3));
    layer0_outputs(774) <= not(inputs(181));
    layer0_outputs(775) <= (inputs(38)) and not (inputs(129));
    layer0_outputs(776) <= not(inputs(240)) or (inputs(127));
    layer0_outputs(777) <= not((inputs(179)) or (inputs(110)));
    layer0_outputs(778) <= (inputs(138)) or (inputs(52));
    layer0_outputs(779) <= not(inputs(163));
    layer0_outputs(780) <= inputs(156);
    layer0_outputs(781) <= not((inputs(91)) or (inputs(57)));
    layer0_outputs(782) <= not((inputs(131)) or (inputs(99)));
    layer0_outputs(783) <= not((inputs(74)) or (inputs(110)));
    layer0_outputs(784) <= (inputs(175)) or (inputs(93));
    layer0_outputs(785) <= not((inputs(217)) or (inputs(223)));
    layer0_outputs(786) <= '1';
    layer0_outputs(787) <= (inputs(183)) xor (inputs(136));
    layer0_outputs(788) <= (inputs(49)) or (inputs(43));
    layer0_outputs(789) <= inputs(150);
    layer0_outputs(790) <= (inputs(198)) or (inputs(255));
    layer0_outputs(791) <= not(inputs(126));
    layer0_outputs(792) <= inputs(150);
    layer0_outputs(793) <= not(inputs(19));
    layer0_outputs(794) <= (inputs(61)) or (inputs(23));
    layer0_outputs(795) <= (inputs(89)) or (inputs(250));
    layer0_outputs(796) <= not(inputs(22)) or (inputs(101));
    layer0_outputs(797) <= inputs(107);
    layer0_outputs(798) <= not((inputs(193)) or (inputs(220)));
    layer0_outputs(799) <= (inputs(194)) and not (inputs(2));
    layer0_outputs(800) <= (inputs(59)) and (inputs(59));
    layer0_outputs(801) <= not((inputs(31)) or (inputs(96)));
    layer0_outputs(802) <= inputs(100);
    layer0_outputs(803) <= not(inputs(132));
    layer0_outputs(804) <= not(inputs(233));
    layer0_outputs(805) <= inputs(201);
    layer0_outputs(806) <= (inputs(159)) or (inputs(29));
    layer0_outputs(807) <= (inputs(209)) and not (inputs(96));
    layer0_outputs(808) <= (inputs(29)) and not (inputs(55));
    layer0_outputs(809) <= not((inputs(1)) and (inputs(46)));
    layer0_outputs(810) <= not(inputs(23));
    layer0_outputs(811) <= not(inputs(85)) or (inputs(190));
    layer0_outputs(812) <= not(inputs(63));
    layer0_outputs(813) <= not(inputs(39));
    layer0_outputs(814) <= inputs(88);
    layer0_outputs(815) <= (inputs(201)) or (inputs(16));
    layer0_outputs(816) <= (inputs(125)) and not (inputs(252));
    layer0_outputs(817) <= inputs(32);
    layer0_outputs(818) <= (inputs(212)) and not (inputs(22));
    layer0_outputs(819) <= not(inputs(162));
    layer0_outputs(820) <= (inputs(92)) and not (inputs(89));
    layer0_outputs(821) <= not((inputs(0)) xor (inputs(57)));
    layer0_outputs(822) <= '1';
    layer0_outputs(823) <= (inputs(101)) and not (inputs(193));
    layer0_outputs(824) <= not((inputs(100)) xor (inputs(120)));
    layer0_outputs(825) <= not((inputs(136)) xor (inputs(147)));
    layer0_outputs(826) <= not((inputs(75)) or (inputs(65)));
    layer0_outputs(827) <= (inputs(192)) or (inputs(92));
    layer0_outputs(828) <= not((inputs(218)) or (inputs(203)));
    layer0_outputs(829) <= inputs(82);
    layer0_outputs(830) <= not(inputs(239));
    layer0_outputs(831) <= not((inputs(10)) xor (inputs(1)));
    layer0_outputs(832) <= not(inputs(68));
    layer0_outputs(833) <= (inputs(88)) and not (inputs(111));
    layer0_outputs(834) <= (inputs(92)) or (inputs(105));
    layer0_outputs(835) <= (inputs(203)) and not (inputs(66));
    layer0_outputs(836) <= not(inputs(136));
    layer0_outputs(837) <= (inputs(118)) and not (inputs(127));
    layer0_outputs(838) <= not((inputs(207)) or (inputs(134)));
    layer0_outputs(839) <= (inputs(87)) and not (inputs(238));
    layer0_outputs(840) <= (inputs(150)) or (inputs(83));
    layer0_outputs(841) <= not(inputs(18));
    layer0_outputs(842) <= (inputs(173)) or (inputs(174));
    layer0_outputs(843) <= not(inputs(121)) or (inputs(155));
    layer0_outputs(844) <= not(inputs(152));
    layer0_outputs(845) <= not(inputs(91));
    layer0_outputs(846) <= not(inputs(121));
    layer0_outputs(847) <= not(inputs(42)) or (inputs(223));
    layer0_outputs(848) <= inputs(135);
    layer0_outputs(849) <= inputs(145);
    layer0_outputs(850) <= not(inputs(183));
    layer0_outputs(851) <= not((inputs(61)) xor (inputs(65)));
    layer0_outputs(852) <= (inputs(162)) or (inputs(251));
    layer0_outputs(853) <= not(inputs(76)) or (inputs(19));
    layer0_outputs(854) <= not(inputs(67));
    layer0_outputs(855) <= (inputs(234)) or (inputs(227));
    layer0_outputs(856) <= (inputs(185)) or (inputs(64));
    layer0_outputs(857) <= (inputs(78)) xor (inputs(223));
    layer0_outputs(858) <= not(inputs(86));
    layer0_outputs(859) <= not((inputs(82)) or (inputs(43)));
    layer0_outputs(860) <= not((inputs(17)) or (inputs(116)));
    layer0_outputs(861) <= (inputs(149)) or (inputs(210));
    layer0_outputs(862) <= not((inputs(32)) or (inputs(225)));
    layer0_outputs(863) <= (inputs(105)) and not (inputs(130));
    layer0_outputs(864) <= inputs(94);
    layer0_outputs(865) <= not(inputs(52)) or (inputs(219));
    layer0_outputs(866) <= not((inputs(172)) xor (inputs(107)));
    layer0_outputs(867) <= inputs(114);
    layer0_outputs(868) <= (inputs(168)) and not (inputs(92));
    layer0_outputs(869) <= (inputs(20)) or (inputs(45));
    layer0_outputs(870) <= not((inputs(138)) xor (inputs(200)));
    layer0_outputs(871) <= not((inputs(56)) or (inputs(245)));
    layer0_outputs(872) <= not((inputs(23)) or (inputs(186)));
    layer0_outputs(873) <= not((inputs(118)) and (inputs(75)));
    layer0_outputs(874) <= not(inputs(226));
    layer0_outputs(875) <= (inputs(14)) or (inputs(169));
    layer0_outputs(876) <= not((inputs(204)) or (inputs(162)));
    layer0_outputs(877) <= not((inputs(95)) or (inputs(190)));
    layer0_outputs(878) <= not((inputs(112)) xor (inputs(241)));
    layer0_outputs(879) <= (inputs(87)) or (inputs(233));
    layer0_outputs(880) <= inputs(193);
    layer0_outputs(881) <= not(inputs(184)) or (inputs(120));
    layer0_outputs(882) <= inputs(41);
    layer0_outputs(883) <= not(inputs(30)) or (inputs(243));
    layer0_outputs(884) <= not((inputs(49)) xor (inputs(88)));
    layer0_outputs(885) <= (inputs(168)) and not (inputs(89));
    layer0_outputs(886) <= not((inputs(197)) xor (inputs(61)));
    layer0_outputs(887) <= not(inputs(137));
    layer0_outputs(888) <= inputs(181);
    layer0_outputs(889) <= not(inputs(13));
    layer0_outputs(890) <= (inputs(139)) or (inputs(7));
    layer0_outputs(891) <= inputs(145);
    layer0_outputs(892) <= inputs(166);
    layer0_outputs(893) <= inputs(217);
    layer0_outputs(894) <= (inputs(195)) and (inputs(184));
    layer0_outputs(895) <= not(inputs(15)) or (inputs(165));
    layer0_outputs(896) <= not((inputs(18)) or (inputs(223)));
    layer0_outputs(897) <= not((inputs(251)) xor (inputs(227)));
    layer0_outputs(898) <= inputs(226);
    layer0_outputs(899) <= not(inputs(5)) or (inputs(72));
    layer0_outputs(900) <= not(inputs(9)) or (inputs(230));
    layer0_outputs(901) <= inputs(215);
    layer0_outputs(902) <= not((inputs(202)) and (inputs(22)));
    layer0_outputs(903) <= not((inputs(99)) xor (inputs(85)));
    layer0_outputs(904) <= (inputs(28)) xor (inputs(46));
    layer0_outputs(905) <= not((inputs(183)) and (inputs(77)));
    layer0_outputs(906) <= not(inputs(195));
    layer0_outputs(907) <= (inputs(199)) or (inputs(144));
    layer0_outputs(908) <= '0';
    layer0_outputs(909) <= inputs(123);
    layer0_outputs(910) <= (inputs(49)) or (inputs(191));
    layer0_outputs(911) <= not((inputs(19)) or (inputs(84)));
    layer0_outputs(912) <= (inputs(42)) or (inputs(159));
    layer0_outputs(913) <= (inputs(25)) xor (inputs(100));
    layer0_outputs(914) <= (inputs(213)) or (inputs(244));
    layer0_outputs(915) <= (inputs(231)) or (inputs(62));
    layer0_outputs(916) <= inputs(249);
    layer0_outputs(917) <= inputs(101);
    layer0_outputs(918) <= not((inputs(219)) or (inputs(132)));
    layer0_outputs(919) <= not(inputs(132));
    layer0_outputs(920) <= inputs(91);
    layer0_outputs(921) <= not(inputs(65)) or (inputs(9));
    layer0_outputs(922) <= not((inputs(201)) or (inputs(90)));
    layer0_outputs(923) <= not((inputs(232)) xor (inputs(202)));
    layer0_outputs(924) <= not((inputs(42)) or (inputs(223)));
    layer0_outputs(925) <= not(inputs(54)) or (inputs(61));
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= not(inputs(159));
    layer0_outputs(928) <= (inputs(28)) or (inputs(75));
    layer0_outputs(929) <= not(inputs(105)) or (inputs(196));
    layer0_outputs(930) <= (inputs(124)) xor (inputs(191));
    layer0_outputs(931) <= (inputs(64)) or (inputs(24));
    layer0_outputs(932) <= (inputs(199)) and not (inputs(45));
    layer0_outputs(933) <= not((inputs(145)) xor (inputs(198)));
    layer0_outputs(934) <= not(inputs(55));
    layer0_outputs(935) <= not(inputs(251)) or (inputs(28));
    layer0_outputs(936) <= not(inputs(166));
    layer0_outputs(937) <= not(inputs(183)) or (inputs(33));
    layer0_outputs(938) <= not((inputs(194)) or (inputs(115)));
    layer0_outputs(939) <= inputs(219);
    layer0_outputs(940) <= not((inputs(177)) or (inputs(248)));
    layer0_outputs(941) <= (inputs(82)) or (inputs(233));
    layer0_outputs(942) <= inputs(234);
    layer0_outputs(943) <= not(inputs(179)) or (inputs(32));
    layer0_outputs(944) <= inputs(235);
    layer0_outputs(945) <= '1';
    layer0_outputs(946) <= (inputs(119)) and not (inputs(206));
    layer0_outputs(947) <= not((inputs(84)) or (inputs(25)));
    layer0_outputs(948) <= (inputs(19)) and not (inputs(205));
    layer0_outputs(949) <= (inputs(119)) or (inputs(47));
    layer0_outputs(950) <= (inputs(148)) xor (inputs(130));
    layer0_outputs(951) <= not((inputs(5)) or (inputs(146)));
    layer0_outputs(952) <= not(inputs(103));
    layer0_outputs(953) <= not((inputs(147)) or (inputs(126)));
    layer0_outputs(954) <= (inputs(56)) xor (inputs(232));
    layer0_outputs(955) <= not(inputs(188));
    layer0_outputs(956) <= inputs(51);
    layer0_outputs(957) <= not(inputs(229)) or (inputs(127));
    layer0_outputs(958) <= (inputs(234)) and not (inputs(170));
    layer0_outputs(959) <= (inputs(232)) or (inputs(130));
    layer0_outputs(960) <= not(inputs(94)) or (inputs(49));
    layer0_outputs(961) <= inputs(158);
    layer0_outputs(962) <= not((inputs(213)) xor (inputs(1)));
    layer0_outputs(963) <= not(inputs(182));
    layer0_outputs(964) <= not(inputs(136)) or (inputs(18));
    layer0_outputs(965) <= (inputs(155)) and not (inputs(125));
    layer0_outputs(966) <= (inputs(184)) or (inputs(21));
    layer0_outputs(967) <= not(inputs(22)) or (inputs(202));
    layer0_outputs(968) <= not(inputs(38)) or (inputs(101));
    layer0_outputs(969) <= (inputs(217)) and (inputs(52));
    layer0_outputs(970) <= (inputs(105)) or (inputs(66));
    layer0_outputs(971) <= (inputs(21)) and not (inputs(162));
    layer0_outputs(972) <= (inputs(139)) and not (inputs(80));
    layer0_outputs(973) <= inputs(35);
    layer0_outputs(974) <= (inputs(139)) and not (inputs(66));
    layer0_outputs(975) <= not(inputs(8)) or (inputs(104));
    layer0_outputs(976) <= not(inputs(166));
    layer0_outputs(977) <= (inputs(68)) and (inputs(184));
    layer0_outputs(978) <= (inputs(179)) and not (inputs(45));
    layer0_outputs(979) <= not(inputs(164));
    layer0_outputs(980) <= '0';
    layer0_outputs(981) <= not(inputs(18)) or (inputs(113));
    layer0_outputs(982) <= (inputs(19)) or (inputs(195));
    layer0_outputs(983) <= not(inputs(232));
    layer0_outputs(984) <= (inputs(192)) or (inputs(149));
    layer0_outputs(985) <= inputs(125);
    layer0_outputs(986) <= not(inputs(26));
    layer0_outputs(987) <= (inputs(247)) xor (inputs(237));
    layer0_outputs(988) <= not(inputs(98)) or (inputs(174));
    layer0_outputs(989) <= inputs(181);
    layer0_outputs(990) <= (inputs(121)) and not (inputs(249));
    layer0_outputs(991) <= (inputs(41)) or (inputs(54));
    layer0_outputs(992) <= inputs(180);
    layer0_outputs(993) <= not(inputs(163));
    layer0_outputs(994) <= (inputs(218)) xor (inputs(193));
    layer0_outputs(995) <= not((inputs(211)) xor (inputs(175)));
    layer0_outputs(996) <= inputs(236);
    layer0_outputs(997) <= not(inputs(184));
    layer0_outputs(998) <= (inputs(79)) or (inputs(212));
    layer0_outputs(999) <= inputs(150);
    layer0_outputs(1000) <= not((inputs(85)) or (inputs(101)));
    layer0_outputs(1001) <= not(inputs(84));
    layer0_outputs(1002) <= (inputs(172)) and not (inputs(0));
    layer0_outputs(1003) <= (inputs(6)) xor (inputs(223));
    layer0_outputs(1004) <= (inputs(199)) or (inputs(47));
    layer0_outputs(1005) <= inputs(97);
    layer0_outputs(1006) <= (inputs(203)) and not (inputs(91));
    layer0_outputs(1007) <= inputs(206);
    layer0_outputs(1008) <= '1';
    layer0_outputs(1009) <= inputs(73);
    layer0_outputs(1010) <= not((inputs(182)) xor (inputs(89)));
    layer0_outputs(1011) <= (inputs(95)) xor (inputs(34));
    layer0_outputs(1012) <= (inputs(148)) and not (inputs(240));
    layer0_outputs(1013) <= inputs(76);
    layer0_outputs(1014) <= not(inputs(163)) or (inputs(74));
    layer0_outputs(1015) <= (inputs(154)) or (inputs(0));
    layer0_outputs(1016) <= not((inputs(25)) or (inputs(241)));
    layer0_outputs(1017) <= (inputs(40)) or (inputs(220));
    layer0_outputs(1018) <= (inputs(156)) or (inputs(82));
    layer0_outputs(1019) <= not((inputs(36)) or (inputs(19)));
    layer0_outputs(1020) <= not(inputs(136));
    layer0_outputs(1021) <= inputs(247);
    layer0_outputs(1022) <= not(inputs(222));
    layer0_outputs(1023) <= (inputs(166)) or (inputs(235));
    layer0_outputs(1024) <= (inputs(8)) xor (inputs(25));
    layer0_outputs(1025) <= not(inputs(228)) or (inputs(110));
    layer0_outputs(1026) <= '0';
    layer0_outputs(1027) <= not((inputs(152)) or (inputs(243)));
    layer0_outputs(1028) <= not((inputs(55)) xor (inputs(34)));
    layer0_outputs(1029) <= (inputs(248)) and (inputs(235));
    layer0_outputs(1030) <= not((inputs(171)) xor (inputs(219)));
    layer0_outputs(1031) <= (inputs(52)) xor (inputs(13));
    layer0_outputs(1032) <= not(inputs(77));
    layer0_outputs(1033) <= (inputs(86)) and (inputs(58));
    layer0_outputs(1034) <= (inputs(169)) xor (inputs(120));
    layer0_outputs(1035) <= not(inputs(149));
    layer0_outputs(1036) <= not(inputs(189));
    layer0_outputs(1037) <= not((inputs(224)) or (inputs(218)));
    layer0_outputs(1038) <= not((inputs(150)) or (inputs(64)));
    layer0_outputs(1039) <= (inputs(51)) and (inputs(253));
    layer0_outputs(1040) <= not((inputs(232)) and (inputs(163)));
    layer0_outputs(1041) <= inputs(247);
    layer0_outputs(1042) <= not((inputs(131)) or (inputs(254)));
    layer0_outputs(1043) <= not(inputs(219));
    layer0_outputs(1044) <= inputs(107);
    layer0_outputs(1045) <= not(inputs(74));
    layer0_outputs(1046) <= (inputs(84)) or (inputs(127));
    layer0_outputs(1047) <= (inputs(244)) or (inputs(3));
    layer0_outputs(1048) <= inputs(207);
    layer0_outputs(1049) <= not(inputs(202));
    layer0_outputs(1050) <= not((inputs(36)) or (inputs(147)));
    layer0_outputs(1051) <= not((inputs(225)) xor (inputs(184)));
    layer0_outputs(1052) <= not(inputs(197));
    layer0_outputs(1053) <= not(inputs(52));
    layer0_outputs(1054) <= inputs(246);
    layer0_outputs(1055) <= (inputs(223)) and not (inputs(32));
    layer0_outputs(1056) <= inputs(163);
    layer0_outputs(1057) <= not(inputs(249));
    layer0_outputs(1058) <= (inputs(34)) or (inputs(27));
    layer0_outputs(1059) <= (inputs(73)) xor (inputs(120));
    layer0_outputs(1060) <= not(inputs(167)) or (inputs(46));
    layer0_outputs(1061) <= inputs(88);
    layer0_outputs(1062) <= (inputs(67)) or (inputs(221));
    layer0_outputs(1063) <= not(inputs(114));
    layer0_outputs(1064) <= (inputs(102)) and not (inputs(222));
    layer0_outputs(1065) <= inputs(22);
    layer0_outputs(1066) <= inputs(37);
    layer0_outputs(1067) <= not(inputs(151));
    layer0_outputs(1068) <= inputs(142);
    layer0_outputs(1069) <= inputs(92);
    layer0_outputs(1070) <= inputs(165);
    layer0_outputs(1071) <= not(inputs(116));
    layer0_outputs(1072) <= (inputs(123)) and not (inputs(236));
    layer0_outputs(1073) <= not((inputs(46)) and (inputs(42)));
    layer0_outputs(1074) <= inputs(158);
    layer0_outputs(1075) <= inputs(248);
    layer0_outputs(1076) <= (inputs(207)) or (inputs(186));
    layer0_outputs(1077) <= inputs(230);
    layer0_outputs(1078) <= not((inputs(81)) or (inputs(254)));
    layer0_outputs(1079) <= not(inputs(69));
    layer0_outputs(1080) <= not((inputs(161)) and (inputs(170)));
    layer0_outputs(1081) <= (inputs(216)) and not (inputs(83));
    layer0_outputs(1082) <= not(inputs(69)) or (inputs(110));
    layer0_outputs(1083) <= (inputs(56)) xor (inputs(24));
    layer0_outputs(1084) <= (inputs(95)) or (inputs(211));
    layer0_outputs(1085) <= not(inputs(93)) or (inputs(59));
    layer0_outputs(1086) <= not(inputs(109));
    layer0_outputs(1087) <= (inputs(160)) and not (inputs(123));
    layer0_outputs(1088) <= not((inputs(45)) or (inputs(123)));
    layer0_outputs(1089) <= not(inputs(65)) or (inputs(58));
    layer0_outputs(1090) <= not(inputs(198)) or (inputs(159));
    layer0_outputs(1091) <= not(inputs(24));
    layer0_outputs(1092) <= inputs(166);
    layer0_outputs(1093) <= not(inputs(60)) or (inputs(238));
    layer0_outputs(1094) <= not(inputs(47));
    layer0_outputs(1095) <= not((inputs(133)) xor (inputs(130)));
    layer0_outputs(1096) <= (inputs(115)) and not (inputs(16));
    layer0_outputs(1097) <= not(inputs(102));
    layer0_outputs(1098) <= not(inputs(191)) or (inputs(83));
    layer0_outputs(1099) <= (inputs(72)) or (inputs(200));
    layer0_outputs(1100) <= (inputs(13)) or (inputs(225));
    layer0_outputs(1101) <= (inputs(75)) or (inputs(253));
    layer0_outputs(1102) <= (inputs(145)) or (inputs(15));
    layer0_outputs(1103) <= not(inputs(88)) or (inputs(108));
    layer0_outputs(1104) <= (inputs(4)) and not (inputs(117));
    layer0_outputs(1105) <= not(inputs(7)) or (inputs(222));
    layer0_outputs(1106) <= (inputs(166)) and not (inputs(177));
    layer0_outputs(1107) <= inputs(158);
    layer0_outputs(1108) <= (inputs(109)) xor (inputs(107));
    layer0_outputs(1109) <= not((inputs(72)) and (inputs(151)));
    layer0_outputs(1110) <= not(inputs(199)) or (inputs(53));
    layer0_outputs(1111) <= inputs(215);
    layer0_outputs(1112) <= not(inputs(155)) or (inputs(155));
    layer0_outputs(1113) <= inputs(231);
    layer0_outputs(1114) <= not(inputs(75)) or (inputs(134));
    layer0_outputs(1115) <= not((inputs(253)) or (inputs(232)));
    layer0_outputs(1116) <= not((inputs(61)) and (inputs(194)));
    layer0_outputs(1117) <= inputs(139);
    layer0_outputs(1118) <= not((inputs(254)) xor (inputs(162)));
    layer0_outputs(1119) <= not((inputs(114)) xor (inputs(85)));
    layer0_outputs(1120) <= not((inputs(94)) or (inputs(86)));
    layer0_outputs(1121) <= not(inputs(227));
    layer0_outputs(1122) <= inputs(180);
    layer0_outputs(1123) <= not(inputs(23));
    layer0_outputs(1124) <= not(inputs(26));
    layer0_outputs(1125) <= inputs(77);
    layer0_outputs(1126) <= not(inputs(174));
    layer0_outputs(1127) <= (inputs(96)) xor (inputs(186));
    layer0_outputs(1128) <= not(inputs(84));
    layer0_outputs(1129) <= not((inputs(245)) or (inputs(204)));
    layer0_outputs(1130) <= not(inputs(150));
    layer0_outputs(1131) <= inputs(216);
    layer0_outputs(1132) <= not(inputs(60)) or (inputs(121));
    layer0_outputs(1133) <= not(inputs(132)) or (inputs(33));
    layer0_outputs(1134) <= (inputs(130)) or (inputs(220));
    layer0_outputs(1135) <= not(inputs(103)) or (inputs(134));
    layer0_outputs(1136) <= (inputs(183)) and not (inputs(79));
    layer0_outputs(1137) <= (inputs(188)) or (inputs(46));
    layer0_outputs(1138) <= (inputs(172)) and not (inputs(127));
    layer0_outputs(1139) <= (inputs(23)) and not (inputs(63));
    layer0_outputs(1140) <= (inputs(17)) or (inputs(106));
    layer0_outputs(1141) <= (inputs(210)) and not (inputs(144));
    layer0_outputs(1142) <= not((inputs(191)) and (inputs(151)));
    layer0_outputs(1143) <= not((inputs(243)) or (inputs(192)));
    layer0_outputs(1144) <= (inputs(1)) and not (inputs(224));
    layer0_outputs(1145) <= (inputs(211)) xor (inputs(128));
    layer0_outputs(1146) <= inputs(246);
    layer0_outputs(1147) <= (inputs(249)) or (inputs(191));
    layer0_outputs(1148) <= (inputs(34)) and not (inputs(123));
    layer0_outputs(1149) <= (inputs(84)) or (inputs(47));
    layer0_outputs(1150) <= not(inputs(115)) or (inputs(205));
    layer0_outputs(1151) <= inputs(223);
    layer0_outputs(1152) <= not(inputs(156)) or (inputs(153));
    layer0_outputs(1153) <= not(inputs(196));
    layer0_outputs(1154) <= inputs(168);
    layer0_outputs(1155) <= (inputs(59)) or (inputs(133));
    layer0_outputs(1156) <= not(inputs(100));
    layer0_outputs(1157) <= not(inputs(14)) or (inputs(244));
    layer0_outputs(1158) <= (inputs(156)) or (inputs(157));
    layer0_outputs(1159) <= (inputs(186)) and not (inputs(238));
    layer0_outputs(1160) <= not((inputs(253)) or (inputs(118)));
    layer0_outputs(1161) <= '0';
    layer0_outputs(1162) <= (inputs(4)) and not (inputs(222));
    layer0_outputs(1163) <= (inputs(204)) or (inputs(142));
    layer0_outputs(1164) <= '1';
    layer0_outputs(1165) <= not((inputs(0)) or (inputs(64)));
    layer0_outputs(1166) <= (inputs(91)) xor (inputs(142));
    layer0_outputs(1167) <= not((inputs(123)) xor (inputs(175)));
    layer0_outputs(1168) <= inputs(244);
    layer0_outputs(1169) <= not((inputs(167)) and (inputs(166)));
    layer0_outputs(1170) <= not(inputs(231));
    layer0_outputs(1171) <= not((inputs(57)) and (inputs(189)));
    layer0_outputs(1172) <= '1';
    layer0_outputs(1173) <= not(inputs(141));
    layer0_outputs(1174) <= not(inputs(122)) or (inputs(196));
    layer0_outputs(1175) <= (inputs(246)) or (inputs(82));
    layer0_outputs(1176) <= (inputs(11)) xor (inputs(60));
    layer0_outputs(1177) <= not(inputs(248));
    layer0_outputs(1178) <= (inputs(21)) and not (inputs(252));
    layer0_outputs(1179) <= not(inputs(196));
    layer0_outputs(1180) <= inputs(64);
    layer0_outputs(1181) <= (inputs(179)) and not (inputs(248));
    layer0_outputs(1182) <= not(inputs(30));
    layer0_outputs(1183) <= not((inputs(204)) xor (inputs(87)));
    layer0_outputs(1184) <= (inputs(38)) and not (inputs(241));
    layer0_outputs(1185) <= (inputs(13)) and not (inputs(208));
    layer0_outputs(1186) <= not((inputs(182)) or (inputs(149)));
    layer0_outputs(1187) <= (inputs(36)) and not (inputs(118));
    layer0_outputs(1188) <= (inputs(83)) and not (inputs(16));
    layer0_outputs(1189) <= (inputs(11)) and (inputs(188));
    layer0_outputs(1190) <= not(inputs(209));
    layer0_outputs(1191) <= (inputs(67)) and not (inputs(232));
    layer0_outputs(1192) <= not(inputs(122)) or (inputs(238));
    layer0_outputs(1193) <= not((inputs(186)) or (inputs(186)));
    layer0_outputs(1194) <= not(inputs(101)) or (inputs(64));
    layer0_outputs(1195) <= not(inputs(67)) or (inputs(55));
    layer0_outputs(1196) <= '0';
    layer0_outputs(1197) <= not((inputs(41)) and (inputs(58)));
    layer0_outputs(1198) <= (inputs(233)) and (inputs(234));
    layer0_outputs(1199) <= not(inputs(29));
    layer0_outputs(1200) <= not((inputs(44)) xor (inputs(73)));
    layer0_outputs(1201) <= (inputs(209)) and not (inputs(15));
    layer0_outputs(1202) <= not((inputs(229)) xor (inputs(25)));
    layer0_outputs(1203) <= not((inputs(111)) or (inputs(241)));
    layer0_outputs(1204) <= '1';
    layer0_outputs(1205) <= not(inputs(166));
    layer0_outputs(1206) <= inputs(24);
    layer0_outputs(1207) <= (inputs(157)) and not (inputs(27));
    layer0_outputs(1208) <= inputs(6);
    layer0_outputs(1209) <= not(inputs(147)) or (inputs(125));
    layer0_outputs(1210) <= inputs(122);
    layer0_outputs(1211) <= (inputs(76)) or (inputs(66));
    layer0_outputs(1212) <= (inputs(2)) or (inputs(45));
    layer0_outputs(1213) <= (inputs(71)) and not (inputs(133));
    layer0_outputs(1214) <= (inputs(118)) and not (inputs(181));
    layer0_outputs(1215) <= (inputs(216)) and not (inputs(40));
    layer0_outputs(1216) <= (inputs(148)) or (inputs(183));
    layer0_outputs(1217) <= (inputs(204)) and not (inputs(1));
    layer0_outputs(1218) <= '0';
    layer0_outputs(1219) <= inputs(217);
    layer0_outputs(1220) <= (inputs(187)) and not (inputs(220));
    layer0_outputs(1221) <= not((inputs(102)) or (inputs(66)));
    layer0_outputs(1222) <= inputs(50);
    layer0_outputs(1223) <= inputs(146);
    layer0_outputs(1224) <= inputs(133);
    layer0_outputs(1225) <= not((inputs(245)) or (inputs(62)));
    layer0_outputs(1226) <= inputs(214);
    layer0_outputs(1227) <= inputs(232);
    layer0_outputs(1228) <= not(inputs(99));
    layer0_outputs(1229) <= (inputs(160)) xor (inputs(188));
    layer0_outputs(1230) <= inputs(185);
    layer0_outputs(1231) <= (inputs(246)) or (inputs(29));
    layer0_outputs(1232) <= not(inputs(110)) or (inputs(48));
    layer0_outputs(1233) <= (inputs(171)) and not (inputs(14));
    layer0_outputs(1234) <= not(inputs(120));
    layer0_outputs(1235) <= (inputs(223)) or (inputs(159));
    layer0_outputs(1236) <= '1';
    layer0_outputs(1237) <= inputs(1);
    layer0_outputs(1238) <= not((inputs(185)) or (inputs(227)));
    layer0_outputs(1239) <= (inputs(40)) and not (inputs(160));
    layer0_outputs(1240) <= (inputs(247)) and not (inputs(122));
    layer0_outputs(1241) <= not(inputs(154));
    layer0_outputs(1242) <= not(inputs(37));
    layer0_outputs(1243) <= (inputs(22)) or (inputs(40));
    layer0_outputs(1244) <= (inputs(39)) or (inputs(33));
    layer0_outputs(1245) <= inputs(76);
    layer0_outputs(1246) <= '0';
    layer0_outputs(1247) <= not((inputs(211)) or (inputs(245)));
    layer0_outputs(1248) <= not(inputs(150));
    layer0_outputs(1249) <= (inputs(146)) and not (inputs(93));
    layer0_outputs(1250) <= not(inputs(88)) or (inputs(94));
    layer0_outputs(1251) <= '1';
    layer0_outputs(1252) <= inputs(51);
    layer0_outputs(1253) <= inputs(135);
    layer0_outputs(1254) <= inputs(172);
    layer0_outputs(1255) <= inputs(245);
    layer0_outputs(1256) <= not(inputs(162));
    layer0_outputs(1257) <= inputs(84);
    layer0_outputs(1258) <= not(inputs(129)) or (inputs(2));
    layer0_outputs(1259) <= not((inputs(195)) or (inputs(158)));
    layer0_outputs(1260) <= (inputs(39)) and not (inputs(178));
    layer0_outputs(1261) <= inputs(5);
    layer0_outputs(1262) <= not(inputs(213)) or (inputs(95));
    layer0_outputs(1263) <= (inputs(224)) and not (inputs(155));
    layer0_outputs(1264) <= inputs(221);
    layer0_outputs(1265) <= (inputs(114)) and not (inputs(12));
    layer0_outputs(1266) <= not((inputs(139)) xor (inputs(172)));
    layer0_outputs(1267) <= not(inputs(44));
    layer0_outputs(1268) <= not(inputs(248));
    layer0_outputs(1269) <= not((inputs(140)) or (inputs(13)));
    layer0_outputs(1270) <= inputs(248);
    layer0_outputs(1271) <= not(inputs(117));
    layer0_outputs(1272) <= not((inputs(79)) or (inputs(38)));
    layer0_outputs(1273) <= (inputs(102)) and not (inputs(192));
    layer0_outputs(1274) <= not(inputs(228));
    layer0_outputs(1275) <= inputs(174);
    layer0_outputs(1276) <= inputs(211);
    layer0_outputs(1277) <= inputs(126);
    layer0_outputs(1278) <= (inputs(198)) and (inputs(0));
    layer0_outputs(1279) <= inputs(232);
    layer0_outputs(1280) <= not(inputs(136)) or (inputs(87));
    layer0_outputs(1281) <= inputs(99);
    layer0_outputs(1282) <= not((inputs(22)) or (inputs(153)));
    layer0_outputs(1283) <= inputs(115);
    layer0_outputs(1284) <= (inputs(96)) and not (inputs(3));
    layer0_outputs(1285) <= not(inputs(39));
    layer0_outputs(1286) <= not(inputs(136));
    layer0_outputs(1287) <= (inputs(22)) and not (inputs(242));
    layer0_outputs(1288) <= not(inputs(120));
    layer0_outputs(1289) <= not(inputs(22)) or (inputs(145));
    layer0_outputs(1290) <= not((inputs(30)) or (inputs(151)));
    layer0_outputs(1291) <= (inputs(21)) and (inputs(145));
    layer0_outputs(1292) <= not((inputs(82)) or (inputs(30)));
    layer0_outputs(1293) <= not((inputs(226)) or (inputs(17)));
    layer0_outputs(1294) <= not(inputs(43));
    layer0_outputs(1295) <= not(inputs(38));
    layer0_outputs(1296) <= (inputs(154)) xor (inputs(205));
    layer0_outputs(1297) <= not(inputs(37));
    layer0_outputs(1298) <= not((inputs(21)) or (inputs(45)));
    layer0_outputs(1299) <= not(inputs(190));
    layer0_outputs(1300) <= not(inputs(205));
    layer0_outputs(1301) <= '1';
    layer0_outputs(1302) <= (inputs(242)) and not (inputs(93));
    layer0_outputs(1303) <= inputs(58);
    layer0_outputs(1304) <= not(inputs(90));
    layer0_outputs(1305) <= not((inputs(202)) or (inputs(144)));
    layer0_outputs(1306) <= (inputs(177)) or (inputs(141));
    layer0_outputs(1307) <= not((inputs(11)) xor (inputs(21)));
    layer0_outputs(1308) <= not(inputs(23)) or (inputs(109));
    layer0_outputs(1309) <= (inputs(82)) xor (inputs(187));
    layer0_outputs(1310) <= not(inputs(109));
    layer0_outputs(1311) <= not(inputs(98));
    layer0_outputs(1312) <= inputs(159);
    layer0_outputs(1313) <= not(inputs(47));
    layer0_outputs(1314) <= (inputs(43)) and not (inputs(209));
    layer0_outputs(1315) <= (inputs(38)) and not (inputs(14));
    layer0_outputs(1316) <= inputs(110);
    layer0_outputs(1317) <= not(inputs(86)) or (inputs(62));
    layer0_outputs(1318) <= not((inputs(145)) xor (inputs(101)));
    layer0_outputs(1319) <= (inputs(230)) and not (inputs(131));
    layer0_outputs(1320) <= not(inputs(22));
    layer0_outputs(1321) <= (inputs(181)) and not (inputs(46));
    layer0_outputs(1322) <= (inputs(125)) or (inputs(179));
    layer0_outputs(1323) <= inputs(143);
    layer0_outputs(1324) <= (inputs(159)) or (inputs(201));
    layer0_outputs(1325) <= (inputs(28)) or (inputs(105));
    layer0_outputs(1326) <= not(inputs(40));
    layer0_outputs(1327) <= (inputs(78)) xor (inputs(238));
    layer0_outputs(1328) <= inputs(245);
    layer0_outputs(1329) <= not(inputs(175));
    layer0_outputs(1330) <= not(inputs(166));
    layer0_outputs(1331) <= not(inputs(121));
    layer0_outputs(1332) <= not((inputs(194)) xor (inputs(220)));
    layer0_outputs(1333) <= '1';
    layer0_outputs(1334) <= inputs(187);
    layer0_outputs(1335) <= not((inputs(145)) xor (inputs(115)));
    layer0_outputs(1336) <= inputs(80);
    layer0_outputs(1337) <= inputs(77);
    layer0_outputs(1338) <= not(inputs(120));
    layer0_outputs(1339) <= not((inputs(150)) or (inputs(204)));
    layer0_outputs(1340) <= not(inputs(130));
    layer0_outputs(1341) <= inputs(231);
    layer0_outputs(1342) <= not(inputs(87)) or (inputs(71));
    layer0_outputs(1343) <= not((inputs(4)) xor (inputs(57)));
    layer0_outputs(1344) <= (inputs(21)) xor (inputs(146));
    layer0_outputs(1345) <= not(inputs(221)) or (inputs(133));
    layer0_outputs(1346) <= (inputs(0)) and not (inputs(162));
    layer0_outputs(1347) <= not((inputs(127)) or (inputs(52)));
    layer0_outputs(1348) <= (inputs(178)) or (inputs(174));
    layer0_outputs(1349) <= not((inputs(90)) or (inputs(150)));
    layer0_outputs(1350) <= (inputs(40)) and not (inputs(24));
    layer0_outputs(1351) <= inputs(213);
    layer0_outputs(1352) <= (inputs(120)) and not (inputs(6));
    layer0_outputs(1353) <= (inputs(181)) or (inputs(79));
    layer0_outputs(1354) <= not(inputs(0));
    layer0_outputs(1355) <= not((inputs(168)) or (inputs(190)));
    layer0_outputs(1356) <= not(inputs(136)) or (inputs(194));
    layer0_outputs(1357) <= (inputs(80)) and (inputs(81));
    layer0_outputs(1358) <= inputs(126);
    layer0_outputs(1359) <= not(inputs(214));
    layer0_outputs(1360) <= not((inputs(129)) or (inputs(155)));
    layer0_outputs(1361) <= not((inputs(213)) or (inputs(221)));
    layer0_outputs(1362) <= not(inputs(217)) or (inputs(34));
    layer0_outputs(1363) <= (inputs(18)) or (inputs(155));
    layer0_outputs(1364) <= not((inputs(193)) xor (inputs(198)));
    layer0_outputs(1365) <= (inputs(172)) and (inputs(201));
    layer0_outputs(1366) <= not((inputs(228)) or (inputs(112)));
    layer0_outputs(1367) <= not((inputs(75)) xor (inputs(34)));
    layer0_outputs(1368) <= inputs(7);
    layer0_outputs(1369) <= (inputs(21)) and (inputs(200));
    layer0_outputs(1370) <= not((inputs(100)) xor (inputs(110)));
    layer0_outputs(1371) <= not(inputs(132));
    layer0_outputs(1372) <= inputs(69);
    layer0_outputs(1373) <= not(inputs(103));
    layer0_outputs(1374) <= inputs(249);
    layer0_outputs(1375) <= inputs(56);
    layer0_outputs(1376) <= inputs(91);
    layer0_outputs(1377) <= not(inputs(95));
    layer0_outputs(1378) <= not(inputs(206));
    layer0_outputs(1379) <= (inputs(45)) and not (inputs(228));
    layer0_outputs(1380) <= not(inputs(180));
    layer0_outputs(1381) <= not((inputs(9)) or (inputs(127)));
    layer0_outputs(1382) <= (inputs(233)) xor (inputs(224));
    layer0_outputs(1383) <= inputs(102);
    layer0_outputs(1384) <= (inputs(216)) or (inputs(16));
    layer0_outputs(1385) <= not(inputs(108));
    layer0_outputs(1386) <= not(inputs(114)) or (inputs(95));
    layer0_outputs(1387) <= not(inputs(89));
    layer0_outputs(1388) <= (inputs(54)) and not (inputs(216));
    layer0_outputs(1389) <= (inputs(99)) and not (inputs(74));
    layer0_outputs(1390) <= not((inputs(245)) or (inputs(124)));
    layer0_outputs(1391) <= not((inputs(1)) xor (inputs(248)));
    layer0_outputs(1392) <= inputs(194);
    layer0_outputs(1393) <= not(inputs(200)) or (inputs(5));
    layer0_outputs(1394) <= not((inputs(68)) or (inputs(15)));
    layer0_outputs(1395) <= '0';
    layer0_outputs(1396) <= (inputs(7)) and not (inputs(140));
    layer0_outputs(1397) <= (inputs(214)) or (inputs(244));
    layer0_outputs(1398) <= not(inputs(201)) or (inputs(119));
    layer0_outputs(1399) <= '0';
    layer0_outputs(1400) <= not(inputs(219)) or (inputs(31));
    layer0_outputs(1401) <= (inputs(25)) and (inputs(101));
    layer0_outputs(1402) <= not(inputs(124));
    layer0_outputs(1403) <= inputs(178);
    layer0_outputs(1404) <= (inputs(162)) or (inputs(177));
    layer0_outputs(1405) <= (inputs(27)) or (inputs(255));
    layer0_outputs(1406) <= inputs(84);
    layer0_outputs(1407) <= not(inputs(91));
    layer0_outputs(1408) <= (inputs(136)) or (inputs(207));
    layer0_outputs(1409) <= (inputs(94)) xor (inputs(168));
    layer0_outputs(1410) <= inputs(228);
    layer0_outputs(1411) <= (inputs(137)) xor (inputs(34));
    layer0_outputs(1412) <= not((inputs(158)) or (inputs(252)));
    layer0_outputs(1413) <= not((inputs(112)) xor (inputs(203)));
    layer0_outputs(1414) <= not((inputs(118)) xor (inputs(81)));
    layer0_outputs(1415) <= not((inputs(17)) or (inputs(242)));
    layer0_outputs(1416) <= not((inputs(139)) or (inputs(54)));
    layer0_outputs(1417) <= not(inputs(178));
    layer0_outputs(1418) <= not(inputs(151));
    layer0_outputs(1419) <= (inputs(37)) xor (inputs(38));
    layer0_outputs(1420) <= not(inputs(10));
    layer0_outputs(1421) <= not(inputs(68)) or (inputs(175));
    layer0_outputs(1422) <= not(inputs(255)) or (inputs(121));
    layer0_outputs(1423) <= not(inputs(104));
    layer0_outputs(1424) <= not(inputs(246)) or (inputs(151));
    layer0_outputs(1425) <= not(inputs(0)) or (inputs(111));
    layer0_outputs(1426) <= inputs(41);
    layer0_outputs(1427) <= (inputs(141)) or (inputs(76));
    layer0_outputs(1428) <= inputs(106);
    layer0_outputs(1429) <= inputs(168);
    layer0_outputs(1430) <= not(inputs(100));
    layer0_outputs(1431) <= not(inputs(60));
    layer0_outputs(1432) <= (inputs(225)) xor (inputs(233));
    layer0_outputs(1433) <= (inputs(239)) and (inputs(198));
    layer0_outputs(1434) <= not((inputs(108)) or (inputs(182)));
    layer0_outputs(1435) <= inputs(145);
    layer0_outputs(1436) <= inputs(233);
    layer0_outputs(1437) <= inputs(88);
    layer0_outputs(1438) <= not(inputs(131)) or (inputs(36));
    layer0_outputs(1439) <= not(inputs(224)) or (inputs(79));
    layer0_outputs(1440) <= not(inputs(142)) or (inputs(2));
    layer0_outputs(1441) <= inputs(0);
    layer0_outputs(1442) <= inputs(32);
    layer0_outputs(1443) <= not(inputs(167));
    layer0_outputs(1444) <= not((inputs(20)) or (inputs(227)));
    layer0_outputs(1445) <= inputs(221);
    layer0_outputs(1446) <= (inputs(13)) and not (inputs(209));
    layer0_outputs(1447) <= (inputs(129)) or (inputs(131));
    layer0_outputs(1448) <= '0';
    layer0_outputs(1449) <= inputs(247);
    layer0_outputs(1450) <= not(inputs(83));
    layer0_outputs(1451) <= not((inputs(253)) xor (inputs(28)));
    layer0_outputs(1452) <= not(inputs(53));
    layer0_outputs(1453) <= inputs(40);
    layer0_outputs(1454) <= (inputs(158)) xor (inputs(172));
    layer0_outputs(1455) <= not(inputs(118));
    layer0_outputs(1456) <= not((inputs(84)) xor (inputs(172)));
    layer0_outputs(1457) <= '1';
    layer0_outputs(1458) <= not(inputs(59));
    layer0_outputs(1459) <= inputs(52);
    layer0_outputs(1460) <= inputs(112);
    layer0_outputs(1461) <= not((inputs(171)) or (inputs(179)));
    layer0_outputs(1462) <= (inputs(199)) or (inputs(214));
    layer0_outputs(1463) <= not((inputs(43)) xor (inputs(191)));
    layer0_outputs(1464) <= (inputs(21)) or (inputs(193));
    layer0_outputs(1465) <= not(inputs(30));
    layer0_outputs(1466) <= '0';
    layer0_outputs(1467) <= not(inputs(41)) or (inputs(254));
    layer0_outputs(1468) <= (inputs(179)) or (inputs(221));
    layer0_outputs(1469) <= (inputs(74)) or (inputs(150));
    layer0_outputs(1470) <= (inputs(17)) and not (inputs(65));
    layer0_outputs(1471) <= not((inputs(218)) and (inputs(16)));
    layer0_outputs(1472) <= (inputs(40)) xor (inputs(243));
    layer0_outputs(1473) <= '0';
    layer0_outputs(1474) <= (inputs(97)) and not (inputs(158));
    layer0_outputs(1475) <= not(inputs(44)) or (inputs(144));
    layer0_outputs(1476) <= inputs(77);
    layer0_outputs(1477) <= not((inputs(32)) or (inputs(151)));
    layer0_outputs(1478) <= not((inputs(178)) or (inputs(114)));
    layer0_outputs(1479) <= not(inputs(201));
    layer0_outputs(1480) <= inputs(89);
    layer0_outputs(1481) <= not(inputs(179)) or (inputs(213));
    layer0_outputs(1482) <= not(inputs(61));
    layer0_outputs(1483) <= (inputs(86)) xor (inputs(24));
    layer0_outputs(1484) <= not(inputs(119)) or (inputs(165));
    layer0_outputs(1485) <= not((inputs(139)) or (inputs(106)));
    layer0_outputs(1486) <= (inputs(18)) xor (inputs(211));
    layer0_outputs(1487) <= not(inputs(5)) or (inputs(158));
    layer0_outputs(1488) <= (inputs(142)) or (inputs(246));
    layer0_outputs(1489) <= (inputs(237)) or (inputs(8));
    layer0_outputs(1490) <= not((inputs(125)) xor (inputs(189)));
    layer0_outputs(1491) <= not((inputs(166)) xor (inputs(229)));
    layer0_outputs(1492) <= (inputs(33)) xor (inputs(45));
    layer0_outputs(1493) <= (inputs(238)) xor (inputs(27));
    layer0_outputs(1494) <= inputs(244);
    layer0_outputs(1495) <= (inputs(246)) and not (inputs(78));
    layer0_outputs(1496) <= not(inputs(223)) or (inputs(159));
    layer0_outputs(1497) <= not((inputs(20)) or (inputs(238)));
    layer0_outputs(1498) <= not((inputs(190)) or (inputs(69)));
    layer0_outputs(1499) <= not((inputs(193)) and (inputs(113)));
    layer0_outputs(1500) <= not((inputs(80)) or (inputs(188)));
    layer0_outputs(1501) <= not((inputs(62)) xor (inputs(50)));
    layer0_outputs(1502) <= not((inputs(26)) or (inputs(225)));
    layer0_outputs(1503) <= (inputs(180)) or (inputs(238));
    layer0_outputs(1504) <= not((inputs(143)) and (inputs(192)));
    layer0_outputs(1505) <= (inputs(102)) or (inputs(183));
    layer0_outputs(1506) <= not(inputs(173)) or (inputs(131));
    layer0_outputs(1507) <= inputs(23);
    layer0_outputs(1508) <= (inputs(87)) or (inputs(191));
    layer0_outputs(1509) <= (inputs(89)) xor (inputs(86));
    layer0_outputs(1510) <= not(inputs(248));
    layer0_outputs(1511) <= not(inputs(199)) or (inputs(141));
    layer0_outputs(1512) <= not(inputs(248)) or (inputs(54));
    layer0_outputs(1513) <= (inputs(49)) or (inputs(66));
    layer0_outputs(1514) <= (inputs(117)) or (inputs(101));
    layer0_outputs(1515) <= not((inputs(77)) and (inputs(140)));
    layer0_outputs(1516) <= (inputs(153)) and (inputs(153));
    layer0_outputs(1517) <= (inputs(193)) xor (inputs(58));
    layer0_outputs(1518) <= not(inputs(116)) or (inputs(206));
    layer0_outputs(1519) <= not((inputs(239)) or (inputs(0)));
    layer0_outputs(1520) <= (inputs(60)) and (inputs(56));
    layer0_outputs(1521) <= inputs(222);
    layer0_outputs(1522) <= inputs(110);
    layer0_outputs(1523) <= not(inputs(215)) or (inputs(0));
    layer0_outputs(1524) <= not(inputs(104)) or (inputs(86));
    layer0_outputs(1525) <= (inputs(184)) and (inputs(122));
    layer0_outputs(1526) <= not((inputs(216)) and (inputs(182)));
    layer0_outputs(1527) <= not(inputs(130));
    layer0_outputs(1528) <= not(inputs(217));
    layer0_outputs(1529) <= not((inputs(57)) or (inputs(43)));
    layer0_outputs(1530) <= not(inputs(248)) or (inputs(254));
    layer0_outputs(1531) <= (inputs(255)) or (inputs(242));
    layer0_outputs(1532) <= not(inputs(192));
    layer0_outputs(1533) <= '1';
    layer0_outputs(1534) <= not(inputs(83));
    layer0_outputs(1535) <= (inputs(30)) and not (inputs(239));
    layer0_outputs(1536) <= not((inputs(12)) xor (inputs(145)));
    layer0_outputs(1537) <= not((inputs(34)) or (inputs(3)));
    layer0_outputs(1538) <= not(inputs(101));
    layer0_outputs(1539) <= (inputs(10)) xor (inputs(190));
    layer0_outputs(1540) <= inputs(25);
    layer0_outputs(1541) <= (inputs(134)) xor (inputs(171));
    layer0_outputs(1542) <= not(inputs(184)) or (inputs(181));
    layer0_outputs(1543) <= not(inputs(48));
    layer0_outputs(1544) <= inputs(193);
    layer0_outputs(1545) <= not(inputs(230)) or (inputs(77));
    layer0_outputs(1546) <= not(inputs(170));
    layer0_outputs(1547) <= not(inputs(231));
    layer0_outputs(1548) <= inputs(45);
    layer0_outputs(1549) <= not((inputs(5)) or (inputs(125)));
    layer0_outputs(1550) <= not((inputs(238)) xor (inputs(251)));
    layer0_outputs(1551) <= (inputs(212)) xor (inputs(144));
    layer0_outputs(1552) <= not((inputs(246)) xor (inputs(154)));
    layer0_outputs(1553) <= (inputs(95)) or (inputs(202));
    layer0_outputs(1554) <= (inputs(149)) or (inputs(147));
    layer0_outputs(1555) <= not(inputs(42)) or (inputs(115));
    layer0_outputs(1556) <= inputs(243);
    layer0_outputs(1557) <= not((inputs(152)) or (inputs(247)));
    layer0_outputs(1558) <= not(inputs(118)) or (inputs(92));
    layer0_outputs(1559) <= (inputs(139)) and not (inputs(132));
    layer0_outputs(1560) <= '0';
    layer0_outputs(1561) <= not(inputs(200));
    layer0_outputs(1562) <= not(inputs(151)) or (inputs(34));
    layer0_outputs(1563) <= not((inputs(217)) and (inputs(208)));
    layer0_outputs(1564) <= not(inputs(206));
    layer0_outputs(1565) <= not(inputs(77));
    layer0_outputs(1566) <= (inputs(92)) or (inputs(104));
    layer0_outputs(1567) <= (inputs(141)) and not (inputs(160));
    layer0_outputs(1568) <= not(inputs(75));
    layer0_outputs(1569) <= not((inputs(97)) xor (inputs(229)));
    layer0_outputs(1570) <= (inputs(118)) and not (inputs(239));
    layer0_outputs(1571) <= (inputs(118)) xor (inputs(168));
    layer0_outputs(1572) <= inputs(233);
    layer0_outputs(1573) <= not((inputs(124)) and (inputs(122)));
    layer0_outputs(1574) <= not(inputs(147));
    layer0_outputs(1575) <= inputs(90);
    layer0_outputs(1576) <= inputs(34);
    layer0_outputs(1577) <= '0';
    layer0_outputs(1578) <= not((inputs(172)) or (inputs(194)));
    layer0_outputs(1579) <= inputs(101);
    layer0_outputs(1580) <= not((inputs(50)) and (inputs(45)));
    layer0_outputs(1581) <= (inputs(229)) and not (inputs(116));
    layer0_outputs(1582) <= not((inputs(137)) xor (inputs(235)));
    layer0_outputs(1583) <= (inputs(132)) and (inputs(164));
    layer0_outputs(1584) <= '0';
    layer0_outputs(1585) <= (inputs(63)) and not (inputs(119));
    layer0_outputs(1586) <= not((inputs(157)) or (inputs(116)));
    layer0_outputs(1587) <= not(inputs(28)) or (inputs(210));
    layer0_outputs(1588) <= not(inputs(118)) or (inputs(49));
    layer0_outputs(1589) <= not(inputs(33));
    layer0_outputs(1590) <= not(inputs(180));
    layer0_outputs(1591) <= (inputs(71)) and not (inputs(151));
    layer0_outputs(1592) <= not(inputs(195)) or (inputs(81));
    layer0_outputs(1593) <= (inputs(174)) xor (inputs(35));
    layer0_outputs(1594) <= not(inputs(91));
    layer0_outputs(1595) <= not(inputs(105)) or (inputs(54));
    layer0_outputs(1596) <= (inputs(239)) or (inputs(93));
    layer0_outputs(1597) <= (inputs(163)) or (inputs(197));
    layer0_outputs(1598) <= '1';
    layer0_outputs(1599) <= (inputs(250)) and not (inputs(175));
    layer0_outputs(1600) <= not((inputs(134)) or (inputs(113)));
    layer0_outputs(1601) <= (inputs(205)) xor (inputs(79));
    layer0_outputs(1602) <= (inputs(129)) or (inputs(5));
    layer0_outputs(1603) <= (inputs(49)) or (inputs(238));
    layer0_outputs(1604) <= inputs(95);
    layer0_outputs(1605) <= (inputs(238)) or (inputs(202));
    layer0_outputs(1606) <= not((inputs(22)) xor (inputs(53)));
    layer0_outputs(1607) <= not((inputs(243)) and (inputs(37)));
    layer0_outputs(1608) <= (inputs(239)) xor (inputs(245));
    layer0_outputs(1609) <= not(inputs(182));
    layer0_outputs(1610) <= (inputs(20)) xor (inputs(48));
    layer0_outputs(1611) <= (inputs(199)) and not (inputs(51));
    layer0_outputs(1612) <= not((inputs(157)) or (inputs(13)));
    layer0_outputs(1613) <= inputs(193);
    layer0_outputs(1614) <= not((inputs(131)) or (inputs(65)));
    layer0_outputs(1615) <= inputs(144);
    layer0_outputs(1616) <= (inputs(229)) xor (inputs(238));
    layer0_outputs(1617) <= (inputs(50)) xor (inputs(76));
    layer0_outputs(1618) <= inputs(129);
    layer0_outputs(1619) <= (inputs(124)) and not (inputs(215));
    layer0_outputs(1620) <= not((inputs(199)) or (inputs(15)));
    layer0_outputs(1621) <= (inputs(211)) xor (inputs(50));
    layer0_outputs(1622) <= inputs(76);
    layer0_outputs(1623) <= (inputs(194)) and not (inputs(17));
    layer0_outputs(1624) <= (inputs(119)) and not (inputs(64));
    layer0_outputs(1625) <= not((inputs(12)) or (inputs(31)));
    layer0_outputs(1626) <= not(inputs(121)) or (inputs(28));
    layer0_outputs(1627) <= not((inputs(179)) or (inputs(35)));
    layer0_outputs(1628) <= inputs(10);
    layer0_outputs(1629) <= not(inputs(147));
    layer0_outputs(1630) <= (inputs(134)) xor (inputs(154));
    layer0_outputs(1631) <= not((inputs(132)) or (inputs(160)));
    layer0_outputs(1632) <= not((inputs(2)) or (inputs(171)));
    layer0_outputs(1633) <= (inputs(143)) and (inputs(56));
    layer0_outputs(1634) <= not((inputs(122)) or (inputs(134)));
    layer0_outputs(1635) <= not(inputs(231));
    layer0_outputs(1636) <= (inputs(253)) or (inputs(68));
    layer0_outputs(1637) <= (inputs(227)) xor (inputs(178));
    layer0_outputs(1638) <= (inputs(245)) and not (inputs(3));
    layer0_outputs(1639) <= not(inputs(218));
    layer0_outputs(1640) <= inputs(74);
    layer0_outputs(1641) <= not((inputs(30)) xor (inputs(58)));
    layer0_outputs(1642) <= inputs(66);
    layer0_outputs(1643) <= inputs(138);
    layer0_outputs(1644) <= inputs(71);
    layer0_outputs(1645) <= not((inputs(102)) xor (inputs(148)));
    layer0_outputs(1646) <= not((inputs(53)) or (inputs(36)));
    layer0_outputs(1647) <= inputs(24);
    layer0_outputs(1648) <= (inputs(47)) and not (inputs(151));
    layer0_outputs(1649) <= '1';
    layer0_outputs(1650) <= not(inputs(126));
    layer0_outputs(1651) <= not(inputs(49));
    layer0_outputs(1652) <= (inputs(30)) and (inputs(165));
    layer0_outputs(1653) <= not(inputs(150)) or (inputs(38));
    layer0_outputs(1654) <= not(inputs(71)) or (inputs(2));
    layer0_outputs(1655) <= inputs(97);
    layer0_outputs(1656) <= not(inputs(95));
    layer0_outputs(1657) <= not(inputs(102));
    layer0_outputs(1658) <= (inputs(169)) and not (inputs(73));
    layer0_outputs(1659) <= inputs(64);
    layer0_outputs(1660) <= not(inputs(211)) or (inputs(97));
    layer0_outputs(1661) <= not(inputs(150));
    layer0_outputs(1662) <= (inputs(33)) xor (inputs(148));
    layer0_outputs(1663) <= not(inputs(102)) or (inputs(114));
    layer0_outputs(1664) <= not(inputs(182)) or (inputs(51));
    layer0_outputs(1665) <= (inputs(12)) or (inputs(132));
    layer0_outputs(1666) <= inputs(25);
    layer0_outputs(1667) <= not((inputs(232)) or (inputs(81)));
    layer0_outputs(1668) <= (inputs(252)) or (inputs(89));
    layer0_outputs(1669) <= inputs(158);
    layer0_outputs(1670) <= (inputs(170)) or (inputs(165));
    layer0_outputs(1671) <= not(inputs(228));
    layer0_outputs(1672) <= (inputs(100)) and not (inputs(183));
    layer0_outputs(1673) <= inputs(180);
    layer0_outputs(1674) <= not((inputs(241)) or (inputs(245)));
    layer0_outputs(1675) <= inputs(55);
    layer0_outputs(1676) <= (inputs(112)) or (inputs(217));
    layer0_outputs(1677) <= not(inputs(77)) or (inputs(143));
    layer0_outputs(1678) <= not((inputs(141)) and (inputs(141)));
    layer0_outputs(1679) <= not(inputs(93));
    layer0_outputs(1680) <= not(inputs(161));
    layer0_outputs(1681) <= not(inputs(231));
    layer0_outputs(1682) <= '1';
    layer0_outputs(1683) <= not(inputs(68)) or (inputs(164));
    layer0_outputs(1684) <= (inputs(112)) xor (inputs(16));
    layer0_outputs(1685) <= inputs(229);
    layer0_outputs(1686) <= not(inputs(102));
    layer0_outputs(1687) <= not(inputs(196)) or (inputs(114));
    layer0_outputs(1688) <= not((inputs(198)) and (inputs(185)));
    layer0_outputs(1689) <= (inputs(246)) and not (inputs(223));
    layer0_outputs(1690) <= (inputs(59)) or (inputs(4));
    layer0_outputs(1691) <= inputs(22);
    layer0_outputs(1692) <= not((inputs(155)) xor (inputs(197)));
    layer0_outputs(1693) <= inputs(167);
    layer0_outputs(1694) <= (inputs(116)) or (inputs(5));
    layer0_outputs(1695) <= (inputs(254)) or (inputs(92));
    layer0_outputs(1696) <= (inputs(241)) and not (inputs(150));
    layer0_outputs(1697) <= not((inputs(189)) or (inputs(208)));
    layer0_outputs(1698) <= not(inputs(163));
    layer0_outputs(1699) <= (inputs(35)) and not (inputs(220));
    layer0_outputs(1700) <= not(inputs(181)) or (inputs(30));
    layer0_outputs(1701) <= (inputs(55)) or (inputs(174));
    layer0_outputs(1702) <= not(inputs(80)) or (inputs(123));
    layer0_outputs(1703) <= (inputs(10)) xor (inputs(163));
    layer0_outputs(1704) <= inputs(106);
    layer0_outputs(1705) <= not(inputs(27)) or (inputs(171));
    layer0_outputs(1706) <= not((inputs(206)) or (inputs(176)));
    layer0_outputs(1707) <= inputs(92);
    layer0_outputs(1708) <= (inputs(40)) xor (inputs(88));
    layer0_outputs(1709) <= (inputs(171)) xor (inputs(98));
    layer0_outputs(1710) <= inputs(11);
    layer0_outputs(1711) <= not(inputs(23));
    layer0_outputs(1712) <= not((inputs(47)) xor (inputs(63)));
    layer0_outputs(1713) <= not((inputs(189)) xor (inputs(10)));
    layer0_outputs(1714) <= not((inputs(197)) or (inputs(225)));
    layer0_outputs(1715) <= inputs(233);
    layer0_outputs(1716) <= not(inputs(144)) or (inputs(241));
    layer0_outputs(1717) <= inputs(23);
    layer0_outputs(1718) <= inputs(137);
    layer0_outputs(1719) <= (inputs(158)) xor (inputs(71));
    layer0_outputs(1720) <= not(inputs(230));
    layer0_outputs(1721) <= not((inputs(29)) xor (inputs(72)));
    layer0_outputs(1722) <= (inputs(74)) or (inputs(91));
    layer0_outputs(1723) <= not(inputs(17));
    layer0_outputs(1724) <= (inputs(24)) and (inputs(232));
    layer0_outputs(1725) <= inputs(254);
    layer0_outputs(1726) <= (inputs(19)) xor (inputs(253));
    layer0_outputs(1727) <= (inputs(243)) or (inputs(104));
    layer0_outputs(1728) <= (inputs(46)) or (inputs(205));
    layer0_outputs(1729) <= (inputs(209)) xor (inputs(171));
    layer0_outputs(1730) <= (inputs(159)) or (inputs(77));
    layer0_outputs(1731) <= inputs(190);
    layer0_outputs(1732) <= not(inputs(218)) or (inputs(52));
    layer0_outputs(1733) <= (inputs(7)) and not (inputs(80));
    layer0_outputs(1734) <= not((inputs(89)) or (inputs(224)));
    layer0_outputs(1735) <= inputs(232);
    layer0_outputs(1736) <= not(inputs(104));
    layer0_outputs(1737) <= (inputs(68)) and not (inputs(180));
    layer0_outputs(1738) <= (inputs(126)) and not (inputs(131));
    layer0_outputs(1739) <= (inputs(5)) or (inputs(233));
    layer0_outputs(1740) <= (inputs(5)) xor (inputs(79));
    layer0_outputs(1741) <= not(inputs(164));
    layer0_outputs(1742) <= inputs(96);
    layer0_outputs(1743) <= not(inputs(59));
    layer0_outputs(1744) <= not(inputs(184));
    layer0_outputs(1745) <= not(inputs(210));
    layer0_outputs(1746) <= not(inputs(127));
    layer0_outputs(1747) <= inputs(181);
    layer0_outputs(1748) <= (inputs(9)) or (inputs(8));
    layer0_outputs(1749) <= not(inputs(8));
    layer0_outputs(1750) <= not(inputs(51));
    layer0_outputs(1751) <= (inputs(134)) and not (inputs(93));
    layer0_outputs(1752) <= (inputs(153)) and not (inputs(16));
    layer0_outputs(1753) <= not(inputs(118));
    layer0_outputs(1754) <= (inputs(44)) and not (inputs(114));
    layer0_outputs(1755) <= not(inputs(90));
    layer0_outputs(1756) <= '0';
    layer0_outputs(1757) <= not(inputs(192));
    layer0_outputs(1758) <= inputs(118);
    layer0_outputs(1759) <= (inputs(150)) and not (inputs(57));
    layer0_outputs(1760) <= not((inputs(200)) xor (inputs(231)));
    layer0_outputs(1761) <= not(inputs(42)) or (inputs(18));
    layer0_outputs(1762) <= not(inputs(156));
    layer0_outputs(1763) <= inputs(229);
    layer0_outputs(1764) <= (inputs(132)) and not (inputs(221));
    layer0_outputs(1765) <= '0';
    layer0_outputs(1766) <= not((inputs(67)) or (inputs(246)));
    layer0_outputs(1767) <= (inputs(24)) and not (inputs(159));
    layer0_outputs(1768) <= not((inputs(241)) xor (inputs(80)));
    layer0_outputs(1769) <= inputs(62);
    layer0_outputs(1770) <= not(inputs(57));
    layer0_outputs(1771) <= not((inputs(237)) xor (inputs(9)));
    layer0_outputs(1772) <= (inputs(125)) or (inputs(214));
    layer0_outputs(1773) <= not(inputs(85));
    layer0_outputs(1774) <= (inputs(67)) or (inputs(79));
    layer0_outputs(1775) <= not((inputs(142)) xor (inputs(224)));
    layer0_outputs(1776) <= not((inputs(212)) or (inputs(175)));
    layer0_outputs(1777) <= not((inputs(26)) or (inputs(191)));
    layer0_outputs(1778) <= inputs(200);
    layer0_outputs(1779) <= not((inputs(58)) and (inputs(250)));
    layer0_outputs(1780) <= not(inputs(173));
    layer0_outputs(1781) <= not(inputs(243)) or (inputs(206));
    layer0_outputs(1782) <= (inputs(98)) xor (inputs(69));
    layer0_outputs(1783) <= not((inputs(185)) or (inputs(190)));
    layer0_outputs(1784) <= not((inputs(26)) or (inputs(38)));
    layer0_outputs(1785) <= (inputs(88)) and not (inputs(110));
    layer0_outputs(1786) <= inputs(172);
    layer0_outputs(1787) <= not(inputs(36));
    layer0_outputs(1788) <= (inputs(238)) and (inputs(54));
    layer0_outputs(1789) <= '1';
    layer0_outputs(1790) <= (inputs(18)) or (inputs(45));
    layer0_outputs(1791) <= not(inputs(211));
    layer0_outputs(1792) <= not((inputs(67)) or (inputs(111)));
    layer0_outputs(1793) <= (inputs(229)) or (inputs(206));
    layer0_outputs(1794) <= inputs(143);
    layer0_outputs(1795) <= not(inputs(91));
    layer0_outputs(1796) <= (inputs(74)) xor (inputs(106));
    layer0_outputs(1797) <= (inputs(250)) and not (inputs(91));
    layer0_outputs(1798) <= inputs(185);
    layer0_outputs(1799) <= (inputs(131)) and not (inputs(16));
    layer0_outputs(1800) <= not(inputs(162));
    layer0_outputs(1801) <= (inputs(203)) and not (inputs(83));
    layer0_outputs(1802) <= not(inputs(58));
    layer0_outputs(1803) <= not(inputs(168)) or (inputs(28));
    layer0_outputs(1804) <= (inputs(151)) and not (inputs(11));
    layer0_outputs(1805) <= not(inputs(248));
    layer0_outputs(1806) <= not((inputs(206)) xor (inputs(251)));
    layer0_outputs(1807) <= not(inputs(154));
    layer0_outputs(1808) <= inputs(196);
    layer0_outputs(1809) <= (inputs(29)) and (inputs(223));
    layer0_outputs(1810) <= not((inputs(43)) or (inputs(59)));
    layer0_outputs(1811) <= (inputs(232)) and not (inputs(99));
    layer0_outputs(1812) <= inputs(169);
    layer0_outputs(1813) <= (inputs(138)) or (inputs(151));
    layer0_outputs(1814) <= not(inputs(189)) or (inputs(125));
    layer0_outputs(1815) <= not(inputs(214)) or (inputs(248));
    layer0_outputs(1816) <= not((inputs(249)) and (inputs(11)));
    layer0_outputs(1817) <= not((inputs(165)) and (inputs(184)));
    layer0_outputs(1818) <= (inputs(194)) or (inputs(242));
    layer0_outputs(1819) <= not(inputs(221)) or (inputs(246));
    layer0_outputs(1820) <= inputs(116);
    layer0_outputs(1821) <= not(inputs(94)) or (inputs(150));
    layer0_outputs(1822) <= not(inputs(36));
    layer0_outputs(1823) <= (inputs(193)) or (inputs(0));
    layer0_outputs(1824) <= not(inputs(118));
    layer0_outputs(1825) <= not((inputs(87)) xor (inputs(122)));
    layer0_outputs(1826) <= (inputs(73)) and (inputs(152));
    layer0_outputs(1827) <= not((inputs(95)) or (inputs(193)));
    layer0_outputs(1828) <= inputs(29);
    layer0_outputs(1829) <= (inputs(116)) and not (inputs(141));
    layer0_outputs(1830) <= inputs(69);
    layer0_outputs(1831) <= not((inputs(250)) xor (inputs(69)));
    layer0_outputs(1832) <= not((inputs(217)) or (inputs(3)));
    layer0_outputs(1833) <= (inputs(58)) and (inputs(53));
    layer0_outputs(1834) <= not((inputs(62)) xor (inputs(218)));
    layer0_outputs(1835) <= not(inputs(168));
    layer0_outputs(1836) <= not((inputs(0)) xor (inputs(94)));
    layer0_outputs(1837) <= (inputs(78)) and not (inputs(221));
    layer0_outputs(1838) <= not((inputs(122)) and (inputs(154)));
    layer0_outputs(1839) <= not(inputs(153));
    layer0_outputs(1840) <= not(inputs(119)) or (inputs(129));
    layer0_outputs(1841) <= not((inputs(146)) or (inputs(43)));
    layer0_outputs(1842) <= not(inputs(89));
    layer0_outputs(1843) <= (inputs(181)) and not (inputs(97));
    layer0_outputs(1844) <= inputs(89);
    layer0_outputs(1845) <= inputs(232);
    layer0_outputs(1846) <= not((inputs(110)) or (inputs(122)));
    layer0_outputs(1847) <= inputs(208);
    layer0_outputs(1848) <= inputs(214);
    layer0_outputs(1849) <= inputs(67);
    layer0_outputs(1850) <= (inputs(163)) and not (inputs(176));
    layer0_outputs(1851) <= inputs(233);
    layer0_outputs(1852) <= (inputs(36)) or (inputs(105));
    layer0_outputs(1853) <= not((inputs(74)) or (inputs(159)));
    layer0_outputs(1854) <= (inputs(87)) xor (inputs(191));
    layer0_outputs(1855) <= (inputs(99)) or (inputs(145));
    layer0_outputs(1856) <= not((inputs(94)) xor (inputs(244)));
    layer0_outputs(1857) <= not(inputs(51)) or (inputs(96));
    layer0_outputs(1858) <= not(inputs(98));
    layer0_outputs(1859) <= not((inputs(187)) xor (inputs(13)));
    layer0_outputs(1860) <= inputs(115);
    layer0_outputs(1861) <= (inputs(52)) and not (inputs(76));
    layer0_outputs(1862) <= (inputs(132)) and not (inputs(143));
    layer0_outputs(1863) <= not((inputs(145)) or (inputs(246)));
    layer0_outputs(1864) <= not(inputs(79));
    layer0_outputs(1865) <= (inputs(179)) or (inputs(147));
    layer0_outputs(1866) <= (inputs(92)) and not (inputs(211));
    layer0_outputs(1867) <= not(inputs(250)) or (inputs(48));
    layer0_outputs(1868) <= inputs(120);
    layer0_outputs(1869) <= inputs(60);
    layer0_outputs(1870) <= (inputs(24)) and not (inputs(114));
    layer0_outputs(1871) <= not((inputs(202)) xor (inputs(111)));
    layer0_outputs(1872) <= not(inputs(200));
    layer0_outputs(1873) <= (inputs(116)) and not (inputs(90));
    layer0_outputs(1874) <= (inputs(145)) or (inputs(14));
    layer0_outputs(1875) <= not(inputs(41)) or (inputs(144));
    layer0_outputs(1876) <= not((inputs(204)) or (inputs(245)));
    layer0_outputs(1877) <= (inputs(71)) or (inputs(229));
    layer0_outputs(1878) <= (inputs(57)) xor (inputs(44));
    layer0_outputs(1879) <= inputs(239);
    layer0_outputs(1880) <= inputs(89);
    layer0_outputs(1881) <= not((inputs(222)) xor (inputs(106)));
    layer0_outputs(1882) <= (inputs(36)) and not (inputs(58));
    layer0_outputs(1883) <= '0';
    layer0_outputs(1884) <= not(inputs(184)) or (inputs(142));
    layer0_outputs(1885) <= not((inputs(130)) or (inputs(235)));
    layer0_outputs(1886) <= not((inputs(176)) and (inputs(83)));
    layer0_outputs(1887) <= not((inputs(144)) or (inputs(186)));
    layer0_outputs(1888) <= inputs(201);
    layer0_outputs(1889) <= inputs(210);
    layer0_outputs(1890) <= (inputs(116)) or (inputs(149));
    layer0_outputs(1891) <= inputs(120);
    layer0_outputs(1892) <= inputs(77);
    layer0_outputs(1893) <= not(inputs(78)) or (inputs(112));
    layer0_outputs(1894) <= not((inputs(135)) or (inputs(207)));
    layer0_outputs(1895) <= not((inputs(201)) or (inputs(70)));
    layer0_outputs(1896) <= (inputs(3)) xor (inputs(51));
    layer0_outputs(1897) <= not((inputs(220)) or (inputs(13)));
    layer0_outputs(1898) <= inputs(197);
    layer0_outputs(1899) <= (inputs(59)) and not (inputs(250));
    layer0_outputs(1900) <= (inputs(114)) xor (inputs(101));
    layer0_outputs(1901) <= inputs(229);
    layer0_outputs(1902) <= (inputs(173)) or (inputs(54));
    layer0_outputs(1903) <= not(inputs(136)) or (inputs(213));
    layer0_outputs(1904) <= not((inputs(142)) xor (inputs(121)));
    layer0_outputs(1905) <= not(inputs(219));
    layer0_outputs(1906) <= not(inputs(180)) or (inputs(63));
    layer0_outputs(1907) <= not((inputs(37)) or (inputs(239)));
    layer0_outputs(1908) <= not((inputs(4)) or (inputs(142)));
    layer0_outputs(1909) <= not((inputs(26)) or (inputs(76)));
    layer0_outputs(1910) <= '1';
    layer0_outputs(1911) <= (inputs(169)) xor (inputs(253));
    layer0_outputs(1912) <= (inputs(121)) and not (inputs(233));
    layer0_outputs(1913) <= not((inputs(108)) or (inputs(152)));
    layer0_outputs(1914) <= not(inputs(193));
    layer0_outputs(1915) <= not((inputs(132)) or (inputs(196)));
    layer0_outputs(1916) <= inputs(188);
    layer0_outputs(1917) <= (inputs(86)) or (inputs(114));
    layer0_outputs(1918) <= (inputs(204)) and not (inputs(65));
    layer0_outputs(1919) <= inputs(41);
    layer0_outputs(1920) <= inputs(209);
    layer0_outputs(1921) <= not((inputs(148)) or (inputs(174)));
    layer0_outputs(1922) <= (inputs(84)) or (inputs(68));
    layer0_outputs(1923) <= (inputs(89)) or (inputs(66));
    layer0_outputs(1924) <= not((inputs(106)) xor (inputs(0)));
    layer0_outputs(1925) <= (inputs(43)) and not (inputs(54));
    layer0_outputs(1926) <= not((inputs(251)) xor (inputs(36)));
    layer0_outputs(1927) <= inputs(180);
    layer0_outputs(1928) <= (inputs(7)) and not (inputs(191));
    layer0_outputs(1929) <= not(inputs(221));
    layer0_outputs(1930) <= (inputs(250)) xor (inputs(29));
    layer0_outputs(1931) <= (inputs(27)) xor (inputs(74));
    layer0_outputs(1932) <= (inputs(132)) or (inputs(138));
    layer0_outputs(1933) <= not(inputs(140)) or (inputs(21));
    layer0_outputs(1934) <= (inputs(186)) and not (inputs(16));
    layer0_outputs(1935) <= not((inputs(146)) or (inputs(108)));
    layer0_outputs(1936) <= not((inputs(116)) and (inputs(73)));
    layer0_outputs(1937) <= not((inputs(135)) xor (inputs(104)));
    layer0_outputs(1938) <= inputs(150);
    layer0_outputs(1939) <= not(inputs(124));
    layer0_outputs(1940) <= inputs(148);
    layer0_outputs(1941) <= (inputs(128)) xor (inputs(135));
    layer0_outputs(1942) <= not((inputs(137)) and (inputs(188)));
    layer0_outputs(1943) <= not(inputs(36)) or (inputs(173));
    layer0_outputs(1944) <= not((inputs(146)) or (inputs(63)));
    layer0_outputs(1945) <= not((inputs(237)) or (inputs(20)));
    layer0_outputs(1946) <= (inputs(131)) or (inputs(68));
    layer0_outputs(1947) <= (inputs(130)) or (inputs(127));
    layer0_outputs(1948) <= not((inputs(200)) or (inputs(240)));
    layer0_outputs(1949) <= not(inputs(238));
    layer0_outputs(1950) <= not((inputs(21)) or (inputs(185)));
    layer0_outputs(1951) <= not(inputs(65));
    layer0_outputs(1952) <= (inputs(86)) or (inputs(170));
    layer0_outputs(1953) <= (inputs(118)) and (inputs(177));
    layer0_outputs(1954) <= (inputs(86)) or (inputs(221));
    layer0_outputs(1955) <= not((inputs(177)) or (inputs(134)));
    layer0_outputs(1956) <= not((inputs(246)) xor (inputs(59)));
    layer0_outputs(1957) <= (inputs(83)) and not (inputs(191));
    layer0_outputs(1958) <= '1';
    layer0_outputs(1959) <= not((inputs(138)) or (inputs(58)));
    layer0_outputs(1960) <= inputs(39);
    layer0_outputs(1961) <= inputs(233);
    layer0_outputs(1962) <= inputs(19);
    layer0_outputs(1963) <= inputs(3);
    layer0_outputs(1964) <= (inputs(157)) and not (inputs(2));
    layer0_outputs(1965) <= (inputs(86)) or (inputs(108));
    layer0_outputs(1966) <= not(inputs(168)) or (inputs(116));
    layer0_outputs(1967) <= not(inputs(74)) or (inputs(183));
    layer0_outputs(1968) <= not(inputs(90));
    layer0_outputs(1969) <= (inputs(183)) xor (inputs(239));
    layer0_outputs(1970) <= not(inputs(9));
    layer0_outputs(1971) <= (inputs(68)) and (inputs(100));
    layer0_outputs(1972) <= not((inputs(106)) and (inputs(169)));
    layer0_outputs(1973) <= inputs(213);
    layer0_outputs(1974) <= not(inputs(125)) or (inputs(205));
    layer0_outputs(1975) <= inputs(228);
    layer0_outputs(1976) <= not(inputs(226));
    layer0_outputs(1977) <= not((inputs(168)) xor (inputs(133)));
    layer0_outputs(1978) <= (inputs(139)) or (inputs(205));
    layer0_outputs(1979) <= not((inputs(184)) or (inputs(56)));
    layer0_outputs(1980) <= (inputs(242)) and not (inputs(30));
    layer0_outputs(1981) <= '0';
    layer0_outputs(1982) <= inputs(72);
    layer0_outputs(1983) <= inputs(94);
    layer0_outputs(1984) <= (inputs(186)) xor (inputs(82));
    layer0_outputs(1985) <= (inputs(109)) and not (inputs(112));
    layer0_outputs(1986) <= inputs(14);
    layer0_outputs(1987) <= not(inputs(232));
    layer0_outputs(1988) <= (inputs(97)) or (inputs(96));
    layer0_outputs(1989) <= not((inputs(165)) or (inputs(205)));
    layer0_outputs(1990) <= not((inputs(131)) or (inputs(34)));
    layer0_outputs(1991) <= not((inputs(14)) or (inputs(235)));
    layer0_outputs(1992) <= (inputs(211)) xor (inputs(226));
    layer0_outputs(1993) <= (inputs(62)) xor (inputs(53));
    layer0_outputs(1994) <= not((inputs(76)) or (inputs(93)));
    layer0_outputs(1995) <= not((inputs(85)) or (inputs(102)));
    layer0_outputs(1996) <= inputs(168);
    layer0_outputs(1997) <= inputs(210);
    layer0_outputs(1998) <= (inputs(74)) xor (inputs(59));
    layer0_outputs(1999) <= inputs(118);
    layer0_outputs(2000) <= inputs(113);
    layer0_outputs(2001) <= inputs(193);
    layer0_outputs(2002) <= inputs(122);
    layer0_outputs(2003) <= '1';
    layer0_outputs(2004) <= (inputs(153)) xor (inputs(116));
    layer0_outputs(2005) <= '1';
    layer0_outputs(2006) <= '1';
    layer0_outputs(2007) <= not(inputs(57));
    layer0_outputs(2008) <= not((inputs(164)) or (inputs(165)));
    layer0_outputs(2009) <= not((inputs(167)) or (inputs(31)));
    layer0_outputs(2010) <= not((inputs(146)) and (inputs(251)));
    layer0_outputs(2011) <= (inputs(244)) and not (inputs(143));
    layer0_outputs(2012) <= (inputs(122)) xor (inputs(212));
    layer0_outputs(2013) <= not(inputs(113));
    layer0_outputs(2014) <= (inputs(47)) or (inputs(189));
    layer0_outputs(2015) <= not((inputs(62)) or (inputs(137)));
    layer0_outputs(2016) <= (inputs(197)) and not (inputs(27));
    layer0_outputs(2017) <= (inputs(21)) xor (inputs(189));
    layer0_outputs(2018) <= not(inputs(228)) or (inputs(254));
    layer0_outputs(2019) <= not(inputs(230));
    layer0_outputs(2020) <= (inputs(238)) xor (inputs(191));
    layer0_outputs(2021) <= not(inputs(235));
    layer0_outputs(2022) <= not((inputs(254)) or (inputs(242)));
    layer0_outputs(2023) <= not((inputs(12)) or (inputs(144)));
    layer0_outputs(2024) <= (inputs(71)) and not (inputs(125));
    layer0_outputs(2025) <= (inputs(174)) or (inputs(54));
    layer0_outputs(2026) <= inputs(77);
    layer0_outputs(2027) <= (inputs(153)) and not (inputs(212));
    layer0_outputs(2028) <= not(inputs(164));
    layer0_outputs(2029) <= not(inputs(24));
    layer0_outputs(2030) <= (inputs(247)) xor (inputs(240));
    layer0_outputs(2031) <= not(inputs(99)) or (inputs(248));
    layer0_outputs(2032) <= not(inputs(142));
    layer0_outputs(2033) <= not(inputs(23)) or (inputs(236));
    layer0_outputs(2034) <= not((inputs(70)) or (inputs(153)));
    layer0_outputs(2035) <= (inputs(189)) xor (inputs(4));
    layer0_outputs(2036) <= not(inputs(44)) or (inputs(218));
    layer0_outputs(2037) <= inputs(135);
    layer0_outputs(2038) <= (inputs(22)) or (inputs(33));
    layer0_outputs(2039) <= (inputs(62)) or (inputs(51));
    layer0_outputs(2040) <= (inputs(230)) and not (inputs(4));
    layer0_outputs(2041) <= not(inputs(136));
    layer0_outputs(2042) <= not(inputs(123));
    layer0_outputs(2043) <= not(inputs(131));
    layer0_outputs(2044) <= not(inputs(172)) or (inputs(36));
    layer0_outputs(2045) <= inputs(77);
    layer0_outputs(2046) <= not(inputs(187)) or (inputs(58));
    layer0_outputs(2047) <= not(inputs(63)) or (inputs(251));
    layer0_outputs(2048) <= not((inputs(195)) xor (inputs(157)));
    layer0_outputs(2049) <= not((inputs(155)) xor (inputs(94)));
    layer0_outputs(2050) <= (inputs(190)) or (inputs(180));
    layer0_outputs(2051) <= (inputs(121)) and not (inputs(38));
    layer0_outputs(2052) <= not(inputs(60));
    layer0_outputs(2053) <= (inputs(159)) or (inputs(105));
    layer0_outputs(2054) <= not(inputs(101)) or (inputs(191));
    layer0_outputs(2055) <= (inputs(132)) or (inputs(148));
    layer0_outputs(2056) <= (inputs(27)) and not (inputs(193));
    layer0_outputs(2057) <= not(inputs(9)) or (inputs(248));
    layer0_outputs(2058) <= not((inputs(4)) or (inputs(187)));
    layer0_outputs(2059) <= inputs(121);
    layer0_outputs(2060) <= inputs(51);
    layer0_outputs(2061) <= inputs(92);
    layer0_outputs(2062) <= (inputs(165)) and (inputs(246));
    layer0_outputs(2063) <= (inputs(229)) xor (inputs(252));
    layer0_outputs(2064) <= inputs(158);
    layer0_outputs(2065) <= not((inputs(186)) xor (inputs(185)));
    layer0_outputs(2066) <= not(inputs(127));
    layer0_outputs(2067) <= not(inputs(227));
    layer0_outputs(2068) <= (inputs(48)) xor (inputs(119));
    layer0_outputs(2069) <= not((inputs(128)) xor (inputs(118)));
    layer0_outputs(2070) <= not((inputs(35)) or (inputs(239)));
    layer0_outputs(2071) <= '0';
    layer0_outputs(2072) <= not(inputs(28));
    layer0_outputs(2073) <= (inputs(23)) and not (inputs(130));
    layer0_outputs(2074) <= not((inputs(171)) or (inputs(227)));
    layer0_outputs(2075) <= (inputs(200)) and not (inputs(243));
    layer0_outputs(2076) <= not((inputs(207)) xor (inputs(212)));
    layer0_outputs(2077) <= (inputs(103)) and not (inputs(201));
    layer0_outputs(2078) <= not(inputs(18));
    layer0_outputs(2079) <= (inputs(131)) or (inputs(158));
    layer0_outputs(2080) <= inputs(179);
    layer0_outputs(2081) <= not(inputs(247));
    layer0_outputs(2082) <= inputs(154);
    layer0_outputs(2083) <= inputs(7);
    layer0_outputs(2084) <= (inputs(104)) or (inputs(46));
    layer0_outputs(2085) <= not(inputs(200)) or (inputs(30));
    layer0_outputs(2086) <= not(inputs(178));
    layer0_outputs(2087) <= not(inputs(198)) or (inputs(77));
    layer0_outputs(2088) <= (inputs(125)) and not (inputs(119));
    layer0_outputs(2089) <= not((inputs(51)) or (inputs(118)));
    layer0_outputs(2090) <= not(inputs(103)) or (inputs(164));
    layer0_outputs(2091) <= inputs(99);
    layer0_outputs(2092) <= (inputs(181)) or (inputs(151));
    layer0_outputs(2093) <= not((inputs(195)) xor (inputs(187)));
    layer0_outputs(2094) <= not(inputs(62));
    layer0_outputs(2095) <= not((inputs(52)) or (inputs(129)));
    layer0_outputs(2096) <= inputs(89);
    layer0_outputs(2097) <= not(inputs(149));
    layer0_outputs(2098) <= not(inputs(196)) or (inputs(240));
    layer0_outputs(2099) <= inputs(132);
    layer0_outputs(2100) <= inputs(14);
    layer0_outputs(2101) <= not(inputs(39));
    layer0_outputs(2102) <= inputs(99);
    layer0_outputs(2103) <= (inputs(214)) and (inputs(119));
    layer0_outputs(2104) <= not(inputs(173));
    layer0_outputs(2105) <= not(inputs(83));
    layer0_outputs(2106) <= not(inputs(62)) or (inputs(239));
    layer0_outputs(2107) <= (inputs(26)) and not (inputs(141));
    layer0_outputs(2108) <= not(inputs(227));
    layer0_outputs(2109) <= inputs(119);
    layer0_outputs(2110) <= not(inputs(70));
    layer0_outputs(2111) <= inputs(44);
    layer0_outputs(2112) <= (inputs(250)) or (inputs(111));
    layer0_outputs(2113) <= inputs(74);
    layer0_outputs(2114) <= not((inputs(127)) or (inputs(200)));
    layer0_outputs(2115) <= inputs(167);
    layer0_outputs(2116) <= not((inputs(222)) or (inputs(103)));
    layer0_outputs(2117) <= inputs(249);
    layer0_outputs(2118) <= inputs(20);
    layer0_outputs(2119) <= not((inputs(186)) or (inputs(6)));
    layer0_outputs(2120) <= not(inputs(180)) or (inputs(97));
    layer0_outputs(2121) <= (inputs(56)) or (inputs(248));
    layer0_outputs(2122) <= inputs(3);
    layer0_outputs(2123) <= not((inputs(139)) and (inputs(20)));
    layer0_outputs(2124) <= not(inputs(115));
    layer0_outputs(2125) <= '0';
    layer0_outputs(2126) <= not(inputs(56)) or (inputs(175));
    layer0_outputs(2127) <= (inputs(92)) and not (inputs(162));
    layer0_outputs(2128) <= (inputs(135)) and not (inputs(160));
    layer0_outputs(2129) <= inputs(181);
    layer0_outputs(2130) <= (inputs(237)) or (inputs(99));
    layer0_outputs(2131) <= (inputs(29)) and not (inputs(254));
    layer0_outputs(2132) <= (inputs(44)) and not (inputs(133));
    layer0_outputs(2133) <= not((inputs(91)) or (inputs(186)));
    layer0_outputs(2134) <= '0';
    layer0_outputs(2135) <= not(inputs(197));
    layer0_outputs(2136) <= not(inputs(197));
    layer0_outputs(2137) <= (inputs(90)) and not (inputs(174));
    layer0_outputs(2138) <= not(inputs(215));
    layer0_outputs(2139) <= inputs(96);
    layer0_outputs(2140) <= (inputs(35)) or (inputs(139));
    layer0_outputs(2141) <= (inputs(49)) xor (inputs(79));
    layer0_outputs(2142) <= (inputs(239)) or (inputs(185));
    layer0_outputs(2143) <= (inputs(115)) or (inputs(164));
    layer0_outputs(2144) <= inputs(87);
    layer0_outputs(2145) <= inputs(7);
    layer0_outputs(2146) <= inputs(153);
    layer0_outputs(2147) <= (inputs(210)) or (inputs(243));
    layer0_outputs(2148) <= (inputs(237)) or (inputs(235));
    layer0_outputs(2149) <= not((inputs(220)) and (inputs(249)));
    layer0_outputs(2150) <= (inputs(155)) xor (inputs(235));
    layer0_outputs(2151) <= '0';
    layer0_outputs(2152) <= (inputs(142)) or (inputs(171));
    layer0_outputs(2153) <= inputs(195);
    layer0_outputs(2154) <= inputs(214);
    layer0_outputs(2155) <= (inputs(139)) and not (inputs(137));
    layer0_outputs(2156) <= not(inputs(227));
    layer0_outputs(2157) <= not((inputs(39)) or (inputs(2)));
    layer0_outputs(2158) <= (inputs(81)) or (inputs(209));
    layer0_outputs(2159) <= inputs(231);
    layer0_outputs(2160) <= inputs(157);
    layer0_outputs(2161) <= not(inputs(107)) or (inputs(47));
    layer0_outputs(2162) <= not(inputs(82));
    layer0_outputs(2163) <= (inputs(197)) or (inputs(211));
    layer0_outputs(2164) <= not(inputs(103));
    layer0_outputs(2165) <= not(inputs(35)) or (inputs(174));
    layer0_outputs(2166) <= inputs(83);
    layer0_outputs(2167) <= (inputs(32)) or (inputs(8));
    layer0_outputs(2168) <= (inputs(218)) or (inputs(236));
    layer0_outputs(2169) <= not(inputs(218));
    layer0_outputs(2170) <= not(inputs(202)) or (inputs(125));
    layer0_outputs(2171) <= (inputs(249)) and not (inputs(127));
    layer0_outputs(2172) <= (inputs(80)) xor (inputs(131));
    layer0_outputs(2173) <= inputs(240);
    layer0_outputs(2174) <= inputs(110);
    layer0_outputs(2175) <= not(inputs(104));
    layer0_outputs(2176) <= (inputs(42)) or (inputs(189));
    layer0_outputs(2177) <= not(inputs(217));
    layer0_outputs(2178) <= not(inputs(130)) or (inputs(48));
    layer0_outputs(2179) <= not((inputs(149)) or (inputs(141)));
    layer0_outputs(2180) <= inputs(93);
    layer0_outputs(2181) <= not(inputs(253)) or (inputs(249));
    layer0_outputs(2182) <= inputs(103);
    layer0_outputs(2183) <= not(inputs(42));
    layer0_outputs(2184) <= not((inputs(81)) or (inputs(203)));
    layer0_outputs(2185) <= not((inputs(208)) or (inputs(35)));
    layer0_outputs(2186) <= (inputs(106)) xor (inputs(93));
    layer0_outputs(2187) <= (inputs(76)) or (inputs(222));
    layer0_outputs(2188) <= not(inputs(23));
    layer0_outputs(2189) <= inputs(227);
    layer0_outputs(2190) <= (inputs(51)) and not (inputs(226));
    layer0_outputs(2191) <= (inputs(87)) or (inputs(222));
    layer0_outputs(2192) <= not(inputs(94));
    layer0_outputs(2193) <= (inputs(54)) or (inputs(249));
    layer0_outputs(2194) <= not(inputs(103));
    layer0_outputs(2195) <= inputs(231);
    layer0_outputs(2196) <= not((inputs(180)) or (inputs(161)));
    layer0_outputs(2197) <= not(inputs(188));
    layer0_outputs(2198) <= not((inputs(76)) or (inputs(75)));
    layer0_outputs(2199) <= inputs(76);
    layer0_outputs(2200) <= inputs(114);
    layer0_outputs(2201) <= not((inputs(209)) or (inputs(244)));
    layer0_outputs(2202) <= (inputs(9)) xor (inputs(174));
    layer0_outputs(2203) <= not(inputs(117));
    layer0_outputs(2204) <= inputs(158);
    layer0_outputs(2205) <= inputs(56);
    layer0_outputs(2206) <= inputs(90);
    layer0_outputs(2207) <= not(inputs(187));
    layer0_outputs(2208) <= inputs(160);
    layer0_outputs(2209) <= inputs(42);
    layer0_outputs(2210) <= (inputs(207)) xor (inputs(25));
    layer0_outputs(2211) <= not((inputs(30)) or (inputs(10)));
    layer0_outputs(2212) <= not((inputs(139)) and (inputs(170)));
    layer0_outputs(2213) <= not(inputs(150)) or (inputs(37));
    layer0_outputs(2214) <= not(inputs(9));
    layer0_outputs(2215) <= inputs(219);
    layer0_outputs(2216) <= not(inputs(122));
    layer0_outputs(2217) <= (inputs(251)) or (inputs(57));
    layer0_outputs(2218) <= inputs(22);
    layer0_outputs(2219) <= (inputs(124)) or (inputs(75));
    layer0_outputs(2220) <= (inputs(43)) and not (inputs(157));
    layer0_outputs(2221) <= not((inputs(110)) or (inputs(107)));
    layer0_outputs(2222) <= (inputs(75)) or (inputs(115));
    layer0_outputs(2223) <= not((inputs(163)) or (inputs(210)));
    layer0_outputs(2224) <= not((inputs(17)) or (inputs(93)));
    layer0_outputs(2225) <= (inputs(4)) xor (inputs(124));
    layer0_outputs(2226) <= (inputs(9)) and not (inputs(214));
    layer0_outputs(2227) <= '1';
    layer0_outputs(2228) <= not(inputs(159));
    layer0_outputs(2229) <= inputs(24);
    layer0_outputs(2230) <= not(inputs(181));
    layer0_outputs(2231) <= (inputs(72)) xor (inputs(185));
    layer0_outputs(2232) <= not(inputs(233));
    layer0_outputs(2233) <= inputs(133);
    layer0_outputs(2234) <= (inputs(46)) or (inputs(99));
    layer0_outputs(2235) <= inputs(38);
    layer0_outputs(2236) <= inputs(15);
    layer0_outputs(2237) <= not(inputs(172));
    layer0_outputs(2238) <= not(inputs(14));
    layer0_outputs(2239) <= inputs(66);
    layer0_outputs(2240) <= (inputs(235)) or (inputs(218));
    layer0_outputs(2241) <= not(inputs(68)) or (inputs(244));
    layer0_outputs(2242) <= not(inputs(26));
    layer0_outputs(2243) <= not((inputs(72)) or (inputs(247)));
    layer0_outputs(2244) <= not((inputs(94)) or (inputs(59)));
    layer0_outputs(2245) <= inputs(212);
    layer0_outputs(2246) <= (inputs(241)) or (inputs(147));
    layer0_outputs(2247) <= (inputs(87)) or (inputs(120));
    layer0_outputs(2248) <= not(inputs(131)) or (inputs(254));
    layer0_outputs(2249) <= (inputs(231)) and not (inputs(46));
    layer0_outputs(2250) <= not(inputs(178)) or (inputs(237));
    layer0_outputs(2251) <= not((inputs(35)) or (inputs(159)));
    layer0_outputs(2252) <= not(inputs(44)) or (inputs(206));
    layer0_outputs(2253) <= inputs(4);
    layer0_outputs(2254) <= inputs(100);
    layer0_outputs(2255) <= not(inputs(108)) or (inputs(175));
    layer0_outputs(2256) <= not(inputs(193));
    layer0_outputs(2257) <= not((inputs(16)) or (inputs(24)));
    layer0_outputs(2258) <= inputs(213);
    layer0_outputs(2259) <= not(inputs(146));
    layer0_outputs(2260) <= inputs(86);
    layer0_outputs(2261) <= (inputs(168)) and not (inputs(132));
    layer0_outputs(2262) <= (inputs(24)) and not (inputs(4));
    layer0_outputs(2263) <= (inputs(195)) or (inputs(248));
    layer0_outputs(2264) <= inputs(191);
    layer0_outputs(2265) <= inputs(164);
    layer0_outputs(2266) <= (inputs(13)) or (inputs(11));
    layer0_outputs(2267) <= not(inputs(219));
    layer0_outputs(2268) <= inputs(27);
    layer0_outputs(2269) <= inputs(185);
    layer0_outputs(2270) <= not(inputs(73));
    layer0_outputs(2271) <= (inputs(61)) xor (inputs(24));
    layer0_outputs(2272) <= not(inputs(92));
    layer0_outputs(2273) <= inputs(166);
    layer0_outputs(2274) <= '1';
    layer0_outputs(2275) <= inputs(66);
    layer0_outputs(2276) <= (inputs(189)) or (inputs(34));
    layer0_outputs(2277) <= not(inputs(198));
    layer0_outputs(2278) <= (inputs(32)) and not (inputs(81));
    layer0_outputs(2279) <= inputs(129);
    layer0_outputs(2280) <= (inputs(119)) or (inputs(30));
    layer0_outputs(2281) <= '0';
    layer0_outputs(2282) <= not(inputs(24)) or (inputs(144));
    layer0_outputs(2283) <= inputs(253);
    layer0_outputs(2284) <= not((inputs(255)) and (inputs(18)));
    layer0_outputs(2285) <= inputs(247);
    layer0_outputs(2286) <= '0';
    layer0_outputs(2287) <= not(inputs(167));
    layer0_outputs(2288) <= not((inputs(173)) xor (inputs(71)));
    layer0_outputs(2289) <= not(inputs(110)) or (inputs(94));
    layer0_outputs(2290) <= not((inputs(32)) or (inputs(63)));
    layer0_outputs(2291) <= not((inputs(168)) or (inputs(13)));
    layer0_outputs(2292) <= not((inputs(202)) and (inputs(1)));
    layer0_outputs(2293) <= (inputs(132)) or (inputs(157));
    layer0_outputs(2294) <= not(inputs(241));
    layer0_outputs(2295) <= inputs(185);
    layer0_outputs(2296) <= (inputs(124)) and not (inputs(194));
    layer0_outputs(2297) <= '1';
    layer0_outputs(2298) <= not(inputs(195)) or (inputs(2));
    layer0_outputs(2299) <= not(inputs(202)) or (inputs(44));
    layer0_outputs(2300) <= not(inputs(89)) or (inputs(73));
    layer0_outputs(2301) <= not(inputs(180));
    layer0_outputs(2302) <= (inputs(120)) and not (inputs(123));
    layer0_outputs(2303) <= not(inputs(37)) or (inputs(130));
    layer0_outputs(2304) <= not(inputs(99));
    layer0_outputs(2305) <= inputs(71);
    layer0_outputs(2306) <= not((inputs(121)) xor (inputs(190)));
    layer0_outputs(2307) <= inputs(178);
    layer0_outputs(2308) <= inputs(80);
    layer0_outputs(2309) <= not(inputs(170)) or (inputs(95));
    layer0_outputs(2310) <= not(inputs(152)) or (inputs(18));
    layer0_outputs(2311) <= not(inputs(202));
    layer0_outputs(2312) <= (inputs(29)) and not (inputs(130));
    layer0_outputs(2313) <= (inputs(25)) or (inputs(147));
    layer0_outputs(2314) <= (inputs(123)) xor (inputs(104));
    layer0_outputs(2315) <= (inputs(26)) and not (inputs(17));
    layer0_outputs(2316) <= not(inputs(127));
    layer0_outputs(2317) <= (inputs(28)) and not (inputs(227));
    layer0_outputs(2318) <= not((inputs(214)) or (inputs(129)));
    layer0_outputs(2319) <= not((inputs(66)) or (inputs(39)));
    layer0_outputs(2320) <= not((inputs(243)) or (inputs(51)));
    layer0_outputs(2321) <= not(inputs(232)) or (inputs(48));
    layer0_outputs(2322) <= not((inputs(67)) and (inputs(215)));
    layer0_outputs(2323) <= inputs(71);
    layer0_outputs(2324) <= not(inputs(167)) or (inputs(65));
    layer0_outputs(2325) <= inputs(208);
    layer0_outputs(2326) <= (inputs(103)) or (inputs(10));
    layer0_outputs(2327) <= not((inputs(55)) xor (inputs(72)));
    layer0_outputs(2328) <= (inputs(10)) or (inputs(127));
    layer0_outputs(2329) <= not(inputs(184));
    layer0_outputs(2330) <= not((inputs(209)) xor (inputs(215)));
    layer0_outputs(2331) <= not(inputs(143));
    layer0_outputs(2332) <= (inputs(149)) or (inputs(70));
    layer0_outputs(2333) <= inputs(58);
    layer0_outputs(2334) <= (inputs(248)) or (inputs(237));
    layer0_outputs(2335) <= not((inputs(176)) xor (inputs(198)));
    layer0_outputs(2336) <= not((inputs(3)) xor (inputs(138)));
    layer0_outputs(2337) <= not(inputs(35)) or (inputs(189));
    layer0_outputs(2338) <= (inputs(218)) and not (inputs(140));
    layer0_outputs(2339) <= not((inputs(120)) and (inputs(135)));
    layer0_outputs(2340) <= (inputs(199)) and not (inputs(60));
    layer0_outputs(2341) <= (inputs(184)) and not (inputs(57));
    layer0_outputs(2342) <= (inputs(183)) and (inputs(238));
    layer0_outputs(2343) <= '0';
    layer0_outputs(2344) <= not(inputs(44)) or (inputs(136));
    layer0_outputs(2345) <= not(inputs(2));
    layer0_outputs(2346) <= (inputs(232)) xor (inputs(40));
    layer0_outputs(2347) <= not((inputs(193)) xor (inputs(173)));
    layer0_outputs(2348) <= (inputs(161)) xor (inputs(135));
    layer0_outputs(2349) <= not(inputs(77)) or (inputs(242));
    layer0_outputs(2350) <= inputs(230);
    layer0_outputs(2351) <= not((inputs(102)) or (inputs(94)));
    layer0_outputs(2352) <= not(inputs(171)) or (inputs(48));
    layer0_outputs(2353) <= (inputs(42)) or (inputs(26));
    layer0_outputs(2354) <= (inputs(124)) and not (inputs(165));
    layer0_outputs(2355) <= not((inputs(180)) xor (inputs(210)));
    layer0_outputs(2356) <= not(inputs(126));
    layer0_outputs(2357) <= not((inputs(216)) or (inputs(131)));
    layer0_outputs(2358) <= inputs(25);
    layer0_outputs(2359) <= (inputs(180)) and not (inputs(140));
    layer0_outputs(2360) <= not(inputs(230));
    layer0_outputs(2361) <= not(inputs(245));
    layer0_outputs(2362) <= not((inputs(78)) or (inputs(133)));
    layer0_outputs(2363) <= not((inputs(175)) and (inputs(13)));
    layer0_outputs(2364) <= not(inputs(221));
    layer0_outputs(2365) <= inputs(95);
    layer0_outputs(2366) <= not(inputs(177));
    layer0_outputs(2367) <= (inputs(255)) or (inputs(7));
    layer0_outputs(2368) <= not(inputs(238));
    layer0_outputs(2369) <= inputs(39);
    layer0_outputs(2370) <= inputs(159);
    layer0_outputs(2371) <= (inputs(42)) and not (inputs(252));
    layer0_outputs(2372) <= (inputs(20)) or (inputs(121));
    layer0_outputs(2373) <= (inputs(165)) or (inputs(200));
    layer0_outputs(2374) <= not(inputs(35));
    layer0_outputs(2375) <= (inputs(190)) or (inputs(5));
    layer0_outputs(2376) <= not(inputs(196)) or (inputs(33));
    layer0_outputs(2377) <= inputs(104);
    layer0_outputs(2378) <= not(inputs(76));
    layer0_outputs(2379) <= (inputs(242)) or (inputs(34));
    layer0_outputs(2380) <= '1';
    layer0_outputs(2381) <= not(inputs(83));
    layer0_outputs(2382) <= not((inputs(83)) and (inputs(16)));
    layer0_outputs(2383) <= not(inputs(120));
    layer0_outputs(2384) <= not((inputs(228)) or (inputs(146)));
    layer0_outputs(2385) <= (inputs(100)) xor (inputs(188));
    layer0_outputs(2386) <= inputs(55);
    layer0_outputs(2387) <= inputs(77);
    layer0_outputs(2388) <= inputs(123);
    layer0_outputs(2389) <= '1';
    layer0_outputs(2390) <= (inputs(250)) xor (inputs(218));
    layer0_outputs(2391) <= not((inputs(203)) or (inputs(84)));
    layer0_outputs(2392) <= inputs(63);
    layer0_outputs(2393) <= (inputs(43)) xor (inputs(238));
    layer0_outputs(2394) <= inputs(20);
    layer0_outputs(2395) <= (inputs(250)) or (inputs(66));
    layer0_outputs(2396) <= not((inputs(141)) or (inputs(144)));
    layer0_outputs(2397) <= (inputs(122)) and not (inputs(101));
    layer0_outputs(2398) <= (inputs(180)) xor (inputs(45));
    layer0_outputs(2399) <= not(inputs(135)) or (inputs(205));
    layer0_outputs(2400) <= not(inputs(215)) or (inputs(205));
    layer0_outputs(2401) <= inputs(193);
    layer0_outputs(2402) <= (inputs(86)) xor (inputs(125));
    layer0_outputs(2403) <= (inputs(24)) or (inputs(93));
    layer0_outputs(2404) <= (inputs(107)) or (inputs(101));
    layer0_outputs(2405) <= (inputs(202)) or (inputs(146));
    layer0_outputs(2406) <= not((inputs(24)) or (inputs(161)));
    layer0_outputs(2407) <= '0';
    layer0_outputs(2408) <= not((inputs(104)) xor (inputs(149)));
    layer0_outputs(2409) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(2410) <= (inputs(190)) and not (inputs(49));
    layer0_outputs(2411) <= (inputs(152)) and not (inputs(39));
    layer0_outputs(2412) <= not(inputs(227));
    layer0_outputs(2413) <= not((inputs(160)) xor (inputs(189)));
    layer0_outputs(2414) <= not(inputs(67));
    layer0_outputs(2415) <= (inputs(167)) and not (inputs(38));
    layer0_outputs(2416) <= (inputs(71)) and not (inputs(57));
    layer0_outputs(2417) <= inputs(229);
    layer0_outputs(2418) <= inputs(130);
    layer0_outputs(2419) <= (inputs(47)) xor (inputs(79));
    layer0_outputs(2420) <= not(inputs(149));
    layer0_outputs(2421) <= (inputs(107)) or (inputs(108));
    layer0_outputs(2422) <= not((inputs(109)) xor (inputs(196)));
    layer0_outputs(2423) <= inputs(146);
    layer0_outputs(2424) <= inputs(120);
    layer0_outputs(2425) <= (inputs(240)) and not (inputs(72));
    layer0_outputs(2426) <= not((inputs(91)) or (inputs(31)));
    layer0_outputs(2427) <= not((inputs(66)) or (inputs(247)));
    layer0_outputs(2428) <= not(inputs(69)) or (inputs(225));
    layer0_outputs(2429) <= (inputs(77)) xor (inputs(173));
    layer0_outputs(2430) <= not((inputs(55)) and (inputs(200)));
    layer0_outputs(2431) <= not(inputs(119));
    layer0_outputs(2432) <= inputs(150);
    layer0_outputs(2433) <= '0';
    layer0_outputs(2434) <= not(inputs(188)) or (inputs(255));
    layer0_outputs(2435) <= not(inputs(205)) or (inputs(248));
    layer0_outputs(2436) <= (inputs(231)) and (inputs(49));
    layer0_outputs(2437) <= not((inputs(121)) or (inputs(126)));
    layer0_outputs(2438) <= not((inputs(213)) or (inputs(253)));
    layer0_outputs(2439) <= (inputs(118)) and not (inputs(6));
    layer0_outputs(2440) <= not((inputs(243)) xor (inputs(234)));
    layer0_outputs(2441) <= not(inputs(156));
    layer0_outputs(2442) <= (inputs(45)) or (inputs(69));
    layer0_outputs(2443) <= (inputs(141)) or (inputs(194));
    layer0_outputs(2444) <= (inputs(78)) or (inputs(116));
    layer0_outputs(2445) <= inputs(253);
    layer0_outputs(2446) <= inputs(189);
    layer0_outputs(2447) <= not((inputs(247)) xor (inputs(219)));
    layer0_outputs(2448) <= inputs(53);
    layer0_outputs(2449) <= (inputs(204)) or (inputs(123));
    layer0_outputs(2450) <= not(inputs(36)) or (inputs(219));
    layer0_outputs(2451) <= inputs(97);
    layer0_outputs(2452) <= not(inputs(83));
    layer0_outputs(2453) <= not(inputs(42));
    layer0_outputs(2454) <= not(inputs(174)) or (inputs(16));
    layer0_outputs(2455) <= (inputs(244)) or (inputs(163));
    layer0_outputs(2456) <= (inputs(54)) and not (inputs(15));
    layer0_outputs(2457) <= (inputs(1)) xor (inputs(8));
    layer0_outputs(2458) <= not((inputs(255)) xor (inputs(87)));
    layer0_outputs(2459) <= (inputs(5)) or (inputs(177));
    layer0_outputs(2460) <= not((inputs(43)) xor (inputs(31)));
    layer0_outputs(2461) <= not(inputs(217)) or (inputs(12));
    layer0_outputs(2462) <= not(inputs(235)) or (inputs(199));
    layer0_outputs(2463) <= inputs(53);
    layer0_outputs(2464) <= not((inputs(69)) and (inputs(19)));
    layer0_outputs(2465) <= not(inputs(92));
    layer0_outputs(2466) <= not(inputs(94));
    layer0_outputs(2467) <= inputs(102);
    layer0_outputs(2468) <= not(inputs(11)) or (inputs(250));
    layer0_outputs(2469) <= (inputs(120)) and not (inputs(178));
    layer0_outputs(2470) <= (inputs(53)) or (inputs(137));
    layer0_outputs(2471) <= not(inputs(89));
    layer0_outputs(2472) <= not(inputs(37));
    layer0_outputs(2473) <= inputs(150);
    layer0_outputs(2474) <= (inputs(189)) or (inputs(65));
    layer0_outputs(2475) <= not((inputs(190)) or (inputs(152)));
    layer0_outputs(2476) <= inputs(73);
    layer0_outputs(2477) <= (inputs(21)) and not (inputs(252));
    layer0_outputs(2478) <= (inputs(214)) and not (inputs(95));
    layer0_outputs(2479) <= not((inputs(22)) or (inputs(140)));
    layer0_outputs(2480) <= (inputs(131)) and not (inputs(95));
    layer0_outputs(2481) <= (inputs(209)) and not (inputs(117));
    layer0_outputs(2482) <= not((inputs(220)) xor (inputs(127)));
    layer0_outputs(2483) <= '0';
    layer0_outputs(2484) <= not(inputs(53));
    layer0_outputs(2485) <= not(inputs(132));
    layer0_outputs(2486) <= (inputs(237)) xor (inputs(12));
    layer0_outputs(2487) <= not((inputs(231)) or (inputs(248)));
    layer0_outputs(2488) <= not((inputs(95)) or (inputs(208)));
    layer0_outputs(2489) <= not(inputs(58)) or (inputs(53));
    layer0_outputs(2490) <= not(inputs(206));
    layer0_outputs(2491) <= (inputs(214)) xor (inputs(137));
    layer0_outputs(2492) <= (inputs(184)) and not (inputs(46));
    layer0_outputs(2493) <= (inputs(181)) xor (inputs(123));
    layer0_outputs(2494) <= (inputs(141)) xor (inputs(86));
    layer0_outputs(2495) <= '0';
    layer0_outputs(2496) <= (inputs(91)) or (inputs(31));
    layer0_outputs(2497) <= (inputs(199)) and not (inputs(78));
    layer0_outputs(2498) <= not(inputs(244)) or (inputs(89));
    layer0_outputs(2499) <= not(inputs(163));
    layer0_outputs(2500) <= not((inputs(45)) or (inputs(38)));
    layer0_outputs(2501) <= inputs(73);
    layer0_outputs(2502) <= not((inputs(78)) or (inputs(246)));
    layer0_outputs(2503) <= not(inputs(35)) or (inputs(112));
    layer0_outputs(2504) <= not(inputs(246)) or (inputs(61));
    layer0_outputs(2505) <= (inputs(149)) and not (inputs(47));
    layer0_outputs(2506) <= not((inputs(211)) or (inputs(217)));
    layer0_outputs(2507) <= not(inputs(106));
    layer0_outputs(2508) <= (inputs(56)) xor (inputs(204));
    layer0_outputs(2509) <= not(inputs(27));
    layer0_outputs(2510) <= not((inputs(139)) xor (inputs(57)));
    layer0_outputs(2511) <= (inputs(144)) or (inputs(156));
    layer0_outputs(2512) <= inputs(166);
    layer0_outputs(2513) <= not((inputs(112)) or (inputs(154)));
    layer0_outputs(2514) <= (inputs(183)) and (inputs(219));
    layer0_outputs(2515) <= (inputs(31)) xor (inputs(236));
    layer0_outputs(2516) <= (inputs(161)) or (inputs(230));
    layer0_outputs(2517) <= (inputs(251)) and (inputs(79));
    layer0_outputs(2518) <= not((inputs(92)) or (inputs(69)));
    layer0_outputs(2519) <= not((inputs(162)) or (inputs(17)));
    layer0_outputs(2520) <= not(inputs(162));
    layer0_outputs(2521) <= not(inputs(152));
    layer0_outputs(2522) <= not(inputs(114)) or (inputs(239));
    layer0_outputs(2523) <= (inputs(36)) and (inputs(132));
    layer0_outputs(2524) <= inputs(20);
    layer0_outputs(2525) <= not(inputs(91)) or (inputs(37));
    layer0_outputs(2526) <= (inputs(97)) or (inputs(53));
    layer0_outputs(2527) <= not((inputs(237)) or (inputs(225)));
    layer0_outputs(2528) <= (inputs(85)) and not (inputs(182));
    layer0_outputs(2529) <= (inputs(43)) or (inputs(125));
    layer0_outputs(2530) <= (inputs(71)) xor (inputs(72));
    layer0_outputs(2531) <= (inputs(73)) or (inputs(86));
    layer0_outputs(2532) <= not((inputs(214)) xor (inputs(161)));
    layer0_outputs(2533) <= not(inputs(204)) or (inputs(209));
    layer0_outputs(2534) <= not(inputs(171)) or (inputs(50));
    layer0_outputs(2535) <= not((inputs(128)) xor (inputs(108)));
    layer0_outputs(2536) <= not((inputs(204)) or (inputs(95)));
    layer0_outputs(2537) <= (inputs(11)) and (inputs(116));
    layer0_outputs(2538) <= not(inputs(41));
    layer0_outputs(2539) <= not((inputs(134)) and (inputs(135)));
    layer0_outputs(2540) <= not((inputs(60)) xor (inputs(37)));
    layer0_outputs(2541) <= not(inputs(37));
    layer0_outputs(2542) <= inputs(66);
    layer0_outputs(2543) <= (inputs(106)) or (inputs(122));
    layer0_outputs(2544) <= not(inputs(88)) or (inputs(60));
    layer0_outputs(2545) <= not((inputs(148)) or (inputs(92)));
    layer0_outputs(2546) <= not(inputs(149));
    layer0_outputs(2547) <= not(inputs(52)) or (inputs(227));
    layer0_outputs(2548) <= inputs(34);
    layer0_outputs(2549) <= (inputs(136)) and not (inputs(53));
    layer0_outputs(2550) <= (inputs(78)) and (inputs(75));
    layer0_outputs(2551) <= (inputs(19)) and not (inputs(129));
    layer0_outputs(2552) <= not(inputs(41)) or (inputs(153));
    layer0_outputs(2553) <= '0';
    layer0_outputs(2554) <= (inputs(204)) xor (inputs(200));
    layer0_outputs(2555) <= (inputs(186)) xor (inputs(99));
    layer0_outputs(2556) <= not(inputs(202)) or (inputs(126));
    layer0_outputs(2557) <= not(inputs(169));
    layer0_outputs(2558) <= not((inputs(183)) xor (inputs(178)));
    layer0_outputs(2559) <= (inputs(116)) and not (inputs(211));
    layer0_outputs(2560) <= (inputs(106)) or (inputs(16));
    layer0_outputs(2561) <= not(inputs(56)) or (inputs(109));
    layer0_outputs(2562) <= (inputs(114)) or (inputs(127));
    layer0_outputs(2563) <= not(inputs(145));
    layer0_outputs(2564) <= not((inputs(111)) or (inputs(196)));
    layer0_outputs(2565) <= (inputs(202)) and not (inputs(32));
    layer0_outputs(2566) <= not(inputs(86)) or (inputs(55));
    layer0_outputs(2567) <= not(inputs(78));
    layer0_outputs(2568) <= not(inputs(228));
    layer0_outputs(2569) <= (inputs(165)) and not (inputs(236));
    layer0_outputs(2570) <= not(inputs(169)) or (inputs(174));
    layer0_outputs(2571) <= not(inputs(89)) or (inputs(180));
    layer0_outputs(2572) <= not((inputs(138)) or (inputs(21)));
    layer0_outputs(2573) <= inputs(145);
    layer0_outputs(2574) <= not(inputs(196));
    layer0_outputs(2575) <= inputs(66);
    layer0_outputs(2576) <= not(inputs(167));
    layer0_outputs(2577) <= not(inputs(170)) or (inputs(105));
    layer0_outputs(2578) <= (inputs(160)) and not (inputs(254));
    layer0_outputs(2579) <= (inputs(252)) and not (inputs(144));
    layer0_outputs(2580) <= not((inputs(243)) xor (inputs(228)));
    layer0_outputs(2581) <= (inputs(135)) and not (inputs(165));
    layer0_outputs(2582) <= not(inputs(234)) or (inputs(107));
    layer0_outputs(2583) <= (inputs(140)) and not (inputs(47));
    layer0_outputs(2584) <= inputs(242);
    layer0_outputs(2585) <= not((inputs(201)) or (inputs(134)));
    layer0_outputs(2586) <= not((inputs(240)) or (inputs(11)));
    layer0_outputs(2587) <= (inputs(204)) or (inputs(197));
    layer0_outputs(2588) <= (inputs(246)) or (inputs(97));
    layer0_outputs(2589) <= inputs(44);
    layer0_outputs(2590) <= not(inputs(102)) or (inputs(178));
    layer0_outputs(2591) <= (inputs(120)) xor (inputs(182));
    layer0_outputs(2592) <= not((inputs(216)) and (inputs(20)));
    layer0_outputs(2593) <= not((inputs(147)) or (inputs(74)));
    layer0_outputs(2594) <= '0';
    layer0_outputs(2595) <= not(inputs(179)) or (inputs(206));
    layer0_outputs(2596) <= '1';
    layer0_outputs(2597) <= not((inputs(195)) or (inputs(247)));
    layer0_outputs(2598) <= not((inputs(188)) or (inputs(65)));
    layer0_outputs(2599) <= not((inputs(78)) or (inputs(213)));
    layer0_outputs(2600) <= (inputs(40)) and not (inputs(137));
    layer0_outputs(2601) <= (inputs(99)) or (inputs(85));
    layer0_outputs(2602) <= (inputs(130)) or (inputs(20));
    layer0_outputs(2603) <= not(inputs(53));
    layer0_outputs(2604) <= not(inputs(78));
    layer0_outputs(2605) <= not(inputs(61));
    layer0_outputs(2606) <= (inputs(10)) and not (inputs(50));
    layer0_outputs(2607) <= not((inputs(177)) xor (inputs(87)));
    layer0_outputs(2608) <= not((inputs(237)) xor (inputs(67)));
    layer0_outputs(2609) <= (inputs(64)) or (inputs(51));
    layer0_outputs(2610) <= inputs(91);
    layer0_outputs(2611) <= not(inputs(134)) or (inputs(1));
    layer0_outputs(2612) <= (inputs(30)) and not (inputs(130));
    layer0_outputs(2613) <= inputs(233);
    layer0_outputs(2614) <= not(inputs(38));
    layer0_outputs(2615) <= not(inputs(55));
    layer0_outputs(2616) <= not(inputs(194));
    layer0_outputs(2617) <= (inputs(165)) xor (inputs(132));
    layer0_outputs(2618) <= (inputs(106)) and (inputs(77));
    layer0_outputs(2619) <= (inputs(11)) xor (inputs(215));
    layer0_outputs(2620) <= (inputs(66)) and not (inputs(185));
    layer0_outputs(2621) <= inputs(106);
    layer0_outputs(2622) <= '0';
    layer0_outputs(2623) <= (inputs(98)) xor (inputs(62));
    layer0_outputs(2624) <= inputs(46);
    layer0_outputs(2625) <= (inputs(90)) and not (inputs(243));
    layer0_outputs(2626) <= not(inputs(50)) or (inputs(224));
    layer0_outputs(2627) <= (inputs(95)) or (inputs(207));
    layer0_outputs(2628) <= not(inputs(60));
    layer0_outputs(2629) <= inputs(56);
    layer0_outputs(2630) <= (inputs(164)) or (inputs(5));
    layer0_outputs(2631) <= not((inputs(212)) xor (inputs(146)));
    layer0_outputs(2632) <= not(inputs(114));
    layer0_outputs(2633) <= (inputs(52)) and not (inputs(4));
    layer0_outputs(2634) <= inputs(153);
    layer0_outputs(2635) <= not(inputs(169)) or (inputs(37));
    layer0_outputs(2636) <= not((inputs(96)) xor (inputs(88)));
    layer0_outputs(2637) <= (inputs(227)) or (inputs(149));
    layer0_outputs(2638) <= not((inputs(132)) or (inputs(146)));
    layer0_outputs(2639) <= not((inputs(76)) or (inputs(43)));
    layer0_outputs(2640) <= not(inputs(130));
    layer0_outputs(2641) <= (inputs(37)) or (inputs(225));
    layer0_outputs(2642) <= not((inputs(35)) or (inputs(32)));
    layer0_outputs(2643) <= inputs(24);
    layer0_outputs(2644) <= inputs(34);
    layer0_outputs(2645) <= not((inputs(201)) or (inputs(255)));
    layer0_outputs(2646) <= (inputs(161)) or (inputs(211));
    layer0_outputs(2647) <= (inputs(220)) and not (inputs(81));
    layer0_outputs(2648) <= not(inputs(130)) or (inputs(76));
    layer0_outputs(2649) <= inputs(155);
    layer0_outputs(2650) <= (inputs(179)) or (inputs(6));
    layer0_outputs(2651) <= not((inputs(82)) or (inputs(145)));
    layer0_outputs(2652) <= (inputs(35)) and not (inputs(203));
    layer0_outputs(2653) <= not((inputs(106)) and (inputs(246)));
    layer0_outputs(2654) <= not(inputs(142)) or (inputs(48));
    layer0_outputs(2655) <= inputs(52);
    layer0_outputs(2656) <= (inputs(164)) or (inputs(246));
    layer0_outputs(2657) <= (inputs(192)) or (inputs(207));
    layer0_outputs(2658) <= (inputs(205)) or (inputs(158));
    layer0_outputs(2659) <= (inputs(189)) and not (inputs(96));
    layer0_outputs(2660) <= (inputs(117)) and not (inputs(185));
    layer0_outputs(2661) <= '0';
    layer0_outputs(2662) <= not((inputs(194)) and (inputs(143)));
    layer0_outputs(2663) <= not((inputs(243)) and (inputs(157)));
    layer0_outputs(2664) <= not(inputs(205)) or (inputs(16));
    layer0_outputs(2665) <= not((inputs(232)) and (inputs(162)));
    layer0_outputs(2666) <= (inputs(79)) or (inputs(214));
    layer0_outputs(2667) <= not((inputs(97)) xor (inputs(165)));
    layer0_outputs(2668) <= not((inputs(223)) xor (inputs(49)));
    layer0_outputs(2669) <= not((inputs(109)) or (inputs(59)));
    layer0_outputs(2670) <= not(inputs(184)) or (inputs(74));
    layer0_outputs(2671) <= not(inputs(93)) or (inputs(30));
    layer0_outputs(2672) <= inputs(225);
    layer0_outputs(2673) <= (inputs(122)) or (inputs(193));
    layer0_outputs(2674) <= not((inputs(255)) or (inputs(219)));
    layer0_outputs(2675) <= (inputs(182)) or (inputs(83));
    layer0_outputs(2676) <= not((inputs(109)) or (inputs(21)));
    layer0_outputs(2677) <= (inputs(228)) and not (inputs(252));
    layer0_outputs(2678) <= not(inputs(149)) or (inputs(227));
    layer0_outputs(2679) <= (inputs(229)) or (inputs(116));
    layer0_outputs(2680) <= not(inputs(253)) or (inputs(225));
    layer0_outputs(2681) <= not((inputs(170)) xor (inputs(69)));
    layer0_outputs(2682) <= (inputs(55)) and not (inputs(162));
    layer0_outputs(2683) <= not(inputs(90)) or (inputs(32));
    layer0_outputs(2684) <= (inputs(124)) xor (inputs(27));
    layer0_outputs(2685) <= not(inputs(211));
    layer0_outputs(2686) <= not(inputs(33));
    layer0_outputs(2687) <= not(inputs(149)) or (inputs(3));
    layer0_outputs(2688) <= not(inputs(181));
    layer0_outputs(2689) <= not(inputs(197));
    layer0_outputs(2690) <= not(inputs(73));
    layer0_outputs(2691) <= not((inputs(11)) xor (inputs(45)));
    layer0_outputs(2692) <= inputs(146);
    layer0_outputs(2693) <= (inputs(59)) and not (inputs(86));
    layer0_outputs(2694) <= inputs(68);
    layer0_outputs(2695) <= inputs(15);
    layer0_outputs(2696) <= not(inputs(120));
    layer0_outputs(2697) <= not(inputs(227));
    layer0_outputs(2698) <= (inputs(80)) xor (inputs(103));
    layer0_outputs(2699) <= not(inputs(21));
    layer0_outputs(2700) <= not(inputs(20));
    layer0_outputs(2701) <= (inputs(142)) and not (inputs(39));
    layer0_outputs(2702) <= not(inputs(243));
    layer0_outputs(2703) <= (inputs(189)) or (inputs(209));
    layer0_outputs(2704) <= not(inputs(106)) or (inputs(148));
    layer0_outputs(2705) <= inputs(141);
    layer0_outputs(2706) <= (inputs(166)) and not (inputs(207));
    layer0_outputs(2707) <= (inputs(172)) and (inputs(183));
    layer0_outputs(2708) <= (inputs(129)) xor (inputs(114));
    layer0_outputs(2709) <= not((inputs(94)) or (inputs(47)));
    layer0_outputs(2710) <= (inputs(252)) or (inputs(103));
    layer0_outputs(2711) <= (inputs(209)) and not (inputs(235));
    layer0_outputs(2712) <= (inputs(111)) xor (inputs(179));
    layer0_outputs(2713) <= not((inputs(1)) or (inputs(50)));
    layer0_outputs(2714) <= (inputs(252)) or (inputs(238));
    layer0_outputs(2715) <= inputs(82);
    layer0_outputs(2716) <= not(inputs(146)) or (inputs(127));
    layer0_outputs(2717) <= (inputs(115)) xor (inputs(187));
    layer0_outputs(2718) <= (inputs(78)) or (inputs(254));
    layer0_outputs(2719) <= (inputs(79)) xor (inputs(105));
    layer0_outputs(2720) <= not((inputs(69)) and (inputs(25)));
    layer0_outputs(2721) <= not((inputs(32)) and (inputs(7)));
    layer0_outputs(2722) <= not((inputs(75)) xor (inputs(192)));
    layer0_outputs(2723) <= not(inputs(39)) or (inputs(150));
    layer0_outputs(2724) <= not(inputs(89)) or (inputs(33));
    layer0_outputs(2725) <= (inputs(219)) and not (inputs(5));
    layer0_outputs(2726) <= not(inputs(227));
    layer0_outputs(2727) <= not(inputs(235));
    layer0_outputs(2728) <= not(inputs(251));
    layer0_outputs(2729) <= (inputs(91)) and not (inputs(186));
    layer0_outputs(2730) <= (inputs(221)) xor (inputs(49));
    layer0_outputs(2731) <= (inputs(84)) or (inputs(160));
    layer0_outputs(2732) <= not(inputs(163));
    layer0_outputs(2733) <= not((inputs(215)) or (inputs(241)));
    layer0_outputs(2734) <= not((inputs(109)) xor (inputs(150)));
    layer0_outputs(2735) <= not((inputs(128)) or (inputs(177)));
    layer0_outputs(2736) <= inputs(196);
    layer0_outputs(2737) <= not(inputs(3));
    layer0_outputs(2738) <= inputs(114);
    layer0_outputs(2739) <= not(inputs(140)) or (inputs(113));
    layer0_outputs(2740) <= (inputs(177)) and not (inputs(223));
    layer0_outputs(2741) <= not((inputs(189)) or (inputs(63)));
    layer0_outputs(2742) <= not((inputs(125)) or (inputs(122)));
    layer0_outputs(2743) <= not(inputs(146));
    layer0_outputs(2744) <= not(inputs(118)) or (inputs(105));
    layer0_outputs(2745) <= not((inputs(21)) or (inputs(0)));
    layer0_outputs(2746) <= inputs(182);
    layer0_outputs(2747) <= inputs(192);
    layer0_outputs(2748) <= not((inputs(106)) or (inputs(73)));
    layer0_outputs(2749) <= not((inputs(81)) or (inputs(60)));
    layer0_outputs(2750) <= inputs(108);
    layer0_outputs(2751) <= inputs(85);
    layer0_outputs(2752) <= (inputs(10)) and not (inputs(102));
    layer0_outputs(2753) <= not(inputs(32));
    layer0_outputs(2754) <= not(inputs(90)) or (inputs(223));
    layer0_outputs(2755) <= not((inputs(5)) xor (inputs(18)));
    layer0_outputs(2756) <= (inputs(211)) and not (inputs(91));
    layer0_outputs(2757) <= not((inputs(17)) or (inputs(235)));
    layer0_outputs(2758) <= (inputs(123)) xor (inputs(104));
    layer0_outputs(2759) <= not(inputs(182)) or (inputs(49));
    layer0_outputs(2760) <= not((inputs(74)) or (inputs(147)));
    layer0_outputs(2761) <= inputs(158);
    layer0_outputs(2762) <= '1';
    layer0_outputs(2763) <= (inputs(116)) xor (inputs(70));
    layer0_outputs(2764) <= not(inputs(104));
    layer0_outputs(2765) <= not(inputs(239)) or (inputs(216));
    layer0_outputs(2766) <= not(inputs(145)) or (inputs(168));
    layer0_outputs(2767) <= not((inputs(20)) or (inputs(4)));
    layer0_outputs(2768) <= not(inputs(64));
    layer0_outputs(2769) <= not((inputs(203)) or (inputs(94)));
    layer0_outputs(2770) <= inputs(13);
    layer0_outputs(2771) <= not((inputs(226)) or (inputs(232)));
    layer0_outputs(2772) <= not(inputs(117));
    layer0_outputs(2773) <= (inputs(192)) or (inputs(226));
    layer0_outputs(2774) <= (inputs(181)) or (inputs(107));
    layer0_outputs(2775) <= not((inputs(6)) or (inputs(124)));
    layer0_outputs(2776) <= (inputs(232)) and not (inputs(95));
    layer0_outputs(2777) <= not(inputs(238)) or (inputs(142));
    layer0_outputs(2778) <= not((inputs(62)) xor (inputs(4)));
    layer0_outputs(2779) <= (inputs(101)) or (inputs(70));
    layer0_outputs(2780) <= not((inputs(214)) xor (inputs(21)));
    layer0_outputs(2781) <= not((inputs(167)) or (inputs(4)));
    layer0_outputs(2782) <= '0';
    layer0_outputs(2783) <= not(inputs(41));
    layer0_outputs(2784) <= not(inputs(194)) or (inputs(201));
    layer0_outputs(2785) <= (inputs(2)) xor (inputs(247));
    layer0_outputs(2786) <= inputs(116);
    layer0_outputs(2787) <= not((inputs(68)) or (inputs(137)));
    layer0_outputs(2788) <= not((inputs(97)) xor (inputs(177)));
    layer0_outputs(2789) <= '1';
    layer0_outputs(2790) <= not(inputs(14));
    layer0_outputs(2791) <= (inputs(30)) or (inputs(97));
    layer0_outputs(2792) <= not((inputs(72)) or (inputs(221)));
    layer0_outputs(2793) <= inputs(40);
    layer0_outputs(2794) <= (inputs(167)) and not (inputs(80));
    layer0_outputs(2795) <= not(inputs(29));
    layer0_outputs(2796) <= inputs(22);
    layer0_outputs(2797) <= not(inputs(247)) or (inputs(144));
    layer0_outputs(2798) <= not((inputs(122)) xor (inputs(60)));
    layer0_outputs(2799) <= not(inputs(176));
    layer0_outputs(2800) <= not(inputs(53));
    layer0_outputs(2801) <= (inputs(59)) or (inputs(70));
    layer0_outputs(2802) <= not((inputs(11)) xor (inputs(91)));
    layer0_outputs(2803) <= inputs(92);
    layer0_outputs(2804) <= not((inputs(226)) or (inputs(35)));
    layer0_outputs(2805) <= inputs(101);
    layer0_outputs(2806) <= (inputs(149)) or (inputs(50));
    layer0_outputs(2807) <= (inputs(220)) or (inputs(97));
    layer0_outputs(2808) <= inputs(146);
    layer0_outputs(2809) <= (inputs(193)) xor (inputs(219));
    layer0_outputs(2810) <= not((inputs(14)) or (inputs(10)));
    layer0_outputs(2811) <= (inputs(204)) and not (inputs(34));
    layer0_outputs(2812) <= inputs(231);
    layer0_outputs(2813) <= (inputs(182)) or (inputs(240));
    layer0_outputs(2814) <= not((inputs(128)) xor (inputs(132)));
    layer0_outputs(2815) <= not((inputs(196)) xor (inputs(216)));
    layer0_outputs(2816) <= not(inputs(228)) or (inputs(148));
    layer0_outputs(2817) <= not((inputs(60)) xor (inputs(46)));
    layer0_outputs(2818) <= not(inputs(70));
    layer0_outputs(2819) <= not(inputs(61));
    layer0_outputs(2820) <= inputs(98);
    layer0_outputs(2821) <= '0';
    layer0_outputs(2822) <= (inputs(152)) or (inputs(137));
    layer0_outputs(2823) <= not((inputs(206)) or (inputs(248)));
    layer0_outputs(2824) <= not((inputs(50)) or (inputs(44)));
    layer0_outputs(2825) <= '1';
    layer0_outputs(2826) <= inputs(179);
    layer0_outputs(2827) <= not((inputs(136)) or (inputs(36)));
    layer0_outputs(2828) <= not(inputs(234)) or (inputs(77));
    layer0_outputs(2829) <= inputs(213);
    layer0_outputs(2830) <= not((inputs(235)) and (inputs(6)));
    layer0_outputs(2831) <= not(inputs(235));
    layer0_outputs(2832) <= (inputs(63)) or (inputs(17));
    layer0_outputs(2833) <= not(inputs(182));
    layer0_outputs(2834) <= not(inputs(55));
    layer0_outputs(2835) <= not((inputs(17)) xor (inputs(124)));
    layer0_outputs(2836) <= (inputs(52)) and not (inputs(249));
    layer0_outputs(2837) <= (inputs(139)) and not (inputs(147));
    layer0_outputs(2838) <= not((inputs(148)) xor (inputs(234)));
    layer0_outputs(2839) <= inputs(62);
    layer0_outputs(2840) <= inputs(104);
    layer0_outputs(2841) <= (inputs(186)) xor (inputs(113));
    layer0_outputs(2842) <= inputs(52);
    layer0_outputs(2843) <= inputs(134);
    layer0_outputs(2844) <= not(inputs(77));
    layer0_outputs(2845) <= not((inputs(224)) xor (inputs(133)));
    layer0_outputs(2846) <= not((inputs(199)) or (inputs(223)));
    layer0_outputs(2847) <= inputs(100);
    layer0_outputs(2848) <= not(inputs(254));
    layer0_outputs(2849) <= inputs(121);
    layer0_outputs(2850) <= (inputs(82)) or (inputs(101));
    layer0_outputs(2851) <= not((inputs(142)) or (inputs(152)));
    layer0_outputs(2852) <= not(inputs(142)) or (inputs(146));
    layer0_outputs(2853) <= not(inputs(162));
    layer0_outputs(2854) <= inputs(153);
    layer0_outputs(2855) <= inputs(86);
    layer0_outputs(2856) <= not((inputs(220)) xor (inputs(188)));
    layer0_outputs(2857) <= inputs(228);
    layer0_outputs(2858) <= inputs(107);
    layer0_outputs(2859) <= not((inputs(132)) xor (inputs(64)));
    layer0_outputs(2860) <= inputs(3);
    layer0_outputs(2861) <= not(inputs(77));
    layer0_outputs(2862) <= (inputs(171)) and not (inputs(67));
    layer0_outputs(2863) <= (inputs(1)) or (inputs(88));
    layer0_outputs(2864) <= not(inputs(176));
    layer0_outputs(2865) <= not(inputs(68));
    layer0_outputs(2866) <= inputs(181);
    layer0_outputs(2867) <= not((inputs(189)) or (inputs(216)));
    layer0_outputs(2868) <= (inputs(116)) and not (inputs(148));
    layer0_outputs(2869) <= not((inputs(205)) and (inputs(205)));
    layer0_outputs(2870) <= not((inputs(198)) or (inputs(5)));
    layer0_outputs(2871) <= not((inputs(15)) or (inputs(110)));
    layer0_outputs(2872) <= (inputs(84)) and not (inputs(1));
    layer0_outputs(2873) <= not((inputs(213)) xor (inputs(157)));
    layer0_outputs(2874) <= inputs(175);
    layer0_outputs(2875) <= (inputs(20)) and not (inputs(144));
    layer0_outputs(2876) <= not((inputs(39)) or (inputs(63)));
    layer0_outputs(2877) <= not(inputs(234)) or (inputs(94));
    layer0_outputs(2878) <= (inputs(1)) or (inputs(36));
    layer0_outputs(2879) <= (inputs(56)) or (inputs(5));
    layer0_outputs(2880) <= '0';
    layer0_outputs(2881) <= '1';
    layer0_outputs(2882) <= (inputs(22)) and not (inputs(249));
    layer0_outputs(2883) <= not((inputs(143)) or (inputs(202)));
    layer0_outputs(2884) <= (inputs(186)) and not (inputs(61));
    layer0_outputs(2885) <= not((inputs(111)) or (inputs(95)));
    layer0_outputs(2886) <= (inputs(151)) or (inputs(194));
    layer0_outputs(2887) <= not(inputs(94));
    layer0_outputs(2888) <= (inputs(150)) or (inputs(114));
    layer0_outputs(2889) <= '0';
    layer0_outputs(2890) <= inputs(82);
    layer0_outputs(2891) <= not(inputs(224)) or (inputs(112));
    layer0_outputs(2892) <= not((inputs(139)) xor (inputs(140)));
    layer0_outputs(2893) <= not(inputs(94));
    layer0_outputs(2894) <= (inputs(57)) and not (inputs(199));
    layer0_outputs(2895) <= not((inputs(206)) or (inputs(166)));
    layer0_outputs(2896) <= (inputs(86)) xor (inputs(8));
    layer0_outputs(2897) <= (inputs(117)) and not (inputs(125));
    layer0_outputs(2898) <= inputs(232);
    layer0_outputs(2899) <= not((inputs(214)) or (inputs(71)));
    layer0_outputs(2900) <= not((inputs(243)) xor (inputs(198)));
    layer0_outputs(2901) <= not(inputs(100));
    layer0_outputs(2902) <= inputs(119);
    layer0_outputs(2903) <= not(inputs(104));
    layer0_outputs(2904) <= not((inputs(204)) or (inputs(50)));
    layer0_outputs(2905) <= inputs(51);
    layer0_outputs(2906) <= inputs(31);
    layer0_outputs(2907) <= not((inputs(49)) or (inputs(236)));
    layer0_outputs(2908) <= (inputs(59)) and (inputs(99));
    layer0_outputs(2909) <= '1';
    layer0_outputs(2910) <= not(inputs(252));
    layer0_outputs(2911) <= '0';
    layer0_outputs(2912) <= not((inputs(31)) or (inputs(20)));
    layer0_outputs(2913) <= (inputs(223)) xor (inputs(11));
    layer0_outputs(2914) <= not(inputs(207));
    layer0_outputs(2915) <= not(inputs(231));
    layer0_outputs(2916) <= not((inputs(33)) or (inputs(177)));
    layer0_outputs(2917) <= (inputs(65)) xor (inputs(165));
    layer0_outputs(2918) <= inputs(166);
    layer0_outputs(2919) <= not((inputs(112)) or (inputs(89)));
    layer0_outputs(2920) <= '0';
    layer0_outputs(2921) <= not(inputs(217));
    layer0_outputs(2922) <= inputs(100);
    layer0_outputs(2923) <= inputs(134);
    layer0_outputs(2924) <= not(inputs(163));
    layer0_outputs(2925) <= (inputs(158)) or (inputs(33));
    layer0_outputs(2926) <= (inputs(232)) and (inputs(197));
    layer0_outputs(2927) <= (inputs(40)) or (inputs(191));
    layer0_outputs(2928) <= (inputs(86)) or (inputs(85));
    layer0_outputs(2929) <= not((inputs(124)) or (inputs(67)));
    layer0_outputs(2930) <= (inputs(28)) xor (inputs(144));
    layer0_outputs(2931) <= '1';
    layer0_outputs(2932) <= '0';
    layer0_outputs(2933) <= inputs(107);
    layer0_outputs(2934) <= not(inputs(228));
    layer0_outputs(2935) <= not(inputs(210));
    layer0_outputs(2936) <= (inputs(5)) or (inputs(190));
    layer0_outputs(2937) <= (inputs(224)) xor (inputs(180));
    layer0_outputs(2938) <= not((inputs(17)) or (inputs(246)));
    layer0_outputs(2939) <= not(inputs(86));
    layer0_outputs(2940) <= not((inputs(241)) or (inputs(3)));
    layer0_outputs(2941) <= not((inputs(221)) or (inputs(209)));
    layer0_outputs(2942) <= not(inputs(243)) or (inputs(50));
    layer0_outputs(2943) <= not(inputs(229));
    layer0_outputs(2944) <= not(inputs(85));
    layer0_outputs(2945) <= inputs(52);
    layer0_outputs(2946) <= (inputs(194)) and not (inputs(112));
    layer0_outputs(2947) <= inputs(248);
    layer0_outputs(2948) <= not((inputs(148)) xor (inputs(79)));
    layer0_outputs(2949) <= (inputs(169)) or (inputs(14));
    layer0_outputs(2950) <= not(inputs(198));
    layer0_outputs(2951) <= (inputs(219)) or (inputs(145));
    layer0_outputs(2952) <= (inputs(66)) and not (inputs(15));
    layer0_outputs(2953) <= not(inputs(40));
    layer0_outputs(2954) <= not((inputs(188)) xor (inputs(99)));
    layer0_outputs(2955) <= not(inputs(142)) or (inputs(42));
    layer0_outputs(2956) <= not((inputs(217)) xor (inputs(25)));
    layer0_outputs(2957) <= inputs(20);
    layer0_outputs(2958) <= not(inputs(24));
    layer0_outputs(2959) <= inputs(23);
    layer0_outputs(2960) <= not(inputs(25)) or (inputs(158));
    layer0_outputs(2961) <= not((inputs(219)) xor (inputs(177)));
    layer0_outputs(2962) <= not(inputs(41));
    layer0_outputs(2963) <= not((inputs(183)) xor (inputs(111)));
    layer0_outputs(2964) <= not(inputs(68));
    layer0_outputs(2965) <= not((inputs(147)) or (inputs(177)));
    layer0_outputs(2966) <= not(inputs(230));
    layer0_outputs(2967) <= not((inputs(247)) or (inputs(147)));
    layer0_outputs(2968) <= not(inputs(137));
    layer0_outputs(2969) <= not(inputs(113));
    layer0_outputs(2970) <= (inputs(204)) or (inputs(179));
    layer0_outputs(2971) <= not(inputs(117)) or (inputs(34));
    layer0_outputs(2972) <= (inputs(245)) and not (inputs(96));
    layer0_outputs(2973) <= not(inputs(219));
    layer0_outputs(2974) <= (inputs(199)) or (inputs(32));
    layer0_outputs(2975) <= (inputs(166)) xor (inputs(78));
    layer0_outputs(2976) <= not(inputs(107)) or (inputs(24));
    layer0_outputs(2977) <= not(inputs(39));
    layer0_outputs(2978) <= not((inputs(57)) and (inputs(247)));
    layer0_outputs(2979) <= inputs(97);
    layer0_outputs(2980) <= not(inputs(117)) or (inputs(162));
    layer0_outputs(2981) <= inputs(248);
    layer0_outputs(2982) <= inputs(164);
    layer0_outputs(2983) <= (inputs(255)) or (inputs(244));
    layer0_outputs(2984) <= not(inputs(24)) or (inputs(158));
    layer0_outputs(2985) <= not((inputs(1)) or (inputs(32)));
    layer0_outputs(2986) <= (inputs(163)) and not (inputs(65));
    layer0_outputs(2987) <= not(inputs(221));
    layer0_outputs(2988) <= not((inputs(225)) xor (inputs(211)));
    layer0_outputs(2989) <= not(inputs(24));
    layer0_outputs(2990) <= (inputs(55)) and not (inputs(149));
    layer0_outputs(2991) <= inputs(158);
    layer0_outputs(2992) <= (inputs(72)) and (inputs(66));
    layer0_outputs(2993) <= inputs(135);
    layer0_outputs(2994) <= (inputs(213)) and (inputs(237));
    layer0_outputs(2995) <= not(inputs(231)) or (inputs(77));
    layer0_outputs(2996) <= not(inputs(71)) or (inputs(254));
    layer0_outputs(2997) <= (inputs(3)) or (inputs(222));
    layer0_outputs(2998) <= not(inputs(96));
    layer0_outputs(2999) <= (inputs(106)) or (inputs(23));
    layer0_outputs(3000) <= not(inputs(94));
    layer0_outputs(3001) <= not(inputs(135));
    layer0_outputs(3002) <= inputs(194);
    layer0_outputs(3003) <= inputs(10);
    layer0_outputs(3004) <= (inputs(135)) and not (inputs(65));
    layer0_outputs(3005) <= inputs(226);
    layer0_outputs(3006) <= (inputs(124)) or (inputs(116));
    layer0_outputs(3007) <= '0';
    layer0_outputs(3008) <= not((inputs(248)) or (inputs(101)));
    layer0_outputs(3009) <= inputs(57);
    layer0_outputs(3010) <= (inputs(62)) xor (inputs(76));
    layer0_outputs(3011) <= (inputs(206)) xor (inputs(78));
    layer0_outputs(3012) <= not(inputs(131));
    layer0_outputs(3013) <= inputs(24);
    layer0_outputs(3014) <= not(inputs(176)) or (inputs(240));
    layer0_outputs(3015) <= inputs(72);
    layer0_outputs(3016) <= not(inputs(240));
    layer0_outputs(3017) <= (inputs(115)) and not (inputs(4));
    layer0_outputs(3018) <= not(inputs(28)) or (inputs(245));
    layer0_outputs(3019) <= not((inputs(206)) xor (inputs(249)));
    layer0_outputs(3020) <= (inputs(172)) and not (inputs(83));
    layer0_outputs(3021) <= (inputs(105)) or (inputs(31));
    layer0_outputs(3022) <= inputs(12);
    layer0_outputs(3023) <= not(inputs(101));
    layer0_outputs(3024) <= inputs(206);
    layer0_outputs(3025) <= not((inputs(152)) or (inputs(93)));
    layer0_outputs(3026) <= not((inputs(112)) xor (inputs(69)));
    layer0_outputs(3027) <= (inputs(232)) and not (inputs(46));
    layer0_outputs(3028) <= not(inputs(21));
    layer0_outputs(3029) <= not(inputs(98));
    layer0_outputs(3030) <= not(inputs(131));
    layer0_outputs(3031) <= (inputs(165)) or (inputs(251));
    layer0_outputs(3032) <= not(inputs(215));
    layer0_outputs(3033) <= (inputs(228)) and not (inputs(132));
    layer0_outputs(3034) <= (inputs(109)) or (inputs(85));
    layer0_outputs(3035) <= inputs(132);
    layer0_outputs(3036) <= inputs(71);
    layer0_outputs(3037) <= (inputs(102)) and not (inputs(252));
    layer0_outputs(3038) <= (inputs(253)) xor (inputs(198));
    layer0_outputs(3039) <= (inputs(35)) or (inputs(146));
    layer0_outputs(3040) <= not((inputs(3)) xor (inputs(26)));
    layer0_outputs(3041) <= not(inputs(114));
    layer0_outputs(3042) <= (inputs(118)) and not (inputs(116));
    layer0_outputs(3043) <= (inputs(98)) or (inputs(239));
    layer0_outputs(3044) <= inputs(48);
    layer0_outputs(3045) <= (inputs(235)) xor (inputs(176));
    layer0_outputs(3046) <= (inputs(70)) and not (inputs(239));
    layer0_outputs(3047) <= not((inputs(196)) or (inputs(61)));
    layer0_outputs(3048) <= not((inputs(63)) or (inputs(80)));
    layer0_outputs(3049) <= not((inputs(189)) or (inputs(148)));
    layer0_outputs(3050) <= not((inputs(205)) or (inputs(40)));
    layer0_outputs(3051) <= '0';
    layer0_outputs(3052) <= (inputs(241)) or (inputs(175));
    layer0_outputs(3053) <= (inputs(182)) xor (inputs(245));
    layer0_outputs(3054) <= (inputs(69)) and not (inputs(94));
    layer0_outputs(3055) <= not((inputs(100)) or (inputs(14)));
    layer0_outputs(3056) <= inputs(187);
    layer0_outputs(3057) <= not(inputs(198));
    layer0_outputs(3058) <= (inputs(206)) or (inputs(14));
    layer0_outputs(3059) <= (inputs(199)) and not (inputs(97));
    layer0_outputs(3060) <= not(inputs(78));
    layer0_outputs(3061) <= (inputs(67)) or (inputs(5));
    layer0_outputs(3062) <= (inputs(153)) and not (inputs(33));
    layer0_outputs(3063) <= inputs(104);
    layer0_outputs(3064) <= not(inputs(62)) or (inputs(129));
    layer0_outputs(3065) <= (inputs(115)) and (inputs(27));
    layer0_outputs(3066) <= not(inputs(43)) or (inputs(34));
    layer0_outputs(3067) <= inputs(215);
    layer0_outputs(3068) <= not(inputs(195)) or (inputs(93));
    layer0_outputs(3069) <= not((inputs(170)) or (inputs(142)));
    layer0_outputs(3070) <= not((inputs(111)) or (inputs(252)));
    layer0_outputs(3071) <= not(inputs(167)) or (inputs(186));
    layer0_outputs(3072) <= (inputs(119)) and not (inputs(26));
    layer0_outputs(3073) <= not((inputs(117)) and (inputs(52)));
    layer0_outputs(3074) <= not(inputs(103));
    layer0_outputs(3075) <= not((inputs(87)) xor (inputs(207)));
    layer0_outputs(3076) <= not((inputs(54)) xor (inputs(23)));
    layer0_outputs(3077) <= not(inputs(10)) or (inputs(191));
    layer0_outputs(3078) <= (inputs(36)) or (inputs(141));
    layer0_outputs(3079) <= inputs(166);
    layer0_outputs(3080) <= not(inputs(87)) or (inputs(76));
    layer0_outputs(3081) <= inputs(26);
    layer0_outputs(3082) <= inputs(169);
    layer0_outputs(3083) <= (inputs(196)) and not (inputs(6));
    layer0_outputs(3084) <= (inputs(93)) and not (inputs(176));
    layer0_outputs(3085) <= not(inputs(231));
    layer0_outputs(3086) <= not(inputs(188));
    layer0_outputs(3087) <= inputs(161);
    layer0_outputs(3088) <= inputs(68);
    layer0_outputs(3089) <= '0';
    layer0_outputs(3090) <= '0';
    layer0_outputs(3091) <= inputs(85);
    layer0_outputs(3092) <= not(inputs(133));
    layer0_outputs(3093) <= not(inputs(234)) or (inputs(54));
    layer0_outputs(3094) <= not(inputs(128));
    layer0_outputs(3095) <= not(inputs(12));
    layer0_outputs(3096) <= not(inputs(211));
    layer0_outputs(3097) <= (inputs(182)) or (inputs(56));
    layer0_outputs(3098) <= not(inputs(168));
    layer0_outputs(3099) <= (inputs(148)) xor (inputs(107));
    layer0_outputs(3100) <= (inputs(74)) xor (inputs(107));
    layer0_outputs(3101) <= inputs(121);
    layer0_outputs(3102) <= not(inputs(95));
    layer0_outputs(3103) <= not((inputs(188)) or (inputs(157)));
    layer0_outputs(3104) <= inputs(222);
    layer0_outputs(3105) <= not((inputs(46)) and (inputs(199)));
    layer0_outputs(3106) <= '0';
    layer0_outputs(3107) <= (inputs(189)) and not (inputs(192));
    layer0_outputs(3108) <= inputs(244);
    layer0_outputs(3109) <= inputs(169);
    layer0_outputs(3110) <= not(inputs(248));
    layer0_outputs(3111) <= not(inputs(126));
    layer0_outputs(3112) <= '1';
    layer0_outputs(3113) <= (inputs(106)) and not (inputs(180));
    layer0_outputs(3114) <= inputs(59);
    layer0_outputs(3115) <= not(inputs(93)) or (inputs(15));
    layer0_outputs(3116) <= (inputs(217)) or (inputs(220));
    layer0_outputs(3117) <= (inputs(245)) xor (inputs(252));
    layer0_outputs(3118) <= inputs(41);
    layer0_outputs(3119) <= inputs(78);
    layer0_outputs(3120) <= not(inputs(107));
    layer0_outputs(3121) <= not((inputs(207)) or (inputs(82)));
    layer0_outputs(3122) <= not((inputs(39)) or (inputs(211)));
    layer0_outputs(3123) <= not((inputs(162)) and (inputs(125)));
    layer0_outputs(3124) <= not(inputs(196));
    layer0_outputs(3125) <= inputs(9);
    layer0_outputs(3126) <= (inputs(140)) and not (inputs(157));
    layer0_outputs(3127) <= not(inputs(75));
    layer0_outputs(3128) <= not(inputs(157));
    layer0_outputs(3129) <= (inputs(195)) xor (inputs(221));
    layer0_outputs(3130) <= (inputs(75)) or (inputs(126));
    layer0_outputs(3131) <= not((inputs(249)) or (inputs(17)));
    layer0_outputs(3132) <= '0';
    layer0_outputs(3133) <= not(inputs(139)) or (inputs(206));
    layer0_outputs(3134) <= not(inputs(113));
    layer0_outputs(3135) <= (inputs(21)) xor (inputs(96));
    layer0_outputs(3136) <= (inputs(225)) and not (inputs(241));
    layer0_outputs(3137) <= (inputs(42)) and not (inputs(147));
    layer0_outputs(3138) <= not((inputs(31)) xor (inputs(11)));
    layer0_outputs(3139) <= inputs(94);
    layer0_outputs(3140) <= not((inputs(186)) or (inputs(80)));
    layer0_outputs(3141) <= (inputs(138)) and (inputs(169));
    layer0_outputs(3142) <= not((inputs(2)) xor (inputs(172)));
    layer0_outputs(3143) <= inputs(174);
    layer0_outputs(3144) <= not((inputs(171)) or (inputs(204)));
    layer0_outputs(3145) <= inputs(170);
    layer0_outputs(3146) <= not(inputs(218));
    layer0_outputs(3147) <= (inputs(124)) or (inputs(42));
    layer0_outputs(3148) <= not((inputs(72)) or (inputs(143)));
    layer0_outputs(3149) <= inputs(113);
    layer0_outputs(3150) <= not(inputs(88));
    layer0_outputs(3151) <= not((inputs(147)) xor (inputs(162)));
    layer0_outputs(3152) <= not(inputs(113));
    layer0_outputs(3153) <= not((inputs(127)) or (inputs(63)));
    layer0_outputs(3154) <= not((inputs(159)) or (inputs(244)));
    layer0_outputs(3155) <= inputs(221);
    layer0_outputs(3156) <= (inputs(185)) or (inputs(48));
    layer0_outputs(3157) <= inputs(163);
    layer0_outputs(3158) <= (inputs(155)) and (inputs(247));
    layer0_outputs(3159) <= not(inputs(210));
    layer0_outputs(3160) <= inputs(202);
    layer0_outputs(3161) <= not(inputs(52)) or (inputs(238));
    layer0_outputs(3162) <= (inputs(85)) and not (inputs(253));
    layer0_outputs(3163) <= not(inputs(128)) or (inputs(61));
    layer0_outputs(3164) <= (inputs(183)) or (inputs(27));
    layer0_outputs(3165) <= (inputs(159)) and not (inputs(173));
    layer0_outputs(3166) <= not((inputs(244)) or (inputs(11)));
    layer0_outputs(3167) <= not((inputs(143)) and (inputs(65)));
    layer0_outputs(3168) <= (inputs(100)) or (inputs(230));
    layer0_outputs(3169) <= (inputs(191)) xor (inputs(126));
    layer0_outputs(3170) <= (inputs(152)) or (inputs(33));
    layer0_outputs(3171) <= not((inputs(216)) xor (inputs(172)));
    layer0_outputs(3172) <= not(inputs(255));
    layer0_outputs(3173) <= inputs(180);
    layer0_outputs(3174) <= inputs(41);
    layer0_outputs(3175) <= not(inputs(220)) or (inputs(51));
    layer0_outputs(3176) <= (inputs(90)) or (inputs(92));
    layer0_outputs(3177) <= (inputs(145)) and not (inputs(64));
    layer0_outputs(3178) <= not(inputs(85)) or (inputs(235));
    layer0_outputs(3179) <= '0';
    layer0_outputs(3180) <= not((inputs(87)) or (inputs(198)));
    layer0_outputs(3181) <= (inputs(62)) xor (inputs(219));
    layer0_outputs(3182) <= inputs(75);
    layer0_outputs(3183) <= not(inputs(42));
    layer0_outputs(3184) <= (inputs(151)) and not (inputs(191));
    layer0_outputs(3185) <= inputs(131);
    layer0_outputs(3186) <= not((inputs(144)) or (inputs(38)));
    layer0_outputs(3187) <= (inputs(204)) xor (inputs(177));
    layer0_outputs(3188) <= (inputs(84)) or (inputs(51));
    layer0_outputs(3189) <= not((inputs(114)) or (inputs(106)));
    layer0_outputs(3190) <= not(inputs(98));
    layer0_outputs(3191) <= inputs(184);
    layer0_outputs(3192) <= not((inputs(123)) or (inputs(151)));
    layer0_outputs(3193) <= not((inputs(246)) xor (inputs(215)));
    layer0_outputs(3194) <= not(inputs(68));
    layer0_outputs(3195) <= inputs(198);
    layer0_outputs(3196) <= not(inputs(25));
    layer0_outputs(3197) <= (inputs(131)) or (inputs(154));
    layer0_outputs(3198) <= not((inputs(213)) xor (inputs(124)));
    layer0_outputs(3199) <= not((inputs(39)) xor (inputs(95)));
    layer0_outputs(3200) <= not((inputs(187)) xor (inputs(248)));
    layer0_outputs(3201) <= inputs(181);
    layer0_outputs(3202) <= (inputs(106)) and not (inputs(203));
    layer0_outputs(3203) <= not((inputs(20)) or (inputs(80)));
    layer0_outputs(3204) <= not(inputs(28)) or (inputs(191));
    layer0_outputs(3205) <= not(inputs(179));
    layer0_outputs(3206) <= (inputs(70)) and not (inputs(229));
    layer0_outputs(3207) <= (inputs(84)) xor (inputs(154));
    layer0_outputs(3208) <= (inputs(63)) or (inputs(13));
    layer0_outputs(3209) <= not((inputs(177)) xor (inputs(223)));
    layer0_outputs(3210) <= inputs(103);
    layer0_outputs(3211) <= not(inputs(8));
    layer0_outputs(3212) <= not(inputs(115));
    layer0_outputs(3213) <= '0';
    layer0_outputs(3214) <= not(inputs(70));
    layer0_outputs(3215) <= not(inputs(51)) or (inputs(1));
    layer0_outputs(3216) <= inputs(227);
    layer0_outputs(3217) <= not(inputs(12));
    layer0_outputs(3218) <= inputs(9);
    layer0_outputs(3219) <= inputs(81);
    layer0_outputs(3220) <= not(inputs(57));
    layer0_outputs(3221) <= not(inputs(105));
    layer0_outputs(3222) <= (inputs(145)) or (inputs(130));
    layer0_outputs(3223) <= not(inputs(68));
    layer0_outputs(3224) <= not((inputs(206)) xor (inputs(178)));
    layer0_outputs(3225) <= inputs(217);
    layer0_outputs(3226) <= not(inputs(100));
    layer0_outputs(3227) <= not(inputs(52)) or (inputs(206));
    layer0_outputs(3228) <= (inputs(63)) xor (inputs(65));
    layer0_outputs(3229) <= not(inputs(105));
    layer0_outputs(3230) <= (inputs(130)) or (inputs(123));
    layer0_outputs(3231) <= not((inputs(42)) or (inputs(35)));
    layer0_outputs(3232) <= not(inputs(169)) or (inputs(44));
    layer0_outputs(3233) <= inputs(58);
    layer0_outputs(3234) <= inputs(118);
    layer0_outputs(3235) <= not((inputs(152)) and (inputs(39)));
    layer0_outputs(3236) <= (inputs(139)) or (inputs(216));
    layer0_outputs(3237) <= not((inputs(198)) and (inputs(166)));
    layer0_outputs(3238) <= not(inputs(246));
    layer0_outputs(3239) <= not((inputs(80)) or (inputs(76)));
    layer0_outputs(3240) <= inputs(199);
    layer0_outputs(3241) <= not((inputs(98)) xor (inputs(10)));
    layer0_outputs(3242) <= inputs(8);
    layer0_outputs(3243) <= not((inputs(55)) or (inputs(31)));
    layer0_outputs(3244) <= (inputs(44)) and not (inputs(146));
    layer0_outputs(3245) <= not(inputs(241));
    layer0_outputs(3246) <= not(inputs(73));
    layer0_outputs(3247) <= not((inputs(100)) or (inputs(65)));
    layer0_outputs(3248) <= inputs(110);
    layer0_outputs(3249) <= not(inputs(26));
    layer0_outputs(3250) <= (inputs(94)) and (inputs(121));
    layer0_outputs(3251) <= not(inputs(100)) or (inputs(80));
    layer0_outputs(3252) <= (inputs(167)) and not (inputs(159));
    layer0_outputs(3253) <= (inputs(105)) or (inputs(58));
    layer0_outputs(3254) <= inputs(93);
    layer0_outputs(3255) <= inputs(82);
    layer0_outputs(3256) <= not(inputs(199));
    layer0_outputs(3257) <= not(inputs(233));
    layer0_outputs(3258) <= '0';
    layer0_outputs(3259) <= inputs(103);
    layer0_outputs(3260) <= (inputs(234)) or (inputs(218));
    layer0_outputs(3261) <= (inputs(106)) or (inputs(34));
    layer0_outputs(3262) <= (inputs(126)) xor (inputs(68));
    layer0_outputs(3263) <= not((inputs(10)) or (inputs(159)));
    layer0_outputs(3264) <= (inputs(74)) or (inputs(174));
    layer0_outputs(3265) <= (inputs(140)) and not (inputs(136));
    layer0_outputs(3266) <= (inputs(133)) and not (inputs(1));
    layer0_outputs(3267) <= inputs(183);
    layer0_outputs(3268) <= not((inputs(253)) or (inputs(226)));
    layer0_outputs(3269) <= inputs(231);
    layer0_outputs(3270) <= inputs(17);
    layer0_outputs(3271) <= (inputs(195)) and not (inputs(31));
    layer0_outputs(3272) <= inputs(135);
    layer0_outputs(3273) <= not((inputs(18)) xor (inputs(80)));
    layer0_outputs(3274) <= inputs(3);
    layer0_outputs(3275) <= not((inputs(138)) or (inputs(33)));
    layer0_outputs(3276) <= not(inputs(151)) or (inputs(190));
    layer0_outputs(3277) <= not(inputs(177)) or (inputs(15));
    layer0_outputs(3278) <= not(inputs(13));
    layer0_outputs(3279) <= (inputs(185)) xor (inputs(177));
    layer0_outputs(3280) <= (inputs(41)) and not (inputs(87));
    layer0_outputs(3281) <= not((inputs(60)) xor (inputs(14)));
    layer0_outputs(3282) <= (inputs(243)) or (inputs(206));
    layer0_outputs(3283) <= not((inputs(64)) and (inputs(247)));
    layer0_outputs(3284) <= (inputs(69)) and not (inputs(171));
    layer0_outputs(3285) <= inputs(113);
    layer0_outputs(3286) <= not(inputs(4)) or (inputs(174));
    layer0_outputs(3287) <= (inputs(114)) xor (inputs(68));
    layer0_outputs(3288) <= not((inputs(220)) xor (inputs(227)));
    layer0_outputs(3289) <= inputs(212);
    layer0_outputs(3290) <= (inputs(116)) or (inputs(102));
    layer0_outputs(3291) <= not((inputs(10)) or (inputs(230)));
    layer0_outputs(3292) <= (inputs(244)) and (inputs(177));
    layer0_outputs(3293) <= not((inputs(247)) xor (inputs(72)));
    layer0_outputs(3294) <= not(inputs(18)) or (inputs(97));
    layer0_outputs(3295) <= not(inputs(190));
    layer0_outputs(3296) <= (inputs(242)) xor (inputs(210));
    layer0_outputs(3297) <= not(inputs(230));
    layer0_outputs(3298) <= (inputs(36)) and not (inputs(175));
    layer0_outputs(3299) <= (inputs(25)) or (inputs(247));
    layer0_outputs(3300) <= not((inputs(46)) or (inputs(86)));
    layer0_outputs(3301) <= not(inputs(188));
    layer0_outputs(3302) <= not(inputs(159)) or (inputs(241));
    layer0_outputs(3303) <= inputs(238);
    layer0_outputs(3304) <= (inputs(74)) and not (inputs(88));
    layer0_outputs(3305) <= not((inputs(246)) or (inputs(227)));
    layer0_outputs(3306) <= not(inputs(225)) or (inputs(80));
    layer0_outputs(3307) <= '0';
    layer0_outputs(3308) <= (inputs(178)) xor (inputs(88));
    layer0_outputs(3309) <= not((inputs(82)) or (inputs(179)));
    layer0_outputs(3310) <= not(inputs(235));
    layer0_outputs(3311) <= not(inputs(98));
    layer0_outputs(3312) <= (inputs(221)) xor (inputs(158));
    layer0_outputs(3313) <= (inputs(172)) xor (inputs(221));
    layer0_outputs(3314) <= not((inputs(187)) or (inputs(101)));
    layer0_outputs(3315) <= not(inputs(237));
    layer0_outputs(3316) <= not(inputs(237));
    layer0_outputs(3317) <= not(inputs(69));
    layer0_outputs(3318) <= not(inputs(229)) or (inputs(49));
    layer0_outputs(3319) <= not(inputs(61)) or (inputs(224));
    layer0_outputs(3320) <= not(inputs(108)) or (inputs(2));
    layer0_outputs(3321) <= inputs(199);
    layer0_outputs(3322) <= not(inputs(218)) or (inputs(238));
    layer0_outputs(3323) <= (inputs(213)) or (inputs(67));
    layer0_outputs(3324) <= inputs(146);
    layer0_outputs(3325) <= not((inputs(102)) and (inputs(22)));
    layer0_outputs(3326) <= inputs(238);
    layer0_outputs(3327) <= (inputs(77)) and not (inputs(160));
    layer0_outputs(3328) <= not((inputs(139)) or (inputs(21)));
    layer0_outputs(3329) <= inputs(167);
    layer0_outputs(3330) <= (inputs(99)) and not (inputs(240));
    layer0_outputs(3331) <= not(inputs(84));
    layer0_outputs(3332) <= inputs(4);
    layer0_outputs(3333) <= inputs(195);
    layer0_outputs(3334) <= inputs(165);
    layer0_outputs(3335) <= not(inputs(57));
    layer0_outputs(3336) <= not(inputs(218));
    layer0_outputs(3337) <= (inputs(95)) and not (inputs(155));
    layer0_outputs(3338) <= not(inputs(83));
    layer0_outputs(3339) <= not((inputs(30)) or (inputs(220)));
    layer0_outputs(3340) <= (inputs(216)) and not (inputs(138));
    layer0_outputs(3341) <= inputs(54);
    layer0_outputs(3342) <= '1';
    layer0_outputs(3343) <= (inputs(20)) and (inputs(165));
    layer0_outputs(3344) <= (inputs(25)) xor (inputs(69));
    layer0_outputs(3345) <= not(inputs(187));
    layer0_outputs(3346) <= '0';
    layer0_outputs(3347) <= inputs(40);
    layer0_outputs(3348) <= not(inputs(152)) or (inputs(234));
    layer0_outputs(3349) <= not(inputs(212)) or (inputs(46));
    layer0_outputs(3350) <= inputs(64);
    layer0_outputs(3351) <= not(inputs(130));
    layer0_outputs(3352) <= not(inputs(151));
    layer0_outputs(3353) <= not(inputs(25));
    layer0_outputs(3354) <= not(inputs(197));
    layer0_outputs(3355) <= (inputs(101)) and not (inputs(18));
    layer0_outputs(3356) <= not((inputs(232)) xor (inputs(215)));
    layer0_outputs(3357) <= not(inputs(31));
    layer0_outputs(3358) <= not((inputs(164)) or (inputs(165)));
    layer0_outputs(3359) <= not((inputs(232)) or (inputs(206)));
    layer0_outputs(3360) <= (inputs(99)) and (inputs(129));
    layer0_outputs(3361) <= not((inputs(129)) xor (inputs(57)));
    layer0_outputs(3362) <= not(inputs(232));
    layer0_outputs(3363) <= (inputs(172)) and not (inputs(122));
    layer0_outputs(3364) <= inputs(179);
    layer0_outputs(3365) <= (inputs(130)) and not (inputs(152));
    layer0_outputs(3366) <= not((inputs(112)) or (inputs(77)));
    layer0_outputs(3367) <= (inputs(205)) and (inputs(61));
    layer0_outputs(3368) <= (inputs(3)) and (inputs(245));
    layer0_outputs(3369) <= not((inputs(211)) or (inputs(96)));
    layer0_outputs(3370) <= (inputs(148)) and not (inputs(17));
    layer0_outputs(3371) <= (inputs(35)) or (inputs(16));
    layer0_outputs(3372) <= (inputs(168)) and not (inputs(63));
    layer0_outputs(3373) <= not(inputs(165));
    layer0_outputs(3374) <= not(inputs(254)) or (inputs(216));
    layer0_outputs(3375) <= not((inputs(24)) or (inputs(79)));
    layer0_outputs(3376) <= (inputs(235)) or (inputs(194));
    layer0_outputs(3377) <= (inputs(73)) and (inputs(101));
    layer0_outputs(3378) <= not((inputs(187)) or (inputs(119)));
    layer0_outputs(3379) <= (inputs(52)) and not (inputs(235));
    layer0_outputs(3380) <= not(inputs(136)) or (inputs(206));
    layer0_outputs(3381) <= not(inputs(204)) or (inputs(112));
    layer0_outputs(3382) <= not(inputs(183));
    layer0_outputs(3383) <= (inputs(103)) and (inputs(234));
    layer0_outputs(3384) <= (inputs(134)) xor (inputs(145));
    layer0_outputs(3385) <= (inputs(119)) and not (inputs(207));
    layer0_outputs(3386) <= not(inputs(181));
    layer0_outputs(3387) <= not(inputs(57)) or (inputs(195));
    layer0_outputs(3388) <= inputs(159);
    layer0_outputs(3389) <= (inputs(194)) xor (inputs(104));
    layer0_outputs(3390) <= (inputs(231)) or (inputs(127));
    layer0_outputs(3391) <= '0';
    layer0_outputs(3392) <= (inputs(92)) xor (inputs(223));
    layer0_outputs(3393) <= (inputs(177)) xor (inputs(161));
    layer0_outputs(3394) <= not(inputs(137));
    layer0_outputs(3395) <= (inputs(56)) and (inputs(91));
    layer0_outputs(3396) <= inputs(48);
    layer0_outputs(3397) <= inputs(124);
    layer0_outputs(3398) <= inputs(74);
    layer0_outputs(3399) <= not((inputs(70)) xor (inputs(49)));
    layer0_outputs(3400) <= '1';
    layer0_outputs(3401) <= inputs(72);
    layer0_outputs(3402) <= (inputs(157)) xor (inputs(112));
    layer0_outputs(3403) <= not(inputs(120)) or (inputs(239));
    layer0_outputs(3404) <= (inputs(208)) or (inputs(116));
    layer0_outputs(3405) <= inputs(115);
    layer0_outputs(3406) <= inputs(192);
    layer0_outputs(3407) <= (inputs(100)) or (inputs(130));
    layer0_outputs(3408) <= not((inputs(163)) or (inputs(34)));
    layer0_outputs(3409) <= inputs(41);
    layer0_outputs(3410) <= not((inputs(179)) or (inputs(249)));
    layer0_outputs(3411) <= not(inputs(50));
    layer0_outputs(3412) <= not(inputs(84));
    layer0_outputs(3413) <= inputs(7);
    layer0_outputs(3414) <= not(inputs(75));
    layer0_outputs(3415) <= not((inputs(175)) or (inputs(203)));
    layer0_outputs(3416) <= inputs(182);
    layer0_outputs(3417) <= not(inputs(128));
    layer0_outputs(3418) <= inputs(114);
    layer0_outputs(3419) <= (inputs(9)) and not (inputs(247));
    layer0_outputs(3420) <= (inputs(11)) and not (inputs(200));
    layer0_outputs(3421) <= not(inputs(217)) or (inputs(46));
    layer0_outputs(3422) <= inputs(153);
    layer0_outputs(3423) <= (inputs(38)) and not (inputs(143));
    layer0_outputs(3424) <= not((inputs(23)) or (inputs(94)));
    layer0_outputs(3425) <= not((inputs(37)) or (inputs(51)));
    layer0_outputs(3426) <= inputs(104);
    layer0_outputs(3427) <= not(inputs(225));
    layer0_outputs(3428) <= not((inputs(110)) xor (inputs(204)));
    layer0_outputs(3429) <= inputs(178);
    layer0_outputs(3430) <= (inputs(116)) and not (inputs(108));
    layer0_outputs(3431) <= (inputs(7)) and not (inputs(175));
    layer0_outputs(3432) <= '1';
    layer0_outputs(3433) <= not((inputs(113)) or (inputs(52)));
    layer0_outputs(3434) <= not((inputs(136)) or (inputs(109)));
    layer0_outputs(3435) <= not(inputs(182));
    layer0_outputs(3436) <= not(inputs(45)) or (inputs(99));
    layer0_outputs(3437) <= not(inputs(189)) or (inputs(80));
    layer0_outputs(3438) <= not((inputs(134)) or (inputs(194)));
    layer0_outputs(3439) <= not(inputs(148)) or (inputs(237));
    layer0_outputs(3440) <= (inputs(12)) xor (inputs(209));
    layer0_outputs(3441) <= not(inputs(122));
    layer0_outputs(3442) <= (inputs(118)) and not (inputs(163));
    layer0_outputs(3443) <= '1';
    layer0_outputs(3444) <= not((inputs(211)) xor (inputs(105)));
    layer0_outputs(3445) <= not((inputs(205)) or (inputs(128)));
    layer0_outputs(3446) <= (inputs(253)) or (inputs(96));
    layer0_outputs(3447) <= (inputs(156)) xor (inputs(174));
    layer0_outputs(3448) <= not(inputs(130));
    layer0_outputs(3449) <= not(inputs(251)) or (inputs(0));
    layer0_outputs(3450) <= inputs(166);
    layer0_outputs(3451) <= (inputs(91)) xor (inputs(240));
    layer0_outputs(3452) <= inputs(183);
    layer0_outputs(3453) <= not(inputs(10)) or (inputs(159));
    layer0_outputs(3454) <= not(inputs(11)) or (inputs(24));
    layer0_outputs(3455) <= not((inputs(190)) or (inputs(87)));
    layer0_outputs(3456) <= not((inputs(189)) or (inputs(229)));
    layer0_outputs(3457) <= (inputs(185)) or (inputs(13));
    layer0_outputs(3458) <= inputs(121);
    layer0_outputs(3459) <= not(inputs(141)) or (inputs(252));
    layer0_outputs(3460) <= (inputs(213)) and not (inputs(142));
    layer0_outputs(3461) <= not((inputs(77)) xor (inputs(173)));
    layer0_outputs(3462) <= not((inputs(20)) or (inputs(196)));
    layer0_outputs(3463) <= (inputs(171)) xor (inputs(125));
    layer0_outputs(3464) <= (inputs(123)) or (inputs(22));
    layer0_outputs(3465) <= not(inputs(116));
    layer0_outputs(3466) <= (inputs(6)) and not (inputs(220));
    layer0_outputs(3467) <= not(inputs(84));
    layer0_outputs(3468) <= not(inputs(47)) or (inputs(240));
    layer0_outputs(3469) <= not((inputs(234)) xor (inputs(173)));
    layer0_outputs(3470) <= not((inputs(251)) xor (inputs(24)));
    layer0_outputs(3471) <= not((inputs(99)) or (inputs(185)));
    layer0_outputs(3472) <= not(inputs(163));
    layer0_outputs(3473) <= (inputs(134)) and not (inputs(220));
    layer0_outputs(3474) <= not(inputs(202)) or (inputs(70));
    layer0_outputs(3475) <= (inputs(219)) or (inputs(236));
    layer0_outputs(3476) <= (inputs(133)) xor (inputs(233));
    layer0_outputs(3477) <= not(inputs(24)) or (inputs(98));
    layer0_outputs(3478) <= not(inputs(56));
    layer0_outputs(3479) <= not(inputs(164));
    layer0_outputs(3480) <= not(inputs(215)) or (inputs(125));
    layer0_outputs(3481) <= (inputs(95)) or (inputs(102));
    layer0_outputs(3482) <= not((inputs(147)) or (inputs(224)));
    layer0_outputs(3483) <= (inputs(139)) and not (inputs(81));
    layer0_outputs(3484) <= not((inputs(33)) or (inputs(31)));
    layer0_outputs(3485) <= not(inputs(93));
    layer0_outputs(3486) <= inputs(179);
    layer0_outputs(3487) <= not(inputs(204));
    layer0_outputs(3488) <= (inputs(78)) or (inputs(23));
    layer0_outputs(3489) <= inputs(194);
    layer0_outputs(3490) <= not(inputs(40));
    layer0_outputs(3491) <= not(inputs(172));
    layer0_outputs(3492) <= inputs(100);
    layer0_outputs(3493) <= (inputs(19)) and not (inputs(87));
    layer0_outputs(3494) <= (inputs(89)) and not (inputs(220));
    layer0_outputs(3495) <= not(inputs(14));
    layer0_outputs(3496) <= (inputs(152)) and not (inputs(248));
    layer0_outputs(3497) <= not((inputs(237)) and (inputs(161)));
    layer0_outputs(3498) <= inputs(74);
    layer0_outputs(3499) <= inputs(101);
    layer0_outputs(3500) <= (inputs(211)) or (inputs(214));
    layer0_outputs(3501) <= not(inputs(181)) or (inputs(104));
    layer0_outputs(3502) <= not(inputs(103)) or (inputs(128));
    layer0_outputs(3503) <= not(inputs(235));
    layer0_outputs(3504) <= not((inputs(198)) and (inputs(37)));
    layer0_outputs(3505) <= not(inputs(235)) or (inputs(158));
    layer0_outputs(3506) <= inputs(157);
    layer0_outputs(3507) <= not(inputs(153)) or (inputs(234));
    layer0_outputs(3508) <= (inputs(16)) xor (inputs(181));
    layer0_outputs(3509) <= '0';
    layer0_outputs(3510) <= not((inputs(1)) or (inputs(76)));
    layer0_outputs(3511) <= not((inputs(154)) or (inputs(17)));
    layer0_outputs(3512) <= not((inputs(2)) and (inputs(147)));
    layer0_outputs(3513) <= not(inputs(198));
    layer0_outputs(3514) <= inputs(164);
    layer0_outputs(3515) <= not(inputs(180));
    layer0_outputs(3516) <= not(inputs(196));
    layer0_outputs(3517) <= (inputs(131)) or (inputs(127));
    layer0_outputs(3518) <= (inputs(190)) or (inputs(157));
    layer0_outputs(3519) <= not(inputs(82)) or (inputs(208));
    layer0_outputs(3520) <= not(inputs(111));
    layer0_outputs(3521) <= inputs(229);
    layer0_outputs(3522) <= not((inputs(191)) or (inputs(35)));
    layer0_outputs(3523) <= not(inputs(206)) or (inputs(254));
    layer0_outputs(3524) <= inputs(135);
    layer0_outputs(3525) <= (inputs(74)) and not (inputs(0));
    layer0_outputs(3526) <= inputs(103);
    layer0_outputs(3527) <= (inputs(119)) xor (inputs(13));
    layer0_outputs(3528) <= not(inputs(173));
    layer0_outputs(3529) <= (inputs(194)) xor (inputs(96));
    layer0_outputs(3530) <= not(inputs(61));
    layer0_outputs(3531) <= not(inputs(164));
    layer0_outputs(3532) <= (inputs(33)) or (inputs(38));
    layer0_outputs(3533) <= not(inputs(216));
    layer0_outputs(3534) <= (inputs(19)) and not (inputs(141));
    layer0_outputs(3535) <= not(inputs(31));
    layer0_outputs(3536) <= inputs(128);
    layer0_outputs(3537) <= (inputs(126)) or (inputs(20));
    layer0_outputs(3538) <= not((inputs(106)) or (inputs(243)));
    layer0_outputs(3539) <= not((inputs(87)) or (inputs(253)));
    layer0_outputs(3540) <= not((inputs(22)) xor (inputs(215)));
    layer0_outputs(3541) <= not(inputs(183));
    layer0_outputs(3542) <= not((inputs(160)) or (inputs(179)));
    layer0_outputs(3543) <= not((inputs(170)) or (inputs(253)));
    layer0_outputs(3544) <= not((inputs(246)) xor (inputs(233)));
    layer0_outputs(3545) <= not((inputs(159)) or (inputs(205)));
    layer0_outputs(3546) <= '1';
    layer0_outputs(3547) <= not((inputs(116)) xor (inputs(145)));
    layer0_outputs(3548) <= (inputs(123)) or (inputs(124));
    layer0_outputs(3549) <= not((inputs(128)) or (inputs(242)));
    layer0_outputs(3550) <= not(inputs(92));
    layer0_outputs(3551) <= not(inputs(237));
    layer0_outputs(3552) <= (inputs(133)) and not (inputs(179));
    layer0_outputs(3553) <= (inputs(213)) xor (inputs(135));
    layer0_outputs(3554) <= not(inputs(70));
    layer0_outputs(3555) <= not(inputs(73)) or (inputs(244));
    layer0_outputs(3556) <= not(inputs(84));
    layer0_outputs(3557) <= (inputs(138)) and not (inputs(9));
    layer0_outputs(3558) <= not(inputs(162)) or (inputs(78));
    layer0_outputs(3559) <= (inputs(67)) xor (inputs(81));
    layer0_outputs(3560) <= (inputs(139)) or (inputs(155));
    layer0_outputs(3561) <= not(inputs(229));
    layer0_outputs(3562) <= inputs(122);
    layer0_outputs(3563) <= not(inputs(208));
    layer0_outputs(3564) <= not(inputs(149));
    layer0_outputs(3565) <= (inputs(107)) and (inputs(5));
    layer0_outputs(3566) <= not(inputs(58));
    layer0_outputs(3567) <= inputs(105);
    layer0_outputs(3568) <= not((inputs(111)) xor (inputs(50)));
    layer0_outputs(3569) <= not((inputs(85)) xor (inputs(255)));
    layer0_outputs(3570) <= not((inputs(160)) xor (inputs(133)));
    layer0_outputs(3571) <= not((inputs(6)) or (inputs(181)));
    layer0_outputs(3572) <= (inputs(139)) and not (inputs(182));
    layer0_outputs(3573) <= not((inputs(209)) xor (inputs(72)));
    layer0_outputs(3574) <= (inputs(238)) and not (inputs(172));
    layer0_outputs(3575) <= not(inputs(173)) or (inputs(48));
    layer0_outputs(3576) <= (inputs(2)) or (inputs(210));
    layer0_outputs(3577) <= not((inputs(197)) and (inputs(199)));
    layer0_outputs(3578) <= not(inputs(190)) or (inputs(98));
    layer0_outputs(3579) <= inputs(7);
    layer0_outputs(3580) <= (inputs(112)) or (inputs(147));
    layer0_outputs(3581) <= not((inputs(252)) or (inputs(116)));
    layer0_outputs(3582) <= inputs(92);
    layer0_outputs(3583) <= (inputs(61)) or (inputs(93));
    layer0_outputs(3584) <= (inputs(38)) and (inputs(138));
    layer0_outputs(3585) <= (inputs(2)) and not (inputs(29));
    layer0_outputs(3586) <= (inputs(124)) and (inputs(36));
    layer0_outputs(3587) <= (inputs(195)) or (inputs(91));
    layer0_outputs(3588) <= not(inputs(113)) or (inputs(192));
    layer0_outputs(3589) <= inputs(115);
    layer0_outputs(3590) <= (inputs(148)) xor (inputs(161));
    layer0_outputs(3591) <= not(inputs(157));
    layer0_outputs(3592) <= not(inputs(131));
    layer0_outputs(3593) <= inputs(114);
    layer0_outputs(3594) <= (inputs(99)) and not (inputs(207));
    layer0_outputs(3595) <= '0';
    layer0_outputs(3596) <= inputs(98);
    layer0_outputs(3597) <= inputs(125);
    layer0_outputs(3598) <= (inputs(98)) xor (inputs(255));
    layer0_outputs(3599) <= not(inputs(228));
    layer0_outputs(3600) <= not(inputs(86));
    layer0_outputs(3601) <= (inputs(79)) and not (inputs(247));
    layer0_outputs(3602) <= (inputs(249)) or (inputs(10));
    layer0_outputs(3603) <= not((inputs(168)) or (inputs(254)));
    layer0_outputs(3604) <= (inputs(192)) or (inputs(46));
    layer0_outputs(3605) <= (inputs(202)) or (inputs(209));
    layer0_outputs(3606) <= not(inputs(47)) or (inputs(99));
    layer0_outputs(3607) <= not(inputs(210));
    layer0_outputs(3608) <= inputs(48);
    layer0_outputs(3609) <= not((inputs(42)) and (inputs(49)));
    layer0_outputs(3610) <= not(inputs(168)) or (inputs(0));
    layer0_outputs(3611) <= not(inputs(210));
    layer0_outputs(3612) <= not(inputs(212));
    layer0_outputs(3613) <= inputs(23);
    layer0_outputs(3614) <= inputs(113);
    layer0_outputs(3615) <= (inputs(191)) or (inputs(18));
    layer0_outputs(3616) <= (inputs(137)) or (inputs(46));
    layer0_outputs(3617) <= not(inputs(254)) or (inputs(106));
    layer0_outputs(3618) <= not(inputs(27)) or (inputs(175));
    layer0_outputs(3619) <= (inputs(189)) and not (inputs(234));
    layer0_outputs(3620) <= not(inputs(99));
    layer0_outputs(3621) <= not((inputs(191)) or (inputs(57)));
    layer0_outputs(3622) <= not(inputs(85));
    layer0_outputs(3623) <= (inputs(43)) or (inputs(42));
    layer0_outputs(3624) <= not(inputs(204)) or (inputs(224));
    layer0_outputs(3625) <= inputs(73);
    layer0_outputs(3626) <= (inputs(138)) and not (inputs(174));
    layer0_outputs(3627) <= (inputs(115)) and not (inputs(56));
    layer0_outputs(3628) <= not((inputs(162)) xor (inputs(8)));
    layer0_outputs(3629) <= not((inputs(65)) or (inputs(162)));
    layer0_outputs(3630) <= not(inputs(122)) or (inputs(86));
    layer0_outputs(3631) <= not((inputs(204)) or (inputs(222)));
    layer0_outputs(3632) <= '0';
    layer0_outputs(3633) <= not((inputs(179)) xor (inputs(250)));
    layer0_outputs(3634) <= not(inputs(124)) or (inputs(163));
    layer0_outputs(3635) <= (inputs(36)) xor (inputs(124));
    layer0_outputs(3636) <= not(inputs(213)) or (inputs(224));
    layer0_outputs(3637) <= not(inputs(158)) or (inputs(49));
    layer0_outputs(3638) <= (inputs(240)) and not (inputs(16));
    layer0_outputs(3639) <= (inputs(227)) and not (inputs(189));
    layer0_outputs(3640) <= not(inputs(245));
    layer0_outputs(3641) <= not((inputs(213)) or (inputs(97)));
    layer0_outputs(3642) <= (inputs(20)) or (inputs(9));
    layer0_outputs(3643) <= not(inputs(137));
    layer0_outputs(3644) <= not(inputs(169)) or (inputs(132));
    layer0_outputs(3645) <= not(inputs(124)) or (inputs(241));
    layer0_outputs(3646) <= not((inputs(193)) or (inputs(217)));
    layer0_outputs(3647) <= not(inputs(170)) or (inputs(104));
    layer0_outputs(3648) <= (inputs(6)) and not (inputs(205));
    layer0_outputs(3649) <= not((inputs(151)) xor (inputs(176)));
    layer0_outputs(3650) <= inputs(23);
    layer0_outputs(3651) <= not((inputs(202)) or (inputs(110)));
    layer0_outputs(3652) <= not((inputs(198)) or (inputs(150)));
    layer0_outputs(3653) <= inputs(105);
    layer0_outputs(3654) <= inputs(60);
    layer0_outputs(3655) <= not((inputs(111)) or (inputs(137)));
    layer0_outputs(3656) <= (inputs(172)) xor (inputs(170));
    layer0_outputs(3657) <= (inputs(34)) xor (inputs(171));
    layer0_outputs(3658) <= not(inputs(137));
    layer0_outputs(3659) <= (inputs(112)) and not (inputs(222));
    layer0_outputs(3660) <= not((inputs(37)) or (inputs(144)));
    layer0_outputs(3661) <= (inputs(71)) and not (inputs(34));
    layer0_outputs(3662) <= (inputs(207)) and not (inputs(15));
    layer0_outputs(3663) <= not(inputs(195)) or (inputs(115));
    layer0_outputs(3664) <= not(inputs(161));
    layer0_outputs(3665) <= (inputs(148)) and not (inputs(225));
    layer0_outputs(3666) <= (inputs(190)) or (inputs(32));
    layer0_outputs(3667) <= (inputs(58)) and not (inputs(95));
    layer0_outputs(3668) <= (inputs(239)) or (inputs(115));
    layer0_outputs(3669) <= not(inputs(187)) or (inputs(28));
    layer0_outputs(3670) <= not((inputs(236)) or (inputs(235)));
    layer0_outputs(3671) <= inputs(47);
    layer0_outputs(3672) <= inputs(17);
    layer0_outputs(3673) <= not((inputs(48)) or (inputs(34)));
    layer0_outputs(3674) <= inputs(7);
    layer0_outputs(3675) <= (inputs(202)) or (inputs(143));
    layer0_outputs(3676) <= inputs(197);
    layer0_outputs(3677) <= (inputs(30)) xor (inputs(1));
    layer0_outputs(3678) <= not(inputs(166));
    layer0_outputs(3679) <= '0';
    layer0_outputs(3680) <= inputs(54);
    layer0_outputs(3681) <= (inputs(124)) or (inputs(180));
    layer0_outputs(3682) <= inputs(220);
    layer0_outputs(3683) <= (inputs(70)) or (inputs(237));
    layer0_outputs(3684) <= not(inputs(190));
    layer0_outputs(3685) <= inputs(241);
    layer0_outputs(3686) <= not(inputs(70)) or (inputs(81));
    layer0_outputs(3687) <= (inputs(110)) or (inputs(169));
    layer0_outputs(3688) <= (inputs(195)) or (inputs(127));
    layer0_outputs(3689) <= not(inputs(191));
    layer0_outputs(3690) <= inputs(114);
    layer0_outputs(3691) <= (inputs(102)) and not (inputs(72));
    layer0_outputs(3692) <= not((inputs(119)) xor (inputs(197)));
    layer0_outputs(3693) <= inputs(24);
    layer0_outputs(3694) <= inputs(12);
    layer0_outputs(3695) <= not(inputs(159));
    layer0_outputs(3696) <= inputs(124);
    layer0_outputs(3697) <= '0';
    layer0_outputs(3698) <= inputs(80);
    layer0_outputs(3699) <= not(inputs(218)) or (inputs(73));
    layer0_outputs(3700) <= not(inputs(10));
    layer0_outputs(3701) <= (inputs(100)) and not (inputs(178));
    layer0_outputs(3702) <= (inputs(204)) and not (inputs(28));
    layer0_outputs(3703) <= (inputs(48)) and not (inputs(96));
    layer0_outputs(3704) <= inputs(105);
    layer0_outputs(3705) <= inputs(232);
    layer0_outputs(3706) <= (inputs(62)) or (inputs(42));
    layer0_outputs(3707) <= inputs(106);
    layer0_outputs(3708) <= (inputs(98)) or (inputs(122));
    layer0_outputs(3709) <= not(inputs(70));
    layer0_outputs(3710) <= (inputs(44)) or (inputs(144));
    layer0_outputs(3711) <= (inputs(137)) xor (inputs(188));
    layer0_outputs(3712) <= not(inputs(77));
    layer0_outputs(3713) <= (inputs(85)) and not (inputs(175));
    layer0_outputs(3714) <= not(inputs(70)) or (inputs(63));
    layer0_outputs(3715) <= inputs(71);
    layer0_outputs(3716) <= (inputs(218)) xor (inputs(37));
    layer0_outputs(3717) <= inputs(45);
    layer0_outputs(3718) <= not((inputs(68)) or (inputs(102)));
    layer0_outputs(3719) <= inputs(206);
    layer0_outputs(3720) <= not((inputs(148)) or (inputs(245)));
    layer0_outputs(3721) <= not(inputs(215));
    layer0_outputs(3722) <= (inputs(156)) xor (inputs(244));
    layer0_outputs(3723) <= inputs(118);
    layer0_outputs(3724) <= not(inputs(131));
    layer0_outputs(3725) <= (inputs(127)) xor (inputs(1));
    layer0_outputs(3726) <= not((inputs(179)) xor (inputs(177)));
    layer0_outputs(3727) <= not(inputs(228));
    layer0_outputs(3728) <= (inputs(42)) and (inputs(40));
    layer0_outputs(3729) <= (inputs(218)) or (inputs(207));
    layer0_outputs(3730) <= not(inputs(64)) or (inputs(238));
    layer0_outputs(3731) <= not(inputs(120));
    layer0_outputs(3732) <= not((inputs(45)) or (inputs(241)));
    layer0_outputs(3733) <= inputs(135);
    layer0_outputs(3734) <= not(inputs(61)) or (inputs(48));
    layer0_outputs(3735) <= inputs(22);
    layer0_outputs(3736) <= not(inputs(84)) or (inputs(53));
    layer0_outputs(3737) <= (inputs(192)) or (inputs(203));
    layer0_outputs(3738) <= (inputs(138)) xor (inputs(11));
    layer0_outputs(3739) <= inputs(161);
    layer0_outputs(3740) <= not((inputs(39)) or (inputs(18)));
    layer0_outputs(3741) <= '0';
    layer0_outputs(3742) <= not(inputs(241)) or (inputs(226));
    layer0_outputs(3743) <= not((inputs(49)) xor (inputs(59)));
    layer0_outputs(3744) <= not(inputs(229)) or (inputs(255));
    layer0_outputs(3745) <= not(inputs(105)) or (inputs(1));
    layer0_outputs(3746) <= (inputs(15)) and not (inputs(192));
    layer0_outputs(3747) <= not(inputs(217)) or (inputs(34));
    layer0_outputs(3748) <= not((inputs(201)) or (inputs(34)));
    layer0_outputs(3749) <= (inputs(8)) or (inputs(49));
    layer0_outputs(3750) <= not(inputs(62)) or (inputs(135));
    layer0_outputs(3751) <= (inputs(176)) and not (inputs(34));
    layer0_outputs(3752) <= (inputs(173)) xor (inputs(31));
    layer0_outputs(3753) <= not(inputs(105));
    layer0_outputs(3754) <= (inputs(198)) xor (inputs(51));
    layer0_outputs(3755) <= not(inputs(77)) or (inputs(51));
    layer0_outputs(3756) <= not(inputs(70)) or (inputs(36));
    layer0_outputs(3757) <= not((inputs(154)) or (inputs(95)));
    layer0_outputs(3758) <= not(inputs(96));
    layer0_outputs(3759) <= (inputs(151)) or (inputs(207));
    layer0_outputs(3760) <= (inputs(174)) or (inputs(197));
    layer0_outputs(3761) <= not(inputs(172)) or (inputs(240));
    layer0_outputs(3762) <= not(inputs(24)) or (inputs(130));
    layer0_outputs(3763) <= inputs(161);
    layer0_outputs(3764) <= not(inputs(111));
    layer0_outputs(3765) <= (inputs(254)) and not (inputs(113));
    layer0_outputs(3766) <= inputs(156);
    layer0_outputs(3767) <= not(inputs(184)) or (inputs(155));
    layer0_outputs(3768) <= inputs(25);
    layer0_outputs(3769) <= not((inputs(19)) xor (inputs(237)));
    layer0_outputs(3770) <= not(inputs(86));
    layer0_outputs(3771) <= not((inputs(18)) or (inputs(186)));
    layer0_outputs(3772) <= not(inputs(69));
    layer0_outputs(3773) <= (inputs(251)) xor (inputs(171));
    layer0_outputs(3774) <= (inputs(90)) or (inputs(73));
    layer0_outputs(3775) <= inputs(119);
    layer0_outputs(3776) <= (inputs(171)) or (inputs(214));
    layer0_outputs(3777) <= (inputs(23)) and not (inputs(124));
    layer0_outputs(3778) <= (inputs(40)) and not (inputs(145));
    layer0_outputs(3779) <= (inputs(35)) and not (inputs(74));
    layer0_outputs(3780) <= (inputs(16)) and not (inputs(83));
    layer0_outputs(3781) <= (inputs(193)) or (inputs(173));
    layer0_outputs(3782) <= (inputs(84)) and not (inputs(176));
    layer0_outputs(3783) <= '0';
    layer0_outputs(3784) <= not((inputs(137)) or (inputs(114)));
    layer0_outputs(3785) <= not((inputs(20)) and (inputs(196)));
    layer0_outputs(3786) <= inputs(208);
    layer0_outputs(3787) <= (inputs(167)) and not (inputs(37));
    layer0_outputs(3788) <= not(inputs(26)) or (inputs(163));
    layer0_outputs(3789) <= not(inputs(226));
    layer0_outputs(3790) <= (inputs(133)) and not (inputs(15));
    layer0_outputs(3791) <= (inputs(156)) or (inputs(46));
    layer0_outputs(3792) <= not(inputs(140));
    layer0_outputs(3793) <= inputs(246);
    layer0_outputs(3794) <= not((inputs(161)) or (inputs(70)));
    layer0_outputs(3795) <= not((inputs(84)) or (inputs(166)));
    layer0_outputs(3796) <= (inputs(27)) and not (inputs(204));
    layer0_outputs(3797) <= (inputs(200)) and (inputs(239));
    layer0_outputs(3798) <= (inputs(88)) and not (inputs(250));
    layer0_outputs(3799) <= not(inputs(164));
    layer0_outputs(3800) <= (inputs(128)) or (inputs(15));
    layer0_outputs(3801) <= not(inputs(90));
    layer0_outputs(3802) <= (inputs(154)) or (inputs(52));
    layer0_outputs(3803) <= inputs(136);
    layer0_outputs(3804) <= not(inputs(22)) or (inputs(250));
    layer0_outputs(3805) <= not(inputs(155)) or (inputs(111));
    layer0_outputs(3806) <= (inputs(242)) or (inputs(222));
    layer0_outputs(3807) <= not((inputs(216)) or (inputs(144)));
    layer0_outputs(3808) <= not(inputs(114));
    layer0_outputs(3809) <= (inputs(78)) or (inputs(115));
    layer0_outputs(3810) <= not(inputs(46));
    layer0_outputs(3811) <= (inputs(251)) or (inputs(150));
    layer0_outputs(3812) <= (inputs(49)) and not (inputs(255));
    layer0_outputs(3813) <= inputs(105);
    layer0_outputs(3814) <= (inputs(83)) or (inputs(239));
    layer0_outputs(3815) <= not((inputs(249)) or (inputs(211)));
    layer0_outputs(3816) <= not((inputs(191)) xor (inputs(237)));
    layer0_outputs(3817) <= (inputs(46)) or (inputs(103));
    layer0_outputs(3818) <= not(inputs(199));
    layer0_outputs(3819) <= not(inputs(64));
    layer0_outputs(3820) <= (inputs(153)) and not (inputs(8));
    layer0_outputs(3821) <= (inputs(40)) or (inputs(87));
    layer0_outputs(3822) <= (inputs(211)) or (inputs(221));
    layer0_outputs(3823) <= (inputs(106)) and not (inputs(209));
    layer0_outputs(3824) <= not(inputs(197));
    layer0_outputs(3825) <= inputs(213);
    layer0_outputs(3826) <= not(inputs(59));
    layer0_outputs(3827) <= not((inputs(112)) or (inputs(110)));
    layer0_outputs(3828) <= not(inputs(103));
    layer0_outputs(3829) <= not(inputs(167)) or (inputs(117));
    layer0_outputs(3830) <= (inputs(188)) or (inputs(160));
    layer0_outputs(3831) <= not(inputs(86));
    layer0_outputs(3832) <= inputs(134);
    layer0_outputs(3833) <= not(inputs(212));
    layer0_outputs(3834) <= '1';
    layer0_outputs(3835) <= (inputs(25)) and not (inputs(203));
    layer0_outputs(3836) <= not(inputs(92));
    layer0_outputs(3837) <= (inputs(156)) or (inputs(111));
    layer0_outputs(3838) <= not(inputs(24)) or (inputs(241));
    layer0_outputs(3839) <= not((inputs(1)) xor (inputs(208)));
    layer0_outputs(3840) <= not(inputs(219));
    layer0_outputs(3841) <= '0';
    layer0_outputs(3842) <= not(inputs(136));
    layer0_outputs(3843) <= not((inputs(123)) or (inputs(19)));
    layer0_outputs(3844) <= not((inputs(197)) xor (inputs(244)));
    layer0_outputs(3845) <= not((inputs(249)) xor (inputs(50)));
    layer0_outputs(3846) <= not((inputs(143)) or (inputs(85)));
    layer0_outputs(3847) <= '1';
    layer0_outputs(3848) <= not(inputs(104));
    layer0_outputs(3849) <= not(inputs(165));
    layer0_outputs(3850) <= not(inputs(90));
    layer0_outputs(3851) <= inputs(76);
    layer0_outputs(3852) <= not(inputs(158));
    layer0_outputs(3853) <= (inputs(178)) xor (inputs(248));
    layer0_outputs(3854) <= not(inputs(191));
    layer0_outputs(3855) <= (inputs(195)) and not (inputs(195));
    layer0_outputs(3856) <= (inputs(63)) and (inputs(38));
    layer0_outputs(3857) <= (inputs(22)) xor (inputs(13));
    layer0_outputs(3858) <= not(inputs(153)) or (inputs(111));
    layer0_outputs(3859) <= inputs(81);
    layer0_outputs(3860) <= not((inputs(206)) or (inputs(190)));
    layer0_outputs(3861) <= not(inputs(212)) or (inputs(16));
    layer0_outputs(3862) <= not(inputs(167));
    layer0_outputs(3863) <= '0';
    layer0_outputs(3864) <= inputs(101);
    layer0_outputs(3865) <= inputs(232);
    layer0_outputs(3866) <= not((inputs(75)) or (inputs(184)));
    layer0_outputs(3867) <= not(inputs(100));
    layer0_outputs(3868) <= not((inputs(83)) xor (inputs(116)));
    layer0_outputs(3869) <= '0';
    layer0_outputs(3870) <= not(inputs(179));
    layer0_outputs(3871) <= (inputs(252)) xor (inputs(226));
    layer0_outputs(3872) <= not(inputs(178)) or (inputs(48));
    layer0_outputs(3873) <= inputs(225);
    layer0_outputs(3874) <= not((inputs(156)) or (inputs(192)));
    layer0_outputs(3875) <= (inputs(149)) or (inputs(252));
    layer0_outputs(3876) <= (inputs(205)) xor (inputs(141));
    layer0_outputs(3877) <= not(inputs(179));
    layer0_outputs(3878) <= (inputs(10)) and (inputs(240));
    layer0_outputs(3879) <= not((inputs(88)) xor (inputs(75)));
    layer0_outputs(3880) <= inputs(113);
    layer0_outputs(3881) <= inputs(148);
    layer0_outputs(3882) <= (inputs(229)) xor (inputs(25));
    layer0_outputs(3883) <= not(inputs(98));
    layer0_outputs(3884) <= not((inputs(92)) xor (inputs(48)));
    layer0_outputs(3885) <= not(inputs(163)) or (inputs(31));
    layer0_outputs(3886) <= not(inputs(249)) or (inputs(207));
    layer0_outputs(3887) <= inputs(28);
    layer0_outputs(3888) <= (inputs(29)) xor (inputs(55));
    layer0_outputs(3889) <= '1';
    layer0_outputs(3890) <= not(inputs(163));
    layer0_outputs(3891) <= not(inputs(68)) or (inputs(210));
    layer0_outputs(3892) <= not(inputs(209));
    layer0_outputs(3893) <= not(inputs(45)) or (inputs(146));
    layer0_outputs(3894) <= not(inputs(104));
    layer0_outputs(3895) <= not((inputs(207)) or (inputs(25)));
    layer0_outputs(3896) <= inputs(105);
    layer0_outputs(3897) <= (inputs(144)) xor (inputs(132));
    layer0_outputs(3898) <= (inputs(54)) and (inputs(57));
    layer0_outputs(3899) <= (inputs(174)) xor (inputs(23));
    layer0_outputs(3900) <= (inputs(242)) and (inputs(17));
    layer0_outputs(3901) <= (inputs(30)) xor (inputs(0));
    layer0_outputs(3902) <= (inputs(70)) or (inputs(227));
    layer0_outputs(3903) <= not((inputs(195)) xor (inputs(88)));
    layer0_outputs(3904) <= (inputs(87)) or (inputs(218));
    layer0_outputs(3905) <= not(inputs(26)) or (inputs(173));
    layer0_outputs(3906) <= not(inputs(93));
    layer0_outputs(3907) <= not(inputs(100)) or (inputs(112));
    layer0_outputs(3908) <= (inputs(230)) and not (inputs(92));
    layer0_outputs(3909) <= not((inputs(220)) or (inputs(51)));
    layer0_outputs(3910) <= (inputs(241)) or (inputs(45));
    layer0_outputs(3911) <= not((inputs(201)) and (inputs(40)));
    layer0_outputs(3912) <= (inputs(49)) and not (inputs(14));
    layer0_outputs(3913) <= not(inputs(141));
    layer0_outputs(3914) <= not(inputs(25));
    layer0_outputs(3915) <= inputs(110);
    layer0_outputs(3916) <= not(inputs(194)) or (inputs(146));
    layer0_outputs(3917) <= inputs(34);
    layer0_outputs(3918) <= not(inputs(142)) or (inputs(177));
    layer0_outputs(3919) <= not(inputs(56));
    layer0_outputs(3920) <= not(inputs(214));
    layer0_outputs(3921) <= not(inputs(120)) or (inputs(207));
    layer0_outputs(3922) <= (inputs(50)) or (inputs(176));
    layer0_outputs(3923) <= not(inputs(239)) or (inputs(207));
    layer0_outputs(3924) <= (inputs(214)) and not (inputs(66));
    layer0_outputs(3925) <= (inputs(75)) or (inputs(88));
    layer0_outputs(3926) <= (inputs(237)) or (inputs(199));
    layer0_outputs(3927) <= (inputs(195)) xor (inputs(176));
    layer0_outputs(3928) <= not(inputs(247));
    layer0_outputs(3929) <= not(inputs(94));
    layer0_outputs(3930) <= not(inputs(106));
    layer0_outputs(3931) <= not(inputs(12)) or (inputs(161));
    layer0_outputs(3932) <= (inputs(5)) or (inputs(141));
    layer0_outputs(3933) <= (inputs(215)) and not (inputs(250));
    layer0_outputs(3934) <= not(inputs(186)) or (inputs(217));
    layer0_outputs(3935) <= (inputs(70)) and not (inputs(99));
    layer0_outputs(3936) <= not((inputs(150)) or (inputs(32)));
    layer0_outputs(3937) <= (inputs(230)) and not (inputs(242));
    layer0_outputs(3938) <= not((inputs(0)) xor (inputs(81)));
    layer0_outputs(3939) <= (inputs(111)) xor (inputs(155));
    layer0_outputs(3940) <= not(inputs(131));
    layer0_outputs(3941) <= not(inputs(27)) or (inputs(225));
    layer0_outputs(3942) <= inputs(107);
    layer0_outputs(3943) <= '0';
    layer0_outputs(3944) <= (inputs(78)) xor (inputs(220));
    layer0_outputs(3945) <= not(inputs(101));
    layer0_outputs(3946) <= (inputs(219)) or (inputs(59));
    layer0_outputs(3947) <= inputs(22);
    layer0_outputs(3948) <= (inputs(251)) and not (inputs(131));
    layer0_outputs(3949) <= (inputs(184)) and not (inputs(209));
    layer0_outputs(3950) <= not(inputs(40));
    layer0_outputs(3951) <= not((inputs(15)) or (inputs(153)));
    layer0_outputs(3952) <= (inputs(230)) xor (inputs(24));
    layer0_outputs(3953) <= not(inputs(55));
    layer0_outputs(3954) <= not((inputs(223)) xor (inputs(133)));
    layer0_outputs(3955) <= not((inputs(143)) or (inputs(138)));
    layer0_outputs(3956) <= inputs(200);
    layer0_outputs(3957) <= (inputs(206)) xor (inputs(155));
    layer0_outputs(3958) <= (inputs(26)) or (inputs(66));
    layer0_outputs(3959) <= (inputs(122)) xor (inputs(240));
    layer0_outputs(3960) <= (inputs(25)) and (inputs(136));
    layer0_outputs(3961) <= (inputs(58)) and not (inputs(208));
    layer0_outputs(3962) <= not(inputs(143));
    layer0_outputs(3963) <= (inputs(73)) xor (inputs(22));
    layer0_outputs(3964) <= not((inputs(154)) or (inputs(129)));
    layer0_outputs(3965) <= (inputs(167)) and not (inputs(143));
    layer0_outputs(3966) <= not((inputs(16)) xor (inputs(176)));
    layer0_outputs(3967) <= not((inputs(188)) and (inputs(99)));
    layer0_outputs(3968) <= inputs(156);
    layer0_outputs(3969) <= not((inputs(199)) and (inputs(203)));
    layer0_outputs(3970) <= inputs(69);
    layer0_outputs(3971) <= not(inputs(83));
    layer0_outputs(3972) <= not(inputs(105));
    layer0_outputs(3973) <= not((inputs(27)) or (inputs(230)));
    layer0_outputs(3974) <= not((inputs(170)) or (inputs(100)));
    layer0_outputs(3975) <= not((inputs(132)) xor (inputs(183)));
    layer0_outputs(3976) <= inputs(113);
    layer0_outputs(3977) <= (inputs(104)) and not (inputs(84));
    layer0_outputs(3978) <= not(inputs(91)) or (inputs(250));
    layer0_outputs(3979) <= not(inputs(197));
    layer0_outputs(3980) <= (inputs(255)) or (inputs(124));
    layer0_outputs(3981) <= inputs(236);
    layer0_outputs(3982) <= (inputs(109)) xor (inputs(19));
    layer0_outputs(3983) <= (inputs(112)) and not (inputs(69));
    layer0_outputs(3984) <= (inputs(231)) and not (inputs(154));
    layer0_outputs(3985) <= not((inputs(121)) xor (inputs(33)));
    layer0_outputs(3986) <= (inputs(66)) or (inputs(242));
    layer0_outputs(3987) <= (inputs(166)) or (inputs(186));
    layer0_outputs(3988) <= not((inputs(59)) or (inputs(96)));
    layer0_outputs(3989) <= not(inputs(115));
    layer0_outputs(3990) <= '1';
    layer0_outputs(3991) <= (inputs(181)) or (inputs(69));
    layer0_outputs(3992) <= inputs(2);
    layer0_outputs(3993) <= (inputs(133)) and not (inputs(32));
    layer0_outputs(3994) <= not(inputs(166));
    layer0_outputs(3995) <= not((inputs(144)) or (inputs(100)));
    layer0_outputs(3996) <= (inputs(23)) or (inputs(240));
    layer0_outputs(3997) <= (inputs(81)) and not (inputs(81));
    layer0_outputs(3998) <= not(inputs(162));
    layer0_outputs(3999) <= (inputs(121)) and not (inputs(78));
    layer0_outputs(4000) <= (inputs(233)) or (inputs(3));
    layer0_outputs(4001) <= not((inputs(118)) xor (inputs(103)));
    layer0_outputs(4002) <= not(inputs(131));
    layer0_outputs(4003) <= not((inputs(108)) or (inputs(104)));
    layer0_outputs(4004) <= not((inputs(171)) xor (inputs(6)));
    layer0_outputs(4005) <= inputs(211);
    layer0_outputs(4006) <= not(inputs(201));
    layer0_outputs(4007) <= not(inputs(25));
    layer0_outputs(4008) <= not(inputs(1)) or (inputs(95));
    layer0_outputs(4009) <= inputs(189);
    layer0_outputs(4010) <= not(inputs(158));
    layer0_outputs(4011) <= (inputs(208)) or (inputs(173));
    layer0_outputs(4012) <= not(inputs(231));
    layer0_outputs(4013) <= not((inputs(144)) xor (inputs(39)));
    layer0_outputs(4014) <= inputs(120);
    layer0_outputs(4015) <= (inputs(236)) and not (inputs(150));
    layer0_outputs(4016) <= not(inputs(15));
    layer0_outputs(4017) <= not(inputs(200)) or (inputs(177));
    layer0_outputs(4018) <= inputs(183);
    layer0_outputs(4019) <= not((inputs(156)) or (inputs(207)));
    layer0_outputs(4020) <= not(inputs(170));
    layer0_outputs(4021) <= (inputs(53)) and not (inputs(190));
    layer0_outputs(4022) <= (inputs(31)) and not (inputs(53));
    layer0_outputs(4023) <= inputs(182);
    layer0_outputs(4024) <= not(inputs(74)) or (inputs(224));
    layer0_outputs(4025) <= inputs(212);
    layer0_outputs(4026) <= not(inputs(143));
    layer0_outputs(4027) <= inputs(44);
    layer0_outputs(4028) <= (inputs(2)) xor (inputs(206));
    layer0_outputs(4029) <= inputs(81);
    layer0_outputs(4030) <= '0';
    layer0_outputs(4031) <= not(inputs(200)) or (inputs(118));
    layer0_outputs(4032) <= (inputs(191)) xor (inputs(28));
    layer0_outputs(4033) <= (inputs(123)) xor (inputs(65));
    layer0_outputs(4034) <= not((inputs(83)) or (inputs(146)));
    layer0_outputs(4035) <= inputs(66);
    layer0_outputs(4036) <= not(inputs(241));
    layer0_outputs(4037) <= not(inputs(110));
    layer0_outputs(4038) <= inputs(28);
    layer0_outputs(4039) <= inputs(230);
    layer0_outputs(4040) <= inputs(103);
    layer0_outputs(4041) <= not(inputs(119));
    layer0_outputs(4042) <= inputs(166);
    layer0_outputs(4043) <= inputs(102);
    layer0_outputs(4044) <= not(inputs(25)) or (inputs(239));
    layer0_outputs(4045) <= not((inputs(208)) or (inputs(173)));
    layer0_outputs(4046) <= not((inputs(219)) xor (inputs(24)));
    layer0_outputs(4047) <= not((inputs(153)) xor (inputs(136)));
    layer0_outputs(4048) <= not(inputs(29));
    layer0_outputs(4049) <= not(inputs(23)) or (inputs(0));
    layer0_outputs(4050) <= not((inputs(216)) or (inputs(33)));
    layer0_outputs(4051) <= (inputs(228)) and (inputs(57));
    layer0_outputs(4052) <= not((inputs(182)) or (inputs(30)));
    layer0_outputs(4053) <= not((inputs(214)) or (inputs(229)));
    layer0_outputs(4054) <= inputs(147);
    layer0_outputs(4055) <= inputs(41);
    layer0_outputs(4056) <= inputs(186);
    layer0_outputs(4057) <= not((inputs(39)) xor (inputs(86)));
    layer0_outputs(4058) <= inputs(230);
    layer0_outputs(4059) <= not((inputs(47)) or (inputs(170)));
    layer0_outputs(4060) <= (inputs(87)) and not (inputs(95));
    layer0_outputs(4061) <= not(inputs(187));
    layer0_outputs(4062) <= (inputs(151)) and not (inputs(102));
    layer0_outputs(4063) <= (inputs(231)) or (inputs(221));
    layer0_outputs(4064) <= not(inputs(246));
    layer0_outputs(4065) <= '1';
    layer0_outputs(4066) <= not(inputs(89)) or (inputs(201));
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= (inputs(15)) and (inputs(2));
    layer0_outputs(4069) <= (inputs(88)) or (inputs(252));
    layer0_outputs(4070) <= (inputs(8)) and not (inputs(164));
    layer0_outputs(4071) <= (inputs(33)) or (inputs(65));
    layer0_outputs(4072) <= not(inputs(35));
    layer0_outputs(4073) <= inputs(81);
    layer0_outputs(4074) <= inputs(234);
    layer0_outputs(4075) <= (inputs(214)) or (inputs(225));
    layer0_outputs(4076) <= (inputs(81)) or (inputs(214));
    layer0_outputs(4077) <= not(inputs(153));
    layer0_outputs(4078) <= inputs(247);
    layer0_outputs(4079) <= (inputs(155)) or (inputs(49));
    layer0_outputs(4080) <= '1';
    layer0_outputs(4081) <= not((inputs(245)) or (inputs(66)));
    layer0_outputs(4082) <= (inputs(90)) or (inputs(4));
    layer0_outputs(4083) <= (inputs(159)) and not (inputs(201));
    layer0_outputs(4084) <= inputs(58);
    layer0_outputs(4085) <= (inputs(238)) xor (inputs(96));
    layer0_outputs(4086) <= not((inputs(97)) xor (inputs(84)));
    layer0_outputs(4087) <= not(inputs(228));
    layer0_outputs(4088) <= '1';
    layer0_outputs(4089) <= not(inputs(162));
    layer0_outputs(4090) <= not((inputs(137)) or (inputs(60)));
    layer0_outputs(4091) <= not((inputs(162)) xor (inputs(60)));
    layer0_outputs(4092) <= not(inputs(135)) or (inputs(143));
    layer0_outputs(4093) <= inputs(232);
    layer0_outputs(4094) <= not((inputs(134)) or (inputs(46)));
    layer0_outputs(4095) <= (inputs(105)) and not (inputs(129));
    layer0_outputs(4096) <= not(inputs(77));
    layer0_outputs(4097) <= inputs(174);
    layer0_outputs(4098) <= not(inputs(98)) or (inputs(170));
    layer0_outputs(4099) <= (inputs(242)) and not (inputs(224));
    layer0_outputs(4100) <= not((inputs(141)) or (inputs(24)));
    layer0_outputs(4101) <= not((inputs(78)) or (inputs(5)));
    layer0_outputs(4102) <= (inputs(93)) or (inputs(35));
    layer0_outputs(4103) <= not(inputs(34));
    layer0_outputs(4104) <= not(inputs(128));
    layer0_outputs(4105) <= not(inputs(216)) or (inputs(89));
    layer0_outputs(4106) <= inputs(185);
    layer0_outputs(4107) <= (inputs(112)) and (inputs(207));
    layer0_outputs(4108) <= (inputs(133)) and not (inputs(111));
    layer0_outputs(4109) <= not((inputs(50)) or (inputs(63)));
    layer0_outputs(4110) <= not(inputs(129));
    layer0_outputs(4111) <= not((inputs(189)) or (inputs(73)));
    layer0_outputs(4112) <= (inputs(33)) or (inputs(248));
    layer0_outputs(4113) <= (inputs(108)) and not (inputs(225));
    layer0_outputs(4114) <= inputs(247);
    layer0_outputs(4115) <= not(inputs(178));
    layer0_outputs(4116) <= inputs(37);
    layer0_outputs(4117) <= not(inputs(200)) or (inputs(129));
    layer0_outputs(4118) <= not(inputs(231)) or (inputs(41));
    layer0_outputs(4119) <= not(inputs(244)) or (inputs(239));
    layer0_outputs(4120) <= not((inputs(38)) xor (inputs(42)));
    layer0_outputs(4121) <= not((inputs(102)) xor (inputs(70)));
    layer0_outputs(4122) <= not((inputs(97)) or (inputs(189)));
    layer0_outputs(4123) <= (inputs(187)) and not (inputs(127));
    layer0_outputs(4124) <= (inputs(38)) and (inputs(73));
    layer0_outputs(4125) <= not(inputs(178));
    layer0_outputs(4126) <= (inputs(57)) xor (inputs(22));
    layer0_outputs(4127) <= (inputs(63)) or (inputs(3));
    layer0_outputs(4128) <= not(inputs(115));
    layer0_outputs(4129) <= not((inputs(234)) xor (inputs(193)));
    layer0_outputs(4130) <= not(inputs(5));
    layer0_outputs(4131) <= (inputs(99)) and not (inputs(10));
    layer0_outputs(4132) <= (inputs(134)) and not (inputs(188));
    layer0_outputs(4133) <= (inputs(173)) and (inputs(109));
    layer0_outputs(4134) <= (inputs(133)) and not (inputs(0));
    layer0_outputs(4135) <= not((inputs(160)) xor (inputs(65)));
    layer0_outputs(4136) <= not(inputs(195)) or (inputs(222));
    layer0_outputs(4137) <= (inputs(181)) and not (inputs(125));
    layer0_outputs(4138) <= not(inputs(7));
    layer0_outputs(4139) <= not(inputs(108));
    layer0_outputs(4140) <= not((inputs(61)) or (inputs(44)));
    layer0_outputs(4141) <= (inputs(210)) and not (inputs(182));
    layer0_outputs(4142) <= not((inputs(153)) and (inputs(183)));
    layer0_outputs(4143) <= not((inputs(248)) or (inputs(208)));
    layer0_outputs(4144) <= not(inputs(198));
    layer0_outputs(4145) <= not((inputs(97)) or (inputs(78)));
    layer0_outputs(4146) <= not(inputs(87)) or (inputs(253));
    layer0_outputs(4147) <= not(inputs(150)) or (inputs(207));
    layer0_outputs(4148) <= not(inputs(47));
    layer0_outputs(4149) <= inputs(232);
    layer0_outputs(4150) <= (inputs(88)) and not (inputs(108));
    layer0_outputs(4151) <= inputs(189);
    layer0_outputs(4152) <= (inputs(246)) and not (inputs(156));
    layer0_outputs(4153) <= not(inputs(120)) or (inputs(49));
    layer0_outputs(4154) <= (inputs(44)) xor (inputs(15));
    layer0_outputs(4155) <= not((inputs(148)) xor (inputs(67)));
    layer0_outputs(4156) <= inputs(212);
    layer0_outputs(4157) <= not(inputs(204)) or (inputs(231));
    layer0_outputs(4158) <= not(inputs(84));
    layer0_outputs(4159) <= '1';
    layer0_outputs(4160) <= not((inputs(143)) xor (inputs(20)));
    layer0_outputs(4161) <= not(inputs(68)) or (inputs(14));
    layer0_outputs(4162) <= '0';
    layer0_outputs(4163) <= not(inputs(139));
    layer0_outputs(4164) <= inputs(192);
    layer0_outputs(4165) <= '1';
    layer0_outputs(4166) <= inputs(37);
    layer0_outputs(4167) <= (inputs(96)) or (inputs(57));
    layer0_outputs(4168) <= inputs(89);
    layer0_outputs(4169) <= not((inputs(231)) and (inputs(62)));
    layer0_outputs(4170) <= (inputs(27)) and (inputs(234));
    layer0_outputs(4171) <= inputs(128);
    layer0_outputs(4172) <= not((inputs(204)) or (inputs(198)));
    layer0_outputs(4173) <= (inputs(165)) or (inputs(97));
    layer0_outputs(4174) <= not(inputs(136)) or (inputs(223));
    layer0_outputs(4175) <= not(inputs(32)) or (inputs(242));
    layer0_outputs(4176) <= inputs(232);
    layer0_outputs(4177) <= not(inputs(214));
    layer0_outputs(4178) <= not((inputs(221)) or (inputs(253)));
    layer0_outputs(4179) <= not(inputs(137));
    layer0_outputs(4180) <= (inputs(22)) and not (inputs(234));
    layer0_outputs(4181) <= '1';
    layer0_outputs(4182) <= (inputs(187)) xor (inputs(222));
    layer0_outputs(4183) <= not((inputs(33)) or (inputs(135)));
    layer0_outputs(4184) <= (inputs(228)) or (inputs(173));
    layer0_outputs(4185) <= not(inputs(155)) or (inputs(14));
    layer0_outputs(4186) <= inputs(99);
    layer0_outputs(4187) <= not(inputs(56));
    layer0_outputs(4188) <= (inputs(145)) or (inputs(37));
    layer0_outputs(4189) <= not(inputs(71)) or (inputs(143));
    layer0_outputs(4190) <= (inputs(28)) xor (inputs(195));
    layer0_outputs(4191) <= not((inputs(21)) or (inputs(194)));
    layer0_outputs(4192) <= inputs(27);
    layer0_outputs(4193) <= not((inputs(186)) xor (inputs(186)));
    layer0_outputs(4194) <= (inputs(197)) or (inputs(226));
    layer0_outputs(4195) <= not(inputs(100));
    layer0_outputs(4196) <= not(inputs(54)) or (inputs(253));
    layer0_outputs(4197) <= inputs(45);
    layer0_outputs(4198) <= not((inputs(9)) and (inputs(32)));
    layer0_outputs(4199) <= not((inputs(7)) or (inputs(240)));
    layer0_outputs(4200) <= inputs(229);
    layer0_outputs(4201) <= not((inputs(141)) or (inputs(212)));
    layer0_outputs(4202) <= (inputs(166)) and not (inputs(204));
    layer0_outputs(4203) <= not((inputs(244)) and (inputs(27)));
    layer0_outputs(4204) <= not((inputs(164)) and (inputs(1)));
    layer0_outputs(4205) <= not((inputs(144)) xor (inputs(132)));
    layer0_outputs(4206) <= not((inputs(224)) xor (inputs(90)));
    layer0_outputs(4207) <= not(inputs(50));
    layer0_outputs(4208) <= inputs(209);
    layer0_outputs(4209) <= (inputs(141)) and (inputs(80));
    layer0_outputs(4210) <= not(inputs(121)) or (inputs(133));
    layer0_outputs(4211) <= inputs(40);
    layer0_outputs(4212) <= not((inputs(36)) xor (inputs(160)));
    layer0_outputs(4213) <= not(inputs(107)) or (inputs(18));
    layer0_outputs(4214) <= not(inputs(107));
    layer0_outputs(4215) <= inputs(250);
    layer0_outputs(4216) <= not((inputs(75)) xor (inputs(110)));
    layer0_outputs(4217) <= not((inputs(205)) or (inputs(190)));
    layer0_outputs(4218) <= (inputs(192)) or (inputs(78));
    layer0_outputs(4219) <= (inputs(225)) or (inputs(244));
    layer0_outputs(4220) <= not(inputs(80));
    layer0_outputs(4221) <= (inputs(144)) and not (inputs(0));
    layer0_outputs(4222) <= not((inputs(61)) xor (inputs(230)));
    layer0_outputs(4223) <= (inputs(149)) xor (inputs(168));
    layer0_outputs(4224) <= not((inputs(126)) xor (inputs(4)));
    layer0_outputs(4225) <= not((inputs(112)) or (inputs(50)));
    layer0_outputs(4226) <= inputs(167);
    layer0_outputs(4227) <= not(inputs(108));
    layer0_outputs(4228) <= inputs(152);
    layer0_outputs(4229) <= '0';
    layer0_outputs(4230) <= not((inputs(253)) or (inputs(5)));
    layer0_outputs(4231) <= not(inputs(39));
    layer0_outputs(4232) <= (inputs(150)) or (inputs(202));
    layer0_outputs(4233) <= (inputs(83)) or (inputs(132));
    layer0_outputs(4234) <= not((inputs(119)) or (inputs(212)));
    layer0_outputs(4235) <= inputs(39);
    layer0_outputs(4236) <= not((inputs(208)) or (inputs(244)));
    layer0_outputs(4237) <= not(inputs(238));
    layer0_outputs(4238) <= (inputs(106)) or (inputs(145));
    layer0_outputs(4239) <= inputs(23);
    layer0_outputs(4240) <= not((inputs(244)) and (inputs(28)));
    layer0_outputs(4241) <= not(inputs(87)) or (inputs(163));
    layer0_outputs(4242) <= (inputs(168)) and not (inputs(189));
    layer0_outputs(4243) <= (inputs(109)) and not (inputs(27));
    layer0_outputs(4244) <= (inputs(30)) and not (inputs(247));
    layer0_outputs(4245) <= not(inputs(86)) or (inputs(65));
    layer0_outputs(4246) <= not(inputs(50)) or (inputs(65));
    layer0_outputs(4247) <= not(inputs(205));
    layer0_outputs(4248) <= not(inputs(176));
    layer0_outputs(4249) <= not((inputs(28)) or (inputs(138)));
    layer0_outputs(4250) <= not(inputs(143));
    layer0_outputs(4251) <= not(inputs(219));
    layer0_outputs(4252) <= '1';
    layer0_outputs(4253) <= inputs(147);
    layer0_outputs(4254) <= not((inputs(53)) xor (inputs(158)));
    layer0_outputs(4255) <= not(inputs(146));
    layer0_outputs(4256) <= not(inputs(139));
    layer0_outputs(4257) <= inputs(105);
    layer0_outputs(4258) <= (inputs(85)) and not (inputs(239));
    layer0_outputs(4259) <= (inputs(201)) and not (inputs(37));
    layer0_outputs(4260) <= not(inputs(62)) or (inputs(47));
    layer0_outputs(4261) <= (inputs(201)) or (inputs(197));
    layer0_outputs(4262) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(4263) <= not((inputs(67)) or (inputs(146)));
    layer0_outputs(4264) <= (inputs(113)) xor (inputs(69));
    layer0_outputs(4265) <= not(inputs(189)) or (inputs(18));
    layer0_outputs(4266) <= not((inputs(169)) and (inputs(155)));
    layer0_outputs(4267) <= (inputs(22)) and not (inputs(183));
    layer0_outputs(4268) <= not(inputs(176));
    layer0_outputs(4269) <= inputs(50);
    layer0_outputs(4270) <= (inputs(227)) and (inputs(199));
    layer0_outputs(4271) <= not((inputs(155)) xor (inputs(20)));
    layer0_outputs(4272) <= inputs(115);
    layer0_outputs(4273) <= inputs(121);
    layer0_outputs(4274) <= not(inputs(73));
    layer0_outputs(4275) <= not(inputs(202)) or (inputs(39));
    layer0_outputs(4276) <= not(inputs(185));
    layer0_outputs(4277) <= inputs(249);
    layer0_outputs(4278) <= not(inputs(38)) or (inputs(190));
    layer0_outputs(4279) <= inputs(82);
    layer0_outputs(4280) <= (inputs(201)) and not (inputs(86));
    layer0_outputs(4281) <= inputs(158);
    layer0_outputs(4282) <= inputs(239);
    layer0_outputs(4283) <= not(inputs(123));
    layer0_outputs(4284) <= inputs(22);
    layer0_outputs(4285) <= (inputs(73)) xor (inputs(65));
    layer0_outputs(4286) <= (inputs(243)) and not (inputs(144));
    layer0_outputs(4287) <= (inputs(245)) and not (inputs(37));
    layer0_outputs(4288) <= not(inputs(190));
    layer0_outputs(4289) <= not((inputs(50)) xor (inputs(45)));
    layer0_outputs(4290) <= (inputs(37)) xor (inputs(45));
    layer0_outputs(4291) <= not(inputs(23));
    layer0_outputs(4292) <= inputs(217);
    layer0_outputs(4293) <= not(inputs(220));
    layer0_outputs(4294) <= inputs(66);
    layer0_outputs(4295) <= not((inputs(5)) or (inputs(134)));
    layer0_outputs(4296) <= not(inputs(39));
    layer0_outputs(4297) <= (inputs(104)) xor (inputs(43));
    layer0_outputs(4298) <= (inputs(138)) and not (inputs(127));
    layer0_outputs(4299) <= not(inputs(28));
    layer0_outputs(4300) <= inputs(198);
    layer0_outputs(4301) <= not(inputs(241));
    layer0_outputs(4302) <= not((inputs(59)) or (inputs(48)));
    layer0_outputs(4303) <= not((inputs(155)) and (inputs(54)));
    layer0_outputs(4304) <= not(inputs(136));
    layer0_outputs(4305) <= (inputs(99)) and not (inputs(117));
    layer0_outputs(4306) <= not((inputs(120)) xor (inputs(255)));
    layer0_outputs(4307) <= not((inputs(89)) and (inputs(38)));
    layer0_outputs(4308) <= not(inputs(17));
    layer0_outputs(4309) <= not((inputs(52)) xor (inputs(34)));
    layer0_outputs(4310) <= (inputs(15)) and not (inputs(110));
    layer0_outputs(4311) <= (inputs(4)) or (inputs(165));
    layer0_outputs(4312) <= inputs(149);
    layer0_outputs(4313) <= not((inputs(115)) or (inputs(29)));
    layer0_outputs(4314) <= not(inputs(236));
    layer0_outputs(4315) <= not(inputs(130));
    layer0_outputs(4316) <= not((inputs(244)) xor (inputs(167)));
    layer0_outputs(4317) <= not((inputs(30)) xor (inputs(213)));
    layer0_outputs(4318) <= not(inputs(82));
    layer0_outputs(4319) <= (inputs(72)) and (inputs(110));
    layer0_outputs(4320) <= not(inputs(86));
    layer0_outputs(4321) <= (inputs(252)) or (inputs(55));
    layer0_outputs(4322) <= (inputs(48)) xor (inputs(80));
    layer0_outputs(4323) <= not((inputs(212)) or (inputs(214)));
    layer0_outputs(4324) <= not(inputs(183)) or (inputs(90));
    layer0_outputs(4325) <= not(inputs(117));
    layer0_outputs(4326) <= not(inputs(85)) or (inputs(125));
    layer0_outputs(4327) <= not(inputs(13)) or (inputs(70));
    layer0_outputs(4328) <= inputs(135);
    layer0_outputs(4329) <= (inputs(162)) and not (inputs(17));
    layer0_outputs(4330) <= inputs(162);
    layer0_outputs(4331) <= (inputs(250)) and not (inputs(108));
    layer0_outputs(4332) <= not((inputs(178)) or (inputs(151)));
    layer0_outputs(4333) <= not(inputs(117)) or (inputs(6));
    layer0_outputs(4334) <= not((inputs(40)) or (inputs(60)));
    layer0_outputs(4335) <= '0';
    layer0_outputs(4336) <= (inputs(11)) or (inputs(34));
    layer0_outputs(4337) <= (inputs(37)) xor (inputs(160));
    layer0_outputs(4338) <= inputs(8);
    layer0_outputs(4339) <= inputs(193);
    layer0_outputs(4340) <= not((inputs(237)) xor (inputs(64)));
    layer0_outputs(4341) <= inputs(156);
    layer0_outputs(4342) <= (inputs(165)) and (inputs(217));
    layer0_outputs(4343) <= '1';
    layer0_outputs(4344) <= not(inputs(223));
    layer0_outputs(4345) <= not((inputs(146)) or (inputs(193)));
    layer0_outputs(4346) <= not(inputs(87)) or (inputs(214));
    layer0_outputs(4347) <= not(inputs(107));
    layer0_outputs(4348) <= not((inputs(18)) xor (inputs(125)));
    layer0_outputs(4349) <= '0';
    layer0_outputs(4350) <= (inputs(91)) xor (inputs(228));
    layer0_outputs(4351) <= not((inputs(153)) or (inputs(153)));
    layer0_outputs(4352) <= not(inputs(77));
    layer0_outputs(4353) <= (inputs(11)) or (inputs(151));
    layer0_outputs(4354) <= not((inputs(27)) or (inputs(81)));
    layer0_outputs(4355) <= inputs(214);
    layer0_outputs(4356) <= not((inputs(26)) xor (inputs(222)));
    layer0_outputs(4357) <= not((inputs(105)) and (inputs(28)));
    layer0_outputs(4358) <= '0';
    layer0_outputs(4359) <= not((inputs(79)) xor (inputs(76)));
    layer0_outputs(4360) <= '1';
    layer0_outputs(4361) <= inputs(52);
    layer0_outputs(4362) <= not((inputs(5)) xor (inputs(207)));
    layer0_outputs(4363) <= not(inputs(190)) or (inputs(152));
    layer0_outputs(4364) <= inputs(98);
    layer0_outputs(4365) <= not((inputs(206)) or (inputs(154)));
    layer0_outputs(4366) <= not(inputs(90)) or (inputs(163));
    layer0_outputs(4367) <= (inputs(74)) or (inputs(35));
    layer0_outputs(4368) <= (inputs(160)) or (inputs(209));
    layer0_outputs(4369) <= inputs(166);
    layer0_outputs(4370) <= not(inputs(6));
    layer0_outputs(4371) <= (inputs(161)) or (inputs(153));
    layer0_outputs(4372) <= '1';
    layer0_outputs(4373) <= not(inputs(221));
    layer0_outputs(4374) <= not((inputs(16)) or (inputs(6)));
    layer0_outputs(4375) <= inputs(160);
    layer0_outputs(4376) <= (inputs(65)) xor (inputs(20));
    layer0_outputs(4377) <= not(inputs(74));
    layer0_outputs(4378) <= (inputs(247)) and not (inputs(111));
    layer0_outputs(4379) <= not((inputs(64)) or (inputs(18)));
    layer0_outputs(4380) <= not(inputs(215));
    layer0_outputs(4381) <= inputs(228);
    layer0_outputs(4382) <= not((inputs(162)) or (inputs(25)));
    layer0_outputs(4383) <= '1';
    layer0_outputs(4384) <= (inputs(75)) or (inputs(17));
    layer0_outputs(4385) <= (inputs(221)) or (inputs(173));
    layer0_outputs(4386) <= not(inputs(226));
    layer0_outputs(4387) <= inputs(157);
    layer0_outputs(4388) <= (inputs(246)) or (inputs(50));
    layer0_outputs(4389) <= inputs(221);
    layer0_outputs(4390) <= inputs(230);
    layer0_outputs(4391) <= not(inputs(136));
    layer0_outputs(4392) <= not(inputs(70)) or (inputs(140));
    layer0_outputs(4393) <= not(inputs(192)) or (inputs(36));
    layer0_outputs(4394) <= (inputs(248)) or (inputs(173));
    layer0_outputs(4395) <= not(inputs(73));
    layer0_outputs(4396) <= inputs(88);
    layer0_outputs(4397) <= not(inputs(201));
    layer0_outputs(4398) <= (inputs(197)) xor (inputs(45));
    layer0_outputs(4399) <= not((inputs(32)) or (inputs(111)));
    layer0_outputs(4400) <= inputs(109);
    layer0_outputs(4401) <= not(inputs(195));
    layer0_outputs(4402) <= (inputs(113)) or (inputs(178));
    layer0_outputs(4403) <= not((inputs(238)) or (inputs(187)));
    layer0_outputs(4404) <= not(inputs(193));
    layer0_outputs(4405) <= inputs(195);
    layer0_outputs(4406) <= not(inputs(147));
    layer0_outputs(4407) <= inputs(129);
    layer0_outputs(4408) <= not((inputs(191)) or (inputs(193)));
    layer0_outputs(4409) <= (inputs(108)) or (inputs(227));
    layer0_outputs(4410) <= (inputs(169)) and not (inputs(227));
    layer0_outputs(4411) <= not((inputs(197)) or (inputs(179)));
    layer0_outputs(4412) <= not(inputs(11));
    layer0_outputs(4413) <= not(inputs(193));
    layer0_outputs(4414) <= (inputs(99)) or (inputs(81));
    layer0_outputs(4415) <= inputs(157);
    layer0_outputs(4416) <= not(inputs(136)) or (inputs(205));
    layer0_outputs(4417) <= inputs(230);
    layer0_outputs(4418) <= inputs(90);
    layer0_outputs(4419) <= (inputs(178)) or (inputs(176));
    layer0_outputs(4420) <= not(inputs(214));
    layer0_outputs(4421) <= not((inputs(225)) xor (inputs(209)));
    layer0_outputs(4422) <= not((inputs(137)) xor (inputs(187)));
    layer0_outputs(4423) <= (inputs(90)) and not (inputs(86));
    layer0_outputs(4424) <= inputs(62);
    layer0_outputs(4425) <= not(inputs(177));
    layer0_outputs(4426) <= not((inputs(2)) xor (inputs(60)));
    layer0_outputs(4427) <= not(inputs(184)) or (inputs(175));
    layer0_outputs(4428) <= not((inputs(99)) xor (inputs(23)));
    layer0_outputs(4429) <= not(inputs(148));
    layer0_outputs(4430) <= (inputs(240)) or (inputs(153));
    layer0_outputs(4431) <= not(inputs(25)) or (inputs(4));
    layer0_outputs(4432) <= (inputs(151)) xor (inputs(167));
    layer0_outputs(4433) <= inputs(219);
    layer0_outputs(4434) <= (inputs(199)) xor (inputs(136));
    layer0_outputs(4435) <= (inputs(190)) or (inputs(228));
    layer0_outputs(4436) <= inputs(43);
    layer0_outputs(4437) <= not(inputs(75));
    layer0_outputs(4438) <= (inputs(61)) or (inputs(74));
    layer0_outputs(4439) <= (inputs(56)) or (inputs(179));
    layer0_outputs(4440) <= not(inputs(27)) or (inputs(219));
    layer0_outputs(4441) <= (inputs(69)) and not (inputs(175));
    layer0_outputs(4442) <= inputs(118);
    layer0_outputs(4443) <= not(inputs(100)) or (inputs(182));
    layer0_outputs(4444) <= not(inputs(211));
    layer0_outputs(4445) <= not((inputs(223)) or (inputs(182)));
    layer0_outputs(4446) <= (inputs(161)) or (inputs(190));
    layer0_outputs(4447) <= inputs(210);
    layer0_outputs(4448) <= not((inputs(17)) or (inputs(106)));
    layer0_outputs(4449) <= not(inputs(25));
    layer0_outputs(4450) <= (inputs(150)) or (inputs(81));
    layer0_outputs(4451) <= not(inputs(129));
    layer0_outputs(4452) <= (inputs(200)) or (inputs(192));
    layer0_outputs(4453) <= (inputs(64)) or (inputs(162));
    layer0_outputs(4454) <= not((inputs(251)) or (inputs(229)));
    layer0_outputs(4455) <= (inputs(134)) xor (inputs(196));
    layer0_outputs(4456) <= inputs(58);
    layer0_outputs(4457) <= inputs(182);
    layer0_outputs(4458) <= not(inputs(147));
    layer0_outputs(4459) <= not(inputs(51));
    layer0_outputs(4460) <= not((inputs(70)) xor (inputs(17)));
    layer0_outputs(4461) <= not(inputs(51));
    layer0_outputs(4462) <= not(inputs(229));
    layer0_outputs(4463) <= not((inputs(123)) or (inputs(97)));
    layer0_outputs(4464) <= not((inputs(226)) or (inputs(191)));
    layer0_outputs(4465) <= not((inputs(14)) or (inputs(132)));
    layer0_outputs(4466) <= not(inputs(22));
    layer0_outputs(4467) <= not(inputs(210));
    layer0_outputs(4468) <= not(inputs(164));
    layer0_outputs(4469) <= inputs(254);
    layer0_outputs(4470) <= not((inputs(154)) or (inputs(244)));
    layer0_outputs(4471) <= (inputs(4)) or (inputs(24));
    layer0_outputs(4472) <= not(inputs(14)) or (inputs(224));
    layer0_outputs(4473) <= inputs(230);
    layer0_outputs(4474) <= inputs(126);
    layer0_outputs(4475) <= (inputs(123)) xor (inputs(237));
    layer0_outputs(4476) <= inputs(239);
    layer0_outputs(4477) <= not(inputs(77));
    layer0_outputs(4478) <= (inputs(139)) or (inputs(84));
    layer0_outputs(4479) <= inputs(107);
    layer0_outputs(4480) <= (inputs(159)) xor (inputs(42));
    layer0_outputs(4481) <= (inputs(124)) or (inputs(72));
    layer0_outputs(4482) <= not(inputs(253));
    layer0_outputs(4483) <= (inputs(13)) or (inputs(195));
    layer0_outputs(4484) <= (inputs(228)) or (inputs(255));
    layer0_outputs(4485) <= '1';
    layer0_outputs(4486) <= not((inputs(147)) xor (inputs(172)));
    layer0_outputs(4487) <= inputs(158);
    layer0_outputs(4488) <= (inputs(43)) or (inputs(251));
    layer0_outputs(4489) <= (inputs(41)) or (inputs(6));
    layer0_outputs(4490) <= (inputs(195)) and not (inputs(140));
    layer0_outputs(4491) <= not((inputs(164)) or (inputs(75)));
    layer0_outputs(4492) <= inputs(151);
    layer0_outputs(4493) <= not((inputs(85)) xor (inputs(116)));
    layer0_outputs(4494) <= (inputs(166)) and (inputs(229));
    layer0_outputs(4495) <= not(inputs(68));
    layer0_outputs(4496) <= not(inputs(221)) or (inputs(134));
    layer0_outputs(4497) <= not((inputs(27)) or (inputs(162)));
    layer0_outputs(4498) <= not((inputs(60)) and (inputs(88)));
    layer0_outputs(4499) <= (inputs(27)) and (inputs(114));
    layer0_outputs(4500) <= inputs(246);
    layer0_outputs(4501) <= not(inputs(92));
    layer0_outputs(4502) <= (inputs(211)) or (inputs(63));
    layer0_outputs(4503) <= not(inputs(103));
    layer0_outputs(4504) <= '1';
    layer0_outputs(4505) <= not(inputs(61));
    layer0_outputs(4506) <= not(inputs(26));
    layer0_outputs(4507) <= not(inputs(93)) or (inputs(64));
    layer0_outputs(4508) <= not(inputs(123)) or (inputs(246));
    layer0_outputs(4509) <= not((inputs(65)) or (inputs(60)));
    layer0_outputs(4510) <= (inputs(150)) xor (inputs(111));
    layer0_outputs(4511) <= (inputs(182)) or (inputs(207));
    layer0_outputs(4512) <= inputs(131);
    layer0_outputs(4513) <= not((inputs(249)) or (inputs(251)));
    layer0_outputs(4514) <= (inputs(40)) or (inputs(204));
    layer0_outputs(4515) <= (inputs(147)) or (inputs(31));
    layer0_outputs(4516) <= (inputs(80)) xor (inputs(144));
    layer0_outputs(4517) <= inputs(27);
    layer0_outputs(4518) <= not((inputs(115)) or (inputs(238)));
    layer0_outputs(4519) <= (inputs(69)) and not (inputs(240));
    layer0_outputs(4520) <= not((inputs(117)) xor (inputs(21)));
    layer0_outputs(4521) <= (inputs(250)) xor (inputs(156));
    layer0_outputs(4522) <= not(inputs(187)) or (inputs(30));
    layer0_outputs(4523) <= (inputs(20)) or (inputs(242));
    layer0_outputs(4524) <= inputs(41);
    layer0_outputs(4525) <= not((inputs(128)) or (inputs(67)));
    layer0_outputs(4526) <= not((inputs(223)) or (inputs(174)));
    layer0_outputs(4527) <= not(inputs(160));
    layer0_outputs(4528) <= inputs(84);
    layer0_outputs(4529) <= inputs(228);
    layer0_outputs(4530) <= not((inputs(106)) or (inputs(109)));
    layer0_outputs(4531) <= not((inputs(236)) or (inputs(148)));
    layer0_outputs(4532) <= not((inputs(21)) xor (inputs(169)));
    layer0_outputs(4533) <= not(inputs(38)) or (inputs(174));
    layer0_outputs(4534) <= (inputs(72)) and (inputs(142));
    layer0_outputs(4535) <= not((inputs(147)) or (inputs(54)));
    layer0_outputs(4536) <= (inputs(236)) xor (inputs(35));
    layer0_outputs(4537) <= not(inputs(90));
    layer0_outputs(4538) <= not(inputs(103));
    layer0_outputs(4539) <= (inputs(80)) or (inputs(194));
    layer0_outputs(4540) <= (inputs(190)) xor (inputs(78));
    layer0_outputs(4541) <= inputs(126);
    layer0_outputs(4542) <= inputs(3);
    layer0_outputs(4543) <= (inputs(90)) xor (inputs(96));
    layer0_outputs(4544) <= not((inputs(110)) xor (inputs(206)));
    layer0_outputs(4545) <= not(inputs(167));
    layer0_outputs(4546) <= (inputs(35)) or (inputs(25));
    layer0_outputs(4547) <= inputs(84);
    layer0_outputs(4548) <= inputs(7);
    layer0_outputs(4549) <= (inputs(104)) and not (inputs(96));
    layer0_outputs(4550) <= not(inputs(72)) or (inputs(138));
    layer0_outputs(4551) <= not(inputs(146)) or (inputs(156));
    layer0_outputs(4552) <= '1';
    layer0_outputs(4553) <= inputs(109);
    layer0_outputs(4554) <= not((inputs(249)) xor (inputs(235)));
    layer0_outputs(4555) <= not((inputs(0)) or (inputs(134)));
    layer0_outputs(4556) <= not(inputs(183));
    layer0_outputs(4557) <= not((inputs(148)) or (inputs(223)));
    layer0_outputs(4558) <= not((inputs(155)) or (inputs(78)));
    layer0_outputs(4559) <= not(inputs(20));
    layer0_outputs(4560) <= not((inputs(187)) or (inputs(202)));
    layer0_outputs(4561) <= inputs(195);
    layer0_outputs(4562) <= '0';
    layer0_outputs(4563) <= inputs(6);
    layer0_outputs(4564) <= not((inputs(76)) and (inputs(116)));
    layer0_outputs(4565) <= (inputs(218)) and not (inputs(25));
    layer0_outputs(4566) <= (inputs(11)) or (inputs(49));
    layer0_outputs(4567) <= not(inputs(9)) or (inputs(18));
    layer0_outputs(4568) <= (inputs(125)) or (inputs(198));
    layer0_outputs(4569) <= not(inputs(76));
    layer0_outputs(4570) <= (inputs(223)) or (inputs(30));
    layer0_outputs(4571) <= not((inputs(174)) xor (inputs(164)));
    layer0_outputs(4572) <= (inputs(31)) xor (inputs(13));
    layer0_outputs(4573) <= not(inputs(92));
    layer0_outputs(4574) <= not(inputs(203)) or (inputs(124));
    layer0_outputs(4575) <= (inputs(132)) and not (inputs(53));
    layer0_outputs(4576) <= (inputs(66)) or (inputs(159));
    layer0_outputs(4577) <= (inputs(214)) and not (inputs(224));
    layer0_outputs(4578) <= not(inputs(233));
    layer0_outputs(4579) <= inputs(67);
    layer0_outputs(4580) <= not(inputs(29));
    layer0_outputs(4581) <= not((inputs(229)) xor (inputs(190)));
    layer0_outputs(4582) <= not((inputs(123)) xor (inputs(4)));
    layer0_outputs(4583) <= (inputs(8)) and not (inputs(221));
    layer0_outputs(4584) <= (inputs(165)) and not (inputs(58));
    layer0_outputs(4585) <= not((inputs(25)) xor (inputs(33)));
    layer0_outputs(4586) <= not(inputs(76));
    layer0_outputs(4587) <= (inputs(156)) and not (inputs(71));
    layer0_outputs(4588) <= (inputs(185)) xor (inputs(121));
    layer0_outputs(4589) <= '0';
    layer0_outputs(4590) <= (inputs(24)) or (inputs(14));
    layer0_outputs(4591) <= (inputs(25)) and not (inputs(201));
    layer0_outputs(4592) <= (inputs(111)) or (inputs(120));
    layer0_outputs(4593) <= not((inputs(78)) or (inputs(238)));
    layer0_outputs(4594) <= not(inputs(18));
    layer0_outputs(4595) <= not((inputs(43)) xor (inputs(89)));
    layer0_outputs(4596) <= (inputs(231)) or (inputs(243));
    layer0_outputs(4597) <= inputs(89);
    layer0_outputs(4598) <= not((inputs(95)) or (inputs(191)));
    layer0_outputs(4599) <= not(inputs(154)) or (inputs(16));
    layer0_outputs(4600) <= not(inputs(226));
    layer0_outputs(4601) <= (inputs(0)) or (inputs(211));
    layer0_outputs(4602) <= (inputs(136)) and not (inputs(111));
    layer0_outputs(4603) <= not(inputs(169)) or (inputs(42));
    layer0_outputs(4604) <= not((inputs(243)) or (inputs(66)));
    layer0_outputs(4605) <= not((inputs(234)) and (inputs(117)));
    layer0_outputs(4606) <= not(inputs(77));
    layer0_outputs(4607) <= (inputs(225)) and not (inputs(4));
    layer0_outputs(4608) <= (inputs(87)) or (inputs(156));
    layer0_outputs(4609) <= inputs(36);
    layer0_outputs(4610) <= not((inputs(11)) or (inputs(43)));
    layer0_outputs(4611) <= not((inputs(84)) or (inputs(234)));
    layer0_outputs(4612) <= inputs(214);
    layer0_outputs(4613) <= (inputs(155)) or (inputs(220));
    layer0_outputs(4614) <= not(inputs(183)) or (inputs(218));
    layer0_outputs(4615) <= (inputs(210)) or (inputs(101));
    layer0_outputs(4616) <= inputs(145);
    layer0_outputs(4617) <= '1';
    layer0_outputs(4618) <= not((inputs(119)) and (inputs(60)));
    layer0_outputs(4619) <= (inputs(220)) xor (inputs(204));
    layer0_outputs(4620) <= inputs(168);
    layer0_outputs(4621) <= not(inputs(72)) or (inputs(82));
    layer0_outputs(4622) <= not(inputs(90)) or (inputs(189));
    layer0_outputs(4623) <= not((inputs(179)) and (inputs(222)));
    layer0_outputs(4624) <= not((inputs(92)) or (inputs(73)));
    layer0_outputs(4625) <= not(inputs(102));
    layer0_outputs(4626) <= not(inputs(252));
    layer0_outputs(4627) <= inputs(111);
    layer0_outputs(4628) <= not(inputs(180));
    layer0_outputs(4629) <= inputs(164);
    layer0_outputs(4630) <= (inputs(10)) xor (inputs(42));
    layer0_outputs(4631) <= not((inputs(185)) and (inputs(211)));
    layer0_outputs(4632) <= (inputs(164)) or (inputs(227));
    layer0_outputs(4633) <= inputs(61);
    layer0_outputs(4634) <= not((inputs(191)) or (inputs(68)));
    layer0_outputs(4635) <= (inputs(76)) and not (inputs(199));
    layer0_outputs(4636) <= (inputs(133)) and not (inputs(185));
    layer0_outputs(4637) <= inputs(166);
    layer0_outputs(4638) <= not(inputs(152)) or (inputs(228));
    layer0_outputs(4639) <= (inputs(255)) or (inputs(184));
    layer0_outputs(4640) <= not(inputs(106)) or (inputs(132));
    layer0_outputs(4641) <= not(inputs(218));
    layer0_outputs(4642) <= not(inputs(181));
    layer0_outputs(4643) <= inputs(76);
    layer0_outputs(4644) <= (inputs(255)) xor (inputs(146));
    layer0_outputs(4645) <= inputs(87);
    layer0_outputs(4646) <= inputs(38);
    layer0_outputs(4647) <= not((inputs(99)) or (inputs(146)));
    layer0_outputs(4648) <= not((inputs(19)) or (inputs(155)));
    layer0_outputs(4649) <= not(inputs(247));
    layer0_outputs(4650) <= (inputs(227)) and (inputs(207));
    layer0_outputs(4651) <= (inputs(203)) or (inputs(107));
    layer0_outputs(4652) <= (inputs(238)) or (inputs(54));
    layer0_outputs(4653) <= not((inputs(7)) or (inputs(114)));
    layer0_outputs(4654) <= (inputs(200)) and (inputs(103));
    layer0_outputs(4655) <= not(inputs(88));
    layer0_outputs(4656) <= not(inputs(199)) or (inputs(118));
    layer0_outputs(4657) <= not(inputs(196));
    layer0_outputs(4658) <= inputs(251);
    layer0_outputs(4659) <= (inputs(209)) and not (inputs(97));
    layer0_outputs(4660) <= (inputs(207)) or (inputs(237));
    layer0_outputs(4661) <= (inputs(236)) or (inputs(239));
    layer0_outputs(4662) <= not(inputs(8)) or (inputs(180));
    layer0_outputs(4663) <= not(inputs(146));
    layer0_outputs(4664) <= not(inputs(178));
    layer0_outputs(4665) <= not((inputs(164)) xor (inputs(103)));
    layer0_outputs(4666) <= (inputs(74)) and not (inputs(112));
    layer0_outputs(4667) <= inputs(210);
    layer0_outputs(4668) <= not((inputs(90)) xor (inputs(122)));
    layer0_outputs(4669) <= (inputs(220)) or (inputs(157));
    layer0_outputs(4670) <= (inputs(113)) or (inputs(203));
    layer0_outputs(4671) <= not(inputs(142));
    layer0_outputs(4672) <= not(inputs(53)) or (inputs(174));
    layer0_outputs(4673) <= inputs(211);
    layer0_outputs(4674) <= '1';
    layer0_outputs(4675) <= not((inputs(175)) and (inputs(98)));
    layer0_outputs(4676) <= not((inputs(46)) xor (inputs(75)));
    layer0_outputs(4677) <= not((inputs(22)) xor (inputs(70)));
    layer0_outputs(4678) <= not((inputs(27)) and (inputs(9)));
    layer0_outputs(4679) <= not((inputs(60)) and (inputs(78)));
    layer0_outputs(4680) <= (inputs(200)) and not (inputs(96));
    layer0_outputs(4681) <= inputs(203);
    layer0_outputs(4682) <= (inputs(202)) xor (inputs(37));
    layer0_outputs(4683) <= not(inputs(99));
    layer0_outputs(4684) <= not((inputs(213)) xor (inputs(206)));
    layer0_outputs(4685) <= not((inputs(177)) or (inputs(133)));
    layer0_outputs(4686) <= not((inputs(202)) or (inputs(241)));
    layer0_outputs(4687) <= not((inputs(253)) xor (inputs(223)));
    layer0_outputs(4688) <= (inputs(207)) or (inputs(103));
    layer0_outputs(4689) <= inputs(46);
    layer0_outputs(4690) <= (inputs(104)) xor (inputs(178));
    layer0_outputs(4691) <= not(inputs(184));
    layer0_outputs(4692) <= not(inputs(229));
    layer0_outputs(4693) <= not(inputs(119));
    layer0_outputs(4694) <= not((inputs(116)) and (inputs(59)));
    layer0_outputs(4695) <= (inputs(39)) xor (inputs(11));
    layer0_outputs(4696) <= not((inputs(63)) or (inputs(229)));
    layer0_outputs(4697) <= (inputs(246)) and not (inputs(5));
    layer0_outputs(4698) <= inputs(231);
    layer0_outputs(4699) <= (inputs(151)) or (inputs(140));
    layer0_outputs(4700) <= not(inputs(152)) or (inputs(206));
    layer0_outputs(4701) <= not((inputs(1)) or (inputs(122)));
    layer0_outputs(4702) <= inputs(71);
    layer0_outputs(4703) <= not(inputs(23)) or (inputs(113));
    layer0_outputs(4704) <= not((inputs(206)) or (inputs(249)));
    layer0_outputs(4705) <= not((inputs(148)) xor (inputs(193)));
    layer0_outputs(4706) <= '1';
    layer0_outputs(4707) <= inputs(217);
    layer0_outputs(4708) <= not(inputs(14));
    layer0_outputs(4709) <= (inputs(194)) xor (inputs(237));
    layer0_outputs(4710) <= not((inputs(102)) or (inputs(142)));
    layer0_outputs(4711) <= inputs(0);
    layer0_outputs(4712) <= inputs(75);
    layer0_outputs(4713) <= (inputs(77)) xor (inputs(247));
    layer0_outputs(4714) <= (inputs(21)) and not (inputs(45));
    layer0_outputs(4715) <= not(inputs(176));
    layer0_outputs(4716) <= not(inputs(144)) or (inputs(173));
    layer0_outputs(4717) <= not(inputs(218)) or (inputs(30));
    layer0_outputs(4718) <= not(inputs(52)) or (inputs(247));
    layer0_outputs(4719) <= (inputs(238)) xor (inputs(68));
    layer0_outputs(4720) <= not(inputs(233)) or (inputs(17));
    layer0_outputs(4721) <= (inputs(131)) xor (inputs(133));
    layer0_outputs(4722) <= not((inputs(108)) xor (inputs(50)));
    layer0_outputs(4723) <= not(inputs(218));
    layer0_outputs(4724) <= not(inputs(91));
    layer0_outputs(4725) <= '1';
    layer0_outputs(4726) <= (inputs(92)) or (inputs(105));
    layer0_outputs(4727) <= (inputs(91)) xor (inputs(158));
    layer0_outputs(4728) <= not(inputs(29)) or (inputs(69));
    layer0_outputs(4729) <= (inputs(171)) or (inputs(8));
    layer0_outputs(4730) <= not((inputs(126)) xor (inputs(12)));
    layer0_outputs(4731) <= (inputs(113)) xor (inputs(161));
    layer0_outputs(4732) <= not(inputs(67));
    layer0_outputs(4733) <= not((inputs(187)) or (inputs(144)));
    layer0_outputs(4734) <= (inputs(55)) or (inputs(233));
    layer0_outputs(4735) <= not(inputs(36));
    layer0_outputs(4736) <= not((inputs(8)) and (inputs(154)));
    layer0_outputs(4737) <= not(inputs(248));
    layer0_outputs(4738) <= not((inputs(224)) and (inputs(42)));
    layer0_outputs(4739) <= '1';
    layer0_outputs(4740) <= not(inputs(232));
    layer0_outputs(4741) <= not((inputs(209)) xor (inputs(205)));
    layer0_outputs(4742) <= inputs(122);
    layer0_outputs(4743) <= not(inputs(19)) or (inputs(13));
    layer0_outputs(4744) <= not(inputs(24));
    layer0_outputs(4745) <= not(inputs(44));
    layer0_outputs(4746) <= inputs(232);
    layer0_outputs(4747) <= not((inputs(174)) xor (inputs(141)));
    layer0_outputs(4748) <= (inputs(28)) or (inputs(116));
    layer0_outputs(4749) <= (inputs(130)) xor (inputs(117));
    layer0_outputs(4750) <= not(inputs(119)) or (inputs(198));
    layer0_outputs(4751) <= (inputs(49)) xor (inputs(139));
    layer0_outputs(4752) <= (inputs(105)) and not (inputs(159));
    layer0_outputs(4753) <= inputs(237);
    layer0_outputs(4754) <= not(inputs(253));
    layer0_outputs(4755) <= (inputs(47)) and (inputs(92));
    layer0_outputs(4756) <= not(inputs(186));
    layer0_outputs(4757) <= not((inputs(47)) xor (inputs(130)));
    layer0_outputs(4758) <= not(inputs(76));
    layer0_outputs(4759) <= inputs(203);
    layer0_outputs(4760) <= not((inputs(8)) xor (inputs(111)));
    layer0_outputs(4761) <= not(inputs(14));
    layer0_outputs(4762) <= not(inputs(136)) or (inputs(0));
    layer0_outputs(4763) <= (inputs(222)) or (inputs(57));
    layer0_outputs(4764) <= (inputs(193)) and not (inputs(88));
    layer0_outputs(4765) <= (inputs(169)) or (inputs(151));
    layer0_outputs(4766) <= not(inputs(107));
    layer0_outputs(4767) <= not(inputs(8)) or (inputs(52));
    layer0_outputs(4768) <= inputs(52);
    layer0_outputs(4769) <= not((inputs(162)) or (inputs(3)));
    layer0_outputs(4770) <= (inputs(153)) xor (inputs(253));
    layer0_outputs(4771) <= inputs(147);
    layer0_outputs(4772) <= (inputs(45)) and not (inputs(235));
    layer0_outputs(4773) <= '1';
    layer0_outputs(4774) <= not(inputs(84)) or (inputs(50));
    layer0_outputs(4775) <= inputs(166);
    layer0_outputs(4776) <= not(inputs(104)) or (inputs(212));
    layer0_outputs(4777) <= (inputs(44)) and not (inputs(216));
    layer0_outputs(4778) <= (inputs(38)) or (inputs(254));
    layer0_outputs(4779) <= inputs(103);
    layer0_outputs(4780) <= not((inputs(20)) or (inputs(203)));
    layer0_outputs(4781) <= not(inputs(232)) or (inputs(226));
    layer0_outputs(4782) <= not(inputs(110));
    layer0_outputs(4783) <= inputs(135);
    layer0_outputs(4784) <= not(inputs(118));
    layer0_outputs(4785) <= not(inputs(229)) or (inputs(16));
    layer0_outputs(4786) <= not(inputs(168));
    layer0_outputs(4787) <= inputs(138);
    layer0_outputs(4788) <= not(inputs(246)) or (inputs(207));
    layer0_outputs(4789) <= not((inputs(158)) or (inputs(146)));
    layer0_outputs(4790) <= (inputs(223)) xor (inputs(242));
    layer0_outputs(4791) <= not(inputs(8)) or (inputs(253));
    layer0_outputs(4792) <= (inputs(134)) and not (inputs(79));
    layer0_outputs(4793) <= inputs(75);
    layer0_outputs(4794) <= inputs(18);
    layer0_outputs(4795) <= (inputs(151)) and not (inputs(51));
    layer0_outputs(4796) <= (inputs(72)) and not (inputs(78));
    layer0_outputs(4797) <= (inputs(2)) or (inputs(175));
    layer0_outputs(4798) <= inputs(85);
    layer0_outputs(4799) <= not((inputs(234)) xor (inputs(145)));
    layer0_outputs(4800) <= inputs(138);
    layer0_outputs(4801) <= not((inputs(7)) or (inputs(171)));
    layer0_outputs(4802) <= (inputs(45)) xor (inputs(106));
    layer0_outputs(4803) <= not(inputs(77));
    layer0_outputs(4804) <= not(inputs(53));
    layer0_outputs(4805) <= (inputs(54)) or (inputs(152));
    layer0_outputs(4806) <= not(inputs(207));
    layer0_outputs(4807) <= (inputs(67)) or (inputs(29));
    layer0_outputs(4808) <= not((inputs(28)) or (inputs(1)));
    layer0_outputs(4809) <= (inputs(5)) and (inputs(44));
    layer0_outputs(4810) <= inputs(8);
    layer0_outputs(4811) <= not((inputs(52)) or (inputs(171)));
    layer0_outputs(4812) <= (inputs(90)) and not (inputs(172));
    layer0_outputs(4813) <= not(inputs(230));
    layer0_outputs(4814) <= (inputs(60)) or (inputs(47));
    layer0_outputs(4815) <= inputs(22);
    layer0_outputs(4816) <= (inputs(212)) or (inputs(203));
    layer0_outputs(4817) <= not(inputs(108)) or (inputs(19));
    layer0_outputs(4818) <= not(inputs(228));
    layer0_outputs(4819) <= not(inputs(232));
    layer0_outputs(4820) <= not(inputs(118));
    layer0_outputs(4821) <= inputs(249);
    layer0_outputs(4822) <= not((inputs(198)) or (inputs(230)));
    layer0_outputs(4823) <= (inputs(192)) or (inputs(86));
    layer0_outputs(4824) <= (inputs(43)) xor (inputs(41));
    layer0_outputs(4825) <= inputs(216);
    layer0_outputs(4826) <= inputs(120);
    layer0_outputs(4827) <= not(inputs(222));
    layer0_outputs(4828) <= (inputs(72)) xor (inputs(8));
    layer0_outputs(4829) <= not(inputs(53));
    layer0_outputs(4830) <= inputs(124);
    layer0_outputs(4831) <= (inputs(82)) xor (inputs(166));
    layer0_outputs(4832) <= not(inputs(124)) or (inputs(154));
    layer0_outputs(4833) <= inputs(119);
    layer0_outputs(4834) <= not(inputs(146));
    layer0_outputs(4835) <= (inputs(3)) or (inputs(17));
    layer0_outputs(4836) <= not((inputs(56)) or (inputs(211)));
    layer0_outputs(4837) <= (inputs(16)) or (inputs(248));
    layer0_outputs(4838) <= not(inputs(60));
    layer0_outputs(4839) <= not((inputs(61)) xor (inputs(119)));
    layer0_outputs(4840) <= inputs(46);
    layer0_outputs(4841) <= inputs(82);
    layer0_outputs(4842) <= not((inputs(92)) xor (inputs(210)));
    layer0_outputs(4843) <= (inputs(209)) or (inputs(69));
    layer0_outputs(4844) <= (inputs(76)) and not (inputs(15));
    layer0_outputs(4845) <= inputs(193);
    layer0_outputs(4846) <= inputs(57);
    layer0_outputs(4847) <= not(inputs(212));
    layer0_outputs(4848) <= inputs(21);
    layer0_outputs(4849) <= inputs(29);
    layer0_outputs(4850) <= not((inputs(136)) and (inputs(60)));
    layer0_outputs(4851) <= inputs(144);
    layer0_outputs(4852) <= inputs(212);
    layer0_outputs(4853) <= (inputs(27)) and not (inputs(148));
    layer0_outputs(4854) <= not((inputs(194)) xor (inputs(78)));
    layer0_outputs(4855) <= not(inputs(194)) or (inputs(241));
    layer0_outputs(4856) <= inputs(30);
    layer0_outputs(4857) <= not(inputs(222));
    layer0_outputs(4858) <= (inputs(117)) and not (inputs(117));
    layer0_outputs(4859) <= not((inputs(196)) xor (inputs(149)));
    layer0_outputs(4860) <= '0';
    layer0_outputs(4861) <= inputs(123);
    layer0_outputs(4862) <= not((inputs(241)) xor (inputs(90)));
    layer0_outputs(4863) <= (inputs(237)) xor (inputs(222));
    layer0_outputs(4864) <= not((inputs(25)) or (inputs(254)));
    layer0_outputs(4865) <= not(inputs(222)) or (inputs(47));
    layer0_outputs(4866) <= not((inputs(14)) or (inputs(52)));
    layer0_outputs(4867) <= not((inputs(148)) and (inputs(56)));
    layer0_outputs(4868) <= inputs(227);
    layer0_outputs(4869) <= not((inputs(32)) xor (inputs(1)));
    layer0_outputs(4870) <= not((inputs(18)) or (inputs(193)));
    layer0_outputs(4871) <= (inputs(250)) or (inputs(160));
    layer0_outputs(4872) <= inputs(24);
    layer0_outputs(4873) <= (inputs(15)) or (inputs(144));
    layer0_outputs(4874) <= not(inputs(109)) or (inputs(152));
    layer0_outputs(4875) <= inputs(230);
    layer0_outputs(4876) <= (inputs(208)) or (inputs(36));
    layer0_outputs(4877) <= not(inputs(32));
    layer0_outputs(4878) <= inputs(84);
    layer0_outputs(4879) <= not(inputs(83));
    layer0_outputs(4880) <= (inputs(203)) or (inputs(34));
    layer0_outputs(4881) <= not(inputs(255)) or (inputs(81));
    layer0_outputs(4882) <= (inputs(224)) or (inputs(62));
    layer0_outputs(4883) <= not(inputs(104)) or (inputs(3));
    layer0_outputs(4884) <= (inputs(9)) or (inputs(64));
    layer0_outputs(4885) <= (inputs(208)) or (inputs(174));
    layer0_outputs(4886) <= not(inputs(207));
    layer0_outputs(4887) <= not(inputs(125));
    layer0_outputs(4888) <= not(inputs(167));
    layer0_outputs(4889) <= (inputs(159)) or (inputs(187));
    layer0_outputs(4890) <= not(inputs(167));
    layer0_outputs(4891) <= (inputs(97)) or (inputs(227));
    layer0_outputs(4892) <= not((inputs(253)) or (inputs(51)));
    layer0_outputs(4893) <= not((inputs(98)) or (inputs(172)));
    layer0_outputs(4894) <= inputs(189);
    layer0_outputs(4895) <= not((inputs(17)) or (inputs(243)));
    layer0_outputs(4896) <= (inputs(246)) or (inputs(193));
    layer0_outputs(4897) <= not(inputs(185)) or (inputs(226));
    layer0_outputs(4898) <= not((inputs(217)) or (inputs(113)));
    layer0_outputs(4899) <= (inputs(134)) or (inputs(226));
    layer0_outputs(4900) <= inputs(232);
    layer0_outputs(4901) <= not(inputs(68)) or (inputs(21));
    layer0_outputs(4902) <= inputs(223);
    layer0_outputs(4903) <= (inputs(23)) xor (inputs(239));
    layer0_outputs(4904) <= inputs(205);
    layer0_outputs(4905) <= inputs(152);
    layer0_outputs(4906) <= not((inputs(212)) or (inputs(129)));
    layer0_outputs(4907) <= inputs(89);
    layer0_outputs(4908) <= (inputs(40)) and not (inputs(12));
    layer0_outputs(4909) <= '1';
    layer0_outputs(4910) <= not((inputs(51)) and (inputs(39)));
    layer0_outputs(4911) <= not(inputs(182));
    layer0_outputs(4912) <= not(inputs(192));
    layer0_outputs(4913) <= not(inputs(229)) or (inputs(105));
    layer0_outputs(4914) <= (inputs(224)) or (inputs(79));
    layer0_outputs(4915) <= not((inputs(19)) xor (inputs(56)));
    layer0_outputs(4916) <= not((inputs(183)) or (inputs(86)));
    layer0_outputs(4917) <= (inputs(222)) or (inputs(67));
    layer0_outputs(4918) <= (inputs(63)) xor (inputs(158));
    layer0_outputs(4919) <= (inputs(165)) or (inputs(116));
    layer0_outputs(4920) <= (inputs(11)) and (inputs(61));
    layer0_outputs(4921) <= not((inputs(228)) or (inputs(47)));
    layer0_outputs(4922) <= not((inputs(220)) or (inputs(148)));
    layer0_outputs(4923) <= (inputs(148)) and not (inputs(236));
    layer0_outputs(4924) <= not(inputs(202)) or (inputs(2));
    layer0_outputs(4925) <= (inputs(83)) or (inputs(84));
    layer0_outputs(4926) <= not((inputs(191)) or (inputs(42)));
    layer0_outputs(4927) <= (inputs(29)) and not (inputs(116));
    layer0_outputs(4928) <= (inputs(243)) or (inputs(65));
    layer0_outputs(4929) <= (inputs(141)) xor (inputs(161));
    layer0_outputs(4930) <= not(inputs(154));
    layer0_outputs(4931) <= not(inputs(59)) or (inputs(98));
    layer0_outputs(4932) <= not((inputs(160)) xor (inputs(229)));
    layer0_outputs(4933) <= (inputs(220)) or (inputs(180));
    layer0_outputs(4934) <= (inputs(6)) and not (inputs(84));
    layer0_outputs(4935) <= not((inputs(64)) or (inputs(46)));
    layer0_outputs(4936) <= not(inputs(7));
    layer0_outputs(4937) <= not(inputs(170));
    layer0_outputs(4938) <= (inputs(23)) and not (inputs(116));
    layer0_outputs(4939) <= (inputs(60)) xor (inputs(88));
    layer0_outputs(4940) <= not((inputs(213)) or (inputs(173)));
    layer0_outputs(4941) <= not(inputs(43));
    layer0_outputs(4942) <= not((inputs(127)) xor (inputs(95)));
    layer0_outputs(4943) <= not((inputs(176)) or (inputs(111)));
    layer0_outputs(4944) <= not((inputs(43)) xor (inputs(29)));
    layer0_outputs(4945) <= not(inputs(172)) or (inputs(122));
    layer0_outputs(4946) <= (inputs(169)) or (inputs(36));
    layer0_outputs(4947) <= (inputs(194)) and (inputs(142));
    layer0_outputs(4948) <= not((inputs(5)) xor (inputs(20)));
    layer0_outputs(4949) <= not(inputs(83));
    layer0_outputs(4950) <= not((inputs(171)) xor (inputs(188)));
    layer0_outputs(4951) <= not(inputs(127));
    layer0_outputs(4952) <= inputs(20);
    layer0_outputs(4953) <= (inputs(146)) xor (inputs(119));
    layer0_outputs(4954) <= (inputs(79)) xor (inputs(168));
    layer0_outputs(4955) <= inputs(79);
    layer0_outputs(4956) <= '0';
    layer0_outputs(4957) <= not(inputs(65)) or (inputs(109));
    layer0_outputs(4958) <= not((inputs(123)) xor (inputs(12)));
    layer0_outputs(4959) <= (inputs(31)) xor (inputs(19));
    layer0_outputs(4960) <= not(inputs(222));
    layer0_outputs(4961) <= not(inputs(29));
    layer0_outputs(4962) <= not((inputs(157)) xor (inputs(170)));
    layer0_outputs(4963) <= not(inputs(179));
    layer0_outputs(4964) <= not(inputs(52));
    layer0_outputs(4965) <= not(inputs(131));
    layer0_outputs(4966) <= not(inputs(123)) or (inputs(159));
    layer0_outputs(4967) <= inputs(134);
    layer0_outputs(4968) <= inputs(171);
    layer0_outputs(4969) <= not((inputs(199)) or (inputs(3)));
    layer0_outputs(4970) <= inputs(91);
    layer0_outputs(4971) <= (inputs(190)) or (inputs(215));
    layer0_outputs(4972) <= inputs(170);
    layer0_outputs(4973) <= inputs(45);
    layer0_outputs(4974) <= not((inputs(196)) or (inputs(66)));
    layer0_outputs(4975) <= inputs(116);
    layer0_outputs(4976) <= not(inputs(25)) or (inputs(158));
    layer0_outputs(4977) <= '1';
    layer0_outputs(4978) <= not((inputs(77)) or (inputs(7)));
    layer0_outputs(4979) <= (inputs(241)) or (inputs(106));
    layer0_outputs(4980) <= not(inputs(89)) or (inputs(1));
    layer0_outputs(4981) <= not(inputs(57)) or (inputs(184));
    layer0_outputs(4982) <= inputs(105);
    layer0_outputs(4983) <= (inputs(194)) and not (inputs(250));
    layer0_outputs(4984) <= not((inputs(81)) or (inputs(230)));
    layer0_outputs(4985) <= not(inputs(2)) or (inputs(32));
    layer0_outputs(4986) <= not((inputs(129)) or (inputs(1)));
    layer0_outputs(4987) <= (inputs(35)) and not (inputs(211));
    layer0_outputs(4988) <= not(inputs(108));
    layer0_outputs(4989) <= not(inputs(236));
    layer0_outputs(4990) <= not((inputs(238)) or (inputs(235)));
    layer0_outputs(4991) <= (inputs(145)) or (inputs(196));
    layer0_outputs(4992) <= inputs(54);
    layer0_outputs(4993) <= not(inputs(196)) or (inputs(159));
    layer0_outputs(4994) <= inputs(246);
    layer0_outputs(4995) <= not((inputs(117)) and (inputs(153)));
    layer0_outputs(4996) <= not(inputs(184)) or (inputs(143));
    layer0_outputs(4997) <= not((inputs(0)) or (inputs(188)));
    layer0_outputs(4998) <= inputs(7);
    layer0_outputs(4999) <= not(inputs(76));
    layer0_outputs(5000) <= (inputs(26)) and (inputs(12));
    layer0_outputs(5001) <= (inputs(157)) or (inputs(30));
    layer0_outputs(5002) <= (inputs(40)) or (inputs(128));
    layer0_outputs(5003) <= (inputs(206)) and not (inputs(117));
    layer0_outputs(5004) <= (inputs(114)) and not (inputs(86));
    layer0_outputs(5005) <= not(inputs(176)) or (inputs(58));
    layer0_outputs(5006) <= not(inputs(61)) or (inputs(21));
    layer0_outputs(5007) <= inputs(48);
    layer0_outputs(5008) <= (inputs(221)) xor (inputs(153));
    layer0_outputs(5009) <= not((inputs(148)) or (inputs(177)));
    layer0_outputs(5010) <= (inputs(216)) xor (inputs(184));
    layer0_outputs(5011) <= (inputs(236)) or (inputs(96));
    layer0_outputs(5012) <= (inputs(3)) or (inputs(121));
    layer0_outputs(5013) <= inputs(7);
    layer0_outputs(5014) <= (inputs(210)) or (inputs(109));
    layer0_outputs(5015) <= not((inputs(100)) or (inputs(173)));
    layer0_outputs(5016) <= (inputs(88)) xor (inputs(31));
    layer0_outputs(5017) <= not(inputs(56)) or (inputs(188));
    layer0_outputs(5018) <= (inputs(3)) xor (inputs(252));
    layer0_outputs(5019) <= not(inputs(117));
    layer0_outputs(5020) <= inputs(133);
    layer0_outputs(5021) <= (inputs(0)) and not (inputs(232));
    layer0_outputs(5022) <= (inputs(124)) or (inputs(161));
    layer0_outputs(5023) <= not((inputs(222)) xor (inputs(8)));
    layer0_outputs(5024) <= not(inputs(97));
    layer0_outputs(5025) <= (inputs(215)) and not (inputs(236));
    layer0_outputs(5026) <= inputs(58);
    layer0_outputs(5027) <= (inputs(248)) or (inputs(57));
    layer0_outputs(5028) <= not((inputs(187)) or (inputs(81)));
    layer0_outputs(5029) <= (inputs(105)) and not (inputs(197));
    layer0_outputs(5030) <= (inputs(103)) xor (inputs(148));
    layer0_outputs(5031) <= inputs(148);
    layer0_outputs(5032) <= (inputs(251)) and not (inputs(191));
    layer0_outputs(5033) <= not((inputs(40)) or (inputs(125)));
    layer0_outputs(5034) <= (inputs(165)) xor (inputs(151));
    layer0_outputs(5035) <= inputs(198);
    layer0_outputs(5036) <= inputs(120);
    layer0_outputs(5037) <= inputs(76);
    layer0_outputs(5038) <= (inputs(8)) and (inputs(253));
    layer0_outputs(5039) <= not(inputs(161)) or (inputs(97));
    layer0_outputs(5040) <= not(inputs(96));
    layer0_outputs(5041) <= not((inputs(49)) xor (inputs(26)));
    layer0_outputs(5042) <= not(inputs(167));
    layer0_outputs(5043) <= (inputs(88)) or (inputs(64));
    layer0_outputs(5044) <= (inputs(42)) or (inputs(46));
    layer0_outputs(5045) <= not(inputs(68)) or (inputs(164));
    layer0_outputs(5046) <= not(inputs(229)) or (inputs(111));
    layer0_outputs(5047) <= (inputs(180)) or (inputs(121));
    layer0_outputs(5048) <= (inputs(237)) xor (inputs(146));
    layer0_outputs(5049) <= not((inputs(207)) or (inputs(37)));
    layer0_outputs(5050) <= not(inputs(49)) or (inputs(92));
    layer0_outputs(5051) <= (inputs(73)) or (inputs(89));
    layer0_outputs(5052) <= (inputs(117)) and not (inputs(158));
    layer0_outputs(5053) <= (inputs(126)) or (inputs(155));
    layer0_outputs(5054) <= inputs(100);
    layer0_outputs(5055) <= '0';
    layer0_outputs(5056) <= (inputs(73)) and not (inputs(160));
    layer0_outputs(5057) <= (inputs(231)) or (inputs(61));
    layer0_outputs(5058) <= (inputs(254)) or (inputs(37));
    layer0_outputs(5059) <= not(inputs(98));
    layer0_outputs(5060) <= inputs(18);
    layer0_outputs(5061) <= (inputs(145)) and not (inputs(42));
    layer0_outputs(5062) <= (inputs(25)) or (inputs(177));
    layer0_outputs(5063) <= inputs(45);
    layer0_outputs(5064) <= inputs(166);
    layer0_outputs(5065) <= not((inputs(248)) or (inputs(69)));
    layer0_outputs(5066) <= (inputs(72)) or (inputs(95));
    layer0_outputs(5067) <= not(inputs(174)) or (inputs(172));
    layer0_outputs(5068) <= inputs(3);
    layer0_outputs(5069) <= inputs(16);
    layer0_outputs(5070) <= not(inputs(59)) or (inputs(173));
    layer0_outputs(5071) <= not((inputs(156)) or (inputs(80)));
    layer0_outputs(5072) <= not((inputs(66)) xor (inputs(9)));
    layer0_outputs(5073) <= inputs(68);
    layer0_outputs(5074) <= (inputs(38)) or (inputs(10));
    layer0_outputs(5075) <= inputs(39);
    layer0_outputs(5076) <= not((inputs(31)) or (inputs(21)));
    layer0_outputs(5077) <= (inputs(4)) and not (inputs(4));
    layer0_outputs(5078) <= (inputs(55)) or (inputs(75));
    layer0_outputs(5079) <= not(inputs(97)) or (inputs(255));
    layer0_outputs(5080) <= '1';
    layer0_outputs(5081) <= (inputs(38)) or (inputs(71));
    layer0_outputs(5082) <= inputs(250);
    layer0_outputs(5083) <= not(inputs(180)) or (inputs(124));
    layer0_outputs(5084) <= not((inputs(212)) or (inputs(43)));
    layer0_outputs(5085) <= '1';
    layer0_outputs(5086) <= not((inputs(57)) or (inputs(113)));
    layer0_outputs(5087) <= not(inputs(101));
    layer0_outputs(5088) <= not(inputs(42));
    layer0_outputs(5089) <= inputs(52);
    layer0_outputs(5090) <= not((inputs(157)) xor (inputs(105)));
    layer0_outputs(5091) <= not((inputs(165)) or (inputs(2)));
    layer0_outputs(5092) <= not(inputs(156));
    layer0_outputs(5093) <= not((inputs(89)) xor (inputs(196)));
    layer0_outputs(5094) <= (inputs(147)) and not (inputs(63));
    layer0_outputs(5095) <= not(inputs(213));
    layer0_outputs(5096) <= not(inputs(134)) or (inputs(18));
    layer0_outputs(5097) <= inputs(245);
    layer0_outputs(5098) <= not((inputs(112)) or (inputs(169)));
    layer0_outputs(5099) <= inputs(205);
    layer0_outputs(5100) <= not(inputs(117)) or (inputs(149));
    layer0_outputs(5101) <= not(inputs(15));
    layer0_outputs(5102) <= (inputs(217)) or (inputs(224));
    layer0_outputs(5103) <= inputs(149);
    layer0_outputs(5104) <= not((inputs(183)) or (inputs(133)));
    layer0_outputs(5105) <= inputs(87);
    layer0_outputs(5106) <= not((inputs(114)) or (inputs(152)));
    layer0_outputs(5107) <= not((inputs(83)) xor (inputs(204)));
    layer0_outputs(5108) <= (inputs(51)) and not (inputs(71));
    layer0_outputs(5109) <= not(inputs(254));
    layer0_outputs(5110) <= (inputs(180)) xor (inputs(158));
    layer0_outputs(5111) <= (inputs(219)) xor (inputs(105));
    layer0_outputs(5112) <= not((inputs(186)) or (inputs(193)));
    layer0_outputs(5113) <= not(inputs(247)) or (inputs(43));
    layer0_outputs(5114) <= not(inputs(116));
    layer0_outputs(5115) <= not(inputs(219)) or (inputs(43));
    layer0_outputs(5116) <= not(inputs(22)) or (inputs(175));
    layer0_outputs(5117) <= not((inputs(235)) or (inputs(3)));
    layer0_outputs(5118) <= not((inputs(27)) or (inputs(46)));
    layer0_outputs(5119) <= not(inputs(91));
    layer0_outputs(5120) <= inputs(132);
    layer0_outputs(5121) <= not(inputs(83));
    layer0_outputs(5122) <= (inputs(143)) or (inputs(19));
    layer0_outputs(5123) <= not((inputs(19)) xor (inputs(221)));
    layer0_outputs(5124) <= not(inputs(47)) or (inputs(145));
    layer0_outputs(5125) <= not(inputs(132));
    layer0_outputs(5126) <= inputs(73);
    layer0_outputs(5127) <= inputs(167);
    layer0_outputs(5128) <= (inputs(10)) and not (inputs(236));
    layer0_outputs(5129) <= not(inputs(136));
    layer0_outputs(5130) <= not((inputs(252)) and (inputs(185)));
    layer0_outputs(5131) <= not((inputs(103)) or (inputs(161)));
    layer0_outputs(5132) <= (inputs(33)) and not (inputs(94));
    layer0_outputs(5133) <= inputs(58);
    layer0_outputs(5134) <= inputs(71);
    layer0_outputs(5135) <= not((inputs(54)) or (inputs(163)));
    layer0_outputs(5136) <= (inputs(137)) and not (inputs(118));
    layer0_outputs(5137) <= not(inputs(219)) or (inputs(136));
    layer0_outputs(5138) <= not(inputs(115));
    layer0_outputs(5139) <= (inputs(192)) or (inputs(144));
    layer0_outputs(5140) <= not(inputs(91));
    layer0_outputs(5141) <= not(inputs(122));
    layer0_outputs(5142) <= inputs(95);
    layer0_outputs(5143) <= (inputs(255)) or (inputs(28));
    layer0_outputs(5144) <= not(inputs(235)) or (inputs(141));
    layer0_outputs(5145) <= not((inputs(166)) and (inputs(205)));
    layer0_outputs(5146) <= inputs(90);
    layer0_outputs(5147) <= not(inputs(233)) or (inputs(127));
    layer0_outputs(5148) <= not(inputs(161)) or (inputs(46));
    layer0_outputs(5149) <= (inputs(39)) and not (inputs(117));
    layer0_outputs(5150) <= inputs(103);
    layer0_outputs(5151) <= inputs(205);
    layer0_outputs(5152) <= (inputs(252)) or (inputs(180));
    layer0_outputs(5153) <= not(inputs(88)) or (inputs(32));
    layer0_outputs(5154) <= not(inputs(232));
    layer0_outputs(5155) <= (inputs(247)) and not (inputs(223));
    layer0_outputs(5156) <= not((inputs(94)) or (inputs(170)));
    layer0_outputs(5157) <= (inputs(74)) or (inputs(131));
    layer0_outputs(5158) <= inputs(222);
    layer0_outputs(5159) <= not(inputs(61));
    layer0_outputs(5160) <= (inputs(102)) or (inputs(247));
    layer0_outputs(5161) <= not(inputs(234)) or (inputs(36));
    layer0_outputs(5162) <= not(inputs(210));
    layer0_outputs(5163) <= (inputs(28)) xor (inputs(91));
    layer0_outputs(5164) <= not(inputs(108)) or (inputs(83));
    layer0_outputs(5165) <= (inputs(71)) xor (inputs(114));
    layer0_outputs(5166) <= not((inputs(48)) or (inputs(210)));
    layer0_outputs(5167) <= inputs(118);
    layer0_outputs(5168) <= inputs(167);
    layer0_outputs(5169) <= not(inputs(211));
    layer0_outputs(5170) <= not(inputs(156));
    layer0_outputs(5171) <= not(inputs(102)) or (inputs(48));
    layer0_outputs(5172) <= inputs(78);
    layer0_outputs(5173) <= inputs(129);
    layer0_outputs(5174) <= (inputs(18)) or (inputs(255));
    layer0_outputs(5175) <= not((inputs(156)) or (inputs(93)));
    layer0_outputs(5176) <= (inputs(147)) xor (inputs(50));
    layer0_outputs(5177) <= not((inputs(152)) xor (inputs(106)));
    layer0_outputs(5178) <= (inputs(10)) or (inputs(234));
    layer0_outputs(5179) <= (inputs(37)) or (inputs(122));
    layer0_outputs(5180) <= not((inputs(36)) or (inputs(229)));
    layer0_outputs(5181) <= not((inputs(203)) or (inputs(35)));
    layer0_outputs(5182) <= inputs(194);
    layer0_outputs(5183) <= not(inputs(253));
    layer0_outputs(5184) <= not((inputs(68)) xor (inputs(255)));
    layer0_outputs(5185) <= inputs(152);
    layer0_outputs(5186) <= inputs(51);
    layer0_outputs(5187) <= inputs(34);
    layer0_outputs(5188) <= (inputs(126)) or (inputs(88));
    layer0_outputs(5189) <= inputs(247);
    layer0_outputs(5190) <= inputs(103);
    layer0_outputs(5191) <= not(inputs(226)) or (inputs(52));
    layer0_outputs(5192) <= inputs(119);
    layer0_outputs(5193) <= not((inputs(197)) and (inputs(3)));
    layer0_outputs(5194) <= (inputs(206)) or (inputs(34));
    layer0_outputs(5195) <= not(inputs(166)) or (inputs(54));
    layer0_outputs(5196) <= (inputs(168)) xor (inputs(31));
    layer0_outputs(5197) <= (inputs(140)) or (inputs(48));
    layer0_outputs(5198) <= not((inputs(161)) xor (inputs(34)));
    layer0_outputs(5199) <= not(inputs(177));
    layer0_outputs(5200) <= not(inputs(164)) or (inputs(255));
    layer0_outputs(5201) <= inputs(38);
    layer0_outputs(5202) <= not(inputs(213)) or (inputs(30));
    layer0_outputs(5203) <= (inputs(239)) and (inputs(50));
    layer0_outputs(5204) <= not((inputs(68)) or (inputs(60)));
    layer0_outputs(5205) <= not((inputs(15)) and (inputs(52)));
    layer0_outputs(5206) <= not(inputs(68));
    layer0_outputs(5207) <= (inputs(135)) or (inputs(251));
    layer0_outputs(5208) <= not(inputs(176));
    layer0_outputs(5209) <= (inputs(87)) xor (inputs(100));
    layer0_outputs(5210) <= (inputs(118)) or (inputs(47));
    layer0_outputs(5211) <= inputs(100);
    layer0_outputs(5212) <= inputs(124);
    layer0_outputs(5213) <= not(inputs(186)) or (inputs(44));
    layer0_outputs(5214) <= inputs(254);
    layer0_outputs(5215) <= (inputs(158)) or (inputs(154));
    layer0_outputs(5216) <= (inputs(59)) or (inputs(181));
    layer0_outputs(5217) <= inputs(82);
    layer0_outputs(5218) <= inputs(191);
    layer0_outputs(5219) <= inputs(181);
    layer0_outputs(5220) <= not(inputs(123));
    layer0_outputs(5221) <= (inputs(182)) or (inputs(15));
    layer0_outputs(5222) <= (inputs(217)) and not (inputs(128));
    layer0_outputs(5223) <= (inputs(102)) and not (inputs(173));
    layer0_outputs(5224) <= (inputs(90)) and not (inputs(174));
    layer0_outputs(5225) <= not(inputs(24));
    layer0_outputs(5226) <= (inputs(75)) or (inputs(145));
    layer0_outputs(5227) <= not(inputs(226));
    layer0_outputs(5228) <= (inputs(43)) and not (inputs(202));
    layer0_outputs(5229) <= (inputs(175)) and (inputs(109));
    layer0_outputs(5230) <= (inputs(45)) and not (inputs(111));
    layer0_outputs(5231) <= not((inputs(70)) and (inputs(86)));
    layer0_outputs(5232) <= not((inputs(210)) or (inputs(75)));
    layer0_outputs(5233) <= inputs(194);
    layer0_outputs(5234) <= (inputs(7)) and not (inputs(125));
    layer0_outputs(5235) <= (inputs(39)) and not (inputs(203));
    layer0_outputs(5236) <= not(inputs(194));
    layer0_outputs(5237) <= not(inputs(22));
    layer0_outputs(5238) <= not((inputs(221)) xor (inputs(212)));
    layer0_outputs(5239) <= not(inputs(116)) or (inputs(20));
    layer0_outputs(5240) <= (inputs(30)) or (inputs(82));
    layer0_outputs(5241) <= inputs(213);
    layer0_outputs(5242) <= (inputs(11)) and not (inputs(201));
    layer0_outputs(5243) <= not(inputs(34));
    layer0_outputs(5244) <= inputs(197);
    layer0_outputs(5245) <= '1';
    layer0_outputs(5246) <= not(inputs(102));
    layer0_outputs(5247) <= '0';
    layer0_outputs(5248) <= inputs(34);
    layer0_outputs(5249) <= '1';
    layer0_outputs(5250) <= not((inputs(158)) or (inputs(173)));
    layer0_outputs(5251) <= (inputs(236)) or (inputs(40));
    layer0_outputs(5252) <= (inputs(190)) xor (inputs(116));
    layer0_outputs(5253) <= not(inputs(247));
    layer0_outputs(5254) <= not((inputs(222)) xor (inputs(227)));
    layer0_outputs(5255) <= (inputs(219)) and not (inputs(160));
    layer0_outputs(5256) <= not((inputs(253)) or (inputs(55)));
    layer0_outputs(5257) <= (inputs(246)) or (inputs(57));
    layer0_outputs(5258) <= (inputs(120)) and (inputs(68));
    layer0_outputs(5259) <= (inputs(121)) or (inputs(148));
    layer0_outputs(5260) <= (inputs(159)) xor (inputs(123));
    layer0_outputs(5261) <= not(inputs(23));
    layer0_outputs(5262) <= (inputs(117)) and not (inputs(112));
    layer0_outputs(5263) <= inputs(139);
    layer0_outputs(5264) <= not(inputs(214)) or (inputs(221));
    layer0_outputs(5265) <= not((inputs(204)) or (inputs(200)));
    layer0_outputs(5266) <= not(inputs(182));
    layer0_outputs(5267) <= not(inputs(97)) or (inputs(224));
    layer0_outputs(5268) <= not(inputs(211));
    layer0_outputs(5269) <= not(inputs(67)) or (inputs(56));
    layer0_outputs(5270) <= not(inputs(35));
    layer0_outputs(5271) <= not((inputs(59)) or (inputs(154)));
    layer0_outputs(5272) <= not(inputs(129));
    layer0_outputs(5273) <= (inputs(143)) or (inputs(144));
    layer0_outputs(5274) <= not(inputs(248)) or (inputs(61));
    layer0_outputs(5275) <= not(inputs(64)) or (inputs(192));
    layer0_outputs(5276) <= (inputs(188)) xor (inputs(195));
    layer0_outputs(5277) <= not((inputs(121)) and (inputs(123)));
    layer0_outputs(5278) <= inputs(165);
    layer0_outputs(5279) <= not(inputs(6));
    layer0_outputs(5280) <= (inputs(82)) and (inputs(233));
    layer0_outputs(5281) <= not(inputs(84)) or (inputs(223));
    layer0_outputs(5282) <= (inputs(26)) and (inputs(203));
    layer0_outputs(5283) <= not((inputs(33)) or (inputs(60)));
    layer0_outputs(5284) <= (inputs(183)) and not (inputs(16));
    layer0_outputs(5285) <= (inputs(233)) and not (inputs(33));
    layer0_outputs(5286) <= (inputs(208)) or (inputs(241));
    layer0_outputs(5287) <= (inputs(127)) or (inputs(10));
    layer0_outputs(5288) <= not(inputs(140)) or (inputs(253));
    layer0_outputs(5289) <= not((inputs(58)) or (inputs(2)));
    layer0_outputs(5290) <= (inputs(170)) or (inputs(142));
    layer0_outputs(5291) <= not((inputs(199)) or (inputs(151)));
    layer0_outputs(5292) <= not((inputs(135)) xor (inputs(173)));
    layer0_outputs(5293) <= not(inputs(195)) or (inputs(17));
    layer0_outputs(5294) <= not(inputs(187)) or (inputs(0));
    layer0_outputs(5295) <= not(inputs(207));
    layer0_outputs(5296) <= not(inputs(183));
    layer0_outputs(5297) <= not(inputs(68)) or (inputs(235));
    layer0_outputs(5298) <= not((inputs(236)) or (inputs(33)));
    layer0_outputs(5299) <= not(inputs(120)) or (inputs(85));
    layer0_outputs(5300) <= (inputs(231)) and not (inputs(170));
    layer0_outputs(5301) <= inputs(85);
    layer0_outputs(5302) <= not(inputs(87));
    layer0_outputs(5303) <= not(inputs(104));
    layer0_outputs(5304) <= not(inputs(144)) or (inputs(221));
    layer0_outputs(5305) <= (inputs(189)) and not (inputs(29));
    layer0_outputs(5306) <= (inputs(167)) xor (inputs(74));
    layer0_outputs(5307) <= (inputs(131)) and not (inputs(250));
    layer0_outputs(5308) <= (inputs(49)) xor (inputs(252));
    layer0_outputs(5309) <= inputs(17);
    layer0_outputs(5310) <= inputs(148);
    layer0_outputs(5311) <= inputs(200);
    layer0_outputs(5312) <= (inputs(215)) and not (inputs(135));
    layer0_outputs(5313) <= (inputs(115)) or (inputs(101));
    layer0_outputs(5314) <= (inputs(84)) and not (inputs(254));
    layer0_outputs(5315) <= (inputs(225)) and not (inputs(187));
    layer0_outputs(5316) <= not((inputs(177)) xor (inputs(37)));
    layer0_outputs(5317) <= (inputs(213)) and (inputs(131));
    layer0_outputs(5318) <= inputs(191);
    layer0_outputs(5319) <= not(inputs(62)) or (inputs(254));
    layer0_outputs(5320) <= (inputs(237)) and not (inputs(43));
    layer0_outputs(5321) <= (inputs(248)) or (inputs(51));
    layer0_outputs(5322) <= not((inputs(82)) or (inputs(73)));
    layer0_outputs(5323) <= inputs(67);
    layer0_outputs(5324) <= '1';
    layer0_outputs(5325) <= not(inputs(149));
    layer0_outputs(5326) <= not(inputs(150)) or (inputs(18));
    layer0_outputs(5327) <= not(inputs(167));
    layer0_outputs(5328) <= (inputs(56)) and not (inputs(237));
    layer0_outputs(5329) <= inputs(102);
    layer0_outputs(5330) <= not(inputs(103));
    layer0_outputs(5331) <= not((inputs(71)) xor (inputs(201)));
    layer0_outputs(5332) <= not(inputs(39));
    layer0_outputs(5333) <= (inputs(55)) or (inputs(126));
    layer0_outputs(5334) <= not(inputs(245)) or (inputs(5));
    layer0_outputs(5335) <= inputs(40);
    layer0_outputs(5336) <= (inputs(195)) or (inputs(144));
    layer0_outputs(5337) <= (inputs(198)) xor (inputs(69));
    layer0_outputs(5338) <= not((inputs(88)) xor (inputs(216)));
    layer0_outputs(5339) <= (inputs(225)) or (inputs(196));
    layer0_outputs(5340) <= not(inputs(236)) or (inputs(157));
    layer0_outputs(5341) <= (inputs(142)) xor (inputs(177));
    layer0_outputs(5342) <= not(inputs(218));
    layer0_outputs(5343) <= inputs(36);
    layer0_outputs(5344) <= not(inputs(74));
    layer0_outputs(5345) <= (inputs(84)) or (inputs(129));
    layer0_outputs(5346) <= inputs(42);
    layer0_outputs(5347) <= not(inputs(234));
    layer0_outputs(5348) <= inputs(131);
    layer0_outputs(5349) <= inputs(229);
    layer0_outputs(5350) <= (inputs(199)) xor (inputs(198));
    layer0_outputs(5351) <= inputs(100);
    layer0_outputs(5352) <= inputs(188);
    layer0_outputs(5353) <= not((inputs(131)) or (inputs(3)));
    layer0_outputs(5354) <= (inputs(68)) and not (inputs(106));
    layer0_outputs(5355) <= (inputs(43)) and not (inputs(217));
    layer0_outputs(5356) <= (inputs(38)) or (inputs(225));
    layer0_outputs(5357) <= (inputs(254)) or (inputs(152));
    layer0_outputs(5358) <= not(inputs(145));
    layer0_outputs(5359) <= (inputs(11)) and not (inputs(212));
    layer0_outputs(5360) <= (inputs(52)) and not (inputs(113));
    layer0_outputs(5361) <= inputs(31);
    layer0_outputs(5362) <= (inputs(178)) or (inputs(152));
    layer0_outputs(5363) <= not((inputs(43)) and (inputs(211)));
    layer0_outputs(5364) <= not(inputs(6));
    layer0_outputs(5365) <= (inputs(71)) xor (inputs(66));
    layer0_outputs(5366) <= not(inputs(135)) or (inputs(249));
    layer0_outputs(5367) <= (inputs(72)) and not (inputs(155));
    layer0_outputs(5368) <= not((inputs(175)) xor (inputs(161)));
    layer0_outputs(5369) <= inputs(7);
    layer0_outputs(5370) <= not(inputs(114));
    layer0_outputs(5371) <= (inputs(227)) or (inputs(202));
    layer0_outputs(5372) <= not(inputs(41));
    layer0_outputs(5373) <= not(inputs(8)) or (inputs(28));
    layer0_outputs(5374) <= (inputs(84)) and not (inputs(196));
    layer0_outputs(5375) <= (inputs(63)) xor (inputs(199));
    layer0_outputs(5376) <= not((inputs(149)) or (inputs(29)));
    layer0_outputs(5377) <= (inputs(230)) and not (inputs(3));
    layer0_outputs(5378) <= inputs(107);
    layer0_outputs(5379) <= (inputs(101)) or (inputs(103));
    layer0_outputs(5380) <= not(inputs(135));
    layer0_outputs(5381) <= (inputs(240)) xor (inputs(55));
    layer0_outputs(5382) <= (inputs(63)) or (inputs(80));
    layer0_outputs(5383) <= (inputs(114)) or (inputs(142));
    layer0_outputs(5384) <= (inputs(17)) and not (inputs(14));
    layer0_outputs(5385) <= not((inputs(162)) or (inputs(191)));
    layer0_outputs(5386) <= inputs(20);
    layer0_outputs(5387) <= not((inputs(80)) or (inputs(188)));
    layer0_outputs(5388) <= (inputs(62)) and not (inputs(114));
    layer0_outputs(5389) <= not((inputs(98)) or (inputs(116)));
    layer0_outputs(5390) <= (inputs(234)) and not (inputs(178));
    layer0_outputs(5391) <= (inputs(41)) and not (inputs(235));
    layer0_outputs(5392) <= (inputs(203)) or (inputs(222));
    layer0_outputs(5393) <= not(inputs(129));
    layer0_outputs(5394) <= not(inputs(82)) or (inputs(16));
    layer0_outputs(5395) <= not((inputs(169)) or (inputs(135)));
    layer0_outputs(5396) <= not(inputs(59));
    layer0_outputs(5397) <= (inputs(174)) or (inputs(5));
    layer0_outputs(5398) <= (inputs(216)) or (inputs(218));
    layer0_outputs(5399) <= (inputs(208)) or (inputs(190));
    layer0_outputs(5400) <= not(inputs(71)) or (inputs(245));
    layer0_outputs(5401) <= not(inputs(7));
    layer0_outputs(5402) <= not(inputs(219));
    layer0_outputs(5403) <= (inputs(121)) xor (inputs(150));
    layer0_outputs(5404) <= not((inputs(179)) or (inputs(84)));
    layer0_outputs(5405) <= not(inputs(222)) or (inputs(170));
    layer0_outputs(5406) <= not((inputs(118)) or (inputs(201)));
    layer0_outputs(5407) <= (inputs(17)) or (inputs(222));
    layer0_outputs(5408) <= not(inputs(62));
    layer0_outputs(5409) <= (inputs(59)) and not (inputs(172));
    layer0_outputs(5410) <= '0';
    layer0_outputs(5411) <= not(inputs(85));
    layer0_outputs(5412) <= (inputs(168)) or (inputs(151));
    layer0_outputs(5413) <= (inputs(85)) xor (inputs(62));
    layer0_outputs(5414) <= not((inputs(10)) xor (inputs(57)));
    layer0_outputs(5415) <= not(inputs(40)) or (inputs(134));
    layer0_outputs(5416) <= not((inputs(81)) or (inputs(177)));
    layer0_outputs(5417) <= (inputs(247)) xor (inputs(190));
    layer0_outputs(5418) <= (inputs(114)) or (inputs(182));
    layer0_outputs(5419) <= inputs(8);
    layer0_outputs(5420) <= (inputs(31)) or (inputs(113));
    layer0_outputs(5421) <= inputs(188);
    layer0_outputs(5422) <= inputs(121);
    layer0_outputs(5423) <= inputs(40);
    layer0_outputs(5424) <= not(inputs(100));
    layer0_outputs(5425) <= (inputs(119)) xor (inputs(168));
    layer0_outputs(5426) <= not(inputs(43));
    layer0_outputs(5427) <= (inputs(185)) xor (inputs(82));
    layer0_outputs(5428) <= not((inputs(217)) or (inputs(158)));
    layer0_outputs(5429) <= (inputs(62)) and (inputs(146));
    layer0_outputs(5430) <= not(inputs(184));
    layer0_outputs(5431) <= not((inputs(175)) xor (inputs(150)));
    layer0_outputs(5432) <= not((inputs(31)) or (inputs(13)));
    layer0_outputs(5433) <= (inputs(9)) and not (inputs(253));
    layer0_outputs(5434) <= (inputs(5)) xor (inputs(42));
    layer0_outputs(5435) <= not((inputs(51)) or (inputs(55)));
    layer0_outputs(5436) <= (inputs(195)) and not (inputs(100));
    layer0_outputs(5437) <= (inputs(197)) or (inputs(93));
    layer0_outputs(5438) <= not(inputs(133)) or (inputs(6));
    layer0_outputs(5439) <= not((inputs(108)) or (inputs(197)));
    layer0_outputs(5440) <= not((inputs(144)) and (inputs(175)));
    layer0_outputs(5441) <= (inputs(140)) and not (inputs(160));
    layer0_outputs(5442) <= not(inputs(33));
    layer0_outputs(5443) <= (inputs(60)) xor (inputs(204));
    layer0_outputs(5444) <= not((inputs(89)) or (inputs(96)));
    layer0_outputs(5445) <= (inputs(89)) and not (inputs(123));
    layer0_outputs(5446) <= not((inputs(204)) or (inputs(192)));
    layer0_outputs(5447) <= (inputs(187)) or (inputs(223));
    layer0_outputs(5448) <= not(inputs(34));
    layer0_outputs(5449) <= (inputs(201)) or (inputs(167));
    layer0_outputs(5450) <= inputs(59);
    layer0_outputs(5451) <= (inputs(53)) or (inputs(165));
    layer0_outputs(5452) <= inputs(53);
    layer0_outputs(5453) <= not(inputs(173)) or (inputs(98));
    layer0_outputs(5454) <= not((inputs(193)) and (inputs(193)));
    layer0_outputs(5455) <= inputs(103);
    layer0_outputs(5456) <= not(inputs(50));
    layer0_outputs(5457) <= not(inputs(25));
    layer0_outputs(5458) <= not((inputs(228)) xor (inputs(197)));
    layer0_outputs(5459) <= '0';
    layer0_outputs(5460) <= not(inputs(53));
    layer0_outputs(5461) <= (inputs(168)) and (inputs(31));
    layer0_outputs(5462) <= not((inputs(83)) or (inputs(131)));
    layer0_outputs(5463) <= (inputs(88)) and (inputs(119));
    layer0_outputs(5464) <= not(inputs(138)) or (inputs(180));
    layer0_outputs(5465) <= inputs(71);
    layer0_outputs(5466) <= not(inputs(107));
    layer0_outputs(5467) <= (inputs(16)) and not (inputs(201));
    layer0_outputs(5468) <= inputs(26);
    layer0_outputs(5469) <= not(inputs(40));
    layer0_outputs(5470) <= '0';
    layer0_outputs(5471) <= '0';
    layer0_outputs(5472) <= not((inputs(126)) or (inputs(44)));
    layer0_outputs(5473) <= (inputs(56)) or (inputs(244));
    layer0_outputs(5474) <= not(inputs(46));
    layer0_outputs(5475) <= (inputs(236)) and not (inputs(126));
    layer0_outputs(5476) <= not(inputs(103));
    layer0_outputs(5477) <= not(inputs(24)) or (inputs(126));
    layer0_outputs(5478) <= (inputs(168)) and not (inputs(91));
    layer0_outputs(5479) <= not((inputs(3)) or (inputs(66)));
    layer0_outputs(5480) <= not((inputs(230)) or (inputs(94)));
    layer0_outputs(5481) <= not((inputs(83)) xor (inputs(113)));
    layer0_outputs(5482) <= (inputs(83)) xor (inputs(188));
    layer0_outputs(5483) <= not((inputs(20)) or (inputs(220)));
    layer0_outputs(5484) <= inputs(101);
    layer0_outputs(5485) <= not(inputs(153)) or (inputs(208));
    layer0_outputs(5486) <= (inputs(177)) or (inputs(119));
    layer0_outputs(5487) <= not(inputs(181));
    layer0_outputs(5488) <= (inputs(231)) and not (inputs(2));
    layer0_outputs(5489) <= (inputs(251)) or (inputs(53));
    layer0_outputs(5490) <= not(inputs(166));
    layer0_outputs(5491) <= not((inputs(222)) or (inputs(151)));
    layer0_outputs(5492) <= (inputs(114)) xor (inputs(83));
    layer0_outputs(5493) <= (inputs(183)) and not (inputs(94));
    layer0_outputs(5494) <= not(inputs(167));
    layer0_outputs(5495) <= not((inputs(98)) or (inputs(98)));
    layer0_outputs(5496) <= not(inputs(2));
    layer0_outputs(5497) <= (inputs(215)) or (inputs(185));
    layer0_outputs(5498) <= not(inputs(119));
    layer0_outputs(5499) <= (inputs(76)) xor (inputs(192));
    layer0_outputs(5500) <= inputs(44);
    layer0_outputs(5501) <= not((inputs(170)) xor (inputs(120)));
    layer0_outputs(5502) <= not(inputs(41)) or (inputs(252));
    layer0_outputs(5503) <= (inputs(7)) or (inputs(66));
    layer0_outputs(5504) <= not(inputs(210));
    layer0_outputs(5505) <= (inputs(31)) or (inputs(8));
    layer0_outputs(5506) <= (inputs(132)) or (inputs(130));
    layer0_outputs(5507) <= not((inputs(242)) or (inputs(127)));
    layer0_outputs(5508) <= inputs(58);
    layer0_outputs(5509) <= inputs(186);
    layer0_outputs(5510) <= not(inputs(212)) or (inputs(102));
    layer0_outputs(5511) <= (inputs(220)) xor (inputs(188));
    layer0_outputs(5512) <= not((inputs(130)) xor (inputs(96)));
    layer0_outputs(5513) <= (inputs(114)) and not (inputs(207));
    layer0_outputs(5514) <= not(inputs(34));
    layer0_outputs(5515) <= not(inputs(54));
    layer0_outputs(5516) <= not(inputs(190));
    layer0_outputs(5517) <= (inputs(53)) and not (inputs(160));
    layer0_outputs(5518) <= not((inputs(132)) and (inputs(202)));
    layer0_outputs(5519) <= inputs(146);
    layer0_outputs(5520) <= not((inputs(121)) xor (inputs(140)));
    layer0_outputs(5521) <= (inputs(44)) and not (inputs(238));
    layer0_outputs(5522) <= (inputs(74)) and not (inputs(118));
    layer0_outputs(5523) <= not(inputs(175)) or (inputs(28));
    layer0_outputs(5524) <= inputs(29);
    layer0_outputs(5525) <= inputs(252);
    layer0_outputs(5526) <= not(inputs(200)) or (inputs(32));
    layer0_outputs(5527) <= (inputs(129)) or (inputs(195));
    layer0_outputs(5528) <= (inputs(72)) and not (inputs(216));
    layer0_outputs(5529) <= (inputs(203)) xor (inputs(139));
    layer0_outputs(5530) <= not(inputs(18));
    layer0_outputs(5531) <= not((inputs(79)) xor (inputs(231)));
    layer0_outputs(5532) <= not(inputs(27)) or (inputs(157));
    layer0_outputs(5533) <= (inputs(204)) or (inputs(203));
    layer0_outputs(5534) <= not((inputs(212)) xor (inputs(142)));
    layer0_outputs(5535) <= not(inputs(68)) or (inputs(207));
    layer0_outputs(5536) <= (inputs(215)) and not (inputs(36));
    layer0_outputs(5537) <= (inputs(78)) xor (inputs(231));
    layer0_outputs(5538) <= not(inputs(179)) or (inputs(48));
    layer0_outputs(5539) <= not(inputs(95));
    layer0_outputs(5540) <= (inputs(241)) xor (inputs(119));
    layer0_outputs(5541) <= (inputs(146)) xor (inputs(49));
    layer0_outputs(5542) <= inputs(162);
    layer0_outputs(5543) <= not((inputs(152)) or (inputs(180)));
    layer0_outputs(5544) <= (inputs(159)) or (inputs(195));
    layer0_outputs(5545) <= inputs(220);
    layer0_outputs(5546) <= not(inputs(184)) or (inputs(16));
    layer0_outputs(5547) <= inputs(39);
    layer0_outputs(5548) <= (inputs(209)) and not (inputs(156));
    layer0_outputs(5549) <= not((inputs(179)) or (inputs(168)));
    layer0_outputs(5550) <= not((inputs(71)) or (inputs(78)));
    layer0_outputs(5551) <= inputs(244);
    layer0_outputs(5552) <= '0';
    layer0_outputs(5553) <= (inputs(23)) xor (inputs(228));
    layer0_outputs(5554) <= not(inputs(154)) or (inputs(227));
    layer0_outputs(5555) <= (inputs(213)) and not (inputs(107));
    layer0_outputs(5556) <= inputs(93);
    layer0_outputs(5557) <= not(inputs(194));
    layer0_outputs(5558) <= '0';
    layer0_outputs(5559) <= (inputs(212)) and not (inputs(128));
    layer0_outputs(5560) <= (inputs(233)) and not (inputs(17));
    layer0_outputs(5561) <= inputs(188);
    layer0_outputs(5562) <= (inputs(163)) and not (inputs(48));
    layer0_outputs(5563) <= (inputs(127)) and (inputs(127));
    layer0_outputs(5564) <= inputs(42);
    layer0_outputs(5565) <= inputs(197);
    layer0_outputs(5566) <= not((inputs(131)) xor (inputs(22)));
    layer0_outputs(5567) <= not((inputs(161)) or (inputs(15)));
    layer0_outputs(5568) <= not(inputs(19));
    layer0_outputs(5569) <= (inputs(82)) and not (inputs(222));
    layer0_outputs(5570) <= (inputs(134)) and not (inputs(93));
    layer0_outputs(5571) <= inputs(106);
    layer0_outputs(5572) <= inputs(142);
    layer0_outputs(5573) <= inputs(121);
    layer0_outputs(5574) <= inputs(40);
    layer0_outputs(5575) <= not((inputs(192)) or (inputs(215)));
    layer0_outputs(5576) <= not((inputs(242)) or (inputs(65)));
    layer0_outputs(5577) <= (inputs(63)) or (inputs(246));
    layer0_outputs(5578) <= not((inputs(211)) or (inputs(254)));
    layer0_outputs(5579) <= (inputs(43)) and not (inputs(192));
    layer0_outputs(5580) <= not((inputs(49)) or (inputs(109)));
    layer0_outputs(5581) <= (inputs(192)) xor (inputs(253));
    layer0_outputs(5582) <= not((inputs(132)) xor (inputs(168)));
    layer0_outputs(5583) <= not(inputs(131));
    layer0_outputs(5584) <= not(inputs(163));
    layer0_outputs(5585) <= '0';
    layer0_outputs(5586) <= not(inputs(246));
    layer0_outputs(5587) <= not(inputs(121));
    layer0_outputs(5588) <= inputs(54);
    layer0_outputs(5589) <= not(inputs(197)) or (inputs(203));
    layer0_outputs(5590) <= not((inputs(143)) or (inputs(238)));
    layer0_outputs(5591) <= (inputs(38)) and not (inputs(232));
    layer0_outputs(5592) <= (inputs(32)) xor (inputs(158));
    layer0_outputs(5593) <= not(inputs(236));
    layer0_outputs(5594) <= '0';
    layer0_outputs(5595) <= (inputs(60)) and not (inputs(14));
    layer0_outputs(5596) <= (inputs(214)) and not (inputs(54));
    layer0_outputs(5597) <= inputs(145);
    layer0_outputs(5598) <= inputs(141);
    layer0_outputs(5599) <= (inputs(22)) and not (inputs(15));
    layer0_outputs(5600) <= (inputs(29)) and not (inputs(70));
    layer0_outputs(5601) <= (inputs(183)) and not (inputs(113));
    layer0_outputs(5602) <= not(inputs(81));
    layer0_outputs(5603) <= inputs(106);
    layer0_outputs(5604) <= (inputs(231)) and (inputs(233));
    layer0_outputs(5605) <= inputs(215);
    layer0_outputs(5606) <= not(inputs(19)) or (inputs(189));
    layer0_outputs(5607) <= (inputs(15)) or (inputs(181));
    layer0_outputs(5608) <= (inputs(222)) or (inputs(215));
    layer0_outputs(5609) <= (inputs(31)) and not (inputs(110));
    layer0_outputs(5610) <= not(inputs(149));
    layer0_outputs(5611) <= not((inputs(132)) or (inputs(159)));
    layer0_outputs(5612) <= inputs(135);
    layer0_outputs(5613) <= inputs(232);
    layer0_outputs(5614) <= not(inputs(151)) or (inputs(28));
    layer0_outputs(5615) <= not((inputs(39)) and (inputs(69)));
    layer0_outputs(5616) <= inputs(45);
    layer0_outputs(5617) <= not(inputs(180)) or (inputs(57));
    layer0_outputs(5618) <= not(inputs(41));
    layer0_outputs(5619) <= not(inputs(104)) or (inputs(109));
    layer0_outputs(5620) <= not((inputs(12)) xor (inputs(37)));
    layer0_outputs(5621) <= (inputs(128)) or (inputs(117));
    layer0_outputs(5622) <= not(inputs(88)) or (inputs(182));
    layer0_outputs(5623) <= not((inputs(32)) or (inputs(227)));
    layer0_outputs(5624) <= not(inputs(203)) or (inputs(33));
    layer0_outputs(5625) <= not(inputs(228));
    layer0_outputs(5626) <= (inputs(155)) or (inputs(113));
    layer0_outputs(5627) <= (inputs(76)) or (inputs(63));
    layer0_outputs(5628) <= not(inputs(102));
    layer0_outputs(5629) <= not(inputs(156)) or (inputs(65));
    layer0_outputs(5630) <= not(inputs(234));
    layer0_outputs(5631) <= not(inputs(99)) or (inputs(212));
    layer0_outputs(5632) <= (inputs(163)) xor (inputs(206));
    layer0_outputs(5633) <= (inputs(205)) xor (inputs(231));
    layer0_outputs(5634) <= not((inputs(80)) and (inputs(13)));
    layer0_outputs(5635) <= (inputs(171)) or (inputs(158));
    layer0_outputs(5636) <= (inputs(164)) or (inputs(126));
    layer0_outputs(5637) <= not(inputs(98));
    layer0_outputs(5638) <= not(inputs(47));
    layer0_outputs(5639) <= not((inputs(2)) and (inputs(92)));
    layer0_outputs(5640) <= not((inputs(7)) or (inputs(110)));
    layer0_outputs(5641) <= not(inputs(109));
    layer0_outputs(5642) <= inputs(23);
    layer0_outputs(5643) <= (inputs(85)) or (inputs(211));
    layer0_outputs(5644) <= not((inputs(173)) xor (inputs(171)));
    layer0_outputs(5645) <= not((inputs(238)) or (inputs(48)));
    layer0_outputs(5646) <= not((inputs(129)) or (inputs(17)));
    layer0_outputs(5647) <= not(inputs(183));
    layer0_outputs(5648) <= (inputs(17)) and (inputs(207));
    layer0_outputs(5649) <= inputs(210);
    layer0_outputs(5650) <= (inputs(91)) and (inputs(196));
    layer0_outputs(5651) <= not(inputs(116));
    layer0_outputs(5652) <= (inputs(12)) or (inputs(32));
    layer0_outputs(5653) <= not((inputs(212)) or (inputs(213)));
    layer0_outputs(5654) <= not((inputs(46)) or (inputs(64)));
    layer0_outputs(5655) <= not(inputs(25)) or (inputs(4));
    layer0_outputs(5656) <= not(inputs(163));
    layer0_outputs(5657) <= (inputs(232)) and not (inputs(34));
    layer0_outputs(5658) <= not((inputs(10)) or (inputs(6)));
    layer0_outputs(5659) <= not(inputs(166));
    layer0_outputs(5660) <= inputs(226);
    layer0_outputs(5661) <= not((inputs(192)) or (inputs(230)));
    layer0_outputs(5662) <= not(inputs(41));
    layer0_outputs(5663) <= not(inputs(244));
    layer0_outputs(5664) <= not(inputs(34));
    layer0_outputs(5665) <= (inputs(41)) xor (inputs(70));
    layer0_outputs(5666) <= inputs(231);
    layer0_outputs(5667) <= inputs(76);
    layer0_outputs(5668) <= inputs(128);
    layer0_outputs(5669) <= not(inputs(218));
    layer0_outputs(5670) <= not(inputs(90));
    layer0_outputs(5671) <= not(inputs(201)) or (inputs(236));
    layer0_outputs(5672) <= (inputs(227)) or (inputs(253));
    layer0_outputs(5673) <= not(inputs(199));
    layer0_outputs(5674) <= not(inputs(10));
    layer0_outputs(5675) <= inputs(181);
    layer0_outputs(5676) <= not((inputs(155)) or (inputs(37)));
    layer0_outputs(5677) <= not((inputs(113)) xor (inputs(48)));
    layer0_outputs(5678) <= (inputs(235)) or (inputs(209));
    layer0_outputs(5679) <= not(inputs(141));
    layer0_outputs(5680) <= not((inputs(227)) xor (inputs(39)));
    layer0_outputs(5681) <= inputs(67);
    layer0_outputs(5682) <= not((inputs(22)) or (inputs(15)));
    layer0_outputs(5683) <= not(inputs(40));
    layer0_outputs(5684) <= inputs(2);
    layer0_outputs(5685) <= not(inputs(22));
    layer0_outputs(5686) <= inputs(171);
    layer0_outputs(5687) <= inputs(104);
    layer0_outputs(5688) <= (inputs(96)) or (inputs(123));
    layer0_outputs(5689) <= inputs(62);
    layer0_outputs(5690) <= not((inputs(182)) xor (inputs(73)));
    layer0_outputs(5691) <= not((inputs(5)) xor (inputs(10)));
    layer0_outputs(5692) <= not(inputs(209));
    layer0_outputs(5693) <= not((inputs(65)) or (inputs(224)));
    layer0_outputs(5694) <= not(inputs(47)) or (inputs(225));
    layer0_outputs(5695) <= not((inputs(42)) and (inputs(76)));
    layer0_outputs(5696) <= not(inputs(134)) or (inputs(127));
    layer0_outputs(5697) <= not((inputs(174)) or (inputs(211)));
    layer0_outputs(5698) <= inputs(68);
    layer0_outputs(5699) <= inputs(108);
    layer0_outputs(5700) <= not((inputs(225)) or (inputs(48)));
    layer0_outputs(5701) <= not(inputs(24));
    layer0_outputs(5702) <= not(inputs(134)) or (inputs(137));
    layer0_outputs(5703) <= (inputs(225)) and not (inputs(69));
    layer0_outputs(5704) <= (inputs(239)) xor (inputs(252));
    layer0_outputs(5705) <= not(inputs(68));
    layer0_outputs(5706) <= inputs(37);
    layer0_outputs(5707) <= not(inputs(25));
    layer0_outputs(5708) <= '1';
    layer0_outputs(5709) <= (inputs(117)) and not (inputs(64));
    layer0_outputs(5710) <= not(inputs(5));
    layer0_outputs(5711) <= (inputs(219)) or (inputs(239));
    layer0_outputs(5712) <= inputs(224);
    layer0_outputs(5713) <= inputs(208);
    layer0_outputs(5714) <= not((inputs(164)) xor (inputs(146)));
    layer0_outputs(5715) <= (inputs(138)) and not (inputs(112));
    layer0_outputs(5716) <= (inputs(52)) xor (inputs(135));
    layer0_outputs(5717) <= not((inputs(153)) xor (inputs(130)));
    layer0_outputs(5718) <= not((inputs(179)) or (inputs(245)));
    layer0_outputs(5719) <= not(inputs(186));
    layer0_outputs(5720) <= inputs(170);
    layer0_outputs(5721) <= (inputs(209)) xor (inputs(145));
    layer0_outputs(5722) <= (inputs(198)) xor (inputs(112));
    layer0_outputs(5723) <= not((inputs(186)) xor (inputs(120)));
    layer0_outputs(5724) <= not(inputs(95)) or (inputs(61));
    layer0_outputs(5725) <= not(inputs(115));
    layer0_outputs(5726) <= not((inputs(204)) or (inputs(171)));
    layer0_outputs(5727) <= not((inputs(163)) or (inputs(85)));
    layer0_outputs(5728) <= (inputs(72)) and (inputs(31));
    layer0_outputs(5729) <= (inputs(217)) and not (inputs(106));
    layer0_outputs(5730) <= not(inputs(77));
    layer0_outputs(5731) <= not((inputs(211)) or (inputs(196)));
    layer0_outputs(5732) <= not((inputs(221)) xor (inputs(172)));
    layer0_outputs(5733) <= (inputs(86)) or (inputs(101));
    layer0_outputs(5734) <= inputs(144);
    layer0_outputs(5735) <= inputs(232);
    layer0_outputs(5736) <= (inputs(174)) and not (inputs(96));
    layer0_outputs(5737) <= (inputs(73)) and (inputs(132));
    layer0_outputs(5738) <= inputs(209);
    layer0_outputs(5739) <= (inputs(63)) or (inputs(78));
    layer0_outputs(5740) <= inputs(83);
    layer0_outputs(5741) <= inputs(150);
    layer0_outputs(5742) <= (inputs(75)) and not (inputs(2));
    layer0_outputs(5743) <= not((inputs(193)) or (inputs(230)));
    layer0_outputs(5744) <= not(inputs(180)) or (inputs(190));
    layer0_outputs(5745) <= not(inputs(198)) or (inputs(197));
    layer0_outputs(5746) <= not(inputs(70));
    layer0_outputs(5747) <= not(inputs(8)) or (inputs(249));
    layer0_outputs(5748) <= inputs(129);
    layer0_outputs(5749) <= not((inputs(223)) or (inputs(91)));
    layer0_outputs(5750) <= '1';
    layer0_outputs(5751) <= not((inputs(157)) or (inputs(230)));
    layer0_outputs(5752) <= not(inputs(130));
    layer0_outputs(5753) <= not((inputs(30)) or (inputs(127)));
    layer0_outputs(5754) <= not((inputs(141)) or (inputs(101)));
    layer0_outputs(5755) <= not(inputs(136)) or (inputs(143));
    layer0_outputs(5756) <= (inputs(24)) and not (inputs(205));
    layer0_outputs(5757) <= (inputs(20)) and not (inputs(158));
    layer0_outputs(5758) <= inputs(90);
    layer0_outputs(5759) <= (inputs(83)) and not (inputs(242));
    layer0_outputs(5760) <= inputs(70);
    layer0_outputs(5761) <= inputs(101);
    layer0_outputs(5762) <= not(inputs(229));
    layer0_outputs(5763) <= not(inputs(164));
    layer0_outputs(5764) <= not((inputs(235)) xor (inputs(46)));
    layer0_outputs(5765) <= not(inputs(202));
    layer0_outputs(5766) <= not((inputs(121)) xor (inputs(111)));
    layer0_outputs(5767) <= inputs(138);
    layer0_outputs(5768) <= not(inputs(182));
    layer0_outputs(5769) <= not(inputs(235)) or (inputs(252));
    layer0_outputs(5770) <= not((inputs(251)) and (inputs(79)));
    layer0_outputs(5771) <= not(inputs(12)) or (inputs(242));
    layer0_outputs(5772) <= inputs(68);
    layer0_outputs(5773) <= (inputs(183)) xor (inputs(134));
    layer0_outputs(5774) <= (inputs(116)) and not (inputs(32));
    layer0_outputs(5775) <= (inputs(149)) or (inputs(162));
    layer0_outputs(5776) <= not(inputs(93)) or (inputs(238));
    layer0_outputs(5777) <= not((inputs(52)) and (inputs(51)));
    layer0_outputs(5778) <= (inputs(72)) xor (inputs(119));
    layer0_outputs(5779) <= (inputs(35)) xor (inputs(87));
    layer0_outputs(5780) <= not(inputs(4)) or (inputs(52));
    layer0_outputs(5781) <= inputs(105);
    layer0_outputs(5782) <= not((inputs(103)) or (inputs(239)));
    layer0_outputs(5783) <= not(inputs(130));
    layer0_outputs(5784) <= not(inputs(136));
    layer0_outputs(5785) <= not((inputs(211)) or (inputs(160)));
    layer0_outputs(5786) <= (inputs(73)) and not (inputs(220));
    layer0_outputs(5787) <= not(inputs(198)) or (inputs(133));
    layer0_outputs(5788) <= inputs(85);
    layer0_outputs(5789) <= inputs(244);
    layer0_outputs(5790) <= not(inputs(8)) or (inputs(191));
    layer0_outputs(5791) <= not((inputs(5)) or (inputs(9)));
    layer0_outputs(5792) <= not((inputs(189)) or (inputs(217)));
    layer0_outputs(5793) <= (inputs(143)) or (inputs(178));
    layer0_outputs(5794) <= (inputs(230)) and not (inputs(129));
    layer0_outputs(5795) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(5796) <= not((inputs(48)) xor (inputs(5)));
    layer0_outputs(5797) <= not(inputs(170)) or (inputs(176));
    layer0_outputs(5798) <= not(inputs(121)) or (inputs(35));
    layer0_outputs(5799) <= (inputs(210)) and not (inputs(122));
    layer0_outputs(5800) <= not((inputs(109)) or (inputs(16)));
    layer0_outputs(5801) <= inputs(151);
    layer0_outputs(5802) <= (inputs(193)) and not (inputs(128));
    layer0_outputs(5803) <= '0';
    layer0_outputs(5804) <= inputs(180);
    layer0_outputs(5805) <= not((inputs(195)) xor (inputs(111)));
    layer0_outputs(5806) <= (inputs(0)) xor (inputs(153));
    layer0_outputs(5807) <= not(inputs(233));
    layer0_outputs(5808) <= (inputs(204)) and not (inputs(144));
    layer0_outputs(5809) <= not(inputs(235)) or (inputs(63));
    layer0_outputs(5810) <= (inputs(195)) and not (inputs(255));
    layer0_outputs(5811) <= not((inputs(70)) xor (inputs(20)));
    layer0_outputs(5812) <= not((inputs(151)) xor (inputs(168)));
    layer0_outputs(5813) <= not(inputs(143));
    layer0_outputs(5814) <= (inputs(251)) and (inputs(218));
    layer0_outputs(5815) <= (inputs(156)) or (inputs(169));
    layer0_outputs(5816) <= inputs(180);
    layer0_outputs(5817) <= (inputs(234)) xor (inputs(248));
    layer0_outputs(5818) <= (inputs(205)) xor (inputs(170));
    layer0_outputs(5819) <= inputs(209);
    layer0_outputs(5820) <= not(inputs(129)) or (inputs(85));
    layer0_outputs(5821) <= (inputs(213)) and (inputs(215));
    layer0_outputs(5822) <= (inputs(27)) and not (inputs(233));
    layer0_outputs(5823) <= (inputs(169)) and not (inputs(117));
    layer0_outputs(5824) <= (inputs(19)) xor (inputs(109));
    layer0_outputs(5825) <= inputs(151);
    layer0_outputs(5826) <= (inputs(18)) or (inputs(32));
    layer0_outputs(5827) <= (inputs(168)) and not (inputs(35));
    layer0_outputs(5828) <= (inputs(141)) or (inputs(111));
    layer0_outputs(5829) <= not((inputs(84)) and (inputs(134)));
    layer0_outputs(5830) <= inputs(99);
    layer0_outputs(5831) <= inputs(17);
    layer0_outputs(5832) <= not((inputs(62)) or (inputs(76)));
    layer0_outputs(5833) <= not(inputs(179)) or (inputs(30));
    layer0_outputs(5834) <= (inputs(165)) xor (inputs(182));
    layer0_outputs(5835) <= (inputs(237)) or (inputs(167));
    layer0_outputs(5836) <= not(inputs(82));
    layer0_outputs(5837) <= not(inputs(194));
    layer0_outputs(5838) <= not((inputs(116)) xor (inputs(123)));
    layer0_outputs(5839) <= (inputs(42)) and not (inputs(242));
    layer0_outputs(5840) <= '1';
    layer0_outputs(5841) <= not((inputs(153)) or (inputs(178)));
    layer0_outputs(5842) <= (inputs(26)) xor (inputs(9));
    layer0_outputs(5843) <= not((inputs(164)) or (inputs(129)));
    layer0_outputs(5844) <= not(inputs(48));
    layer0_outputs(5845) <= inputs(13);
    layer0_outputs(5846) <= (inputs(25)) or (inputs(55));
    layer0_outputs(5847) <= not(inputs(106)) or (inputs(251));
    layer0_outputs(5848) <= not((inputs(170)) xor (inputs(108)));
    layer0_outputs(5849) <= not((inputs(196)) xor (inputs(47)));
    layer0_outputs(5850) <= (inputs(113)) or (inputs(205));
    layer0_outputs(5851) <= not((inputs(177)) and (inputs(160)));
    layer0_outputs(5852) <= not(inputs(149)) or (inputs(122));
    layer0_outputs(5853) <= (inputs(21)) and not (inputs(163));
    layer0_outputs(5854) <= not((inputs(79)) xor (inputs(4)));
    layer0_outputs(5855) <= (inputs(142)) or (inputs(190));
    layer0_outputs(5856) <= (inputs(134)) and not (inputs(172));
    layer0_outputs(5857) <= inputs(16);
    layer0_outputs(5858) <= not(inputs(32));
    layer0_outputs(5859) <= not((inputs(53)) xor (inputs(177)));
    layer0_outputs(5860) <= not(inputs(25)) or (inputs(95));
    layer0_outputs(5861) <= (inputs(51)) or (inputs(228));
    layer0_outputs(5862) <= not(inputs(28)) or (inputs(171));
    layer0_outputs(5863) <= not((inputs(248)) xor (inputs(121)));
    layer0_outputs(5864) <= (inputs(133)) and not (inputs(222));
    layer0_outputs(5865) <= not(inputs(50)) or (inputs(63));
    layer0_outputs(5866) <= inputs(176);
    layer0_outputs(5867) <= not((inputs(12)) and (inputs(142)));
    layer0_outputs(5868) <= (inputs(222)) xor (inputs(85));
    layer0_outputs(5869) <= (inputs(179)) xor (inputs(240));
    layer0_outputs(5870) <= not(inputs(247));
    layer0_outputs(5871) <= not(inputs(134)) or (inputs(197));
    layer0_outputs(5872) <= not(inputs(59));
    layer0_outputs(5873) <= not(inputs(157));
    layer0_outputs(5874) <= not(inputs(23));
    layer0_outputs(5875) <= (inputs(161)) xor (inputs(169));
    layer0_outputs(5876) <= inputs(188);
    layer0_outputs(5877) <= inputs(39);
    layer0_outputs(5878) <= (inputs(86)) xor (inputs(8));
    layer0_outputs(5879) <= not((inputs(183)) xor (inputs(230)));
    layer0_outputs(5880) <= not((inputs(141)) or (inputs(90)));
    layer0_outputs(5881) <= (inputs(142)) or (inputs(142));
    layer0_outputs(5882) <= (inputs(168)) and (inputs(93));
    layer0_outputs(5883) <= not(inputs(26));
    layer0_outputs(5884) <= not((inputs(227)) xor (inputs(130)));
    layer0_outputs(5885) <= not((inputs(159)) and (inputs(82)));
    layer0_outputs(5886) <= (inputs(96)) xor (inputs(92));
    layer0_outputs(5887) <= inputs(178);
    layer0_outputs(5888) <= not(inputs(180));
    layer0_outputs(5889) <= inputs(246);
    layer0_outputs(5890) <= (inputs(3)) and not (inputs(99));
    layer0_outputs(5891) <= (inputs(26)) and not (inputs(142));
    layer0_outputs(5892) <= not(inputs(170));
    layer0_outputs(5893) <= '1';
    layer0_outputs(5894) <= not(inputs(218));
    layer0_outputs(5895) <= (inputs(186)) and not (inputs(122));
    layer0_outputs(5896) <= inputs(241);
    layer0_outputs(5897) <= not((inputs(111)) or (inputs(147)));
    layer0_outputs(5898) <= inputs(65);
    layer0_outputs(5899) <= not(inputs(4));
    layer0_outputs(5900) <= inputs(121);
    layer0_outputs(5901) <= not(inputs(21)) or (inputs(127));
    layer0_outputs(5902) <= (inputs(160)) or (inputs(11));
    layer0_outputs(5903) <= not(inputs(201));
    layer0_outputs(5904) <= inputs(216);
    layer0_outputs(5905) <= inputs(248);
    layer0_outputs(5906) <= (inputs(106)) and not (inputs(178));
    layer0_outputs(5907) <= (inputs(234)) and not (inputs(128));
    layer0_outputs(5908) <= not((inputs(137)) and (inputs(139)));
    layer0_outputs(5909) <= (inputs(57)) and not (inputs(47));
    layer0_outputs(5910) <= (inputs(160)) or (inputs(128));
    layer0_outputs(5911) <= not(inputs(219)) or (inputs(61));
    layer0_outputs(5912) <= not(inputs(66));
    layer0_outputs(5913) <= not(inputs(121));
    layer0_outputs(5914) <= (inputs(245)) xor (inputs(206));
    layer0_outputs(5915) <= not(inputs(181));
    layer0_outputs(5916) <= not((inputs(89)) or (inputs(78)));
    layer0_outputs(5917) <= not((inputs(75)) xor (inputs(88)));
    layer0_outputs(5918) <= (inputs(14)) or (inputs(43));
    layer0_outputs(5919) <= (inputs(208)) or (inputs(226));
    layer0_outputs(5920) <= inputs(217);
    layer0_outputs(5921) <= not(inputs(232));
    layer0_outputs(5922) <= (inputs(68)) and not (inputs(223));
    layer0_outputs(5923) <= (inputs(66)) xor (inputs(104));
    layer0_outputs(5924) <= not(inputs(147));
    layer0_outputs(5925) <= not((inputs(180)) or (inputs(239)));
    layer0_outputs(5926) <= not(inputs(213)) or (inputs(117));
    layer0_outputs(5927) <= (inputs(4)) xor (inputs(101));
    layer0_outputs(5928) <= inputs(127);
    layer0_outputs(5929) <= (inputs(9)) and not (inputs(17));
    layer0_outputs(5930) <= (inputs(96)) and (inputs(183));
    layer0_outputs(5931) <= (inputs(70)) xor (inputs(131));
    layer0_outputs(5932) <= (inputs(42)) or (inputs(19));
    layer0_outputs(5933) <= not(inputs(62)) or (inputs(155));
    layer0_outputs(5934) <= not(inputs(193));
    layer0_outputs(5935) <= (inputs(199)) and not (inputs(18));
    layer0_outputs(5936) <= (inputs(151)) and not (inputs(162));
    layer0_outputs(5937) <= inputs(86);
    layer0_outputs(5938) <= inputs(75);
    layer0_outputs(5939) <= (inputs(119)) or (inputs(29));
    layer0_outputs(5940) <= '1';
    layer0_outputs(5941) <= not((inputs(11)) xor (inputs(61)));
    layer0_outputs(5942) <= not((inputs(104)) xor (inputs(254)));
    layer0_outputs(5943) <= not(inputs(129));
    layer0_outputs(5944) <= (inputs(200)) and not (inputs(250));
    layer0_outputs(5945) <= (inputs(196)) or (inputs(221));
    layer0_outputs(5946) <= (inputs(12)) or (inputs(139));
    layer0_outputs(5947) <= inputs(221);
    layer0_outputs(5948) <= not(inputs(40));
    layer0_outputs(5949) <= not(inputs(60));
    layer0_outputs(5950) <= not((inputs(124)) xor (inputs(190)));
    layer0_outputs(5951) <= (inputs(71)) xor (inputs(11));
    layer0_outputs(5952) <= inputs(110);
    layer0_outputs(5953) <= (inputs(0)) or (inputs(250));
    layer0_outputs(5954) <= (inputs(11)) xor (inputs(143));
    layer0_outputs(5955) <= not(inputs(131)) or (inputs(12));
    layer0_outputs(5956) <= inputs(52);
    layer0_outputs(5957) <= not(inputs(138)) or (inputs(190));
    layer0_outputs(5958) <= inputs(213);
    layer0_outputs(5959) <= not((inputs(190)) or (inputs(176)));
    layer0_outputs(5960) <= (inputs(252)) or (inputs(243));
    layer0_outputs(5961) <= not((inputs(164)) or (inputs(134)));
    layer0_outputs(5962) <= not(inputs(113));
    layer0_outputs(5963) <= (inputs(182)) and not (inputs(255));
    layer0_outputs(5964) <= inputs(183);
    layer0_outputs(5965) <= not((inputs(187)) or (inputs(212)));
    layer0_outputs(5966) <= not(inputs(180));
    layer0_outputs(5967) <= (inputs(117)) or (inputs(245));
    layer0_outputs(5968) <= (inputs(138)) and not (inputs(189));
    layer0_outputs(5969) <= not(inputs(146)) or (inputs(254));
    layer0_outputs(5970) <= not((inputs(66)) or (inputs(131)));
    layer0_outputs(5971) <= not((inputs(219)) or (inputs(244)));
    layer0_outputs(5972) <= (inputs(247)) and not (inputs(21));
    layer0_outputs(5973) <= inputs(208);
    layer0_outputs(5974) <= not((inputs(71)) or (inputs(29)));
    layer0_outputs(5975) <= not((inputs(193)) or (inputs(223)));
    layer0_outputs(5976) <= inputs(143);
    layer0_outputs(5977) <= not((inputs(208)) or (inputs(4)));
    layer0_outputs(5978) <= not((inputs(160)) xor (inputs(251)));
    layer0_outputs(5979) <= (inputs(212)) and not (inputs(76));
    layer0_outputs(5980) <= (inputs(26)) xor (inputs(130));
    layer0_outputs(5981) <= not(inputs(175));
    layer0_outputs(5982) <= inputs(168);
    layer0_outputs(5983) <= not(inputs(229));
    layer0_outputs(5984) <= not(inputs(68));
    layer0_outputs(5985) <= (inputs(131)) and not (inputs(239));
    layer0_outputs(5986) <= not(inputs(26));
    layer0_outputs(5987) <= '1';
    layer0_outputs(5988) <= not((inputs(91)) or (inputs(5)));
    layer0_outputs(5989) <= not((inputs(9)) or (inputs(34)));
    layer0_outputs(5990) <= not(inputs(65));
    layer0_outputs(5991) <= inputs(171);
    layer0_outputs(5992) <= (inputs(157)) or (inputs(79));
    layer0_outputs(5993) <= inputs(140);
    layer0_outputs(5994) <= (inputs(52)) and not (inputs(62));
    layer0_outputs(5995) <= '0';
    layer0_outputs(5996) <= (inputs(169)) and not (inputs(225));
    layer0_outputs(5997) <= not((inputs(27)) xor (inputs(103)));
    layer0_outputs(5998) <= not((inputs(86)) xor (inputs(67)));
    layer0_outputs(5999) <= not((inputs(86)) xor (inputs(36)));
    layer0_outputs(6000) <= not((inputs(105)) or (inputs(205)));
    layer0_outputs(6001) <= not((inputs(57)) or (inputs(166)));
    layer0_outputs(6002) <= '1';
    layer0_outputs(6003) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(6004) <= (inputs(32)) xor (inputs(203));
    layer0_outputs(6005) <= not(inputs(148));
    layer0_outputs(6006) <= not(inputs(41));
    layer0_outputs(6007) <= not(inputs(229));
    layer0_outputs(6008) <= (inputs(35)) and not (inputs(172));
    layer0_outputs(6009) <= not(inputs(190));
    layer0_outputs(6010) <= not(inputs(81));
    layer0_outputs(6011) <= inputs(213);
    layer0_outputs(6012) <= inputs(6);
    layer0_outputs(6013) <= inputs(232);
    layer0_outputs(6014) <= not(inputs(1));
    layer0_outputs(6015) <= inputs(197);
    layer0_outputs(6016) <= not((inputs(11)) or (inputs(206)));
    layer0_outputs(6017) <= not(inputs(7));
    layer0_outputs(6018) <= '1';
    layer0_outputs(6019) <= '0';
    layer0_outputs(6020) <= inputs(144);
    layer0_outputs(6021) <= inputs(226);
    layer0_outputs(6022) <= not(inputs(164)) or (inputs(78));
    layer0_outputs(6023) <= (inputs(126)) or (inputs(213));
    layer0_outputs(6024) <= not(inputs(203)) or (inputs(107));
    layer0_outputs(6025) <= (inputs(195)) xor (inputs(72));
    layer0_outputs(6026) <= inputs(191);
    layer0_outputs(6027) <= (inputs(234)) or (inputs(41));
    layer0_outputs(6028) <= inputs(149);
    layer0_outputs(6029) <= '1';
    layer0_outputs(6030) <= not(inputs(7));
    layer0_outputs(6031) <= (inputs(163)) and not (inputs(47));
    layer0_outputs(6032) <= not((inputs(241)) xor (inputs(167)));
    layer0_outputs(6033) <= inputs(16);
    layer0_outputs(6034) <= (inputs(157)) xor (inputs(60));
    layer0_outputs(6035) <= inputs(204);
    layer0_outputs(6036) <= not(inputs(163));
    layer0_outputs(6037) <= not((inputs(117)) xor (inputs(103)));
    layer0_outputs(6038) <= not(inputs(21));
    layer0_outputs(6039) <= not((inputs(204)) or (inputs(157)));
    layer0_outputs(6040) <= not(inputs(193));
    layer0_outputs(6041) <= inputs(40);
    layer0_outputs(6042) <= not(inputs(228)) or (inputs(135));
    layer0_outputs(6043) <= not((inputs(107)) or (inputs(57)));
    layer0_outputs(6044) <= (inputs(184)) and (inputs(146));
    layer0_outputs(6045) <= not(inputs(10)) or (inputs(173));
    layer0_outputs(6046) <= not((inputs(200)) or (inputs(201)));
    layer0_outputs(6047) <= (inputs(1)) or (inputs(51));
    layer0_outputs(6048) <= (inputs(94)) or (inputs(253));
    layer0_outputs(6049) <= not(inputs(117)) or (inputs(146));
    layer0_outputs(6050) <= not(inputs(191));
    layer0_outputs(6051) <= not(inputs(193));
    layer0_outputs(6052) <= (inputs(16)) xor (inputs(38));
    layer0_outputs(6053) <= not(inputs(72));
    layer0_outputs(6054) <= (inputs(82)) and not (inputs(72));
    layer0_outputs(6055) <= (inputs(174)) xor (inputs(8));
    layer0_outputs(6056) <= inputs(171);
    layer0_outputs(6057) <= inputs(198);
    layer0_outputs(6058) <= not(inputs(49));
    layer0_outputs(6059) <= (inputs(61)) xor (inputs(233));
    layer0_outputs(6060) <= (inputs(212)) and not (inputs(13));
    layer0_outputs(6061) <= (inputs(234)) and not (inputs(144));
    layer0_outputs(6062) <= not(inputs(13));
    layer0_outputs(6063) <= inputs(65);
    layer0_outputs(6064) <= not((inputs(176)) xor (inputs(112)));
    layer0_outputs(6065) <= (inputs(136)) and not (inputs(215));
    layer0_outputs(6066) <= (inputs(194)) or (inputs(210));
    layer0_outputs(6067) <= inputs(244);
    layer0_outputs(6068) <= inputs(230);
    layer0_outputs(6069) <= not(inputs(154)) or (inputs(150));
    layer0_outputs(6070) <= (inputs(249)) or (inputs(210));
    layer0_outputs(6071) <= not(inputs(105));
    layer0_outputs(6072) <= not(inputs(51)) or (inputs(243));
    layer0_outputs(6073) <= not(inputs(55));
    layer0_outputs(6074) <= inputs(132);
    layer0_outputs(6075) <= not(inputs(242));
    layer0_outputs(6076) <= (inputs(85)) and not (inputs(204));
    layer0_outputs(6077) <= inputs(130);
    layer0_outputs(6078) <= (inputs(215)) or (inputs(195));
    layer0_outputs(6079) <= (inputs(162)) xor (inputs(76));
    layer0_outputs(6080) <= not((inputs(56)) xor (inputs(100)));
    layer0_outputs(6081) <= not((inputs(152)) xor (inputs(197)));
    layer0_outputs(6082) <= not(inputs(71)) or (inputs(239));
    layer0_outputs(6083) <= (inputs(108)) and (inputs(140));
    layer0_outputs(6084) <= not((inputs(219)) or (inputs(30)));
    layer0_outputs(6085) <= not(inputs(100)) or (inputs(127));
    layer0_outputs(6086) <= not(inputs(45));
    layer0_outputs(6087) <= not((inputs(152)) or (inputs(134)));
    layer0_outputs(6088) <= (inputs(255)) and not (inputs(236));
    layer0_outputs(6089) <= not(inputs(107));
    layer0_outputs(6090) <= '1';
    layer0_outputs(6091) <= inputs(130);
    layer0_outputs(6092) <= not(inputs(145)) or (inputs(103));
    layer0_outputs(6093) <= (inputs(193)) and not (inputs(253));
    layer0_outputs(6094) <= inputs(136);
    layer0_outputs(6095) <= not(inputs(36));
    layer0_outputs(6096) <= (inputs(204)) or (inputs(245));
    layer0_outputs(6097) <= not((inputs(143)) or (inputs(55)));
    layer0_outputs(6098) <= not(inputs(61)) or (inputs(194));
    layer0_outputs(6099) <= inputs(116);
    layer0_outputs(6100) <= not((inputs(30)) or (inputs(128)));
    layer0_outputs(6101) <= (inputs(67)) or (inputs(255));
    layer0_outputs(6102) <= (inputs(255)) and not (inputs(224));
    layer0_outputs(6103) <= (inputs(98)) and not (inputs(48));
    layer0_outputs(6104) <= (inputs(250)) and not (inputs(4));
    layer0_outputs(6105) <= not((inputs(80)) or (inputs(86)));
    layer0_outputs(6106) <= inputs(178);
    layer0_outputs(6107) <= (inputs(151)) and not (inputs(13));
    layer0_outputs(6108) <= not((inputs(10)) or (inputs(26)));
    layer0_outputs(6109) <= not((inputs(210)) or (inputs(174)));
    layer0_outputs(6110) <= inputs(148);
    layer0_outputs(6111) <= (inputs(176)) or (inputs(213));
    layer0_outputs(6112) <= inputs(21);
    layer0_outputs(6113) <= not(inputs(222)) or (inputs(31));
    layer0_outputs(6114) <= (inputs(94)) or (inputs(28));
    layer0_outputs(6115) <= inputs(117);
    layer0_outputs(6116) <= not((inputs(77)) xor (inputs(188)));
    layer0_outputs(6117) <= not((inputs(203)) or (inputs(127)));
    layer0_outputs(6118) <= not(inputs(147));
    layer0_outputs(6119) <= inputs(149);
    layer0_outputs(6120) <= not(inputs(24)) or (inputs(195));
    layer0_outputs(6121) <= (inputs(6)) or (inputs(104));
    layer0_outputs(6122) <= (inputs(224)) and not (inputs(163));
    layer0_outputs(6123) <= inputs(99);
    layer0_outputs(6124) <= not((inputs(53)) xor (inputs(48)));
    layer0_outputs(6125) <= (inputs(41)) or (inputs(46));
    layer0_outputs(6126) <= not((inputs(208)) xor (inputs(18)));
    layer0_outputs(6127) <= not(inputs(124));
    layer0_outputs(6128) <= (inputs(78)) or (inputs(110));
    layer0_outputs(6129) <= not(inputs(47));
    layer0_outputs(6130) <= not(inputs(72)) or (inputs(249));
    layer0_outputs(6131) <= not((inputs(199)) xor (inputs(167)));
    layer0_outputs(6132) <= not(inputs(209)) or (inputs(225));
    layer0_outputs(6133) <= inputs(39);
    layer0_outputs(6134) <= inputs(112);
    layer0_outputs(6135) <= not(inputs(23)) or (inputs(157));
    layer0_outputs(6136) <= (inputs(18)) or (inputs(164));
    layer0_outputs(6137) <= (inputs(220)) xor (inputs(55));
    layer0_outputs(6138) <= inputs(113);
    layer0_outputs(6139) <= (inputs(202)) and (inputs(142));
    layer0_outputs(6140) <= (inputs(90)) and (inputs(233));
    layer0_outputs(6141) <= not((inputs(208)) or (inputs(117)));
    layer0_outputs(6142) <= not(inputs(248)) or (inputs(75));
    layer0_outputs(6143) <= (inputs(42)) and not (inputs(182));
    layer0_outputs(6144) <= not((inputs(158)) or (inputs(111)));
    layer0_outputs(6145) <= (inputs(30)) xor (inputs(174));
    layer0_outputs(6146) <= inputs(169);
    layer0_outputs(6147) <= (inputs(200)) and not (inputs(170));
    layer0_outputs(6148) <= not(inputs(211));
    layer0_outputs(6149) <= not(inputs(191));
    layer0_outputs(6150) <= '0';
    layer0_outputs(6151) <= not((inputs(92)) or (inputs(252)));
    layer0_outputs(6152) <= not(inputs(152)) or (inputs(193));
    layer0_outputs(6153) <= inputs(176);
    layer0_outputs(6154) <= inputs(105);
    layer0_outputs(6155) <= not(inputs(26));
    layer0_outputs(6156) <= not(inputs(29)) or (inputs(205));
    layer0_outputs(6157) <= inputs(147);
    layer0_outputs(6158) <= not((inputs(225)) and (inputs(255)));
    layer0_outputs(6159) <= inputs(129);
    layer0_outputs(6160) <= inputs(177);
    layer0_outputs(6161) <= not((inputs(7)) xor (inputs(52)));
    layer0_outputs(6162) <= not((inputs(79)) and (inputs(90)));
    layer0_outputs(6163) <= inputs(121);
    layer0_outputs(6164) <= not((inputs(65)) or (inputs(234)));
    layer0_outputs(6165) <= not(inputs(78));
    layer0_outputs(6166) <= not((inputs(157)) xor (inputs(174)));
    layer0_outputs(6167) <= not(inputs(105));
    layer0_outputs(6168) <= (inputs(216)) and not (inputs(77));
    layer0_outputs(6169) <= (inputs(115)) or (inputs(115));
    layer0_outputs(6170) <= (inputs(44)) and not (inputs(253));
    layer0_outputs(6171) <= (inputs(138)) or (inputs(17));
    layer0_outputs(6172) <= inputs(124);
    layer0_outputs(6173) <= not((inputs(62)) or (inputs(239)));
    layer0_outputs(6174) <= inputs(54);
    layer0_outputs(6175) <= inputs(75);
    layer0_outputs(6176) <= not((inputs(226)) or (inputs(163)));
    layer0_outputs(6177) <= not((inputs(15)) or (inputs(42)));
    layer0_outputs(6178) <= (inputs(149)) and not (inputs(184));
    layer0_outputs(6179) <= not(inputs(143)) or (inputs(52));
    layer0_outputs(6180) <= not(inputs(174));
    layer0_outputs(6181) <= not((inputs(0)) or (inputs(234)));
    layer0_outputs(6182) <= inputs(230);
    layer0_outputs(6183) <= not(inputs(56)) or (inputs(126));
    layer0_outputs(6184) <= (inputs(28)) and not (inputs(187));
    layer0_outputs(6185) <= not((inputs(231)) or (inputs(63)));
    layer0_outputs(6186) <= (inputs(247)) xor (inputs(192));
    layer0_outputs(6187) <= (inputs(82)) or (inputs(135));
    layer0_outputs(6188) <= not((inputs(224)) or (inputs(245)));
    layer0_outputs(6189) <= (inputs(151)) or (inputs(160));
    layer0_outputs(6190) <= (inputs(93)) or (inputs(73));
    layer0_outputs(6191) <= not((inputs(238)) or (inputs(64)));
    layer0_outputs(6192) <= (inputs(247)) and not (inputs(122));
    layer0_outputs(6193) <= not(inputs(5)) or (inputs(175));
    layer0_outputs(6194) <= inputs(18);
    layer0_outputs(6195) <= (inputs(198)) xor (inputs(175));
    layer0_outputs(6196) <= not((inputs(67)) or (inputs(228)));
    layer0_outputs(6197) <= not(inputs(72));
    layer0_outputs(6198) <= (inputs(27)) and (inputs(148));
    layer0_outputs(6199) <= (inputs(172)) or (inputs(157));
    layer0_outputs(6200) <= not(inputs(184));
    layer0_outputs(6201) <= not((inputs(181)) or (inputs(13)));
    layer0_outputs(6202) <= not((inputs(14)) or (inputs(126)));
    layer0_outputs(6203) <= not(inputs(152));
    layer0_outputs(6204) <= (inputs(149)) and not (inputs(255));
    layer0_outputs(6205) <= (inputs(30)) and not (inputs(102));
    layer0_outputs(6206) <= not(inputs(3)) or (inputs(47));
    layer0_outputs(6207) <= (inputs(87)) xor (inputs(75));
    layer0_outputs(6208) <= not(inputs(159)) or (inputs(103));
    layer0_outputs(6209) <= not(inputs(40)) or (inputs(145));
    layer0_outputs(6210) <= not(inputs(245));
    layer0_outputs(6211) <= not(inputs(26));
    layer0_outputs(6212) <= not((inputs(76)) xor (inputs(156)));
    layer0_outputs(6213) <= not(inputs(198)) or (inputs(154));
    layer0_outputs(6214) <= (inputs(115)) xor (inputs(24));
    layer0_outputs(6215) <= (inputs(148)) or (inputs(131));
    layer0_outputs(6216) <= not((inputs(107)) xor (inputs(160)));
    layer0_outputs(6217) <= inputs(202);
    layer0_outputs(6218) <= not(inputs(28)) or (inputs(193));
    layer0_outputs(6219) <= (inputs(50)) xor (inputs(109));
    layer0_outputs(6220) <= not(inputs(103)) or (inputs(48));
    layer0_outputs(6221) <= (inputs(246)) and not (inputs(220));
    layer0_outputs(6222) <= '1';
    layer0_outputs(6223) <= (inputs(119)) and not (inputs(140));
    layer0_outputs(6224) <= not(inputs(137));
    layer0_outputs(6225) <= (inputs(2)) and (inputs(39));
    layer0_outputs(6226) <= inputs(201);
    layer0_outputs(6227) <= not(inputs(148));
    layer0_outputs(6228) <= (inputs(227)) or (inputs(33));
    layer0_outputs(6229) <= not((inputs(31)) or (inputs(191)));
    layer0_outputs(6230) <= not((inputs(142)) xor (inputs(171)));
    layer0_outputs(6231) <= not(inputs(125)) or (inputs(163));
    layer0_outputs(6232) <= (inputs(162)) and not (inputs(92));
    layer0_outputs(6233) <= not((inputs(17)) or (inputs(241)));
    layer0_outputs(6234) <= not(inputs(104));
    layer0_outputs(6235) <= not(inputs(243)) or (inputs(80));
    layer0_outputs(6236) <= (inputs(118)) xor (inputs(127));
    layer0_outputs(6237) <= not(inputs(29)) or (inputs(70));
    layer0_outputs(6238) <= not((inputs(229)) or (inputs(245)));
    layer0_outputs(6239) <= (inputs(21)) or (inputs(43));
    layer0_outputs(6240) <= not(inputs(216));
    layer0_outputs(6241) <= (inputs(2)) and not (inputs(191));
    layer0_outputs(6242) <= not((inputs(88)) xor (inputs(13)));
    layer0_outputs(6243) <= not((inputs(32)) or (inputs(152)));
    layer0_outputs(6244) <= not((inputs(45)) xor (inputs(60)));
    layer0_outputs(6245) <= (inputs(212)) xor (inputs(65));
    layer0_outputs(6246) <= inputs(200);
    layer0_outputs(6247) <= (inputs(209)) or (inputs(63));
    layer0_outputs(6248) <= (inputs(58)) xor (inputs(176));
    layer0_outputs(6249) <= not(inputs(247));
    layer0_outputs(6250) <= (inputs(154)) and not (inputs(72));
    layer0_outputs(6251) <= inputs(130);
    layer0_outputs(6252) <= not(inputs(82));
    layer0_outputs(6253) <= (inputs(84)) and not (inputs(195));
    layer0_outputs(6254) <= not((inputs(146)) xor (inputs(100)));
    layer0_outputs(6255) <= (inputs(183)) xor (inputs(105));
    layer0_outputs(6256) <= (inputs(177)) and (inputs(147));
    layer0_outputs(6257) <= inputs(91);
    layer0_outputs(6258) <= '0';
    layer0_outputs(6259) <= (inputs(64)) and not (inputs(31));
    layer0_outputs(6260) <= (inputs(202)) or (inputs(173));
    layer0_outputs(6261) <= not(inputs(57));
    layer0_outputs(6262) <= (inputs(155)) and not (inputs(12));
    layer0_outputs(6263) <= not(inputs(188)) or (inputs(170));
    layer0_outputs(6264) <= inputs(255);
    layer0_outputs(6265) <= not((inputs(68)) xor (inputs(102)));
    layer0_outputs(6266) <= (inputs(25)) and not (inputs(162));
    layer0_outputs(6267) <= not((inputs(236)) xor (inputs(228)));
    layer0_outputs(6268) <= not((inputs(145)) and (inputs(218)));
    layer0_outputs(6269) <= (inputs(151)) or (inputs(68));
    layer0_outputs(6270) <= inputs(120);
    layer0_outputs(6271) <= not(inputs(104));
    layer0_outputs(6272) <= inputs(38);
    layer0_outputs(6273) <= not(inputs(12)) or (inputs(132));
    layer0_outputs(6274) <= (inputs(218)) and not (inputs(168));
    layer0_outputs(6275) <= inputs(19);
    layer0_outputs(6276) <= (inputs(97)) and not (inputs(61));
    layer0_outputs(6277) <= inputs(158);
    layer0_outputs(6278) <= not((inputs(90)) or (inputs(148)));
    layer0_outputs(6279) <= not(inputs(6)) or (inputs(69));
    layer0_outputs(6280) <= inputs(118);
    layer0_outputs(6281) <= inputs(141);
    layer0_outputs(6282) <= not(inputs(91)) or (inputs(245));
    layer0_outputs(6283) <= (inputs(248)) and (inputs(61));
    layer0_outputs(6284) <= (inputs(117)) and not (inputs(110));
    layer0_outputs(6285) <= not(inputs(209));
    layer0_outputs(6286) <= inputs(66);
    layer0_outputs(6287) <= inputs(194);
    layer0_outputs(6288) <= not((inputs(53)) xor (inputs(55)));
    layer0_outputs(6289) <= not((inputs(77)) or (inputs(30)));
    layer0_outputs(6290) <= not((inputs(144)) or (inputs(247)));
    layer0_outputs(6291) <= not((inputs(228)) or (inputs(101)));
    layer0_outputs(6292) <= not((inputs(64)) or (inputs(119)));
    layer0_outputs(6293) <= (inputs(209)) xor (inputs(6));
    layer0_outputs(6294) <= not(inputs(41)) or (inputs(36));
    layer0_outputs(6295) <= not(inputs(3));
    layer0_outputs(6296) <= not(inputs(208)) or (inputs(0));
    layer0_outputs(6297) <= (inputs(139)) and not (inputs(69));
    layer0_outputs(6298) <= inputs(139);
    layer0_outputs(6299) <= not(inputs(4));
    layer0_outputs(6300) <= inputs(228);
    layer0_outputs(6301) <= inputs(9);
    layer0_outputs(6302) <= (inputs(52)) or (inputs(14));
    layer0_outputs(6303) <= not((inputs(234)) xor (inputs(68)));
    layer0_outputs(6304) <= inputs(9);
    layer0_outputs(6305) <= inputs(21);
    layer0_outputs(6306) <= not(inputs(247)) or (inputs(7));
    layer0_outputs(6307) <= inputs(98);
    layer0_outputs(6308) <= not(inputs(27));
    layer0_outputs(6309) <= not(inputs(167));
    layer0_outputs(6310) <= '1';
    layer0_outputs(6311) <= (inputs(227)) xor (inputs(175));
    layer0_outputs(6312) <= not(inputs(62));
    layer0_outputs(6313) <= (inputs(134)) and not (inputs(4));
    layer0_outputs(6314) <= inputs(36);
    layer0_outputs(6315) <= not((inputs(169)) and (inputs(195)));
    layer0_outputs(6316) <= (inputs(23)) or (inputs(174));
    layer0_outputs(6317) <= (inputs(145)) or (inputs(150));
    layer0_outputs(6318) <= not((inputs(85)) or (inputs(113)));
    layer0_outputs(6319) <= inputs(130);
    layer0_outputs(6320) <= not(inputs(153)) or (inputs(93));
    layer0_outputs(6321) <= (inputs(246)) and not (inputs(15));
    layer0_outputs(6322) <= (inputs(122)) and not (inputs(84));
    layer0_outputs(6323) <= not(inputs(219));
    layer0_outputs(6324) <= (inputs(188)) and not (inputs(71));
    layer0_outputs(6325) <= not(inputs(167));
    layer0_outputs(6326) <= (inputs(174)) and not (inputs(161));
    layer0_outputs(6327) <= not(inputs(186)) or (inputs(116));
    layer0_outputs(6328) <= not(inputs(166)) or (inputs(223));
    layer0_outputs(6329) <= '0';
    layer0_outputs(6330) <= not(inputs(152));
    layer0_outputs(6331) <= not(inputs(75));
    layer0_outputs(6332) <= not((inputs(33)) or (inputs(14)));
    layer0_outputs(6333) <= (inputs(148)) or (inputs(99));
    layer0_outputs(6334) <= not(inputs(50));
    layer0_outputs(6335) <= not(inputs(23)) or (inputs(204));
    layer0_outputs(6336) <= not(inputs(1));
    layer0_outputs(6337) <= (inputs(115)) and not (inputs(11));
    layer0_outputs(6338) <= not((inputs(234)) or (inputs(147)));
    layer0_outputs(6339) <= inputs(130);
    layer0_outputs(6340) <= inputs(138);
    layer0_outputs(6341) <= inputs(19);
    layer0_outputs(6342) <= inputs(102);
    layer0_outputs(6343) <= not((inputs(190)) or (inputs(228)));
    layer0_outputs(6344) <= not(inputs(4));
    layer0_outputs(6345) <= (inputs(59)) xor (inputs(43));
    layer0_outputs(6346) <= inputs(219);
    layer0_outputs(6347) <= inputs(39);
    layer0_outputs(6348) <= inputs(210);
    layer0_outputs(6349) <= (inputs(180)) and (inputs(247));
    layer0_outputs(6350) <= not((inputs(113)) or (inputs(106)));
    layer0_outputs(6351) <= not((inputs(176)) or (inputs(70)));
    layer0_outputs(6352) <= inputs(93);
    layer0_outputs(6353) <= (inputs(14)) or (inputs(170));
    layer0_outputs(6354) <= (inputs(226)) or (inputs(157));
    layer0_outputs(6355) <= (inputs(40)) and not (inputs(92));
    layer0_outputs(6356) <= not(inputs(23)) or (inputs(146));
    layer0_outputs(6357) <= (inputs(73)) xor (inputs(241));
    layer0_outputs(6358) <= not((inputs(43)) xor (inputs(143)));
    layer0_outputs(6359) <= not(inputs(198)) or (inputs(208));
    layer0_outputs(6360) <= inputs(197);
    layer0_outputs(6361) <= not(inputs(210));
    layer0_outputs(6362) <= (inputs(163)) and not (inputs(17));
    layer0_outputs(6363) <= not(inputs(122)) or (inputs(32));
    layer0_outputs(6364) <= inputs(173);
    layer0_outputs(6365) <= (inputs(230)) and not (inputs(45));
    layer0_outputs(6366) <= (inputs(117)) xor (inputs(160));
    layer0_outputs(6367) <= '0';
    layer0_outputs(6368) <= (inputs(42)) and (inputs(25));
    layer0_outputs(6369) <= '0';
    layer0_outputs(6370) <= (inputs(225)) and not (inputs(169));
    layer0_outputs(6371) <= (inputs(239)) or (inputs(105));
    layer0_outputs(6372) <= not(inputs(165)) or (inputs(175));
    layer0_outputs(6373) <= not(inputs(68));
    layer0_outputs(6374) <= (inputs(227)) and not (inputs(97));
    layer0_outputs(6375) <= not(inputs(149));
    layer0_outputs(6376) <= '0';
    layer0_outputs(6377) <= not((inputs(252)) or (inputs(155)));
    layer0_outputs(6378) <= (inputs(127)) and not (inputs(207));
    layer0_outputs(6379) <= not((inputs(178)) or (inputs(191)));
    layer0_outputs(6380) <= (inputs(152)) or (inputs(245));
    layer0_outputs(6381) <= (inputs(203)) or (inputs(4));
    layer0_outputs(6382) <= '1';
    layer0_outputs(6383) <= not(inputs(101));
    layer0_outputs(6384) <= (inputs(204)) and not (inputs(98));
    layer0_outputs(6385) <= not((inputs(12)) or (inputs(132)));
    layer0_outputs(6386) <= '1';
    layer0_outputs(6387) <= not(inputs(145)) or (inputs(104));
    layer0_outputs(6388) <= inputs(151);
    layer0_outputs(6389) <= (inputs(92)) xor (inputs(139));
    layer0_outputs(6390) <= inputs(9);
    layer0_outputs(6391) <= not(inputs(244)) or (inputs(234));
    layer0_outputs(6392) <= (inputs(224)) and not (inputs(250));
    layer0_outputs(6393) <= (inputs(120)) xor (inputs(50));
    layer0_outputs(6394) <= not(inputs(166));
    layer0_outputs(6395) <= not((inputs(146)) xor (inputs(88)));
    layer0_outputs(6396) <= not(inputs(232)) or (inputs(37));
    layer0_outputs(6397) <= not(inputs(55)) or (inputs(122));
    layer0_outputs(6398) <= inputs(92);
    layer0_outputs(6399) <= (inputs(113)) or (inputs(209));
    layer0_outputs(6400) <= not(inputs(104)) or (inputs(35));
    layer0_outputs(6401) <= (inputs(30)) or (inputs(145));
    layer0_outputs(6402) <= not(inputs(96));
    layer0_outputs(6403) <= not(inputs(51)) or (inputs(130));
    layer0_outputs(6404) <= inputs(91);
    layer0_outputs(6405) <= (inputs(118)) and not (inputs(239));
    layer0_outputs(6406) <= not((inputs(191)) and (inputs(14)));
    layer0_outputs(6407) <= (inputs(22)) and not (inputs(161));
    layer0_outputs(6408) <= not(inputs(19));
    layer0_outputs(6409) <= not(inputs(55)) or (inputs(109));
    layer0_outputs(6410) <= inputs(196);
    layer0_outputs(6411) <= not(inputs(157));
    layer0_outputs(6412) <= (inputs(188)) and not (inputs(17));
    layer0_outputs(6413) <= not(inputs(176));
    layer0_outputs(6414) <= not(inputs(88));
    layer0_outputs(6415) <= not(inputs(180));
    layer0_outputs(6416) <= (inputs(133)) and not (inputs(137));
    layer0_outputs(6417) <= not(inputs(107));
    layer0_outputs(6418) <= not(inputs(133));
    layer0_outputs(6419) <= not(inputs(168)) or (inputs(207));
    layer0_outputs(6420) <= not(inputs(5)) or (inputs(94));
    layer0_outputs(6421) <= inputs(242);
    layer0_outputs(6422) <= inputs(193);
    layer0_outputs(6423) <= (inputs(184)) and (inputs(249));
    layer0_outputs(6424) <= (inputs(115)) and not (inputs(220));
    layer0_outputs(6425) <= (inputs(231)) and not (inputs(79));
    layer0_outputs(6426) <= not(inputs(29));
    layer0_outputs(6427) <= (inputs(213)) and (inputs(112));
    layer0_outputs(6428) <= not(inputs(59));
    layer0_outputs(6429) <= not(inputs(215));
    layer0_outputs(6430) <= (inputs(151)) and not (inputs(143));
    layer0_outputs(6431) <= inputs(176);
    layer0_outputs(6432) <= not(inputs(38));
    layer0_outputs(6433) <= not((inputs(165)) or (inputs(49)));
    layer0_outputs(6434) <= (inputs(236)) or (inputs(32));
    layer0_outputs(6435) <= not(inputs(30)) or (inputs(129));
    layer0_outputs(6436) <= (inputs(77)) or (inputs(118));
    layer0_outputs(6437) <= not(inputs(188));
    layer0_outputs(6438) <= inputs(117);
    layer0_outputs(6439) <= (inputs(120)) or (inputs(90));
    layer0_outputs(6440) <= not(inputs(53)) or (inputs(224));
    layer0_outputs(6441) <= (inputs(124)) and not (inputs(54));
    layer0_outputs(6442) <= (inputs(102)) and not (inputs(12));
    layer0_outputs(6443) <= not(inputs(168)) or (inputs(47));
    layer0_outputs(6444) <= (inputs(196)) or (inputs(173));
    layer0_outputs(6445) <= (inputs(0)) or (inputs(103));
    layer0_outputs(6446) <= not((inputs(60)) or (inputs(141)));
    layer0_outputs(6447) <= not(inputs(234));
    layer0_outputs(6448) <= not((inputs(6)) xor (inputs(53)));
    layer0_outputs(6449) <= not((inputs(12)) or (inputs(114)));
    layer0_outputs(6450) <= (inputs(144)) and not (inputs(118));
    layer0_outputs(6451) <= (inputs(168)) and not (inputs(69));
    layer0_outputs(6452) <= not((inputs(160)) xor (inputs(102)));
    layer0_outputs(6453) <= (inputs(27)) and not (inputs(249));
    layer0_outputs(6454) <= (inputs(58)) and not (inputs(225));
    layer0_outputs(6455) <= (inputs(176)) or (inputs(187));
    layer0_outputs(6456) <= (inputs(84)) and not (inputs(160));
    layer0_outputs(6457) <= '0';
    layer0_outputs(6458) <= (inputs(166)) or (inputs(96));
    layer0_outputs(6459) <= not((inputs(106)) xor (inputs(16)));
    layer0_outputs(6460) <= not((inputs(230)) or (inputs(87)));
    layer0_outputs(6461) <= not(inputs(28)) or (inputs(255));
    layer0_outputs(6462) <= inputs(82);
    layer0_outputs(6463) <= not(inputs(14));
    layer0_outputs(6464) <= (inputs(85)) and not (inputs(32));
    layer0_outputs(6465) <= (inputs(78)) or (inputs(211));
    layer0_outputs(6466) <= inputs(25);
    layer0_outputs(6467) <= inputs(165);
    layer0_outputs(6468) <= not((inputs(196)) or (inputs(204)));
    layer0_outputs(6469) <= inputs(106);
    layer0_outputs(6470) <= not((inputs(180)) xor (inputs(225)));
    layer0_outputs(6471) <= (inputs(207)) and not (inputs(134));
    layer0_outputs(6472) <= not((inputs(140)) or (inputs(145)));
    layer0_outputs(6473) <= inputs(19);
    layer0_outputs(6474) <= not((inputs(173)) or (inputs(20)));
    layer0_outputs(6475) <= not((inputs(198)) or (inputs(236)));
    layer0_outputs(6476) <= (inputs(23)) or (inputs(207));
    layer0_outputs(6477) <= not(inputs(145)) or (inputs(239));
    layer0_outputs(6478) <= not(inputs(230));
    layer0_outputs(6479) <= (inputs(69)) and not (inputs(242));
    layer0_outputs(6480) <= (inputs(142)) and not (inputs(175));
    layer0_outputs(6481) <= (inputs(167)) xor (inputs(119));
    layer0_outputs(6482) <= '1';
    layer0_outputs(6483) <= (inputs(16)) xor (inputs(77));
    layer0_outputs(6484) <= (inputs(32)) xor (inputs(102));
    layer0_outputs(6485) <= '0';
    layer0_outputs(6486) <= inputs(18);
    layer0_outputs(6487) <= (inputs(51)) and not (inputs(8));
    layer0_outputs(6488) <= inputs(35);
    layer0_outputs(6489) <= not(inputs(161));
    layer0_outputs(6490) <= not((inputs(163)) xor (inputs(100)));
    layer0_outputs(6491) <= (inputs(32)) or (inputs(156));
    layer0_outputs(6492) <= (inputs(39)) and not (inputs(240));
    layer0_outputs(6493) <= (inputs(163)) and not (inputs(80));
    layer0_outputs(6494) <= (inputs(169)) and not (inputs(108));
    layer0_outputs(6495) <= inputs(66);
    layer0_outputs(6496) <= (inputs(199)) xor (inputs(180));
    layer0_outputs(6497) <= not(inputs(8));
    layer0_outputs(6498) <= not((inputs(133)) and (inputs(197)));
    layer0_outputs(6499) <= (inputs(55)) xor (inputs(67));
    layer0_outputs(6500) <= not(inputs(60));
    layer0_outputs(6501) <= not(inputs(105));
    layer0_outputs(6502) <= not(inputs(98));
    layer0_outputs(6503) <= (inputs(65)) xor (inputs(49));
    layer0_outputs(6504) <= (inputs(79)) and not (inputs(173));
    layer0_outputs(6505) <= (inputs(112)) and not (inputs(237));
    layer0_outputs(6506) <= not(inputs(138));
    layer0_outputs(6507) <= not(inputs(138));
    layer0_outputs(6508) <= (inputs(65)) or (inputs(202));
    layer0_outputs(6509) <= (inputs(80)) or (inputs(112));
    layer0_outputs(6510) <= not(inputs(69)) or (inputs(208));
    layer0_outputs(6511) <= not((inputs(29)) and (inputs(75)));
    layer0_outputs(6512) <= not(inputs(118)) or (inputs(63));
    layer0_outputs(6513) <= (inputs(33)) xor (inputs(226));
    layer0_outputs(6514) <= not(inputs(74)) or (inputs(215));
    layer0_outputs(6515) <= not((inputs(161)) and (inputs(91)));
    layer0_outputs(6516) <= (inputs(81)) or (inputs(221));
    layer0_outputs(6517) <= not((inputs(249)) xor (inputs(160)));
    layer0_outputs(6518) <= (inputs(56)) and not (inputs(77));
    layer0_outputs(6519) <= (inputs(67)) or (inputs(222));
    layer0_outputs(6520) <= not(inputs(72));
    layer0_outputs(6521) <= not(inputs(44)) or (inputs(175));
    layer0_outputs(6522) <= (inputs(72)) xor (inputs(202));
    layer0_outputs(6523) <= inputs(232);
    layer0_outputs(6524) <= inputs(162);
    layer0_outputs(6525) <= not(inputs(196));
    layer0_outputs(6526) <= not(inputs(129));
    layer0_outputs(6527) <= not((inputs(208)) xor (inputs(239)));
    layer0_outputs(6528) <= not((inputs(130)) xor (inputs(181)));
    layer0_outputs(6529) <= inputs(229);
    layer0_outputs(6530) <= not((inputs(19)) xor (inputs(10)));
    layer0_outputs(6531) <= inputs(18);
    layer0_outputs(6532) <= (inputs(57)) xor (inputs(50));
    layer0_outputs(6533) <= inputs(112);
    layer0_outputs(6534) <= (inputs(121)) xor (inputs(115));
    layer0_outputs(6535) <= not((inputs(82)) and (inputs(134)));
    layer0_outputs(6536) <= inputs(138);
    layer0_outputs(6537) <= (inputs(140)) and not (inputs(51));
    layer0_outputs(6538) <= not((inputs(44)) or (inputs(218)));
    layer0_outputs(6539) <= inputs(115);
    layer0_outputs(6540) <= not(inputs(103));
    layer0_outputs(6541) <= not((inputs(120)) or (inputs(137)));
    layer0_outputs(6542) <= not((inputs(80)) xor (inputs(83)));
    layer0_outputs(6543) <= not((inputs(249)) xor (inputs(183)));
    layer0_outputs(6544) <= not((inputs(58)) xor (inputs(61)));
    layer0_outputs(6545) <= (inputs(85)) and not (inputs(72));
    layer0_outputs(6546) <= not(inputs(79)) or (inputs(152));
    layer0_outputs(6547) <= (inputs(40)) and (inputs(67));
    layer0_outputs(6548) <= inputs(183);
    layer0_outputs(6549) <= not((inputs(138)) or (inputs(15)));
    layer0_outputs(6550) <= not((inputs(235)) xor (inputs(251)));
    layer0_outputs(6551) <= inputs(182);
    layer0_outputs(6552) <= (inputs(96)) or (inputs(225));
    layer0_outputs(6553) <= not((inputs(172)) xor (inputs(62)));
    layer0_outputs(6554) <= not((inputs(149)) xor (inputs(17)));
    layer0_outputs(6555) <= (inputs(194)) or (inputs(84));
    layer0_outputs(6556) <= (inputs(110)) xor (inputs(238));
    layer0_outputs(6557) <= inputs(195);
    layer0_outputs(6558) <= (inputs(216)) and not (inputs(109));
    layer0_outputs(6559) <= not((inputs(169)) or (inputs(49)));
    layer0_outputs(6560) <= not(inputs(94));
    layer0_outputs(6561) <= '1';
    layer0_outputs(6562) <= inputs(161);
    layer0_outputs(6563) <= '0';
    layer0_outputs(6564) <= inputs(224);
    layer0_outputs(6565) <= not((inputs(175)) xor (inputs(122)));
    layer0_outputs(6566) <= not((inputs(215)) or (inputs(223)));
    layer0_outputs(6567) <= not((inputs(177)) xor (inputs(88)));
    layer0_outputs(6568) <= inputs(217);
    layer0_outputs(6569) <= '1';
    layer0_outputs(6570) <= (inputs(47)) and not (inputs(254));
    layer0_outputs(6571) <= not(inputs(97));
    layer0_outputs(6572) <= not((inputs(74)) or (inputs(49)));
    layer0_outputs(6573) <= not(inputs(74));
    layer0_outputs(6574) <= (inputs(106)) and not (inputs(249));
    layer0_outputs(6575) <= not((inputs(47)) or (inputs(95)));
    layer0_outputs(6576) <= not(inputs(120)) or (inputs(204));
    layer0_outputs(6577) <= inputs(81);
    layer0_outputs(6578) <= (inputs(89)) and not (inputs(4));
    layer0_outputs(6579) <= inputs(148);
    layer0_outputs(6580) <= inputs(119);
    layer0_outputs(6581) <= (inputs(85)) and not (inputs(125));
    layer0_outputs(6582) <= not((inputs(72)) or (inputs(2)));
    layer0_outputs(6583) <= not(inputs(80));
    layer0_outputs(6584) <= not((inputs(198)) xor (inputs(134)));
    layer0_outputs(6585) <= not(inputs(166));
    layer0_outputs(6586) <= not((inputs(30)) or (inputs(223)));
    layer0_outputs(6587) <= '1';
    layer0_outputs(6588) <= (inputs(160)) and not (inputs(8));
    layer0_outputs(6589) <= not((inputs(100)) or (inputs(83)));
    layer0_outputs(6590) <= not(inputs(213)) or (inputs(109));
    layer0_outputs(6591) <= not(inputs(99));
    layer0_outputs(6592) <= (inputs(206)) and not (inputs(246));
    layer0_outputs(6593) <= not(inputs(188)) or (inputs(67));
    layer0_outputs(6594) <= (inputs(254)) or (inputs(165));
    layer0_outputs(6595) <= '0';
    layer0_outputs(6596) <= (inputs(65)) or (inputs(64));
    layer0_outputs(6597) <= (inputs(129)) or (inputs(114));
    layer0_outputs(6598) <= not(inputs(140)) or (inputs(195));
    layer0_outputs(6599) <= not(inputs(91));
    layer0_outputs(6600) <= inputs(245);
    layer0_outputs(6601) <= (inputs(63)) or (inputs(136));
    layer0_outputs(6602) <= inputs(164);
    layer0_outputs(6603) <= not((inputs(138)) or (inputs(23)));
    layer0_outputs(6604) <= not(inputs(134));
    layer0_outputs(6605) <= inputs(104);
    layer0_outputs(6606) <= not((inputs(31)) or (inputs(18)));
    layer0_outputs(6607) <= inputs(74);
    layer0_outputs(6608) <= not(inputs(225));
    layer0_outputs(6609) <= (inputs(164)) xor (inputs(118));
    layer0_outputs(6610) <= (inputs(65)) or (inputs(150));
    layer0_outputs(6611) <= inputs(177);
    layer0_outputs(6612) <= (inputs(231)) and not (inputs(241));
    layer0_outputs(6613) <= not(inputs(187)) or (inputs(238));
    layer0_outputs(6614) <= (inputs(9)) and (inputs(37));
    layer0_outputs(6615) <= (inputs(170)) or (inputs(199));
    layer0_outputs(6616) <= (inputs(53)) and (inputs(141));
    layer0_outputs(6617) <= (inputs(26)) and (inputs(107));
    layer0_outputs(6618) <= not(inputs(51));
    layer0_outputs(6619) <= not((inputs(106)) or (inputs(129)));
    layer0_outputs(6620) <= inputs(221);
    layer0_outputs(6621) <= inputs(0);
    layer0_outputs(6622) <= (inputs(165)) and not (inputs(99));
    layer0_outputs(6623) <= '1';
    layer0_outputs(6624) <= (inputs(193)) xor (inputs(255));
    layer0_outputs(6625) <= not((inputs(157)) or (inputs(216)));
    layer0_outputs(6626) <= (inputs(243)) xor (inputs(208));
    layer0_outputs(6627) <= not((inputs(72)) or (inputs(139)));
    layer0_outputs(6628) <= (inputs(228)) and (inputs(74));
    layer0_outputs(6629) <= not((inputs(133)) or (inputs(46)));
    layer0_outputs(6630) <= (inputs(174)) or (inputs(43));
    layer0_outputs(6631) <= not(inputs(209));
    layer0_outputs(6632) <= inputs(76);
    layer0_outputs(6633) <= not((inputs(244)) xor (inputs(109)));
    layer0_outputs(6634) <= (inputs(49)) xor (inputs(197));
    layer0_outputs(6635) <= not(inputs(55));
    layer0_outputs(6636) <= (inputs(179)) or (inputs(220));
    layer0_outputs(6637) <= not(inputs(97)) or (inputs(31));
    layer0_outputs(6638) <= not(inputs(192));
    layer0_outputs(6639) <= inputs(113);
    layer0_outputs(6640) <= (inputs(230)) and not (inputs(237));
    layer0_outputs(6641) <= (inputs(185)) and not (inputs(133));
    layer0_outputs(6642) <= (inputs(232)) xor (inputs(169));
    layer0_outputs(6643) <= inputs(206);
    layer0_outputs(6644) <= (inputs(98)) or (inputs(155));
    layer0_outputs(6645) <= inputs(12);
    layer0_outputs(6646) <= not(inputs(233));
    layer0_outputs(6647) <= not(inputs(199));
    layer0_outputs(6648) <= inputs(222);
    layer0_outputs(6649) <= (inputs(215)) and not (inputs(104));
    layer0_outputs(6650) <= not(inputs(127));
    layer0_outputs(6651) <= (inputs(233)) and not (inputs(79));
    layer0_outputs(6652) <= (inputs(61)) xor (inputs(58));
    layer0_outputs(6653) <= (inputs(201)) and not (inputs(33));
    layer0_outputs(6654) <= not((inputs(231)) or (inputs(141)));
    layer0_outputs(6655) <= not((inputs(191)) xor (inputs(115)));
    layer0_outputs(6656) <= (inputs(74)) and not (inputs(245));
    layer0_outputs(6657) <= not(inputs(38)) or (inputs(112));
    layer0_outputs(6658) <= inputs(170);
    layer0_outputs(6659) <= not(inputs(253)) or (inputs(156));
    layer0_outputs(6660) <= (inputs(13)) xor (inputs(130));
    layer0_outputs(6661) <= not(inputs(246)) or (inputs(66));
    layer0_outputs(6662) <= not(inputs(247)) or (inputs(242));
    layer0_outputs(6663) <= not(inputs(100)) or (inputs(63));
    layer0_outputs(6664) <= not((inputs(199)) and (inputs(136)));
    layer0_outputs(6665) <= inputs(214);
    layer0_outputs(6666) <= not(inputs(179)) or (inputs(138));
    layer0_outputs(6667) <= not(inputs(83));
    layer0_outputs(6668) <= not((inputs(107)) and (inputs(30)));
    layer0_outputs(6669) <= not((inputs(46)) xor (inputs(167)));
    layer0_outputs(6670) <= not((inputs(135)) xor (inputs(242)));
    layer0_outputs(6671) <= not(inputs(120)) or (inputs(64));
    layer0_outputs(6672) <= (inputs(32)) or (inputs(52));
    layer0_outputs(6673) <= not(inputs(167));
    layer0_outputs(6674) <= inputs(11);
    layer0_outputs(6675) <= inputs(105);
    layer0_outputs(6676) <= not(inputs(74));
    layer0_outputs(6677) <= not((inputs(226)) or (inputs(115)));
    layer0_outputs(6678) <= (inputs(74)) or (inputs(101));
    layer0_outputs(6679) <= (inputs(195)) and not (inputs(11));
    layer0_outputs(6680) <= not((inputs(7)) or (inputs(244)));
    layer0_outputs(6681) <= (inputs(3)) or (inputs(14));
    layer0_outputs(6682) <= not(inputs(4));
    layer0_outputs(6683) <= not(inputs(102));
    layer0_outputs(6684) <= inputs(151);
    layer0_outputs(6685) <= (inputs(35)) and not (inputs(135));
    layer0_outputs(6686) <= (inputs(181)) and not (inputs(79));
    layer0_outputs(6687) <= not((inputs(117)) xor (inputs(235)));
    layer0_outputs(6688) <= not(inputs(238));
    layer0_outputs(6689) <= not(inputs(80)) or (inputs(248));
    layer0_outputs(6690) <= not(inputs(247));
    layer0_outputs(6691) <= (inputs(19)) xor (inputs(78));
    layer0_outputs(6692) <= (inputs(207)) xor (inputs(163));
    layer0_outputs(6693) <= (inputs(181)) and not (inputs(183));
    layer0_outputs(6694) <= (inputs(111)) and not (inputs(232));
    layer0_outputs(6695) <= inputs(147);
    layer0_outputs(6696) <= not(inputs(9)) or (inputs(224));
    layer0_outputs(6697) <= not(inputs(230));
    layer0_outputs(6698) <= not(inputs(162));
    layer0_outputs(6699) <= (inputs(10)) or (inputs(53));
    layer0_outputs(6700) <= not(inputs(115));
    layer0_outputs(6701) <= (inputs(221)) or (inputs(220));
    layer0_outputs(6702) <= not((inputs(34)) or (inputs(40)));
    layer0_outputs(6703) <= not((inputs(238)) xor (inputs(7)));
    layer0_outputs(6704) <= not((inputs(79)) xor (inputs(9)));
    layer0_outputs(6705) <= not(inputs(229));
    layer0_outputs(6706) <= inputs(19);
    layer0_outputs(6707) <= (inputs(82)) or (inputs(123));
    layer0_outputs(6708) <= (inputs(115)) or (inputs(115));
    layer0_outputs(6709) <= (inputs(202)) xor (inputs(13));
    layer0_outputs(6710) <= (inputs(13)) and not (inputs(112));
    layer0_outputs(6711) <= not((inputs(90)) and (inputs(93)));
    layer0_outputs(6712) <= not(inputs(63)) or (inputs(1));
    layer0_outputs(6713) <= inputs(115);
    layer0_outputs(6714) <= inputs(37);
    layer0_outputs(6715) <= not((inputs(176)) or (inputs(161)));
    layer0_outputs(6716) <= not((inputs(126)) or (inputs(178)));
    layer0_outputs(6717) <= (inputs(237)) or (inputs(49));
    layer0_outputs(6718) <= not(inputs(70)) or (inputs(78));
    layer0_outputs(6719) <= (inputs(141)) and not (inputs(149));
    layer0_outputs(6720) <= not(inputs(20));
    layer0_outputs(6721) <= not(inputs(76));
    layer0_outputs(6722) <= inputs(91);
    layer0_outputs(6723) <= not(inputs(35)) or (inputs(62));
    layer0_outputs(6724) <= (inputs(45)) and not (inputs(210));
    layer0_outputs(6725) <= (inputs(247)) or (inputs(161));
    layer0_outputs(6726) <= not(inputs(100)) or (inputs(231));
    layer0_outputs(6727) <= not(inputs(209));
    layer0_outputs(6728) <= not(inputs(147));
    layer0_outputs(6729) <= inputs(184);
    layer0_outputs(6730) <= (inputs(8)) or (inputs(25));
    layer0_outputs(6731) <= (inputs(3)) xor (inputs(70));
    layer0_outputs(6732) <= (inputs(215)) and not (inputs(240));
    layer0_outputs(6733) <= not(inputs(175));
    layer0_outputs(6734) <= inputs(60);
    layer0_outputs(6735) <= not((inputs(71)) xor (inputs(225)));
    layer0_outputs(6736) <= inputs(98);
    layer0_outputs(6737) <= (inputs(10)) or (inputs(58));
    layer0_outputs(6738) <= not(inputs(72)) or (inputs(177));
    layer0_outputs(6739) <= (inputs(29)) xor (inputs(209));
    layer0_outputs(6740) <= not((inputs(126)) xor (inputs(18)));
    layer0_outputs(6741) <= not(inputs(180)) or (inputs(46));
    layer0_outputs(6742) <= (inputs(75)) and not (inputs(236));
    layer0_outputs(6743) <= not((inputs(138)) or (inputs(14)));
    layer0_outputs(6744) <= not(inputs(226)) or (inputs(144));
    layer0_outputs(6745) <= not(inputs(160));
    layer0_outputs(6746) <= inputs(105);
    layer0_outputs(6747) <= not(inputs(64));
    layer0_outputs(6748) <= not((inputs(80)) or (inputs(105)));
    layer0_outputs(6749) <= inputs(204);
    layer0_outputs(6750) <= not(inputs(120)) or (inputs(176));
    layer0_outputs(6751) <= inputs(111);
    layer0_outputs(6752) <= not(inputs(101));
    layer0_outputs(6753) <= not(inputs(86));
    layer0_outputs(6754) <= (inputs(166)) and not (inputs(147));
    layer0_outputs(6755) <= '1';
    layer0_outputs(6756) <= not(inputs(25)) or (inputs(244));
    layer0_outputs(6757) <= (inputs(174)) and not (inputs(125));
    layer0_outputs(6758) <= not(inputs(229)) or (inputs(46));
    layer0_outputs(6759) <= (inputs(143)) and (inputs(19));
    layer0_outputs(6760) <= not(inputs(167)) or (inputs(38));
    layer0_outputs(6761) <= inputs(154);
    layer0_outputs(6762) <= (inputs(182)) xor (inputs(250));
    layer0_outputs(6763) <= not(inputs(104));
    layer0_outputs(6764) <= (inputs(149)) or (inputs(148));
    layer0_outputs(6765) <= inputs(55);
    layer0_outputs(6766) <= not(inputs(202)) or (inputs(111));
    layer0_outputs(6767) <= not((inputs(23)) xor (inputs(50)));
    layer0_outputs(6768) <= not((inputs(218)) xor (inputs(107)));
    layer0_outputs(6769) <= not((inputs(33)) xor (inputs(62)));
    layer0_outputs(6770) <= not((inputs(39)) or (inputs(110)));
    layer0_outputs(6771) <= not(inputs(135));
    layer0_outputs(6772) <= (inputs(220)) or (inputs(113));
    layer0_outputs(6773) <= not((inputs(109)) xor (inputs(91)));
    layer0_outputs(6774) <= (inputs(144)) or (inputs(217));
    layer0_outputs(6775) <= inputs(233);
    layer0_outputs(6776) <= not(inputs(9)) or (inputs(188));
    layer0_outputs(6777) <= not((inputs(131)) or (inputs(97)));
    layer0_outputs(6778) <= inputs(67);
    layer0_outputs(6779) <= not((inputs(250)) or (inputs(172)));
    layer0_outputs(6780) <= '0';
    layer0_outputs(6781) <= not(inputs(25));
    layer0_outputs(6782) <= not((inputs(174)) or (inputs(212)));
    layer0_outputs(6783) <= not((inputs(255)) or (inputs(106)));
    layer0_outputs(6784) <= (inputs(145)) xor (inputs(142));
    layer0_outputs(6785) <= not(inputs(214)) or (inputs(35));
    layer0_outputs(6786) <= (inputs(234)) or (inputs(175));
    layer0_outputs(6787) <= not((inputs(35)) or (inputs(180)));
    layer0_outputs(6788) <= inputs(94);
    layer0_outputs(6789) <= not(inputs(164));
    layer0_outputs(6790) <= (inputs(95)) or (inputs(130));
    layer0_outputs(6791) <= (inputs(25)) and not (inputs(14));
    layer0_outputs(6792) <= inputs(217);
    layer0_outputs(6793) <= not(inputs(212));
    layer0_outputs(6794) <= not(inputs(183));
    layer0_outputs(6795) <= inputs(12);
    layer0_outputs(6796) <= (inputs(90)) and (inputs(54));
    layer0_outputs(6797) <= inputs(115);
    layer0_outputs(6798) <= (inputs(227)) or (inputs(3));
    layer0_outputs(6799) <= not(inputs(213)) or (inputs(81));
    layer0_outputs(6800) <= not(inputs(213)) or (inputs(15));
    layer0_outputs(6801) <= not(inputs(121));
    layer0_outputs(6802) <= (inputs(97)) or (inputs(35));
    layer0_outputs(6803) <= not(inputs(22));
    layer0_outputs(6804) <= (inputs(121)) and (inputs(186));
    layer0_outputs(6805) <= not(inputs(70));
    layer0_outputs(6806) <= (inputs(89)) or (inputs(32));
    layer0_outputs(6807) <= (inputs(117)) and not (inputs(2));
    layer0_outputs(6808) <= not((inputs(41)) or (inputs(175)));
    layer0_outputs(6809) <= not((inputs(108)) or (inputs(254)));
    layer0_outputs(6810) <= (inputs(236)) xor (inputs(253));
    layer0_outputs(6811) <= not(inputs(110)) or (inputs(176));
    layer0_outputs(6812) <= not(inputs(198)) or (inputs(149));
    layer0_outputs(6813) <= not((inputs(47)) and (inputs(8)));
    layer0_outputs(6814) <= not(inputs(82));
    layer0_outputs(6815) <= not(inputs(149));
    layer0_outputs(6816) <= (inputs(163)) or (inputs(32));
    layer0_outputs(6817) <= (inputs(222)) and not (inputs(241));
    layer0_outputs(6818) <= (inputs(119)) or (inputs(120));
    layer0_outputs(6819) <= inputs(176);
    layer0_outputs(6820) <= not((inputs(23)) and (inputs(99)));
    layer0_outputs(6821) <= (inputs(108)) and not (inputs(160));
    layer0_outputs(6822) <= (inputs(103)) and not (inputs(109));
    layer0_outputs(6823) <= (inputs(71)) xor (inputs(84));
    layer0_outputs(6824) <= not(inputs(230)) or (inputs(168));
    layer0_outputs(6825) <= (inputs(156)) and not (inputs(148));
    layer0_outputs(6826) <= (inputs(154)) or (inputs(112));
    layer0_outputs(6827) <= not(inputs(195)) or (inputs(159));
    layer0_outputs(6828) <= not(inputs(64));
    layer0_outputs(6829) <= not(inputs(74)) or (inputs(255));
    layer0_outputs(6830) <= (inputs(34)) and not (inputs(235));
    layer0_outputs(6831) <= (inputs(3)) or (inputs(71));
    layer0_outputs(6832) <= (inputs(209)) or (inputs(124));
    layer0_outputs(6833) <= not(inputs(21));
    layer0_outputs(6834) <= not(inputs(227));
    layer0_outputs(6835) <= not(inputs(230)) or (inputs(5));
    layer0_outputs(6836) <= inputs(43);
    layer0_outputs(6837) <= not((inputs(44)) xor (inputs(17)));
    layer0_outputs(6838) <= not(inputs(156)) or (inputs(97));
    layer0_outputs(6839) <= not((inputs(211)) or (inputs(24)));
    layer0_outputs(6840) <= (inputs(76)) or (inputs(91));
    layer0_outputs(6841) <= not(inputs(26)) or (inputs(1));
    layer0_outputs(6842) <= (inputs(151)) and not (inputs(62));
    layer0_outputs(6843) <= not((inputs(93)) xor (inputs(154)));
    layer0_outputs(6844) <= not((inputs(6)) or (inputs(179)));
    layer0_outputs(6845) <= not(inputs(90)) or (inputs(85));
    layer0_outputs(6846) <= not((inputs(102)) and (inputs(218)));
    layer0_outputs(6847) <= inputs(36);
    layer0_outputs(6848) <= not(inputs(114));
    layer0_outputs(6849) <= (inputs(167)) and not (inputs(125));
    layer0_outputs(6850) <= not(inputs(231)) or (inputs(47));
    layer0_outputs(6851) <= not((inputs(228)) and (inputs(66)));
    layer0_outputs(6852) <= (inputs(230)) and not (inputs(20));
    layer0_outputs(6853) <= not(inputs(249)) or (inputs(99));
    layer0_outputs(6854) <= (inputs(7)) or (inputs(94));
    layer0_outputs(6855) <= (inputs(192)) and not (inputs(20));
    layer0_outputs(6856) <= (inputs(117)) and not (inputs(8));
    layer0_outputs(6857) <= not((inputs(42)) and (inputs(181)));
    layer0_outputs(6858) <= not(inputs(167)) or (inputs(228));
    layer0_outputs(6859) <= not(inputs(31));
    layer0_outputs(6860) <= (inputs(32)) or (inputs(180));
    layer0_outputs(6861) <= not(inputs(107));
    layer0_outputs(6862) <= (inputs(69)) xor (inputs(89));
    layer0_outputs(6863) <= (inputs(239)) xor (inputs(138));
    layer0_outputs(6864) <= (inputs(199)) and not (inputs(79));
    layer0_outputs(6865) <= not((inputs(164)) xor (inputs(240)));
    layer0_outputs(6866) <= not(inputs(227)) or (inputs(253));
    layer0_outputs(6867) <= not((inputs(118)) xor (inputs(88)));
    layer0_outputs(6868) <= (inputs(87)) and not (inputs(108));
    layer0_outputs(6869) <= inputs(116);
    layer0_outputs(6870) <= not(inputs(119));
    layer0_outputs(6871) <= '1';
    layer0_outputs(6872) <= (inputs(108)) and (inputs(1));
    layer0_outputs(6873) <= (inputs(17)) xor (inputs(130));
    layer0_outputs(6874) <= not(inputs(88)) or (inputs(78));
    layer0_outputs(6875) <= inputs(179);
    layer0_outputs(6876) <= not((inputs(158)) or (inputs(67)));
    layer0_outputs(6877) <= not(inputs(69));
    layer0_outputs(6878) <= inputs(220);
    layer0_outputs(6879) <= not(inputs(137)) or (inputs(53));
    layer0_outputs(6880) <= (inputs(137)) and not (inputs(128));
    layer0_outputs(6881) <= not(inputs(167)) or (inputs(29));
    layer0_outputs(6882) <= inputs(75);
    layer0_outputs(6883) <= not(inputs(73));
    layer0_outputs(6884) <= not(inputs(49)) or (inputs(237));
    layer0_outputs(6885) <= not((inputs(150)) xor (inputs(88)));
    layer0_outputs(6886) <= (inputs(87)) or (inputs(171));
    layer0_outputs(6887) <= not(inputs(120)) or (inputs(191));
    layer0_outputs(6888) <= '1';
    layer0_outputs(6889) <= not((inputs(141)) xor (inputs(246)));
    layer0_outputs(6890) <= not(inputs(89)) or (inputs(93));
    layer0_outputs(6891) <= (inputs(16)) or (inputs(123));
    layer0_outputs(6892) <= (inputs(74)) and not (inputs(6));
    layer0_outputs(6893) <= (inputs(168)) xor (inputs(87));
    layer0_outputs(6894) <= inputs(149);
    layer0_outputs(6895) <= not((inputs(203)) xor (inputs(246)));
    layer0_outputs(6896) <= not(inputs(114));
    layer0_outputs(6897) <= not(inputs(166)) or (inputs(12));
    layer0_outputs(6898) <= not(inputs(89)) or (inputs(103));
    layer0_outputs(6899) <= (inputs(5)) xor (inputs(76));
    layer0_outputs(6900) <= (inputs(192)) or (inputs(81));
    layer0_outputs(6901) <= (inputs(72)) xor (inputs(7));
    layer0_outputs(6902) <= not(inputs(71)) or (inputs(251));
    layer0_outputs(6903) <= not((inputs(114)) or (inputs(42)));
    layer0_outputs(6904) <= inputs(254);
    layer0_outputs(6905) <= (inputs(153)) and not (inputs(192));
    layer0_outputs(6906) <= not(inputs(0)) or (inputs(160));
    layer0_outputs(6907) <= (inputs(58)) or (inputs(81));
    layer0_outputs(6908) <= (inputs(19)) or (inputs(208));
    layer0_outputs(6909) <= inputs(247);
    layer0_outputs(6910) <= not((inputs(84)) and (inputs(201)));
    layer0_outputs(6911) <= not((inputs(77)) or (inputs(203)));
    layer0_outputs(6912) <= not(inputs(195));
    layer0_outputs(6913) <= not((inputs(105)) or (inputs(160)));
    layer0_outputs(6914) <= not((inputs(79)) or (inputs(177)));
    layer0_outputs(6915) <= not((inputs(33)) or (inputs(142)));
    layer0_outputs(6916) <= (inputs(133)) and not (inputs(17));
    layer0_outputs(6917) <= '1';
    layer0_outputs(6918) <= (inputs(48)) or (inputs(43));
    layer0_outputs(6919) <= not((inputs(166)) or (inputs(137)));
    layer0_outputs(6920) <= not(inputs(119)) or (inputs(2));
    layer0_outputs(6921) <= not((inputs(199)) or (inputs(207)));
    layer0_outputs(6922) <= inputs(90);
    layer0_outputs(6923) <= (inputs(49)) xor (inputs(77));
    layer0_outputs(6924) <= (inputs(197)) xor (inputs(217));
    layer0_outputs(6925) <= not((inputs(5)) or (inputs(214)));
    layer0_outputs(6926) <= inputs(69);
    layer0_outputs(6927) <= not(inputs(102));
    layer0_outputs(6928) <= inputs(6);
    layer0_outputs(6929) <= not((inputs(139)) and (inputs(171)));
    layer0_outputs(6930) <= not((inputs(162)) xor (inputs(224)));
    layer0_outputs(6931) <= (inputs(25)) or (inputs(7));
    layer0_outputs(6932) <= (inputs(151)) or (inputs(199));
    layer0_outputs(6933) <= inputs(106);
    layer0_outputs(6934) <= (inputs(122)) and not (inputs(129));
    layer0_outputs(6935) <= not(inputs(219));
    layer0_outputs(6936) <= (inputs(185)) and not (inputs(241));
    layer0_outputs(6937) <= inputs(20);
    layer0_outputs(6938) <= not(inputs(220)) or (inputs(96));
    layer0_outputs(6939) <= inputs(88);
    layer0_outputs(6940) <= not((inputs(106)) or (inputs(124)));
    layer0_outputs(6941) <= not((inputs(233)) xor (inputs(225)));
    layer0_outputs(6942) <= not(inputs(62)) or (inputs(9));
    layer0_outputs(6943) <= (inputs(149)) and not (inputs(90));
    layer0_outputs(6944) <= inputs(162);
    layer0_outputs(6945) <= (inputs(24)) and not (inputs(211));
    layer0_outputs(6946) <= (inputs(178)) or (inputs(93));
    layer0_outputs(6947) <= inputs(57);
    layer0_outputs(6948) <= not(inputs(250));
    layer0_outputs(6949) <= not((inputs(50)) or (inputs(46)));
    layer0_outputs(6950) <= inputs(94);
    layer0_outputs(6951) <= inputs(50);
    layer0_outputs(6952) <= not((inputs(190)) or (inputs(17)));
    layer0_outputs(6953) <= (inputs(255)) or (inputs(199));
    layer0_outputs(6954) <= not((inputs(227)) or (inputs(212)));
    layer0_outputs(6955) <= inputs(60);
    layer0_outputs(6956) <= inputs(178);
    layer0_outputs(6957) <= not(inputs(196));
    layer0_outputs(6958) <= not(inputs(188)) or (inputs(2));
    layer0_outputs(6959) <= not((inputs(28)) or (inputs(165)));
    layer0_outputs(6960) <= not((inputs(240)) or (inputs(236)));
    layer0_outputs(6961) <= inputs(152);
    layer0_outputs(6962) <= not((inputs(107)) xor (inputs(193)));
    layer0_outputs(6963) <= not(inputs(208));
    layer0_outputs(6964) <= not((inputs(212)) or (inputs(128)));
    layer0_outputs(6965) <= '0';
    layer0_outputs(6966) <= inputs(73);
    layer0_outputs(6967) <= (inputs(77)) xor (inputs(29));
    layer0_outputs(6968) <= (inputs(187)) and not (inputs(112));
    layer0_outputs(6969) <= inputs(114);
    layer0_outputs(6970) <= not(inputs(76));
    layer0_outputs(6971) <= not((inputs(194)) or (inputs(125)));
    layer0_outputs(6972) <= not((inputs(254)) or (inputs(223)));
    layer0_outputs(6973) <= not((inputs(2)) or (inputs(160)));
    layer0_outputs(6974) <= not((inputs(191)) xor (inputs(194)));
    layer0_outputs(6975) <= not((inputs(168)) or (inputs(89)));
    layer0_outputs(6976) <= not(inputs(41));
    layer0_outputs(6977) <= (inputs(128)) or (inputs(4));
    layer0_outputs(6978) <= not((inputs(196)) or (inputs(216)));
    layer0_outputs(6979) <= (inputs(112)) and (inputs(190));
    layer0_outputs(6980) <= not(inputs(5));
    layer0_outputs(6981) <= inputs(189);
    layer0_outputs(6982) <= (inputs(141)) or (inputs(161));
    layer0_outputs(6983) <= not(inputs(224));
    layer0_outputs(6984) <= inputs(14);
    layer0_outputs(6985) <= not((inputs(235)) or (inputs(211)));
    layer0_outputs(6986) <= not(inputs(22));
    layer0_outputs(6987) <= inputs(94);
    layer0_outputs(6988) <= not((inputs(38)) xor (inputs(146)));
    layer0_outputs(6989) <= (inputs(129)) and not (inputs(192));
    layer0_outputs(6990) <= not(inputs(21)) or (inputs(140));
    layer0_outputs(6991) <= not(inputs(228)) or (inputs(107));
    layer0_outputs(6992) <= inputs(135);
    layer0_outputs(6993) <= inputs(115);
    layer0_outputs(6994) <= not(inputs(90)) or (inputs(176));
    layer0_outputs(6995) <= not(inputs(249));
    layer0_outputs(6996) <= not(inputs(101));
    layer0_outputs(6997) <= not(inputs(217));
    layer0_outputs(6998) <= not(inputs(27)) or (inputs(117));
    layer0_outputs(6999) <= not((inputs(209)) and (inputs(43)));
    layer0_outputs(7000) <= not(inputs(165));
    layer0_outputs(7001) <= not((inputs(157)) or (inputs(98)));
    layer0_outputs(7002) <= not(inputs(229));
    layer0_outputs(7003) <= not((inputs(57)) and (inputs(182)));
    layer0_outputs(7004) <= inputs(149);
    layer0_outputs(7005) <= (inputs(222)) or (inputs(138));
    layer0_outputs(7006) <= (inputs(166)) and not (inputs(34));
    layer0_outputs(7007) <= (inputs(49)) xor (inputs(4));
    layer0_outputs(7008) <= (inputs(210)) and not (inputs(125));
    layer0_outputs(7009) <= not(inputs(101));
    layer0_outputs(7010) <= inputs(90);
    layer0_outputs(7011) <= (inputs(201)) or (inputs(196));
    layer0_outputs(7012) <= not((inputs(177)) xor (inputs(197)));
    layer0_outputs(7013) <= (inputs(57)) or (inputs(17));
    layer0_outputs(7014) <= inputs(109);
    layer0_outputs(7015) <= (inputs(15)) and not (inputs(217));
    layer0_outputs(7016) <= (inputs(42)) and not (inputs(96));
    layer0_outputs(7017) <= inputs(107);
    layer0_outputs(7018) <= inputs(132);
    layer0_outputs(7019) <= (inputs(245)) or (inputs(219));
    layer0_outputs(7020) <= inputs(156);
    layer0_outputs(7021) <= inputs(3);
    layer0_outputs(7022) <= inputs(145);
    layer0_outputs(7023) <= not((inputs(30)) or (inputs(85)));
    layer0_outputs(7024) <= not(inputs(240));
    layer0_outputs(7025) <= inputs(163);
    layer0_outputs(7026) <= not((inputs(222)) xor (inputs(106)));
    layer0_outputs(7027) <= '0';
    layer0_outputs(7028) <= inputs(99);
    layer0_outputs(7029) <= inputs(167);
    layer0_outputs(7030) <= not((inputs(176)) xor (inputs(27)));
    layer0_outputs(7031) <= not((inputs(51)) xor (inputs(197)));
    layer0_outputs(7032) <= not((inputs(175)) or (inputs(218)));
    layer0_outputs(7033) <= inputs(132);
    layer0_outputs(7034) <= (inputs(148)) and not (inputs(8));
    layer0_outputs(7035) <= not(inputs(44));
    layer0_outputs(7036) <= (inputs(19)) and not (inputs(129));
    layer0_outputs(7037) <= '1';
    layer0_outputs(7038) <= (inputs(222)) or (inputs(212));
    layer0_outputs(7039) <= not(inputs(149));
    layer0_outputs(7040) <= not(inputs(53)) or (inputs(56));
    layer0_outputs(7041) <= (inputs(77)) and (inputs(43));
    layer0_outputs(7042) <= (inputs(111)) and not (inputs(140));
    layer0_outputs(7043) <= not(inputs(38));
    layer0_outputs(7044) <= inputs(194);
    layer0_outputs(7045) <= not(inputs(99));
    layer0_outputs(7046) <= (inputs(124)) and (inputs(162));
    layer0_outputs(7047) <= not((inputs(96)) xor (inputs(228)));
    layer0_outputs(7048) <= inputs(233);
    layer0_outputs(7049) <= (inputs(226)) and not (inputs(27));
    layer0_outputs(7050) <= (inputs(206)) or (inputs(49));
    layer0_outputs(7051) <= not((inputs(157)) xor (inputs(154)));
    layer0_outputs(7052) <= not(inputs(89)) or (inputs(51));
    layer0_outputs(7053) <= not(inputs(7)) or (inputs(218));
    layer0_outputs(7054) <= (inputs(94)) xor (inputs(128));
    layer0_outputs(7055) <= not(inputs(114));
    layer0_outputs(7056) <= not((inputs(59)) or (inputs(160)));
    layer0_outputs(7057) <= (inputs(67)) or (inputs(97));
    layer0_outputs(7058) <= inputs(208);
    layer0_outputs(7059) <= inputs(181);
    layer0_outputs(7060) <= inputs(42);
    layer0_outputs(7061) <= (inputs(63)) or (inputs(38));
    layer0_outputs(7062) <= (inputs(165)) and not (inputs(205));
    layer0_outputs(7063) <= inputs(107);
    layer0_outputs(7064) <= not(inputs(74)) or (inputs(178));
    layer0_outputs(7065) <= not((inputs(144)) or (inputs(226)));
    layer0_outputs(7066) <= not((inputs(96)) or (inputs(101)));
    layer0_outputs(7067) <= not(inputs(100));
    layer0_outputs(7068) <= not((inputs(108)) or (inputs(75)));
    layer0_outputs(7069) <= not(inputs(46)) or (inputs(159));
    layer0_outputs(7070) <= not((inputs(251)) xor (inputs(11)));
    layer0_outputs(7071) <= (inputs(210)) and not (inputs(16));
    layer0_outputs(7072) <= (inputs(67)) and not (inputs(110));
    layer0_outputs(7073) <= not(inputs(114)) or (inputs(102));
    layer0_outputs(7074) <= not((inputs(66)) and (inputs(184)));
    layer0_outputs(7075) <= '1';
    layer0_outputs(7076) <= not(inputs(167)) or (inputs(128));
    layer0_outputs(7077) <= not((inputs(143)) or (inputs(131)));
    layer0_outputs(7078) <= inputs(164);
    layer0_outputs(7079) <= inputs(135);
    layer0_outputs(7080) <= inputs(113);
    layer0_outputs(7081) <= '1';
    layer0_outputs(7082) <= not(inputs(137)) or (inputs(160));
    layer0_outputs(7083) <= not((inputs(107)) xor (inputs(117)));
    layer0_outputs(7084) <= not((inputs(85)) or (inputs(157)));
    layer0_outputs(7085) <= not((inputs(93)) or (inputs(233)));
    layer0_outputs(7086) <= not(inputs(166));
    layer0_outputs(7087) <= not(inputs(229)) or (inputs(59));
    layer0_outputs(7088) <= inputs(115);
    layer0_outputs(7089) <= not(inputs(105));
    layer0_outputs(7090) <= not((inputs(131)) or (inputs(2)));
    layer0_outputs(7091) <= not(inputs(213)) or (inputs(127));
    layer0_outputs(7092) <= not(inputs(76)) or (inputs(190));
    layer0_outputs(7093) <= not(inputs(61));
    layer0_outputs(7094) <= not(inputs(230));
    layer0_outputs(7095) <= (inputs(73)) and (inputs(103));
    layer0_outputs(7096) <= not(inputs(172));
    layer0_outputs(7097) <= (inputs(226)) xor (inputs(222));
    layer0_outputs(7098) <= inputs(85);
    layer0_outputs(7099) <= (inputs(48)) or (inputs(47));
    layer0_outputs(7100) <= not((inputs(135)) xor (inputs(243)));
    layer0_outputs(7101) <= (inputs(95)) and not (inputs(34));
    layer0_outputs(7102) <= (inputs(124)) and not (inputs(226));
    layer0_outputs(7103) <= not((inputs(246)) and (inputs(228)));
    layer0_outputs(7104) <= (inputs(116)) or (inputs(253));
    layer0_outputs(7105) <= not(inputs(63)) or (inputs(16));
    layer0_outputs(7106) <= not(inputs(63));
    layer0_outputs(7107) <= not((inputs(198)) xor (inputs(23)));
    layer0_outputs(7108) <= inputs(101);
    layer0_outputs(7109) <= inputs(13);
    layer0_outputs(7110) <= not((inputs(31)) xor (inputs(165)));
    layer0_outputs(7111) <= not(inputs(212));
    layer0_outputs(7112) <= inputs(248);
    layer0_outputs(7113) <= (inputs(120)) or (inputs(47));
    layer0_outputs(7114) <= not((inputs(95)) or (inputs(86)));
    layer0_outputs(7115) <= not((inputs(7)) or (inputs(242)));
    layer0_outputs(7116) <= (inputs(36)) and not (inputs(156));
    layer0_outputs(7117) <= (inputs(104)) and not (inputs(1));
    layer0_outputs(7118) <= not(inputs(107));
    layer0_outputs(7119) <= (inputs(233)) or (inputs(87));
    layer0_outputs(7120) <= not((inputs(124)) xor (inputs(88)));
    layer0_outputs(7121) <= not(inputs(197)) or (inputs(223));
    layer0_outputs(7122) <= (inputs(29)) xor (inputs(62));
    layer0_outputs(7123) <= (inputs(125)) or (inputs(208));
    layer0_outputs(7124) <= not(inputs(104)) or (inputs(31));
    layer0_outputs(7125) <= (inputs(194)) and not (inputs(15));
    layer0_outputs(7126) <= not((inputs(168)) or (inputs(251)));
    layer0_outputs(7127) <= inputs(22);
    layer0_outputs(7128) <= not((inputs(180)) or (inputs(229)));
    layer0_outputs(7129) <= not(inputs(102));
    layer0_outputs(7130) <= (inputs(217)) xor (inputs(6));
    layer0_outputs(7131) <= (inputs(45)) xor (inputs(157));
    layer0_outputs(7132) <= not(inputs(59)) or (inputs(250));
    layer0_outputs(7133) <= '1';
    layer0_outputs(7134) <= not((inputs(126)) and (inputs(237)));
    layer0_outputs(7135) <= not((inputs(160)) or (inputs(178)));
    layer0_outputs(7136) <= not((inputs(128)) xor (inputs(84)));
    layer0_outputs(7137) <= inputs(85);
    layer0_outputs(7138) <= not(inputs(229)) or (inputs(74));
    layer0_outputs(7139) <= not((inputs(48)) or (inputs(23)));
    layer0_outputs(7140) <= (inputs(0)) xor (inputs(170));
    layer0_outputs(7141) <= not(inputs(133));
    layer0_outputs(7142) <= inputs(233);
    layer0_outputs(7143) <= not(inputs(165));
    layer0_outputs(7144) <= not(inputs(95)) or (inputs(62));
    layer0_outputs(7145) <= (inputs(235)) and not (inputs(145));
    layer0_outputs(7146) <= (inputs(13)) or (inputs(220));
    layer0_outputs(7147) <= not(inputs(162));
    layer0_outputs(7148) <= not((inputs(55)) and (inputs(70)));
    layer0_outputs(7149) <= not(inputs(22)) or (inputs(238));
    layer0_outputs(7150) <= not(inputs(101));
    layer0_outputs(7151) <= not(inputs(23));
    layer0_outputs(7152) <= not(inputs(7));
    layer0_outputs(7153) <= inputs(115);
    layer0_outputs(7154) <= (inputs(26)) and (inputs(27));
    layer0_outputs(7155) <= not(inputs(165));
    layer0_outputs(7156) <= inputs(24);
    layer0_outputs(7157) <= not((inputs(72)) or (inputs(159)));
    layer0_outputs(7158) <= inputs(24);
    layer0_outputs(7159) <= '0';
    layer0_outputs(7160) <= not(inputs(112));
    layer0_outputs(7161) <= (inputs(214)) and not (inputs(110));
    layer0_outputs(7162) <= not(inputs(138)) or (inputs(214));
    layer0_outputs(7163) <= (inputs(54)) xor (inputs(58));
    layer0_outputs(7164) <= not((inputs(216)) or (inputs(113)));
    layer0_outputs(7165) <= inputs(150);
    layer0_outputs(7166) <= not(inputs(209)) or (inputs(160));
    layer0_outputs(7167) <= not((inputs(42)) and (inputs(45)));
    layer0_outputs(7168) <= (inputs(254)) and not (inputs(241));
    layer0_outputs(7169) <= (inputs(43)) xor (inputs(18));
    layer0_outputs(7170) <= (inputs(28)) xor (inputs(13));
    layer0_outputs(7171) <= not((inputs(131)) xor (inputs(31)));
    layer0_outputs(7172) <= not(inputs(62)) or (inputs(20));
    layer0_outputs(7173) <= inputs(154);
    layer0_outputs(7174) <= (inputs(87)) or (inputs(37));
    layer0_outputs(7175) <= (inputs(0)) xor (inputs(32));
    layer0_outputs(7176) <= not((inputs(144)) or (inputs(107)));
    layer0_outputs(7177) <= (inputs(151)) and not (inputs(116));
    layer0_outputs(7178) <= not(inputs(76));
    layer0_outputs(7179) <= inputs(191);
    layer0_outputs(7180) <= not(inputs(157)) or (inputs(239));
    layer0_outputs(7181) <= (inputs(88)) and not (inputs(208));
    layer0_outputs(7182) <= (inputs(128)) and not (inputs(240));
    layer0_outputs(7183) <= '1';
    layer0_outputs(7184) <= (inputs(28)) and not (inputs(201));
    layer0_outputs(7185) <= not(inputs(27)) or (inputs(33));
    layer0_outputs(7186) <= not((inputs(96)) or (inputs(69)));
    layer0_outputs(7187) <= (inputs(159)) and not (inputs(128));
    layer0_outputs(7188) <= not((inputs(189)) or (inputs(232)));
    layer0_outputs(7189) <= not((inputs(49)) or (inputs(185)));
    layer0_outputs(7190) <= (inputs(250)) xor (inputs(210));
    layer0_outputs(7191) <= (inputs(175)) xor (inputs(222));
    layer0_outputs(7192) <= not((inputs(223)) or (inputs(122)));
    layer0_outputs(7193) <= not(inputs(212));
    layer0_outputs(7194) <= not((inputs(243)) or (inputs(167)));
    layer0_outputs(7195) <= not(inputs(87));
    layer0_outputs(7196) <= inputs(45);
    layer0_outputs(7197) <= not(inputs(215));
    layer0_outputs(7198) <= (inputs(108)) xor (inputs(135));
    layer0_outputs(7199) <= not(inputs(182));
    layer0_outputs(7200) <= not(inputs(102)) or (inputs(147));
    layer0_outputs(7201) <= not(inputs(74));
    layer0_outputs(7202) <= (inputs(101)) and (inputs(201));
    layer0_outputs(7203) <= inputs(121);
    layer0_outputs(7204) <= inputs(115);
    layer0_outputs(7205) <= inputs(147);
    layer0_outputs(7206) <= inputs(164);
    layer0_outputs(7207) <= '0';
    layer0_outputs(7208) <= (inputs(133)) and not (inputs(17));
    layer0_outputs(7209) <= not(inputs(114));
    layer0_outputs(7210) <= (inputs(112)) xor (inputs(209));
    layer0_outputs(7211) <= not((inputs(191)) xor (inputs(20)));
    layer0_outputs(7212) <= (inputs(133)) or (inputs(247));
    layer0_outputs(7213) <= not((inputs(171)) or (inputs(5)));
    layer0_outputs(7214) <= not(inputs(182)) or (inputs(85));
    layer0_outputs(7215) <= inputs(146);
    layer0_outputs(7216) <= not((inputs(80)) xor (inputs(70)));
    layer0_outputs(7217) <= (inputs(50)) and not (inputs(243));
    layer0_outputs(7218) <= (inputs(59)) or (inputs(63));
    layer0_outputs(7219) <= not(inputs(81));
    layer0_outputs(7220) <= (inputs(243)) and not (inputs(2));
    layer0_outputs(7221) <= not((inputs(162)) or (inputs(33)));
    layer0_outputs(7222) <= (inputs(189)) xor (inputs(115));
    layer0_outputs(7223) <= not(inputs(67));
    layer0_outputs(7224) <= not(inputs(72)) or (inputs(221));
    layer0_outputs(7225) <= (inputs(80)) or (inputs(52));
    layer0_outputs(7226) <= not(inputs(253));
    layer0_outputs(7227) <= inputs(100);
    layer0_outputs(7228) <= not(inputs(227));
    layer0_outputs(7229) <= '0';
    layer0_outputs(7230) <= (inputs(253)) xor (inputs(202));
    layer0_outputs(7231) <= inputs(186);
    layer0_outputs(7232) <= not((inputs(118)) xor (inputs(93)));
    layer0_outputs(7233) <= not((inputs(122)) xor (inputs(86)));
    layer0_outputs(7234) <= inputs(138);
    layer0_outputs(7235) <= inputs(57);
    layer0_outputs(7236) <= not(inputs(151)) or (inputs(179));
    layer0_outputs(7237) <= not(inputs(220));
    layer0_outputs(7238) <= (inputs(37)) xor (inputs(6));
    layer0_outputs(7239) <= (inputs(210)) and not (inputs(46));
    layer0_outputs(7240) <= (inputs(168)) and not (inputs(35));
    layer0_outputs(7241) <= (inputs(18)) and not (inputs(118));
    layer0_outputs(7242) <= inputs(153);
    layer0_outputs(7243) <= '0';
    layer0_outputs(7244) <= inputs(214);
    layer0_outputs(7245) <= inputs(82);
    layer0_outputs(7246) <= not((inputs(182)) xor (inputs(55)));
    layer0_outputs(7247) <= not(inputs(24)) or (inputs(141));
    layer0_outputs(7248) <= not(inputs(44));
    layer0_outputs(7249) <= inputs(216);
    layer0_outputs(7250) <= inputs(201);
    layer0_outputs(7251) <= not(inputs(17));
    layer0_outputs(7252) <= inputs(25);
    layer0_outputs(7253) <= not(inputs(47));
    layer0_outputs(7254) <= (inputs(232)) and not (inputs(112));
    layer0_outputs(7255) <= inputs(136);
    layer0_outputs(7256) <= not((inputs(221)) xor (inputs(105)));
    layer0_outputs(7257) <= (inputs(152)) and not (inputs(221));
    layer0_outputs(7258) <= '1';
    layer0_outputs(7259) <= not((inputs(251)) or (inputs(242)));
    layer0_outputs(7260) <= inputs(117);
    layer0_outputs(7261) <= not(inputs(233)) or (inputs(128));
    layer0_outputs(7262) <= not(inputs(64)) or (inputs(185));
    layer0_outputs(7263) <= inputs(207);
    layer0_outputs(7264) <= (inputs(10)) or (inputs(14));
    layer0_outputs(7265) <= (inputs(21)) and not (inputs(128));
    layer0_outputs(7266) <= (inputs(14)) or (inputs(213));
    layer0_outputs(7267) <= inputs(163);
    layer0_outputs(7268) <= not(inputs(200));
    layer0_outputs(7269) <= (inputs(233)) and not (inputs(73));
    layer0_outputs(7270) <= not(inputs(34)) or (inputs(16));
    layer0_outputs(7271) <= not(inputs(83)) or (inputs(234));
    layer0_outputs(7272) <= (inputs(146)) or (inputs(89));
    layer0_outputs(7273) <= not(inputs(195));
    layer0_outputs(7274) <= (inputs(105)) xor (inputs(173));
    layer0_outputs(7275) <= not(inputs(103));
    layer0_outputs(7276) <= not((inputs(116)) xor (inputs(81)));
    layer0_outputs(7277) <= (inputs(92)) or (inputs(178));
    layer0_outputs(7278) <= not((inputs(50)) xor (inputs(234)));
    layer0_outputs(7279) <= not(inputs(70)) or (inputs(94));
    layer0_outputs(7280) <= not(inputs(215));
    layer0_outputs(7281) <= (inputs(219)) or (inputs(218));
    layer0_outputs(7282) <= not(inputs(239));
    layer0_outputs(7283) <= not(inputs(87));
    layer0_outputs(7284) <= not((inputs(13)) xor (inputs(87)));
    layer0_outputs(7285) <= not(inputs(230));
    layer0_outputs(7286) <= not(inputs(179));
    layer0_outputs(7287) <= not((inputs(53)) xor (inputs(71)));
    layer0_outputs(7288) <= (inputs(59)) and not (inputs(220));
    layer0_outputs(7289) <= not(inputs(83)) or (inputs(111));
    layer0_outputs(7290) <= (inputs(105)) xor (inputs(167));
    layer0_outputs(7291) <= not(inputs(105));
    layer0_outputs(7292) <= not((inputs(79)) xor (inputs(175)));
    layer0_outputs(7293) <= (inputs(225)) xor (inputs(36));
    layer0_outputs(7294) <= not(inputs(158));
    layer0_outputs(7295) <= (inputs(63)) or (inputs(43));
    layer0_outputs(7296) <= inputs(89);
    layer0_outputs(7297) <= not((inputs(23)) xor (inputs(219)));
    layer0_outputs(7298) <= inputs(21);
    layer0_outputs(7299) <= not((inputs(64)) or (inputs(242)));
    layer0_outputs(7300) <= (inputs(194)) and not (inputs(36));
    layer0_outputs(7301) <= not((inputs(71)) and (inputs(234)));
    layer0_outputs(7302) <= not(inputs(170)) or (inputs(28));
    layer0_outputs(7303) <= not(inputs(81)) or (inputs(70));
    layer0_outputs(7304) <= not(inputs(174)) or (inputs(19));
    layer0_outputs(7305) <= inputs(98);
    layer0_outputs(7306) <= not(inputs(235)) or (inputs(0));
    layer0_outputs(7307) <= inputs(60);
    layer0_outputs(7308) <= not((inputs(6)) xor (inputs(175)));
    layer0_outputs(7309) <= not(inputs(189));
    layer0_outputs(7310) <= (inputs(87)) and not (inputs(0));
    layer0_outputs(7311) <= not(inputs(75)) or (inputs(127));
    layer0_outputs(7312) <= not(inputs(90)) or (inputs(196));
    layer0_outputs(7313) <= inputs(98);
    layer0_outputs(7314) <= not(inputs(165));
    layer0_outputs(7315) <= (inputs(94)) and not (inputs(32));
    layer0_outputs(7316) <= (inputs(254)) or (inputs(111));
    layer0_outputs(7317) <= inputs(177);
    layer0_outputs(7318) <= (inputs(139)) or (inputs(2));
    layer0_outputs(7319) <= (inputs(52)) or (inputs(106));
    layer0_outputs(7320) <= (inputs(216)) and (inputs(175));
    layer0_outputs(7321) <= inputs(161);
    layer0_outputs(7322) <= (inputs(203)) or (inputs(21));
    layer0_outputs(7323) <= (inputs(164)) or (inputs(33));
    layer0_outputs(7324) <= not(inputs(96));
    layer0_outputs(7325) <= inputs(212);
    layer0_outputs(7326) <= inputs(217);
    layer0_outputs(7327) <= (inputs(140)) or (inputs(56));
    layer0_outputs(7328) <= (inputs(24)) and not (inputs(193));
    layer0_outputs(7329) <= (inputs(116)) and not (inputs(108));
    layer0_outputs(7330) <= (inputs(136)) and (inputs(134));
    layer0_outputs(7331) <= inputs(179);
    layer0_outputs(7332) <= not(inputs(98));
    layer0_outputs(7333) <= not(inputs(205));
    layer0_outputs(7334) <= (inputs(8)) and (inputs(90));
    layer0_outputs(7335) <= '0';
    layer0_outputs(7336) <= (inputs(16)) or (inputs(164));
    layer0_outputs(7337) <= not((inputs(189)) xor (inputs(87)));
    layer0_outputs(7338) <= not(inputs(199)) or (inputs(80));
    layer0_outputs(7339) <= (inputs(139)) and not (inputs(39));
    layer0_outputs(7340) <= (inputs(100)) and not (inputs(126));
    layer0_outputs(7341) <= '1';
    layer0_outputs(7342) <= (inputs(56)) xor (inputs(20));
    layer0_outputs(7343) <= inputs(119);
    layer0_outputs(7344) <= not((inputs(73)) or (inputs(226)));
    layer0_outputs(7345) <= not((inputs(104)) or (inputs(135)));
    layer0_outputs(7346) <= not(inputs(237));
    layer0_outputs(7347) <= not(inputs(216));
    layer0_outputs(7348) <= not(inputs(98));
    layer0_outputs(7349) <= inputs(211);
    layer0_outputs(7350) <= (inputs(194)) and not (inputs(47));
    layer0_outputs(7351) <= not(inputs(75)) or (inputs(160));
    layer0_outputs(7352) <= (inputs(136)) and not (inputs(217));
    layer0_outputs(7353) <= not(inputs(214));
    layer0_outputs(7354) <= not((inputs(118)) or (inputs(30)));
    layer0_outputs(7355) <= (inputs(219)) and not (inputs(50));
    layer0_outputs(7356) <= inputs(120);
    layer0_outputs(7357) <= not(inputs(64));
    layer0_outputs(7358) <= inputs(162);
    layer0_outputs(7359) <= (inputs(105)) xor (inputs(93));
    layer0_outputs(7360) <= not(inputs(106));
    layer0_outputs(7361) <= not(inputs(251));
    layer0_outputs(7362) <= inputs(27);
    layer0_outputs(7363) <= not((inputs(127)) or (inputs(238)));
    layer0_outputs(7364) <= not(inputs(88));
    layer0_outputs(7365) <= not(inputs(101));
    layer0_outputs(7366) <= (inputs(26)) xor (inputs(0));
    layer0_outputs(7367) <= (inputs(122)) xor (inputs(111));
    layer0_outputs(7368) <= not((inputs(169)) and (inputs(70)));
    layer0_outputs(7369) <= not((inputs(4)) or (inputs(202)));
    layer0_outputs(7370) <= (inputs(244)) and not (inputs(240));
    layer0_outputs(7371) <= not(inputs(78));
    layer0_outputs(7372) <= (inputs(36)) or (inputs(228));
    layer0_outputs(7373) <= inputs(242);
    layer0_outputs(7374) <= (inputs(38)) and not (inputs(250));
    layer0_outputs(7375) <= (inputs(133)) and not (inputs(22));
    layer0_outputs(7376) <= (inputs(9)) and not (inputs(64));
    layer0_outputs(7377) <= (inputs(248)) or (inputs(163));
    layer0_outputs(7378) <= not(inputs(90));
    layer0_outputs(7379) <= not((inputs(252)) or (inputs(239)));
    layer0_outputs(7380) <= (inputs(121)) and not (inputs(202));
    layer0_outputs(7381) <= (inputs(58)) and not (inputs(171));
    layer0_outputs(7382) <= not((inputs(89)) or (inputs(16)));
    layer0_outputs(7383) <= (inputs(203)) and (inputs(163));
    layer0_outputs(7384) <= inputs(129);
    layer0_outputs(7385) <= not((inputs(54)) and (inputs(41)));
    layer0_outputs(7386) <= (inputs(132)) and not (inputs(89));
    layer0_outputs(7387) <= not((inputs(152)) xor (inputs(145)));
    layer0_outputs(7388) <= not(inputs(87));
    layer0_outputs(7389) <= not(inputs(240));
    layer0_outputs(7390) <= not(inputs(124)) or (inputs(235));
    layer0_outputs(7391) <= inputs(47);
    layer0_outputs(7392) <= (inputs(147)) or (inputs(9));
    layer0_outputs(7393) <= not(inputs(165));
    layer0_outputs(7394) <= not(inputs(122)) or (inputs(143));
    layer0_outputs(7395) <= inputs(68);
    layer0_outputs(7396) <= not(inputs(128)) or (inputs(240));
    layer0_outputs(7397) <= (inputs(68)) and not (inputs(177));
    layer0_outputs(7398) <= (inputs(133)) and not (inputs(96));
    layer0_outputs(7399) <= not(inputs(194));
    layer0_outputs(7400) <= not((inputs(174)) or (inputs(110)));
    layer0_outputs(7401) <= (inputs(202)) and not (inputs(128));
    layer0_outputs(7402) <= inputs(18);
    layer0_outputs(7403) <= (inputs(156)) or (inputs(159));
    layer0_outputs(7404) <= inputs(210);
    layer0_outputs(7405) <= not((inputs(252)) and (inputs(113)));
    layer0_outputs(7406) <= not(inputs(159));
    layer0_outputs(7407) <= not((inputs(138)) or (inputs(16)));
    layer0_outputs(7408) <= (inputs(7)) or (inputs(24));
    layer0_outputs(7409) <= not(inputs(141));
    layer0_outputs(7410) <= not((inputs(112)) or (inputs(209)));
    layer0_outputs(7411) <= inputs(146);
    layer0_outputs(7412) <= not((inputs(79)) xor (inputs(31)));
    layer0_outputs(7413) <= (inputs(216)) or (inputs(56));
    layer0_outputs(7414) <= not(inputs(81));
    layer0_outputs(7415) <= inputs(91);
    layer0_outputs(7416) <= not(inputs(55)) or (inputs(177));
    layer0_outputs(7417) <= not(inputs(228));
    layer0_outputs(7418) <= (inputs(236)) or (inputs(181));
    layer0_outputs(7419) <= inputs(109);
    layer0_outputs(7420) <= inputs(77);
    layer0_outputs(7421) <= not(inputs(152));
    layer0_outputs(7422) <= not(inputs(137));
    layer0_outputs(7423) <= inputs(151);
    layer0_outputs(7424) <= not(inputs(171)) or (inputs(13));
    layer0_outputs(7425) <= not((inputs(169)) or (inputs(48)));
    layer0_outputs(7426) <= not((inputs(201)) and (inputs(216)));
    layer0_outputs(7427) <= inputs(45);
    layer0_outputs(7428) <= (inputs(41)) xor (inputs(119));
    layer0_outputs(7429) <= (inputs(38)) or (inputs(125));
    layer0_outputs(7430) <= not(inputs(83));
    layer0_outputs(7431) <= (inputs(197)) and (inputs(9));
    layer0_outputs(7432) <= (inputs(95)) or (inputs(60));
    layer0_outputs(7433) <= (inputs(4)) xor (inputs(108));
    layer0_outputs(7434) <= not(inputs(196)) or (inputs(69));
    layer0_outputs(7435) <= not((inputs(102)) xor (inputs(150)));
    layer0_outputs(7436) <= not(inputs(84));
    layer0_outputs(7437) <= (inputs(214)) or (inputs(14));
    layer0_outputs(7438) <= inputs(124);
    layer0_outputs(7439) <= (inputs(98)) and not (inputs(55));
    layer0_outputs(7440) <= inputs(101);
    layer0_outputs(7441) <= (inputs(118)) or (inputs(188));
    layer0_outputs(7442) <= not(inputs(163));
    layer0_outputs(7443) <= not((inputs(51)) or (inputs(173)));
    layer0_outputs(7444) <= (inputs(15)) or (inputs(124));
    layer0_outputs(7445) <= not(inputs(162));
    layer0_outputs(7446) <= (inputs(216)) xor (inputs(178));
    layer0_outputs(7447) <= not((inputs(100)) or (inputs(85)));
    layer0_outputs(7448) <= (inputs(80)) or (inputs(225));
    layer0_outputs(7449) <= not((inputs(236)) xor (inputs(203)));
    layer0_outputs(7450) <= not(inputs(102)) or (inputs(255));
    layer0_outputs(7451) <= (inputs(99)) and (inputs(137));
    layer0_outputs(7452) <= (inputs(45)) xor (inputs(34));
    layer0_outputs(7453) <= not(inputs(156)) or (inputs(80));
    layer0_outputs(7454) <= not((inputs(204)) or (inputs(155)));
    layer0_outputs(7455) <= not((inputs(230)) xor (inputs(90)));
    layer0_outputs(7456) <= inputs(140);
    layer0_outputs(7457) <= inputs(229);
    layer0_outputs(7458) <= inputs(230);
    layer0_outputs(7459) <= not(inputs(202));
    layer0_outputs(7460) <= inputs(209);
    layer0_outputs(7461) <= not((inputs(176)) or (inputs(212)));
    layer0_outputs(7462) <= not(inputs(171)) or (inputs(98));
    layer0_outputs(7463) <= (inputs(90)) xor (inputs(63));
    layer0_outputs(7464) <= (inputs(210)) xor (inputs(219));
    layer0_outputs(7465) <= (inputs(124)) xor (inputs(190));
    layer0_outputs(7466) <= (inputs(179)) xor (inputs(113));
    layer0_outputs(7467) <= (inputs(68)) and (inputs(193));
    layer0_outputs(7468) <= '0';
    layer0_outputs(7469) <= not(inputs(210));
    layer0_outputs(7470) <= not((inputs(48)) or (inputs(36)));
    layer0_outputs(7471) <= not((inputs(117)) or (inputs(252)));
    layer0_outputs(7472) <= inputs(147);
    layer0_outputs(7473) <= (inputs(206)) or (inputs(171));
    layer0_outputs(7474) <= inputs(37);
    layer0_outputs(7475) <= not((inputs(206)) xor (inputs(47)));
    layer0_outputs(7476) <= not((inputs(117)) or (inputs(81)));
    layer0_outputs(7477) <= not((inputs(29)) or (inputs(110)));
    layer0_outputs(7478) <= not(inputs(156));
    layer0_outputs(7479) <= inputs(113);
    layer0_outputs(7480) <= not(inputs(60));
    layer0_outputs(7481) <= (inputs(136)) and not (inputs(210));
    layer0_outputs(7482) <= not(inputs(105)) or (inputs(0));
    layer0_outputs(7483) <= not(inputs(77));
    layer0_outputs(7484) <= (inputs(24)) or (inputs(1));
    layer0_outputs(7485) <= not(inputs(239)) or (inputs(188));
    layer0_outputs(7486) <= not(inputs(55));
    layer0_outputs(7487) <= not(inputs(103));
    layer0_outputs(7488) <= (inputs(36)) xor (inputs(75));
    layer0_outputs(7489) <= inputs(23);
    layer0_outputs(7490) <= (inputs(245)) or (inputs(112));
    layer0_outputs(7491) <= not(inputs(174));
    layer0_outputs(7492) <= inputs(62);
    layer0_outputs(7493) <= (inputs(153)) or (inputs(127));
    layer0_outputs(7494) <= not((inputs(236)) or (inputs(140)));
    layer0_outputs(7495) <= not(inputs(147));
    layer0_outputs(7496) <= not(inputs(140));
    layer0_outputs(7497) <= (inputs(232)) xor (inputs(90));
    layer0_outputs(7498) <= not((inputs(73)) or (inputs(54)));
    layer0_outputs(7499) <= not((inputs(140)) xor (inputs(88)));
    layer0_outputs(7500) <= '1';
    layer0_outputs(7501) <= not(inputs(114)) or (inputs(89));
    layer0_outputs(7502) <= not((inputs(215)) xor (inputs(254)));
    layer0_outputs(7503) <= (inputs(39)) or (inputs(33));
    layer0_outputs(7504) <= (inputs(12)) and not (inputs(95));
    layer0_outputs(7505) <= (inputs(82)) and not (inputs(223));
    layer0_outputs(7506) <= inputs(84);
    layer0_outputs(7507) <= (inputs(29)) and not (inputs(109));
    layer0_outputs(7508) <= inputs(86);
    layer0_outputs(7509) <= not(inputs(122)) or (inputs(196));
    layer0_outputs(7510) <= not(inputs(109)) or (inputs(198));
    layer0_outputs(7511) <= (inputs(26)) and (inputs(110));
    layer0_outputs(7512) <= not(inputs(58));
    layer0_outputs(7513) <= not(inputs(203)) or (inputs(202));
    layer0_outputs(7514) <= not(inputs(153));
    layer0_outputs(7515) <= (inputs(119)) and not (inputs(235));
    layer0_outputs(7516) <= not(inputs(198));
    layer0_outputs(7517) <= inputs(187);
    layer0_outputs(7518) <= (inputs(151)) and not (inputs(82));
    layer0_outputs(7519) <= not((inputs(188)) or (inputs(212)));
    layer0_outputs(7520) <= (inputs(205)) and not (inputs(134));
    layer0_outputs(7521) <= (inputs(235)) and (inputs(183));
    layer0_outputs(7522) <= not((inputs(169)) or (inputs(69)));
    layer0_outputs(7523) <= (inputs(83)) and not (inputs(194));
    layer0_outputs(7524) <= (inputs(209)) xor (inputs(43));
    layer0_outputs(7525) <= (inputs(231)) and (inputs(180));
    layer0_outputs(7526) <= (inputs(19)) or (inputs(225));
    layer0_outputs(7527) <= (inputs(204)) or (inputs(226));
    layer0_outputs(7528) <= (inputs(136)) and not (inputs(140));
    layer0_outputs(7529) <= not(inputs(207));
    layer0_outputs(7530) <= not((inputs(151)) or (inputs(101)));
    layer0_outputs(7531) <= inputs(198);
    layer0_outputs(7532) <= not((inputs(64)) or (inputs(62)));
    layer0_outputs(7533) <= inputs(169);
    layer0_outputs(7534) <= not(inputs(58));
    layer0_outputs(7535) <= not(inputs(247));
    layer0_outputs(7536) <= (inputs(161)) or (inputs(65));
    layer0_outputs(7537) <= not(inputs(162));
    layer0_outputs(7538) <= not((inputs(75)) or (inputs(77)));
    layer0_outputs(7539) <= (inputs(240)) or (inputs(203));
    layer0_outputs(7540) <= not((inputs(45)) and (inputs(76)));
    layer0_outputs(7541) <= not((inputs(251)) or (inputs(161)));
    layer0_outputs(7542) <= (inputs(47)) xor (inputs(189));
    layer0_outputs(7543) <= inputs(59);
    layer0_outputs(7544) <= (inputs(75)) and (inputs(200));
    layer0_outputs(7545) <= (inputs(34)) or (inputs(234));
    layer0_outputs(7546) <= inputs(146);
    layer0_outputs(7547) <= '1';
    layer0_outputs(7548) <= not(inputs(178));
    layer0_outputs(7549) <= (inputs(148)) or (inputs(95));
    layer0_outputs(7550) <= inputs(53);
    layer0_outputs(7551) <= not((inputs(205)) or (inputs(31)));
    layer0_outputs(7552) <= (inputs(237)) xor (inputs(188));
    layer0_outputs(7553) <= (inputs(231)) and (inputs(83));
    layer0_outputs(7554) <= inputs(113);
    layer0_outputs(7555) <= not((inputs(169)) xor (inputs(177)));
    layer0_outputs(7556) <= inputs(198);
    layer0_outputs(7557) <= not(inputs(54));
    layer0_outputs(7558) <= (inputs(65)) and not (inputs(225));
    layer0_outputs(7559) <= inputs(186);
    layer0_outputs(7560) <= not(inputs(167)) or (inputs(81));
    layer0_outputs(7561) <= (inputs(14)) or (inputs(215));
    layer0_outputs(7562) <= not((inputs(62)) xor (inputs(243)));
    layer0_outputs(7563) <= not(inputs(165)) or (inputs(186));
    layer0_outputs(7564) <= not((inputs(122)) xor (inputs(224)));
    layer0_outputs(7565) <= not(inputs(117)) or (inputs(12));
    layer0_outputs(7566) <= not((inputs(33)) or (inputs(54)));
    layer0_outputs(7567) <= (inputs(74)) and (inputs(211));
    layer0_outputs(7568) <= not(inputs(26));
    layer0_outputs(7569) <= not(inputs(123));
    layer0_outputs(7570) <= (inputs(139)) or (inputs(136));
    layer0_outputs(7571) <= '0';
    layer0_outputs(7572) <= inputs(193);
    layer0_outputs(7573) <= (inputs(132)) and not (inputs(243));
    layer0_outputs(7574) <= (inputs(158)) and not (inputs(30));
    layer0_outputs(7575) <= inputs(38);
    layer0_outputs(7576) <= not((inputs(214)) or (inputs(156)));
    layer0_outputs(7577) <= inputs(180);
    layer0_outputs(7578) <= inputs(76);
    layer0_outputs(7579) <= not(inputs(9));
    layer0_outputs(7580) <= not((inputs(250)) or (inputs(176)));
    layer0_outputs(7581) <= not(inputs(84));
    layer0_outputs(7582) <= not((inputs(67)) or (inputs(181)));
    layer0_outputs(7583) <= inputs(9);
    layer0_outputs(7584) <= not(inputs(173)) or (inputs(31));
    layer0_outputs(7585) <= not((inputs(224)) xor (inputs(194)));
    layer0_outputs(7586) <= (inputs(235)) and not (inputs(19));
    layer0_outputs(7587) <= not((inputs(24)) xor (inputs(53)));
    layer0_outputs(7588) <= (inputs(149)) xor (inputs(238));
    layer0_outputs(7589) <= inputs(165);
    layer0_outputs(7590) <= inputs(144);
    layer0_outputs(7591) <= (inputs(168)) xor (inputs(115));
    layer0_outputs(7592) <= not(inputs(66));
    layer0_outputs(7593) <= inputs(111);
    layer0_outputs(7594) <= (inputs(86)) and not (inputs(150));
    layer0_outputs(7595) <= (inputs(245)) and not (inputs(93));
    layer0_outputs(7596) <= not(inputs(252)) or (inputs(1));
    layer0_outputs(7597) <= not(inputs(8)) or (inputs(162));
    layer0_outputs(7598) <= inputs(244);
    layer0_outputs(7599) <= (inputs(162)) or (inputs(154));
    layer0_outputs(7600) <= '0';
    layer0_outputs(7601) <= not(inputs(97));
    layer0_outputs(7602) <= (inputs(3)) or (inputs(201));
    layer0_outputs(7603) <= not((inputs(254)) or (inputs(248)));
    layer0_outputs(7604) <= not(inputs(137)) or (inputs(111));
    layer0_outputs(7605) <= not(inputs(91));
    layer0_outputs(7606) <= inputs(189);
    layer0_outputs(7607) <= inputs(147);
    layer0_outputs(7608) <= (inputs(38)) and not (inputs(180));
    layer0_outputs(7609) <= (inputs(19)) and not (inputs(239));
    layer0_outputs(7610) <= not(inputs(44)) or (inputs(254));
    layer0_outputs(7611) <= (inputs(252)) and not (inputs(97));
    layer0_outputs(7612) <= (inputs(0)) xor (inputs(60));
    layer0_outputs(7613) <= (inputs(166)) and (inputs(207));
    layer0_outputs(7614) <= '1';
    layer0_outputs(7615) <= (inputs(241)) or (inputs(131));
    layer0_outputs(7616) <= not((inputs(106)) xor (inputs(125)));
    layer0_outputs(7617) <= not(inputs(100));
    layer0_outputs(7618) <= not(inputs(79));
    layer0_outputs(7619) <= not((inputs(16)) and (inputs(95)));
    layer0_outputs(7620) <= not(inputs(146));
    layer0_outputs(7621) <= not(inputs(191)) or (inputs(243));
    layer0_outputs(7622) <= not((inputs(66)) or (inputs(9)));
    layer0_outputs(7623) <= (inputs(230)) and not (inputs(104));
    layer0_outputs(7624) <= not(inputs(57));
    layer0_outputs(7625) <= inputs(121);
    layer0_outputs(7626) <= not((inputs(180)) or (inputs(19)));
    layer0_outputs(7627) <= not(inputs(29)) or (inputs(192));
    layer0_outputs(7628) <= not((inputs(9)) or (inputs(61)));
    layer0_outputs(7629) <= (inputs(178)) or (inputs(205));
    layer0_outputs(7630) <= (inputs(155)) and not (inputs(76));
    layer0_outputs(7631) <= (inputs(232)) and not (inputs(51));
    layer0_outputs(7632) <= inputs(244);
    layer0_outputs(7633) <= (inputs(220)) and not (inputs(211));
    layer0_outputs(7634) <= not((inputs(85)) xor (inputs(100)));
    layer0_outputs(7635) <= not(inputs(40)) or (inputs(236));
    layer0_outputs(7636) <= (inputs(208)) xor (inputs(11));
    layer0_outputs(7637) <= (inputs(176)) or (inputs(224));
    layer0_outputs(7638) <= (inputs(133)) and not (inputs(64));
    layer0_outputs(7639) <= not(inputs(164));
    layer0_outputs(7640) <= (inputs(215)) xor (inputs(185));
    layer0_outputs(7641) <= not(inputs(186));
    layer0_outputs(7642) <= not(inputs(217)) or (inputs(231));
    layer0_outputs(7643) <= not(inputs(194));
    layer0_outputs(7644) <= not(inputs(152)) or (inputs(129));
    layer0_outputs(7645) <= (inputs(200)) or (inputs(69));
    layer0_outputs(7646) <= (inputs(91)) or (inputs(43));
    layer0_outputs(7647) <= (inputs(64)) or (inputs(163));
    layer0_outputs(7648) <= (inputs(237)) xor (inputs(5));
    layer0_outputs(7649) <= inputs(56);
    layer0_outputs(7650) <= not(inputs(102));
    layer0_outputs(7651) <= not(inputs(208)) or (inputs(16));
    layer0_outputs(7652) <= not(inputs(23));
    layer0_outputs(7653) <= not(inputs(82));
    layer0_outputs(7654) <= (inputs(71)) and not (inputs(204));
    layer0_outputs(7655) <= inputs(159);
    layer0_outputs(7656) <= not((inputs(76)) or (inputs(146)));
    layer0_outputs(7657) <= (inputs(202)) or (inputs(52));
    layer0_outputs(7658) <= not(inputs(61));
    layer0_outputs(7659) <= (inputs(98)) and not (inputs(159));
    layer0_outputs(7660) <= (inputs(15)) and not (inputs(78));
    layer0_outputs(7661) <= not((inputs(74)) and (inputs(198)));
    layer0_outputs(7662) <= not(inputs(122));
    layer0_outputs(7663) <= inputs(86);
    layer0_outputs(7664) <= inputs(179);
    layer0_outputs(7665) <= '1';
    layer0_outputs(7666) <= (inputs(177)) or (inputs(85));
    layer0_outputs(7667) <= not(inputs(245));
    layer0_outputs(7668) <= not((inputs(83)) or (inputs(229)));
    layer0_outputs(7669) <= not(inputs(100));
    layer0_outputs(7670) <= not(inputs(204));
    layer0_outputs(7671) <= not(inputs(53));
    layer0_outputs(7672) <= not((inputs(100)) or (inputs(155)));
    layer0_outputs(7673) <= not(inputs(186));
    layer0_outputs(7674) <= not(inputs(150));
    layer0_outputs(7675) <= not(inputs(58)) or (inputs(51));
    layer0_outputs(7676) <= '1';
    layer0_outputs(7677) <= not(inputs(27)) or (inputs(225));
    layer0_outputs(7678) <= not(inputs(115));
    layer0_outputs(7679) <= not(inputs(211)) or (inputs(207));
    outputs(0) <= layer0_outputs(998);
    outputs(1) <= not(layer0_outputs(2266)) or (layer0_outputs(7598));
    outputs(2) <= (layer0_outputs(3511)) or (layer0_outputs(7220));
    outputs(3) <= (layer0_outputs(7360)) xor (layer0_outputs(380));
    outputs(4) <= not((layer0_outputs(649)) and (layer0_outputs(3694)));
    outputs(5) <= not((layer0_outputs(2843)) or (layer0_outputs(6893)));
    outputs(6) <= not(layer0_outputs(1656)) or (layer0_outputs(510));
    outputs(7) <= not(layer0_outputs(4042));
    outputs(8) <= not(layer0_outputs(6739));
    outputs(9) <= not(layer0_outputs(3967)) or (layer0_outputs(3378));
    outputs(10) <= (layer0_outputs(7475)) and not (layer0_outputs(2018));
    outputs(11) <= not(layer0_outputs(1225));
    outputs(12) <= not(layer0_outputs(7165)) or (layer0_outputs(3265));
    outputs(13) <= layer0_outputs(816);
    outputs(14) <= not((layer0_outputs(5518)) or (layer0_outputs(6728)));
    outputs(15) <= (layer0_outputs(6098)) and not (layer0_outputs(1797));
    outputs(16) <= not(layer0_outputs(5540));
    outputs(17) <= not(layer0_outputs(4765));
    outputs(18) <= not(layer0_outputs(741));
    outputs(19) <= layer0_outputs(6134);
    outputs(20) <= layer0_outputs(1894);
    outputs(21) <= (layer0_outputs(4561)) or (layer0_outputs(908));
    outputs(22) <= layer0_outputs(4156);
    outputs(23) <= not((layer0_outputs(3506)) xor (layer0_outputs(3389)));
    outputs(24) <= (layer0_outputs(3484)) and not (layer0_outputs(3383));
    outputs(25) <= not(layer0_outputs(4161)) or (layer0_outputs(4513));
    outputs(26) <= layer0_outputs(5592);
    outputs(27) <= layer0_outputs(2216);
    outputs(28) <= not((layer0_outputs(5641)) and (layer0_outputs(3178)));
    outputs(29) <= (layer0_outputs(3102)) xor (layer0_outputs(3886));
    outputs(30) <= not(layer0_outputs(2059));
    outputs(31) <= (layer0_outputs(3225)) xor (layer0_outputs(2865));
    outputs(32) <= not(layer0_outputs(6481));
    outputs(33) <= not(layer0_outputs(2654));
    outputs(34) <= not(layer0_outputs(1463)) or (layer0_outputs(1608));
    outputs(35) <= (layer0_outputs(6554)) xor (layer0_outputs(3331));
    outputs(36) <= not(layer0_outputs(7678));
    outputs(37) <= layer0_outputs(2150);
    outputs(38) <= (layer0_outputs(4793)) and not (layer0_outputs(2905));
    outputs(39) <= not((layer0_outputs(1007)) or (layer0_outputs(1499)));
    outputs(40) <= not(layer0_outputs(238));
    outputs(41) <= layer0_outputs(4749);
    outputs(42) <= not(layer0_outputs(3820));
    outputs(43) <= not(layer0_outputs(2384));
    outputs(44) <= not(layer0_outputs(2018));
    outputs(45) <= not((layer0_outputs(1499)) and (layer0_outputs(1987)));
    outputs(46) <= layer0_outputs(2692);
    outputs(47) <= layer0_outputs(5696);
    outputs(48) <= (layer0_outputs(4316)) or (layer0_outputs(5010));
    outputs(49) <= not(layer0_outputs(4328));
    outputs(50) <= layer0_outputs(6901);
    outputs(51) <= (layer0_outputs(1589)) xor (layer0_outputs(6992));
    outputs(52) <= not(layer0_outputs(5814)) or (layer0_outputs(3388));
    outputs(53) <= (layer0_outputs(4969)) and (layer0_outputs(5664));
    outputs(54) <= not((layer0_outputs(2860)) or (layer0_outputs(6877)));
    outputs(55) <= (layer0_outputs(2285)) or (layer0_outputs(5866));
    outputs(56) <= not(layer0_outputs(5671)) or (layer0_outputs(3894));
    outputs(57) <= (layer0_outputs(6035)) or (layer0_outputs(7202));
    outputs(58) <= layer0_outputs(6901);
    outputs(59) <= layer0_outputs(6167);
    outputs(60) <= not(layer0_outputs(2299)) or (layer0_outputs(4601));
    outputs(61) <= layer0_outputs(5107);
    outputs(62) <= layer0_outputs(7411);
    outputs(63) <= (layer0_outputs(7125)) and (layer0_outputs(7590));
    outputs(64) <= (layer0_outputs(4077)) and not (layer0_outputs(2523));
    outputs(65) <= not(layer0_outputs(5849));
    outputs(66) <= (layer0_outputs(5106)) or (layer0_outputs(5073));
    outputs(67) <= (layer0_outputs(5490)) and (layer0_outputs(500));
    outputs(68) <= not(layer0_outputs(2520));
    outputs(69) <= not(layer0_outputs(4906));
    outputs(70) <= not(layer0_outputs(6092));
    outputs(71) <= not(layer0_outputs(1150));
    outputs(72) <= not(layer0_outputs(3272));
    outputs(73) <= not(layer0_outputs(3475));
    outputs(74) <= (layer0_outputs(6378)) or (layer0_outputs(5380));
    outputs(75) <= layer0_outputs(6987);
    outputs(76) <= (layer0_outputs(630)) or (layer0_outputs(5292));
    outputs(77) <= not(layer0_outputs(5138));
    outputs(78) <= not(layer0_outputs(2923)) or (layer0_outputs(1982));
    outputs(79) <= not((layer0_outputs(693)) or (layer0_outputs(1578)));
    outputs(80) <= (layer0_outputs(189)) xor (layer0_outputs(3935));
    outputs(81) <= not(layer0_outputs(6429));
    outputs(82) <= not((layer0_outputs(7210)) and (layer0_outputs(2563)));
    outputs(83) <= layer0_outputs(7233);
    outputs(84) <= not((layer0_outputs(3397)) xor (layer0_outputs(6807)));
    outputs(85) <= not((layer0_outputs(4747)) and (layer0_outputs(2499)));
    outputs(86) <= (layer0_outputs(7314)) and (layer0_outputs(6562));
    outputs(87) <= (layer0_outputs(6330)) and (layer0_outputs(1415));
    outputs(88) <= not(layer0_outputs(4856));
    outputs(89) <= not((layer0_outputs(6939)) or (layer0_outputs(2822)));
    outputs(90) <= (layer0_outputs(3551)) and not (layer0_outputs(4549));
    outputs(91) <= not(layer0_outputs(2988));
    outputs(92) <= not(layer0_outputs(4805)) or (layer0_outputs(84));
    outputs(93) <= (layer0_outputs(5938)) and not (layer0_outputs(2621));
    outputs(94) <= not((layer0_outputs(2949)) or (layer0_outputs(6244)));
    outputs(95) <= not(layer0_outputs(6528));
    outputs(96) <= not(layer0_outputs(5466)) or (layer0_outputs(7583));
    outputs(97) <= not(layer0_outputs(1173));
    outputs(98) <= layer0_outputs(4285);
    outputs(99) <= not(layer0_outputs(4609));
    outputs(100) <= layer0_outputs(7577);
    outputs(101) <= not(layer0_outputs(50));
    outputs(102) <= (layer0_outputs(3306)) or (layer0_outputs(5944));
    outputs(103) <= not(layer0_outputs(2396));
    outputs(104) <= (layer0_outputs(514)) and (layer0_outputs(5509));
    outputs(105) <= not((layer0_outputs(858)) xor (layer0_outputs(7141)));
    outputs(106) <= not(layer0_outputs(2545));
    outputs(107) <= not(layer0_outputs(2474));
    outputs(108) <= (layer0_outputs(6529)) and not (layer0_outputs(3586));
    outputs(109) <= not(layer0_outputs(6439));
    outputs(110) <= not(layer0_outputs(4494));
    outputs(111) <= not((layer0_outputs(6126)) xor (layer0_outputs(4596)));
    outputs(112) <= not(layer0_outputs(4095));
    outputs(113) <= not(layer0_outputs(1236)) or (layer0_outputs(3017));
    outputs(114) <= layer0_outputs(772);
    outputs(115) <= not(layer0_outputs(2244));
    outputs(116) <= (layer0_outputs(7026)) xor (layer0_outputs(5478));
    outputs(117) <= layer0_outputs(2583);
    outputs(118) <= layer0_outputs(5941);
    outputs(119) <= layer0_outputs(4786);
    outputs(120) <= layer0_outputs(3658);
    outputs(121) <= not(layer0_outputs(3995));
    outputs(122) <= layer0_outputs(3010);
    outputs(123) <= (layer0_outputs(7321)) xor (layer0_outputs(4923));
    outputs(124) <= not(layer0_outputs(4660));
    outputs(125) <= not(layer0_outputs(9));
    outputs(126) <= not((layer0_outputs(3957)) xor (layer0_outputs(955)));
    outputs(127) <= (layer0_outputs(329)) and not (layer0_outputs(7528));
    outputs(128) <= not((layer0_outputs(3965)) or (layer0_outputs(5038)));
    outputs(129) <= not((layer0_outputs(6216)) and (layer0_outputs(2498)));
    outputs(130) <= not(layer0_outputs(5127));
    outputs(131) <= not(layer0_outputs(2109)) or (layer0_outputs(3395));
    outputs(132) <= (layer0_outputs(6237)) and (layer0_outputs(6665));
    outputs(133) <= not((layer0_outputs(1210)) or (layer0_outputs(3123)));
    outputs(134) <= not(layer0_outputs(2461)) or (layer0_outputs(7574));
    outputs(135) <= layer0_outputs(2040);
    outputs(136) <= not((layer0_outputs(4570)) or (layer0_outputs(5135)));
    outputs(137) <= (layer0_outputs(7086)) and (layer0_outputs(7312));
    outputs(138) <= layer0_outputs(887);
    outputs(139) <= not(layer0_outputs(3170));
    outputs(140) <= not(layer0_outputs(3808));
    outputs(141) <= (layer0_outputs(1439)) or (layer0_outputs(5792));
    outputs(142) <= layer0_outputs(319);
    outputs(143) <= (layer0_outputs(475)) and not (layer0_outputs(3291));
    outputs(144) <= (layer0_outputs(6693)) xor (layer0_outputs(3536));
    outputs(145) <= not(layer0_outputs(5272)) or (layer0_outputs(707));
    outputs(146) <= not((layer0_outputs(7385)) or (layer0_outputs(3608)));
    outputs(147) <= not((layer0_outputs(1521)) or (layer0_outputs(6962)));
    outputs(148) <= not(layer0_outputs(5741));
    outputs(149) <= layer0_outputs(6394);
    outputs(150) <= layer0_outputs(5002);
    outputs(151) <= layer0_outputs(5155);
    outputs(152) <= not(layer0_outputs(5806));
    outputs(153) <= (layer0_outputs(5927)) or (layer0_outputs(5976));
    outputs(154) <= not(layer0_outputs(4733));
    outputs(155) <= layer0_outputs(1443);
    outputs(156) <= (layer0_outputs(7320)) or (layer0_outputs(7623));
    outputs(157) <= not(layer0_outputs(5825));
    outputs(158) <= not((layer0_outputs(5656)) and (layer0_outputs(3214)));
    outputs(159) <= not(layer0_outputs(1259));
    outputs(160) <= not(layer0_outputs(5680));
    outputs(161) <= layer0_outputs(1432);
    outputs(162) <= not(layer0_outputs(2743));
    outputs(163) <= not(layer0_outputs(4939));
    outputs(164) <= not(layer0_outputs(6270));
    outputs(165) <= layer0_outputs(5569);
    outputs(166) <= not((layer0_outputs(3774)) and (layer0_outputs(3642)));
    outputs(167) <= (layer0_outputs(6243)) and not (layer0_outputs(3288));
    outputs(168) <= (layer0_outputs(7304)) xor (layer0_outputs(7442));
    outputs(169) <= not(layer0_outputs(64));
    outputs(170) <= layer0_outputs(4888);
    outputs(171) <= (layer0_outputs(627)) and (layer0_outputs(799));
    outputs(172) <= not(layer0_outputs(48));
    outputs(173) <= layer0_outputs(60);
    outputs(174) <= not(layer0_outputs(4792));
    outputs(175) <= (layer0_outputs(436)) and not (layer0_outputs(637));
    outputs(176) <= not((layer0_outputs(5970)) or (layer0_outputs(4201)));
    outputs(177) <= not(layer0_outputs(206));
    outputs(178) <= layer0_outputs(3676);
    outputs(179) <= (layer0_outputs(6960)) and not (layer0_outputs(4621));
    outputs(180) <= not(layer0_outputs(2769));
    outputs(181) <= layer0_outputs(3365);
    outputs(182) <= (layer0_outputs(5513)) and not (layer0_outputs(358));
    outputs(183) <= not(layer0_outputs(4765));
    outputs(184) <= not((layer0_outputs(470)) and (layer0_outputs(1173)));
    outputs(185) <= (layer0_outputs(5171)) xor (layer0_outputs(4138));
    outputs(186) <= not((layer0_outputs(5370)) or (layer0_outputs(7159)));
    outputs(187) <= not(layer0_outputs(4069));
    outputs(188) <= not(layer0_outputs(7228));
    outputs(189) <= layer0_outputs(7126);
    outputs(190) <= not(layer0_outputs(2723));
    outputs(191) <= layer0_outputs(3643);
    outputs(192) <= not(layer0_outputs(5480));
    outputs(193) <= not(layer0_outputs(4836));
    outputs(194) <= layer0_outputs(2204);
    outputs(195) <= not((layer0_outputs(6208)) and (layer0_outputs(211)));
    outputs(196) <= not(layer0_outputs(3356));
    outputs(197) <= (layer0_outputs(6813)) and not (layer0_outputs(2835));
    outputs(198) <= layer0_outputs(2186);
    outputs(199) <= not(layer0_outputs(5478));
    outputs(200) <= not((layer0_outputs(4037)) or (layer0_outputs(2543)));
    outputs(201) <= (layer0_outputs(7291)) and not (layer0_outputs(6793));
    outputs(202) <= not(layer0_outputs(7242));
    outputs(203) <= not(layer0_outputs(4858)) or (layer0_outputs(4208));
    outputs(204) <= not(layer0_outputs(1667));
    outputs(205) <= not(layer0_outputs(4705));
    outputs(206) <= layer0_outputs(2475);
    outputs(207) <= (layer0_outputs(6913)) and not (layer0_outputs(5870));
    outputs(208) <= (layer0_outputs(54)) and not (layer0_outputs(808));
    outputs(209) <= (layer0_outputs(2132)) xor (layer0_outputs(2256));
    outputs(210) <= layer0_outputs(1839);
    outputs(211) <= layer0_outputs(1349);
    outputs(212) <= not(layer0_outputs(7224));
    outputs(213) <= layer0_outputs(7435);
    outputs(214) <= not(layer0_outputs(3115));
    outputs(215) <= (layer0_outputs(4141)) and not (layer0_outputs(1081));
    outputs(216) <= not(layer0_outputs(1095));
    outputs(217) <= not(layer0_outputs(675)) or (layer0_outputs(2184));
    outputs(218) <= layer0_outputs(5491);
    outputs(219) <= (layer0_outputs(5270)) and not (layer0_outputs(7029));
    outputs(220) <= layer0_outputs(6011);
    outputs(221) <= (layer0_outputs(1618)) or (layer0_outputs(7642));
    outputs(222) <= (layer0_outputs(4066)) and (layer0_outputs(399));
    outputs(223) <= layer0_outputs(2539);
    outputs(224) <= (layer0_outputs(5035)) xor (layer0_outputs(2083));
    outputs(225) <= layer0_outputs(4691);
    outputs(226) <= not(layer0_outputs(2638));
    outputs(227) <= not(layer0_outputs(242));
    outputs(228) <= not((layer0_outputs(5206)) xor (layer0_outputs(1611)));
    outputs(229) <= not(layer0_outputs(2316));
    outputs(230) <= layer0_outputs(4211);
    outputs(231) <= not((layer0_outputs(2981)) xor (layer0_outputs(6647)));
    outputs(232) <= not(layer0_outputs(4313));
    outputs(233) <= layer0_outputs(1240);
    outputs(234) <= not(layer0_outputs(4228));
    outputs(235) <= layer0_outputs(5129);
    outputs(236) <= not((layer0_outputs(1663)) xor (layer0_outputs(3922)));
    outputs(237) <= not(layer0_outputs(4664));
    outputs(238) <= (layer0_outputs(1884)) and not (layer0_outputs(1141));
    outputs(239) <= not((layer0_outputs(682)) xor (layer0_outputs(7306)));
    outputs(240) <= layer0_outputs(2757);
    outputs(241) <= layer0_outputs(2287);
    outputs(242) <= not((layer0_outputs(4639)) and (layer0_outputs(2485)));
    outputs(243) <= (layer0_outputs(4241)) and not (layer0_outputs(4800));
    outputs(244) <= not((layer0_outputs(2032)) or (layer0_outputs(1796)));
    outputs(245) <= not(layer0_outputs(3962)) or (layer0_outputs(4920));
    outputs(246) <= (layer0_outputs(6074)) xor (layer0_outputs(7182));
    outputs(247) <= not((layer0_outputs(3877)) or (layer0_outputs(7109)));
    outputs(248) <= not((layer0_outputs(7538)) or (layer0_outputs(4454)));
    outputs(249) <= layer0_outputs(2371);
    outputs(250) <= not((layer0_outputs(1152)) and (layer0_outputs(3127)));
    outputs(251) <= layer0_outputs(5491);
    outputs(252) <= layer0_outputs(430);
    outputs(253) <= not(layer0_outputs(7148));
    outputs(254) <= not(layer0_outputs(2110)) or (layer0_outputs(7142));
    outputs(255) <= (layer0_outputs(6076)) and not (layer0_outputs(1815));
    outputs(256) <= not(layer0_outputs(2567)) or (layer0_outputs(5619));
    outputs(257) <= layer0_outputs(4416);
    outputs(258) <= (layer0_outputs(4487)) or (layer0_outputs(1833));
    outputs(259) <= not(layer0_outputs(201));
    outputs(260) <= not(layer0_outputs(259));
    outputs(261) <= not(layer0_outputs(5801));
    outputs(262) <= not(layer0_outputs(4248)) or (layer0_outputs(6298));
    outputs(263) <= (layer0_outputs(5120)) or (layer0_outputs(2042));
    outputs(264) <= not(layer0_outputs(5661));
    outputs(265) <= not(layer0_outputs(4125)) or (layer0_outputs(389));
    outputs(266) <= layer0_outputs(4194);
    outputs(267) <= not((layer0_outputs(5414)) and (layer0_outputs(4737)));
    outputs(268) <= not((layer0_outputs(3508)) xor (layer0_outputs(5933)));
    outputs(269) <= layer0_outputs(1069);
    outputs(270) <= not(layer0_outputs(3259));
    outputs(271) <= not(layer0_outputs(2743));
    outputs(272) <= not(layer0_outputs(5743));
    outputs(273) <= (layer0_outputs(765)) and not (layer0_outputs(817));
    outputs(274) <= not(layer0_outputs(72));
    outputs(275) <= not((layer0_outputs(572)) or (layer0_outputs(6896)));
    outputs(276) <= (layer0_outputs(7336)) and not (layer0_outputs(1390));
    outputs(277) <= layer0_outputs(317);
    outputs(278) <= not((layer0_outputs(2452)) and (layer0_outputs(790)));
    outputs(279) <= not((layer0_outputs(6117)) and (layer0_outputs(2735)));
    outputs(280) <= not(layer0_outputs(1800));
    outputs(281) <= not(layer0_outputs(5156));
    outputs(282) <= not((layer0_outputs(886)) and (layer0_outputs(1340)));
    outputs(283) <= not((layer0_outputs(5565)) xor (layer0_outputs(7319)));
    outputs(284) <= not((layer0_outputs(4581)) and (layer0_outputs(3520)));
    outputs(285) <= layer0_outputs(4039);
    outputs(286) <= layer0_outputs(1248);
    outputs(287) <= layer0_outputs(2507);
    outputs(288) <= (layer0_outputs(6218)) and not (layer0_outputs(3584));
    outputs(289) <= not(layer0_outputs(6883)) or (layer0_outputs(1620));
    outputs(290) <= not(layer0_outputs(719));
    outputs(291) <= not(layer0_outputs(6970));
    outputs(292) <= layer0_outputs(3951);
    outputs(293) <= not((layer0_outputs(4817)) or (layer0_outputs(3878)));
    outputs(294) <= not(layer0_outputs(7031)) or (layer0_outputs(6114));
    outputs(295) <= not(layer0_outputs(5897));
    outputs(296) <= (layer0_outputs(380)) xor (layer0_outputs(793));
    outputs(297) <= not((layer0_outputs(2624)) and (layer0_outputs(2223)));
    outputs(298) <= (layer0_outputs(2123)) and not (layer0_outputs(4794));
    outputs(299) <= not(layer0_outputs(2854));
    outputs(300) <= not((layer0_outputs(6283)) xor (layer0_outputs(1114)));
    outputs(301) <= not((layer0_outputs(4192)) and (layer0_outputs(5386)));
    outputs(302) <= layer0_outputs(6673);
    outputs(303) <= layer0_outputs(7664);
    outputs(304) <= not(layer0_outputs(5939));
    outputs(305) <= not(layer0_outputs(4564));
    outputs(306) <= layer0_outputs(257);
    outputs(307) <= layer0_outputs(6743);
    outputs(308) <= layer0_outputs(836);
    outputs(309) <= layer0_outputs(7194);
    outputs(310) <= layer0_outputs(729);
    outputs(311) <= layer0_outputs(2670);
    outputs(312) <= not((layer0_outputs(361)) xor (layer0_outputs(7265)));
    outputs(313) <= not((layer0_outputs(5980)) or (layer0_outputs(791)));
    outputs(314) <= layer0_outputs(2781);
    outputs(315) <= not(layer0_outputs(3058));
    outputs(316) <= not((layer0_outputs(6999)) and (layer0_outputs(7111)));
    outputs(317) <= (layer0_outputs(3232)) and (layer0_outputs(5027));
    outputs(318) <= layer0_outputs(1286);
    outputs(319) <= layer0_outputs(4221);
    outputs(320) <= not((layer0_outputs(1345)) xor (layer0_outputs(3766)));
    outputs(321) <= (layer0_outputs(5246)) xor (layer0_outputs(6497));
    outputs(322) <= (layer0_outputs(1012)) or (layer0_outputs(4163));
    outputs(323) <= layer0_outputs(1435);
    outputs(324) <= layer0_outputs(6801);
    outputs(325) <= (layer0_outputs(686)) or (layer0_outputs(2457));
    outputs(326) <= not(layer0_outputs(709));
    outputs(327) <= layer0_outputs(3506);
    outputs(328) <= not(layer0_outputs(5232));
    outputs(329) <= not((layer0_outputs(5003)) or (layer0_outputs(770)));
    outputs(330) <= not((layer0_outputs(5647)) xor (layer0_outputs(1455)));
    outputs(331) <= not((layer0_outputs(7176)) and (layer0_outputs(4874)));
    outputs(332) <= not(layer0_outputs(5289)) or (layer0_outputs(5333));
    outputs(333) <= (layer0_outputs(527)) or (layer0_outputs(917));
    outputs(334) <= layer0_outputs(3763);
    outputs(335) <= (layer0_outputs(6231)) xor (layer0_outputs(7008));
    outputs(336) <= not((layer0_outputs(2819)) xor (layer0_outputs(7102)));
    outputs(337) <= (layer0_outputs(1378)) and not (layer0_outputs(3459));
    outputs(338) <= layer0_outputs(3936);
    outputs(339) <= layer0_outputs(6679);
    outputs(340) <= layer0_outputs(1423);
    outputs(341) <= layer0_outputs(4908);
    outputs(342) <= (layer0_outputs(4081)) xor (layer0_outputs(1645));
    outputs(343) <= (layer0_outputs(5233)) or (layer0_outputs(2016));
    outputs(344) <= layer0_outputs(4052);
    outputs(345) <= layer0_outputs(4640);
    outputs(346) <= (layer0_outputs(6771)) and (layer0_outputs(2759));
    outputs(347) <= not(layer0_outputs(7353));
    outputs(348) <= not((layer0_outputs(745)) and (layer0_outputs(4876)));
    outputs(349) <= not((layer0_outputs(531)) xor (layer0_outputs(6249)));
    outputs(350) <= (layer0_outputs(764)) and not (layer0_outputs(4775));
    outputs(351) <= (layer0_outputs(1544)) or (layer0_outputs(5742));
    outputs(352) <= not(layer0_outputs(5185));
    outputs(353) <= (layer0_outputs(6595)) or (layer0_outputs(4640));
    outputs(354) <= not(layer0_outputs(207));
    outputs(355) <= not(layer0_outputs(3772));
    outputs(356) <= layer0_outputs(5572);
    outputs(357) <= not((layer0_outputs(2802)) or (layer0_outputs(5043)));
    outputs(358) <= not((layer0_outputs(7079)) or (layer0_outputs(3416)));
    outputs(359) <= not(layer0_outputs(5109)) or (layer0_outputs(7278));
    outputs(360) <= layer0_outputs(43);
    outputs(361) <= not(layer0_outputs(2902));
    outputs(362) <= (layer0_outputs(6158)) and not (layer0_outputs(2893));
    outputs(363) <= layer0_outputs(5300);
    outputs(364) <= not(layer0_outputs(2861));
    outputs(365) <= not(layer0_outputs(6724));
    outputs(366) <= not((layer0_outputs(1758)) and (layer0_outputs(5205)));
    outputs(367) <= (layer0_outputs(7436)) and not (layer0_outputs(3032));
    outputs(368) <= (layer0_outputs(5878)) and (layer0_outputs(7076));
    outputs(369) <= (layer0_outputs(5177)) and (layer0_outputs(1558));
    outputs(370) <= layer0_outputs(7028);
    outputs(371) <= not((layer0_outputs(7150)) xor (layer0_outputs(4807)));
    outputs(372) <= layer0_outputs(3394);
    outputs(373) <= not(layer0_outputs(2859));
    outputs(374) <= not(layer0_outputs(5570)) or (layer0_outputs(2354));
    outputs(375) <= layer0_outputs(1869);
    outputs(376) <= (layer0_outputs(6129)) and not (layer0_outputs(2326));
    outputs(377) <= (layer0_outputs(4969)) and not (layer0_outputs(3104));
    outputs(378) <= not(layer0_outputs(7396)) or (layer0_outputs(5172));
    outputs(379) <= layer0_outputs(7654);
    outputs(380) <= layer0_outputs(6287);
    outputs(381) <= layer0_outputs(3119);
    outputs(382) <= (layer0_outputs(6952)) and not (layer0_outputs(773));
    outputs(383) <= (layer0_outputs(6484)) xor (layer0_outputs(7471));
    outputs(384) <= (layer0_outputs(290)) and (layer0_outputs(5117));
    outputs(385) <= (layer0_outputs(3541)) and not (layer0_outputs(2695));
    outputs(386) <= layer0_outputs(1418);
    outputs(387) <= not(layer0_outputs(2591));
    outputs(388) <= (layer0_outputs(2412)) xor (layer0_outputs(6703));
    outputs(389) <= (layer0_outputs(4500)) xor (layer0_outputs(3240));
    outputs(390) <= layer0_outputs(3514);
    outputs(391) <= not((layer0_outputs(487)) xor (layer0_outputs(3420)));
    outputs(392) <= not(layer0_outputs(3085));
    outputs(393) <= (layer0_outputs(5442)) and not (layer0_outputs(473));
    outputs(394) <= not(layer0_outputs(5781));
    outputs(395) <= (layer0_outputs(7514)) and not (layer0_outputs(3038));
    outputs(396) <= not(layer0_outputs(2775)) or (layer0_outputs(5824));
    outputs(397) <= layer0_outputs(5650);
    outputs(398) <= not(layer0_outputs(519)) or (layer0_outputs(1992));
    outputs(399) <= not(layer0_outputs(2671));
    outputs(400) <= not(layer0_outputs(3059)) or (layer0_outputs(1774));
    outputs(401) <= layer0_outputs(4307);
    outputs(402) <= layer0_outputs(5774);
    outputs(403) <= not((layer0_outputs(6860)) xor (layer0_outputs(7303)));
    outputs(404) <= not(layer0_outputs(1716)) or (layer0_outputs(1685));
    outputs(405) <= not(layer0_outputs(859));
    outputs(406) <= layer0_outputs(2398);
    outputs(407) <= layer0_outputs(306);
    outputs(408) <= not((layer0_outputs(3135)) or (layer0_outputs(3031)));
    outputs(409) <= not(layer0_outputs(5059));
    outputs(410) <= layer0_outputs(6349);
    outputs(411) <= not(layer0_outputs(3351));
    outputs(412) <= (layer0_outputs(4880)) and not (layer0_outputs(4429));
    outputs(413) <= layer0_outputs(6239);
    outputs(414) <= not(layer0_outputs(840)) or (layer0_outputs(5698));
    outputs(415) <= layer0_outputs(3514);
    outputs(416) <= not(layer0_outputs(6042));
    outputs(417) <= not(layer0_outputs(7648));
    outputs(418) <= layer0_outputs(480);
    outputs(419) <= not(layer0_outputs(975));
    outputs(420) <= layer0_outputs(1087);
    outputs(421) <= (layer0_outputs(3074)) or (layer0_outputs(2303));
    outputs(422) <= (layer0_outputs(1714)) xor (layer0_outputs(4119));
    outputs(423) <= (layer0_outputs(1877)) and (layer0_outputs(1707));
    outputs(424) <= not(layer0_outputs(2356));
    outputs(425) <= not((layer0_outputs(7191)) or (layer0_outputs(2409)));
    outputs(426) <= (layer0_outputs(4445)) or (layer0_outputs(6774));
    outputs(427) <= not(layer0_outputs(906));
    outputs(428) <= (layer0_outputs(2021)) or (layer0_outputs(4243));
    outputs(429) <= layer0_outputs(5328);
    outputs(430) <= (layer0_outputs(136)) and (layer0_outputs(2290));
    outputs(431) <= not(layer0_outputs(7234));
    outputs(432) <= not((layer0_outputs(3369)) and (layer0_outputs(3142)));
    outputs(433) <= layer0_outputs(1794);
    outputs(434) <= layer0_outputs(117);
    outputs(435) <= layer0_outputs(7315);
    outputs(436) <= not((layer0_outputs(3159)) xor (layer0_outputs(5052)));
    outputs(437) <= (layer0_outputs(5338)) or (layer0_outputs(1005));
    outputs(438) <= not(layer0_outputs(6154));
    outputs(439) <= not(layer0_outputs(4507));
    outputs(440) <= not((layer0_outputs(4084)) xor (layer0_outputs(6712)));
    outputs(441) <= layer0_outputs(4456);
    outputs(442) <= not((layer0_outputs(573)) xor (layer0_outputs(3682)));
    outputs(443) <= layer0_outputs(6794);
    outputs(444) <= (layer0_outputs(5423)) and not (layer0_outputs(3029));
    outputs(445) <= not((layer0_outputs(1952)) xor (layer0_outputs(1554)));
    outputs(446) <= (layer0_outputs(1850)) or (layer0_outputs(548));
    outputs(447) <= not((layer0_outputs(35)) and (layer0_outputs(3000)));
    outputs(448) <= (layer0_outputs(213)) or (layer0_outputs(4615));
    outputs(449) <= (layer0_outputs(1406)) or (layer0_outputs(7655));
    outputs(450) <= not(layer0_outputs(553));
    outputs(451) <= (layer0_outputs(5124)) and not (layer0_outputs(2518));
    outputs(452) <= (layer0_outputs(2557)) and not (layer0_outputs(6932));
    outputs(453) <= not(layer0_outputs(1751));
    outputs(454) <= (layer0_outputs(4394)) and (layer0_outputs(3181));
    outputs(455) <= not(layer0_outputs(4010)) or (layer0_outputs(687));
    outputs(456) <= not(layer0_outputs(7114)) or (layer0_outputs(2890));
    outputs(457) <= layer0_outputs(478);
    outputs(458) <= not(layer0_outputs(698));
    outputs(459) <= not(layer0_outputs(6470)) or (layer0_outputs(4407));
    outputs(460) <= (layer0_outputs(2417)) and (layer0_outputs(1991));
    outputs(461) <= not(layer0_outputs(1727));
    outputs(462) <= layer0_outputs(1331);
    outputs(463) <= not(layer0_outputs(198)) or (layer0_outputs(3525));
    outputs(464) <= not((layer0_outputs(3320)) and (layer0_outputs(1836)));
    outputs(465) <= (layer0_outputs(3872)) xor (layer0_outputs(3479));
    outputs(466) <= layer0_outputs(3991);
    outputs(467) <= not(layer0_outputs(6684));
    outputs(468) <= not(layer0_outputs(5207));
    outputs(469) <= not(layer0_outputs(4034)) or (layer0_outputs(7297));
    outputs(470) <= layer0_outputs(7089);
    outputs(471) <= layer0_outputs(3392);
    outputs(472) <= layer0_outputs(6606);
    outputs(473) <= not((layer0_outputs(582)) or (layer0_outputs(5018)));
    outputs(474) <= not(layer0_outputs(5422));
    outputs(475) <= (layer0_outputs(5527)) and (layer0_outputs(1573));
    outputs(476) <= not((layer0_outputs(2231)) or (layer0_outputs(5874)));
    outputs(477) <= not(layer0_outputs(1197));
    outputs(478) <= not(layer0_outputs(1528));
    outputs(479) <= not((layer0_outputs(3137)) or (layer0_outputs(5363)));
    outputs(480) <= not(layer0_outputs(96)) or (layer0_outputs(1337));
    outputs(481) <= layer0_outputs(4092);
    outputs(482) <= not(layer0_outputs(3066));
    outputs(483) <= not(layer0_outputs(6902));
    outputs(484) <= not(layer0_outputs(593));
    outputs(485) <= layer0_outputs(2972);
    outputs(486) <= layer0_outputs(5233);
    outputs(487) <= not((layer0_outputs(70)) or (layer0_outputs(4789)));
    outputs(488) <= layer0_outputs(4241);
    outputs(489) <= not(layer0_outputs(2502));
    outputs(490) <= (layer0_outputs(7467)) or (layer0_outputs(7016));
    outputs(491) <= not(layer0_outputs(7512));
    outputs(492) <= not(layer0_outputs(2224)) or (layer0_outputs(5427));
    outputs(493) <= not(layer0_outputs(3178)) or (layer0_outputs(5004));
    outputs(494) <= not(layer0_outputs(1128)) or (layer0_outputs(1591));
    outputs(495) <= (layer0_outputs(4379)) and not (layer0_outputs(971));
    outputs(496) <= (layer0_outputs(2626)) and not (layer0_outputs(7148));
    outputs(497) <= (layer0_outputs(414)) or (layer0_outputs(5544));
    outputs(498) <= not(layer0_outputs(3350));
    outputs(499) <= (layer0_outputs(6077)) and not (layer0_outputs(6781));
    outputs(500) <= layer0_outputs(6091);
    outputs(501) <= not(layer0_outputs(2084));
    outputs(502) <= layer0_outputs(3517);
    outputs(503) <= not(layer0_outputs(1086)) or (layer0_outputs(1315));
    outputs(504) <= (layer0_outputs(6192)) or (layer0_outputs(1122));
    outputs(505) <= layer0_outputs(4546);
    outputs(506) <= not(layer0_outputs(3917));
    outputs(507) <= not(layer0_outputs(1932));
    outputs(508) <= not((layer0_outputs(166)) and (layer0_outputs(3212)));
    outputs(509) <= (layer0_outputs(2781)) and not (layer0_outputs(2593));
    outputs(510) <= not((layer0_outputs(6336)) and (layer0_outputs(1266)));
    outputs(511) <= layer0_outputs(5595);
    outputs(512) <= not(layer0_outputs(6964));
    outputs(513) <= not(layer0_outputs(1687)) or (layer0_outputs(1309));
    outputs(514) <= (layer0_outputs(1084)) and not (layer0_outputs(1438));
    outputs(515) <= layer0_outputs(1595);
    outputs(516) <= not(layer0_outputs(5949));
    outputs(517) <= not(layer0_outputs(6829));
    outputs(518) <= (layer0_outputs(7562)) or (layer0_outputs(2142));
    outputs(519) <= not((layer0_outputs(7636)) xor (layer0_outputs(5733)));
    outputs(520) <= (layer0_outputs(7468)) or (layer0_outputs(1616));
    outputs(521) <= layer0_outputs(3500);
    outputs(522) <= not(layer0_outputs(390));
    outputs(523) <= not((layer0_outputs(4972)) xor (layer0_outputs(3345)));
    outputs(524) <= not(layer0_outputs(3807));
    outputs(525) <= layer0_outputs(5377);
    outputs(526) <= not(layer0_outputs(6773));
    outputs(527) <= not(layer0_outputs(5680)) or (layer0_outputs(7411));
    outputs(528) <= layer0_outputs(2696);
    outputs(529) <= (layer0_outputs(1537)) and not (layer0_outputs(428));
    outputs(530) <= layer0_outputs(7162);
    outputs(531) <= not(layer0_outputs(1886));
    outputs(532) <= not(layer0_outputs(7096));
    outputs(533) <= not(layer0_outputs(681));
    outputs(534) <= layer0_outputs(1010);
    outputs(535) <= not(layer0_outputs(1183));
    outputs(536) <= not(layer0_outputs(868));
    outputs(537) <= not(layer0_outputs(3277));
    outputs(538) <= layer0_outputs(77);
    outputs(539) <= not(layer0_outputs(2361));
    outputs(540) <= layer0_outputs(7422);
    outputs(541) <= layer0_outputs(6532);
    outputs(542) <= not(layer0_outputs(655));
    outputs(543) <= not((layer0_outputs(5607)) xor (layer0_outputs(2223)));
    outputs(544) <= not(layer0_outputs(4155));
    outputs(545) <= not((layer0_outputs(6739)) or (layer0_outputs(3615)));
    outputs(546) <= not(layer0_outputs(3998));
    outputs(547) <= (layer0_outputs(991)) and (layer0_outputs(4712));
    outputs(548) <= (layer0_outputs(4227)) xor (layer0_outputs(4096));
    outputs(549) <= layer0_outputs(1280);
    outputs(550) <= not(layer0_outputs(4951));
    outputs(551) <= not(layer0_outputs(6073));
    outputs(552) <= layer0_outputs(976);
    outputs(553) <= layer0_outputs(914);
    outputs(554) <= not(layer0_outputs(5741));
    outputs(555) <= not((layer0_outputs(3458)) or (layer0_outputs(2037)));
    outputs(556) <= (layer0_outputs(276)) and not (layer0_outputs(4334));
    outputs(557) <= layer0_outputs(2592);
    outputs(558) <= layer0_outputs(2801);
    outputs(559) <= not((layer0_outputs(1180)) or (layer0_outputs(1938)));
    outputs(560) <= not(layer0_outputs(1197));
    outputs(561) <= (layer0_outputs(3505)) and not (layer0_outputs(3703));
    outputs(562) <= (layer0_outputs(5645)) and not (layer0_outputs(1680));
    outputs(563) <= (layer0_outputs(3606)) and (layer0_outputs(1186));
    outputs(564) <= (layer0_outputs(1855)) and not (layer0_outputs(2889));
    outputs(565) <= not(layer0_outputs(5923));
    outputs(566) <= layer0_outputs(6221);
    outputs(567) <= not(layer0_outputs(5322));
    outputs(568) <= (layer0_outputs(5395)) and not (layer0_outputs(3210));
    outputs(569) <= not(layer0_outputs(2993));
    outputs(570) <= not(layer0_outputs(5194));
    outputs(571) <= not(layer0_outputs(3113));
    outputs(572) <= not(layer0_outputs(2722));
    outputs(573) <= not(layer0_outputs(2538));
    outputs(574) <= (layer0_outputs(6013)) and not (layer0_outputs(2913));
    outputs(575) <= layer0_outputs(1719);
    outputs(576) <= not(layer0_outputs(2331));
    outputs(577) <= not((layer0_outputs(1521)) or (layer0_outputs(4795)));
    outputs(578) <= (layer0_outputs(1522)) and not (layer0_outputs(1180));
    outputs(579) <= (layer0_outputs(1147)) or (layer0_outputs(4948));
    outputs(580) <= not((layer0_outputs(342)) and (layer0_outputs(4300)));
    outputs(581) <= not((layer0_outputs(6382)) and (layer0_outputs(2817)));
    outputs(582) <= layer0_outputs(1709);
    outputs(583) <= (layer0_outputs(1860)) and (layer0_outputs(6765));
    outputs(584) <= (layer0_outputs(805)) xor (layer0_outputs(1572));
    outputs(585) <= layer0_outputs(6339);
    outputs(586) <= layer0_outputs(4436);
    outputs(587) <= layer0_outputs(167);
    outputs(588) <= layer0_outputs(25);
    outputs(589) <= (layer0_outputs(844)) and not (layer0_outputs(7391));
    outputs(590) <= layer0_outputs(7543);
    outputs(591) <= not((layer0_outputs(4772)) xor (layer0_outputs(6281)));
    outputs(592) <= not(layer0_outputs(534)) or (layer0_outputs(1973));
    outputs(593) <= not(layer0_outputs(6176)) or (layer0_outputs(6977));
    outputs(594) <= not((layer0_outputs(4740)) xor (layer0_outputs(1920)));
    outputs(595) <= layer0_outputs(4066);
    outputs(596) <= not((layer0_outputs(6979)) xor (layer0_outputs(1198)));
    outputs(597) <= not(layer0_outputs(2192)) or (layer0_outputs(2016));
    outputs(598) <= (layer0_outputs(3870)) xor (layer0_outputs(2005));
    outputs(599) <= (layer0_outputs(5390)) xor (layer0_outputs(1014));
    outputs(600) <= not(layer0_outputs(7051));
    outputs(601) <= layer0_outputs(5587);
    outputs(602) <= not((layer0_outputs(3531)) or (layer0_outputs(4463)));
    outputs(603) <= not((layer0_outputs(5112)) or (layer0_outputs(554)));
    outputs(604) <= (layer0_outputs(1964)) or (layer0_outputs(980));
    outputs(605) <= layer0_outputs(4852);
    outputs(606) <= not(layer0_outputs(3111));
    outputs(607) <= (layer0_outputs(1646)) or (layer0_outputs(2145));
    outputs(608) <= not(layer0_outputs(5086));
    outputs(609) <= not(layer0_outputs(3113));
    outputs(610) <= not((layer0_outputs(1682)) and (layer0_outputs(3803)));
    outputs(611) <= not((layer0_outputs(1817)) xor (layer0_outputs(6087)));
    outputs(612) <= (layer0_outputs(357)) and (layer0_outputs(247));
    outputs(613) <= not(layer0_outputs(6402)) or (layer0_outputs(2393));
    outputs(614) <= not(layer0_outputs(4783));
    outputs(615) <= not(layer0_outputs(2595));
    outputs(616) <= (layer0_outputs(3067)) and (layer0_outputs(5243));
    outputs(617) <= not((layer0_outputs(1918)) xor (layer0_outputs(5830)));
    outputs(618) <= (layer0_outputs(5104)) or (layer0_outputs(7549));
    outputs(619) <= layer0_outputs(6907);
    outputs(620) <= not((layer0_outputs(3868)) or (layer0_outputs(977)));
    outputs(621) <= (layer0_outputs(2181)) and (layer0_outputs(5101));
    outputs(622) <= (layer0_outputs(4341)) and not (layer0_outputs(204));
    outputs(623) <= (layer0_outputs(4882)) xor (layer0_outputs(4344));
    outputs(624) <= not((layer0_outputs(6645)) and (layer0_outputs(732)));
    outputs(625) <= layer0_outputs(5499);
    outputs(626) <= layer0_outputs(6143);
    outputs(627) <= not(layer0_outputs(733)) or (layer0_outputs(1155));
    outputs(628) <= not((layer0_outputs(1691)) and (layer0_outputs(4108)));
    outputs(629) <= not(layer0_outputs(2103));
    outputs(630) <= not(layer0_outputs(3426));
    outputs(631) <= not(layer0_outputs(1256)) or (layer0_outputs(6695));
    outputs(632) <= not((layer0_outputs(7015)) or (layer0_outputs(7113)));
    outputs(633) <= not(layer0_outputs(4527)) or (layer0_outputs(747));
    outputs(634) <= not((layer0_outputs(5924)) or (layer0_outputs(313)));
    outputs(635) <= (layer0_outputs(6454)) or (layer0_outputs(5564));
    outputs(636) <= not(layer0_outputs(2724)) or (layer0_outputs(270));
    outputs(637) <= not(layer0_outputs(283));
    outputs(638) <= (layer0_outputs(95)) xor (layer0_outputs(5376));
    outputs(639) <= not((layer0_outputs(4290)) xor (layer0_outputs(3857)));
    outputs(640) <= not(layer0_outputs(2397));
    outputs(641) <= not(layer0_outputs(1232));
    outputs(642) <= not(layer0_outputs(5785)) or (layer0_outputs(1633));
    outputs(643) <= layer0_outputs(6080);
    outputs(644) <= not(layer0_outputs(4637));
    outputs(645) <= not(layer0_outputs(6477)) or (layer0_outputs(2159));
    outputs(646) <= not(layer0_outputs(6024));
    outputs(647) <= not(layer0_outputs(2479));
    outputs(648) <= not(layer0_outputs(2860));
    outputs(649) <= not(layer0_outputs(3047));
    outputs(650) <= not(layer0_outputs(6498)) or (layer0_outputs(5280));
    outputs(651) <= (layer0_outputs(4825)) and not (layer0_outputs(749));
    outputs(652) <= not(layer0_outputs(2493));
    outputs(653) <= not(layer0_outputs(4584));
    outputs(654) <= (layer0_outputs(7666)) or (layer0_outputs(1350));
    outputs(655) <= layer0_outputs(164);
    outputs(656) <= layer0_outputs(6919);
    outputs(657) <= not(layer0_outputs(3099));
    outputs(658) <= (layer0_outputs(2664)) and not (layer0_outputs(4507));
    outputs(659) <= (layer0_outputs(2767)) and (layer0_outputs(4721));
    outputs(660) <= not(layer0_outputs(1446));
    outputs(661) <= not(layer0_outputs(1377));
    outputs(662) <= layer0_outputs(1925);
    outputs(663) <= not(layer0_outputs(3459));
    outputs(664) <= (layer0_outputs(4878)) and not (layer0_outputs(4585));
    outputs(665) <= not(layer0_outputs(6818));
    outputs(666) <= (layer0_outputs(1022)) and (layer0_outputs(6224));
    outputs(667) <= not(layer0_outputs(7537)) or (layer0_outputs(3842));
    outputs(668) <= (layer0_outputs(326)) and (layer0_outputs(5483));
    outputs(669) <= not(layer0_outputs(1305));
    outputs(670) <= (layer0_outputs(6475)) and (layer0_outputs(4489));
    outputs(671) <= not(layer0_outputs(6413)) or (layer0_outputs(5723));
    outputs(672) <= (layer0_outputs(5297)) or (layer0_outputs(4670));
    outputs(673) <= (layer0_outputs(6234)) or (layer0_outputs(5558));
    outputs(674) <= not(layer0_outputs(3870));
    outputs(675) <= not(layer0_outputs(2322)) or (layer0_outputs(1497));
    outputs(676) <= layer0_outputs(5630);
    outputs(677) <= not(layer0_outputs(322));
    outputs(678) <= not(layer0_outputs(953));
    outputs(679) <= not(layer0_outputs(5482));
    outputs(680) <= not(layer0_outputs(2783));
    outputs(681) <= not((layer0_outputs(1325)) xor (layer0_outputs(1784)));
    outputs(682) <= not(layer0_outputs(96));
    outputs(683) <= layer0_outputs(891);
    outputs(684) <= layer0_outputs(5745);
    outputs(685) <= (layer0_outputs(1692)) and not (layer0_outputs(6943));
    outputs(686) <= layer0_outputs(5643);
    outputs(687) <= not((layer0_outputs(1310)) and (layer0_outputs(6158)));
    outputs(688) <= not(layer0_outputs(4867));
    outputs(689) <= (layer0_outputs(6506)) and (layer0_outputs(1068));
    outputs(690) <= not((layer0_outputs(1253)) or (layer0_outputs(3677)));
    outputs(691) <= layer0_outputs(7022);
    outputs(692) <= not(layer0_outputs(3458));
    outputs(693) <= not(layer0_outputs(3344));
    outputs(694) <= layer0_outputs(3248);
    outputs(695) <= layer0_outputs(6823);
    outputs(696) <= not(layer0_outputs(4145));
    outputs(697) <= not(layer0_outputs(2366));
    outputs(698) <= (layer0_outputs(3606)) and (layer0_outputs(3541));
    outputs(699) <= not((layer0_outputs(6573)) and (layer0_outputs(3134)));
    outputs(700) <= (layer0_outputs(1801)) or (layer0_outputs(6947));
    outputs(701) <= (layer0_outputs(3970)) xor (layer0_outputs(5424));
    outputs(702) <= not(layer0_outputs(2301));
    outputs(703) <= not(layer0_outputs(16)) or (layer0_outputs(5828));
    outputs(704) <= (layer0_outputs(4324)) and not (layer0_outputs(779));
    outputs(705) <= layer0_outputs(7499);
    outputs(706) <= layer0_outputs(3821);
    outputs(707) <= not((layer0_outputs(1285)) or (layer0_outputs(1402)));
    outputs(708) <= (layer0_outputs(3665)) or (layer0_outputs(5381));
    outputs(709) <= not((layer0_outputs(4326)) xor (layer0_outputs(3669)));
    outputs(710) <= layer0_outputs(3087);
    outputs(711) <= (layer0_outputs(6636)) and not (layer0_outputs(3338));
    outputs(712) <= layer0_outputs(75);
    outputs(713) <= layer0_outputs(552);
    outputs(714) <= layer0_outputs(6553);
    outputs(715) <= not(layer0_outputs(5231)) or (layer0_outputs(1087));
    outputs(716) <= (layer0_outputs(496)) or (layer0_outputs(992));
    outputs(717) <= layer0_outputs(4304);
    outputs(718) <= (layer0_outputs(4373)) and not (layer0_outputs(3140));
    outputs(719) <= not(layer0_outputs(310));
    outputs(720) <= layer0_outputs(3876);
    outputs(721) <= not(layer0_outputs(3759));
    outputs(722) <= layer0_outputs(3222);
    outputs(723) <= (layer0_outputs(1907)) and (layer0_outputs(4754));
    outputs(724) <= not(layer0_outputs(6746));
    outputs(725) <= layer0_outputs(6882);
    outputs(726) <= not((layer0_outputs(4855)) or (layer0_outputs(5677)));
    outputs(727) <= layer0_outputs(1622);
    outputs(728) <= not((layer0_outputs(5103)) and (layer0_outputs(3075)));
    outputs(729) <= layer0_outputs(5818);
    outputs(730) <= layer0_outputs(500);
    outputs(731) <= not(layer0_outputs(4023));
    outputs(732) <= layer0_outputs(2174);
    outputs(733) <= layer0_outputs(1288);
    outputs(734) <= (layer0_outputs(5181)) or (layer0_outputs(7553));
    outputs(735) <= not(layer0_outputs(6697)) or (layer0_outputs(1997));
    outputs(736) <= not(layer0_outputs(521));
    outputs(737) <= (layer0_outputs(7574)) or (layer0_outputs(4330));
    outputs(738) <= layer0_outputs(6303);
    outputs(739) <= not((layer0_outputs(1096)) xor (layer0_outputs(149)));
    outputs(740) <= (layer0_outputs(4605)) and (layer0_outputs(3630));
    outputs(741) <= not(layer0_outputs(7287));
    outputs(742) <= (layer0_outputs(5787)) and not (layer0_outputs(5603));
    outputs(743) <= (layer0_outputs(5909)) and (layer0_outputs(4486));
    outputs(744) <= not(layer0_outputs(1760));
    outputs(745) <= (layer0_outputs(2448)) and not (layer0_outputs(5190));
    outputs(746) <= not(layer0_outputs(1352));
    outputs(747) <= not(layer0_outputs(6936)) or (layer0_outputs(7071));
    outputs(748) <= (layer0_outputs(574)) xor (layer0_outputs(227));
    outputs(749) <= not(layer0_outputs(4979));
    outputs(750) <= not(layer0_outputs(4062));
    outputs(751) <= not(layer0_outputs(798)) or (layer0_outputs(1055));
    outputs(752) <= layer0_outputs(1477);
    outputs(753) <= not(layer0_outputs(4423));
    outputs(754) <= not(layer0_outputs(4747));
    outputs(755) <= (layer0_outputs(2337)) and not (layer0_outputs(554));
    outputs(756) <= layer0_outputs(2143);
    outputs(757) <= (layer0_outputs(3357)) and (layer0_outputs(7083));
    outputs(758) <= (layer0_outputs(2686)) and not (layer0_outputs(316));
    outputs(759) <= (layer0_outputs(2208)) or (layer0_outputs(1945));
    outputs(760) <= not((layer0_outputs(5676)) and (layer0_outputs(5753)));
    outputs(761) <= not((layer0_outputs(309)) xor (layer0_outputs(4590)));
    outputs(762) <= (layer0_outputs(4603)) or (layer0_outputs(3015));
    outputs(763) <= layer0_outputs(6023);
    outputs(764) <= layer0_outputs(4324);
    outputs(765) <= not(layer0_outputs(2965));
    outputs(766) <= not(layer0_outputs(1151));
    outputs(767) <= layer0_outputs(3656);
    outputs(768) <= (layer0_outputs(3556)) and not (layer0_outputs(5609));
    outputs(769) <= (layer0_outputs(5148)) and not (layer0_outputs(7339));
    outputs(770) <= not((layer0_outputs(174)) xor (layer0_outputs(3847)));
    outputs(771) <= not((layer0_outputs(3480)) or (layer0_outputs(6399)));
    outputs(772) <= (layer0_outputs(3086)) and (layer0_outputs(4544));
    outputs(773) <= (layer0_outputs(375)) and not (layer0_outputs(5407));
    outputs(774) <= not((layer0_outputs(788)) or (layer0_outputs(3751)));
    outputs(775) <= (layer0_outputs(2683)) xor (layer0_outputs(3080));
    outputs(776) <= (layer0_outputs(1518)) and (layer0_outputs(3060));
    outputs(777) <= (layer0_outputs(4574)) and (layer0_outputs(3203));
    outputs(778) <= not(layer0_outputs(4290));
    outputs(779) <= (layer0_outputs(2095)) and not (layer0_outputs(4746));
    outputs(780) <= not(layer0_outputs(3791));
    outputs(781) <= layer0_outputs(3004);
    outputs(782) <= (layer0_outputs(7053)) and not (layer0_outputs(849));
    outputs(783) <= not(layer0_outputs(2014));
    outputs(784) <= (layer0_outputs(5629)) and not (layer0_outputs(5688));
    outputs(785) <= not(layer0_outputs(5757));
    outputs(786) <= (layer0_outputs(3311)) and not (layer0_outputs(5286));
    outputs(787) <= layer0_outputs(4034);
    outputs(788) <= not(layer0_outputs(4875));
    outputs(789) <= (layer0_outputs(553)) and (layer0_outputs(2883));
    outputs(790) <= (layer0_outputs(6958)) and not (layer0_outputs(5588));
    outputs(791) <= not(layer0_outputs(7054));
    outputs(792) <= (layer0_outputs(1857)) and not (layer0_outputs(4513));
    outputs(793) <= not(layer0_outputs(263)) or (layer0_outputs(1950));
    outputs(794) <= not((layer0_outputs(5546)) or (layer0_outputs(7527)));
    outputs(795) <= not((layer0_outputs(990)) xor (layer0_outputs(1405)));
    outputs(796) <= not(layer0_outputs(7120));
    outputs(797) <= (layer0_outputs(7117)) and (layer0_outputs(5121));
    outputs(798) <= (layer0_outputs(1863)) and not (layer0_outputs(364));
    outputs(799) <= (layer0_outputs(3417)) and (layer0_outputs(672));
    outputs(800) <= not((layer0_outputs(5617)) xor (layer0_outputs(2795)));
    outputs(801) <= (layer0_outputs(6949)) and not (layer0_outputs(290));
    outputs(802) <= layer0_outputs(4271);
    outputs(803) <= (layer0_outputs(760)) and (layer0_outputs(4038));
    outputs(804) <= (layer0_outputs(4725)) xor (layer0_outputs(4904));
    outputs(805) <= (layer0_outputs(2070)) and (layer0_outputs(5726));
    outputs(806) <= (layer0_outputs(3816)) and (layer0_outputs(1501));
    outputs(807) <= (layer0_outputs(3856)) and not (layer0_outputs(340));
    outputs(808) <= (layer0_outputs(602)) xor (layer0_outputs(256));
    outputs(809) <= (layer0_outputs(1990)) and not (layer0_outputs(7224));
    outputs(810) <= (layer0_outputs(7669)) and not (layer0_outputs(6576));
    outputs(811) <= not((layer0_outputs(5496)) xor (layer0_outputs(1079)));
    outputs(812) <= not((layer0_outputs(4385)) or (layer0_outputs(2872)));
    outputs(813) <= (layer0_outputs(5821)) and (layer0_outputs(7556));
    outputs(814) <= layer0_outputs(6025);
    outputs(815) <= (layer0_outputs(4251)) and not (layer0_outputs(1769));
    outputs(816) <= (layer0_outputs(5989)) and not (layer0_outputs(6134));
    outputs(817) <= not((layer0_outputs(5967)) or (layer0_outputs(973)));
    outputs(818) <= (layer0_outputs(4251)) xor (layer0_outputs(5498));
    outputs(819) <= (layer0_outputs(4922)) and (layer0_outputs(5480));
    outputs(820) <= not((layer0_outputs(1315)) xor (layer0_outputs(5134)));
    outputs(821) <= (layer0_outputs(5300)) xor (layer0_outputs(127));
    outputs(822) <= layer0_outputs(5387);
    outputs(823) <= layer0_outputs(7163);
    outputs(824) <= layer0_outputs(5034);
    outputs(825) <= layer0_outputs(4953);
    outputs(826) <= (layer0_outputs(4288)) and not (layer0_outputs(3529));
    outputs(827) <= (layer0_outputs(6843)) and (layer0_outputs(454));
    outputs(828) <= not((layer0_outputs(2399)) or (layer0_outputs(3593)));
    outputs(829) <= (layer0_outputs(6874)) xor (layer0_outputs(5710));
    outputs(830) <= not((layer0_outputs(2779)) or (layer0_outputs(1076)));
    outputs(831) <= not((layer0_outputs(3131)) and (layer0_outputs(106)));
    outputs(832) <= (layer0_outputs(2722)) xor (layer0_outputs(5282));
    outputs(833) <= (layer0_outputs(3212)) and (layer0_outputs(4057));
    outputs(834) <= (layer0_outputs(7090)) and (layer0_outputs(4525));
    outputs(835) <= (layer0_outputs(4893)) and not (layer0_outputs(5592));
    outputs(836) <= not(layer0_outputs(1931));
    outputs(837) <= (layer0_outputs(7251)) and not (layer0_outputs(1562));
    outputs(838) <= not((layer0_outputs(4182)) or (layer0_outputs(4210)));
    outputs(839) <= layer0_outputs(7112);
    outputs(840) <= not((layer0_outputs(3549)) xor (layer0_outputs(2420)));
    outputs(841) <= (layer0_outputs(5817)) and not (layer0_outputs(4054));
    outputs(842) <= (layer0_outputs(7470)) and not (layer0_outputs(6305));
    outputs(843) <= not(layer0_outputs(1729));
    outputs(844) <= (layer0_outputs(29)) and (layer0_outputs(6618));
    outputs(845) <= (layer0_outputs(658)) and not (layer0_outputs(7265));
    outputs(846) <= (layer0_outputs(3338)) and not (layer0_outputs(2313));
    outputs(847) <= layer0_outputs(6754);
    outputs(848) <= not(layer0_outputs(2878));
    outputs(849) <= not(layer0_outputs(1595));
    outputs(850) <= (layer0_outputs(6207)) and not (layer0_outputs(2254));
    outputs(851) <= (layer0_outputs(2767)) and not (layer0_outputs(73));
    outputs(852) <= not((layer0_outputs(731)) or (layer0_outputs(730)));
    outputs(853) <= not((layer0_outputs(6319)) or (layer0_outputs(1275)));
    outputs(854) <= not((layer0_outputs(5014)) or (layer0_outputs(5468)));
    outputs(855) <= not((layer0_outputs(5366)) xor (layer0_outputs(7199)));
    outputs(856) <= (layer0_outputs(7147)) and not (layer0_outputs(5290));
    outputs(857) <= not((layer0_outputs(3289)) xor (layer0_outputs(6557)));
    outputs(858) <= not((layer0_outputs(7225)) or (layer0_outputs(2191)));
    outputs(859) <= (layer0_outputs(4702)) and not (layer0_outputs(6694));
    outputs(860) <= not(layer0_outputs(3623));
    outputs(861) <= (layer0_outputs(5605)) and (layer0_outputs(66));
    outputs(862) <= layer0_outputs(2581);
    outputs(863) <= not(layer0_outputs(6853));
    outputs(864) <= (layer0_outputs(2954)) and not (layer0_outputs(4123));
    outputs(865) <= not((layer0_outputs(216)) or (layer0_outputs(2946)));
    outputs(866) <= (layer0_outputs(5646)) and not (layer0_outputs(6247));
    outputs(867) <= (layer0_outputs(277)) and (layer0_outputs(2497));
    outputs(868) <= not(layer0_outputs(4188));
    outputs(869) <= (layer0_outputs(7564)) and (layer0_outputs(5841));
    outputs(870) <= '0';
    outputs(871) <= not(layer0_outputs(4704));
    outputs(872) <= (layer0_outputs(1980)) and not (layer0_outputs(275));
    outputs(873) <= not((layer0_outputs(7003)) or (layer0_outputs(425)));
    outputs(874) <= (layer0_outputs(2859)) and not (layer0_outputs(6900));
    outputs(875) <= (layer0_outputs(7672)) and not (layer0_outputs(4124));
    outputs(876) <= (layer0_outputs(684)) and not (layer0_outputs(961));
    outputs(877) <= not((layer0_outputs(6760)) or (layer0_outputs(6157)));
    outputs(878) <= not(layer0_outputs(457));
    outputs(879) <= layer0_outputs(2058);
    outputs(880) <= not(layer0_outputs(83));
    outputs(881) <= (layer0_outputs(2598)) and (layer0_outputs(7399));
    outputs(882) <= not((layer0_outputs(4050)) xor (layer0_outputs(53)));
    outputs(883) <= not(layer0_outputs(4872));
    outputs(884) <= not((layer0_outputs(1204)) or (layer0_outputs(912)));
    outputs(885) <= not((layer0_outputs(6812)) or (layer0_outputs(1761)));
    outputs(886) <= (layer0_outputs(1099)) and (layer0_outputs(6940));
    outputs(887) <= not((layer0_outputs(6340)) or (layer0_outputs(6785)));
    outputs(888) <= (layer0_outputs(6862)) and not (layer0_outputs(6214));
    outputs(889) <= (layer0_outputs(5116)) and not (layer0_outputs(1322));
    outputs(890) <= (layer0_outputs(7348)) and not (layer0_outputs(7301));
    outputs(891) <= (layer0_outputs(1725)) and not (layer0_outputs(5992));
    outputs(892) <= (layer0_outputs(5725)) and (layer0_outputs(5368));
    outputs(893) <= (layer0_outputs(5957)) and not (layer0_outputs(2202));
    outputs(894) <= not((layer0_outputs(464)) or (layer0_outputs(1665)));
    outputs(895) <= (layer0_outputs(2317)) xor (layer0_outputs(5150));
    outputs(896) <= layer0_outputs(93);
    outputs(897) <= (layer0_outputs(4060)) and not (layer0_outputs(6183));
    outputs(898) <= (layer0_outputs(4122)) and not (layer0_outputs(6886));
    outputs(899) <= not(layer0_outputs(4041));
    outputs(900) <= not((layer0_outputs(1695)) or (layer0_outputs(6826)));
    outputs(901) <= layer0_outputs(4040);
    outputs(902) <= (layer0_outputs(661)) and not (layer0_outputs(1774));
    outputs(903) <= '0';
    outputs(904) <= '0';
    outputs(905) <= not(layer0_outputs(2847));
    outputs(906) <= (layer0_outputs(2309)) and (layer0_outputs(3121));
    outputs(907) <= (layer0_outputs(6410)) xor (layer0_outputs(4745));
    outputs(908) <= (layer0_outputs(6914)) and not (layer0_outputs(6146));
    outputs(909) <= (layer0_outputs(5278)) and not (layer0_outputs(4680));
    outputs(910) <= (layer0_outputs(6526)) and (layer0_outputs(4191));
    outputs(911) <= not((layer0_outputs(6678)) or (layer0_outputs(2899)));
    outputs(912) <= (layer0_outputs(6924)) and not (layer0_outputs(5591));
    outputs(913) <= (layer0_outputs(2530)) and not (layer0_outputs(1324));
    outputs(914) <= (layer0_outputs(7121)) and not (layer0_outputs(519));
    outputs(915) <= (layer0_outputs(4295)) and (layer0_outputs(2735));
    outputs(916) <= not((layer0_outputs(3651)) xor (layer0_outputs(7566)));
    outputs(917) <= (layer0_outputs(5825)) and not (layer0_outputs(6750));
    outputs(918) <= not((layer0_outputs(4718)) xor (layer0_outputs(3945)));
    outputs(919) <= (layer0_outputs(5981)) and (layer0_outputs(2500));
    outputs(920) <= not((layer0_outputs(622)) or (layer0_outputs(3922)));
    outputs(921) <= layer0_outputs(2800);
    outputs(922) <= (layer0_outputs(1766)) and (layer0_outputs(2043));
    outputs(923) <= not((layer0_outputs(4739)) or (layer0_outputs(7007)));
    outputs(924) <= (layer0_outputs(3977)) and not (layer0_outputs(5886));
    outputs(925) <= (layer0_outputs(2834)) and not (layer0_outputs(685));
    outputs(926) <= layer0_outputs(3874);
    outputs(927) <= not((layer0_outputs(5824)) or (layer0_outputs(1219)));
    outputs(928) <= not((layer0_outputs(7246)) or (layer0_outputs(4700)));
    outputs(929) <= (layer0_outputs(1787)) and (layer0_outputs(2929));
    outputs(930) <= (layer0_outputs(841)) and not (layer0_outputs(3605));
    outputs(931) <= (layer0_outputs(3956)) and not (layer0_outputs(3944));
    outputs(932) <= layer0_outputs(6369);
    outputs(933) <= (layer0_outputs(725)) and not (layer0_outputs(4860));
    outputs(934) <= not((layer0_outputs(5787)) or (layer0_outputs(7661)));
    outputs(935) <= (layer0_outputs(1299)) and (layer0_outputs(2362));
    outputs(936) <= (layer0_outputs(3199)) and not (layer0_outputs(6832));
    outputs(937) <= layer0_outputs(6072);
    outputs(938) <= (layer0_outputs(6447)) xor (layer0_outputs(1205));
    outputs(939) <= (layer0_outputs(1750)) and not (layer0_outputs(1368));
    outputs(940) <= not(layer0_outputs(4613));
    outputs(941) <= '0';
    outputs(942) <= not((layer0_outputs(1300)) or (layer0_outputs(1484)));
    outputs(943) <= (layer0_outputs(1944)) xor (layer0_outputs(987));
    outputs(944) <= (layer0_outputs(1496)) and not (layer0_outputs(5533));
    outputs(945) <= not((layer0_outputs(3661)) xor (layer0_outputs(859)));
    outputs(946) <= not((layer0_outputs(1110)) xor (layer0_outputs(3348)));
    outputs(947) <= (layer0_outputs(1631)) and not (layer0_outputs(4888));
    outputs(948) <= (layer0_outputs(3209)) and (layer0_outputs(4796));
    outputs(949) <= (layer0_outputs(1586)) and not (layer0_outputs(3185));
    outputs(950) <= (layer0_outputs(2533)) and not (layer0_outputs(3483));
    outputs(951) <= '0';
    outputs(952) <= (layer0_outputs(59)) and not (layer0_outputs(6015));
    outputs(953) <= (layer0_outputs(5691)) and not (layer0_outputs(559));
    outputs(954) <= (layer0_outputs(870)) and not (layer0_outputs(6276));
    outputs(955) <= (layer0_outputs(2178)) and not (layer0_outputs(2264));
    outputs(956) <= not(layer0_outputs(186));
    outputs(957) <= (layer0_outputs(2381)) and not (layer0_outputs(5345));
    outputs(958) <= not((layer0_outputs(3791)) or (layer0_outputs(5299)));
    outputs(959) <= (layer0_outputs(6613)) and (layer0_outputs(162));
    outputs(960) <= (layer0_outputs(6824)) and not (layer0_outputs(5252));
    outputs(961) <= not(layer0_outputs(756));
    outputs(962) <= (layer0_outputs(4645)) xor (layer0_outputs(1638));
    outputs(963) <= (layer0_outputs(6002)) xor (layer0_outputs(5161));
    outputs(964) <= not((layer0_outputs(2416)) xor (layer0_outputs(509)));
    outputs(965) <= (layer0_outputs(1251)) and not (layer0_outputs(2346));
    outputs(966) <= layer0_outputs(2912);
    outputs(967) <= not(layer0_outputs(720));
    outputs(968) <= (layer0_outputs(6147)) and (layer0_outputs(4426));
    outputs(969) <= not((layer0_outputs(5163)) or (layer0_outputs(4863)));
    outputs(970) <= (layer0_outputs(7570)) and not (layer0_outputs(6221));
    outputs(971) <= (layer0_outputs(3050)) and (layer0_outputs(5009));
    outputs(972) <= not(layer0_outputs(5374));
    outputs(973) <= (layer0_outputs(1461)) and (layer0_outputs(7443));
    outputs(974) <= (layer0_outputs(2302)) and (layer0_outputs(530));
    outputs(975) <= (layer0_outputs(7622)) and not (layer0_outputs(1818));
    outputs(976) <= not((layer0_outputs(6052)) or (layer0_outputs(5561)));
    outputs(977) <= not(layer0_outputs(3991));
    outputs(978) <= (layer0_outputs(5854)) and not (layer0_outputs(5818));
    outputs(979) <= (layer0_outputs(5342)) xor (layer0_outputs(592));
    outputs(980) <= (layer0_outputs(3473)) and not (layer0_outputs(6128));
    outputs(981) <= (layer0_outputs(3140)) and not (layer0_outputs(4083));
    outputs(982) <= not((layer0_outputs(4361)) or (layer0_outputs(7012)));
    outputs(983) <= '0';
    outputs(984) <= layer0_outputs(2415);
    outputs(985) <= (layer0_outputs(1831)) and (layer0_outputs(1939));
    outputs(986) <= layer0_outputs(5367);
    outputs(987) <= '0';
    outputs(988) <= not((layer0_outputs(5167)) or (layer0_outputs(569)));
    outputs(989) <= (layer0_outputs(1822)) and (layer0_outputs(4634));
    outputs(990) <= layer0_outputs(938);
    outputs(991) <= (layer0_outputs(3097)) and (layer0_outputs(5843));
    outputs(992) <= not((layer0_outputs(3678)) or (layer0_outputs(520)));
    outputs(993) <= not((layer0_outputs(1542)) or (layer0_outputs(1978)));
    outputs(994) <= (layer0_outputs(1887)) and not (layer0_outputs(567));
    outputs(995) <= not((layer0_outputs(6891)) xor (layer0_outputs(6738)));
    outputs(996) <= not((layer0_outputs(436)) xor (layer0_outputs(5318)));
    outputs(997) <= not((layer0_outputs(3150)) or (layer0_outputs(1006)));
    outputs(998) <= (layer0_outputs(4954)) and (layer0_outputs(7497));
    outputs(999) <= (layer0_outputs(4811)) and not (layer0_outputs(3795));
    outputs(1000) <= layer0_outputs(58);
    outputs(1001) <= not((layer0_outputs(3985)) or (layer0_outputs(433)));
    outputs(1002) <= layer0_outputs(3433);
    outputs(1003) <= (layer0_outputs(1384)) xor (layer0_outputs(2975));
    outputs(1004) <= not((layer0_outputs(6079)) xor (layer0_outputs(2219)));
    outputs(1005) <= not((layer0_outputs(2055)) or (layer0_outputs(154)));
    outputs(1006) <= not((layer0_outputs(2945)) xor (layer0_outputs(1823)));
    outputs(1007) <= (layer0_outputs(2985)) and not (layer0_outputs(7398));
    outputs(1008) <= (layer0_outputs(6594)) and not (layer0_outputs(229));
    outputs(1009) <= layer0_outputs(4634);
    outputs(1010) <= layer0_outputs(1614);
    outputs(1011) <= (layer0_outputs(2422)) and not (layer0_outputs(4566));
    outputs(1012) <= not((layer0_outputs(7299)) or (layer0_outputs(2728)));
    outputs(1013) <= (layer0_outputs(4532)) and (layer0_outputs(723));
    outputs(1014) <= not(layer0_outputs(3596));
    outputs(1015) <= (layer0_outputs(4705)) and not (layer0_outputs(6644));
    outputs(1016) <= (layer0_outputs(6420)) and not (layer0_outputs(4919));
    outputs(1017) <= (layer0_outputs(6986)) and (layer0_outputs(1651));
    outputs(1018) <= not((layer0_outputs(3196)) xor (layer0_outputs(6769)));
    outputs(1019) <= (layer0_outputs(4892)) and (layer0_outputs(4703));
    outputs(1020) <= (layer0_outputs(4965)) and not (layer0_outputs(6062));
    outputs(1021) <= (layer0_outputs(2479)) and not (layer0_outputs(4281));
    outputs(1022) <= not((layer0_outputs(6333)) or (layer0_outputs(3250)));
    outputs(1023) <= not((layer0_outputs(1155)) or (layer0_outputs(557)));
    outputs(1024) <= layer0_outputs(3282);
    outputs(1025) <= (layer0_outputs(626)) and (layer0_outputs(4461));
    outputs(1026) <= not(layer0_outputs(5085)) or (layer0_outputs(2281));
    outputs(1027) <= (layer0_outputs(5316)) and (layer0_outputs(5050));
    outputs(1028) <= (layer0_outputs(7478)) and (layer0_outputs(5185));
    outputs(1029) <= not((layer0_outputs(5008)) or (layer0_outputs(3056)));
    outputs(1030) <= (layer0_outputs(739)) xor (layer0_outputs(6338));
    outputs(1031) <= (layer0_outputs(149)) and not (layer0_outputs(6226));
    outputs(1032) <= layer0_outputs(5676);
    outputs(1033) <= not(layer0_outputs(1396));
    outputs(1034) <= (layer0_outputs(1400)) and not (layer0_outputs(3168));
    outputs(1035) <= not((layer0_outputs(6935)) xor (layer0_outputs(3964)));
    outputs(1036) <= (layer0_outputs(2015)) and not (layer0_outputs(5681));
    outputs(1037) <= (layer0_outputs(5611)) and not (layer0_outputs(3393));
    outputs(1038) <= (layer0_outputs(4362)) and not (layer0_outputs(711));
    outputs(1039) <= layer0_outputs(3787);
    outputs(1040) <= (layer0_outputs(6377)) and (layer0_outputs(4086));
    outputs(1041) <= (layer0_outputs(3300)) and not (layer0_outputs(7341));
    outputs(1042) <= (layer0_outputs(4864)) and not (layer0_outputs(357));
    outputs(1043) <= (layer0_outputs(3687)) xor (layer0_outputs(818));
    outputs(1044) <= (layer0_outputs(2119)) and not (layer0_outputs(1018));
    outputs(1045) <= not((layer0_outputs(7429)) or (layer0_outputs(5251)));
    outputs(1046) <= layer0_outputs(6603);
    outputs(1047) <= (layer0_outputs(7167)) and (layer0_outputs(125));
    outputs(1048) <= layer0_outputs(5082);
    outputs(1049) <= (layer0_outputs(6252)) and (layer0_outputs(3507));
    outputs(1050) <= (layer0_outputs(2552)) xor (layer0_outputs(3538));
    outputs(1051) <= not(layer0_outputs(2601));
    outputs(1052) <= (layer0_outputs(7255)) and not (layer0_outputs(7222));
    outputs(1053) <= layer0_outputs(3356);
    outputs(1054) <= (layer0_outputs(3468)) and not (layer0_outputs(4961));
    outputs(1055) <= layer0_outputs(5939);
    outputs(1056) <= (layer0_outputs(6442)) and not (layer0_outputs(5736));
    outputs(1057) <= layer0_outputs(1827);
    outputs(1058) <= (layer0_outputs(7425)) and not (layer0_outputs(6830));
    outputs(1059) <= (layer0_outputs(329)) and not (layer0_outputs(3326));
    outputs(1060) <= (layer0_outputs(5966)) and (layer0_outputs(4205));
    outputs(1061) <= (layer0_outputs(3570)) and (layer0_outputs(5833));
    outputs(1062) <= layer0_outputs(2944);
    outputs(1063) <= not((layer0_outputs(837)) or (layer0_outputs(2163)));
    outputs(1064) <= not(layer0_outputs(1504));
    outputs(1065) <= (layer0_outputs(3999)) and not (layer0_outputs(6435));
    outputs(1066) <= not(layer0_outputs(2041));
    outputs(1067) <= (layer0_outputs(1123)) and (layer0_outputs(2101));
    outputs(1068) <= not((layer0_outputs(6474)) xor (layer0_outputs(5162)));
    outputs(1069) <= layer0_outputs(2391);
    outputs(1070) <= (layer0_outputs(5893)) and not (layer0_outputs(4566));
    outputs(1071) <= layer0_outputs(7297);
    outputs(1072) <= (layer0_outputs(2757)) xor (layer0_outputs(6422));
    outputs(1073) <= (layer0_outputs(2357)) and not (layer0_outputs(587));
    outputs(1074) <= (layer0_outputs(1561)) and not (layer0_outputs(3617));
    outputs(1075) <= (layer0_outputs(6500)) xor (layer0_outputs(7005));
    outputs(1076) <= not((layer0_outputs(508)) or (layer0_outputs(4076)));
    outputs(1077) <= (layer0_outputs(6127)) and (layer0_outputs(6766));
    outputs(1078) <= (layer0_outputs(121)) and not (layer0_outputs(3848));
    outputs(1079) <= (layer0_outputs(1926)) and not (layer0_outputs(229));
    outputs(1080) <= (layer0_outputs(5455)) and not (layer0_outputs(170));
    outputs(1081) <= layer0_outputs(5184);
    outputs(1082) <= (layer0_outputs(709)) and not (layer0_outputs(4571));
    outputs(1083) <= (layer0_outputs(924)) and (layer0_outputs(7342));
    outputs(1084) <= (layer0_outputs(7450)) and not (layer0_outputs(6744));
    outputs(1085) <= not((layer0_outputs(3492)) or (layer0_outputs(461)));
    outputs(1086) <= not((layer0_outputs(4524)) or (layer0_outputs(6636)));
    outputs(1087) <= not((layer0_outputs(5186)) or (layer0_outputs(1999)));
    outputs(1088) <= (layer0_outputs(1926)) and (layer0_outputs(3962));
    outputs(1089) <= (layer0_outputs(3467)) and (layer0_outputs(3700));
    outputs(1090) <= (layer0_outputs(2264)) and not (layer0_outputs(3217));
    outputs(1091) <= (layer0_outputs(3354)) and not (layer0_outputs(4033));
    outputs(1092) <= not(layer0_outputs(1327));
    outputs(1093) <= layer0_outputs(4354);
    outputs(1094) <= not((layer0_outputs(4803)) xor (layer0_outputs(130)));
    outputs(1095) <= not(layer0_outputs(4729));
    outputs(1096) <= not(layer0_outputs(1041));
    outputs(1097) <= layer0_outputs(6238);
    outputs(1098) <= (layer0_outputs(2250)) and not (layer0_outputs(4336));
    outputs(1099) <= layer0_outputs(762);
    outputs(1100) <= layer0_outputs(2989);
    outputs(1101) <= (layer0_outputs(447)) and (layer0_outputs(5832));
    outputs(1102) <= (layer0_outputs(4653)) and not (layer0_outputs(4478));
    outputs(1103) <= not(layer0_outputs(1372));
    outputs(1104) <= (layer0_outputs(6913)) xor (layer0_outputs(7452));
    outputs(1105) <= (layer0_outputs(6296)) and not (layer0_outputs(2494));
    outputs(1106) <= (layer0_outputs(7129)) and (layer0_outputs(3764));
    outputs(1107) <= (layer0_outputs(7626)) and not (layer0_outputs(5634));
    outputs(1108) <= not(layer0_outputs(4455));
    outputs(1109) <= (layer0_outputs(2614)) and not (layer0_outputs(6640));
    outputs(1110) <= layer0_outputs(6283);
    outputs(1111) <= (layer0_outputs(2466)) xor (layer0_outputs(5058));
    outputs(1112) <= (layer0_outputs(5837)) and (layer0_outputs(1611));
    outputs(1113) <= '0';
    outputs(1114) <= not((layer0_outputs(6174)) or (layer0_outputs(4359)));
    outputs(1115) <= (layer0_outputs(4468)) xor (layer0_outputs(3037));
    outputs(1116) <= (layer0_outputs(1071)) and not (layer0_outputs(7098));
    outputs(1117) <= not((layer0_outputs(612)) or (layer0_outputs(794)));
    outputs(1118) <= not(layer0_outputs(7214));
    outputs(1119) <= (layer0_outputs(5315)) xor (layer0_outputs(6844));
    outputs(1120) <= (layer0_outputs(6224)) xor (layer0_outputs(3946));
    outputs(1121) <= not(layer0_outputs(1137));
    outputs(1122) <= (layer0_outputs(7449)) and not (layer0_outputs(834));
    outputs(1123) <= (layer0_outputs(2435)) and not (layer0_outputs(6812));
    outputs(1124) <= not(layer0_outputs(4632));
    outputs(1125) <= not((layer0_outputs(7056)) xor (layer0_outputs(7455)));
    outputs(1126) <= (layer0_outputs(4352)) and (layer0_outputs(3843));
    outputs(1127) <= (layer0_outputs(6980)) and not (layer0_outputs(6778));
    outputs(1128) <= (layer0_outputs(2513)) and not (layer0_outputs(2882));
    outputs(1129) <= not(layer0_outputs(5264));
    outputs(1130) <= (layer0_outputs(4041)) and not (layer0_outputs(3972));
    outputs(1131) <= not(layer0_outputs(4031));
    outputs(1132) <= (layer0_outputs(2580)) and (layer0_outputs(1914));
    outputs(1133) <= not(layer0_outputs(1027));
    outputs(1134) <= (layer0_outputs(3341)) xor (layer0_outputs(663));
    outputs(1135) <= (layer0_outputs(1534)) and (layer0_outputs(3252));
    outputs(1136) <= not(layer0_outputs(3078));
    outputs(1137) <= (layer0_outputs(1448)) and not (layer0_outputs(1296));
    outputs(1138) <= (layer0_outputs(2100)) and not (layer0_outputs(5863));
    outputs(1139) <= not((layer0_outputs(1261)) or (layer0_outputs(337)));
    outputs(1140) <= not((layer0_outputs(1764)) or (layer0_outputs(5793)));
    outputs(1141) <= (layer0_outputs(851)) and not (layer0_outputs(55));
    outputs(1142) <= not(layer0_outputs(3016)) or (layer0_outputs(4856));
    outputs(1143) <= not(layer0_outputs(453));
    outputs(1144) <= (layer0_outputs(2034)) xor (layer0_outputs(2631));
    outputs(1145) <= layer0_outputs(947);
    outputs(1146) <= (layer0_outputs(876)) and not (layer0_outputs(1984));
    outputs(1147) <= not((layer0_outputs(1452)) xor (layer0_outputs(432)));
    outputs(1148) <= not((layer0_outputs(7361)) xor (layer0_outputs(5071)));
    outputs(1149) <= (layer0_outputs(3097)) and (layer0_outputs(6040));
    outputs(1150) <= (layer0_outputs(1397)) and not (layer0_outputs(2005));
    outputs(1151) <= (layer0_outputs(4535)) and not (layer0_outputs(668));
    outputs(1152) <= not((layer0_outputs(1998)) or (layer0_outputs(3197)));
    outputs(1153) <= not((layer0_outputs(3731)) xor (layer0_outputs(4174)));
    outputs(1154) <= not((layer0_outputs(3192)) or (layer0_outputs(5292)));
    outputs(1155) <= (layer0_outputs(2427)) and (layer0_outputs(3511));
    outputs(1156) <= layer0_outputs(4470);
    outputs(1157) <= not(layer0_outputs(1103));
    outputs(1158) <= not(layer0_outputs(5324));
    outputs(1159) <= (layer0_outputs(4075)) xor (layer0_outputs(1797));
    outputs(1160) <= not((layer0_outputs(5927)) or (layer0_outputs(6476)));
    outputs(1161) <= not(layer0_outputs(4633));
    outputs(1162) <= (layer0_outputs(1789)) and not (layer0_outputs(5519));
    outputs(1163) <= (layer0_outputs(2427)) and (layer0_outputs(7445));
    outputs(1164) <= (layer0_outputs(6212)) and not (layer0_outputs(7474));
    outputs(1165) <= (layer0_outputs(7086)) xor (layer0_outputs(923));
    outputs(1166) <= (layer0_outputs(1819)) and not (layer0_outputs(6183));
    outputs(1167) <= (layer0_outputs(5118)) and (layer0_outputs(6490));
    outputs(1168) <= not(layer0_outputs(1664));
    outputs(1169) <= (layer0_outputs(1375)) and not (layer0_outputs(2092));
    outputs(1170) <= (layer0_outputs(2484)) and not (layer0_outputs(6664));
    outputs(1171) <= not((layer0_outputs(6517)) xor (layer0_outputs(3424)));
    outputs(1172) <= (layer0_outputs(2566)) and (layer0_outputs(1858));
    outputs(1173) <= not(layer0_outputs(6725));
    outputs(1174) <= not(layer0_outputs(630));
    outputs(1175) <= (layer0_outputs(2798)) and not (layer0_outputs(3773));
    outputs(1176) <= not((layer0_outputs(4122)) xor (layer0_outputs(4520)));
    outputs(1177) <= not((layer0_outputs(2587)) or (layer0_outputs(7392)));
    outputs(1178) <= (layer0_outputs(698)) and not (layer0_outputs(5022));
    outputs(1179) <= (layer0_outputs(657)) and not (layer0_outputs(1503));
    outputs(1180) <= not((layer0_outputs(7358)) or (layer0_outputs(1654)));
    outputs(1181) <= not(layer0_outputs(7227));
    outputs(1182) <= (layer0_outputs(1632)) and not (layer0_outputs(7374));
    outputs(1183) <= not((layer0_outputs(4812)) xor (layer0_outputs(5302)));
    outputs(1184) <= (layer0_outputs(2610)) and not (layer0_outputs(5268));
    outputs(1185) <= (layer0_outputs(5136)) and (layer0_outputs(93));
    outputs(1186) <= (layer0_outputs(442)) and not (layer0_outputs(3177));
    outputs(1187) <= layer0_outputs(2518);
    outputs(1188) <= (layer0_outputs(7424)) and not (layer0_outputs(6708));
    outputs(1189) <= not(layer0_outputs(4980));
    outputs(1190) <= (layer0_outputs(4491)) and not (layer0_outputs(956));
    outputs(1191) <= not((layer0_outputs(4795)) xor (layer0_outputs(3432)));
    outputs(1192) <= not((layer0_outputs(4991)) or (layer0_outputs(5713)));
    outputs(1193) <= (layer0_outputs(3142)) and (layer0_outputs(5236));
    outputs(1194) <= layer0_outputs(6423);
    outputs(1195) <= (layer0_outputs(4118)) and not (layer0_outputs(4239));
    outputs(1196) <= not((layer0_outputs(1901)) or (layer0_outputs(1662)));
    outputs(1197) <= (layer0_outputs(6114)) xor (layer0_outputs(1529));
    outputs(1198) <= (layer0_outputs(4497)) and not (layer0_outputs(1188));
    outputs(1199) <= layer0_outputs(3771);
    outputs(1200) <= layer0_outputs(298);
    outputs(1201) <= (layer0_outputs(6085)) and (layer0_outputs(1091));
    outputs(1202) <= layer0_outputs(6824);
    outputs(1203) <= (layer0_outputs(4411)) and not (layer0_outputs(1900));
    outputs(1204) <= (layer0_outputs(863)) and not (layer0_outputs(1046));
    outputs(1205) <= (layer0_outputs(843)) xor (layer0_outputs(4261));
    outputs(1206) <= (layer0_outputs(4478)) xor (layer0_outputs(4671));
    outputs(1207) <= not(layer0_outputs(4337));
    outputs(1208) <= (layer0_outputs(3846)) and not (layer0_outputs(6099));
    outputs(1209) <= not((layer0_outputs(5248)) or (layer0_outputs(5399)));
    outputs(1210) <= (layer0_outputs(1088)) and (layer0_outputs(3366));
    outputs(1211) <= layer0_outputs(2089);
    outputs(1212) <= (layer0_outputs(7656)) and not (layer0_outputs(5433));
    outputs(1213) <= (layer0_outputs(4870)) and not (layer0_outputs(2253));
    outputs(1214) <= not(layer0_outputs(7204));
    outputs(1215) <= (layer0_outputs(994)) xor (layer0_outputs(3645));
    outputs(1216) <= not((layer0_outputs(776)) or (layer0_outputs(7439)));
    outputs(1217) <= not(layer0_outputs(6219));
    outputs(1218) <= not((layer0_outputs(6505)) or (layer0_outputs(3266)));
    outputs(1219) <= not((layer0_outputs(5301)) or (layer0_outputs(7560)));
    outputs(1220) <= (layer0_outputs(6811)) and (layer0_outputs(536));
    outputs(1221) <= (layer0_outputs(4594)) and not (layer0_outputs(5057));
    outputs(1222) <= (layer0_outputs(3535)) and (layer0_outputs(1360));
    outputs(1223) <= (layer0_outputs(3639)) and not (layer0_outputs(1301));
    outputs(1224) <= not((layer0_outputs(3235)) or (layer0_outputs(6513)));
    outputs(1225) <= layer0_outputs(3846);
    outputs(1226) <= (layer0_outputs(328)) and (layer0_outputs(3021));
    outputs(1227) <= not((layer0_outputs(829)) or (layer0_outputs(6465)));
    outputs(1228) <= (layer0_outputs(3066)) and (layer0_outputs(5156));
    outputs(1229) <= (layer0_outputs(2529)) xor (layer0_outputs(3566));
    outputs(1230) <= layer0_outputs(2487);
    outputs(1231) <= (layer0_outputs(1320)) xor (layer0_outputs(1701));
    outputs(1232) <= (layer0_outputs(3494)) xor (layer0_outputs(5931));
    outputs(1233) <= (layer0_outputs(342)) and not (layer0_outputs(6199));
    outputs(1234) <= (layer0_outputs(1434)) xor (layer0_outputs(3473));
    outputs(1235) <= (layer0_outputs(5414)) and not (layer0_outputs(2555));
    outputs(1236) <= not(layer0_outputs(4274)) or (layer0_outputs(6661));
    outputs(1237) <= not(layer0_outputs(7550));
    outputs(1238) <= not(layer0_outputs(1721));
    outputs(1239) <= (layer0_outputs(1936)) and (layer0_outputs(6051));
    outputs(1240) <= (layer0_outputs(1053)) and not (layer0_outputs(2271));
    outputs(1241) <= (layer0_outputs(3804)) and (layer0_outputs(3408));
    outputs(1242) <= (layer0_outputs(5174)) xor (layer0_outputs(3522));
    outputs(1243) <= (layer0_outputs(354)) and not (layer0_outputs(6316));
    outputs(1244) <= layer0_outputs(5175);
    outputs(1245) <= (layer0_outputs(4121)) and not (layer0_outputs(5108));
    outputs(1246) <= (layer0_outputs(2929)) and not (layer0_outputs(1924));
    outputs(1247) <= (layer0_outputs(7138)) and not (layer0_outputs(5991));
    outputs(1248) <= not((layer0_outputs(3812)) or (layer0_outputs(3262)));
    outputs(1249) <= (layer0_outputs(6177)) and not (layer0_outputs(4350));
    outputs(1250) <= not(layer0_outputs(3958));
    outputs(1251) <= not((layer0_outputs(1960)) or (layer0_outputs(4357)));
    outputs(1252) <= (layer0_outputs(6729)) and (layer0_outputs(6930));
    outputs(1253) <= not((layer0_outputs(856)) or (layer0_outputs(5855)));
    outputs(1254) <= (layer0_outputs(5714)) xor (layer0_outputs(6520));
    outputs(1255) <= (layer0_outputs(100)) and (layer0_outputs(1716));
    outputs(1256) <= not((layer0_outputs(1283)) or (layer0_outputs(7657)));
    outputs(1257) <= not(layer0_outputs(3469));
    outputs(1258) <= '0';
    outputs(1259) <= (layer0_outputs(4984)) and (layer0_outputs(4315));
    outputs(1260) <= not(layer0_outputs(1163));
    outputs(1261) <= layer0_outputs(86);
    outputs(1262) <= layer0_outputs(2151);
    outputs(1263) <= (layer0_outputs(6415)) and not (layer0_outputs(2615));
    outputs(1264) <= (layer0_outputs(3954)) and not (layer0_outputs(7364));
    outputs(1265) <= layer0_outputs(5975);
    outputs(1266) <= not(layer0_outputs(6567));
    outputs(1267) <= layer0_outputs(782);
    outputs(1268) <= (layer0_outputs(5551)) and (layer0_outputs(472));
    outputs(1269) <= (layer0_outputs(5140)) and not (layer0_outputs(4851));
    outputs(1270) <= layer0_outputs(1711);
    outputs(1271) <= layer0_outputs(6971);
    outputs(1272) <= (layer0_outputs(995)) and not (layer0_outputs(4670));
    outputs(1273) <= layer0_outputs(6710);
    outputs(1274) <= (layer0_outputs(6654)) and (layer0_outputs(746));
    outputs(1275) <= (layer0_outputs(927)) and not (layer0_outputs(784));
    outputs(1276) <= not((layer0_outputs(2370)) xor (layer0_outputs(3932)));
    outputs(1277) <= (layer0_outputs(6862)) and not (layer0_outputs(778));
    outputs(1278) <= (layer0_outputs(6702)) and (layer0_outputs(957));
    outputs(1279) <= not((layer0_outputs(3156)) or (layer0_outputs(79)));
    outputs(1280) <= layer0_outputs(6687);
    outputs(1281) <= layer0_outputs(6563);
    outputs(1282) <= not(layer0_outputs(7563));
    outputs(1283) <= not((layer0_outputs(1305)) xor (layer0_outputs(3556)));
    outputs(1284) <= not(layer0_outputs(3579));
    outputs(1285) <= not(layer0_outputs(2339));
    outputs(1286) <= not((layer0_outputs(2602)) or (layer0_outputs(2717)));
    outputs(1287) <= (layer0_outputs(1050)) and (layer0_outputs(2844));
    outputs(1288) <= (layer0_outputs(1498)) and (layer0_outputs(1133));
    outputs(1289) <= layer0_outputs(5009);
    outputs(1290) <= (layer0_outputs(171)) and not (layer0_outputs(6099));
    outputs(1291) <= (layer0_outputs(4090)) and (layer0_outputs(7640));
    outputs(1292) <= (layer0_outputs(2530)) xor (layer0_outputs(1982));
    outputs(1293) <= (layer0_outputs(3757)) and not (layer0_outputs(313));
    outputs(1294) <= not(layer0_outputs(569));
    outputs(1295) <= (layer0_outputs(3069)) and (layer0_outputs(5844));
    outputs(1296) <= (layer0_outputs(3856)) xor (layer0_outputs(5936));
    outputs(1297) <= not((layer0_outputs(935)) xor (layer0_outputs(6270)));
    outputs(1298) <= (layer0_outputs(43)) xor (layer0_outputs(3308));
    outputs(1299) <= (layer0_outputs(1123)) xor (layer0_outputs(7511));
    outputs(1300) <= (layer0_outputs(5873)) and (layer0_outputs(6667));
    outputs(1301) <= (layer0_outputs(6064)) and not (layer0_outputs(2647));
    outputs(1302) <= (layer0_outputs(3146)) xor (layer0_outputs(4751));
    outputs(1303) <= not((layer0_outputs(7657)) or (layer0_outputs(690)));
    outputs(1304) <= (layer0_outputs(988)) and not (layer0_outputs(1911));
    outputs(1305) <= (layer0_outputs(4539)) xor (layer0_outputs(5337));
    outputs(1306) <= not((layer0_outputs(7123)) or (layer0_outputs(282)));
    outputs(1307) <= (layer0_outputs(3966)) and not (layer0_outputs(7545));
    outputs(1308) <= (layer0_outputs(935)) and (layer0_outputs(2432));
    outputs(1309) <= (layer0_outputs(4782)) and not (layer0_outputs(1060));
    outputs(1310) <= not(layer0_outputs(1977));
    outputs(1311) <= layer0_outputs(5463);
    outputs(1312) <= (layer0_outputs(1370)) xor (layer0_outputs(7490));
    outputs(1313) <= (layer0_outputs(3121)) and not (layer0_outputs(264));
    outputs(1314) <= (layer0_outputs(5695)) and (layer0_outputs(1371));
    outputs(1315) <= not(layer0_outputs(7088));
    outputs(1316) <= not((layer0_outputs(1740)) or (layer0_outputs(7057)));
    outputs(1317) <= (layer0_outputs(103)) and not (layer0_outputs(2060));
    outputs(1318) <= not((layer0_outputs(3393)) xor (layer0_outputs(7239)));
    outputs(1319) <= not((layer0_outputs(3045)) or (layer0_outputs(3082)));
    outputs(1320) <= (layer0_outputs(48)) and not (layer0_outputs(478));
    outputs(1321) <= (layer0_outputs(1145)) xor (layer0_outputs(4571));
    outputs(1322) <= not(layer0_outputs(4021));
    outputs(1323) <= layer0_outputs(2482);
    outputs(1324) <= not((layer0_outputs(2697)) xor (layer0_outputs(4770)));
    outputs(1325) <= not((layer0_outputs(7491)) xor (layer0_outputs(7476)));
    outputs(1326) <= (layer0_outputs(5613)) and not (layer0_outputs(5307));
    outputs(1327) <= not((layer0_outputs(5400)) or (layer0_outputs(6370)));
    outputs(1328) <= not(layer0_outputs(3834));
    outputs(1329) <= (layer0_outputs(3799)) and (layer0_outputs(896));
    outputs(1330) <= (layer0_outputs(7385)) and not (layer0_outputs(3382));
    outputs(1331) <= (layer0_outputs(5841)) and not (layer0_outputs(2808));
    outputs(1332) <= (layer0_outputs(5611)) and (layer0_outputs(5084));
    outputs(1333) <= (layer0_outputs(3422)) and not (layer0_outputs(3481));
    outputs(1334) <= not((layer0_outputs(3866)) or (layer0_outputs(4929)));
    outputs(1335) <= (layer0_outputs(6344)) and not (layer0_outputs(1287));
    outputs(1336) <= layer0_outputs(860);
    outputs(1337) <= (layer0_outputs(3647)) and not (layer0_outputs(4655));
    outputs(1338) <= (layer0_outputs(1783)) and not (layer0_outputs(5581));
    outputs(1339) <= (layer0_outputs(4909)) and not (layer0_outputs(3118));
    outputs(1340) <= not((layer0_outputs(5025)) xor (layer0_outputs(7481)));
    outputs(1341) <= (layer0_outputs(176)) xor (layer0_outputs(2481));
    outputs(1342) <= not((layer0_outputs(3695)) xor (layer0_outputs(4927)));
    outputs(1343) <= not((layer0_outputs(6365)) or (layer0_outputs(5988)));
    outputs(1344) <= (layer0_outputs(2242)) and (layer0_outputs(7634));
    outputs(1345) <= not((layer0_outputs(7456)) or (layer0_outputs(6167)));
    outputs(1346) <= (layer0_outputs(2248)) and not (layer0_outputs(2262));
    outputs(1347) <= (layer0_outputs(4247)) and (layer0_outputs(5690));
    outputs(1348) <= layer0_outputs(4654);
    outputs(1349) <= not((layer0_outputs(6419)) or (layer0_outputs(3480)));
    outputs(1350) <= not(layer0_outputs(7301));
    outputs(1351) <= not((layer0_outputs(396)) or (layer0_outputs(4339)));
    outputs(1352) <= layer0_outputs(49);
    outputs(1353) <= not((layer0_outputs(716)) or (layer0_outputs(4531)));
    outputs(1354) <= (layer0_outputs(7476)) and not (layer0_outputs(3900));
    outputs(1355) <= (layer0_outputs(2536)) and not (layer0_outputs(1928));
    outputs(1356) <= layer0_outputs(2);
    outputs(1357) <= (layer0_outputs(3309)) and not (layer0_outputs(7095));
    outputs(1358) <= layer0_outputs(6490);
    outputs(1359) <= layer0_outputs(648);
    outputs(1360) <= (layer0_outputs(2678)) and not (layer0_outputs(7525));
    outputs(1361) <= not(layer0_outputs(2588));
    outputs(1362) <= layer0_outputs(5158);
    outputs(1363) <= (layer0_outputs(5277)) xor (layer0_outputs(7250));
    outputs(1364) <= (layer0_outputs(2492)) and (layer0_outputs(4248));
    outputs(1365) <= layer0_outputs(2406);
    outputs(1366) <= (layer0_outputs(305)) and (layer0_outputs(886));
    outputs(1367) <= not((layer0_outputs(4342)) or (layer0_outputs(6453)));
    outputs(1368) <= (layer0_outputs(3700)) and not (layer0_outputs(1847));
    outputs(1369) <= (layer0_outputs(2699)) and (layer0_outputs(6911));
    outputs(1370) <= (layer0_outputs(2072)) and (layer0_outputs(5941));
    outputs(1371) <= (layer0_outputs(1826)) and (layer0_outputs(570));
    outputs(1372) <= not((layer0_outputs(4533)) xor (layer0_outputs(365)));
    outputs(1373) <= not(layer0_outputs(2158));
    outputs(1374) <= layer0_outputs(2569);
    outputs(1375) <= not(layer0_outputs(4204));
    outputs(1376) <= not(layer0_outputs(3053));
    outputs(1377) <= layer0_outputs(2519);
    outputs(1378) <= not(layer0_outputs(6213));
    outputs(1379) <= not((layer0_outputs(3317)) xor (layer0_outputs(5796)));
    outputs(1380) <= not((layer0_outputs(1623)) or (layer0_outputs(1055)));
    outputs(1381) <= layer0_outputs(2411);
    outputs(1382) <= layer0_outputs(5479);
    outputs(1383) <= (layer0_outputs(5293)) and not (layer0_outputs(3400));
    outputs(1384) <= (layer0_outputs(6810)) and (layer0_outputs(1955));
    outputs(1385) <= not(layer0_outputs(3693));
    outputs(1386) <= (layer0_outputs(2065)) and not (layer0_outputs(6817));
    outputs(1387) <= not((layer0_outputs(6790)) or (layer0_outputs(2268)));
    outputs(1388) <= (layer0_outputs(2221)) and not (layer0_outputs(2516));
    outputs(1389) <= (layer0_outputs(1242)) and not (layer0_outputs(260));
    outputs(1390) <= (layer0_outputs(7496)) and not (layer0_outputs(541));
    outputs(1391) <= not(layer0_outputs(1017));
    outputs(1392) <= not(layer0_outputs(4776));
    outputs(1393) <= (layer0_outputs(6478)) and not (layer0_outputs(5366));
    outputs(1394) <= not((layer0_outputs(6572)) xor (layer0_outputs(6549)));
    outputs(1395) <= (layer0_outputs(5362)) and not (layer0_outputs(2882));
    outputs(1396) <= not(layer0_outputs(5778));
    outputs(1397) <= (layer0_outputs(4558)) and (layer0_outputs(5100));
    outputs(1398) <= (layer0_outputs(758)) xor (layer0_outputs(4448));
    outputs(1399) <= '0';
    outputs(1400) <= (layer0_outputs(3038)) and not (layer0_outputs(7089));
    outputs(1401) <= (layer0_outputs(826)) xor (layer0_outputs(4084));
    outputs(1402) <= (layer0_outputs(6893)) and not (layer0_outputs(1703));
    outputs(1403) <= (layer0_outputs(372)) and (layer0_outputs(4730));
    outputs(1404) <= (layer0_outputs(946)) and not (layer0_outputs(5735));
    outputs(1405) <= not((layer0_outputs(3313)) or (layer0_outputs(4055)));
    outputs(1406) <= not(layer0_outputs(2559));
    outputs(1407) <= (layer0_outputs(5583)) and not (layer0_outputs(244));
    outputs(1408) <= (layer0_outputs(2572)) and not (layer0_outputs(2190));
    outputs(1409) <= '0';
    outputs(1410) <= (layer0_outputs(2366)) and not (layer0_outputs(5197));
    outputs(1411) <= (layer0_outputs(31)) and not (layer0_outputs(4823));
    outputs(1412) <= (layer0_outputs(4440)) and not (layer0_outputs(5556));
    outputs(1413) <= layer0_outputs(2676);
    outputs(1414) <= not((layer0_outputs(6289)) xor (layer0_outputs(6565)));
    outputs(1415) <= (layer0_outputs(479)) and (layer0_outputs(6417));
    outputs(1416) <= (layer0_outputs(1263)) xor (layer0_outputs(1571));
    outputs(1417) <= (layer0_outputs(1413)) and not (layer0_outputs(5287));
    outputs(1418) <= not((layer0_outputs(7655)) xor (layer0_outputs(5980)));
    outputs(1419) <= (layer0_outputs(2114)) xor (layer0_outputs(5084));
    outputs(1420) <= (layer0_outputs(5015)) and not (layer0_outputs(3790));
    outputs(1421) <= (layer0_outputs(1961)) and not (layer0_outputs(2437));
    outputs(1422) <= (layer0_outputs(1351)) xor (layer0_outputs(1705));
    outputs(1423) <= (layer0_outputs(2314)) and not (layer0_outputs(4446));
    outputs(1424) <= layer0_outputs(4328);
    outputs(1425) <= not((layer0_outputs(4550)) or (layer0_outputs(1283)));
    outputs(1426) <= (layer0_outputs(1213)) and not (layer0_outputs(983));
    outputs(1427) <= (layer0_outputs(828)) and not (layer0_outputs(4120));
    outputs(1428) <= not((layer0_outputs(304)) or (layer0_outputs(6400)));
    outputs(1429) <= not(layer0_outputs(2887)) or (layer0_outputs(3743));
    outputs(1430) <= (layer0_outputs(771)) and not (layer0_outputs(1840));
    outputs(1431) <= (layer0_outputs(1132)) and (layer0_outputs(4501));
    outputs(1432) <= not((layer0_outputs(3524)) xor (layer0_outputs(4150)));
    outputs(1433) <= (layer0_outputs(5385)) and not (layer0_outputs(6275));
    outputs(1434) <= '0';
    outputs(1435) <= layer0_outputs(459);
    outputs(1436) <= not(layer0_outputs(4116));
    outputs(1437) <= not((layer0_outputs(7281)) or (layer0_outputs(3564)));
    outputs(1438) <= (layer0_outputs(3190)) and (layer0_outputs(1221));
    outputs(1439) <= '0';
    outputs(1440) <= (layer0_outputs(675)) and not (layer0_outputs(2922));
    outputs(1441) <= (layer0_outputs(6574)) xor (layer0_outputs(839));
    outputs(1442) <= (layer0_outputs(1657)) and not (layer0_outputs(5642));
    outputs(1443) <= (layer0_outputs(7641)) and (layer0_outputs(3048));
    outputs(1444) <= (layer0_outputs(6803)) and not (layer0_outputs(6047));
    outputs(1445) <= (layer0_outputs(3186)) xor (layer0_outputs(3826));
    outputs(1446) <= not(layer0_outputs(1184));
    outputs(1447) <= (layer0_outputs(3720)) and not (layer0_outputs(2321));
    outputs(1448) <= (layer0_outputs(7646)) xor (layer0_outputs(1451));
    outputs(1449) <= (layer0_outputs(6285)) and (layer0_outputs(4981));
    outputs(1450) <= not(layer0_outputs(2430));
    outputs(1451) <= not((layer0_outputs(4727)) xor (layer0_outputs(5720)));
    outputs(1452) <= not((layer0_outputs(2928)) xor (layer0_outputs(6802)));
    outputs(1453) <= (layer0_outputs(3468)) and (layer0_outputs(6318));
    outputs(1454) <= (layer0_outputs(3792)) and not (layer0_outputs(4883));
    outputs(1455) <= (layer0_outputs(6665)) xor (layer0_outputs(3048));
    outputs(1456) <= (layer0_outputs(269)) and not (layer0_outputs(253));
    outputs(1457) <= '0';
    outputs(1458) <= not((layer0_outputs(4682)) xor (layer0_outputs(5850)));
    outputs(1459) <= (layer0_outputs(6801)) and not (layer0_outputs(2359));
    outputs(1460) <= (layer0_outputs(2938)) and (layer0_outputs(3611));
    outputs(1461) <= (layer0_outputs(1300)) and not (layer0_outputs(5215));
    outputs(1462) <= (layer0_outputs(171)) and not (layer0_outputs(2375));
    outputs(1463) <= (layer0_outputs(3545)) and not (layer0_outputs(3604));
    outputs(1464) <= (layer0_outputs(1000)) and not (layer0_outputs(1327));
    outputs(1465) <= not((layer0_outputs(911)) xor (layer0_outputs(2961)));
    outputs(1466) <= not(layer0_outputs(6397));
    outputs(1467) <= (layer0_outputs(6446)) and not (layer0_outputs(867));
    outputs(1468) <= (layer0_outputs(6144)) and not (layer0_outputs(3781));
    outputs(1469) <= not(layer0_outputs(73));
    outputs(1470) <= (layer0_outputs(4552)) and not (layer0_outputs(4079));
    outputs(1471) <= not((layer0_outputs(1027)) or (layer0_outputs(3809)));
    outputs(1472) <= not(layer0_outputs(2694));
    outputs(1473) <= (layer0_outputs(6857)) and not (layer0_outputs(6136));
    outputs(1474) <= (layer0_outputs(3999)) and (layer0_outputs(6061));
    outputs(1475) <= (layer0_outputs(2597)) and not (layer0_outputs(2131));
    outputs(1476) <= (layer0_outputs(2619)) and not (layer0_outputs(1108));
    outputs(1477) <= (layer0_outputs(5076)) and (layer0_outputs(4458));
    outputs(1478) <= (layer0_outputs(4687)) and (layer0_outputs(6131));
    outputs(1479) <= layer0_outputs(3072);
    outputs(1480) <= not(layer0_outputs(3776));
    outputs(1481) <= (layer0_outputs(5014)) and not (layer0_outputs(2146));
    outputs(1482) <= (layer0_outputs(1641)) and not (layer0_outputs(7523));
    outputs(1483) <= (layer0_outputs(7077)) and not (layer0_outputs(4180));
    outputs(1484) <= not((layer0_outputs(7130)) or (layer0_outputs(1489)));
    outputs(1485) <= not(layer0_outputs(2353));
    outputs(1486) <= (layer0_outputs(4398)) and not (layer0_outputs(4250));
    outputs(1487) <= not((layer0_outputs(1694)) or (layer0_outputs(6672)));
    outputs(1488) <= not(layer0_outputs(4621));
    outputs(1489) <= (layer0_outputs(6629)) and not (layer0_outputs(6381));
    outputs(1490) <= (layer0_outputs(3046)) and not (layer0_outputs(7457));
    outputs(1491) <= (layer0_outputs(3241)) and not (layer0_outputs(3117));
    outputs(1492) <= (layer0_outputs(4648)) and not (layer0_outputs(4810));
    outputs(1493) <= layer0_outputs(4859);
    outputs(1494) <= (layer0_outputs(4059)) and not (layer0_outputs(1998));
    outputs(1495) <= (layer0_outputs(6930)) and not (layer0_outputs(1127));
    outputs(1496) <= not((layer0_outputs(896)) xor (layer0_outputs(4695)));
    outputs(1497) <= (layer0_outputs(5528)) xor (layer0_outputs(1420));
    outputs(1498) <= not((layer0_outputs(6063)) or (layer0_outputs(5542)));
    outputs(1499) <= (layer0_outputs(4426)) and not (layer0_outputs(3946));
    outputs(1500) <= (layer0_outputs(5481)) and (layer0_outputs(7176));
    outputs(1501) <= layer0_outputs(6548);
    outputs(1502) <= (layer0_outputs(3688)) and not (layer0_outputs(1301));
    outputs(1503) <= (layer0_outputs(6782)) and not (layer0_outputs(425));
    outputs(1504) <= (layer0_outputs(3452)) and not (layer0_outputs(7663));
    outputs(1505) <= (layer0_outputs(1876)) and not (layer0_outputs(6248));
    outputs(1506) <= layer0_outputs(1509);
    outputs(1507) <= not((layer0_outputs(4921)) xor (layer0_outputs(653)));
    outputs(1508) <= not(layer0_outputs(1137));
    outputs(1509) <= (layer0_outputs(5458)) and (layer0_outputs(1417));
    outputs(1510) <= (layer0_outputs(2062)) xor (layer0_outputs(137));
    outputs(1511) <= (layer0_outputs(6530)) and (layer0_outputs(7380));
    outputs(1512) <= (layer0_outputs(4557)) and not (layer0_outputs(1694));
    outputs(1513) <= (layer0_outputs(4467)) and not (layer0_outputs(360));
    outputs(1514) <= (layer0_outputs(2133)) and not (layer0_outputs(6763));
    outputs(1515) <= (layer0_outputs(577)) and (layer0_outputs(5462));
    outputs(1516) <= (layer0_outputs(5389)) and not (layer0_outputs(5436));
    outputs(1517) <= not((layer0_outputs(1872)) xor (layer0_outputs(2806)));
    outputs(1518) <= (layer0_outputs(75)) and (layer0_outputs(2512));
    outputs(1519) <= (layer0_outputs(1332)) and (layer0_outputs(7068));
    outputs(1520) <= not((layer0_outputs(189)) or (layer0_outputs(3478)));
    outputs(1521) <= (layer0_outputs(4769)) and not (layer0_outputs(1337));
    outputs(1522) <= not((layer0_outputs(3080)) and (layer0_outputs(6890)));
    outputs(1523) <= (layer0_outputs(4526)) and not (layer0_outputs(6771));
    outputs(1524) <= (layer0_outputs(6849)) and not (layer0_outputs(7052));
    outputs(1525) <= not((layer0_outputs(6435)) or (layer0_outputs(1265)));
    outputs(1526) <= not((layer0_outputs(5566)) xor (layer0_outputs(7557)));
    outputs(1527) <= (layer0_outputs(3213)) and not (layer0_outputs(3845));
    outputs(1528) <= not((layer0_outputs(5002)) or (layer0_outputs(351)));
    outputs(1529) <= not((layer0_outputs(258)) or (layer0_outputs(6119)));
    outputs(1530) <= (layer0_outputs(6363)) or (layer0_outputs(4068));
    outputs(1531) <= not((layer0_outputs(5075)) xor (layer0_outputs(6959)));
    outputs(1532) <= layer0_outputs(1880);
    outputs(1533) <= not(layer0_outputs(2099));
    outputs(1534) <= (layer0_outputs(3907)) and (layer0_outputs(2501));
    outputs(1535) <= (layer0_outputs(2675)) and (layer0_outputs(344));
    outputs(1536) <= not(layer0_outputs(5340));
    outputs(1537) <= (layer0_outputs(4629)) or (layer0_outputs(3570));
    outputs(1538) <= layer0_outputs(3321);
    outputs(1539) <= layer0_outputs(429);
    outputs(1540) <= (layer0_outputs(2364)) xor (layer0_outputs(7541));
    outputs(1541) <= layer0_outputs(6111);
    outputs(1542) <= not((layer0_outputs(7427)) or (layer0_outputs(5683)));
    outputs(1543) <= not(layer0_outputs(1037));
    outputs(1544) <= layer0_outputs(5276);
    outputs(1545) <= (layer0_outputs(5903)) xor (layer0_outputs(6887));
    outputs(1546) <= not(layer0_outputs(506)) or (layer0_outputs(4282));
    outputs(1547) <= layer0_outputs(348);
    outputs(1548) <= not(layer0_outputs(4576));
    outputs(1549) <= not(layer0_outputs(1966));
    outputs(1550) <= not(layer0_outputs(5573));
    outputs(1551) <= not(layer0_outputs(5041)) or (layer0_outputs(362));
    outputs(1552) <= not(layer0_outputs(6852));
    outputs(1553) <= layer0_outputs(3008);
    outputs(1554) <= not(layer0_outputs(4006));
    outputs(1555) <= layer0_outputs(6348);
    outputs(1556) <= not(layer0_outputs(7356)) or (layer0_outputs(3401));
    outputs(1557) <= (layer0_outputs(5474)) and (layer0_outputs(4832));
    outputs(1558) <= (layer0_outputs(5)) or (layer0_outputs(5392));
    outputs(1559) <= (layer0_outputs(6878)) xor (layer0_outputs(3968));
    outputs(1560) <= layer0_outputs(297);
    outputs(1561) <= (layer0_outputs(2401)) and not (layer0_outputs(5488));
    outputs(1562) <= not(layer0_outputs(3614));
    outputs(1563) <= not(layer0_outputs(6897));
    outputs(1564) <= layer0_outputs(1512);
    outputs(1565) <= layer0_outputs(4433);
    outputs(1566) <= (layer0_outputs(6202)) xor (layer0_outputs(5731));
    outputs(1567) <= not(layer0_outputs(5365));
    outputs(1568) <= layer0_outputs(6576);
    outputs(1569) <= layer0_outputs(6641);
    outputs(1570) <= layer0_outputs(5451);
    outputs(1571) <= not(layer0_outputs(740)) or (layer0_outputs(735));
    outputs(1572) <= not(layer0_outputs(3230));
    outputs(1573) <= not((layer0_outputs(1669)) xor (layer0_outputs(4348)));
    outputs(1574) <= not((layer0_outputs(1358)) xor (layer0_outputs(199)));
    outputs(1575) <= not((layer0_outputs(2390)) xor (layer0_outputs(5512)));
    outputs(1576) <= not(layer0_outputs(5759));
    outputs(1577) <= layer0_outputs(366);
    outputs(1578) <= not((layer0_outputs(6253)) xor (layer0_outputs(5273)));
    outputs(1579) <= not(layer0_outputs(5905));
    outputs(1580) <= not((layer0_outputs(560)) and (layer0_outputs(405)));
    outputs(1581) <= layer0_outputs(3587);
    outputs(1582) <= not(layer0_outputs(6776)) or (layer0_outputs(4611));
    outputs(1583) <= not(layer0_outputs(6608));
    outputs(1584) <= layer0_outputs(6753);
    outputs(1585) <= (layer0_outputs(2994)) or (layer0_outputs(4368));
    outputs(1586) <= (layer0_outputs(4671)) and not (layer0_outputs(1979));
    outputs(1587) <= (layer0_outputs(7428)) or (layer0_outputs(3026));
    outputs(1588) <= not((layer0_outputs(1794)) or (layer0_outputs(4990)));
    outputs(1589) <= not(layer0_outputs(5057)) or (layer0_outputs(954));
    outputs(1590) <= layer0_outputs(5436);
    outputs(1591) <= not((layer0_outputs(4127)) xor (layer0_outputs(5198)));
    outputs(1592) <= layer0_outputs(7093);
    outputs(1593) <= layer0_outputs(1670);
    outputs(1594) <= not(layer0_outputs(3268));
    outputs(1595) <= layer0_outputs(6903);
    outputs(1596) <= (layer0_outputs(6071)) or (layer0_outputs(6060));
    outputs(1597) <= (layer0_outputs(1234)) or (layer0_outputs(6107));
    outputs(1598) <= layer0_outputs(4781);
    outputs(1599) <= layer0_outputs(7418);
    outputs(1600) <= layer0_outputs(2974);
    outputs(1601) <= layer0_outputs(7401);
    outputs(1602) <= (layer0_outputs(5802)) and (layer0_outputs(632));
    outputs(1603) <= not((layer0_outputs(6345)) xor (layer0_outputs(5882)));
    outputs(1604) <= layer0_outputs(1150);
    outputs(1605) <= (layer0_outputs(4232)) xor (layer0_outputs(6536));
    outputs(1606) <= layer0_outputs(6060);
    outputs(1607) <= not(layer0_outputs(5716));
    outputs(1608) <= not(layer0_outputs(4340));
    outputs(1609) <= (layer0_outputs(5318)) or (layer0_outputs(7191));
    outputs(1610) <= layer0_outputs(1571);
    outputs(1611) <= (layer0_outputs(3899)) xor (layer0_outputs(3007));
    outputs(1612) <= (layer0_outputs(7107)) and (layer0_outputs(2349));
    outputs(1613) <= not(layer0_outputs(4827)) or (layer0_outputs(5447));
    outputs(1614) <= not(layer0_outputs(2254));
    outputs(1615) <= (layer0_outputs(5773)) and (layer0_outputs(3403));
    outputs(1616) <= layer0_outputs(6502);
    outputs(1617) <= (layer0_outputs(194)) xor (layer0_outputs(6102));
    outputs(1618) <= not(layer0_outputs(68)) or (layer0_outputs(6395));
    outputs(1619) <= (layer0_outputs(1940)) or (layer0_outputs(7448));
    outputs(1620) <= not(layer0_outputs(2170));
    outputs(1621) <= not(layer0_outputs(7108));
    outputs(1622) <= (layer0_outputs(5820)) xor (layer0_outputs(802));
    outputs(1623) <= not((layer0_outputs(415)) xor (layer0_outputs(4673)));
    outputs(1624) <= not(layer0_outputs(3035));
    outputs(1625) <= (layer0_outputs(3982)) or (layer0_outputs(3574));
    outputs(1626) <= layer0_outputs(6156);
    outputs(1627) <= layer0_outputs(6086);
    outputs(1628) <= (layer0_outputs(672)) and not (layer0_outputs(7504));
    outputs(1629) <= not((layer0_outputs(164)) or (layer0_outputs(6916)));
    outputs(1630) <= (layer0_outputs(3882)) xor (layer0_outputs(5006));
    outputs(1631) <= not(layer0_outputs(4953)) or (layer0_outputs(5475));
    outputs(1632) <= not(layer0_outputs(1828));
    outputs(1633) <= layer0_outputs(4610);
    outputs(1634) <= not(layer0_outputs(5456)) or (layer0_outputs(1062));
    outputs(1635) <= not(layer0_outputs(151)) or (layer0_outputs(588));
    outputs(1636) <= layer0_outputs(2049);
    outputs(1637) <= not(layer0_outputs(2037));
    outputs(1638) <= not(layer0_outputs(1511));
    outputs(1639) <= not((layer0_outputs(2435)) and (layer0_outputs(5709)));
    outputs(1640) <= layer0_outputs(2452);
    outputs(1641) <= not(layer0_outputs(5327));
    outputs(1642) <= layer0_outputs(1135);
    outputs(1643) <= (layer0_outputs(5489)) or (layer0_outputs(2903));
    outputs(1644) <= not(layer0_outputs(1948));
    outputs(1645) <= (layer0_outputs(914)) xor (layer0_outputs(7550));
    outputs(1646) <= layer0_outputs(5678);
    outputs(1647) <= layer0_outputs(3055);
    outputs(1648) <= layer0_outputs(4158);
    outputs(1649) <= layer0_outputs(728);
    outputs(1650) <= not(layer0_outputs(5774));
    outputs(1651) <= not(layer0_outputs(1514));
    outputs(1652) <= not(layer0_outputs(5687));
    outputs(1653) <= not(layer0_outputs(156));
    outputs(1654) <= layer0_outputs(1530);
    outputs(1655) <= (layer0_outputs(3729)) xor (layer0_outputs(891));
    outputs(1656) <= not(layer0_outputs(823));
    outputs(1657) <= layer0_outputs(4208);
    outputs(1658) <= not(layer0_outputs(5291)) or (layer0_outputs(6932));
    outputs(1659) <= (layer0_outputs(7209)) and (layer0_outputs(4625));
    outputs(1660) <= not(layer0_outputs(1500)) or (layer0_outputs(3703));
    outputs(1661) <= not((layer0_outputs(3233)) xor (layer0_outputs(1615)));
    outputs(1662) <= not(layer0_outputs(3612));
    outputs(1663) <= layer0_outputs(6848);
    outputs(1664) <= layer0_outputs(3313);
    outputs(1665) <= layer0_outputs(1544);
    outputs(1666) <= (layer0_outputs(466)) or (layer0_outputs(4389));
    outputs(1667) <= not(layer0_outputs(5166)) or (layer0_outputs(7611));
    outputs(1668) <= layer0_outputs(6350);
    outputs(1669) <= not(layer0_outputs(2310)) or (layer0_outputs(4714));
    outputs(1670) <= not(layer0_outputs(4556));
    outputs(1671) <= layer0_outputs(3941);
    outputs(1672) <= layer0_outputs(5407);
    outputs(1673) <= not(layer0_outputs(1655));
    outputs(1674) <= (layer0_outputs(6026)) or (layer0_outputs(5396));
    outputs(1675) <= not((layer0_outputs(4402)) xor (layer0_outputs(2969)));
    outputs(1676) <= not((layer0_outputs(2066)) and (layer0_outputs(7290)));
    outputs(1677) <= not(layer0_outputs(6404)) or (layer0_outputs(1812));
    outputs(1678) <= (layer0_outputs(932)) or (layer0_outputs(7331));
    outputs(1679) <= (layer0_outputs(6056)) xor (layer0_outputs(7145));
    outputs(1680) <= not((layer0_outputs(7054)) xor (layer0_outputs(7646)));
    outputs(1681) <= not((layer0_outputs(320)) or (layer0_outputs(5430)));
    outputs(1682) <= not(layer0_outputs(2008));
    outputs(1683) <= (layer0_outputs(4153)) or (layer0_outputs(562));
    outputs(1684) <= not(layer0_outputs(1374));
    outputs(1685) <= (layer0_outputs(6161)) xor (layer0_outputs(1440));
    outputs(1686) <= not((layer0_outputs(6461)) xor (layer0_outputs(6185)));
    outputs(1687) <= layer0_outputs(2997);
    outputs(1688) <= not((layer0_outputs(946)) and (layer0_outputs(4628)));
    outputs(1689) <= layer0_outputs(5799);
    outputs(1690) <= layer0_outputs(352);
    outputs(1691) <= not(layer0_outputs(3349));
    outputs(1692) <= not(layer0_outputs(4859));
    outputs(1693) <= layer0_outputs(7084);
    outputs(1694) <= not((layer0_outputs(7375)) and (layer0_outputs(1013)));
    outputs(1695) <= not(layer0_outputs(3572));
    outputs(1696) <= not(layer0_outputs(4869)) or (layer0_outputs(5153));
    outputs(1697) <= not(layer0_outputs(682));
    outputs(1698) <= (layer0_outputs(514)) and not (layer0_outputs(389));
    outputs(1699) <= layer0_outputs(6592);
    outputs(1700) <= not(layer0_outputs(3330));
    outputs(1701) <= not(layer0_outputs(7237));
    outputs(1702) <= not(layer0_outputs(7642)) or (layer0_outputs(1812));
    outputs(1703) <= not(layer0_outputs(1400));
    outputs(1704) <= (layer0_outputs(801)) xor (layer0_outputs(4358));
    outputs(1705) <= layer0_outputs(7125);
    outputs(1706) <= (layer0_outputs(5908)) and not (layer0_outputs(5623));
    outputs(1707) <= not(layer0_outputs(2280));
    outputs(1708) <= (layer0_outputs(4469)) or (layer0_outputs(2379));
    outputs(1709) <= not(layer0_outputs(5543));
    outputs(1710) <= not(layer0_outputs(5925));
    outputs(1711) <= not(layer0_outputs(2895));
    outputs(1712) <= layer0_outputs(7348);
    outputs(1713) <= not(layer0_outputs(143));
    outputs(1714) <= not((layer0_outputs(5415)) xor (layer0_outputs(315)));
    outputs(1715) <= not(layer0_outputs(159));
    outputs(1716) <= layer0_outputs(1414);
    outputs(1717) <= (layer0_outputs(7460)) or (layer0_outputs(2714));
    outputs(1718) <= not(layer0_outputs(2921)) or (layer0_outputs(4896));
    outputs(1719) <= layer0_outputs(196);
    outputs(1720) <= (layer0_outputs(973)) or (layer0_outputs(2431));
    outputs(1721) <= not(layer0_outputs(7131));
    outputs(1722) <= not((layer0_outputs(882)) xor (layer0_outputs(4459)));
    outputs(1723) <= not((layer0_outputs(4932)) or (layer0_outputs(4697)));
    outputs(1724) <= layer0_outputs(3029);
    outputs(1725) <= layer0_outputs(7453);
    outputs(1726) <= (layer0_outputs(4774)) and not (layer0_outputs(3469));
    outputs(1727) <= not(layer0_outputs(6997));
    outputs(1728) <= not(layer0_outputs(4272));
    outputs(1729) <= not(layer0_outputs(6881));
    outputs(1730) <= not((layer0_outputs(872)) or (layer0_outputs(1660)));
    outputs(1731) <= not(layer0_outputs(2589));
    outputs(1732) <= not((layer0_outputs(7126)) and (layer0_outputs(4348)));
    outputs(1733) <= layer0_outputs(3160);
    outputs(1734) <= (layer0_outputs(6899)) and not (layer0_outputs(2602));
    outputs(1735) <= not((layer0_outputs(3562)) and (layer0_outputs(5188)));
    outputs(1736) <= not(layer0_outputs(3817));
    outputs(1737) <= layer0_outputs(5962);
    outputs(1738) <= not(layer0_outputs(6895));
    outputs(1739) <= layer0_outputs(1228);
    outputs(1740) <= not((layer0_outputs(5142)) xor (layer0_outputs(2165)));
    outputs(1741) <= not(layer0_outputs(5748));
    outputs(1742) <= not(layer0_outputs(2834));
    outputs(1743) <= layer0_outputs(944);
    outputs(1744) <= (layer0_outputs(218)) xor (layer0_outputs(7038));
    outputs(1745) <= layer0_outputs(3682);
    outputs(1746) <= not(layer0_outputs(2404));
    outputs(1747) <= not((layer0_outputs(2950)) or (layer0_outputs(2890)));
    outputs(1748) <= (layer0_outputs(2268)) xor (layer0_outputs(4578));
    outputs(1749) <= layer0_outputs(7577);
    outputs(1750) <= not(layer0_outputs(4631));
    outputs(1751) <= not(layer0_outputs(7393));
    outputs(1752) <= (layer0_outputs(2453)) or (layer0_outputs(1108));
    outputs(1753) <= (layer0_outputs(3193)) and not (layer0_outputs(6988));
    outputs(1754) <= not(layer0_outputs(7088));
    outputs(1755) <= layer0_outputs(5281);
    outputs(1756) <= not(layer0_outputs(4807));
    outputs(1757) <= (layer0_outputs(2826)) or (layer0_outputs(5149));
    outputs(1758) <= not(layer0_outputs(4993));
    outputs(1759) <= layer0_outputs(3758);
    outputs(1760) <= not(layer0_outputs(6689)) or (layer0_outputs(1581));
    outputs(1761) <= layer0_outputs(1605);
    outputs(1762) <= layer0_outputs(111);
    outputs(1763) <= (layer0_outputs(1913)) or (layer0_outputs(533));
    outputs(1764) <= not(layer0_outputs(4574));
    outputs(1765) <= (layer0_outputs(81)) or (layer0_outputs(3622));
    outputs(1766) <= layer0_outputs(3304);
    outputs(1767) <= (layer0_outputs(3139)) xor (layer0_outputs(4668));
    outputs(1768) <= (layer0_outputs(6086)) and (layer0_outputs(5241));
    outputs(1769) <= (layer0_outputs(4200)) xor (layer0_outputs(4281));
    outputs(1770) <= (layer0_outputs(5330)) and (layer0_outputs(4484));
    outputs(1771) <= not(layer0_outputs(2873)) or (layer0_outputs(3370));
    outputs(1772) <= not(layer0_outputs(3670)) or (layer0_outputs(7034));
    outputs(1773) <= (layer0_outputs(5021)) xor (layer0_outputs(7447));
    outputs(1774) <= not((layer0_outputs(660)) or (layer0_outputs(5361)));
    outputs(1775) <= (layer0_outputs(2327)) and (layer0_outputs(2273));
    outputs(1776) <= layer0_outputs(1097);
    outputs(1777) <= (layer0_outputs(5424)) xor (layer0_outputs(6645));
    outputs(1778) <= layer0_outputs(4683);
    outputs(1779) <= layer0_outputs(4538);
    outputs(1780) <= layer0_outputs(7559);
    outputs(1781) <= (layer0_outputs(5789)) and not (layer0_outputs(4192));
    outputs(1782) <= layer0_outputs(6434);
    outputs(1783) <= not((layer0_outputs(2705)) or (layer0_outputs(2234)));
    outputs(1784) <= layer0_outputs(5829);
    outputs(1785) <= not((layer0_outputs(3261)) xor (layer0_outputs(3460)));
    outputs(1786) <= layer0_outputs(6671);
    outputs(1787) <= not(layer0_outputs(2726));
    outputs(1788) <= not(layer0_outputs(2786));
    outputs(1789) <= not(layer0_outputs(4723)) or (layer0_outputs(528));
    outputs(1790) <= layer0_outputs(7336);
    outputs(1791) <= not(layer0_outputs(2686)) or (layer0_outputs(1139));
    outputs(1792) <= layer0_outputs(6662);
    outputs(1793) <= layer0_outputs(7677);
    outputs(1794) <= not(layer0_outputs(7076)) or (layer0_outputs(1249));
    outputs(1795) <= not((layer0_outputs(4552)) xor (layer0_outputs(7503)));
    outputs(1796) <= layer0_outputs(6449);
    outputs(1797) <= layer0_outputs(520);
    outputs(1798) <= not(layer0_outputs(7529)) or (layer0_outputs(7431));
    outputs(1799) <= not((layer0_outputs(1344)) xor (layer0_outputs(584)));
    outputs(1800) <= not(layer0_outputs(4780));
    outputs(1801) <= not(layer0_outputs(1224));
    outputs(1802) <= layer0_outputs(7450);
    outputs(1803) <= not(layer0_outputs(6533));
    outputs(1804) <= not(layer0_outputs(2222));
    outputs(1805) <= layer0_outputs(2636);
    outputs(1806) <= not((layer0_outputs(7625)) or (layer0_outputs(4238)));
    outputs(1807) <= layer0_outputs(6100);
    outputs(1808) <= not(layer0_outputs(5923));
    outputs(1809) <= layer0_outputs(4632);
    outputs(1810) <= (layer0_outputs(6448)) xor (layer0_outputs(6003));
    outputs(1811) <= not(layer0_outputs(1706));
    outputs(1812) <= not((layer0_outputs(4415)) and (layer0_outputs(287)));
    outputs(1813) <= layer0_outputs(1997);
    outputs(1814) <= (layer0_outputs(1066)) xor (layer0_outputs(3397));
    outputs(1815) <= not(layer0_outputs(5791)) or (layer0_outputs(7116));
    outputs(1816) <= (layer0_outputs(5180)) xor (layer0_outputs(4417));
    outputs(1817) <= not(layer0_outputs(6251));
    outputs(1818) <= layer0_outputs(4803);
    outputs(1819) <= not((layer0_outputs(5362)) xor (layer0_outputs(7532)));
    outputs(1820) <= not((layer0_outputs(6892)) and (layer0_outputs(1314)));
    outputs(1821) <= not(layer0_outputs(1640)) or (layer0_outputs(2252));
    outputs(1822) <= not((layer0_outputs(2828)) xor (layer0_outputs(1539)));
    outputs(1823) <= (layer0_outputs(5541)) xor (layer0_outputs(2367));
    outputs(1824) <= layer0_outputs(4899);
    outputs(1825) <= not(layer0_outputs(7553));
    outputs(1826) <= not(layer0_outputs(5566));
    outputs(1827) <= layer0_outputs(807);
    outputs(1828) <= layer0_outputs(1047);
    outputs(1829) <= (layer0_outputs(3948)) xor (layer0_outputs(7517));
    outputs(1830) <= layer0_outputs(2050);
    outputs(1831) <= (layer0_outputs(7556)) and (layer0_outputs(1194));
    outputs(1832) <= layer0_outputs(5895);
    outputs(1833) <= layer0_outputs(3547);
    outputs(1834) <= layer0_outputs(3773);
    outputs(1835) <= not(layer0_outputs(1930));
    outputs(1836) <= layer0_outputs(4249);
    outputs(1837) <= not(layer0_outputs(4857));
    outputs(1838) <= not((layer0_outputs(7357)) and (layer0_outputs(4045)));
    outputs(1839) <= layer0_outputs(5823);
    outputs(1840) <= not((layer0_outputs(219)) and (layer0_outputs(6117)));
    outputs(1841) <= layer0_outputs(5754);
    outputs(1842) <= not(layer0_outputs(3268)) or (layer0_outputs(7287));
    outputs(1843) <= not(layer0_outputs(1814));
    outputs(1844) <= (layer0_outputs(4880)) and (layer0_outputs(4104));
    outputs(1845) <= not(layer0_outputs(7143)) or (layer0_outputs(4297));
    outputs(1846) <= not(layer0_outputs(2196));
    outputs(1847) <= not(layer0_outputs(4996));
    outputs(1848) <= layer0_outputs(488);
    outputs(1849) <= not(layer0_outputs(3386));
    outputs(1850) <= not(layer0_outputs(3381)) or (layer0_outputs(884));
    outputs(1851) <= not(layer0_outputs(3979));
    outputs(1852) <= not(layer0_outputs(979));
    outputs(1853) <= layer0_outputs(6929);
    outputs(1854) <= not((layer0_outputs(2910)) and (layer0_outputs(3063)));
    outputs(1855) <= not(layer0_outputs(2166));
    outputs(1856) <= not((layer0_outputs(2916)) and (layer0_outputs(4217)));
    outputs(1857) <= layer0_outputs(2587);
    outputs(1858) <= not(layer0_outputs(6184));
    outputs(1859) <= (layer0_outputs(7055)) and (layer0_outputs(1938));
    outputs(1860) <= (layer0_outputs(6081)) and (layer0_outputs(4761));
    outputs(1861) <= not(layer0_outputs(6040));
    outputs(1862) <= not(layer0_outputs(3382)) or (layer0_outputs(7518));
    outputs(1863) <= layer0_outputs(4416);
    outputs(1864) <= (layer0_outputs(2630)) and not (layer0_outputs(6533));
    outputs(1865) <= not(layer0_outputs(6530));
    outputs(1866) <= not(layer0_outputs(3543)) or (layer0_outputs(5605));
    outputs(1867) <= not(layer0_outputs(4591)) or (layer0_outputs(1841));
    outputs(1868) <= not(layer0_outputs(963));
    outputs(1869) <= not((layer0_outputs(810)) or (layer0_outputs(5510)));
    outputs(1870) <= not((layer0_outputs(2712)) xor (layer0_outputs(949)));
    outputs(1871) <= not(layer0_outputs(220)) or (layer0_outputs(2432));
    outputs(1872) <= layer0_outputs(5602);
    outputs(1873) <= not(layer0_outputs(7314));
    outputs(1874) <= (layer0_outputs(273)) or (layer0_outputs(7631));
    outputs(1875) <= not(layer0_outputs(1511)) or (layer0_outputs(2516));
    outputs(1876) <= layer0_outputs(484);
    outputs(1877) <= not(layer0_outputs(4799)) or (layer0_outputs(3368));
    outputs(1878) <= not(layer0_outputs(2044)) or (layer0_outputs(4661));
    outputs(1879) <= not(layer0_outputs(2451));
    outputs(1880) <= layer0_outputs(3045);
    outputs(1881) <= (layer0_outputs(5007)) or (layer0_outputs(5489));
    outputs(1882) <= layer0_outputs(3030);
    outputs(1883) <= not(layer0_outputs(5879));
    outputs(1884) <= layer0_outputs(3227);
    outputs(1885) <= (layer0_outputs(4310)) xor (layer0_outputs(7216));
    outputs(1886) <= not(layer0_outputs(4271));
    outputs(1887) <= not(layer0_outputs(5978));
    outputs(1888) <= layer0_outputs(1865);
    outputs(1889) <= (layer0_outputs(395)) or (layer0_outputs(1483));
    outputs(1890) <= layer0_outputs(7064);
    outputs(1891) <= layer0_outputs(4681);
    outputs(1892) <= not((layer0_outputs(2230)) and (layer0_outputs(5780)));
    outputs(1893) <= layer0_outputs(3540);
    outputs(1894) <= (layer0_outputs(4802)) and (layer0_outputs(323));
    outputs(1895) <= not((layer0_outputs(6443)) and (layer0_outputs(5161)));
    outputs(1896) <= not(layer0_outputs(3315));
    outputs(1897) <= (layer0_outputs(2304)) and (layer0_outputs(3553));
    outputs(1898) <= not(layer0_outputs(5965));
    outputs(1899) <= not(layer0_outputs(6689)) or (layer0_outputs(5286));
    outputs(1900) <= not((layer0_outputs(3245)) and (layer0_outputs(128)));
    outputs(1901) <= not(layer0_outputs(4826));
    outputs(1902) <= not((layer0_outputs(2920)) or (layer0_outputs(665)));
    outputs(1903) <= (layer0_outputs(6845)) xor (layer0_outputs(1677));
    outputs(1904) <= layer0_outputs(2976);
    outputs(1905) <= layer0_outputs(1927);
    outputs(1906) <= (layer0_outputs(6885)) or (layer0_outputs(105));
    outputs(1907) <= layer0_outputs(3109);
    outputs(1908) <= layer0_outputs(2248);
    outputs(1909) <= layer0_outputs(978);
    outputs(1910) <= layer0_outputs(6306);
    outputs(1911) <= not((layer0_outputs(5531)) xor (layer0_outputs(4805)));
    outputs(1912) <= layer0_outputs(2772);
    outputs(1913) <= layer0_outputs(3087);
    outputs(1914) <= not(layer0_outputs(4798));
    outputs(1915) <= not(layer0_outputs(2933));
    outputs(1916) <= not(layer0_outputs(2051));
    outputs(1917) <= layer0_outputs(455);
    outputs(1918) <= (layer0_outputs(5250)) xor (layer0_outputs(6666));
    outputs(1919) <= not((layer0_outputs(2139)) xor (layer0_outputs(367)));
    outputs(1920) <= not(layer0_outputs(4912));
    outputs(1921) <= not((layer0_outputs(7137)) or (layer0_outputs(7047)));
    outputs(1922) <= not((layer0_outputs(367)) xor (layer0_outputs(3405)));
    outputs(1923) <= (layer0_outputs(7413)) xor (layer0_outputs(1284));
    outputs(1924) <= not(layer0_outputs(3849));
    outputs(1925) <= not((layer0_outputs(3937)) xor (layer0_outputs(6670)));
    outputs(1926) <= (layer0_outputs(1063)) and not (layer0_outputs(2527));
    outputs(1927) <= layer0_outputs(1721);
    outputs(1928) <= layer0_outputs(4580);
    outputs(1929) <= layer0_outputs(6252);
    outputs(1930) <= not((layer0_outputs(3130)) and (layer0_outputs(7091)));
    outputs(1931) <= layer0_outputs(7323);
    outputs(1932) <= not(layer0_outputs(5162));
    outputs(1933) <= not(layer0_outputs(7616));
    outputs(1934) <= layer0_outputs(6622);
    outputs(1935) <= not(layer0_outputs(2418));
    outputs(1936) <= not(layer0_outputs(7479));
    outputs(1937) <= layer0_outputs(5244);
    outputs(1938) <= layer0_outputs(3251);
    outputs(1939) <= not(layer0_outputs(4464));
    outputs(1940) <= (layer0_outputs(1538)) and not (layer0_outputs(6707));
    outputs(1941) <= not(layer0_outputs(44));
    outputs(1942) <= not(layer0_outputs(6905)) or (layer0_outputs(1847));
    outputs(1943) <= not(layer0_outputs(2201));
    outputs(1944) <= not((layer0_outputs(6082)) xor (layer0_outputs(4964)));
    outputs(1945) <= not(layer0_outputs(1570));
    outputs(1946) <= (layer0_outputs(4852)) and (layer0_outputs(1792));
    outputs(1947) <= not(layer0_outputs(1266)) or (layer0_outputs(6970));
    outputs(1948) <= not((layer0_outputs(301)) or (layer0_outputs(795)));
    outputs(1949) <= not(layer0_outputs(2442));
    outputs(1950) <= layer0_outputs(1795);
    outputs(1951) <= (layer0_outputs(7322)) and not (layer0_outputs(1514));
    outputs(1952) <= layer0_outputs(6346);
    outputs(1953) <= not(layer0_outputs(4827)) or (layer0_outputs(4492));
    outputs(1954) <= not(layer0_outputs(4144)) or (layer0_outputs(1007));
    outputs(1955) <= (layer0_outputs(5798)) and (layer0_outputs(4205));
    outputs(1956) <= not(layer0_outputs(7181));
    outputs(1957) <= layer0_outputs(803);
    outputs(1958) <= not(layer0_outputs(137)) or (layer0_outputs(6842));
    outputs(1959) <= not(layer0_outputs(2087));
    outputs(1960) <= layer0_outputs(3921);
    outputs(1961) <= not(layer0_outputs(1158));
    outputs(1962) <= layer0_outputs(4146);
    outputs(1963) <= not((layer0_outputs(1030)) or (layer0_outputs(3594)));
    outputs(1964) <= not(layer0_outputs(6161));
    outputs(1965) <= not((layer0_outputs(5477)) and (layer0_outputs(941)));
    outputs(1966) <= not((layer0_outputs(5263)) or (layer0_outputs(359)));
    outputs(1967) <= layer0_outputs(2405);
    outputs(1968) <= layer0_outputs(6246);
    outputs(1969) <= layer0_outputs(2813);
    outputs(1970) <= not(layer0_outputs(3864));
    outputs(1971) <= layer0_outputs(3642);
    outputs(1972) <= (layer0_outputs(4465)) and not (layer0_outputs(213));
    outputs(1973) <= (layer0_outputs(6466)) xor (layer0_outputs(7248));
    outputs(1974) <= (layer0_outputs(285)) xor (layer0_outputs(1808));
    outputs(1975) <= (layer0_outputs(22)) xor (layer0_outputs(7261));
    outputs(1976) <= not((layer0_outputs(1310)) and (layer0_outputs(6405)));
    outputs(1977) <= not(layer0_outputs(2079));
    outputs(1978) <= not(layer0_outputs(1257)) or (layer0_outputs(3303));
    outputs(1979) <= not(layer0_outputs(4722)) or (layer0_outputs(3270));
    outputs(1980) <= not(layer0_outputs(3202));
    outputs(1981) <= (layer0_outputs(4067)) and not (layer0_outputs(1460));
    outputs(1982) <= not(layer0_outputs(6356));
    outputs(1983) <= layer0_outputs(2730);
    outputs(1984) <= not(layer0_outputs(2200));
    outputs(1985) <= layer0_outputs(462);
    outputs(1986) <= (layer0_outputs(188)) and (layer0_outputs(1120));
    outputs(1987) <= not((layer0_outputs(6288)) xor (layer0_outputs(2778)));
    outputs(1988) <= not(layer0_outputs(2293));
    outputs(1989) <= not(layer0_outputs(1827));
    outputs(1990) <= not((layer0_outputs(5543)) or (layer0_outputs(6076)));
    outputs(1991) <= layer0_outputs(3376);
    outputs(1992) <= layer0_outputs(2359);
    outputs(1993) <= layer0_outputs(1805);
    outputs(1994) <= layer0_outputs(4280);
    outputs(1995) <= not(layer0_outputs(4131));
    outputs(1996) <= not(layer0_outputs(2048));
    outputs(1997) <= layer0_outputs(6701);
    outputs(1998) <= not(layer0_outputs(4117));
    outputs(1999) <= not(layer0_outputs(2592));
    outputs(2000) <= (layer0_outputs(5724)) xor (layer0_outputs(3171));
    outputs(2001) <= not(layer0_outputs(590));
    outputs(2002) <= (layer0_outputs(3033)) or (layer0_outputs(1276));
    outputs(2003) <= not(layer0_outputs(660));
    outputs(2004) <= not(layer0_outputs(2853)) or (layer0_outputs(1985));
    outputs(2005) <= layer0_outputs(6602);
    outputs(2006) <= not(layer0_outputs(3542));
    outputs(2007) <= (layer0_outputs(1753)) and (layer0_outputs(3412));
    outputs(2008) <= not((layer0_outputs(2088)) xor (layer0_outputs(6607)));
    outputs(2009) <= not(layer0_outputs(1547)) or (layer0_outputs(585));
    outputs(2010) <= layer0_outputs(5998);
    outputs(2011) <= not(layer0_outputs(1487));
    outputs(2012) <= not((layer0_outputs(2022)) and (layer0_outputs(2442)));
    outputs(2013) <= not(layer0_outputs(5852));
    outputs(2014) <= (layer0_outputs(1628)) xor (layer0_outputs(4096));
    outputs(2015) <= (layer0_outputs(6711)) and not (layer0_outputs(6236));
    outputs(2016) <= not(layer0_outputs(6115));
    outputs(2017) <= not(layer0_outputs(3390)) or (layer0_outputs(5308));
    outputs(2018) <= not((layer0_outputs(7211)) and (layer0_outputs(4399)));
    outputs(2019) <= layer0_outputs(2129);
    outputs(2020) <= not((layer0_outputs(6952)) xor (layer0_outputs(5604)));
    outputs(2021) <= not(layer0_outputs(132));
    outputs(2022) <= not(layer0_outputs(63)) or (layer0_outputs(952));
    outputs(2023) <= not(layer0_outputs(460));
    outputs(2024) <= not(layer0_outputs(2786));
    outputs(2025) <= not(layer0_outputs(5510));
    outputs(2026) <= not(layer0_outputs(2267));
    outputs(2027) <= not(layer0_outputs(6187));
    outputs(2028) <= not(layer0_outputs(6109)) or (layer0_outputs(3326));
    outputs(2029) <= not((layer0_outputs(6450)) or (layer0_outputs(4798)));
    outputs(2030) <= layer0_outputs(4320);
    outputs(2031) <= layer0_outputs(517);
    outputs(2032) <= layer0_outputs(5019);
    outputs(2033) <= (layer0_outputs(2225)) xor (layer0_outputs(3779));
    outputs(2034) <= not((layer0_outputs(3103)) and (layer0_outputs(289)));
    outputs(2035) <= layer0_outputs(116);
    outputs(2036) <= not((layer0_outputs(5488)) xor (layer0_outputs(2867)));
    outputs(2037) <= not(layer0_outputs(1903)) or (layer0_outputs(7448));
    outputs(2038) <= layer0_outputs(892);
    outputs(2039) <= layer0_outputs(6619);
    outputs(2040) <= not((layer0_outputs(4293)) xor (layer0_outputs(6250)));
    outputs(2041) <= layer0_outputs(1597);
    outputs(2042) <= layer0_outputs(4511);
    outputs(2043) <= not(layer0_outputs(2131));
    outputs(2044) <= (layer0_outputs(4276)) xor (layer0_outputs(7614));
    outputs(2045) <= layer0_outputs(7049);
    outputs(2046) <= layer0_outputs(1148);
    outputs(2047) <= not(layer0_outputs(5484));
    outputs(2048) <= not((layer0_outputs(4627)) xor (layer0_outputs(4154)));
    outputs(2049) <= not(layer0_outputs(2560));
    outputs(2050) <= (layer0_outputs(3260)) or (layer0_outputs(609));
    outputs(2051) <= not((layer0_outputs(3504)) and (layer0_outputs(7560)));
    outputs(2052) <= not((layer0_outputs(7317)) xor (layer0_outputs(2846)));
    outputs(2053) <= not((layer0_outputs(606)) or (layer0_outputs(1444)));
    outputs(2054) <= layer0_outputs(6620);
    outputs(2055) <= not(layer0_outputs(2444));
    outputs(2056) <= (layer0_outputs(2563)) and not (layer0_outputs(2067));
    outputs(2057) <= not((layer0_outputs(1593)) xor (layer0_outputs(6650)));
    outputs(2058) <= not(layer0_outputs(5453)) or (layer0_outputs(1577));
    outputs(2059) <= not((layer0_outputs(4597)) and (layer0_outputs(39)));
    outputs(2060) <= layer0_outputs(3921);
    outputs(2061) <= not(layer0_outputs(677));
    outputs(2062) <= (layer0_outputs(717)) and not (layer0_outputs(3421));
    outputs(2063) <= (layer0_outputs(1683)) and (layer0_outputs(4995));
    outputs(2064) <= layer0_outputs(1202);
    outputs(2065) <= not(layer0_outputs(3315));
    outputs(2066) <= not(layer0_outputs(1854));
    outputs(2067) <= not(layer0_outputs(7516)) or (layer0_outputs(2401));
    outputs(2068) <= not(layer0_outputs(3536));
    outputs(2069) <= not((layer0_outputs(5635)) and (layer0_outputs(5727)));
    outputs(2070) <= (layer0_outputs(5087)) and (layer0_outputs(5216));
    outputs(2071) <= not(layer0_outputs(1064));
    outputs(2072) <= (layer0_outputs(6889)) and not (layer0_outputs(711));
    outputs(2073) <= layer0_outputs(3079);
    outputs(2074) <= not(layer0_outputs(446));
    outputs(2075) <= not(layer0_outputs(2731)) or (layer0_outputs(2295));
    outputs(2076) <= not(layer0_outputs(6912));
    outputs(2077) <= not(layer0_outputs(4598));
    outputs(2078) <= not(layer0_outputs(7585)) or (layer0_outputs(6015));
    outputs(2079) <= layer0_outputs(2020);
    outputs(2080) <= (layer0_outputs(5031)) xor (layer0_outputs(6451));
    outputs(2081) <= not((layer0_outputs(6744)) and (layer0_outputs(1273)));
    outputs(2082) <= not(layer0_outputs(2745));
    outputs(2083) <= not(layer0_outputs(5833)) or (layer0_outputs(1562));
    outputs(2084) <= (layer0_outputs(491)) and not (layer0_outputs(1837));
    outputs(2085) <= layer0_outputs(4056);
    outputs(2086) <= layer0_outputs(2013);
    outputs(2087) <= not(layer0_outputs(7268));
    outputs(2088) <= layer0_outputs(7195);
    outputs(2089) <= not(layer0_outputs(5350));
    outputs(2090) <= not(layer0_outputs(1592));
    outputs(2091) <= not(layer0_outputs(5842));
    outputs(2092) <= not(layer0_outputs(2053));
    outputs(2093) <= layer0_outputs(6300);
    outputs(2094) <= layer0_outputs(6021);
    outputs(2095) <= layer0_outputs(5444);
    outputs(2096) <= not(layer0_outputs(7184));
    outputs(2097) <= layer0_outputs(6648);
    outputs(2098) <= (layer0_outputs(5705)) xor (layer0_outputs(5150));
    outputs(2099) <= layer0_outputs(5651);
    outputs(2100) <= not(layer0_outputs(4314));
    outputs(2101) <= layer0_outputs(6876);
    outputs(2102) <= layer0_outputs(4659);
    outputs(2103) <= not((layer0_outputs(555)) xor (layer0_outputs(3671)));
    outputs(2104) <= not(layer0_outputs(4626)) or (layer0_outputs(4778));
    outputs(2105) <= layer0_outputs(3540);
    outputs(2106) <= not(layer0_outputs(922));
    outputs(2107) <= not(layer0_outputs(7638));
    outputs(2108) <= not(layer0_outputs(6170));
    outputs(2109) <= not((layer0_outputs(237)) xor (layer0_outputs(5045)));
    outputs(2110) <= not(layer0_outputs(5578)) or (layer0_outputs(5309));
    outputs(2111) <= not(layer0_outputs(1687));
    outputs(2112) <= layer0_outputs(2590);
    outputs(2113) <= layer0_outputs(3417);
    outputs(2114) <= layer0_outputs(3333);
    outputs(2115) <= not(layer0_outputs(4545)) or (layer0_outputs(1416));
    outputs(2116) <= not((layer0_outputs(4378)) or (layer0_outputs(4027)));
    outputs(2117) <= (layer0_outputs(5904)) xor (layer0_outputs(4446));
    outputs(2118) <= (layer0_outputs(1273)) xor (layer0_outputs(4910));
    outputs(2119) <= layer0_outputs(5462);
    outputs(2120) <= not(layer0_outputs(4531));
    outputs(2121) <= not((layer0_outputs(205)) xor (layer0_outputs(526)));
    outputs(2122) <= layer0_outputs(1353);
    outputs(2123) <= not(layer0_outputs(6688));
    outputs(2124) <= layer0_outputs(1148);
    outputs(2125) <= not(layer0_outputs(7310));
    outputs(2126) <= (layer0_outputs(2036)) and (layer0_outputs(3450));
    outputs(2127) <= layer0_outputs(1000);
    outputs(2128) <= not(layer0_outputs(3699)) or (layer0_outputs(1336));
    outputs(2129) <= layer0_outputs(6649);
    outputs(2130) <= not(layer0_outputs(949)) or (layer0_outputs(6599));
    outputs(2131) <= layer0_outputs(414);
    outputs(2132) <= (layer0_outputs(3760)) and not (layer0_outputs(6825));
    outputs(2133) <= not(layer0_outputs(6479)) or (layer0_outputs(7610));
    outputs(2134) <= layer0_outputs(2780);
    outputs(2135) <= not(layer0_outputs(4870));
    outputs(2136) <= not(layer0_outputs(3503)) or (layer0_outputs(2724));
    outputs(2137) <= layer0_outputs(3784);
    outputs(2138) <= not(layer0_outputs(1142)) or (layer0_outputs(3873));
    outputs(2139) <= layer0_outputs(1804);
    outputs(2140) <= not(layer0_outputs(7095));
    outputs(2141) <= not(layer0_outputs(3663));
    outputs(2142) <= not(layer0_outputs(7393));
    outputs(2143) <= layer0_outputs(746);
    outputs(2144) <= not(layer0_outputs(1401));
    outputs(2145) <= layer0_outputs(7239);
    outputs(2146) <= (layer0_outputs(4685)) and not (layer0_outputs(1884));
    outputs(2147) <= (layer0_outputs(1818)) and not (layer0_outputs(6342));
    outputs(2148) <= (layer0_outputs(1588)) or (layer0_outputs(2644));
    outputs(2149) <= (layer0_outputs(7365)) and not (layer0_outputs(7245));
    outputs(2150) <= layer0_outputs(6374);
    outputs(2151) <= not(layer0_outputs(5446));
    outputs(2152) <= not(layer0_outputs(5329));
    outputs(2153) <= not((layer0_outputs(692)) xor (layer0_outputs(6492)));
    outputs(2154) <= not(layer0_outputs(921)) or (layer0_outputs(3926));
    outputs(2155) <= not(layer0_outputs(1488));
    outputs(2156) <= layer0_outputs(5253);
    outputs(2157) <= not((layer0_outputs(251)) xor (layer0_outputs(6056)));
    outputs(2158) <= not((layer0_outputs(1923)) xor (layer0_outputs(3196)));
    outputs(2159) <= (layer0_outputs(3143)) xor (layer0_outputs(5096));
    outputs(2160) <= not(layer0_outputs(3969)) or (layer0_outputs(4299));
    outputs(2161) <= not((layer0_outputs(4656)) xor (layer0_outputs(644)));
    outputs(2162) <= not(layer0_outputs(2488)) or (layer0_outputs(893));
    outputs(2163) <= layer0_outputs(2861);
    outputs(2164) <= (layer0_outputs(1269)) and not (layer0_outputs(393));
    outputs(2165) <= not(layer0_outputs(6727));
    outputs(2166) <= layer0_outputs(5138);
    outputs(2167) <= layer0_outputs(815);
    outputs(2168) <= layer0_outputs(4708);
    outputs(2169) <= not(layer0_outputs(6272)) or (layer0_outputs(146));
    outputs(2170) <= not(layer0_outputs(302)) or (layer0_outputs(1181));
    outputs(2171) <= (layer0_outputs(7487)) and not (layer0_outputs(1719));
    outputs(2172) <= (layer0_outputs(2367)) or (layer0_outputs(1516));
    outputs(2173) <= not((layer0_outputs(4950)) xor (layer0_outputs(6360)));
    outputs(2174) <= (layer0_outputs(7249)) and not (layer0_outputs(5230));
    outputs(2175) <= (layer0_outputs(207)) or (layer0_outputs(3777));
    outputs(2176) <= not(layer0_outputs(1121)) or (layer0_outputs(6594));
    outputs(2177) <= (layer0_outputs(4894)) or (layer0_outputs(3899));
    outputs(2178) <= layer0_outputs(5665);
    outputs(2179) <= not((layer0_outputs(5128)) and (layer0_outputs(2372)));
    outputs(2180) <= not(layer0_outputs(4425)) or (layer0_outputs(7559));
    outputs(2181) <= (layer0_outputs(4432)) and not (layer0_outputs(6138));
    outputs(2182) <= not(layer0_outputs(614));
    outputs(2183) <= not((layer0_outputs(2051)) or (layer0_outputs(3336)));
    outputs(2184) <= not(layer0_outputs(485));
    outputs(2185) <= not(layer0_outputs(1768)) or (layer0_outputs(482));
    outputs(2186) <= not(layer0_outputs(7459)) or (layer0_outputs(1442));
    outputs(2187) <= not(layer0_outputs(1796));
    outputs(2188) <= not(layer0_outputs(165));
    outputs(2189) <= not((layer0_outputs(2674)) and (layer0_outputs(719)));
    outputs(2190) <= not(layer0_outputs(72)) or (layer0_outputs(4620));
    outputs(2191) <= not(layer0_outputs(3829));
    outputs(2192) <= layer0_outputs(1001);
    outputs(2193) <= not(layer0_outputs(4043));
    outputs(2194) <= (layer0_outputs(1318)) and (layer0_outputs(7678));
    outputs(2195) <= '1';
    outputs(2196) <= not(layer0_outputs(2660));
    outputs(2197) <= not((layer0_outputs(6935)) and (layer0_outputs(3854)));
    outputs(2198) <= not((layer0_outputs(5295)) and (layer0_outputs(4617)));
    outputs(2199) <= layer0_outputs(7482);
    outputs(2200) <= not(layer0_outputs(5975));
    outputs(2201) <= not(layer0_outputs(2684));
    outputs(2202) <= not(layer0_outputs(583)) or (layer0_outputs(2754));
    outputs(2203) <= not((layer0_outputs(1293)) xor (layer0_outputs(1784)));
    outputs(2204) <= not(layer0_outputs(11)) or (layer0_outputs(3074));
    outputs(2205) <= not(layer0_outputs(4108));
    outputs(2206) <= not(layer0_outputs(5166));
    outputs(2207) <= layer0_outputs(919);
    outputs(2208) <= not((layer0_outputs(7127)) xor (layer0_outputs(5555)));
    outputs(2209) <= not((layer0_outputs(850)) or (layer0_outputs(1986)));
    outputs(2210) <= not(layer0_outputs(1782)) or (layer0_outputs(4465));
    outputs(2211) <= not(layer0_outputs(2236));
    outputs(2212) <= layer0_outputs(4503);
    outputs(2213) <= layer0_outputs(6174);
    outputs(2214) <= not(layer0_outputs(6285)) or (layer0_outputs(343));
    outputs(2215) <= not((layer0_outputs(5948)) and (layer0_outputs(1480)));
    outputs(2216) <= (layer0_outputs(5020)) xor (layer0_outputs(5836));
    outputs(2217) <= (layer0_outputs(1778)) or (layer0_outputs(2307));
    outputs(2218) <= not(layer0_outputs(5534));
    outputs(2219) <= (layer0_outputs(6271)) and (layer0_outputs(5969));
    outputs(2220) <= layer0_outputs(2023);
    outputs(2221) <= not(layer0_outputs(2789)) or (layer0_outputs(1264));
    outputs(2222) <= (layer0_outputs(3813)) xor (layer0_outputs(5372));
    outputs(2223) <= layer0_outputs(7011);
    outputs(2224) <= not(layer0_outputs(2574)) or (layer0_outputs(1793));
    outputs(2225) <= layer0_outputs(7527);
    outputs(2226) <= layer0_outputs(741);
    outputs(2227) <= (layer0_outputs(6095)) xor (layer0_outputs(7211));
    outputs(2228) <= layer0_outputs(5062);
    outputs(2229) <= (layer0_outputs(2881)) and not (layer0_outputs(4772));
    outputs(2230) <= (layer0_outputs(1540)) xor (layer0_outputs(1280));
    outputs(2231) <= layer0_outputs(5086);
    outputs(2232) <= not((layer0_outputs(6244)) and (layer0_outputs(5261)));
    outputs(2233) <= (layer0_outputs(1527)) and not (layer0_outputs(5577));
    outputs(2234) <= (layer0_outputs(286)) or (layer0_outputs(1841));
    outputs(2235) <= not(layer0_outputs(432)) or (layer0_outputs(3992));
    outputs(2236) <= not(layer0_outputs(1274)) or (layer0_outputs(3024));
    outputs(2237) <= not(layer0_outputs(2438)) or (layer0_outputs(3988));
    outputs(2238) <= not(layer0_outputs(7308)) or (layer0_outputs(6908));
    outputs(2239) <= not(layer0_outputs(4186));
    outputs(2240) <= layer0_outputs(638);
    outputs(2241) <= not(layer0_outputs(3442));
    outputs(2242) <= layer0_outputs(6388);
    outputs(2243) <= (layer0_outputs(297)) and not (layer0_outputs(5860));
    outputs(2244) <= (layer0_outputs(7413)) and not (layer0_outputs(4073));
    outputs(2245) <= not((layer0_outputs(4801)) or (layer0_outputs(5323)));
    outputs(2246) <= (layer0_outputs(3088)) xor (layer0_outputs(5269));
    outputs(2247) <= layer0_outputs(4824);
    outputs(2248) <= not(layer0_outputs(4316)) or (layer0_outputs(579));
    outputs(2249) <= not(layer0_outputs(2532));
    outputs(2250) <= layer0_outputs(402);
    outputs(2251) <= (layer0_outputs(2288)) and (layer0_outputs(4555));
    outputs(2252) <= (layer0_outputs(464)) and not (layer0_outputs(3690));
    outputs(2253) <= layer0_outputs(3247);
    outputs(2254) <= not((layer0_outputs(1999)) xor (layer0_outputs(926)));
    outputs(2255) <= layer0_outputs(1658);
    outputs(2256) <= not((layer0_outputs(1988)) xor (layer0_outputs(3632)));
    outputs(2257) <= not(layer0_outputs(4975));
    outputs(2258) <= not(layer0_outputs(1044));
    outputs(2259) <= layer0_outputs(3238);
    outputs(2260) <= (layer0_outputs(6306)) and not (layer0_outputs(4911));
    outputs(2261) <= not(layer0_outputs(1005));
    outputs(2262) <= not((layer0_outputs(2118)) xor (layer0_outputs(750)));
    outputs(2263) <= not(layer0_outputs(6397));
    outputs(2264) <= layer0_outputs(5725);
    outputs(2265) <= not((layer0_outputs(7605)) xor (layer0_outputs(6861)));
    outputs(2266) <= (layer0_outputs(7383)) or (layer0_outputs(4062));
    outputs(2267) <= not(layer0_outputs(1669));
    outputs(2268) <= layer0_outputs(3229);
    outputs(2269) <= layer0_outputs(3454);
    outputs(2270) <= '1';
    outputs(2271) <= layer0_outputs(671);
    outputs(2272) <= not(layer0_outputs(6191)) or (layer0_outputs(1230));
    outputs(2273) <= not(layer0_outputs(4626));
    outputs(2274) <= (layer0_outputs(632)) xor (layer0_outputs(1917));
    outputs(2275) <= not(layer0_outputs(7508));
    outputs(2276) <= not((layer0_outputs(2308)) xor (layer0_outputs(5347)));
    outputs(2277) <= not(layer0_outputs(968)) or (layer0_outputs(4106));
    outputs(2278) <= not(layer0_outputs(1479)) or (layer0_outputs(6641));
    outputs(2279) <= layer0_outputs(2073);
    outputs(2280) <= layer0_outputs(5649);
    outputs(2281) <= not(layer0_outputs(2940)) or (layer0_outputs(1264));
    outputs(2282) <= not(layer0_outputs(2545)) or (layer0_outputs(5907));
    outputs(2283) <= not(layer0_outputs(780));
    outputs(2284) <= not(layer0_outputs(5657)) or (layer0_outputs(51));
    outputs(2285) <= layer0_outputs(5846);
    outputs(2286) <= not(layer0_outputs(3816));
    outputs(2287) <= not((layer0_outputs(6799)) or (layer0_outputs(3250)));
    outputs(2288) <= not((layer0_outputs(6749)) xor (layer0_outputs(2728)));
    outputs(2289) <= (layer0_outputs(7175)) or (layer0_outputs(2605));
    outputs(2290) <= not(layer0_outputs(1713));
    outputs(2291) <= not(layer0_outputs(2085));
    outputs(2292) <= not((layer0_outputs(5137)) and (layer0_outputs(5911)));
    outputs(2293) <= (layer0_outputs(3945)) and not (layer0_outputs(5965));
    outputs(2294) <= not(layer0_outputs(5900));
    outputs(2295) <= (layer0_outputs(7231)) and not (layer0_outputs(3774));
    outputs(2296) <= (layer0_outputs(1396)) or (layer0_outputs(6615));
    outputs(2297) <= (layer0_outputs(318)) and not (layer0_outputs(2451));
    outputs(2298) <= not(layer0_outputs(1149));
    outputs(2299) <= not((layer0_outputs(2249)) xor (layer0_outputs(6559)));
    outputs(2300) <= not(layer0_outputs(5022));
    outputs(2301) <= (layer0_outputs(4194)) or (layer0_outputs(2826));
    outputs(2302) <= not(layer0_outputs(4886)) or (layer0_outputs(1726));
    outputs(2303) <= layer0_outputs(2919);
    outputs(2304) <= not(layer0_outputs(7085)) or (layer0_outputs(4387));
    outputs(2305) <= layer0_outputs(3933);
    outputs(2306) <= not(layer0_outputs(1102));
    outputs(2307) <= not((layer0_outputs(2856)) or (layer0_outputs(1459)));
    outputs(2308) <= not((layer0_outputs(3845)) xor (layer0_outputs(600)));
    outputs(2309) <= not(layer0_outputs(3978));
    outputs(2310) <= not(layer0_outputs(7157)) or (layer0_outputs(7520));
    outputs(2311) <= layer0_outputs(3925);
    outputs(2312) <= (layer0_outputs(2551)) and not (layer0_outputs(3833));
    outputs(2313) <= not((layer0_outputs(5952)) or (layer0_outputs(6411)));
    outputs(2314) <= (layer0_outputs(3607)) xor (layer0_outputs(3147));
    outputs(2315) <= not(layer0_outputs(4247));
    outputs(2316) <= (layer0_outputs(6239)) xor (layer0_outputs(6516));
    outputs(2317) <= not(layer0_outputs(2917));
    outputs(2318) <= layer0_outputs(3890);
    outputs(2319) <= not(layer0_outputs(3474));
    outputs(2320) <= layer0_outputs(4318);
    outputs(2321) <= (layer0_outputs(6375)) and not (layer0_outputs(2151));
    outputs(2322) <= not(layer0_outputs(3255));
    outputs(2323) <= not(layer0_outputs(846)) or (layer0_outputs(5320));
    outputs(2324) <= not(layer0_outputs(1856));
    outputs(2325) <= (layer0_outputs(7601)) and (layer0_outputs(7530));
    outputs(2326) <= not(layer0_outputs(4294));
    outputs(2327) <= not(layer0_outputs(7345));
    outputs(2328) <= (layer0_outputs(6880)) and not (layer0_outputs(2535));
    outputs(2329) <= not(layer0_outputs(5623));
    outputs(2330) <= (layer0_outputs(1733)) and (layer0_outputs(7541));
    outputs(2331) <= not(layer0_outputs(616));
    outputs(2332) <= (layer0_outputs(5473)) and (layer0_outputs(6991));
    outputs(2333) <= (layer0_outputs(3073)) and (layer0_outputs(6475));
    outputs(2334) <= not(layer0_outputs(404));
    outputs(2335) <= (layer0_outputs(5961)) and not (layer0_outputs(4900));
    outputs(2336) <= not((layer0_outputs(3828)) and (layer0_outputs(7284)));
    outputs(2337) <= (layer0_outputs(7528)) xor (layer0_outputs(2984));
    outputs(2338) <= not(layer0_outputs(1431));
    outputs(2339) <= (layer0_outputs(2853)) and (layer0_outputs(2329));
    outputs(2340) <= layer0_outputs(5416);
    outputs(2341) <= (layer0_outputs(7674)) and (layer0_outputs(347));
    outputs(2342) <= not((layer0_outputs(5221)) or (layer0_outputs(4650)));
    outputs(2343) <= (layer0_outputs(7274)) xor (layer0_outputs(4470));
    outputs(2344) <= layer0_outputs(2096);
    outputs(2345) <= layer0_outputs(850);
    outputs(2346) <= not(layer0_outputs(812)) or (layer0_outputs(2647));
    outputs(2347) <= layer0_outputs(3223);
    outputs(2348) <= layer0_outputs(1347);
    outputs(2349) <= not(layer0_outputs(2175));
    outputs(2350) <= (layer0_outputs(3971)) and (layer0_outputs(211));
    outputs(2351) <= not(layer0_outputs(7029));
    outputs(2352) <= not(layer0_outputs(2778));
    outputs(2353) <= (layer0_outputs(5993)) or (layer0_outputs(835));
    outputs(2354) <= (layer0_outputs(794)) and (layer0_outputs(443));
    outputs(2355) <= layer0_outputs(3129);
    outputs(2356) <= not(layer0_outputs(4743)) or (layer0_outputs(3270));
    outputs(2357) <= not((layer0_outputs(57)) xor (layer0_outputs(1147)));
    outputs(2358) <= not(layer0_outputs(5365));
    outputs(2359) <= not(layer0_outputs(3267));
    outputs(2360) <= (layer0_outputs(6936)) xor (layer0_outputs(462));
    outputs(2361) <= not((layer0_outputs(1304)) xor (layer0_outputs(2002)));
    outputs(2362) <= (layer0_outputs(4189)) and not (layer0_outputs(6210));
    outputs(2363) <= layer0_outputs(936);
    outputs(2364) <= layer0_outputs(2858);
    outputs(2365) <= (layer0_outputs(4673)) and not (layer0_outputs(201));
    outputs(2366) <= not(layer0_outputs(7589));
    outputs(2367) <= not((layer0_outputs(5913)) or (layer0_outputs(6343)));
    outputs(2368) <= layer0_outputs(5573);
    outputs(2369) <= not(layer0_outputs(4111));
    outputs(2370) <= layer0_outputs(3772);
    outputs(2371) <= not(layer0_outputs(3681));
    outputs(2372) <= not(layer0_outputs(7115));
    outputs(2373) <= layer0_outputs(1417);
    outputs(2374) <= layer0_outputs(3767);
    outputs(2375) <= layer0_outputs(795);
    outputs(2376) <= (layer0_outputs(966)) or (layer0_outputs(697));
    outputs(2377) <= layer0_outputs(5789);
    outputs(2378) <= not(layer0_outputs(1742));
    outputs(2379) <= (layer0_outputs(1078)) and not (layer0_outputs(2384));
    outputs(2380) <= not(layer0_outputs(7213));
    outputs(2381) <= layer0_outputs(3299);
    outputs(2382) <= layer0_outputs(1690);
    outputs(2383) <= not((layer0_outputs(4226)) or (layer0_outputs(5299)));
    outputs(2384) <= (layer0_outputs(1906)) and (layer0_outputs(1398));
    outputs(2385) <= layer0_outputs(2335);
    outputs(2386) <= not((layer0_outputs(2653)) or (layer0_outputs(2033)));
    outputs(2387) <= layer0_outputs(835);
    outputs(2388) <= layer0_outputs(6528);
    outputs(2389) <= not((layer0_outputs(76)) or (layer0_outputs(5235)));
    outputs(2390) <= not(layer0_outputs(1908)) or (layer0_outputs(4389));
    outputs(2391) <= not(layer0_outputs(3474)) or (layer0_outputs(7334));
    outputs(2392) <= (layer0_outputs(7324)) and not (layer0_outputs(5196));
    outputs(2393) <= not(layer0_outputs(3913));
    outputs(2394) <= layer0_outputs(7203);
    outputs(2395) <= layer0_outputs(6027);
    outputs(2396) <= layer0_outputs(90);
    outputs(2397) <= (layer0_outputs(765)) and not (layer0_outputs(2706));
    outputs(2398) <= not(layer0_outputs(358));
    outputs(2399) <= not(layer0_outputs(5959));
    outputs(2400) <= not(layer0_outputs(5971));
    outputs(2401) <= (layer0_outputs(4556)) and not (layer0_outputs(1855));
    outputs(2402) <= (layer0_outputs(2901)) or (layer0_outputs(487));
    outputs(2403) <= not(layer0_outputs(6551));
    outputs(2404) <= not((layer0_outputs(6949)) and (layer0_outputs(2142)));
    outputs(2405) <= not((layer0_outputs(1016)) xor (layer0_outputs(1433)));
    outputs(2406) <= layer0_outputs(6716);
    outputs(2407) <= not(layer0_outputs(413));
    outputs(2408) <= (layer0_outputs(1089)) and not (layer0_outputs(1947));
    outputs(2409) <= not(layer0_outputs(4676));
    outputs(2410) <= (layer0_outputs(7045)) and not (layer0_outputs(6057));
    outputs(2411) <= not(layer0_outputs(640)) or (layer0_outputs(6257));
    outputs(2412) <= not(layer0_outputs(233));
    outputs(2413) <= layer0_outputs(4257);
    outputs(2414) <= not(layer0_outputs(7167)) or (layer0_outputs(1229));
    outputs(2415) <= (layer0_outputs(2802)) and not (layer0_outputs(3328));
    outputs(2416) <= layer0_outputs(3678);
    outputs(2417) <= (layer0_outputs(7066)) and (layer0_outputs(6186));
    outputs(2418) <= layer0_outputs(6036);
    outputs(2419) <= (layer0_outputs(2640)) and (layer0_outputs(5087));
    outputs(2420) <= layer0_outputs(1878);
    outputs(2421) <= layer0_outputs(2981);
    outputs(2422) <= not(layer0_outputs(2607));
    outputs(2423) <= (layer0_outputs(7377)) xor (layer0_outputs(4914));
    outputs(2424) <= layer0_outputs(3560);
    outputs(2425) <= (layer0_outputs(3433)) and (layer0_outputs(4915));
    outputs(2426) <= not(layer0_outputs(6829));
    outputs(2427) <= not(layer0_outputs(5238));
    outputs(2428) <= not(layer0_outputs(6593)) or (layer0_outputs(3180));
    outputs(2429) <= not(layer0_outputs(1389));
    outputs(2430) <= layer0_outputs(4691);
    outputs(2431) <= (layer0_outputs(7592)) and (layer0_outputs(634));
    outputs(2432) <= (layer0_outputs(6673)) and not (layer0_outputs(1947));
    outputs(2433) <= not((layer0_outputs(2573)) xor (layer0_outputs(2579)));
    outputs(2434) <= not(layer0_outputs(7309));
    outputs(2435) <= not(layer0_outputs(5816));
    outputs(2436) <= (layer0_outputs(5843)) and not (layer0_outputs(6000));
    outputs(2437) <= (layer0_outputs(2564)) and not (layer0_outputs(4183));
    outputs(2438) <= layer0_outputs(4804);
    outputs(2439) <= not(layer0_outputs(5357)) or (layer0_outputs(3722));
    outputs(2440) <= (layer0_outputs(7155)) and not (layer0_outputs(528));
    outputs(2441) <= (layer0_outputs(7326)) and not (layer0_outputs(7062));
    outputs(2442) <= not(layer0_outputs(200));
    outputs(2443) <= not((layer0_outputs(1875)) xor (layer0_outputs(2398)));
    outputs(2444) <= not(layer0_outputs(1406));
    outputs(2445) <= layer0_outputs(6341);
    outputs(2446) <= not((layer0_outputs(524)) xor (layer0_outputs(3523)));
    outputs(2447) <= (layer0_outputs(1629)) and not (layer0_outputs(1560));
    outputs(2448) <= not(layer0_outputs(7588));
    outputs(2449) <= layer0_outputs(6741);
    outputs(2450) <= (layer0_outputs(6352)) or (layer0_outputs(6822));
    outputs(2451) <= layer0_outputs(7452);
    outputs(2452) <= layer0_outputs(3603);
    outputs(2453) <= not(layer0_outputs(2283));
    outputs(2454) <= not(layer0_outputs(1853));
    outputs(2455) <= (layer0_outputs(1343)) and not (layer0_outputs(4745));
    outputs(2456) <= not(layer0_outputs(5240));
    outputs(2457) <= layer0_outputs(1364);
    outputs(2458) <= not(layer0_outputs(755));
    outputs(2459) <= not((layer0_outputs(4758)) or (layer0_outputs(3229)));
    outputs(2460) <= not(layer0_outputs(6539));
    outputs(2461) <= layer0_outputs(4427);
    outputs(2462) <= not((layer0_outputs(225)) or (layer0_outputs(5214)));
    outputs(2463) <= not(layer0_outputs(1372));
    outputs(2464) <= not(layer0_outputs(6129));
    outputs(2465) <= (layer0_outputs(5341)) or (layer0_outputs(5397));
    outputs(2466) <= not(layer0_outputs(5994));
    outputs(2467) <= not(layer0_outputs(5141));
    outputs(2468) <= not(layer0_outputs(7407));
    outputs(2469) <= not(layer0_outputs(3690));
    outputs(2470) <= not(layer0_outputs(7652)) or (layer0_outputs(827));
    outputs(2471) <= not(layer0_outputs(6540)) or (layer0_outputs(2397));
    outputs(2472) <= (layer0_outputs(4190)) or (layer0_outputs(515));
    outputs(2473) <= not(layer0_outputs(6414));
    outputs(2474) <= (layer0_outputs(4892)) and (layer0_outputs(3317));
    outputs(2475) <= not(layer0_outputs(2490));
    outputs(2476) <= not(layer0_outputs(2850));
    outputs(2477) <= (layer0_outputs(3633)) and not (layer0_outputs(7347));
    outputs(2478) <= layer0_outputs(2204);
    outputs(2479) <= not(layer0_outputs(2739));
    outputs(2480) <= layer0_outputs(1698);
    outputs(2481) <= layer0_outputs(442);
    outputs(2482) <= not(layer0_outputs(3001)) or (layer0_outputs(6366));
    outputs(2483) <= (layer0_outputs(2501)) and not (layer0_outputs(3173));
    outputs(2484) <= not(layer0_outputs(82));
    outputs(2485) <= layer0_outputs(6357);
    outputs(2486) <= not(layer0_outputs(3918)) or (layer0_outputs(1075));
    outputs(2487) <= not((layer0_outputs(3713)) or (layer0_outputs(6378)));
    outputs(2488) <= (layer0_outputs(5900)) and not (layer0_outputs(6178));
    outputs(2489) <= not(layer0_outputs(1234));
    outputs(2490) <= (layer0_outputs(6336)) xor (layer0_outputs(3727));
    outputs(2491) <= (layer0_outputs(7650)) and (layer0_outputs(1109));
    outputs(2492) <= not(layer0_outputs(6944));
    outputs(2493) <= layer0_outputs(7058);
    outputs(2494) <= (layer0_outputs(2244)) xor (layer0_outputs(3387));
    outputs(2495) <= not((layer0_outputs(3573)) or (layer0_outputs(4457)));
    outputs(2496) <= not(layer0_outputs(3295)) or (layer0_outputs(331));
    outputs(2497) <= not(layer0_outputs(7018));
    outputs(2498) <= (layer0_outputs(6293)) and not (layer0_outputs(852));
    outputs(2499) <= not(layer0_outputs(2228)) or (layer0_outputs(699));
    outputs(2500) <= (layer0_outputs(4945)) and not (layer0_outputs(6842));
    outputs(2501) <= (layer0_outputs(1590)) and not (layer0_outputs(7536));
    outputs(2502) <= not(layer0_outputs(407)) or (layer0_outputs(6614));
    outputs(2503) <= not(layer0_outputs(620)) or (layer0_outputs(2385));
    outputs(2504) <= (layer0_outputs(7117)) and not (layer0_outputs(114));
    outputs(2505) <= (layer0_outputs(4225)) and not (layer0_outputs(7059));
    outputs(2506) <= (layer0_outputs(4683)) and not (layer0_outputs(1971));
    outputs(2507) <= layer0_outputs(3187);
    outputs(2508) <= (layer0_outputs(7637)) or (layer0_outputs(1560));
    outputs(2509) <= not(layer0_outputs(7462));
    outputs(2510) <= not(layer0_outputs(6123));
    outputs(2511) <= layer0_outputs(2576);
    outputs(2512) <= (layer0_outputs(7276)) and (layer0_outputs(6537));
    outputs(2513) <= (layer0_outputs(7414)) and not (layer0_outputs(1216));
    outputs(2514) <= layer0_outputs(7031);
    outputs(2515) <= not((layer0_outputs(6791)) xor (layer0_outputs(4849)));
    outputs(2516) <= not(layer0_outputs(6269));
    outputs(2517) <= (layer0_outputs(5781)) and not (layer0_outputs(4932));
    outputs(2518) <= not(layer0_outputs(1143));
    outputs(2519) <= not(layer0_outputs(3755)) or (layer0_outputs(6211));
    outputs(2520) <= (layer0_outputs(5197)) xor (layer0_outputs(1153));
    outputs(2521) <= layer0_outputs(235);
    outputs(2522) <= (layer0_outputs(2560)) xor (layer0_outputs(6148));
    outputs(2523) <= (layer0_outputs(334)) xor (layer0_outputs(230));
    outputs(2524) <= layer0_outputs(3947);
    outputs(2525) <= (layer0_outputs(3860)) xor (layer0_outputs(4020));
    outputs(2526) <= (layer0_outputs(5559)) xor (layer0_outputs(848));
    outputs(2527) <= not((layer0_outputs(3052)) xor (layer0_outputs(1533)));
    outputs(2528) <= not(layer0_outputs(6501)) or (layer0_outputs(396));
    outputs(2529) <= not(layer0_outputs(3627));
    outputs(2530) <= layer0_outputs(6326);
    outputs(2531) <= layer0_outputs(4642);
    outputs(2532) <= layer0_outputs(1318);
    outputs(2533) <= not(layer0_outputs(3221));
    outputs(2534) <= not(layer0_outputs(3499));
    outputs(2535) <= not(layer0_outputs(1187)) or (layer0_outputs(3783));
    outputs(2536) <= layer0_outputs(4834);
    outputs(2537) <= layer0_outputs(3885);
    outputs(2538) <= layer0_outputs(7318);
    outputs(2539) <= not((layer0_outputs(6126)) and (layer0_outputs(3973)));
    outputs(2540) <= layer0_outputs(7530);
    outputs(2541) <= (layer0_outputs(3827)) and (layer0_outputs(4189));
    outputs(2542) <= layer0_outputs(4263);
    outputs(2543) <= (layer0_outputs(1744)) and not (layer0_outputs(3814));
    outputs(2544) <= layer0_outputs(2689);
    outputs(2545) <= not((layer0_outputs(3215)) xor (layer0_outputs(6691)));
    outputs(2546) <= (layer0_outputs(5304)) and not (layer0_outputs(108));
    outputs(2547) <= not(layer0_outputs(7025));
    outputs(2548) <= not(layer0_outputs(6969));
    outputs(2549) <= not(layer0_outputs(114));
    outputs(2550) <= layer0_outputs(20);
    outputs(2551) <= not(layer0_outputs(6545));
    outputs(2552) <= (layer0_outputs(5727)) and not (layer0_outputs(5722));
    outputs(2553) <= (layer0_outputs(6409)) xor (layer0_outputs(3392));
    outputs(2554) <= layer0_outputs(6389);
    outputs(2555) <= layer0_outputs(4451);
    outputs(2556) <= not(layer0_outputs(6661));
    outputs(2557) <= layer0_outputs(7552);
    outputs(2558) <= layer0_outputs(2840);
    outputs(2559) <= (layer0_outputs(1773)) and not (layer0_outputs(471));
    outputs(2560) <= (layer0_outputs(1763)) and (layer0_outputs(6777));
    outputs(2561) <= not(layer0_outputs(4054));
    outputs(2562) <= (layer0_outputs(2554)) and not (layer0_outputs(3040));
    outputs(2563) <= (layer0_outputs(2289)) and not (layer0_outputs(3660));
    outputs(2564) <= layer0_outputs(3198);
    outputs(2565) <= not(layer0_outputs(5453));
    outputs(2566) <= layer0_outputs(3358);
    outputs(2567) <= layer0_outputs(1643);
    outputs(2568) <= not((layer0_outputs(984)) or (layer0_outputs(346)));
    outputs(2569) <= layer0_outputs(505);
    outputs(2570) <= not((layer0_outputs(2176)) xor (layer0_outputs(300)));
    outputs(2571) <= layer0_outputs(1453);
    outputs(2572) <= not((layer0_outputs(581)) and (layer0_outputs(6561)));
    outputs(2573) <= not(layer0_outputs(6703));
    outputs(2574) <= (layer0_outputs(6128)) xor (layer0_outputs(6978));
    outputs(2575) <= (layer0_outputs(3512)) and not (layer0_outputs(485));
    outputs(2576) <= not(layer0_outputs(5764));
    outputs(2577) <= layer0_outputs(1119);
    outputs(2578) <= not(layer0_outputs(4750)) or (layer0_outputs(1081));
    outputs(2579) <= (layer0_outputs(1714)) and not (layer0_outputs(1674));
    outputs(2580) <= layer0_outputs(2546);
    outputs(2581) <= layer0_outputs(2376);
    outputs(2582) <= layer0_outputs(265);
    outputs(2583) <= not(layer0_outputs(2275));
    outputs(2584) <= (layer0_outputs(4147)) and not (layer0_outputs(6672));
    outputs(2585) <= not(layer0_outputs(1865));
    outputs(2586) <= not((layer0_outputs(1106)) or (layer0_outputs(128)));
    outputs(2587) <= layer0_outputs(5121);
    outputs(2588) <= not(layer0_outputs(6209));
    outputs(2589) <= (layer0_outputs(3071)) and not (layer0_outputs(256));
    outputs(2590) <= not(layer0_outputs(6883));
    outputs(2591) <= (layer0_outputs(5271)) xor (layer0_outputs(4026));
    outputs(2592) <= layer0_outputs(336);
    outputs(2593) <= (layer0_outputs(3362)) xor (layer0_outputs(2846));
    outputs(2594) <= layer0_outputs(1637);
    outputs(2595) <= not(layer0_outputs(2047));
    outputs(2596) <= layer0_outputs(1992);
    outputs(2597) <= (layer0_outputs(7631)) and not (layer0_outputs(6447));
    outputs(2598) <= layer0_outputs(2105);
    outputs(2599) <= not((layer0_outputs(2979)) or (layer0_outputs(3146)));
    outputs(2600) <= not((layer0_outputs(6603)) or (layer0_outputs(5345)));
    outputs(2601) <= layer0_outputs(179);
    outputs(2602) <= layer0_outputs(7209);
    outputs(2603) <= layer0_outputs(4396);
    outputs(2604) <= not(layer0_outputs(4541));
    outputs(2605) <= layer0_outputs(933);
    outputs(2606) <= layer0_outputs(3723);
    outputs(2607) <= (layer0_outputs(7522)) and (layer0_outputs(5358));
    outputs(2608) <= not((layer0_outputs(58)) or (layer0_outputs(4087)));
    outputs(2609) <= not(layer0_outputs(7024)) or (layer0_outputs(4438));
    outputs(2610) <= layer0_outputs(191);
    outputs(2611) <= (layer0_outputs(5497)) xor (layer0_outputs(4581));
    outputs(2612) <= layer0_outputs(1159);
    outputs(2613) <= (layer0_outputs(6035)) xor (layer0_outputs(1189));
    outputs(2614) <= layer0_outputs(94);
    outputs(2615) <= (layer0_outputs(3827)) and (layer0_outputs(3068));
    outputs(2616) <= not((layer0_outputs(1171)) and (layer0_outputs(5670)));
    outputs(2617) <= not(layer0_outputs(1636));
    outputs(2618) <= not(layer0_outputs(2080));
    outputs(2619) <= not((layer0_outputs(3425)) xor (layer0_outputs(2521)));
    outputs(2620) <= not(layer0_outputs(2844));
    outputs(2621) <= (layer0_outputs(3738)) and not (layer0_outputs(7049));
    outputs(2622) <= not(layer0_outputs(4350));
    outputs(2623) <= layer0_outputs(1575);
    outputs(2624) <= (layer0_outputs(6005)) and (layer0_outputs(3448));
    outputs(2625) <= layer0_outputs(1421);
    outputs(2626) <= not((layer0_outputs(4288)) and (layer0_outputs(6837)));
    outputs(2627) <= not(layer0_outputs(6231));
    outputs(2628) <= (layer0_outputs(4184)) and not (layer0_outputs(4629));
    outputs(2629) <= not(layer0_outputs(6031));
    outputs(2630) <= (layer0_outputs(2837)) and (layer0_outputs(5958));
    outputs(2631) <= (layer0_outputs(6203)) xor (layer0_outputs(6761));
    outputs(2632) <= (layer0_outputs(5494)) and not (layer0_outputs(829));
    outputs(2633) <= (layer0_outputs(2688)) and not (layer0_outputs(6499));
    outputs(2634) <= layer0_outputs(155);
    outputs(2635) <= layer0_outputs(4787);
    outputs(2636) <= (layer0_outputs(3592)) and (layer0_outputs(4052));
    outputs(2637) <= not(layer0_outputs(2402));
    outputs(2638) <= layer0_outputs(4284);
    outputs(2639) <= (layer0_outputs(4993)) and (layer0_outputs(6700));
    outputs(2640) <= (layer0_outputs(1540)) and not (layer0_outputs(1861));
    outputs(2641) <= layer0_outputs(615);
    outputs(2642) <= (layer0_outputs(4879)) and not (layer0_outputs(5921));
    outputs(2643) <= layer0_outputs(2381);
    outputs(2644) <= not(layer0_outputs(377));
    outputs(2645) <= not(layer0_outputs(2888));
    outputs(2646) <= not((layer0_outputs(4437)) xor (layer0_outputs(5066)));
    outputs(2647) <= (layer0_outputs(3706)) and not (layer0_outputs(1388));
    outputs(2648) <= not((layer0_outputs(1720)) or (layer0_outputs(992)));
    outputs(2649) <= not((layer0_outputs(2568)) or (layer0_outputs(738)));
    outputs(2650) <= not((layer0_outputs(2648)) xor (layer0_outputs(265)));
    outputs(2651) <= (layer0_outputs(5044)) and not (layer0_outputs(3842));
    outputs(2652) <= (layer0_outputs(5109)) and (layer0_outputs(7671));
    outputs(2653) <= (layer0_outputs(332)) and not (layer0_outputs(2448));
    outputs(2654) <= (layer0_outputs(5599)) and not (layer0_outputs(2383));
    outputs(2655) <= not((layer0_outputs(875)) or (layer0_outputs(5856)));
    outputs(2656) <= not((layer0_outputs(4791)) or (layer0_outputs(3628)));
    outputs(2657) <= (layer0_outputs(1724)) or (layer0_outputs(2147));
    outputs(2658) <= layer0_outputs(3795);
    outputs(2659) <= (layer0_outputs(3849)) and not (layer0_outputs(1321));
    outputs(2660) <= (layer0_outputs(2378)) xor (layer0_outputs(3887));
    outputs(2661) <= not(layer0_outputs(1506));
    outputs(2662) <= not(layer0_outputs(6711)) or (layer0_outputs(5599));
    outputs(2663) <= layer0_outputs(5970);
    outputs(2664) <= layer0_outputs(5914);
    outputs(2665) <= not(layer0_outputs(6495));
    outputs(2666) <= layer0_outputs(3108);
    outputs(2667) <= layer0_outputs(6825);
    outputs(2668) <= not(layer0_outputs(6467));
    outputs(2669) <= not(layer0_outputs(792));
    outputs(2670) <= (layer0_outputs(2217)) xor (layer0_outputs(2246));
    outputs(2671) <= (layer0_outputs(5305)) and not (layer0_outputs(3754));
    outputs(2672) <= layer0_outputs(800);
    outputs(2673) <= not(layer0_outputs(6188));
    outputs(2674) <= not((layer0_outputs(3238)) and (layer0_outputs(1908)));
    outputs(2675) <= not(layer0_outputs(3762));
    outputs(2676) <= layer0_outputs(4824);
    outputs(2677) <= (layer0_outputs(777)) and not (layer0_outputs(3219));
    outputs(2678) <= (layer0_outputs(2677)) or (layer0_outputs(6376));
    outputs(2679) <= layer0_outputs(2999);
    outputs(2680) <= (layer0_outputs(3799)) and not (layer0_outputs(4579));
    outputs(2681) <= (layer0_outputs(250)) and not (layer0_outputs(3489));
    outputs(2682) <= not(layer0_outputs(604));
    outputs(2683) <= (layer0_outputs(5495)) and (layer0_outputs(7445));
    outputs(2684) <= not(layer0_outputs(1568));
    outputs(2685) <= not(layer0_outputs(4365)) or (layer0_outputs(91));
    outputs(2686) <= not((layer0_outputs(6868)) xor (layer0_outputs(3014)));
    outputs(2687) <= (layer0_outputs(2121)) and not (layer0_outputs(6539));
    outputs(2688) <= (layer0_outputs(854)) and (layer0_outputs(6433));
    outputs(2689) <= (layer0_outputs(6266)) and not (layer0_outputs(2979));
    outputs(2690) <= not((layer0_outputs(1338)) and (layer0_outputs(4762)));
    outputs(2691) <= (layer0_outputs(1690)) and (layer0_outputs(1715));
    outputs(2692) <= (layer0_outputs(814)) xor (layer0_outputs(4840));
    outputs(2693) <= (layer0_outputs(1753)) xor (layer0_outputs(2216));
    outputs(2694) <= layer0_outputs(832);
    outputs(2695) <= not((layer0_outputs(1329)) and (layer0_outputs(5401)));
    outputs(2696) <= layer0_outputs(769);
    outputs(2697) <= (layer0_outputs(4435)) or (layer0_outputs(3793));
    outputs(2698) <= not((layer0_outputs(7638)) or (layer0_outputs(6198)));
    outputs(2699) <= not(layer0_outputs(6307));
    outputs(2700) <= not(layer0_outputs(7454));
    outputs(2701) <= not((layer0_outputs(6927)) or (layer0_outputs(984)));
    outputs(2702) <= not(layer0_outputs(401));
    outputs(2703) <= (layer0_outputs(288)) or (layer0_outputs(6749));
    outputs(2704) <= layer0_outputs(6354);
    outputs(2705) <= layer0_outputs(4182);
    outputs(2706) <= not(layer0_outputs(7426));
    outputs(2707) <= not(layer0_outputs(3800));
    outputs(2708) <= layer0_outputs(3158);
    outputs(2709) <= layer0_outputs(3123);
    outputs(2710) <= (layer0_outputs(6405)) and (layer0_outputs(6207));
    outputs(2711) <= layer0_outputs(1661);
    outputs(2712) <= not(layer0_outputs(5475)) or (layer0_outputs(369));
    outputs(2713) <= not(layer0_outputs(4185));
    outputs(2714) <= layer0_outputs(2291);
    outputs(2715) <= not(layer0_outputs(6946));
    outputs(2716) <= layer0_outputs(5398);
    outputs(2717) <= not((layer0_outputs(2307)) xor (layer0_outputs(3150)));
    outputs(2718) <= not(layer0_outputs(2133));
    outputs(2719) <= not(layer0_outputs(2746));
    outputs(2720) <= not(layer0_outputs(6619));
    outputs(2721) <= layer0_outputs(997);
    outputs(2722) <= not(layer0_outputs(3164)) or (layer0_outputs(6163));
    outputs(2723) <= not(layer0_outputs(1512));
    outputs(2724) <= (layer0_outputs(3448)) and not (layer0_outputs(6524));
    outputs(2725) <= not(layer0_outputs(4279));
    outputs(2726) <= (layer0_outputs(6067)) xor (layer0_outputs(5802));
    outputs(2727) <= not(layer0_outputs(1482));
    outputs(2728) <= not(layer0_outputs(3375));
    outputs(2729) <= layer0_outputs(5068);
    outputs(2730) <= layer0_outputs(3775);
    outputs(2731) <= not(layer0_outputs(618)) or (layer0_outputs(144));
    outputs(2732) <= not((layer0_outputs(7472)) or (layer0_outputs(2779)));
    outputs(2733) <= not(layer0_outputs(2888));
    outputs(2734) <= (layer0_outputs(4920)) or (layer0_outputs(6385));
    outputs(2735) <= not(layer0_outputs(721));
    outputs(2736) <= (layer0_outputs(7343)) or (layer0_outputs(2659));
    outputs(2737) <= layer0_outputs(7012);
    outputs(2738) <= (layer0_outputs(2002)) and not (layer0_outputs(3496));
    outputs(2739) <= not((layer0_outputs(7293)) or (layer0_outputs(7042)));
    outputs(2740) <= not(layer0_outputs(4767));
    outputs(2741) <= (layer0_outputs(4756)) and (layer0_outputs(7121));
    outputs(2742) <= not((layer0_outputs(716)) xor (layer0_outputs(7177)));
    outputs(2743) <= (layer0_outputs(2187)) and (layer0_outputs(7620));
    outputs(2744) <= layer0_outputs(7322);
    outputs(2745) <= not(layer0_outputs(7345));
    outputs(2746) <= not((layer0_outputs(4240)) xor (layer0_outputs(4565)));
    outputs(2747) <= (layer0_outputs(7665)) xor (layer0_outputs(3643));
    outputs(2748) <= not(layer0_outputs(4931));
    outputs(2749) <= (layer0_outputs(2441)) xor (layer0_outputs(4997));
    outputs(2750) <= (layer0_outputs(7346)) xor (layer0_outputs(293));
    outputs(2751) <= layer0_outputs(2160);
    outputs(2752) <= layer0_outputs(7279);
    outputs(2753) <= not(layer0_outputs(2164)) or (layer0_outputs(86));
    outputs(2754) <= (layer0_outputs(4116)) and not (layer0_outputs(2004));
    outputs(2755) <= layer0_outputs(5667);
    outputs(2756) <= layer0_outputs(3616);
    outputs(2757) <= not(layer0_outputs(2413));
    outputs(2758) <= (layer0_outputs(1925)) and not (layer0_outputs(3895));
    outputs(2759) <= (layer0_outputs(7101)) or (layer0_outputs(2972));
    outputs(2760) <= not(layer0_outputs(4010));
    outputs(2761) <= not(layer0_outputs(4050));
    outputs(2762) <= layer0_outputs(5589);
    outputs(2763) <= not((layer0_outputs(7313)) or (layer0_outputs(3538)));
    outputs(2764) <= not((layer0_outputs(1874)) or (layer0_outputs(6905)));
    outputs(2765) <= layer0_outputs(6571);
    outputs(2766) <= not(layer0_outputs(2099));
    outputs(2767) <= not(layer0_outputs(2961)) or (layer0_outputs(4479));
    outputs(2768) <= not(layer0_outputs(5523)) or (layer0_outputs(451));
    outputs(2769) <= (layer0_outputs(1138)) or (layer0_outputs(1395));
    outputs(2770) <= not(layer0_outputs(4353)) or (layer0_outputs(6891));
    outputs(2771) <= not(layer0_outputs(1780));
    outputs(2772) <= (layer0_outputs(5404)) and not (layer0_outputs(4242));
    outputs(2773) <= not(layer0_outputs(892));
    outputs(2774) <= not(layer0_outputs(6845));
    outputs(2775) <= not(layer0_outputs(1671));
    outputs(2776) <= not(layer0_outputs(5942)) or (layer0_outputs(5135));
    outputs(2777) <= not((layer0_outputs(2512)) or (layer0_outputs(2847)));
    outputs(2778) <= not((layer0_outputs(7391)) xor (layer0_outputs(376)));
    outputs(2779) <= not(layer0_outputs(3040)) or (layer0_outputs(4218));
    outputs(2780) <= not(layer0_outputs(704));
    outputs(2781) <= not(layer0_outputs(5088)) or (layer0_outputs(531));
    outputs(2782) <= layer0_outputs(9);
    outputs(2783) <= (layer0_outputs(4039)) and not (layer0_outputs(385));
    outputs(2784) <= not(layer0_outputs(3743));
    outputs(2785) <= not(layer0_outputs(5250));
    outputs(2786) <= not((layer0_outputs(7065)) xor (layer0_outputs(2894)));
    outputs(2787) <= layer0_outputs(1803);
    outputs(2788) <= not(layer0_outputs(1565)) or (layer0_outputs(583));
    outputs(2789) <= not(layer0_outputs(2332));
    outputs(2790) <= not(layer0_outputs(4236));
    outputs(2791) <= not(layer0_outputs(7260));
    outputs(2792) <= (layer0_outputs(3633)) or (layer0_outputs(74));
    outputs(2793) <= not((layer0_outputs(2869)) and (layer0_outputs(4213)));
    outputs(2794) <= not(layer0_outputs(6969));
    outputs(2795) <= not(layer0_outputs(3297));
    outputs(2796) <= not(layer0_outputs(2029));
    outputs(2797) <= (layer0_outputs(1801)) and not (layer0_outputs(4391));
    outputs(2798) <= not(layer0_outputs(2852));
    outputs(2799) <= layer0_outputs(4123);
    outputs(2800) <= (layer0_outputs(1014)) xor (layer0_outputs(2486));
    outputs(2801) <= not(layer0_outputs(5776)) or (layer0_outputs(4322));
    outputs(2802) <= (layer0_outputs(6912)) and not (layer0_outputs(4258));
    outputs(2803) <= layer0_outputs(1518);
    outputs(2804) <= not(layer0_outputs(2748));
    outputs(2805) <= not((layer0_outputs(7397)) and (layer0_outputs(7551)));
    outputs(2806) <= not((layer0_outputs(4364)) or (layer0_outputs(3034)));
    outputs(2807) <= not(layer0_outputs(3598));
    outputs(2808) <= not(layer0_outputs(4686));
    outputs(2809) <= layer0_outputs(3198);
    outputs(2810) <= (layer0_outputs(257)) or (layer0_outputs(6347));
    outputs(2811) <= not((layer0_outputs(5216)) xor (layer0_outputs(6301)));
    outputs(2812) <= not(layer0_outputs(6951));
    outputs(2813) <= not(layer0_outputs(624));
    outputs(2814) <= not(layer0_outputs(6317));
    outputs(2815) <= not(layer0_outputs(3157));
    outputs(2816) <= (layer0_outputs(5231)) xor (layer0_outputs(3914));
    outputs(2817) <= (layer0_outputs(6168)) xor (layer0_outputs(6770));
    outputs(2818) <= not((layer0_outputs(2683)) and (layer0_outputs(2490)));
    outputs(2819) <= not(layer0_outputs(6925));
    outputs(2820) <= layer0_outputs(6227);
    outputs(2821) <= not((layer0_outputs(3321)) xor (layer0_outputs(4568)));
    outputs(2822) <= not((layer0_outputs(223)) xor (layer0_outputs(3757)));
    outputs(2823) <= layer0_outputs(4317);
    outputs(2824) <= (layer0_outputs(3735)) and not (layer0_outputs(7554));
    outputs(2825) <= not(layer0_outputs(1745));
    outputs(2826) <= (layer0_outputs(5820)) and not (layer0_outputs(4841));
    outputs(2827) <= layer0_outputs(2521);
    outputs(2828) <= not(layer0_outputs(2855));
    outputs(2829) <= layer0_outputs(3442);
    outputs(2830) <= (layer0_outputs(3707)) xor (layer0_outputs(7093));
    outputs(2831) <= (layer0_outputs(3259)) or (layer0_outputs(3101));
    outputs(2832) <= (layer0_outputs(412)) and (layer0_outputs(601));
    outputs(2833) <= layer0_outputs(4815);
    outputs(2834) <= (layer0_outputs(4255)) and (layer0_outputs(7270));
    outputs(2835) <= (layer0_outputs(3092)) xor (layer0_outputs(3765));
    outputs(2836) <= not(layer0_outputs(6833)) or (layer0_outputs(4563));
    outputs(2837) <= (layer0_outputs(5580)) xor (layer0_outputs(7587));
    outputs(2838) <= layer0_outputs(5966);
    outputs(2839) <= not(layer0_outputs(7206));
    outputs(2840) <= not((layer0_outputs(6709)) xor (layer0_outputs(1088)));
    outputs(2841) <= not(layer0_outputs(7232)) or (layer0_outputs(2429));
    outputs(2842) <= not(layer0_outputs(1697));
    outputs(2843) <= not((layer0_outputs(4744)) xor (layer0_outputs(7668)));
    outputs(2844) <= (layer0_outputs(1336)) or (layer0_outputs(5800));
    outputs(2845) <= layer0_outputs(2259);
    outputs(2846) <= layer0_outputs(2152);
    outputs(2847) <= not(layer0_outputs(6764));
    outputs(2848) <= not(layer0_outputs(840));
    outputs(2849) <= not(layer0_outputs(3103)) or (layer0_outputs(2419));
    outputs(2850) <= (layer0_outputs(338)) xor (layer0_outputs(67));
    outputs(2851) <= not(layer0_outputs(6538));
    outputs(2852) <= not(layer0_outputs(4140));
    outputs(2853) <= (layer0_outputs(1093)) xor (layer0_outputs(6942));
    outputs(2854) <= not(layer0_outputs(5176));
    outputs(2855) <= not((layer0_outputs(3497)) and (layer0_outputs(1440)));
    outputs(2856) <= (layer0_outputs(5653)) xor (layer0_outputs(5182));
    outputs(2857) <= not(layer0_outputs(6838)) or (layer0_outputs(2030));
    outputs(2858) <= layer0_outputs(4907);
    outputs(2859) <= (layer0_outputs(1481)) and not (layer0_outputs(5729));
    outputs(2860) <= not((layer0_outputs(3455)) or (layer0_outputs(5873)));
    outputs(2861) <= not(layer0_outputs(5636));
    outputs(2862) <= layer0_outputs(3890);
    outputs(2863) <= not(layer0_outputs(4410));
    outputs(2864) <= (layer0_outputs(6010)) and (layer0_outputs(6445));
    outputs(2865) <= not(layer0_outputs(3076));
    outputs(2866) <= (layer0_outputs(3603)) and not (layer0_outputs(5337));
    outputs(2867) <= not(layer0_outputs(3436));
    outputs(2868) <= layer0_outputs(814);
    outputs(2869) <= not((layer0_outputs(4008)) and (layer0_outputs(5669)));
    outputs(2870) <= not((layer0_outputs(4636)) xor (layer0_outputs(7354)));
    outputs(2871) <= not(layer0_outputs(3731));
    outputs(2872) <= layer0_outputs(4063);
    outputs(2873) <= (layer0_outputs(6663)) and not (layer0_outputs(917));
    outputs(2874) <= not(layer0_outputs(5303));
    outputs(2875) <= (layer0_outputs(596)) xor (layer0_outputs(3057));
    outputs(2876) <= (layer0_outputs(1206)) and not (layer0_outputs(6900));
    outputs(2877) <= not(layer0_outputs(1842));
    outputs(2878) <= layer0_outputs(1792);
    outputs(2879) <= not(layer0_outputs(3692));
    outputs(2880) <= not(layer0_outputs(1682)) or (layer0_outputs(6617));
    outputs(2881) <= layer0_outputs(6322);
    outputs(2882) <= (layer0_outputs(2469)) and not (layer0_outputs(2261));
    outputs(2883) <= not(layer0_outputs(2953)) or (layer0_outputs(6570));
    outputs(2884) <= (layer0_outputs(5637)) and not (layer0_outputs(7395));
    outputs(2885) <= layer0_outputs(5098);
    outputs(2886) <= not(layer0_outputs(6479));
    outputs(2887) <= not(layer0_outputs(6738));
    outputs(2888) <= layer0_outputs(4815);
    outputs(2889) <= not(layer0_outputs(3290)) or (layer0_outputs(1740));
    outputs(2890) <= (layer0_outputs(1382)) and not (layer0_outputs(2791));
    outputs(2891) <= not((layer0_outputs(6532)) or (layer0_outputs(6790)));
    outputs(2892) <= layer0_outputs(2577);
    outputs(2893) <= layer0_outputs(1689);
    outputs(2894) <= not((layer0_outputs(6695)) or (layer0_outputs(2675)));
    outputs(2895) <= not(layer0_outputs(1216));
    outputs(2896) <= not(layer0_outputs(2538)) or (layer0_outputs(3107));
    outputs(2897) <= (layer0_outputs(5263)) and not (layer0_outputs(4512));
    outputs(2898) <= not((layer0_outputs(3009)) xor (layer0_outputs(5798)));
    outputs(2899) <= not(layer0_outputs(3219));
    outputs(2900) <= not((layer0_outputs(7033)) xor (layer0_outputs(2086)));
    outputs(2901) <= (layer0_outputs(5455)) and not (layer0_outputs(34));
    outputs(2902) <= not(layer0_outputs(6704));
    outputs(2903) <= layer0_outputs(2651);
    outputs(2904) <= (layer0_outputs(1698)) and (layer0_outputs(303));
    outputs(2905) <= not(layer0_outputs(1020)) or (layer0_outputs(2874));
    outputs(2906) <= (layer0_outputs(5148)) and not (layer0_outputs(781));
    outputs(2907) <= not(layer0_outputs(1693));
    outputs(2908) <= not((layer0_outputs(525)) or (layer0_outputs(4813)));
    outputs(2909) <= (layer0_outputs(6140)) and not (layer0_outputs(4030));
    outputs(2910) <= layer0_outputs(700);
    outputs(2911) <= not((layer0_outputs(1655)) xor (layer0_outputs(1056)));
    outputs(2912) <= not(layer0_outputs(6396)) or (layer0_outputs(842));
    outputs(2913) <= (layer0_outputs(246)) or (layer0_outputs(1704));
    outputs(2914) <= layer0_outputs(4959);
    outputs(2915) <= layer0_outputs(2447);
    outputs(2916) <= not(layer0_outputs(5119)) or (layer0_outputs(2549));
    outputs(2917) <= layer0_outputs(5924);
    outputs(2918) <= not(layer0_outputs(7233));
    outputs(2919) <= not(layer0_outputs(2463));
    outputs(2920) <= (layer0_outputs(4040)) and not (layer0_outputs(4021));
    outputs(2921) <= not(layer0_outputs(2163)) or (layer0_outputs(6145));
    outputs(2922) <= not(layer0_outputs(3916));
    outputs(2923) <= not(layer0_outputs(5073));
    outputs(2924) <= (layer0_outputs(1178)) and not (layer0_outputs(3381));
    outputs(2925) <= not((layer0_outputs(82)) xor (layer0_outputs(1466)));
    outputs(2926) <= not(layer0_outputs(4111));
    outputs(2927) <= not(layer0_outputs(5277));
    outputs(2928) <= layer0_outputs(542);
    outputs(2929) <= layer0_outputs(2999);
    outputs(2930) <= not((layer0_outputs(888)) or (layer0_outputs(4655)));
    outputs(2931) <= layer0_outputs(603);
    outputs(2932) <= not(layer0_outputs(960)) or (layer0_outputs(5876));
    outputs(2933) <= not(layer0_outputs(6437)) or (layer0_outputs(5904));
    outputs(2934) <= not(layer0_outputs(1338)) or (layer0_outputs(6194));
    outputs(2935) <= not(layer0_outputs(188));
    outputs(2936) <= (layer0_outputs(1120)) and not (layer0_outputs(6625));
    outputs(2937) <= not(layer0_outputs(4169));
    outputs(2938) <= (layer0_outputs(5969)) and (layer0_outputs(4429));
    outputs(2939) <= (layer0_outputs(1275)) or (layer0_outputs(7298));
    outputs(2940) <= (layer0_outputs(1436)) and not (layer0_outputs(6039));
    outputs(2941) <= not(layer0_outputs(4962));
    outputs(2942) <= layer0_outputs(3519);
    outputs(2943) <= not(layer0_outputs(2041)) or (layer0_outputs(5855));
    outputs(2944) <= layer0_outputs(6628);
    outputs(2945) <= (layer0_outputs(6904)) xor (layer0_outputs(3388));
    outputs(2946) <= (layer0_outputs(2983)) xor (layer0_outputs(445));
    outputs(2947) <= not((layer0_outputs(4799)) or (layer0_outputs(5729)));
    outputs(2948) <= not(layer0_outputs(3875));
    outputs(2949) <= not((layer0_outputs(5716)) or (layer0_outputs(7579)));
    outputs(2950) <= layer0_outputs(4996);
    outputs(2951) <= layer0_outputs(88);
    outputs(2952) <= not(layer0_outputs(636)) or (layer0_outputs(1559));
    outputs(2953) <= layer0_outputs(3629);
    outputs(2954) <= layer0_outputs(7473);
    outputs(2955) <= not((layer0_outputs(4312)) xor (layer0_outputs(4616)));
    outputs(2956) <= (layer0_outputs(4136)) and (layer0_outputs(6698));
    outputs(2957) <= layer0_outputs(5582);
    outputs(2958) <= (layer0_outputs(17)) and not (layer0_outputs(6509));
    outputs(2959) <= not(layer0_outputs(4831));
    outputs(2960) <= not(layer0_outputs(6292));
    outputs(2961) <= not((layer0_outputs(871)) or (layer0_outputs(6496)));
    outputs(2962) <= (layer0_outputs(495)) and (layer0_outputs(6394));
    outputs(2963) <= (layer0_outputs(7282)) and not (layer0_outputs(6993));
    outputs(2964) <= layer0_outputs(4842);
    outputs(2965) <= (layer0_outputs(611)) and (layer0_outputs(3071));
    outputs(2966) <= layer0_outputs(4596);
    outputs(2967) <= not(layer0_outputs(677));
    outputs(2968) <= not(layer0_outputs(3032));
    outputs(2969) <= (layer0_outputs(4460)) and not (layer0_outputs(3753));
    outputs(2970) <= not(layer0_outputs(2953));
    outputs(2971) <= not((layer0_outputs(6457)) or (layer0_outputs(6635)));
    outputs(2972) <= not((layer0_outputs(4036)) xor (layer0_outputs(6070)));
    outputs(2973) <= (layer0_outputs(1424)) xor (layer0_outputs(5507));
    outputs(2974) <= layer0_outputs(3518);
    outputs(2975) <= not((layer0_outputs(4119)) or (layer0_outputs(6020)));
    outputs(2976) <= (layer0_outputs(701)) or (layer0_outputs(961));
    outputs(2977) <= (layer0_outputs(6419)) and (layer0_outputs(3269));
    outputs(2978) <= not(layer0_outputs(4019));
    outputs(2979) <= layer0_outputs(1328);
    outputs(2980) <= (layer0_outputs(3423)) xor (layer0_outputs(4854));
    outputs(2981) <= not(layer0_outputs(2138)) or (layer0_outputs(3777));
    outputs(2982) <= not(layer0_outputs(4223));
    outputs(2983) <= not(layer0_outputs(5835));
    outputs(2984) <= not(layer0_outputs(706));
    outputs(2985) <= (layer0_outputs(7226)) and not (layer0_outputs(4074));
    outputs(2986) <= (layer0_outputs(5999)) or (layer0_outputs(268));
    outputs(2987) <= (layer0_outputs(919)) and not (layer0_outputs(3561));
    outputs(2988) <= (layer0_outputs(4351)) xor (layer0_outputs(5645));
    outputs(2989) <= not(layer0_outputs(6141)) or (layer0_outputs(2991));
    outputs(2990) <= not(layer0_outputs(1192));
    outputs(2991) <= layer0_outputs(3276);
    outputs(2992) <= (layer0_outputs(7500)) and (layer0_outputs(7286));
    outputs(2993) <= layer0_outputs(1099);
    outputs(2994) <= not(layer0_outputs(5804));
    outputs(2995) <= not(layer0_outputs(364));
    outputs(2996) <= not(layer0_outputs(2000));
    outputs(2997) <= not((layer0_outputs(6486)) xor (layer0_outputs(1482)));
    outputs(2998) <= not(layer0_outputs(6555));
    outputs(2999) <= layer0_outputs(1053);
    outputs(3000) <= layer0_outputs(579);
    outputs(3001) <= not(layer0_outputs(2926)) or (layer0_outputs(985));
    outputs(3002) <= not((layer0_outputs(5795)) or (layer0_outputs(4476)));
    outputs(3003) <= (layer0_outputs(5111)) xor (layer0_outputs(3836));
    outputs(3004) <= not((layer0_outputs(2237)) and (layer0_outputs(6229)));
    outputs(3005) <= not(layer0_outputs(2741));
    outputs(3006) <= not(layer0_outputs(6054));
    outputs(3007) <= not((layer0_outputs(841)) and (layer0_outputs(1385)));
    outputs(3008) <= not((layer0_outputs(6687)) or (layer0_outputs(3200)));
    outputs(3009) <= layer0_outputs(3467);
    outputs(3010) <= not(layer0_outputs(4173));
    outputs(3011) <= (layer0_outputs(3138)) and not (layer0_outputs(1026));
    outputs(3012) <= not(layer0_outputs(4414));
    outputs(3013) <= (layer0_outputs(3883)) and (layer0_outputs(2230));
    outputs(3014) <= not(layer0_outputs(378));
    outputs(3015) <= (layer0_outputs(5584)) or (layer0_outputs(4068));
    outputs(3016) <= not((layer0_outputs(4994)) xor (layer0_outputs(252)));
    outputs(3017) <= not(layer0_outputs(657)) or (layer0_outputs(7555));
    outputs(3018) <= (layer0_outputs(7171)) and not (layer0_outputs(4905));
    outputs(3019) <= layer0_outputs(5390);
    outputs(3020) <= layer0_outputs(4677);
    outputs(3021) <= not(layer0_outputs(6889));
    outputs(3022) <= not(layer0_outputs(1967));
    outputs(3023) <= layer0_outputs(5200);
    outputs(3024) <= not((layer0_outputs(1697)) or (layer0_outputs(7505)));
    outputs(3025) <= layer0_outputs(7582);
    outputs(3026) <= (layer0_outputs(3472)) and not (layer0_outputs(6577));
    outputs(3027) <= not(layer0_outputs(5330));
    outputs(3028) <= not(layer0_outputs(5412));
    outputs(3029) <= layer0_outputs(5266);
    outputs(3030) <= not((layer0_outputs(4356)) and (layer0_outputs(5147)));
    outputs(3031) <= (layer0_outputs(7561)) xor (layer0_outputs(996));
    outputs(3032) <= layer0_outputs(1478);
    outputs(3033) <= not(layer0_outputs(6767));
    outputs(3034) <= layer0_outputs(5097);
    outputs(3035) <= (layer0_outputs(3562)) xor (layer0_outputs(5319));
    outputs(3036) <= not(layer0_outputs(2106));
    outputs(3037) <= (layer0_outputs(69)) and (layer0_outputs(3527));
    outputs(3038) <= (layer0_outputs(1785)) or (layer0_outputs(3282));
    outputs(3039) <= not(layer0_outputs(824));
    outputs(3040) <= not((layer0_outputs(2027)) and (layer0_outputs(4061)));
    outputs(3041) <= not((layer0_outputs(4264)) or (layer0_outputs(439)));
    outputs(3042) <= layer0_outputs(4151);
    outputs(3043) <= (layer0_outputs(4907)) and (layer0_outputs(3435));
    outputs(3044) <= (layer0_outputs(2998)) xor (layer0_outputs(7652));
    outputs(3045) <= not(layer0_outputs(5173));
    outputs(3046) <= (layer0_outputs(7187)) or (layer0_outputs(2001));
    outputs(3047) <= not((layer0_outputs(7645)) or (layer0_outputs(3043)));
    outputs(3048) <= (layer0_outputs(8)) xor (layer0_outputs(3387));
    outputs(3049) <= not(layer0_outputs(2945));
    outputs(3050) <= (layer0_outputs(680)) and not (layer0_outputs(2267));
    outputs(3051) <= not((layer0_outputs(2439)) or (layer0_outputs(6610)));
    outputs(3052) <= (layer0_outputs(3237)) and not (layer0_outputs(2746));
    outputs(3053) <= layer0_outputs(3831);
    outputs(3054) <= not((layer0_outputs(7367)) xor (layer0_outputs(4377)));
    outputs(3055) <= layer0_outputs(4471);
    outputs(3056) <= layer0_outputs(7244);
    outputs(3057) <= (layer0_outputs(890)) and (layer0_outputs(7669));
    outputs(3058) <= not((layer0_outputs(6362)) or (layer0_outputs(5177)));
    outputs(3059) <= not(layer0_outputs(2694));
    outputs(3060) <= layer0_outputs(1260);
    outputs(3061) <= (layer0_outputs(597)) and (layer0_outputs(498));
    outputs(3062) <= (layer0_outputs(2477)) and not (layer0_outputs(1882));
    outputs(3063) <= not(layer0_outputs(5937));
    outputs(3064) <= (layer0_outputs(4488)) and (layer0_outputs(4583));
    outputs(3065) <= (layer0_outputs(2671)) xor (layer0_outputs(1678));
    outputs(3066) <= layer0_outputs(5326);
    outputs(3067) <= (layer0_outputs(6934)) and not (layer0_outputs(513));
    outputs(3068) <= not(layer0_outputs(1046));
    outputs(3069) <= not(layer0_outputs(3428));
    outputs(3070) <= (layer0_outputs(3443)) xor (layer0_outputs(1419));
    outputs(3071) <= not((layer0_outputs(6017)) xor (layer0_outputs(6759)));
    outputs(3072) <= not(layer0_outputs(6390));
    outputs(3073) <= not(layer0_outputs(1851));
    outputs(3074) <= layer0_outputs(3149);
    outputs(3075) <= not(layer0_outputs(7325));
    outputs(3076) <= (layer0_outputs(3125)) xor (layer0_outputs(7299));
    outputs(3077) <= layer0_outputs(3006);
    outputs(3078) <= layer0_outputs(1491);
    outputs(3079) <= not(layer0_outputs(2793));
    outputs(3080) <= layer0_outputs(1828);
    outputs(3081) <= not(layer0_outputs(3724));
    outputs(3082) <= (layer0_outputs(1281)) or (layer0_outputs(6736));
    outputs(3083) <= layer0_outputs(940);
    outputs(3084) <= not((layer0_outputs(1348)) or (layer0_outputs(3280)));
    outputs(3085) <= layer0_outputs(7475);
    outputs(3086) <= not(layer0_outputs(4070));
    outputs(3087) <= (layer0_outputs(5694)) xor (layer0_outputs(1407));
    outputs(3088) <= not((layer0_outputs(1043)) xor (layer0_outputs(2311)));
    outputs(3089) <= (layer0_outputs(6933)) and (layer0_outputs(3203));
    outputs(3090) <= not(layer0_outputs(6383));
    outputs(3091) <= not((layer0_outputs(6105)) and (layer0_outputs(2913)));
    outputs(3092) <= (layer0_outputs(2997)) xor (layer0_outputs(2599));
    outputs(3093) <= not((layer0_outputs(6844)) xor (layer0_outputs(853)));
    outputs(3094) <= layer0_outputs(7562);
    outputs(3095) <= not(layer0_outputs(5945));
    outputs(3096) <= layer0_outputs(4510);
    outputs(3097) <= not(layer0_outputs(713));
    outputs(3098) <= not((layer0_outputs(6774)) xor (layer0_outputs(726)));
    outputs(3099) <= not(layer0_outputs(3380));
    outputs(3100) <= layer0_outputs(1307);
    outputs(3101) <= not(layer0_outputs(5464));
    outputs(3102) <= not(layer0_outputs(2641));
    outputs(3103) <= not(layer0_outputs(5201)) or (layer0_outputs(5827));
    outputs(3104) <= not((layer0_outputs(493)) or (layer0_outputs(4022)));
    outputs(3105) <= (layer0_outputs(7344)) or (layer0_outputs(628));
    outputs(3106) <= not((layer0_outputs(2449)) xor (layer0_outputs(7653)));
    outputs(3107) <= (layer0_outputs(4715)) and not (layer0_outputs(732));
    outputs(3108) <= not(layer0_outputs(1464));
    outputs(3109) <= not(layer0_outputs(7050));
    outputs(3110) <= layer0_outputs(4370);
    outputs(3111) <= not(layer0_outputs(809)) or (layer0_outputs(363));
    outputs(3112) <= layer0_outputs(6680);
    outputs(3113) <= not((layer0_outputs(6918)) xor (layer0_outputs(7600)));
    outputs(3114) <= (layer0_outputs(5954)) xor (layer0_outputs(7282));
    outputs(3115) <= not(layer0_outputs(4128));
    outputs(3116) <= (layer0_outputs(5575)) and (layer0_outputs(2823));
    outputs(3117) <= not(layer0_outputs(4966));
    outputs(3118) <= (layer0_outputs(6097)) and (layer0_outputs(4684));
    outputs(3119) <= not(layer0_outputs(6777));
    outputs(3120) <= layer0_outputs(5168);
    outputs(3121) <= layer0_outputs(4475);
    outputs(3122) <= layer0_outputs(509);
    outputs(3123) <= not(layer0_outputs(4897));
    outputs(3124) <= not(layer0_outputs(7158));
    outputs(3125) <= layer0_outputs(2820);
    outputs(3126) <= not(layer0_outputs(216));
    outputs(3127) <= (layer0_outputs(2828)) xor (layer0_outputs(5134));
    outputs(3128) <= (layer0_outputs(653)) and not (layer0_outputs(1835));
    outputs(3129) <= (layer0_outputs(5428)) and not (layer0_outputs(4245));
    outputs(3130) <= not((layer0_outputs(5501)) or (layer0_outputs(6786)));
    outputs(3131) <= (layer0_outputs(4212)) and (layer0_outputs(224));
    outputs(3132) <= not(layer0_outputs(4070)) or (layer0_outputs(4400));
    outputs(3133) <= not((layer0_outputs(3133)) or (layer0_outputs(2711)));
    outputs(3134) <= not(layer0_outputs(2588)) or (layer0_outputs(6189));
    outputs(3135) <= (layer0_outputs(5739)) xor (layer0_outputs(6299));
    outputs(3136) <= not(layer0_outputs(3013));
    outputs(3137) <= (layer0_outputs(5986)) xor (layer0_outputs(4419));
    outputs(3138) <= not((layer0_outputs(2678)) and (layer0_outputs(6809)));
    outputs(3139) <= not(layer0_outputs(1426));
    outputs(3140) <= not((layer0_outputs(3825)) or (layer0_outputs(2203)));
    outputs(3141) <= (layer0_outputs(47)) xor (layer0_outputs(6328));
    outputs(3142) <= (layer0_outputs(4242)) and (layer0_outputs(1946));
    outputs(3143) <= not((layer0_outputs(4882)) or (layer0_outputs(2358)));
    outputs(3144) <= not(layer0_outputs(5880));
    outputs(3145) <= (layer0_outputs(7283)) xor (layer0_outputs(6351));
    outputs(3146) <= not(layer0_outputs(3228));
    outputs(3147) <= layer0_outputs(975);
    outputs(3148) <= not(layer0_outputs(2681));
    outputs(3149) <= (layer0_outputs(4428)) xor (layer0_outputs(5213));
    outputs(3150) <= (layer0_outputs(2610)) and (layer0_outputs(7483));
    outputs(3151) <= (layer0_outputs(4168)) and not (layer0_outputs(4071));
    outputs(3152) <= not(layer0_outputs(4896));
    outputs(3153) <= not(layer0_outputs(3005));
    outputs(3154) <= not(layer0_outputs(5411));
    outputs(3155) <= not(layer0_outputs(3441));
    outputs(3156) <= layer0_outputs(5211);
    outputs(3157) <= not((layer0_outputs(7099)) or (layer0_outputs(383)));
    outputs(3158) <= (layer0_outputs(6782)) and not (layer0_outputs(5574));
    outputs(3159) <= not((layer0_outputs(6143)) xor (layer0_outputs(2052)));
    outputs(3160) <= layer0_outputs(6941);
    outputs(3161) <= (layer0_outputs(1415)) xor (layer0_outputs(5728));
    outputs(3162) <= layer0_outputs(5626);
    outputs(3163) <= not(layer0_outputs(6858));
    outputs(3164) <= not(layer0_outputs(2353));
    outputs(3165) <= not((layer0_outputs(3281)) xor (layer0_outputs(5809)));
    outputs(3166) <= (layer0_outputs(2406)) and not (layer0_outputs(751));
    outputs(3167) <= not((layer0_outputs(3311)) or (layer0_outputs(5110)));
    outputs(3168) <= (layer0_outputs(4298)) and (layer0_outputs(7663));
    outputs(3169) <= not(layer0_outputs(4368));
    outputs(3170) <= (layer0_outputs(7515)) or (layer0_outputs(3621));
    outputs(3171) <= layer0_outputs(3050);
    outputs(3172) <= layer0_outputs(3252);
    outputs(3173) <= not((layer0_outputs(4917)) or (layer0_outputs(3858)));
    outputs(3174) <= not(layer0_outputs(4983));
    outputs(3175) <= (layer0_outputs(7618)) xor (layer0_outputs(116));
    outputs(3176) <= (layer0_outputs(4657)) and not (layer0_outputs(6449));
    outputs(3177) <= not(layer0_outputs(819)) or (layer0_outputs(1681));
    outputs(3178) <= not((layer0_outputs(5641)) and (layer0_outputs(40)));
    outputs(3179) <= not(layer0_outputs(4390));
    outputs(3180) <= not(layer0_outputs(6815)) or (layer0_outputs(3054));
    outputs(3181) <= layer0_outputs(1170);
    outputs(3182) <= not(layer0_outputs(4995)) or (layer0_outputs(1191));
    outputs(3183) <= (layer0_outputs(2792)) and not (layer0_outputs(5257));
    outputs(3184) <= not(layer0_outputs(3581));
    outputs(3185) <= not((layer0_outputs(4099)) xor (layer0_outputs(5546)));
    outputs(3186) <= not(layer0_outputs(7252));
    outputs(3187) <= layer0_outputs(460);
    outputs(3188) <= (layer0_outputs(7101)) xor (layer0_outputs(3427));
    outputs(3189) <= not((layer0_outputs(875)) xor (layer0_outputs(6069)));
    outputs(3190) <= (layer0_outputs(416)) and not (layer0_outputs(1138));
    outputs(3191) <= (layer0_outputs(3577)) and not (layer0_outputs(5917));
    outputs(3192) <= layer0_outputs(4404);
    outputs(3193) <= not(layer0_outputs(2510)) or (layer0_outputs(1639));
    outputs(3194) <= not(layer0_outputs(179));
    outputs(3195) <= (layer0_outputs(3501)) and (layer0_outputs(4268));
    outputs(3196) <= (layer0_outputs(3723)) and not (layer0_outputs(845));
    outputs(3197) <= not(layer0_outputs(1960));
    outputs(3198) <= (layer0_outputs(233)) xor (layer0_outputs(273));
    outputs(3199) <= not((layer0_outputs(5442)) xor (layer0_outputs(6866)));
    outputs(3200) <= layer0_outputs(6432);
    outputs(3201) <= layer0_outputs(3844);
    outputs(3202) <= not((layer0_outputs(4844)) xor (layer0_outputs(4286)));
    outputs(3203) <= layer0_outputs(3976);
    outputs(3204) <= (layer0_outputs(274)) and not (layer0_outputs(2171));
    outputs(3205) <= (layer0_outputs(19)) and (layer0_outputs(3552));
    outputs(3206) <= not(layer0_outputs(5797));
    outputs(3207) <= not(layer0_outputs(7569));
    outputs(3208) <= not(layer0_outputs(5358)) or (layer0_outputs(768));
    outputs(3209) <= layer0_outputs(4822);
    outputs(3210) <= (layer0_outputs(7339)) or (layer0_outputs(3691));
    outputs(3211) <= not((layer0_outputs(601)) and (layer0_outputs(113)));
    outputs(3212) <= not(layer0_outputs(7256));
    outputs(3213) <= layer0_outputs(5673);
    outputs(3214) <= (layer0_outputs(1606)) and not (layer0_outputs(2011));
    outputs(3215) <= not(layer0_outputs(5554));
    outputs(3216) <= layer0_outputs(3950);
    outputs(3217) <= layer0_outputs(5049);
    outputs(3218) <= not(layer0_outputs(3189));
    outputs(3219) <= layer0_outputs(2082);
    outputs(3220) <= (layer0_outputs(2755)) and (layer0_outputs(5284));
    outputs(3221) <= layer0_outputs(4370);
    outputs(3222) <= layer0_outputs(3461);
    outputs(3223) <= layer0_outputs(7153);
    outputs(3224) <= (layer0_outputs(6408)) xor (layer0_outputs(221));
    outputs(3225) <= layer0_outputs(5883);
    outputs(3226) <= not((layer0_outputs(5091)) xor (layer0_outputs(3385)));
    outputs(3227) <= layer0_outputs(3305);
    outputs(3228) <= layer0_outputs(2504);
    outputs(3229) <= (layer0_outputs(7506)) and not (layer0_outputs(3218));
    outputs(3230) <= (layer0_outputs(3874)) and not (layer0_outputs(7583));
    outputs(3231) <= layer0_outputs(4641);
    outputs(3232) <= (layer0_outputs(7677)) and (layer0_outputs(4679));
    outputs(3233) <= (layer0_outputs(2093)) and not (layer0_outputs(2550));
    outputs(3234) <= layer0_outputs(3122);
    outputs(3235) <= layer0_outputs(7285);
    outputs(3236) <= layer0_outputs(4238);
    outputs(3237) <= not((layer0_outputs(1466)) xor (layer0_outputs(757)));
    outputs(3238) <= not(layer0_outputs(5485));
    outputs(3239) <= layer0_outputs(2388);
    outputs(3240) <= not((layer0_outputs(7365)) or (layer0_outputs(4424)));
    outputs(3241) <= not((layer0_outputs(2440)) xor (layer0_outputs(5245)));
    outputs(3242) <= (layer0_outputs(2430)) and not (layer0_outputs(7526));
    outputs(3243) <= not(layer0_outputs(1717));
    outputs(3244) <= not(layer0_outputs(2369));
    outputs(3245) <= (layer0_outputs(3499)) and not (layer0_outputs(2970));
    outputs(3246) <= not(layer0_outputs(865));
    outputs(3247) <= not(layer0_outputs(2213));
    outputs(3248) <= not(layer0_outputs(6100));
    outputs(3249) <= layer0_outputs(3895);
    outputs(3250) <= (layer0_outputs(759)) and not (layer0_outputs(5065));
    outputs(3251) <= layer0_outputs(1411);
    outputs(3252) <= not((layer0_outputs(5239)) or (layer0_outputs(5803)));
    outputs(3253) <= (layer0_outputs(5692)) or (layer0_outputs(5441));
    outputs(3254) <= not(layer0_outputs(6870));
    outputs(3255) <= (layer0_outputs(5777)) and (layer0_outputs(6733));
    outputs(3256) <= (layer0_outputs(3987)) and not (layer0_outputs(6459));
    outputs(3257) <= layer0_outputs(3290);
    outputs(3258) <= (layer0_outputs(2580)) and not (layer0_outputs(5107));
    outputs(3259) <= not(layer0_outputs(6465));
    outputs(3260) <= (layer0_outputs(393)) and not (layer0_outputs(4287));
    outputs(3261) <= (layer0_outputs(157)) and not (layer0_outputs(5631));
    outputs(3262) <= layer0_outputs(5259);
    outputs(3263) <= not(layer0_outputs(4546));
    outputs(3264) <= layer0_outputs(7152);
    outputs(3265) <= not(layer0_outputs(2632));
    outputs(3266) <= (layer0_outputs(2750)) and not (layer0_outputs(2083));
    outputs(3267) <= not((layer0_outputs(3011)) or (layer0_outputs(6975)));
    outputs(3268) <= not((layer0_outputs(7127)) xor (layer0_outputs(6855)));
    outputs(3269) <= (layer0_outputs(1930)) and not (layer0_outputs(5172));
    outputs(3270) <= layer0_outputs(5709);
    outputs(3271) <= not(layer0_outputs(286));
    outputs(3272) <= (layer0_outputs(7375)) xor (layer0_outputs(4329));
    outputs(3273) <= (layer0_outputs(7135)) and not (layer0_outputs(1432));
    outputs(3274) <= not(layer0_outputs(708));
    outputs(3275) <= layer0_outputs(3820);
    outputs(3276) <= not(layer0_outputs(7581));
    outputs(3277) <= (layer0_outputs(158)) xor (layer0_outputs(3030));
    outputs(3278) <= (layer0_outputs(3817)) and not (layer0_outputs(4139));
    outputs(3279) <= (layer0_outputs(5530)) and not (layer0_outputs(4709));
    outputs(3280) <= not((layer0_outputs(7379)) xor (layer0_outputs(2075)));
    outputs(3281) <= not(layer0_outputs(4897));
    outputs(3282) <= layer0_outputs(1117);
    outputs(3283) <= (layer0_outputs(1179)) and not (layer0_outputs(147));
    outputs(3284) <= not((layer0_outputs(7361)) xor (layer0_outputs(1253)));
    outputs(3285) <= not(layer0_outputs(3116)) or (layer0_outputs(5944));
    outputs(3286) <= layer0_outputs(76);
    outputs(3287) <= layer0_outputs(2715);
    outputs(3288) <= not((layer0_outputs(5826)) or (layer0_outputs(6311)));
    outputs(3289) <= layer0_outputs(7523);
    outputs(3290) <= not((layer0_outputs(6653)) or (layer0_outputs(645)));
    outputs(3291) <= layer0_outputs(1509);
    outputs(3292) <= not((layer0_outputs(142)) or (layer0_outputs(146)));
    outputs(3293) <= not(layer0_outputs(4422));
    outputs(3294) <= not(layer0_outputs(2658));
    outputs(3295) <= not(layer0_outputs(1493));
    outputs(3296) <= not(layer0_outputs(5961));
    outputs(3297) <= layer0_outputs(104);
    outputs(3298) <= layer0_outputs(1752);
    outputs(3299) <= layer0_outputs(2574);
    outputs(3300) <= not(layer0_outputs(2031));
    outputs(3301) <= layer0_outputs(5968);
    outputs(3302) <= layer0_outputs(6856);
    outputs(3303) <= not(layer0_outputs(6534)) or (layer0_outputs(1015));
    outputs(3304) <= not(layer0_outputs(6752));
    outputs(3305) <= (layer0_outputs(99)) and (layer0_outputs(5338));
    outputs(3306) <= not(layer0_outputs(2946));
    outputs(3307) <= (layer0_outputs(5516)) and not (layer0_outputs(4866));
    outputs(3308) <= layer0_outputs(378);
    outputs(3309) <= layer0_outputs(5788);
    outputs(3310) <= not(layer0_outputs(4391));
    outputs(3311) <= not(layer0_outputs(5321));
    outputs(3312) <= not(layer0_outputs(3331));
    outputs(3313) <= not(layer0_outputs(4862));
    outputs(3314) <= not((layer0_outputs(3105)) xor (layer0_outputs(24)));
    outputs(3315) <= layer0_outputs(6312);
    outputs(3316) <= layer0_outputs(7546);
    outputs(3317) <= (layer0_outputs(5145)) and (layer0_outputs(2143));
    outputs(3318) <= (layer0_outputs(4578)) xor (layer0_outputs(2080));
    outputs(3319) <= (layer0_outputs(3246)) xor (layer0_outputs(1795));
    outputs(3320) <= (layer0_outputs(7138)) and not (layer0_outputs(1456));
    outputs(3321) <= not(layer0_outputs(7372));
    outputs(3322) <= not(layer0_outputs(1083));
    outputs(3323) <= layer0_outputs(1813);
    outputs(3324) <= not(layer0_outputs(5249)) or (layer0_outputs(4037));
    outputs(3325) <= (layer0_outputs(650)) and not (layer0_outputs(5465));
    outputs(3326) <= layer0_outputs(7028);
    outputs(3327) <= layer0_outputs(3017);
    outputs(3328) <= layer0_outputs(4441);
    outputs(3329) <= layer0_outputs(3548);
    outputs(3330) <= not(layer0_outputs(3974));
    outputs(3331) <= (layer0_outputs(6222)) xor (layer0_outputs(2666));
    outputs(3332) <= (layer0_outputs(1813)) and not (layer0_outputs(97));
    outputs(3333) <= not(layer0_outputs(5754));
    outputs(3334) <= (layer0_outputs(3580)) and not (layer0_outputs(391));
    outputs(3335) <= (layer0_outputs(1171)) and not (layer0_outputs(3026));
    outputs(3336) <= layer0_outputs(652);
    outputs(3337) <= (layer0_outputs(5934)) and (layer0_outputs(6016));
    outputs(3338) <= (layer0_outputs(7173)) and not (layer0_outputs(440));
    outputs(3339) <= not((layer0_outputs(6153)) or (layer0_outputs(5389)));
    outputs(3340) <= not(layer0_outputs(3251));
    outputs(3341) <= not(layer0_outputs(3479)) or (layer0_outputs(1742));
    outputs(3342) <= not((layer0_outputs(634)) or (layer0_outputs(5651)));
    outputs(3343) <= layer0_outputs(6989);
    outputs(3344) <= not(layer0_outputs(5670)) or (layer0_outputs(7359));
    outputs(3345) <= layer0_outputs(4136);
    outputs(3346) <= not(layer0_outputs(1382));
    outputs(3347) <= layer0_outputs(3557);
    outputs(3348) <= layer0_outputs(3953);
    outputs(3349) <= layer0_outputs(6976);
    outputs(3350) <= layer0_outputs(3335);
    outputs(3351) <= (layer0_outputs(1889)) xor (layer0_outputs(4105));
    outputs(3352) <= layer0_outputs(3410);
    outputs(3353) <= not((layer0_outputs(1617)) xor (layer0_outputs(1029)));
    outputs(3354) <= not(layer0_outputs(3937));
    outputs(3355) <= layer0_outputs(3970);
    outputs(3356) <= not(layer0_outputs(2249));
    outputs(3357) <= (layer0_outputs(4744)) and not (layer0_outputs(2429));
    outputs(3358) <= not(layer0_outputs(522));
    outputs(3359) <= not((layer0_outputs(4935)) xor (layer0_outputs(237)));
    outputs(3360) <= not(layer0_outputs(7572));
    outputs(3361) <= (layer0_outputs(513)) or (layer0_outputs(4171));
    outputs(3362) <= (layer0_outputs(3953)) and (layer0_outputs(3035));
    outputs(3363) <= layer0_outputs(4134);
    outputs(3364) <= not(layer0_outputs(4816));
    outputs(3365) <= not(layer0_outputs(1083));
    outputs(3366) <= not(layer0_outputs(4834));
    outputs(3367) <= not(layer0_outputs(2001));
    outputs(3368) <= not(layer0_outputs(5920)) or (layer0_outputs(3310));
    outputs(3369) <= not(layer0_outputs(4622));
    outputs(3370) <= not(layer0_outputs(5752));
    outputs(3371) <= not(layer0_outputs(2038));
    outputs(3372) <= (layer0_outputs(2419)) xor (layer0_outputs(6998));
    outputs(3373) <= layer0_outputs(4602);
    outputs(3374) <= layer0_outputs(1541);
    outputs(3375) <= not(layer0_outputs(4603));
    outputs(3376) <= (layer0_outputs(4312)) xor (layer0_outputs(6163));
    outputs(3377) <= (layer0_outputs(4943)) and not (layer0_outputs(7201));
    outputs(3378) <= not(layer0_outputs(4667));
    outputs(3379) <= layer0_outputs(3782);
    outputs(3380) <= not(layer0_outputs(486));
    outputs(3381) <= layer0_outputs(6356);
    outputs(3382) <= not(layer0_outputs(2959));
    outputs(3383) <= not(layer0_outputs(4816));
    outputs(3384) <= (layer0_outputs(6169)) and (layer0_outputs(5005));
    outputs(3385) <= not(layer0_outputs(3041));
    outputs(3386) <= not(layer0_outputs(3129));
    outputs(3387) <= layer0_outputs(2102);
    outputs(3388) <= (layer0_outputs(2595)) and not (layer0_outputs(6754));
    outputs(3389) <= not((layer0_outputs(7326)) xor (layer0_outputs(4277)));
    outputs(3390) <= not((layer0_outputs(1823)) xor (layer0_outputs(4500)));
    outputs(3391) <= not(layer0_outputs(6152));
    outputs(3392) <= layer0_outputs(5830);
    outputs(3393) <= layer0_outputs(904);
    outputs(3394) <= not(layer0_outputs(540));
    outputs(3395) <= (layer0_outputs(780)) or (layer0_outputs(3206));
    outputs(3396) <= not((layer0_outputs(3364)) or (layer0_outputs(5356)));
    outputs(3397) <= not(layer0_outputs(587));
    outputs(3398) <= (layer0_outputs(6519)) or (layer0_outputs(421));
    outputs(3399) <= not(layer0_outputs(7404));
    outputs(3400) <= not((layer0_outputs(2362)) and (layer0_outputs(1739)));
    outputs(3401) <= (layer0_outputs(6705)) and not (layer0_outputs(1353));
    outputs(3402) <= not(layer0_outputs(4266));
    outputs(3403) <= (layer0_outputs(4018)) xor (layer0_outputs(7197));
    outputs(3404) <= (layer0_outputs(4374)) and not (layer0_outputs(5092));
    outputs(3405) <= not((layer0_outputs(3003)) or (layer0_outputs(6012)));
    outputs(3406) <= layer0_outputs(112);
    outputs(3407) <= layer0_outputs(6456);
    outputs(3408) <= not(layer0_outputs(2167));
    outputs(3409) <= layer0_outputs(4466);
    outputs(3410) <= layer0_outputs(705);
    outputs(3411) <= (layer0_outputs(3415)) and not (layer0_outputs(3519));
    outputs(3412) <= (layer0_outputs(7013)) xor (layer0_outputs(5005));
    outputs(3413) <= not(layer0_outputs(6112));
    outputs(3414) <= (layer0_outputs(3767)) xor (layer0_outputs(5376));
    outputs(3415) <= not(layer0_outputs(6634));
    outputs(3416) <= (layer0_outputs(2807)) and not (layer0_outputs(452));
    outputs(3417) <= (layer0_outputs(650)) and not (layer0_outputs(3507));
    outputs(3418) <= (layer0_outputs(3288)) and not (layer0_outputs(55));
    outputs(3419) <= not(layer0_outputs(3502));
    outputs(3420) <= (layer0_outputs(6769)) and (layer0_outputs(3517));
    outputs(3421) <= not(layer0_outputs(2324));
    outputs(3422) <= (layer0_outputs(2904)) xor (layer0_outputs(5037));
    outputs(3423) <= (layer0_outputs(6973)) and (layer0_outputs(6113));
    outputs(3424) <= (layer0_outputs(4203)) and not (layer0_outputs(4164));
    outputs(3425) <= (layer0_outputs(655)) xor (layer0_outputs(5713));
    outputs(3426) <= (layer0_outputs(5726)) xor (layer0_outputs(5226));
    outputs(3427) <= layer0_outputs(1034);
    outputs(3428) <= (layer0_outputs(1554)) and not (layer0_outputs(5660));
    outputs(3429) <= not((layer0_outputs(3653)) xor (layer0_outputs(981)));
    outputs(3430) <= (layer0_outputs(6631)) and not (layer0_outputs(5537));
    outputs(3431) <= not(layer0_outputs(6417));
    outputs(3432) <= not(layer0_outputs(1243));
    outputs(3433) <= layer0_outputs(986);
    outputs(3434) <= not((layer0_outputs(4093)) xor (layer0_outputs(1633)));
    outputs(3435) <= not(layer0_outputs(175));
    outputs(3436) <= layer0_outputs(5653);
    outputs(3437) <= not((layer0_outputs(6102)) or (layer0_outputs(5317)));
    outputs(3438) <= (layer0_outputs(4869)) xor (layer0_outputs(6444));
    outputs(3439) <= not(layer0_outputs(5222));
    outputs(3440) <= not((layer0_outputs(3806)) xor (layer0_outputs(7187)));
    outputs(3441) <= layer0_outputs(140);
    outputs(3442) <= not(layer0_outputs(1488));
    outputs(3443) <= layer0_outputs(1383);
    outputs(3444) <= layer0_outputs(7371);
    outputs(3445) <= layer0_outputs(1091);
    outputs(3446) <= not(layer0_outputs(6859)) or (layer0_outputs(499));
    outputs(3447) <= not((layer0_outputs(1392)) or (layer0_outputs(1201)));
    outputs(3448) <= not(layer0_outputs(1168));
    outputs(3449) <= layer0_outputs(5029);
    outputs(3450) <= not(layer0_outputs(7351));
    outputs(3451) <= (layer0_outputs(3982)) and not (layer0_outputs(6329));
    outputs(3452) <= layer0_outputs(669);
    outputs(3453) <= (layer0_outputs(1210)) xor (layer0_outputs(395));
    outputs(3454) <= not(layer0_outputs(1311));
    outputs(3455) <= not(layer0_outputs(1666));
    outputs(3456) <= not(layer0_outputs(2304)) or (layer0_outputs(1900));
    outputs(3457) <= layer0_outputs(2082);
    outputs(3458) <= not((layer0_outputs(2650)) and (layer0_outputs(3351)));
    outputs(3459) <= not(layer0_outputs(3613));
    outputs(3460) <= not(layer0_outputs(3081));
    outputs(3461) <= not(layer0_outputs(7617));
    outputs(3462) <= (layer0_outputs(5124)) or (layer0_outputs(5018));
    outputs(3463) <= layer0_outputs(934);
    outputs(3464) <= (layer0_outputs(3638)) or (layer0_outputs(325));
    outputs(3465) <= layer0_outputs(4957);
    outputs(3466) <= not(layer0_outputs(7232)) or (layer0_outputs(2377));
    outputs(3467) <= (layer0_outputs(6639)) and not (layer0_outputs(3680));
    outputs(3468) <= not(layer0_outputs(4601));
    outputs(3469) <= not((layer0_outputs(3460)) or (layer0_outputs(7039)));
    outputs(3470) <= layer0_outputs(3593);
    outputs(3471) <= layer0_outputs(3708);
    outputs(3472) <= not(layer0_outputs(2896));
    outputs(3473) <= not((layer0_outputs(7400)) xor (layer0_outputs(1834)));
    outputs(3474) <= not((layer0_outputs(4351)) or (layer0_outputs(230)));
    outputs(3475) <= not((layer0_outputs(5195)) or (layer0_outputs(7331)));
    outputs(3476) <= not((layer0_outputs(4537)) xor (layer0_outputs(6840)));
    outputs(3477) <= (layer0_outputs(5922)) and not (layer0_outputs(5423));
    outputs(3478) <= not((layer0_outputs(736)) xor (layer0_outputs(1166)));
    outputs(3479) <= (layer0_outputs(5385)) and not (layer0_outputs(2983));
    outputs(3480) <= layer0_outputs(1102);
    outputs(3481) <= layer0_outputs(2186);
    outputs(3482) <= not(layer0_outputs(725));
    outputs(3483) <= layer0_outputs(5849);
    outputs(3484) <= not((layer0_outputs(1916)) xor (layer0_outputs(6079)));
    outputs(3485) <= layer0_outputs(4677);
    outputs(3486) <= not(layer0_outputs(3471));
    outputs(3487) <= layer0_outputs(6778);
    outputs(3488) <= not(layer0_outputs(7154));
    outputs(3489) <= layer0_outputs(2685);
    outputs(3490) <= layer0_outputs(5425);
    outputs(3491) <= (layer0_outputs(2668)) and not (layer0_outputs(6584));
    outputs(3492) <= (layer0_outputs(2183)) and not (layer0_outputs(2851));
    outputs(3493) <= not(layer0_outputs(232)) or (layer0_outputs(1526));
    outputs(3494) <= not(layer0_outputs(4338));
    outputs(3495) <= not(layer0_outputs(599));
    outputs(3496) <= not(layer0_outputs(4665));
    outputs(3497) <= (layer0_outputs(3673)) and (layer0_outputs(178));
    outputs(3498) <= layer0_outputs(3291);
    outputs(3499) <= layer0_outputs(6154);
    outputs(3500) <= not(layer0_outputs(1422)) or (layer0_outputs(5217));
    outputs(3501) <= not(layer0_outputs(2054));
    outputs(3502) <= layer0_outputs(1016);
    outputs(3503) <= not(layer0_outputs(429));
    outputs(3504) <= not((layer0_outputs(1735)) or (layer0_outputs(7404)));
    outputs(3505) <= (layer0_outputs(1232)) and (layer0_outputs(4572));
    outputs(3506) <= not(layer0_outputs(7124)) or (layer0_outputs(6639));
    outputs(3507) <= (layer0_outputs(4637)) or (layer0_outputs(2201));
    outputs(3508) <= layer0_outputs(2243);
    outputs(3509) <= layer0_outputs(924);
    outputs(3510) <= layer0_outputs(3815);
    outputs(3511) <= not(layer0_outputs(2030));
    outputs(3512) <= not(layer0_outputs(6455));
    outputs(3513) <= layer0_outputs(1970);
    outputs(3514) <= not(layer0_outputs(3005));
    outputs(3515) <= not(layer0_outputs(5114));
    outputs(3516) <= (layer0_outputs(3494)) and not (layer0_outputs(4152));
    outputs(3517) <= not(layer0_outputs(194));
    outputs(3518) <= not(layer0_outputs(1678));
    outputs(3519) <= (layer0_outputs(5621)) and not (layer0_outputs(1485));
    outputs(3520) <= layer0_outputs(5761);
    outputs(3521) <= not((layer0_outputs(3662)) xor (layer0_outputs(6186)));
    outputs(3522) <= not(layer0_outputs(5178));
    outputs(3523) <= not(layer0_outputs(155)) or (layer0_outputs(1643));
    outputs(3524) <= layer0_outputs(5313);
    outputs(3525) <= layer0_outputs(3211);
    outputs(3526) <= (layer0_outputs(388)) and (layer0_outputs(5655));
    outputs(3527) <= layer0_outputs(1912);
    outputs(3528) <= layer0_outputs(6116);
    outputs(3529) <= not(layer0_outputs(7150));
    outputs(3530) <= layer0_outputs(4849);
    outputs(3531) <= not((layer0_outputs(6354)) xor (layer0_outputs(85)));
    outputs(3532) <= not(layer0_outputs(5794));
    outputs(3533) <= layer0_outputs(6298);
    outputs(3534) <= (layer0_outputs(1535)) or (layer0_outputs(1624));
    outputs(3535) <= layer0_outputs(1569);
    outputs(3536) <= not(layer0_outputs(3853));
    outputs(3537) <= not((layer0_outputs(2149)) xor (layer0_outputs(4485)));
    outputs(3538) <= (layer0_outputs(1905)) and (layer0_outputs(1668));
    outputs(3539) <= layer0_outputs(3109);
    outputs(3540) <= not((layer0_outputs(1060)) and (layer0_outputs(4850)));
    outputs(3541) <= not((layer0_outputs(1031)) xor (layer0_outputs(1125)));
    outputs(3542) <= not((layer0_outputs(6556)) or (layer0_outputs(2670)));
    outputs(3543) <= layer0_outputs(2995);
    outputs(3544) <= (layer0_outputs(7406)) and (layer0_outputs(7532));
    outputs(3545) <= not(layer0_outputs(6683));
    outputs(3546) <= not(layer0_outputs(1901));
    outputs(3547) <= not(layer0_outputs(2716));
    outputs(3548) <= (layer0_outputs(5320)) and (layer0_outputs(3522));
    outputs(3549) <= (layer0_outputs(1423)) xor (layer0_outputs(1193));
    outputs(3550) <= (layer0_outputs(6132)) xor (layer0_outputs(6552));
    outputs(3551) <= layer0_outputs(3598);
    outputs(3552) <= layer0_outputs(5685);
    outputs(3553) <= not(layer0_outputs(3812));
    outputs(3554) <= not(layer0_outputs(7256));
    outputs(3555) <= not(layer0_outputs(916));
    outputs(3556) <= not(layer0_outputs(7376));
    outputs(3557) <= not((layer0_outputs(6718)) xor (layer0_outputs(4536)));
    outputs(3558) <= not(layer0_outputs(7097));
    outputs(3559) <= not(layer0_outputs(1386));
    outputs(3560) <= layer0_outputs(6704);
    outputs(3561) <= (layer0_outputs(1545)) and (layer0_outputs(5862));
    outputs(3562) <= layer0_outputs(2214);
    outputs(3563) <= not((layer0_outputs(805)) or (layer0_outputs(5866)));
    outputs(3564) <= (layer0_outputs(1820)) and (layer0_outputs(5658));
    outputs(3565) <= not(layer0_outputs(1401));
    outputs(3566) <= (layer0_outputs(5854)) and (layer0_outputs(3246));
    outputs(3567) <= not(layer0_outputs(6511));
    outputs(3568) <= (layer0_outputs(5243)) xor (layer0_outputs(7210));
    outputs(3569) <= not((layer0_outputs(6788)) xor (layer0_outputs(7349)));
    outputs(3570) <= not(layer0_outputs(7009)) or (layer0_outputs(6215));
    outputs(3571) <= not(layer0_outputs(664));
    outputs(3572) <= not(layer0_outputs(4539));
    outputs(3573) <= not(layer0_outputs(14));
    outputs(3574) <= not(layer0_outputs(1484));
    outputs(3575) <= layer0_outputs(6438);
    outputs(3576) <= (layer0_outputs(1392)) xor (layer0_outputs(401));
    outputs(3577) <= not(layer0_outputs(4315));
    outputs(3578) <= layer0_outputs(4466);
    outputs(3579) <= not((layer0_outputs(982)) xor (layer0_outputs(3841)));
    outputs(3580) <= not(layer0_outputs(6321));
    outputs(3581) <= layer0_outputs(6839);
    outputs(3582) <= not((layer0_outputs(3119)) or (layer0_outputs(680)));
    outputs(3583) <= not(layer0_outputs(5942)) or (layer0_outputs(3880));
    outputs(3584) <= not(layer0_outputs(6291));
    outputs(3585) <= layer0_outputs(5484);
    outputs(3586) <= not(layer0_outputs(6726));
    outputs(3587) <= not(layer0_outputs(7653));
    outputs(3588) <= layer0_outputs(7078);
    outputs(3589) <= not((layer0_outputs(7498)) xor (layer0_outputs(6982)));
    outputs(3590) <= not(layer0_outputs(7484));
    outputs(3591) <= not((layer0_outputs(6160)) or (layer0_outputs(5354)));
    outputs(3592) <= not(layer0_outputs(2682));
    outputs(3593) <= layer0_outputs(7643);
    outputs(3594) <= (layer0_outputs(3561)) and (layer0_outputs(5695));
    outputs(3595) <= not((layer0_outputs(6757)) xor (layer0_outputs(5341)));
    outputs(3596) <= layer0_outputs(3149);
    outputs(3597) <= layer0_outputs(7018);
    outputs(3598) <= layer0_outputs(5874);
    outputs(3599) <= layer0_outputs(7047);
    outputs(3600) <= layer0_outputs(5111);
    outputs(3601) <= not(layer0_outputs(1995));
    outputs(3602) <= (layer0_outputs(3294)) and (layer0_outputs(2819));
    outputs(3603) <= not((layer0_outputs(713)) or (layer0_outputs(504)));
    outputs(3604) <= not(layer0_outputs(4309));
    outputs(3605) <= not((layer0_outputs(2663)) xor (layer0_outputs(5618)));
    outputs(3606) <= not((layer0_outputs(4166)) xor (layer0_outputs(6023)));
    outputs(3607) <= not(layer0_outputs(5099)) or (layer0_outputs(7544));
    outputs(3608) <= (layer0_outputs(3802)) and not (layer0_outputs(1848));
    outputs(3609) <= not((layer0_outputs(5393)) and (layer0_outputs(4333)));
    outputs(3610) <= layer0_outputs(6045);
    outputs(3611) <= not((layer0_outputs(7041)) or (layer0_outputs(1241)));
    outputs(3612) <= (layer0_outputs(4380)) or (layer0_outputs(4723));
    outputs(3613) <= (layer0_outputs(1329)) and (layer0_outputs(5989));
    outputs(3614) <= not((layer0_outputs(2845)) and (layer0_outputs(2031)));
    outputs(3615) <= not(layer0_outputs(7302));
    outputs(3616) <= layer0_outputs(4657);
    outputs(3617) <= not(layer0_outputs(5577));
    outputs(3618) <= not(layer0_outputs(1169));
    outputs(3619) <= not(layer0_outputs(6382)) or (layer0_outputs(1547));
    outputs(3620) <= layer0_outputs(6188);
    outputs(3621) <= (layer0_outputs(2830)) and (layer0_outputs(6644));
    outputs(3622) <= layer0_outputs(3626);
    outputs(3623) <= not((layer0_outputs(5913)) or (layer0_outputs(6400)));
    outputs(3624) <= layer0_outputs(7215);
    outputs(3625) <= not((layer0_outputs(6580)) xor (layer0_outputs(2300)));
    outputs(3626) <= (layer0_outputs(6678)) and not (layer0_outputs(2485));
    outputs(3627) <= not((layer0_outputs(163)) or (layer0_outputs(6626)));
    outputs(3628) <= (layer0_outputs(218)) xor (layer0_outputs(6964));
    outputs(3629) <= layer0_outputs(6333);
    outputs(3630) <= not((layer0_outputs(6701)) xor (layer0_outputs(6512)));
    outputs(3631) <= layer0_outputs(6579);
    outputs(3632) <= not(layer0_outputs(7500)) or (layer0_outputs(7285));
    outputs(3633) <= layer0_outputs(3285);
    outputs(3634) <= not(layer0_outputs(2968));
    outputs(3635) <= layer0_outputs(4544);
    outputs(3636) <= layer0_outputs(5348);
    outputs(3637) <= not(layer0_outputs(1128));
    outputs(3638) <= layer0_outputs(1044);
    outputs(3639) <= (layer0_outputs(1996)) and (layer0_outputs(2806));
    outputs(3640) <= not(layer0_outputs(5657));
    outputs(3641) <= (layer0_outputs(7193)) xor (layer0_outputs(172));
    outputs(3642) <= not(layer0_outputs(2189));
    outputs(3643) <= (layer0_outputs(2912)) and not (layer0_outputs(2147));
    outputs(3644) <= not(layer0_outputs(5783));
    outputs(3645) <= (layer0_outputs(4199)) and not (layer0_outputs(5887));
    outputs(3646) <= layer0_outputs(3193);
    outputs(3647) <= layer0_outputs(972);
    outputs(3648) <= layer0_outputs(1297);
    outputs(3649) <= not(layer0_outputs(7001));
    outputs(3650) <= layer0_outputs(2076);
    outputs(3651) <= layer0_outputs(5372);
    outputs(3652) <= (layer0_outputs(6430)) and not (layer0_outputs(2672));
    outputs(3653) <= (layer0_outputs(3347)) xor (layer0_outputs(4165));
    outputs(3654) <= layer0_outputs(7257);
    outputs(3655) <= layer0_outputs(2616);
    outputs(3656) <= not(layer0_outputs(5503));
    outputs(3657) <= layer0_outputs(5054);
    outputs(3658) <= not(layer0_outputs(7067));
    outputs(3659) <= not(layer0_outputs(753));
    outputs(3660) <= not(layer0_outputs(4176));
    outputs(3661) <= not((layer0_outputs(7619)) and (layer0_outputs(468)));
    outputs(3662) <= layer0_outputs(2634);
    outputs(3663) <= layer0_outputs(398);
    outputs(3664) <= not(layer0_outputs(183));
    outputs(3665) <= not(layer0_outputs(6642));
    outputs(3666) <= not((layer0_outputs(1365)) or (layer0_outputs(2289)));
    outputs(3667) <= layer0_outputs(3166);
    outputs(3668) <= not(layer0_outputs(6300));
    outputs(3669) <= not(layer0_outputs(5943)) or (layer0_outputs(4777));
    outputs(3670) <= not((layer0_outputs(5985)) xor (layer0_outputs(2566)));
    outputs(3671) <= not(layer0_outputs(5178));
    outputs(3672) <= not(layer0_outputs(3));
    outputs(3673) <= layer0_outputs(234);
    outputs(3674) <= (layer0_outputs(434)) and (layer0_outputs(6456));
    outputs(3675) <= layer0_outputs(4515);
    outputs(3676) <= layer0_outputs(7533);
    outputs(3677) <= not(layer0_outputs(1710));
    outputs(3678) <= layer0_outputs(4479);
    outputs(3679) <= layer0_outputs(489);
    outputs(3680) <= not(layer0_outputs(4025));
    outputs(3681) <= not(layer0_outputs(1020));
    outputs(3682) <= (layer0_outputs(5502)) and (layer0_outputs(3501));
    outputs(3683) <= layer0_outputs(6053);
    outputs(3684) <= not(layer0_outputs(1097));
    outputs(3685) <= layer0_outputs(6290);
    outputs(3686) <= (layer0_outputs(5882)) xor (layer0_outputs(1665));
    outputs(3687) <= not(layer0_outputs(3600));
    outputs(3688) <= not(layer0_outputs(3120));
    outputs(3689) <= layer0_outputs(2502);
    outputs(3690) <= layer0_outputs(1970);
    outputs(3691) <= layer0_outputs(6030);
    outputs(3692) <= layer0_outputs(3144);
    outputs(3693) <= layer0_outputs(6424);
    outputs(3694) <= not(layer0_outputs(2240)) or (layer0_outputs(416));
    outputs(3695) <= (layer0_outputs(4130)) and not (layer0_outputs(2748));
    outputs(3696) <= (layer0_outputs(210)) and not (layer0_outputs(6078));
    outputs(3697) <= (layer0_outputs(387)) and not (layer0_outputs(6798));
    outputs(3698) <= not(layer0_outputs(3314)) or (layer0_outputs(6441));
    outputs(3699) <= not(layer0_outputs(6466));
    outputs(3700) <= layer0_outputs(773);
    outputs(3701) <= (layer0_outputs(1647)) xor (layer0_outputs(355));
    outputs(3702) <= not((layer0_outputs(4254)) xor (layer0_outputs(5784)));
    outputs(3703) <= not((layer0_outputs(6112)) or (layer0_outputs(169)));
    outputs(3704) <= layer0_outputs(4492);
    outputs(3705) <= (layer0_outputs(2714)) xor (layer0_outputs(2137));
    outputs(3706) <= (layer0_outputs(7260)) and not (layer0_outputs(1582));
    outputs(3707) <= not((layer0_outputs(574)) and (layer0_outputs(1686)));
    outputs(3708) <= (layer0_outputs(5674)) and not (layer0_outputs(2103));
    outputs(3709) <= not((layer0_outputs(5765)) xor (layer0_outputs(4690)));
    outputs(3710) <= layer0_outputs(3422);
    outputs(3711) <= layer0_outputs(4444);
    outputs(3712) <= layer0_outputs(3330);
    outputs(3713) <= not(layer0_outputs(2202));
    outputs(3714) <= layer0_outputs(5351);
    outputs(3715) <= layer0_outputs(6279);
    outputs(3716) <= layer0_outputs(2114);
    outputs(3717) <= (layer0_outputs(4957)) and (layer0_outputs(140));
    outputs(3718) <= not(layer0_outputs(1430));
    outputs(3719) <= not((layer0_outputs(6499)) xor (layer0_outputs(6263)));
    outputs(3720) <= not(layer0_outputs(5257)) or (layer0_outputs(2096));
    outputs(3721) <= not(layer0_outputs(857));
    outputs(3722) <= layer0_outputs(7274);
    outputs(3723) <= not(layer0_outputs(2386));
    outputs(3724) <= layer0_outputs(5697);
    outputs(3725) <= (layer0_outputs(2598)) and not (layer0_outputs(4078));
    outputs(3726) <= not(layer0_outputs(2205));
    outputs(3727) <= layer0_outputs(537);
    outputs(3728) <= not(layer0_outputs(6011));
    outputs(3729) <= not(layer0_outputs(6540)) or (layer0_outputs(3580));
    outputs(3730) <= not(layer0_outputs(5559));
    outputs(3731) <= not((layer0_outputs(1045)) or (layer0_outputs(2020)));
    outputs(3732) <= layer0_outputs(4233);
    outputs(3733) <= not(layer0_outputs(2752));
    outputs(3734) <= not(layer0_outputs(6444));
    outputs(3735) <= (layer0_outputs(4430)) and (layer0_outputs(4704));
    outputs(3736) <= not(layer0_outputs(5495));
    outputs(3737) <= not(layer0_outputs(2790));
    outputs(3738) <= not(layer0_outputs(3152)) or (layer0_outputs(4081));
    outputs(3739) <= not(layer0_outputs(491));
    outputs(3740) <= layer0_outputs(2849);
    outputs(3741) <= not(layer0_outputs(44)) or (layer0_outputs(3567));
    outputs(3742) <= not(layer0_outputs(3792));
    outputs(3743) <= (layer0_outputs(3919)) and not (layer0_outputs(287));
    outputs(3744) <= layer0_outputs(4298);
    outputs(3745) <= not(layer0_outputs(643));
    outputs(3746) <= not(layer0_outputs(3867));
    outputs(3747) <= (layer0_outputs(5974)) xor (layer0_outputs(2796));
    outputs(3748) <= layer0_outputs(6660);
    outputs(3749) <= not(layer0_outputs(1919));
    outputs(3750) <= layer0_outputs(4771);
    outputs(3751) <= (layer0_outputs(556)) and (layer0_outputs(6123));
    outputs(3752) <= layer0_outputs(6361);
    outputs(3753) <= layer0_outputs(3513);
    outputs(3754) <= layer0_outputs(6438);
    outputs(3755) <= not(layer0_outputs(3715));
    outputs(3756) <= layer0_outputs(7607);
    outputs(3757) <= layer0_outputs(2101);
    outputs(3758) <= not(layer0_outputs(3853)) or (layer0_outputs(3082));
    outputs(3759) <= layer0_outputs(6800);
    outputs(3760) <= layer0_outputs(1862);
    outputs(3761) <= not(layer0_outputs(3752));
    outputs(3762) <= not((layer0_outputs(3350)) or (layer0_outputs(5861)));
    outputs(3763) <= (layer0_outputs(2140)) xor (layer0_outputs(6314));
    outputs(3764) <= (layer0_outputs(1090)) and (layer0_outputs(3154));
    outputs(3765) <= layer0_outputs(7292);
    outputs(3766) <= layer0_outputs(4132);
    outputs(3767) <= (layer0_outputs(6961)) and not (layer0_outputs(4853));
    outputs(3768) <= layer0_outputs(902);
    outputs(3769) <= not(layer0_outputs(2927));
    outputs(3770) <= (layer0_outputs(7002)) and not (layer0_outputs(438));
    outputs(3771) <= layer0_outputs(6826);
    outputs(3772) <= layer0_outputs(3762);
    outputs(3773) <= layer0_outputs(4131);
    outputs(3774) <= layer0_outputs(62);
    outputs(3775) <= (layer0_outputs(7632)) xor (layer0_outputs(7582));
    outputs(3776) <= (layer0_outputs(2559)) and (layer0_outputs(2482));
    outputs(3777) <= not((layer0_outputs(782)) or (layer0_outputs(84)));
    outputs(3778) <= layer0_outputs(4411);
    outputs(3779) <= not(layer0_outputs(135));
    outputs(3780) <= layer0_outputs(5254);
    outputs(3781) <= not(layer0_outputs(584));
    outputs(3782) <= not(layer0_outputs(727));
    outputs(3783) <= not((layer0_outputs(5335)) or (layer0_outputs(6245)));
    outputs(3784) <= not(layer0_outputs(7271));
    outputs(3785) <= layer0_outputs(6608);
    outputs(3786) <= not(layer0_outputs(4269));
    outputs(3787) <= not(layer0_outputs(6488));
    outputs(3788) <= layer0_outputs(2738);
    outputs(3789) <= not(layer0_outputs(6589));
    outputs(3790) <= not(layer0_outputs(7360));
    outputs(3791) <= not(layer0_outputs(2205));
    outputs(3792) <= not((layer0_outputs(7129)) and (layer0_outputs(5535)));
    outputs(3793) <= (layer0_outputs(348)) xor (layer0_outputs(4877));
    outputs(3794) <= layer0_outputs(4418);
    outputs(3795) <= (layer0_outputs(5639)) and (layer0_outputs(4547));
    outputs(3796) <= (layer0_outputs(1624)) xor (layer0_outputs(6204));
    outputs(3797) <= (layer0_outputs(6715)) xor (layer0_outputs(2164));
    outputs(3798) <= not((layer0_outputs(7633)) xor (layer0_outputs(7604)));
    outputs(3799) <= (layer0_outputs(1683)) xor (layer0_outputs(1817));
    outputs(3800) <= not((layer0_outputs(6585)) or (layer0_outputs(3685)));
    outputs(3801) <= not((layer0_outputs(2795)) or (layer0_outputs(6427)));
    outputs(3802) <= layer0_outputs(63);
    outputs(3803) <= not(layer0_outputs(4110));
    outputs(3804) <= not(layer0_outputs(5957));
    outputs(3805) <= layer0_outputs(138);
    outputs(3806) <= (layer0_outputs(1295)) xor (layer0_outputs(4689));
    outputs(3807) <= (layer0_outputs(3384)) and not (layer0_outputs(910));
    outputs(3808) <= not(layer0_outputs(4002));
    outputs(3809) <= (layer0_outputs(1770)) and not (layer0_outputs(3118));
    outputs(3810) <= not(layer0_outputs(5846));
    outputs(3811) <= not((layer0_outputs(6787)) xor (layer0_outputs(4732)));
    outputs(3812) <= (layer0_outputs(139)) and not (layer0_outputs(2276));
    outputs(3813) <= not(layer0_outputs(1472));
    outputs(3814) <= not(layer0_outputs(1339)) or (layer0_outputs(6926));
    outputs(3815) <= layer0_outputs(558);
    outputs(3816) <= not((layer0_outputs(3413)) or (layer0_outputs(5106)));
    outputs(3817) <= layer0_outputs(1296);
    outputs(3818) <= (layer0_outputs(6517)) and (layer0_outputs(1295));
    outputs(3819) <= not(layer0_outputs(5182));
    outputs(3820) <= layer0_outputs(7573);
    outputs(3821) <= not(layer0_outputs(3271));
    outputs(3822) <= layer0_outputs(5618);
    outputs(3823) <= layer0_outputs(131);
    outputs(3824) <= not(layer0_outputs(1601));
    outputs(3825) <= not(layer0_outputs(2176));
    outputs(3826) <= not((layer0_outputs(41)) or (layer0_outputs(3680)));
    outputs(3827) <= not((layer0_outputs(565)) or (layer0_outputs(3900)));
    outputs(3828) <= (layer0_outputs(1073)) and not (layer0_outputs(2145));
    outputs(3829) <= (layer0_outputs(5569)) and not (layer0_outputs(7249));
    outputs(3830) <= not((layer0_outputs(1644)) or (layer0_outputs(3912)));
    outputs(3831) <= not(layer0_outputs(5880));
    outputs(3832) <= not(layer0_outputs(1708));
    outputs(3833) <= layer0_outputs(586);
    outputs(3834) <= not(layer0_outputs(6472));
    outputs(3835) <= (layer0_outputs(3359)) and not (layer0_outputs(7649));
    outputs(3836) <= layer0_outputs(5146);
    outputs(3837) <= (layer0_outputs(7180)) xor (layer0_outputs(1626));
    outputs(3838) <= layer0_outputs(4044);
    outputs(3839) <= not((layer0_outputs(1244)) xor (layer0_outputs(4858)));
    outputs(3840) <= not(layer0_outputs(291));
    outputs(3841) <= not((layer0_outputs(948)) xor (layer0_outputs(3243)));
    outputs(3842) <= layer0_outputs(1913);
    outputs(3843) <= not((layer0_outputs(1152)) xor (layer0_outputs(621)));
    outputs(3844) <= layer0_outputs(4731);
    outputs(3845) <= not(layer0_outputs(2162)) or (layer0_outputs(1350));
    outputs(3846) <= (layer0_outputs(1746)) and not (layer0_outputs(2045));
    outputs(3847) <= not((layer0_outputs(4871)) xor (layer0_outputs(5012)));
    outputs(3848) <= layer0_outputs(2260);
    outputs(3849) <= not((layer0_outputs(5498)) xor (layer0_outputs(1079)));
    outputs(3850) <= layer0_outputs(5772);
    outputs(3851) <= not(layer0_outputs(7219)) or (layer0_outputs(3470));
    outputs(3852) <= layer0_outputs(3713);
    outputs(3853) <= layer0_outputs(6059);
    outputs(3854) <= not((layer0_outputs(4132)) xor (layer0_outputs(6763)));
    outputs(3855) <= (layer0_outputs(3510)) and not (layer0_outputs(2816));
    outputs(3856) <= not(layer0_outputs(4444));
    outputs(3857) <= layer0_outputs(6915);
    outputs(3858) <= layer0_outputs(1214);
    outputs(3859) <= layer0_outputs(6588);
    outputs(3860) <= not((layer0_outputs(3096)) xor (layer0_outputs(1168)));
    outputs(3861) <= (layer0_outputs(6598)) xor (layer0_outputs(7377));
    outputs(3862) <= layer0_outputs(5090);
    outputs(3863) <= not(layer0_outputs(3339));
    outputs(3864) <= not((layer0_outputs(2471)) xor (layer0_outputs(5036)));
    outputs(3865) <= (layer0_outputs(2930)) and (layer0_outputs(6917));
    outputs(3866) <= (layer0_outputs(1257)) and (layer0_outputs(7390));
    outputs(3867) <= not(layer0_outputs(3704));
    outputs(3868) <= not(layer0_outputs(7186));
    outputs(3869) <= layer0_outputs(2760);
    outputs(3870) <= not(layer0_outputs(594));
    outputs(3871) <= layer0_outputs(5420);
    outputs(3872) <= (layer0_outputs(1045)) and not (layer0_outputs(173));
    outputs(3873) <= layer0_outputs(7072);
    outputs(3874) <= not(layer0_outputs(2273));
    outputs(3875) <= layer0_outputs(915);
    outputs(3876) <= layer0_outputs(4743);
    outputs(3877) <= not(layer0_outputs(3813));
    outputs(3878) <= (layer0_outputs(3664)) and not (layer0_outputs(5962));
    outputs(3879) <= not((layer0_outputs(339)) or (layer0_outputs(3324)));
    outputs(3880) <= (layer0_outputs(5508)) xor (layer0_outputs(133));
    outputs(3881) <= not(layer0_outputs(3716));
    outputs(3882) <= not((layer0_outputs(1596)) or (layer0_outputs(4028)));
    outputs(3883) <= layer0_outputs(457);
    outputs(3884) <= layer0_outputs(1829);
    outputs(3885) <= not(layer0_outputs(4392));
    outputs(3886) <= (layer0_outputs(700)) and not (layer0_outputs(3869));
    outputs(3887) <= not((layer0_outputs(7465)) or (layer0_outputs(5103)));
    outputs(3888) <= not((layer0_outputs(254)) xor (layer0_outputs(2064)));
    outputs(3889) <= not(layer0_outputs(3141));
    outputs(3890) <= not((layer0_outputs(6316)) xor (layer0_outputs(1222)));
    outputs(3891) <= (layer0_outputs(951)) and not (layer0_outputs(3718));
    outputs(3892) <= not((layer0_outputs(2509)) xor (layer0_outputs(2578)));
    outputs(3893) <= layer0_outputs(2817);
    outputs(3894) <= layer0_outputs(5710);
    outputs(3895) <= not((layer0_outputs(1791)) xor (layer0_outputs(5122)));
    outputs(3896) <= not(layer0_outputs(7272));
    outputs(3897) <= (layer0_outputs(6303)) xor (layer0_outputs(7595));
    outputs(3898) <= not(layer0_outputs(5110));
    outputs(3899) <= layer0_outputs(15);
    outputs(3900) <= (layer0_outputs(2870)) and not (layer0_outputs(6007));
    outputs(3901) <= not(layer0_outputs(2348));
    outputs(3902) <= (layer0_outputs(898)) and not (layer0_outputs(1144));
    outputs(3903) <= not((layer0_outputs(5420)) xor (layer0_outputs(2464)));
    outputs(3904) <= not((layer0_outputs(5564)) xor (layer0_outputs(4027)));
    outputs(3905) <= not((layer0_outputs(3098)) xor (layer0_outputs(282)));
    outputs(3906) <= layer0_outputs(5723);
    outputs(3907) <= not((layer0_outputs(2799)) xor (layer0_outputs(4011)));
    outputs(3908) <= not(layer0_outputs(3031));
    outputs(3909) <= not((layer0_outputs(4631)) and (layer0_outputs(7283)));
    outputs(3910) <= layer0_outputs(7161);
    outputs(3911) <= not((layer0_outputs(6599)) xor (layer0_outputs(2604)));
    outputs(3912) <= not((layer0_outputs(4384)) xor (layer0_outputs(1788)));
    outputs(3913) <= (layer0_outputs(6443)) or (layer0_outputs(5760));
    outputs(3914) <= (layer0_outputs(2611)) xor (layer0_outputs(6334));
    outputs(3915) <= not(layer0_outputs(3370));
    outputs(3916) <= not((layer0_outputs(7427)) xor (layer0_outputs(2531)));
    outputs(3917) <= (layer0_outputs(5751)) and (layer0_outputs(1248));
    outputs(3918) <= layer0_outputs(2554);
    outputs(3919) <= not(layer0_outputs(2901));
    outputs(3920) <= layer0_outputs(4179);
    outputs(3921) <= not((layer0_outputs(5476)) or (layer0_outputs(6706)));
    outputs(3922) <= not(layer0_outputs(3308)) or (layer0_outputs(363));
    outputs(3923) <= not(layer0_outputs(6652));
    outputs(3924) <= not((layer0_outputs(3840)) xor (layer0_outputs(4153)));
    outputs(3925) <= not(layer0_outputs(6352));
    outputs(3926) <= layer0_outputs(7594);
    outputs(3927) <= not(layer0_outputs(1816)) or (layer0_outputs(7401));
    outputs(3928) <= not((layer0_outputs(2276)) xor (layer0_outputs(4837)));
    outputs(3929) <= not(layer0_outputs(7091));
    outputs(3930) <= not((layer0_outputs(562)) xor (layer0_outputs(6870)));
    outputs(3931) <= layer0_outputs(1492);
    outputs(3932) <= layer0_outputs(3627);
    outputs(3933) <= layer0_outputs(276);
    outputs(3934) <= not((layer0_outputs(1799)) xor (layer0_outputs(4386)));
    outputs(3935) <= not(layer0_outputs(2750));
    outputs(3936) <= not((layer0_outputs(3528)) xor (layer0_outputs(1349)));
    outputs(3937) <= not((layer0_outputs(4649)) xor (layer0_outputs(1043)));
    outputs(3938) <= layer0_outputs(5240);
    outputs(3939) <= not(layer0_outputs(2408));
    outputs(3940) <= not(layer0_outputs(1517));
    outputs(3941) <= not(layer0_outputs(5531));
    outputs(3942) <= not(layer0_outputs(3293));
    outputs(3943) <= layer0_outputs(5950);
    outputs(3944) <= not((layer0_outputs(7298)) xor (layer0_outputs(5598)));
    outputs(3945) <= (layer0_outputs(4473)) xor (layer0_outputs(5375));
    outputs(3946) <= not(layer0_outputs(2618));
    outputs(3947) <= layer0_outputs(2312);
    outputs(3948) <= not(layer0_outputs(2347));
    outputs(3949) <= (layer0_outputs(2669)) and (layer0_outputs(2582));
    outputs(3950) <= layer0_outputs(3884);
    outputs(3951) <= (layer0_outputs(774)) and (layer0_outputs(7605));
    outputs(3952) <= not(layer0_outputs(7149)) or (layer0_outputs(115));
    outputs(3953) <= (layer0_outputs(540)) and not (layer0_outputs(2365));
    outputs(3954) <= (layer0_outputs(4590)) and not (layer0_outputs(7296));
    outputs(3955) <= (layer0_outputs(4200)) xor (layer0_outputs(4249));
    outputs(3956) <= layer0_outputs(7201);
    outputs(3957) <= not(layer0_outputs(1604));
    outputs(3958) <= (layer0_outputs(4817)) xor (layer0_outputs(490));
    outputs(3959) <= layer0_outputs(3903);
    outputs(3960) <= (layer0_outputs(1621)) or (layer0_outputs(5211));
    outputs(3961) <= (layer0_outputs(3801)) and not (layer0_outputs(3340));
    outputs(3962) <= (layer0_outputs(7071)) xor (layer0_outputs(1334));
    outputs(3963) <= (layer0_outputs(3652)) and not (layer0_outputs(1403));
    outputs(3964) <= (layer0_outputs(2122)) xor (layer0_outputs(6411));
    outputs(3965) <= not(layer0_outputs(1182));
    outputs(3966) <= layer0_outputs(349);
    outputs(3967) <= not((layer0_outputs(5230)) xor (layer0_outputs(5457)));
    outputs(3968) <= not(layer0_outputs(4592)) or (layer0_outputs(2443));
    outputs(3969) <= (layer0_outputs(5343)) and not (layer0_outputs(1760));
    outputs(3970) <= layer0_outputs(6768);
    outputs(3971) <= not(layer0_outputs(6493)) or (layer0_outputs(6054));
    outputs(3972) <= layer0_outputs(1594);
    outputs(3973) <= not(layer0_outputs(2918));
    outputs(3974) <= not(layer0_outputs(5236)) or (layer0_outputs(1074));
    outputs(3975) <= (layer0_outputs(2542)) or (layer0_outputs(2324));
    outputs(3976) <= not(layer0_outputs(1880));
    outputs(3977) <= layer0_outputs(1319);
    outputs(3978) <= layer0_outputs(5768);
    outputs(3979) <= (layer0_outputs(7604)) and not (layer0_outputs(4326));
    outputs(3980) <= not((layer0_outputs(4820)) or (layer0_outputs(3372)));
    outputs(3981) <= layer0_outputs(2465);
    outputs(3982) <= (layer0_outputs(2311)) xor (layer0_outputs(6489));
    outputs(3983) <= layer0_outputs(4447);
    outputs(3984) <= (layer0_outputs(4480)) xor (layer0_outputs(766));
    outputs(3985) <= not(layer0_outputs(3194)) or (layer0_outputs(3859));
    outputs(3986) <= not((layer0_outputs(4117)) xor (layer0_outputs(255)));
    outputs(3987) <= layer0_outputs(2014);
    outputs(3988) <= not(layer0_outputs(5363));
    outputs(3989) <= not((layer0_outputs(1453)) xor (layer0_outputs(2017)));
    outputs(3990) <= (layer0_outputs(5987)) and not (layer0_outputs(613));
    outputs(3991) <= layer0_outputs(2742);
    outputs(3992) <= layer0_outputs(6247);
    outputs(3993) <= (layer0_outputs(4435)) xor (layer0_outputs(1898));
    outputs(3994) <= (layer0_outputs(6095)) xor (layer0_outputs(1206));
    outputs(3995) <= not(layer0_outputs(3896));
    outputs(3996) <= layer0_outputs(936);
    outputs(3997) <= layer0_outputs(2623);
    outputs(3998) <= layer0_outputs(6424);
    outputs(3999) <= (layer0_outputs(2526)) or (layer0_outputs(3136));
    outputs(4000) <= layer0_outputs(5988);
    outputs(4001) <= (layer0_outputs(5361)) xor (layer0_outputs(7305));
    outputs(4002) <= (layer0_outputs(6267)) xor (layer0_outputs(708));
    outputs(4003) <= (layer0_outputs(6182)) and not (layer0_outputs(7420));
    outputs(4004) <= not(layer0_outputs(851));
    outputs(4005) <= not((layer0_outputs(1500)) xor (layer0_outputs(28)));
    outputs(4006) <= not(layer0_outputs(1625)) or (layer0_outputs(2385));
    outputs(4007) <= layer0_outputs(5779);
    outputs(4008) <= layer0_outputs(245);
    outputs(4009) <= not(layer0_outputs(2333)) or (layer0_outputs(1381));
    outputs(4010) <= (layer0_outputs(2950)) or (layer0_outputs(6808));
    outputs(4011) <= layer0_outputs(6967);
    outputs(4012) <= (layer0_outputs(1096)) and not (layer0_outputs(3925));
    outputs(4013) <= not(layer0_outputs(6894));
    outputs(4014) <= layer0_outputs(6043);
    outputs(4015) <= layer0_outputs(1972);
    outputs(4016) <= layer0_outputs(6993);
    outputs(4017) <= (layer0_outputs(661)) and not (layer0_outputs(2627));
    outputs(4018) <= layer0_outputs(6596);
    outputs(4019) <= not(layer0_outputs(4523));
    outputs(4020) <= (layer0_outputs(4291)) xor (layer0_outputs(3014));
    outputs(4021) <= not((layer0_outputs(789)) xor (layer0_outputs(3325)));
    outputs(4022) <= (layer0_outputs(4371)) xor (layer0_outputs(2458));
    outputs(4023) <= not((layer0_outputs(5615)) xor (layer0_outputs(6038)));
    outputs(4024) <= layer0_outputs(2809);
    outputs(4025) <= not((layer0_outputs(1369)) or (layer0_outputs(7593)));
    outputs(4026) <= not((layer0_outputs(2589)) xor (layer0_outputs(214)));
    outputs(4027) <= not((layer0_outputs(102)) or (layer0_outputs(7580)));
    outputs(4028) <= not(layer0_outputs(1538));
    outputs(4029) <= not(layer0_outputs(4830));
    outputs(4030) <= not(layer0_outputs(3770));
    outputs(4031) <= layer0_outputs(2841);
    outputs(4032) <= not(layer0_outputs(4939));
    outputs(4033) <= not((layer0_outputs(2770)) xor (layer0_outputs(6165)));
    outputs(4034) <= (layer0_outputs(629)) xor (layer0_outputs(7096));
    outputs(4035) <= not((layer0_outputs(4933)) and (layer0_outputs(4741)));
    outputs(4036) <= (layer0_outputs(7453)) xor (layer0_outputs(1715));
    outputs(4037) <= (layer0_outputs(5712)) or (layer0_outputs(5678));
    outputs(4038) <= not(layer0_outputs(1566));
    outputs(4039) <= not((layer0_outputs(4754)) xor (layer0_outputs(1910)));
    outputs(4040) <= layer0_outputs(3434);
    outputs(4041) <= (layer0_outputs(5920)) xor (layer0_outputs(3614));
    outputs(4042) <= not((layer0_outputs(5876)) xor (layer0_outputs(5368)));
    outputs(4043) <= not(layer0_outputs(1956));
    outputs(4044) <= not(layer0_outputs(4222));
    outputs(4045) <= not((layer0_outputs(4847)) and (layer0_outputs(5722)));
    outputs(4046) <= not(layer0_outputs(5095));
    outputs(4047) <= not(layer0_outputs(619)) or (layer0_outputs(2548));
    outputs(4048) <= not(layer0_outputs(811)) or (layer0_outputs(6462));
    outputs(4049) <= not(layer0_outputs(7066));
    outputs(4050) <= layer0_outputs(1535);
    outputs(4051) <= not((layer0_outputs(2824)) xor (layer0_outputs(1892)));
    outputs(4052) <= (layer0_outputs(2682)) and not (layer0_outputs(1600));
    outputs(4053) <= not(layer0_outputs(5206));
    outputs(4054) <= not(layer0_outputs(3161));
    outputs(4055) <= layer0_outputs(7505);
    outputs(4056) <= (layer0_outputs(3851)) xor (layer0_outputs(1802));
    outputs(4057) <= not(layer0_outputs(1094));
    outputs(4058) <= not(layer0_outputs(950));
    outputs(4059) <= not(layer0_outputs(30));
    outputs(4060) <= layer0_outputs(4573);
    outputs(4061) <= not(layer0_outputs(5968));
    outputs(4062) <= layer0_outputs(1920);
    outputs(4063) <= layer0_outputs(1825);
    outputs(4064) <= not((layer0_outputs(3948)) xor (layer0_outputs(6985)));
    outputs(4065) <= not((layer0_outputs(1237)) or (layer0_outputs(7316)));
    outputs(4066) <= (layer0_outputs(3386)) or (layer0_outputs(3477));
    outputs(4067) <= (layer0_outputs(5523)) and not (layer0_outputs(5875));
    outputs(4068) <= (layer0_outputs(1130)) and (layer0_outputs(4038));
    outputs(4069) <= not(layer0_outputs(1072));
    outputs(4070) <= layer0_outputs(1713);
    outputs(4071) <= layer0_outputs(7246);
    outputs(4072) <= (layer0_outputs(2026)) xor (layer0_outputs(6331));
    outputs(4073) <= layer0_outputs(4004);
    outputs(4074) <= not(layer0_outputs(2265));
    outputs(4075) <= layer0_outputs(4537);
    outputs(4076) <= layer0_outputs(4638);
    outputs(4077) <= not(layer0_outputs(4222));
    outputs(4078) <= not((layer0_outputs(3368)) xor (layer0_outputs(6105)));
    outputs(4079) <= not(layer0_outputs(5136)) or (layer0_outputs(6783));
    outputs(4080) <= not((layer0_outputs(6032)) xor (layer0_outputs(21)));
    outputs(4081) <= not(layer0_outputs(2975));
    outputs(4082) <= not(layer0_outputs(3227));
    outputs(4083) <= not(layer0_outputs(1366));
    outputs(4084) <= not(layer0_outputs(1469));
    outputs(4085) <= not(layer0_outputs(439));
    outputs(4086) <= (layer0_outputs(6075)) and (layer0_outputs(4046));
    outputs(4087) <= not(layer0_outputs(152)) or (layer0_outputs(3296));
    outputs(4088) <= (layer0_outputs(1853)) and not (layer0_outputs(2184));
    outputs(4089) <= layer0_outputs(4891);
    outputs(4090) <= not(layer0_outputs(3654)) or (layer0_outputs(6581));
    outputs(4091) <= layer0_outputs(1931);
    outputs(4092) <= (layer0_outputs(50)) xor (layer0_outputs(4526));
    outputs(4093) <= (layer0_outputs(2710)) or (layer0_outputs(4887));
    outputs(4094) <= layer0_outputs(5659);
    outputs(4095) <= (layer0_outputs(4502)) and not (layer0_outputs(7517));
    outputs(4096) <= not((layer0_outputs(3022)) xor (layer0_outputs(2036)));
    outputs(4097) <= (layer0_outputs(577)) and not (layer0_outputs(3756));
    outputs(4098) <= not(layer0_outputs(3537));
    outputs(4099) <= not(layer0_outputs(328));
    outputs(4100) <= not(layer0_outputs(729));
    outputs(4101) <= (layer0_outputs(7340)) and (layer0_outputs(3454));
    outputs(4102) <= (layer0_outputs(7624)) xor (layer0_outputs(4354));
    outputs(4103) <= layer0_outputs(7312);
    outputs(4104) <= not((layer0_outputs(1532)) xor (layer0_outputs(5748)));
    outputs(4105) <= (layer0_outputs(3811)) xor (layer0_outputs(1974));
    outputs(4106) <= not((layer0_outputs(3987)) and (layer0_outputs(6745)));
    outputs(4107) <= (layer0_outputs(4887)) and not (layer0_outputs(336));
    outputs(4108) <= not((layer0_outputs(3420)) xor (layer0_outputs(4056)));
    outputs(4109) <= layer0_outputs(4442);
    outputs(4110) <= not((layer0_outputs(3098)) xor (layer0_outputs(2561)));
    outputs(4111) <= not((layer0_outputs(6373)) or (layer0_outputs(7203)));
    outputs(4112) <= not(layer0_outputs(5048));
    outputs(4113) <= not((layer0_outputs(2785)) xor (layer0_outputs(5102)));
    outputs(4114) <= layer0_outputs(4839);
    outputs(4115) <= not((layer0_outputs(5405)) xor (layer0_outputs(494)));
    outputs(4116) <= not((layer0_outputs(5400)) xor (layer0_outputs(5706)));
    outputs(4117) <= layer0_outputs(4091);
    outputs(4118) <= not(layer0_outputs(2849)) or (layer0_outputs(7026));
    outputs(4119) <= layer0_outputs(6895);
    outputs(4120) <= (layer0_outputs(3158)) xor (layer0_outputs(5527));
    outputs(4121) <= '0';
    outputs(4122) <= (layer0_outputs(2119)) xor (layer0_outputs(5192));
    outputs(4123) <= not((layer0_outputs(625)) xor (layer0_outputs(2899)));
    outputs(4124) <= not(layer0_outputs(467));
    outputs(4125) <= layer0_outputs(4517);
    outputs(4126) <= (layer0_outputs(877)) and (layer0_outputs(7407));
    outputs(4127) <= not((layer0_outputs(6986)) xor (layer0_outputs(3788)));
    outputs(4128) <= layer0_outputs(3070);
    outputs(4129) <= not(layer0_outputs(6248));
    outputs(4130) <= not(layer0_outputs(4961));
    outputs(4131) <= not((layer0_outputs(1219)) xor (layer0_outputs(5642)));
    outputs(4132) <= not(layer0_outputs(1517));
    outputs(4133) <= not((layer0_outputs(4690)) or (layer0_outputs(2199)));
    outputs(4134) <= (layer0_outputs(5336)) xor (layer0_outputs(271));
    outputs(4135) <= layer0_outputs(4554);
    outputs(4136) <= not(layer0_outputs(3620));
    outputs(4137) <= not(layer0_outputs(5152));
    outputs(4138) <= layer0_outputs(6137);
    outputs(4139) <= not(layer0_outputs(6065));
    outputs(4140) <= not((layer0_outputs(5590)) xor (layer0_outputs(6506)));
    outputs(4141) <= not((layer0_outputs(5666)) xor (layer0_outputs(5255)));
    outputs(4142) <= not((layer0_outputs(2794)) or (layer0_outputs(6866)));
    outputs(4143) <= layer0_outputs(1490);
    outputs(4144) <= not(layer0_outputs(3600));
    outputs(4145) <= not(layer0_outputs(3357));
    outputs(4146) <= not((layer0_outputs(191)) xor (layer0_outputs(1205)));
    outputs(4147) <= not((layer0_outputs(431)) or (layer0_outputs(4541)));
    outputs(4148) <= not(layer0_outputs(2174));
    outputs(4149) <= not((layer0_outputs(3278)) xor (layer0_outputs(4356)));
    outputs(4150) <= layer0_outputs(2467);
    outputs(4151) <= (layer0_outputs(7373)) xor (layer0_outputs(7464));
    outputs(4152) <= not(layer0_outputs(6085));
    outputs(4153) <= not(layer0_outputs(3447));
    outputs(4154) <= not((layer0_outputs(6992)) xor (layer0_outputs(7140)));
    outputs(4155) <= not((layer0_outputs(1622)) xor (layer0_outputs(1429)));
    outputs(4156) <= layer0_outputs(6274);
    outputs(4157) <= not(layer0_outputs(864));
    outputs(4158) <= layer0_outputs(3879);
    outputs(4159) <= not(layer0_outputs(1654));
    outputs(4160) <= not(layer0_outputs(4459));
    outputs(4161) <= not(layer0_outputs(5804)) or (layer0_outputs(3604));
    outputs(4162) <= (layer0_outputs(2662)) xor (layer0_outputs(1003));
    outputs(4163) <= not((layer0_outputs(6318)) or (layer0_outputs(3312)));
    outputs(4164) <= not(layer0_outputs(3202));
    outputs(4165) <= layer0_outputs(2835);
    outputs(4166) <= (layer0_outputs(1975)) and (layer0_outputs(4406));
    outputs(4167) <= not((layer0_outputs(2980)) or (layer0_outputs(4970)));
    outputs(4168) <= layer0_outputs(4224);
    outputs(4169) <= layer0_outputs(5717);
    outputs(4170) <= (layer0_outputs(6903)) xor (layer0_outputs(2193));
    outputs(4171) <= not((layer0_outputs(4620)) xor (layer0_outputs(3491)));
    outputs(4172) <= not(layer0_outputs(3412));
    outputs(4173) <= (layer0_outputs(6362)) xor (layer0_outputs(1580));
    outputs(4174) <= (layer0_outputs(4659)) and (layer0_outputs(5951));
    outputs(4175) <= layer0_outputs(6355);
    outputs(4176) <= not(layer0_outputs(4511)) or (layer0_outputs(2624));
    outputs(4177) <= not(layer0_outputs(101)) or (layer0_outputs(702));
    outputs(4178) <= not(layer0_outputs(6875));
    outputs(4179) <= (layer0_outputs(2396)) xor (layer0_outputs(1208));
    outputs(4180) <= layer0_outputs(4713);
    outputs(4181) <= (layer0_outputs(2576)) and not (layer0_outputs(5064));
    outputs(4182) <= layer0_outputs(2272);
    outputs(4183) <= not((layer0_outputs(2076)) or (layer0_outputs(962)));
    outputs(4184) <= layer0_outputs(3694);
    outputs(4185) <= (layer0_outputs(7152)) and not (layer0_outputs(7415));
    outputs(4186) <= layer0_outputs(1463);
    outputs(4187) <= not(layer0_outputs(4742));
    outputs(4188) <= not(layer0_outputs(2492));
    outputs(4189) <= (layer0_outputs(2978)) and (layer0_outputs(4767));
    outputs(4190) <= not((layer0_outputs(1028)) xor (layer0_outputs(1261)));
    outputs(4191) <= layer0_outputs(1380);
    outputs(4192) <= not((layer0_outputs(2068)) xor (layer0_outputs(1384)));
    outputs(4193) <= layer0_outputs(1176);
    outputs(4194) <= layer0_outputs(4255);
    outputs(4195) <= not((layer0_outputs(572)) xor (layer0_outputs(3837)));
    outputs(4196) <= not((layer0_outputs(6671)) xor (layer0_outputs(1009)));
    outputs(4197) <= not(layer0_outputs(5775));
    outputs(4198) <= not(layer0_outputs(3611));
    outputs(4199) <= (layer0_outputs(1038)) xor (layer0_outputs(5597));
    outputs(4200) <= (layer0_outputs(5443)) and not (layer0_outputs(5720));
    outputs(4201) <= not(layer0_outputs(3167)) or (layer0_outputs(2708));
    outputs(4202) <= not(layer0_outputs(6064)) or (layer0_outputs(5799));
    outputs(4203) <= (layer0_outputs(6294)) and not (layer0_outputs(7373));
    outputs(4204) <= (layer0_outputs(5633)) xor (layer0_outputs(2251));
    outputs(4205) <= (layer0_outputs(5622)) and not (layer0_outputs(4518));
    outputs(4206) <= layer0_outputs(4748);
    outputs(4207) <= layer0_outputs(1281);
    outputs(4208) <= (layer0_outputs(3701)) xor (layer0_outputs(1154));
    outputs(4209) <= not((layer0_outputs(2125)) or (layer0_outputs(834)));
    outputs(4210) <= layer0_outputs(7338);
    outputs(4211) <= not(layer0_outputs(1940));
    outputs(4212) <= layer0_outputs(1800);
    outputs(4213) <= layer0_outputs(4186);
    outputs(4214) <= not(layer0_outputs(1015));
    outputs(4215) <= layer0_outputs(7329);
    outputs(4216) <= not(layer0_outputs(6950));
    outputs(4217) <= layer0_outputs(7221);
    outputs(4218) <= (layer0_outputs(4075)) and not (layer0_outputs(6177));
    outputs(4219) <= not(layer0_outputs(6049));
    outputs(4220) <= (layer0_outputs(3929)) and not (layer0_outputs(7589));
    outputs(4221) <= not(layer0_outputs(6351));
    outputs(4222) <= not(layer0_outputs(2606));
    outputs(4223) <= layer0_outputs(5721);
    outputs(4224) <= (layer0_outputs(4951)) and not (layer0_outputs(1136));
    outputs(4225) <= (layer0_outputs(3374)) and (layer0_outputs(3972));
    outputs(4226) <= not((layer0_outputs(2884)) xor (layer0_outputs(3225)));
    outputs(4227) <= layer0_outputs(5439);
    outputs(4228) <= (layer0_outputs(2863)) xor (layer0_outputs(1804));
    outputs(4229) <= (layer0_outputs(2144)) xor (layer0_outputs(6286));
    outputs(4230) <= (layer0_outputs(5255)) xor (layer0_outputs(620));
    outputs(4231) <= not((layer0_outputs(5553)) xor (layer0_outputs(3365)));
    outputs(4232) <= (layer0_outputs(7437)) and not (layer0_outputs(4898));
    outputs(4233) <= not((layer0_outputs(4165)) xor (layer0_outputs(1434)));
    outputs(4234) <= not(layer0_outputs(7074));
    outputs(4235) <= not(layer0_outputs(5838));
    outputs(4236) <= not(layer0_outputs(7417));
    outputs(4237) <= not(layer0_outputs(3961));
    outputs(4238) <= not(layer0_outputs(3915));
    outputs(4239) <= not(layer0_outputs(3620)) or (layer0_outputs(5868));
    outputs(4240) <= (layer0_outputs(1179)) xor (layer0_outputs(3710));
    outputs(4241) <= (layer0_outputs(5550)) xor (layer0_outputs(5528));
    outputs(4242) <= (layer0_outputs(867)) xor (layer0_outputs(5139));
    outputs(4243) <= (layer0_outputs(3019)) and not (layer0_outputs(1470));
    outputs(4244) <= (layer0_outputs(4144)) xor (layer0_outputs(3185));
    outputs(4245) <= not((layer0_outputs(7578)) or (layer0_outputs(5612)));
    outputs(4246) <= not(layer0_outputs(7200));
    outputs(4247) <= not((layer0_outputs(4695)) and (layer0_outputs(2762)));
    outputs(4248) <= layer0_outputs(506);
    outputs(4249) <= layer0_outputs(4731);
    outputs(4250) <= layer0_outputs(639);
    outputs(4251) <= (layer0_outputs(7667)) xor (layer0_outputs(2902));
    outputs(4252) <= not((layer0_outputs(2649)) xor (layer0_outputs(6975)));
    outputs(4253) <= (layer0_outputs(7085)) and (layer0_outputs(1877));
    outputs(4254) <= not((layer0_outputs(2804)) xor (layer0_outputs(3476)));
    outputs(4255) <= not(layer0_outputs(91));
    outputs(4256) <= not(layer0_outputs(4727));
    outputs(4257) <= (layer0_outputs(4187)) and (layer0_outputs(5761));
    outputs(4258) <= not(layer0_outputs(2491));
    outputs(4259) <= not((layer0_outputs(5274)) and (layer0_outputs(895)));
    outputs(4260) <= not((layer0_outputs(4613)) xor (layer0_outputs(5327)));
    outputs(4261) <= not(layer0_outputs(6308)) or (layer0_outputs(7208));
    outputs(4262) <= not(layer0_outputs(6863));
    outputs(4263) <= not((layer0_outputs(4699)) and (layer0_outputs(3101)));
    outputs(4264) <= (layer0_outputs(2437)) and not (layer0_outputs(2377));
    outputs(4265) <= not(layer0_outputs(5246));
    outputs(4266) <= not(layer0_outputs(5049));
    outputs(4267) <= layer0_outputs(4058);
    outputs(4268) <= not(layer0_outputs(1631));
    outputs(4269) <= layer0_outputs(4823);
    outputs(4270) <= layer0_outputs(6669);
    outputs(4271) <= (layer0_outputs(5808)) xor (layer0_outputs(6504));
    outputs(4272) <= not(layer0_outputs(6157));
    outputs(4273) <= layer0_outputs(2872);
    outputs(4274) <= (layer0_outputs(6408)) and not (layer0_outputs(2038));
    outputs(4275) <= not((layer0_outputs(6828)) xor (layer0_outputs(7259)));
    outputs(4276) <= layer0_outputs(280);
    outputs(4277) <= (layer0_outputs(4766)) or (layer0_outputs(2906));
    outputs(4278) <= layer0_outputs(1729);
    outputs(4279) <= not(layer0_outputs(6463)) or (layer0_outputs(4490));
    outputs(4280) <= layer0_outputs(5620);
    outputs(4281) <= not((layer0_outputs(6311)) xor (layer0_outputs(5179)));
    outputs(4282) <= not(layer0_outputs(3169));
    outputs(4283) <= layer0_outputs(7269);
    outputs(4284) <= layer0_outputs(6731);
    outputs(4285) <= (layer0_outputs(373)) and not (layer0_outputs(6746));
    outputs(4286) <= (layer0_outputs(403)) or (layer0_outputs(5547));
    outputs(4287) <= not(layer0_outputs(1501));
    outputs(4288) <= (layer0_outputs(2837)) xor (layer0_outputs(3928));
    outputs(4289) <= (layer0_outputs(6050)) xor (layer0_outputs(3554));
    outputs(4290) <= not(layer0_outputs(4013)) or (layer0_outputs(450));
    outputs(4291) <= not(layer0_outputs(1450));
    outputs(4292) <= layer0_outputs(3529);
    outputs(4293) <= not(layer0_outputs(1335));
    outputs(4294) <= not(layer0_outputs(166)) or (layer0_outputs(6284));
    outputs(4295) <= layer0_outputs(1741);
    outputs(4296) <= not(layer0_outputs(1718));
    outputs(4297) <= (layer0_outputs(6455)) xor (layer0_outputs(2562));
    outputs(4298) <= layer0_outputs(2887);
    outputs(4299) <= not(layer0_outputs(952));
    outputs(4300) <= (layer0_outputs(3818)) xor (layer0_outputs(78));
    outputs(4301) <= not(layer0_outputs(5572));
    outputs(4302) <= not(layer0_outputs(7017));
    outputs(4303) <= not((layer0_outputs(4785)) or (layer0_outputs(6409)));
    outputs(4304) <= layer0_outputs(6001);
    outputs(4305) <= (layer0_outputs(6425)) and (layer0_outputs(3414));
    outputs(4306) <= layer0_outputs(52);
    outputs(4307) <= (layer0_outputs(3578)) xor (layer0_outputs(2424));
    outputs(4308) <= not(layer0_outputs(5350));
    outputs(4309) <= not((layer0_outputs(1238)) and (layer0_outputs(3742)));
    outputs(4310) <= not(layer0_outputs(5822));
    outputs(4311) <= layer0_outputs(5931);
    outputs(4312) <= not(layer0_outputs(1028));
    outputs(4313) <= layer0_outputs(5548);
    outputs(4314) <= not(layer0_outputs(7105)) or (layer0_outputs(3822));
    outputs(4315) <= layer0_outputs(4554);
    outputs(4316) <= not(layer0_outputs(5126));
    outputs(4317) <= (layer0_outputs(4179)) and (layer0_outputs(4317));
    outputs(4318) <= not(layer0_outputs(3995));
    outputs(4319) <= layer0_outputs(4256);
    outputs(4320) <= (layer0_outputs(4214)) and not (layer0_outputs(6471));
    outputs(4321) <= layer0_outputs(4089);
    outputs(4322) <= (layer0_outputs(5589)) xor (layer0_outputs(1390));
    outputs(4323) <= not(layer0_outputs(7004));
    outputs(4324) <= layer0_outputs(4157);
    outputs(4325) <= not((layer0_outputs(4830)) or (layer0_outputs(5859)));
    outputs(4326) <= (layer0_outputs(3298)) xor (layer0_outputs(609));
    outputs(4327) <= not(layer0_outputs(6591)) or (layer0_outputs(5558));
    outputs(4328) <= not((layer0_outputs(1358)) or (layer0_outputs(5449)));
    outputs(4329) <= layer0_outputs(4944);
    outputs(4330) <= not(layer0_outputs(7277));
    outputs(4331) <= not((layer0_outputs(2944)) and (layer0_outputs(263)));
    outputs(4332) <= not(layer0_outputs(2933));
    outputs(4333) <= (layer0_outputs(3734)) xor (layer0_outputs(1831));
    outputs(4334) <= (layer0_outputs(5187)) xor (layer0_outputs(3036));
    outputs(4335) <= (layer0_outputs(6196)) xor (layer0_outputs(4757));
    outputs(4336) <= not((layer0_outputs(4400)) or (layer0_outputs(2803)));
    outputs(4337) <= (layer0_outputs(1951)) xor (layer0_outputs(5434));
    outputs(4338) <= layer0_outputs(4843);
    outputs(4339) <= layer0_outputs(2439);
    outputs(4340) <= (layer0_outputs(3162)) and not (layer0_outputs(1686));
    outputs(4341) <= (layer0_outputs(7020)) xor (layer0_outputs(3175));
    outputs(4342) <= not(layer0_outputs(4696));
    outputs(4343) <= not((layer0_outputs(7431)) or (layer0_outputs(6816)));
    outputs(4344) <= (layer0_outputs(1118)) and not (layer0_outputs(3426));
    outputs(4345) <= (layer0_outputs(1666)) and not (layer0_outputs(1001));
    outputs(4346) <= not(layer0_outputs(5699));
    outputs(4347) <= layer0_outputs(1917);
    outputs(4348) <= layer0_outputs(368);
    outputs(4349) <= (layer0_outputs(717)) or (layer0_outputs(6504));
    outputs(4350) <= (layer0_outputs(2227)) and (layer0_outputs(7072));
    outputs(4351) <= (layer0_outputs(4314)) xor (layer0_outputs(5158));
    outputs(4352) <= layer0_outputs(6773);
    outputs(4353) <= layer0_outputs(2956);
    outputs(4354) <= not(layer0_outputs(2347));
    outputs(4355) <= not(layer0_outputs(4042));
    outputs(4356) <= not(layer0_outputs(4771));
    outputs(4357) <= (layer0_outputs(5191)) xor (layer0_outputs(1941));
    outputs(4358) <= not(layer0_outputs(6553));
    outputs(4359) <= layer0_outputs(3188);
    outputs(4360) <= not(layer0_outputs(27));
    outputs(4361) <= not(layer0_outputs(5024));
    outputs(4362) <= (layer0_outputs(3923)) xor (layer0_outputs(2226));
    outputs(4363) <= not(layer0_outputs(6434)) or (layer0_outputs(6393));
    outputs(4364) <= not(layer0_outputs(2980));
    outputs(4365) <= (layer0_outputs(3975)) xor (layer0_outputs(241));
    outputs(4366) <= (layer0_outputs(6363)) or (layer0_outputs(5336));
    outputs(4367) <= (layer0_outputs(6485)) or (layer0_outputs(4719));
    outputs(4368) <= layer0_outputs(2822);
    outputs(4369) <= not(layer0_outputs(2414));
    outputs(4370) <= (layer0_outputs(6664)) and not (layer0_outputs(3254));
    outputs(4371) <= layer0_outputs(2120);
    outputs(4372) <= not(layer0_outputs(5688)) or (layer0_outputs(1994));
    outputs(4373) <= not(layer0_outputs(4421)) or (layer0_outputs(4889));
    outputs(4374) <= (layer0_outputs(6650)) and not (layer0_outputs(3130));
    outputs(4375) <= not((layer0_outputs(1254)) xor (layer0_outputs(4166)));
    outputs(4376) <= not((layer0_outputs(4790)) xor (layer0_outputs(107)));
    outputs(4377) <= (layer0_outputs(6495)) or (layer0_outputs(6337));
    outputs(4378) <= not(layer0_outputs(7493));
    outputs(4379) <= not((layer0_outputs(1951)) and (layer0_outputs(6938)));
    outputs(4380) <= not((layer0_outputs(3819)) xor (layer0_outputs(2224)));
    outputs(4381) <= layer0_outputs(3764);
    outputs(4382) <= (layer0_outputs(5973)) or (layer0_outputs(2668));
    outputs(4383) <= not((layer0_outputs(617)) xor (layer0_outputs(6031)));
    outputs(4384) <= not((layer0_outputs(2284)) and (layer0_outputs(7289)));
    outputs(4385) <= (layer0_outputs(3663)) xor (layer0_outputs(5663));
    outputs(4386) <= (layer0_outputs(7540)) and (layer0_outputs(538));
    outputs(4387) <= not(layer0_outputs(1313)) or (layer0_outputs(1474));
    outputs(4388) <= not(layer0_outputs(1465)) or (layer0_outputs(2102));
    outputs(4389) <= not(layer0_outputs(5817));
    outputs(4390) <= layer0_outputs(3531);
    outputs(4391) <= not(layer0_outputs(26));
    outputs(4392) <= (layer0_outputs(2604)) xor (layer0_outputs(2321));
    outputs(4393) <= not(layer0_outputs(6922));
    outputs(4394) <= not(layer0_outputs(4453));
    outputs(4395) <= not((layer0_outputs(6974)) xor (layer0_outputs(143)));
    outputs(4396) <= layer0_outputs(5656);
    outputs(4397) <= not(layer0_outputs(6625));
    outputs(4398) <= not(layer0_outputs(5437)) or (layer0_outputs(2208));
    outputs(4399) <= (layer0_outputs(767)) xor (layer0_outputs(1047));
    outputs(4400) <= not((layer0_outputs(5105)) xor (layer0_outputs(5568)));
    outputs(4401) <= not(layer0_outputs(5996));
    outputs(4402) <= layer0_outputs(5812);
    outputs(4403) <= (layer0_outputs(5485)) xor (layer0_outputs(864));
    outputs(4404) <= (layer0_outputs(7542)) or (layer0_outputs(5077));
    outputs(4405) <= layer0_outputs(3200);
    outputs(4406) <= (layer0_outputs(3512)) and (layer0_outputs(1574));
    outputs(4407) <= (layer0_outputs(17)) and (layer0_outputs(1935));
    outputs(4408) <= (layer0_outputs(6484)) and (layer0_outputs(7214));
    outputs(4409) <= layer0_outputs(5888);
    outputs(4410) <= layer0_outputs(503);
    outputs(4411) <= (layer0_outputs(508)) and (layer0_outputs(7061));
    outputs(4412) <= layer0_outputs(7264);
    outputs(4413) <= not(layer0_outputs(558));
    outputs(4414) <= layer0_outputs(4925);
    outputs(4415) <= (layer0_outputs(3931)) xor (layer0_outputs(6568));
    outputs(4416) <= not(layer0_outputs(1878));
    outputs(4417) <= not(layer0_outputs(557));
    outputs(4418) <= not(layer0_outputs(7067)) or (layer0_outputs(3855));
    outputs(4419) <= not((layer0_outputs(4460)) and (layer0_outputs(2603)));
    outputs(4420) <= (layer0_outputs(2274)) and (layer0_outputs(3472));
    outputs(4421) <= not(layer0_outputs(6722));
    outputs(4422) <= (layer0_outputs(7080)) or (layer0_outputs(5744));
    outputs(4423) <= not(layer0_outputs(5051)) or (layer0_outputs(4871));
    outputs(4424) <= (layer0_outputs(1679)) and not (layer0_outputs(6256));
    outputs(4425) <= not(layer0_outputs(3254));
    outputs(4426) <= not((layer0_outputs(1757)) and (layer0_outputs(7543)));
    outputs(4427) <= not((layer0_outputs(7412)) and (layer0_outputs(497)));
    outputs(4428) <= not(layer0_outputs(1223));
    outputs(4429) <= (layer0_outputs(6345)) or (layer0_outputs(1731));
    outputs(4430) <= (layer0_outputs(2948)) and not (layer0_outputs(7611));
    outputs(4431) <= layer0_outputs(5001);
    outputs(4432) <= (layer0_outputs(5772)) xor (layer0_outputs(5493));
    outputs(4433) <= (layer0_outputs(2399)) and not (layer0_outputs(6062));
    outputs(4434) <= (layer0_outputs(775)) and not (layer0_outputs(6796));
    outputs(4435) <= layer0_outputs(4126);
    outputs(4436) <= not(layer0_outputs(6590));
    outputs(4437) <= not((layer0_outputs(6779)) xor (layer0_outputs(5117)));
    outputs(4438) <= not(layer0_outputs(3248));
    outputs(4439) <= not(layer0_outputs(5412));
    outputs(4440) <= (layer0_outputs(3601)) xor (layer0_outputs(2793));
    outputs(4441) <= not(layer0_outputs(4325));
    outputs(4442) <= layer0_outputs(7529);
    outputs(4443) <= layer0_outputs(5796);
    outputs(4444) <= layer0_outputs(4491);
    outputs(4445) <= not((layer0_outputs(2740)) xor (layer0_outputs(3329)));
    outputs(4446) <= layer0_outputs(4190);
    outputs(4447) <= layer0_outputs(2471);
    outputs(4448) <= (layer0_outputs(5921)) xor (layer0_outputs(756));
    outputs(4449) <= not(layer0_outputs(4385));
    outputs(4450) <= not(layer0_outputs(1816)) or (layer0_outputs(2754));
    outputs(4451) <= (layer0_outputs(5344)) xor (layer0_outputs(2183));
    outputs(4452) <= not(layer0_outputs(5316));
    outputs(4453) <= not((layer0_outputs(158)) xor (layer0_outputs(1214)));
    outputs(4454) <= not(layer0_outputs(4905));
    outputs(4455) <= (layer0_outputs(3771)) and (layer0_outputs(37));
    outputs(4456) <= not((layer0_outputs(906)) and (layer0_outputs(4846)));
    outputs(4457) <= (layer0_outputs(6511)) and (layer0_outputs(269));
    outputs(4458) <= not(layer0_outputs(5758));
    outputs(4459) <= not((layer0_outputs(190)) or (layer0_outputs(6996)));
    outputs(4460) <= not((layer0_outputs(1667)) xor (layer0_outputs(1467)));
    outputs(4461) <= layer0_outputs(56);
    outputs(4462) <= not(layer0_outputs(4313));
    outputs(4463) <= (layer0_outputs(2614)) xor (layer0_outputs(5089));
    outputs(4464) <= not((layer0_outputs(6390)) xor (layer0_outputs(6745)));
    outputs(4465) <= (layer0_outputs(6407)) and not (layer0_outputs(4443));
    outputs(4466) <= (layer0_outputs(7147)) and (layer0_outputs(5321));
    outputs(4467) <= layer0_outputs(6307);
    outputs(4468) <= not(layer0_outputs(7136));
    outputs(4469) <= not(layer0_outputs(6788));
    outputs(4470) <= (layer0_outputs(4369)) xor (layer0_outputs(5415));
    outputs(4471) <= not((layer0_outputs(5704)) or (layer0_outputs(2718)));
    outputs(4472) <= not((layer0_outputs(4863)) or (layer0_outputs(2387)));
    outputs(4473) <= not(layer0_outputs(4954));
    outputs(4474) <= (layer0_outputs(7660)) or (layer0_outputs(1579));
    outputs(4475) <= layer0_outputs(6750);
    outputs(4476) <= layer0_outputs(2499);
    outputs(4477) <= layer0_outputs(4483);
    outputs(4478) <= not(layer0_outputs(1824));
    outputs(4479) <= not(layer0_outputs(6432)) or (layer0_outputs(2235));
    outputs(4480) <= not(layer0_outputs(6996)) or (layer0_outputs(1829));
    outputs(4481) <= not((layer0_outputs(5183)) xor (layer0_outputs(2528)));
    outputs(4482) <= layer0_outputs(5091);
    outputs(4483) <= (layer0_outputs(6063)) xor (layer0_outputs(2751));
    outputs(4484) <= (layer0_outputs(1993)) and (layer0_outputs(2654));
    outputs(4485) <= not(layer0_outputs(3455));
    outputs(4486) <= (layer0_outputs(6659)) and (layer0_outputs(4532));
    outputs(4487) <= not(layer0_outputs(6398));
    outputs(4488) <= not(layer0_outputs(7668));
    outputs(4489) <= not((layer0_outputs(1647)) xor (layer0_outputs(4707)));
    outputs(4490) <= not(layer0_outputs(2691));
    outputs(4491) <= layer0_outputs(4519);
    outputs(4492) <= layer0_outputs(6507);
    outputs(4493) <= layer0_outputs(3287);
    outputs(4494) <= not((layer0_outputs(3361)) xor (layer0_outputs(2250)));
    outputs(4495) <= not(layer0_outputs(1166));
    outputs(4496) <= (layer0_outputs(5919)) or (layer0_outputs(2907));
    outputs(4497) <= not((layer0_outputs(833)) xor (layer0_outputs(3696)));
    outputs(4498) <= (layer0_outputs(5160)) and not (layer0_outputs(6107));
    outputs(4499) <= not(layer0_outputs(1645));
    outputs(4500) <= not(layer0_outputs(3831));
    outputs(4501) <= (layer0_outputs(5433)) xor (layer0_outputs(4384));
    outputs(4502) <= not(layer0_outputs(5259));
    outputs(4503) <= layer0_outputs(2120);
    outputs(4504) <= (layer0_outputs(182)) and (layer0_outputs(4582));
    outputs(4505) <= not(layer0_outputs(1822));
    outputs(4506) <= not((layer0_outputs(1447)) xor (layer0_outputs(4536)));
    outputs(4507) <= layer0_outputs(525);
    outputs(4508) <= not(layer0_outputs(2061));
    outputs(4509) <= layer0_outputs(643);
    outputs(4510) <= (layer0_outputs(6276)) xor (layer0_outputs(504));
    outputs(4511) <= not(layer0_outputs(4597)) or (layer0_outputs(1524));
    outputs(4512) <= layer0_outputs(3404);
    outputs(4513) <= (layer0_outputs(666)) and (layer0_outputs(5617));
    outputs(4514) <= (layer0_outputs(2486)) and not (layer0_outputs(6080));
    outputs(4515) <= not(layer0_outputs(535));
    outputs(4516) <= layer0_outputs(5314);
    outputs(4517) <= (layer0_outputs(905)) xor (layer0_outputs(1693));
    outputs(4518) <= layer0_outputs(5925);
    outputs(4519) <= not((layer0_outputs(2508)) xor (layer0_outputs(1832)));
    outputs(4520) <= not(layer0_outputs(710));
    outputs(4521) <= (layer0_outputs(6523)) and (layer0_outputs(3373));
    outputs(4522) <= (layer0_outputs(6135)) and not (layer0_outputs(3537));
    outputs(4523) <= not(layer0_outputs(4619));
    outputs(4524) <= not((layer0_outputs(6559)) xor (layer0_outputs(3276)));
    outputs(4525) <= layer0_outputs(2919);
    outputs(4526) <= not((layer0_outputs(228)) and (layer0_outputs(4846)));
    outputs(4527) <= layer0_outputs(3440);
    outputs(4528) <= (layer0_outputs(980)) or (layer0_outputs(4748));
    outputs(4529) <= not((layer0_outputs(3766)) xor (layer0_outputs(7570)));
    outputs(4530) <= not(layer0_outputs(6049));
    outputs(4531) <= layer0_outputs(7302);
    outputs(4532) <= layer0_outputs(696);
    outputs(4533) <= not(layer0_outputs(6404));
    outputs(4534) <= not(layer0_outputs(3085));
    outputs(4535) <= not(layer0_outputs(3319)) or (layer0_outputs(2056));
    outputs(4536) <= layer0_outputs(3418);
    outputs(4537) <= layer0_outputs(2179);
    outputs(4538) <= not(layer0_outputs(6896)) or (layer0_outputs(6660));
    outputs(4539) <= layer0_outputs(1977);
    outputs(4540) <= (layer0_outputs(6379)) and not (layer0_outputs(6531));
    outputs(4541) <= not((layer0_outputs(5283)) xor (layer0_outputs(135)));
    outputs(4542) <= layer0_outputs(5590);
    outputs(4543) <= not(layer0_outputs(3588)) or (layer0_outputs(2820));
    outputs(4544) <= not((layer0_outputs(3334)) or (layer0_outputs(751)));
    outputs(4545) <= not(layer0_outputs(6944));
    outputs(4546) <= not(layer0_outputs(6806));
    outputs(4547) <= (layer0_outputs(1279)) xor (layer0_outputs(7235));
    outputs(4548) <= not(layer0_outputs(7435));
    outputs(4549) <= not(layer0_outputs(7023));
    outputs(4550) <= layer0_outputs(5030);
    outputs(4551) <= (layer0_outputs(1515)) and not (layer0_outputs(4644));
    outputs(4552) <= not(layer0_outputs(3681));
    outputs(4553) <= layer0_outputs(7122);
    outputs(4554) <= layer0_outputs(2306);
    outputs(4555) <= not(layer0_outputs(6010));
    outputs(4556) <= (layer0_outputs(1832)) xor (layer0_outputs(4273));
    outputs(4557) <= layer0_outputs(665);
    outputs(4558) <= not((layer0_outputs(3416)) and (layer0_outputs(6968)));
    outputs(4559) <= not((layer0_outputs(5571)) or (layer0_outputs(6605)));
    outputs(4560) <= not(layer0_outputs(705));
    outputs(4561) <= not(layer0_outputs(4970));
    outputs(4562) <= layer0_outputs(748);
    outputs(4563) <= not((layer0_outputs(4759)) and (layer0_outputs(4785)));
    outputs(4564) <= layer0_outputs(7137);
    outputs(4565) <= not((layer0_outputs(3993)) xor (layer0_outputs(4728)));
    outputs(4566) <= not((layer0_outputs(2989)) xor (layer0_outputs(1170)));
    outputs(4567) <= layer0_outputs(3430);
    outputs(4568) <= not(layer0_outputs(1223));
    outputs(4569) <= not((layer0_outputs(423)) xor (layer0_outputs(2104)));
    outputs(4570) <= not(layer0_outputs(6950));
    outputs(4571) <= not((layer0_outputs(4735)) or (layer0_outputs(6164)));
    outputs(4572) <= not(layer0_outputs(7664));
    outputs(4573) <= not(layer0_outputs(2816));
    outputs(4574) <= not((layer0_outputs(3463)) xor (layer0_outputs(1077)));
    outputs(4575) <= layer0_outputs(2742);
    outputs(4576) <= not(layer0_outputs(267));
    outputs(4577) <= layer0_outputs(492);
    outputs(4578) <= (layer0_outputs(595)) and not (layer0_outputs(5157));
    outputs(4579) <= not(layer0_outputs(3699)) or (layer0_outputs(1));
    outputs(4580) <= layer0_outputs(1755);
    outputs(4581) <= not(layer0_outputs(445));
    outputs(4582) <= (layer0_outputs(320)) xor (layer0_outputs(774));
    outputs(4583) <= (layer0_outputs(2504)) xor (layer0_outputs(4498));
    outputs(4584) <= not(layer0_outputs(6851));
    outputs(4585) <= not((layer0_outputs(5260)) xor (layer0_outputs(2639)));
    outputs(4586) <= layer0_outputs(7387);
    outputs(4587) <= (layer0_outputs(6833)) xor (layer0_outputs(1692));
    outputs(4588) <= not(layer0_outputs(2692));
    outputs(4589) <= (layer0_outputs(4779)) xor (layer0_outputs(3993));
    outputs(4590) <= layer0_outputs(2679);
    outputs(4591) <= layer0_outputs(7616);
    outputs(4592) <= not(layer0_outputs(5015));
    outputs(4593) <= not((layer0_outputs(7275)) or (layer0_outputs(7240)));
    outputs(4594) <= not((layer0_outputs(7521)) xor (layer0_outputs(2062)));
    outputs(4595) <= not(layer0_outputs(4289));
    outputs(4596) <= not(layer0_outputs(1409));
    outputs(4597) <= (layer0_outputs(1486)) and not (layer0_outputs(2509));
    outputs(4598) <= layer0_outputs(2271);
    outputs(4599) <= layer0_outputs(2922);
    outputs(4600) <= layer0_outputs(6166);
    outputs(4601) <= (layer0_outputs(465)) and not (layer0_outputs(3915));
    outputs(4602) <= layer0_outputs(1861);
    outputs(4603) <= (layer0_outputs(7058)) and not (layer0_outputs(4952));
    outputs(4604) <= layer0_outputs(5140);
    outputs(4605) <= not(layer0_outputs(2788));
    outputs(4606) <= not(layer0_outputs(3389));
    outputs(4607) <= not((layer0_outputs(1134)) xor (layer0_outputs(1887)));
    outputs(4608) <= not((layer0_outputs(3439)) and (layer0_outputs(4965)));
    outputs(4609) <= not(layer0_outputs(6439));
    outputs(4610) <= not(layer0_outputs(3551)) or (layer0_outputs(2505));
    outputs(4611) <= (layer0_outputs(4274)) and not (layer0_outputs(7079));
    outputs(4612) <= not(layer0_outputs(3646));
    outputs(4613) <= not(layer0_outputs(330));
    outputs(4614) <= layer0_outputs(5256);
    outputs(4615) <= not(layer0_outputs(3377));
    outputs(4616) <= not(layer0_outputs(3013));
    outputs(4617) <= layer0_outputs(7006);
    outputs(4618) <= layer0_outputs(1454);
    outputs(4619) <= (layer0_outputs(5654)) and (layer0_outputs(4261));
    outputs(4620) <= not(layer0_outputs(2167)) or (layer0_outputs(5173));
    outputs(4621) <= (layer0_outputs(2775)) and not (layer0_outputs(5760));
    outputs(4622) <= not((layer0_outputs(2003)) xor (layer0_outputs(799)));
    outputs(4623) <= layer0_outputs(4216);
    outputs(4624) <= not(layer0_outputs(1172)) or (layer0_outputs(6953));
    outputs(4625) <= not(layer0_outputs(248));
    outputs(4626) <= not(layer0_outputs(4652)) or (layer0_outputs(2166));
    outputs(4627) <= not(layer0_outputs(1492));
    outputs(4628) <= not(layer0_outputs(3650));
    outputs(4629) <= (layer0_outputs(7451)) or (layer0_outputs(3363));
    outputs(4630) <= not(layer0_outputs(3823));
    outputs(4631) <= layer0_outputs(2511);
    outputs(4632) <= not((layer0_outputs(3585)) or (layer0_outputs(5063)));
    outputs(4633) <= not(layer0_outputs(5840)) or (layer0_outputs(4407));
    outputs(4634) <= (layer0_outputs(5859)) and not (layer0_outputs(7429));
    outputs(4635) <= not(layer0_outputs(3959)) or (layer0_outputs(922));
    outputs(4636) <= not(layer0_outputs(6200));
    outputs(4637) <= (layer0_outputs(6575)) and (layer0_outputs(6982));
    outputs(4638) <= not(layer0_outputs(451));
    outputs(4639) <= layer0_outputs(1462);
    outputs(4640) <= (layer0_outputs(6990)) and not (layer0_outputs(2894));
    outputs(4641) <= not(layer0_outputs(6995));
    outputs(4642) <= (layer0_outputs(141)) and not (layer0_outputs(4218));
    outputs(4643) <= not((layer0_outputs(5932)) or (layer0_outputs(1125)));
    outputs(4644) <= not(layer0_outputs(501));
    outputs(4645) <= (layer0_outputs(7236)) and not (layer0_outputs(2436));
    outputs(4646) <= (layer0_outputs(7371)) and not (layer0_outputs(3084));
    outputs(4647) <= layer0_outputs(3500);
    outputs(4648) <= layer0_outputs(4864);
    outputs(4649) <= not(layer0_outputs(6469));
    outputs(4650) <= not(layer0_outputs(1052));
    outputs(4651) <= layer0_outputs(4352);
    outputs(4652) <= not(layer0_outputs(2693)) or (layer0_outputs(4966));
    outputs(4653) <= not(layer0_outputs(6646));
    outputs(4654) <= (layer0_outputs(1272)) and not (layer0_outputs(3942));
    outputs(4655) <= not(layer0_outputs(1790));
    outputs(4656) <= not((layer0_outputs(4244)) or (layer0_outputs(6923)));
    outputs(4657) <= not((layer0_outputs(6794)) or (layer0_outputs(6556)));
    outputs(4658) <= not(layer0_outputs(523)) or (layer0_outputs(5118));
    outputs(4659) <= not((layer0_outputs(2247)) xor (layer0_outputs(4804)));
    outputs(4660) <= layer0_outputs(6324);
    outputs(4661) <= not(layer0_outputs(5098));
    outputs(4662) <= layer0_outputs(2562);
    outputs(4663) <= (layer0_outputs(7014)) xor (layer0_outputs(552));
    outputs(4664) <= not(layer0_outputs(2469));
    outputs(4665) <= not(layer0_outputs(6368));
    outputs(4666) <= (layer0_outputs(6403)) and not (layer0_outputs(6534));
    outputs(4667) <= layer0_outputs(2776);
    outputs(4668) <= not(layer0_outputs(7198));
    outputs(4669) <= layer0_outputs(3292);
    outputs(4670) <= (layer0_outputs(5116)) and not (layer0_outputs(1211));
    outputs(4671) <= not(layer0_outputs(7396)) or (layer0_outputs(241));
    outputs(4672) <= not(layer0_outputs(4666));
    outputs(4673) <= (layer0_outputs(5204)) and not (layer0_outputs(7492));
    outputs(4674) <= (layer0_outputs(1945)) and not (layer0_outputs(1868));
    outputs(4675) <= layer0_outputs(5997);
    outputs(4676) <= not(layer0_outputs(798));
    outputs(4677) <= not((layer0_outputs(6083)) or (layer0_outputs(5126)));
    outputs(4678) <= layer0_outputs(3281);
    outputs(4679) <= not(layer0_outputs(2199));
    outputs(4680) <= not(layer0_outputs(1664));
    outputs(4681) <= not(layer0_outputs(3498));
    outputs(4682) <= not((layer0_outputs(3644)) and (layer0_outputs(3824)));
    outputs(4683) <= not(layer0_outputs(1617));
    outputs(4684) <= not(layer0_outputs(761));
    outputs(4685) <= (layer0_outputs(2706)) and not (layer0_outputs(5721));
    outputs(4686) <= (layer0_outputs(4135)) and (layer0_outputs(5621));
    outputs(4687) <= (layer0_outputs(3563)) xor (layer0_outputs(70));
    outputs(4688) <= layer0_outputs(6558);
    outputs(4689) <= (layer0_outputs(42)) and (layer0_outputs(1565));
    outputs(4690) <= layer0_outputs(2926);
    outputs(4691) <= (layer0_outputs(2669)) and (layer0_outputs(4678));
    outputs(4692) <= (layer0_outputs(4894)) and not (layer0_outputs(5952));
    outputs(4693) <= (layer0_outputs(2984)) and not (layer0_outputs(7087));
    outputs(4694) <= layer0_outputs(5948);
    outputs(4695) <= (layer0_outputs(1810)) and not (layer0_outputs(5918));
    outputs(4696) <= not(layer0_outputs(197)) or (layer0_outputs(2659));
    outputs(4697) <= not(layer0_outputs(3567));
    outputs(4698) <= not(layer0_outputs(200));
    outputs(4699) <= not(layer0_outputs(6429));
    outputs(4700) <= layer0_outputs(6713);
    outputs(4701) <= not(layer0_outputs(6320));
    outputs(4702) <= not((layer0_outputs(3445)) and (layer0_outputs(4266)));
    outputs(4703) <= not((layer0_outputs(3587)) xor (layer0_outputs(1684)));
    outputs(4704) <= layer0_outputs(2547);
    outputs(4705) <= (layer0_outputs(341)) and not (layer0_outputs(6048));
    outputs(4706) <= layer0_outputs(3279);
    outputs(4707) <= (layer0_outputs(4176)) and (layer0_outputs(1936));
    outputs(4708) <= layer0_outputs(5285);
    outputs(4709) <= (layer0_outputs(3236)) and not (layer0_outputs(4633));
    outputs(4710) <= (layer0_outputs(1858)) xor (layer0_outputs(2069));
    outputs(4711) <= not(layer0_outputs(3466));
    outputs(4712) <= (layer0_outputs(3675)) and not (layer0_outputs(2218));
    outputs(4713) <= layer0_outputs(2857);
    outputs(4714) <= layer0_outputs(3414);
    outputs(4715) <= not((layer0_outputs(6253)) or (layer0_outputs(5089)));
    outputs(4716) <= (layer0_outputs(1705)) and not (layer0_outputs(496));
    outputs(4717) <= not(layer0_outputs(2814));
    outputs(4718) <= layer0_outputs(4359);
    outputs(4719) <= not(layer0_outputs(5078));
    outputs(4720) <= not((layer0_outputs(4642)) or (layer0_outputs(1379)));
    outputs(4721) <= not(layer0_outputs(6758));
    outputs(4722) <= not(layer0_outputs(6730));
    outputs(4723) <= (layer0_outputs(4160)) and not (layer0_outputs(5083));
    outputs(4724) <= not(layer0_outputs(4560));
    outputs(4725) <= not(layer0_outputs(2326));
    outputs(4726) <= not(layer0_outputs(7612));
    outputs(4727) <= not(layer0_outputs(4543));
    outputs(4728) <= (layer0_outputs(2811)) and not (layer0_outputs(6092));
    outputs(4729) <= layer0_outputs(177);
    outputs(4730) <= not((layer0_outputs(2463)) or (layer0_outputs(6626)));
    outputs(4731) <= not(layer0_outputs(6705));
    outputs(4732) <= layer0_outputs(1495);
    outputs(4733) <= not((layer0_outputs(6643)) or (layer0_outputs(209)));
    outputs(4734) <= (layer0_outputs(2160)) and not (layer0_outputs(266));
    outputs(4735) <= (layer0_outputs(5418)) and not (layer0_outputs(6048));
    outputs(4736) <= layer0_outputs(6611);
    outputs(4737) <= not((layer0_outputs(6637)) and (layer0_outputs(5210)));
    outputs(4738) <= not(layer0_outputs(187)) or (layer0_outputs(4375));
    outputs(4739) <= not(layer0_outputs(931));
    outputs(4740) <= layer0_outputs(5793);
    outputs(4741) <= (layer0_outputs(3286)) xor (layer0_outputs(538));
    outputs(4742) <= layer0_outputs(3908);
    outputs(4743) <= layer0_outputs(4910);
    outputs(4744) <= not((layer0_outputs(3300)) xor (layer0_outputs(4044)));
    outputs(4745) <= not(layer0_outputs(6590));
    outputs(4746) <= (layer0_outputs(581)) xor (layer0_outputs(61));
    outputs(4747) <= not(layer0_outputs(3488));
    outputs(4748) <= not((layer0_outputs(6047)) or (layer0_outputs(1441)));
    outputs(4749) <= layer0_outputs(4484);
    outputs(4750) <= not(layer0_outputs(4599));
    outputs(4751) <= layer0_outputs(4212);
    outputs(4752) <= not(layer0_outputs(6806));
    outputs(4753) <= not(layer0_outputs(4802));
    outputs(4754) <= not(layer0_outputs(4570));
    outputs(4755) <= layer0_outputs(4976);
    outputs(4756) <= layer0_outputs(1407);
    outputs(4757) <= not(layer0_outputs(1852));
    outputs(4758) <= layer0_outputs(5555);
    outputs(4759) <= not(layer0_outputs(4522)) or (layer0_outputs(366));
    outputs(4760) <= not(layer0_outputs(536));
    outputs(4761) <= layer0_outputs(2541);
    outputs(4762) <= layer0_outputs(3952);
    outputs(4763) <= (layer0_outputs(918)) xor (layer0_outputs(6960));
    outputs(4764) <= layer0_outputs(2094);
    outputs(4765) <= (layer0_outputs(92)) and (layer0_outputs(3027));
    outputs(4766) <= (layer0_outputs(5916)) and (layer0_outputs(2776));
    outputs(4767) <= not(layer0_outputs(4814));
    outputs(4768) <= not((layer0_outputs(4337)) or (layer0_outputs(6205)));
    outputs(4769) <= (layer0_outputs(4227)) and not (layer0_outputs(5669));
    outputs(4770) <= (layer0_outputs(4942)) xor (layer0_outputs(7367));
    outputs(4771) <= (layer0_outputs(5979)) and not (layer0_outputs(5133));
    outputs(4772) <= not(layer0_outputs(1238)) or (layer0_outputs(6653));
    outputs(4773) <= (layer0_outputs(193)) and not (layer0_outputs(2727));
    outputs(4774) <= (layer0_outputs(19)) or (layer0_outputs(2154));
    outputs(4775) <= not((layer0_outputs(1864)) xor (layer0_outputs(5119)));
    outputs(4776) <= not(layer0_outputs(971));
    outputs(4777) <= layer0_outputs(1736);
    outputs(4778) <= not(layer0_outputs(5163));
    outputs(4779) <= not((layer0_outputs(6899)) or (layer0_outputs(3805)));
    outputs(4780) <= layer0_outputs(648);
    outputs(4781) <= not(layer0_outputs(3487));
    outputs(4782) <= not(layer0_outputs(6249));
    outputs(4783) <= layer0_outputs(4001);
    outputs(4784) <= not(layer0_outputs(248));
    outputs(4785) <= not(layer0_outputs(2533));
    outputs(4786) <= layer0_outputs(6006);
    outputs(4787) <= layer0_outputs(5545);
    outputs(4788) <= not(layer0_outputs(701));
    outputs(4789) <= layer0_outputs(2808);
    outputs(4790) <= not(layer0_outputs(5938));
    outputs(4791) <= (layer0_outputs(1907)) and not (layer0_outputs(4822));
    outputs(4792) <= not(layer0_outputs(3558));
    outputs(4793) <= layer0_outputs(2493);
    outputs(4794) <= not(layer0_outputs(2207));
    outputs(4795) <= not((layer0_outputs(2836)) or (layer0_outputs(763)));
    outputs(4796) <= not(layer0_outputs(351));
    outputs(4797) <= not(layer0_outputs(1707));
    outputs(4798) <= not(layer0_outputs(1260)) or (layer0_outputs(4506));
    outputs(4799) <= (layer0_outputs(1367)) and not (layer0_outputs(5785));
    outputs(4800) <= not(layer0_outputs(4733));
    outputs(4801) <= not((layer0_outputs(5044)) or (layer0_outputs(4102)));
    outputs(4802) <= (layer0_outputs(3741)) or (layer0_outputs(6020));
    outputs(4803) <= layer0_outputs(5730);
    outputs(4804) <= layer0_outputs(561);
    outputs(4805) <= (layer0_outputs(2510)) xor (layer0_outputs(2680));
    outputs(4806) <= (layer0_outputs(4216)) and not (layer0_outputs(5143));
    outputs(4807) <= layer0_outputs(1215);
    outputs(4808) <= (layer0_outputs(6865)) xor (layer0_outputs(7537));
    outputs(4809) <= layer0_outputs(625);
    outputs(4810) <= not((layer0_outputs(6721)) xor (layer0_outputs(7389)));
    outputs(4811) <= not((layer0_outputs(1362)) or (layer0_outputs(2394)));
    outputs(4812) <= (layer0_outputs(4109)) and not (layer0_outputs(3301));
    outputs(4813) <= not((layer0_outputs(4007)) xor (layer0_outputs(4674)));
    outputs(4814) <= not(layer0_outputs(4373)) or (layer0_outputs(2373));
    outputs(4815) <= layer0_outputs(671);
    outputs(4816) <= layer0_outputs(42);
    outputs(4817) <= not(layer0_outputs(441));
    outputs(4818) <= not(layer0_outputs(3582));
    outputs(4819) <= not((layer0_outputs(4032)) or (layer0_outputs(4934)));
    outputs(4820) <= layer0_outputs(4622);
    outputs(4821) <= (layer0_outputs(5640)) and not (layer0_outputs(2232));
    outputs(4822) <= (layer0_outputs(3165)) or (layer0_outputs(6094));
    outputs(4823) <= (layer0_outputs(1199)) and (layer0_outputs(3425));
    outputs(4824) <= layer0_outputs(5312);
    outputs(4825) <= (layer0_outputs(160)) xor (layer0_outputs(5983));
    outputs(4826) <= (layer0_outputs(4302)) and not (layer0_outputs(7511));
    outputs(4827) <= layer0_outputs(7599);
    outputs(4828) <= not((layer0_outputs(937)) and (layer0_outputs(2210)));
    outputs(4829) <= not(layer0_outputs(6928));
    outputs(4830) <= not(layer0_outputs(6947));
    outputs(4831) <= layer0_outputs(6523);
    outputs(4832) <= (layer0_outputs(3555)) and not (layer0_outputs(7196));
    outputs(4833) <= not(layer0_outputs(2496));
    outputs(4834) <= not(layer0_outputs(209));
    outputs(4835) <= not((layer0_outputs(7620)) or (layer0_outputs(4125)));
    outputs(4836) <= (layer0_outputs(6649)) and not (layer0_outputs(6519));
    outputs(4837) <= layer0_outputs(6612);
    outputs(4838) <= not((layer0_outputs(3548)) or (layer0_outputs(2111)));
    outputs(4839) <= layer0_outputs(563);
    outputs(4840) <= (layer0_outputs(1298)) and (layer0_outputs(1135));
    outputs(4841) <= (layer0_outputs(5261)) xor (layer0_outputs(4711));
    outputs(4842) <= layer0_outputs(2157);
    outputs(4843) <= not((layer0_outputs(2665)) and (layer0_outputs(1040)));
    outputs(4844) <= layer0_outputs(5284);
    outputs(4845) <= layer0_outputs(6106);
    outputs(4846) <= not((layer0_outputs(1124)) xor (layer0_outputs(6197)));
    outputs(4847) <= layer0_outputs(2415);
    outputs(4848) <= (layer0_outputs(6527)) xor (layer0_outputs(6605));
    outputs(4849) <= layer0_outputs(267);
    outputs(4850) <= not(layer0_outputs(2180));
    outputs(4851) <= (layer0_outputs(6326)) xor (layer0_outputs(1356));
    outputs(4852) <= (layer0_outputs(2428)) and not (layer0_outputs(5739));
    outputs(4853) <= (layer0_outputs(6747)) and not (layer0_outputs(4031));
    outputs(4854) <= not(layer0_outputs(5334));
    outputs(4855) <= layer0_outputs(3983);
    outputs(4856) <= (layer0_outputs(203)) and not (layer0_outputs(1741));
    outputs(4857) <= layer0_outputs(6748);
    outputs(4858) <= (layer0_outputs(4758)) and not (layer0_outputs(1278));
    outputs(4859) <= (layer0_outputs(1113)) and not (layer0_outputs(1603));
    outputs(4860) <= (layer0_outputs(7037)) and not (layer0_outputs(3464));
    outputs(4861) <= layer0_outputs(6232);
    outputs(4862) <= not(layer0_outputs(3491)) or (layer0_outputs(7046));
    outputs(4863) <= layer0_outputs(6573);
    outputs(4864) <= (layer0_outputs(928)) xor (layer0_outputs(646));
    outputs(4865) <= not(layer0_outputs(6210));
    outputs(4866) <= not(layer0_outputs(5500));
    outputs(4867) <= not((layer0_outputs(820)) or (layer0_outputs(2643)));
    outputs(4868) <= layer0_outputs(1019);
    outputs(4869) <= (layer0_outputs(2185)) and not (layer0_outputs(3624));
    outputs(4870) <= (layer0_outputs(1519)) and not (layer0_outputs(6393));
    outputs(4871) <= not(layer0_outputs(1783));
    outputs(4872) <= layer0_outputs(6215);
    outputs(4873) <= (layer0_outputs(6898)) and not (layer0_outputs(1186));
    outputs(4874) <= layer0_outputs(2245);
    outputs(4875) <= not(layer0_outputs(2196));
    outputs(4876) <= not(layer0_outputs(4592)) or (layer0_outputs(7271));
    outputs(4877) <= not((layer0_outputs(3211)) xor (layer0_outputs(4614)));
    outputs(4878) <= layer0_outputs(3688);
    outputs(4879) <= (layer0_outputs(392)) or (layer0_outputs(2539));
    outputs(4880) <= layer0_outputs(6287);
    outputs(4881) <= (layer0_outputs(3328)) or (layer0_outputs(38));
    outputs(4882) <= layer0_outputs(225);
    outputs(4883) <= not((layer0_outputs(4934)) or (layer0_outputs(5797)));
    outputs(4884) <= not(layer0_outputs(66));
    outputs(4885) <= not((layer0_outputs(7593)) xor (layer0_outputs(449)));
    outputs(4886) <= (layer0_outputs(4374)) and not (layer0_outputs(3727));
    outputs(4887) <= (layer0_outputs(295)) and (layer0_outputs(885));
    outputs(4888) <= (layer0_outputs(2777)) xor (layer0_outputs(34));
    outputs(4889) <= (layer0_outputs(2309)) xor (layer0_outputs(4725));
    outputs(4890) <= not(layer0_outputs(2875));
    outputs(4891) <= not(layer0_outputs(827));
    outputs(4892) <= not((layer0_outputs(7405)) and (layer0_outputs(2664)));
    outputs(4893) <= not((layer0_outputs(6406)) xor (layer0_outputs(4103)));
    outputs(4894) <= (layer0_outputs(3094)) xor (layer0_outputs(6741));
    outputs(4895) <= (layer0_outputs(5560)) and (layer0_outputs(6686));
    outputs(4896) <= (layer0_outputs(1375)) xor (layer0_outputs(18));
    outputs(4897) <= not(layer0_outputs(47));
    outputs(4898) <= layer0_outputs(1968);
    outputs(4899) <= not(layer0_outputs(23));
    outputs(4900) <= (layer0_outputs(3530)) and not (layer0_outputs(6241));
    outputs(4901) <= (layer0_outputs(4994)) and not (layer0_outputs(3942));
    outputs(4902) <= not(layer0_outputs(5813)) or (layer0_outputs(885));
    outputs(4903) <= not(layer0_outputs(3343));
    outputs(4904) <= layer0_outputs(4405);
    outputs(4905) <= layer0_outputs(1497);
    outputs(4906) <= not((layer0_outputs(1618)) xor (layer0_outputs(4142)));
    outputs(4907) <= not(layer0_outputs(943));
    outputs(4908) <= not(layer0_outputs(3253));
    outputs(4909) <= (layer0_outputs(427)) and not (layer0_outputs(5218));
    outputs(4910) <= layer0_outputs(1529);
    outputs(4911) <= not((layer0_outputs(110)) xor (layer0_outputs(5696)));
    outputs(4912) <= not(layer0_outputs(2357));
    outputs(4913) <= layer0_outputs(5872);
    outputs(4914) <= not(layer0_outputs(3435));
    outputs(4915) <= not((layer0_outputs(3515)) and (layer0_outputs(5245)));
    outputs(4916) <= not((layer0_outputs(3746)) or (layer0_outputs(6850)));
    outputs(4917) <= layer0_outputs(7250);
    outputs(4918) <= not(layer0_outputs(7433));
    outputs(4919) <= (layer0_outputs(5916)) and not (layer0_outputs(3084));
    outputs(4920) <= not(layer0_outputs(5492));
    outputs(4921) <= not(layer0_outputs(3516));
    outputs(4922) <= layer0_outputs(2172);
    outputs(4923) <= not((layer0_outputs(1428)) xor (layer0_outputs(2180)));
    outputs(4924) <= (layer0_outputs(549)) and (layer0_outputs(2165));
    outputs(4925) <= not(layer0_outputs(7258)) or (layer0_outputs(1502));
    outputs(4926) <= layer0_outputs(2466);
    outputs(4927) <= layer0_outputs(4494);
    outputs(4928) <= layer0_outputs(4926);
    outputs(4929) <= (layer0_outputs(5471)) or (layer0_outputs(580));
    outputs(4930) <= not(layer0_outputs(253));
    outputs(4931) <= layer0_outputs(2390);
    outputs(4932) <= (layer0_outputs(4477)) and not (layer0_outputs(2097));
    outputs(4933) <= not(layer0_outputs(6991));
    outputs(4934) <= (layer0_outputs(7247)) and (layer0_outputs(3390));
    outputs(4935) <= not((layer0_outputs(2098)) or (layer0_outputs(6225)));
    outputs(4936) <= (layer0_outputs(2715)) xor (layer0_outputs(5864));
    outputs(4937) <= (layer0_outputs(5640)) and not (layer0_outputs(4903));
    outputs(4938) <= not((layer0_outputs(2524)) and (layer0_outputs(153)));
    outputs(4939) <= (layer0_outputs(2876)) xor (layer0_outputs(2751));
    outputs(4940) <= (layer0_outputs(3169)) xor (layer0_outputs(1890));
    outputs(4941) <= not(layer0_outputs(3721));
    outputs(4942) <= not(layer0_outputs(592)) or (layer0_outputs(1207));
    outputs(4943) <= (layer0_outputs(1994)) and not (layer0_outputs(2206));
    outputs(4944) <= layer0_outputs(5791);
    outputs(4945) <= not((layer0_outputs(6208)) and (layer0_outputs(1781)));
    outputs(4946) <= (layer0_outputs(4663)) xor (layer0_outputs(2234));
    outputs(4947) <= layer0_outputs(3273);
    outputs(4948) <= (layer0_outputs(4593)) and not (layer0_outputs(477));
    outputs(4949) <= not((layer0_outputs(4973)) or (layer0_outputs(833)));
    outputs(4950) <= layer0_outputs(7490);
    outputs(4951) <= layer0_outputs(5613);
    outputs(4952) <= layer0_outputs(124);
    outputs(4953) <= (layer0_outputs(419)) and not (layer0_outputs(2434));
    outputs(4954) <= not((layer0_outputs(3163)) xor (layer0_outputs(6616)));
    outputs(4955) <= not(layer0_outputs(5627));
    outputs(4956) <= layer0_outputs(5189);
    outputs(4957) <= not(layer0_outputs(5783));
    outputs(4958) <= layer0_outputs(831);
    outputs(4959) <= (layer0_outputs(2198)) and not (layer0_outputs(1720));
    outputs(4960) <= layer0_outputs(3825);
    outputs(4961) <= not((layer0_outputs(797)) or (layer0_outputs(3833)));
    outputs(4962) <= (layer0_outputs(5444)) and not (layer0_outputs(6359));
    outputs(4963) <= layer0_outputs(818);
    outputs(4964) <= (layer0_outputs(5847)) and (layer0_outputs(1702));
    outputs(4965) <= layer0_outputs(4565);
    outputs(4966) <= layer0_outputs(4533);
    outputs(4967) <= not(layer0_outputs(6834));
    outputs(4968) <= not(layer0_outputs(4649));
    outputs(4969) <= not(layer0_outputs(2557)) or (layer0_outputs(1220));
    outputs(4970) <= (layer0_outputs(7006)) and not (layer0_outputs(3765));
    outputs(4971) <= not(layer0_outputs(3398));
    outputs(4972) <= not(layer0_outputs(2607));
    outputs(4973) <= not(layer0_outputs(3862));
    outputs(4974) <= (layer0_outputs(938)) xor (layer0_outputs(2570));
    outputs(4975) <= not((layer0_outputs(147)) xor (layer0_outputs(4567)));
    outputs(4976) <= (layer0_outputs(7008)) or (layer0_outputs(5794));
    outputs(4977) <= not(layer0_outputs(476));
    outputs(4978) <= not((layer0_outputs(3409)) or (layer0_outputs(7094)));
    outputs(4979) <= layer0_outputs(1404);
    outputs(4980) <= layer0_outputs(3668);
    outputs(4981) <= not(layer0_outputs(4265));
    outputs(4982) <= (layer0_outputs(4156)) and not (layer0_outputs(940));
    outputs(4983) <= (layer0_outputs(1516)) or (layer0_outputs(4311));
    outputs(4984) <= (layer0_outputs(1294)) and not (layer0_outputs(5055));
    outputs(4985) <= not(layer0_outputs(3979));
    outputs(4986) <= (layer0_outputs(318)) and (layer0_outputs(4594));
    outputs(4987) <= not(layer0_outputs(2966));
    outputs(4988) <= layer0_outputs(1131);
    outputs(4989) <= not((layer0_outputs(510)) or (layer0_outputs(5016)));
    outputs(4990) <= not(layer0_outputs(4666));
    outputs(4991) <= not(layer0_outputs(2310));
    outputs(4992) <= layer0_outputs(1200);
    outputs(4993) <= (layer0_outputs(2651)) xor (layer0_outputs(2772));
    outputs(4994) <= not(layer0_outputs(4924));
    outputs(4995) <= not(layer0_outputs(7169));
    outputs(4996) <= (layer0_outputs(1165)) and not (layer0_outputs(2061));
    outputs(4997) <= (layer0_outputs(4559)) and (layer0_outputs(5159));
    outputs(4998) <= layer0_outputs(202);
    outputs(4999) <= not(layer0_outputs(5614)) or (layer0_outputs(6548));
    outputs(5000) <= (layer0_outputs(6916)) and (layer0_outputs(4100));
    outputs(5001) <= (layer0_outputs(6254)) and (layer0_outputs(4214));
    outputs(5002) <= not((layer0_outputs(1606)) xor (layer0_outputs(6413)));
    outputs(5003) <= not((layer0_outputs(2454)) and (layer0_outputs(5518)));
    outputs(5004) <= not((layer0_outputs(7362)) or (layer0_outputs(3674)));
    outputs(5005) <= not(layer0_outputs(2421)) or (layer0_outputs(6597));
    outputs(5006) <= not(layer0_outputs(3318));
    outputs(5007) <= not(layer0_outputs(1380));
    outputs(5008) <= (layer0_outputs(6972)) xor (layer0_outputs(4164));
    outputs(5009) <= not(layer0_outputs(3610));
    outputs(5010) <= not((layer0_outputs(1871)) or (layer0_outputs(222)));
    outputs(5011) <= not(layer0_outputs(7087));
    outputs(5012) <= layer0_outputs(192);
    outputs(5013) <= not(layer0_outputs(5877));
    outputs(5014) <= not(layer0_outputs(5630));
    outputs(5015) <= not((layer0_outputs(5746)) xor (layer0_outputs(1941)));
    outputs(5016) <= not((layer0_outputs(4979)) or (layer0_outputs(5616)));
    outputs(5017) <= not(layer0_outputs(6951));
    outputs(5018) <= not((layer0_outputs(3371)) or (layer0_outputs(6418)));
    outputs(5019) <= layer0_outputs(6423);
    outputs(5020) <= not((layer0_outputs(4501)) xor (layer0_outputs(7134)));
    outputs(5021) <= layer0_outputs(6168);
    outputs(5022) <= (layer0_outputs(480)) and not (layer0_outputs(1290));
    outputs(5023) <= layer0_outputs(2350);
    outputs(5024) <= not(layer0_outputs(0));
    outputs(5025) <= not((layer0_outputs(2641)) or (layer0_outputs(2839)));
    outputs(5026) <= (layer0_outputs(4972)) or (layer0_outputs(5887));
    outputs(5027) <= layer0_outputs(752);
    outputs(5028) <= not(layer0_outputs(1268));
    outputs(5029) <= layer0_outputs(5700);
    outputs(5030) <= (layer0_outputs(309)) and not (layer0_outputs(5995));
    outputs(5031) <= not(layer0_outputs(4819));
    outputs(5032) <= (layer0_outputs(1451)) and (layer0_outputs(2540));
    outputs(5033) <= (layer0_outputs(1431)) and (layer0_outputs(4577));
    outputs(5034) <= not(layer0_outputs(937));
    outputs(5035) <= not(layer0_outputs(5296));
    outputs(5036) <= layer0_outputs(2258);
    outputs(5037) <= layer0_outputs(3897);
    outputs(5038) <= (layer0_outputs(3930)) and (layer0_outputs(7630));
    outputs(5039) <= (layer0_outputs(6327)) xor (layer0_outputs(6007));
    outputs(5040) <= not(layer0_outputs(3768));
    outputs(5041) <= layer0_outputs(3195);
    outputs(5042) <= layer0_outputs(5408);
    outputs(5043) <= (layer0_outputs(5476)) and not (layer0_outputs(5450));
    outputs(5044) <= not((layer0_outputs(6181)) or (layer0_outputs(4524)));
    outputs(5045) <= layer0_outputs(7248);
    outputs(5046) <= not((layer0_outputs(656)) xor (layer0_outputs(4358)));
    outputs(5047) <= not(layer0_outputs(3728));
    outputs(5048) <= layer0_outputs(4624);
    outputs(5049) <= (layer0_outputs(6939)) xor (layer0_outputs(3168));
    outputs(5050) <= not(layer0_outputs(6032));
    outputs(5051) <= not(layer0_outputs(6483));
    outputs(5052) <= not(layer0_outputs(2759));
    outputs(5053) <= (layer0_outputs(1092)) or (layer0_outputs(2827));
    outputs(5054) <= not(layer0_outputs(6190));
    outputs(5055) <= not(layer0_outputs(4436));
    outputs(5056) <= not(layer0_outputs(5624));
    outputs(5057) <= not(layer0_outputs(7116));
    outputs(5058) <= layer0_outputs(883);
    outputs(5059) <= not(layer0_outputs(3761));
    outputs(5060) <= (layer0_outputs(5313)) and not (layer0_outputs(1140));
    outputs(5061) <= layer0_outputs(1436);
    outputs(5062) <= layer0_outputs(3590);
    outputs(5063) <= (layer0_outputs(6331)) and not (layer0_outputs(4740));
    outputs(5064) <= (layer0_outputs(1023)) and not (layer0_outputs(5369));
    outputs(5065) <= not(layer0_outputs(7359));
    outputs(5066) <= layer0_outputs(3665);
    outputs(5067) <= layer0_outputs(813);
    outputs(5068) <= layer0_outputs(3424);
    outputs(5069) <= not((layer0_outputs(4716)) xor (layer0_outputs(4988)));
    outputs(5070) <= not(layer0_outputs(4517));
    outputs(5071) <= (layer0_outputs(4199)) and not (layer0_outputs(7526));
    outputs(5072) <= not((layer0_outputs(1470)) xor (layer0_outputs(3001)));
    outputs(5073) <= not((layer0_outputs(5553)) xor (layer0_outputs(3432)));
    outputs(5074) <= not((layer0_outputs(2190)) and (layer0_outputs(2760)));
    outputs(5075) <= layer0_outputs(5889);
    outputs(5076) <= (layer0_outputs(5990)) and not (layer0_outputs(125));
    outputs(5077) <= (layer0_outputs(4672)) and (layer0_outputs(6783));
    outputs(5078) <= layer0_outputs(3908);
    outputs(5079) <= not(layer0_outputs(5940)) or (layer0_outputs(2195));
    outputs(5080) <= not(layer0_outputs(6799));
    outputs(5081) <= not((layer0_outputs(7311)) xor (layer0_outputs(6828)));
    outputs(5082) <= not(layer0_outputs(6840));
    outputs(5083) <= layer0_outputs(4509);
    outputs(5084) <= not(layer0_outputs(4297));
    outputs(5085) <= not(layer0_outputs(4717)) or (layer0_outputs(619));
    outputs(5086) <= layer0_outputs(6410);
    outputs(5087) <= (layer0_outputs(649)) and not (layer0_outputs(3208));
    outputs(5088) <= (layer0_outputs(3126)) xor (layer0_outputs(5977));
    outputs(5089) <= not(layer0_outputs(7535));
    outputs(5090) <= not((layer0_outputs(2135)) and (layer0_outputs(5130)));
    outputs(5091) <= not(layer0_outputs(7474));
    outputs(5092) <= not(layer0_outputs(6908));
    outputs(5093) <= layer0_outputs(2977);
    outputs(5094) <= not(layer0_outputs(4197));
    outputs(5095) <= (layer0_outputs(855)) and not (layer0_outputs(2758));
    outputs(5096) <= layer0_outputs(3334);
    outputs(5097) <= not((layer0_outputs(6266)) xor (layer0_outputs(1675)));
    outputs(5098) <= not(layer0_outputs(7196));
    outputs(5099) <= (layer0_outputs(4981)) and not (layer0_outputs(112));
    outputs(5100) <= not(layer0_outputs(6800));
    outputs(5101) <= layer0_outputs(5176);
    outputs(5102) <= layer0_outputs(4926);
    outputs(5103) <= not((layer0_outputs(5574)) or (layer0_outputs(7679)));
    outputs(5104) <= (layer0_outputs(4612)) and (layer0_outputs(7269));
    outputs(5105) <= layer0_outputs(5198);
    outputs(5106) <= not(layer0_outputs(4293));
    outputs(5107) <= (layer0_outputs(4079)) and not (layer0_outputs(3339));
    outputs(5108) <= layer0_outputs(7038);
    outputs(5109) <= layer0_outputs(2736);
    outputs(5110) <= layer0_outputs(5560);
    outputs(5111) <= (layer0_outputs(3060)) and not (layer0_outputs(5037));
    outputs(5112) <= not(layer0_outputs(7494));
    outputs(5113) <= layer0_outputs(7418);
    outputs(5114) <= not(layer0_outputs(4937));
    outputs(5115) <= layer0_outputs(421);
    outputs(5116) <= not(layer0_outputs(3636));
    outputs(5117) <= layer0_outputs(4698);
    outputs(5118) <= layer0_outputs(1409);
    outputs(5119) <= layer0_outputs(4569);
    outputs(5120) <= not(layer0_outputs(742));
    outputs(5121) <= layer0_outputs(3411);
    outputs(5122) <= (layer0_outputs(6615)) and (layer0_outputs(7281));
    outputs(5123) <= layer0_outputs(60);
    outputs(5124) <= not(layer0_outputs(1545));
    outputs(5125) <= layer0_outputs(1227);
    outputs(5126) <= not(layer0_outputs(943));
    outputs(5127) <= not(layer0_outputs(1671));
    outputs(5128) <= (layer0_outputs(575)) and not (layer0_outputs(4818));
    outputs(5129) <= layer0_outputs(843);
    outputs(5130) <= not((layer0_outputs(7123)) xor (layer0_outputs(6706)));
    outputs(5131) <= (layer0_outputs(1285)) and not (layer0_outputs(2229));
    outputs(5132) <= (layer0_outputs(5139)) xor (layer0_outputs(3239));
    outputs(5133) <= layer0_outputs(1747);
    outputs(5134) <= layer0_outputs(3107);
    outputs(5135) <= not((layer0_outputs(4323)) or (layer0_outputs(1011)));
    outputs(5136) <= not((layer0_outputs(2236)) xor (layer0_outputs(3298)));
    outputs(5137) <= not(layer0_outputs(5268)) or (layer0_outputs(5668));
    outputs(5138) <= (layer0_outputs(1064)) or (layer0_outputs(7350));
    outputs(5139) <= (layer0_outputs(6075)) and not (layer0_outputs(2179));
    outputs(5140) <= not((layer0_outputs(3095)) xor (layer0_outputs(3837)));
    outputs(5141) <= (layer0_outputs(1983)) xor (layer0_outputs(6990));
    outputs(5142) <= layer0_outputs(942);
    outputs(5143) <= (layer0_outputs(1555)) and not (layer0_outputs(5113));
    outputs(5144) <= not((layer0_outputs(1870)) xor (layer0_outputs(6225)));
    outputs(5145) <= not((layer0_outputs(863)) xor (layer0_outputs(6187)));
    outputs(5146) <= not(layer0_outputs(311));
    outputs(5147) <= not(layer0_outputs(3344));
    outputs(5148) <= layer0_outputs(4588);
    outputs(5149) <= not((layer0_outputs(3379)) xor (layer0_outputs(4742)));
    outputs(5150) <= not((layer0_outputs(3439)) and (layer0_outputs(4545)));
    outputs(5151) <= (layer0_outputs(6242)) xor (layer0_outputs(3534));
    outputs(5152) <= (layer0_outputs(2374)) and (layer0_outputs(7132));
    outputs(5153) <= not(layer0_outputs(532));
    outputs(5154) <= not(layer0_outputs(1025));
    outputs(5155) <= not((layer0_outputs(6607)) or (layer0_outputs(5807)));
    outputs(5156) <= layer0_outputs(3590);
    outputs(5157) <= not(layer0_outputs(1340)) or (layer0_outputs(6803));
    outputs(5158) <= layer0_outputs(2241);
    outputs(5159) <= not((layer0_outputs(2672)) or (layer0_outputs(2393)));
    outputs(5160) <= not(layer0_outputs(2187));
    outputs(5161) <= layer0_outputs(6898);
    outputs(5162) <= not((layer0_outputs(356)) xor (layer0_outputs(2158)));
    outputs(5163) <= layer0_outputs(7525);
    outputs(5164) <= not(layer0_outputs(6357));
    outputs(5165) <= not((layer0_outputs(3051)) or (layer0_outputs(3527)));
    outputs(5166) <= not(layer0_outputs(529));
    outputs(5167) <= not((layer0_outputs(3863)) or (layer0_outputs(3885)));
    outputs(5168) <= not(layer0_outputs(1355));
    outputs(5169) <= layer0_outputs(3675);
    outputs(5170) <= not(layer0_outputs(953));
    outputs(5171) <= not(layer0_outputs(2915));
    outputs(5172) <= layer0_outputs(6861);
    outputs(5173) <= (layer0_outputs(4206)) and not (layer0_outputs(1548));
    outputs(5174) <= not((layer0_outputs(737)) xor (layer0_outputs(734)));
    outputs(5175) <= layer0_outputs(7048);
    outputs(5176) <= not((layer0_outputs(2546)) and (layer0_outputs(523)));
    outputs(5177) <= layer0_outputs(3729);
    outputs(5178) <= not((layer0_outputs(3044)) or (layer0_outputs(1325)));
    outputs(5179) <= not((layer0_outputs(1129)) xor (layer0_outputs(361)));
    outputs(5180) <= layer0_outputs(1111);
    outputs(5181) <= (layer0_outputs(4230)) and not (layer0_outputs(5133));
    outputs(5182) <= not(layer0_outputs(3818));
    outputs(5183) <= not(layer0_outputs(4267));
    outputs(5184) <= layer0_outputs(5392);
    outputs(5185) <= layer0_outputs(7378);
    outputs(5186) <= not((layer0_outputs(6700)) and (layer0_outputs(5906)));
    outputs(5187) <= not((layer0_outputs(4191)) xor (layer0_outputs(3630)));
    outputs(5188) <= not((layer0_outputs(2054)) and (layer0_outputs(6926)));
    outputs(5189) <= layer0_outputs(3353);
    outputs(5190) <= (layer0_outputs(7651)) and (layer0_outputs(1594));
    outputs(5191) <= layer0_outputs(1458);
    outputs(5192) <= not(layer0_outputs(4848));
    outputs(5193) <= not(layer0_outputs(3437)) or (layer0_outputs(1836));
    outputs(5194) <= (layer0_outputs(6312)) and not (layer0_outputs(2085));
    outputs(5195) <= (layer0_outputs(3832)) xor (layer0_outputs(208));
    outputs(5196) <= layer0_outputs(7386);
    outputs(5197) <= (layer0_outputs(5766)) and not (layer0_outputs(204));
    outputs(5198) <= not(layer0_outputs(2074));
    outputs(5199) <= layer0_outputs(2514);
    outputs(5200) <= (layer0_outputs(7439)) or (layer0_outputs(4947));
    outputs(5201) <= layer0_outputs(1904);
    outputs(5202) <= not(layer0_outputs(6452)) or (layer0_outputs(3143));
    outputs(5203) <= not(layer0_outputs(5191)) or (layer0_outputs(821));
    outputs(5204) <= layer0_outputs(3463);
    outputs(5205) <= not(layer0_outputs(3683));
    outputs(5206) <= (layer0_outputs(2212)) xor (layer0_outputs(4756));
    outputs(5207) <= not(layer0_outputs(1510));
    outputs(5208) <= layer0_outputs(7539);
    outputs(5209) <= not(layer0_outputs(5888));
    outputs(5210) <= layer0_outputs(2426);
    outputs(5211) <= layer0_outputs(550);
    outputs(5212) <= layer0_outputs(4724);
    outputs(5213) <= not(layer0_outputs(7608));
    outputs(5214) <= (layer0_outputs(2500)) and (layer0_outputs(2608));
    outputs(5215) <= (layer0_outputs(5529)) xor (layer0_outputs(7419));
    outputs(5216) <= not(layer0_outputs(5308)) or (layer0_outputs(1874));
    outputs(5217) <= not(layer0_outputs(3635));
    outputs(5218) <= layer0_outputs(5349);
    outputs(5219) <= (layer0_outputs(7390)) and not (layer0_outputs(1011));
    outputs(5220) <= not((layer0_outputs(2104)) xor (layer0_outputs(1233)));
    outputs(5221) <= layer0_outputs(4058);
    outputs(5222) <= (layer0_outputs(1864)) and not (layer0_outputs(7010));
    outputs(5223) <= (layer0_outputs(5995)) and not (layer0_outputs(6441));
    outputs(5224) <= (layer0_outputs(5520)) and not (layer0_outputs(3135));
    outputs(5225) <= layer0_outputs(7586);
    outputs(5226) <= layer0_outputs(3429);
    outputs(5227) <= (layer0_outputs(419)) and (layer0_outputs(2306));
    outputs(5228) <= layer0_outputs(3260);
    outputs(5229) <= not(layer0_outputs(1989));
    outputs(5230) <= not((layer0_outputs(2007)) xor (layer0_outputs(4625)));
    outputs(5231) <= not(layer0_outputs(1598)) or (layer0_outputs(3832));
    outputs(5232) <= (layer0_outputs(6365)) and (layer0_outputs(6233));
    outputs(5233) <= not(layer0_outputs(3805));
    outputs(5234) <= (layer0_outputs(408)) xor (layer0_outputs(6542));
    outputs(5235) <= (layer0_outputs(876)) xor (layer0_outputs(5990));
    outputs(5236) <= not((layer0_outputs(6042)) and (layer0_outputs(6613)));
    outputs(5237) <= layer0_outputs(1242);
    outputs(5238) <= not(layer0_outputs(2209));
    outputs(5239) <= layer0_outputs(6494);
    outputs(5240) <= not((layer0_outputs(7208)) xor (layer0_outputs(2632)));
    outputs(5241) <= layer0_outputs(1070);
    outputs(5242) <= not(layer0_outputs(1876));
    outputs(5243) <= layer0_outputs(193);
    outputs(5244) <= not(layer0_outputs(3726));
    outputs(5245) <= (layer0_outputs(407)) and not (layer0_outputs(4630));
    outputs(5246) <= layer0_outputs(3521);
    outputs(5247) <= layer0_outputs(3220);
    outputs(5248) <= not(layer0_outputs(322));
    outputs(5249) <= not((layer0_outputs(4377)) xor (layer0_outputs(1387)));
    outputs(5250) <= not(layer0_outputs(2957));
    outputs(5251) <= layer0_outputs(7205);
    outputs(5252) <= not(layer0_outputs(4124));
    outputs(5253) <= not((layer0_outputs(2732)) xor (layer0_outputs(1156)));
    outputs(5254) <= (layer0_outputs(7013)) xor (layer0_outputs(4412));
    outputs(5255) <= (layer0_outputs(4608)) or (layer0_outputs(3006));
    outputs(5256) <= not((layer0_outputs(6204)) xor (layer0_outputs(6598)));
    outputs(5257) <= not(layer0_outputs(2814));
    outputs(5258) <= not(layer0_outputs(5291));
    outputs(5259) <= (layer0_outputs(3028)) and not (layer0_outputs(4982));
    outputs(5260) <= layer0_outputs(4862);
    outputs(5261) <= not(layer0_outputs(1013));
    outputs(5262) <= layer0_outputs(7534);
    outputs(5263) <= not(layer0_outputs(2225));
    outputs(5264) <= layer0_outputs(4595);
    outputs(5265) <= layer0_outputs(2917);
    outputs(5266) <= layer0_outputs(1734);
    outputs(5267) <= layer0_outputs(1641);
    outputs(5268) <= layer0_outputs(7068);
    outputs(5269) <= not((layer0_outputs(6)) xor (layer0_outputs(2690)));
    outputs(5270) <= (layer0_outputs(6226)) and not (layer0_outputs(5388));
    outputs(5271) <= not(layer0_outputs(101));
    outputs(5272) <= (layer0_outputs(826)) or (layer0_outputs(3702));
    outputs(5273) <= (layer0_outputs(5677)) xor (layer0_outputs(6675));
    outputs(5274) <= layer0_outputs(5701);
    outputs(5275) <= (layer0_outputs(2153)) or (layer0_outputs(1029));
    outputs(5276) <= not(layer0_outputs(3829)) or (layer0_outputs(1194));
    outputs(5277) <= not(layer0_outputs(4285));
    outputs(5278) <= (layer0_outputs(3271)) or (layer0_outputs(4342));
    outputs(5279) <= layer0_outputs(1324);
    outputs(5280) <= not((layer0_outputs(6734)) or (layer0_outputs(3671)));
    outputs(5281) <= not(layer0_outputs(4938));
    outputs(5282) <= (layer0_outputs(6719)) or (layer0_outputs(6004));
    outputs(5283) <= (layer0_outputs(1826)) xor (layer0_outputs(3539));
    outputs(5284) <= (layer0_outputs(684)) and not (layer0_outputs(2973));
    outputs(5285) <= (layer0_outputs(6058)) and not (layer0_outputs(178));
    outputs(5286) <= not(layer0_outputs(930));
    outputs(5287) <= not((layer0_outputs(6121)) or (layer0_outputs(1837)));
    outputs(5288) <= not(layer0_outputs(5264));
    outputs(5289) <= layer0_outputs(5241);
    outputs(5290) <= not(layer0_outputs(3861));
    outputs(5291) <= layer0_outputs(111);
    outputs(5292) <= not(layer0_outputs(2454));
    outputs(5293) <= (layer0_outputs(4919)) and not (layer0_outputs(551));
    outputs(5294) <= (layer0_outputs(3927)) or (layer0_outputs(1201));
    outputs(5295) <= not(layer0_outputs(5192)) or (layer0_outputs(2907));
    outputs(5296) <= not(layer0_outputs(6937)) or (layer0_outputs(2279));
    outputs(5297) <= not(layer0_outputs(6219));
    outputs(5298) <= layer0_outputs(4334);
    outputs(5299) <= not((layer0_outputs(6214)) or (layer0_outputs(743)));
    outputs(5300) <= not(layer0_outputs(7164));
    outputs(5301) <= (layer0_outputs(6864)) and (layer0_outputs(2525));
    outputs(5302) <= (layer0_outputs(5949)) and not (layer0_outputs(81));
    outputs(5303) <= (layer0_outputs(499)) or (layer0_outputs(5196));
    outputs(5304) <= (layer0_outputs(1601)) and not (layer0_outputs(3935));
    outputs(5305) <= layer0_outputs(1279);
    outputs(5306) <= layer0_outputs(571);
    outputs(5307) <= not(layer0_outputs(6022));
    outputs(5308) <= not(layer0_outputs(6699));
    outputs(5309) <= (layer0_outputs(5982)) and (layer0_outputs(5295));
    outputs(5310) <= not(layer0_outputs(3205)) or (layer0_outputs(2725));
    outputs(5311) <= layer0_outputs(4437);
    outputs(5312) <= (layer0_outputs(7154)) xor (layer0_outputs(3112));
    outputs(5313) <= not((layer0_outputs(686)) xor (layer0_outputs(6541)));
    outputs(5314) <= not((layer0_outputs(3674)) or (layer0_outputs(89)));
    outputs(5315) <= layer0_outputs(2866);
    outputs(5316) <= not(layer0_outputs(4403));
    outputs(5317) <= not((layer0_outputs(2394)) or (layer0_outputs(2582)));
    outputs(5318) <= (layer0_outputs(5100)) and (layer0_outputs(46));
    outputs(5319) <= (layer0_outputs(2511)) or (layer0_outputs(4074));
    outputs(5320) <= (layer0_outputs(4262)) and not (layer0_outputs(4095));
    outputs(5321) <= not((layer0_outputs(2971)) and (layer0_outputs(7276)));
    outputs(5322) <= not(layer0_outputs(6601)) or (layer0_outputs(4094));
    outputs(5323) <= layer0_outputs(3760);
    outputs(5324) <= not((layer0_outputs(2457)) and (layer0_outputs(221)));
    outputs(5325) <= layer0_outputs(5536);
    outputs(5326) <= layer0_outputs(1778);
    outputs(5327) <= layer0_outputs(7120);
    outputs(5328) <= (layer0_outputs(3660)) xor (layer0_outputs(3986));
    outputs(5329) <= not(layer0_outputs(6190));
    outputs(5330) <= not(layer0_outputs(7679));
    outputs(5331) <= layer0_outputs(7364);
    outputs(5332) <= not(layer0_outputs(1362));
    outputs(5333) <= layer0_outputs(2115);
    outputs(5334) <= not(layer0_outputs(4855));
    outputs(5335) <= not(layer0_outputs(6343));
    outputs(5336) <= layer0_outputs(3364);
    outputs(5337) <= not(layer0_outputs(4793));
    outputs(5338) <= not(layer0_outputs(3796));
    outputs(5339) <= layer0_outputs(4347);
    outputs(5340) <= not((layer0_outputs(2218)) or (layer0_outputs(5522)));
    outputs(5341) <= (layer0_outputs(3884)) and not (layer0_outputs(2551));
    outputs(5342) <= not(layer0_outputs(98)) or (layer0_outputs(5061));
    outputs(5343) <= not(layer0_outputs(7495)) or (layer0_outputs(314));
    outputs(5344) <= not(layer0_outputs(775));
    outputs(5345) <= not((layer0_outputs(5229)) or (layer0_outputs(4275)));
    outputs(5346) <= not((layer0_outputs(6222)) and (layer0_outputs(740)));
    outputs(5347) <= not(layer0_outputs(5687)) or (layer0_outputs(2408));
    outputs(5348) <= (layer0_outputs(1789)) and not (layer0_outputs(5911));
    outputs(5349) <= layer0_outputs(4417);
    outputs(5350) <= (layer0_outputs(1757)) and not (layer0_outputs(4959));
    outputs(5351) <= not((layer0_outputs(6265)) or (layer0_outputs(4319)));
    outputs(5352) <= (layer0_outputs(4644)) and not (layer0_outputs(4643));
    outputs(5353) <= not((layer0_outputs(7628)) xor (layer0_outputs(654)));
    outputs(5354) <= not(layer0_outputs(2635));
    outputs(5355) <= not(layer0_outputs(5179)) or (layer0_outputs(548));
    outputs(5356) <= (layer0_outputs(7659)) xor (layer0_outputs(139));
    outputs(5357) <= (layer0_outputs(5972)) and not (layer0_outputs(5369));
    outputs(5358) <= (layer0_outputs(7382)) and not (layer0_outputs(1065));
    outputs(5359) <= layer0_outputs(6676);
    outputs(5360) <= not(layer0_outputs(2667));
    outputs(5361) <= layer0_outputs(4606);
    outputs(5362) <= not((layer0_outputs(1245)) or (layer0_outputs(869)));
    outputs(5363) <= layer0_outputs(5418);
    outputs(5364) <= layer0_outputs(2569);
    outputs(5365) <= not((layer0_outputs(3114)) or (layer0_outputs(3619)));
    outputs(5366) <= layer0_outputs(4329);
    outputs(5367) <= not((layer0_outputs(1153)) or (layer0_outputs(2747)));
    outputs(5368) <= layer0_outputs(5035);
    outputs(5369) <= (layer0_outputs(2168)) and not (layer0_outputs(5471));
    outputs(5370) <= layer0_outputs(3062);
    outputs(5371) <= (layer0_outputs(4977)) and not (layer0_outputs(5757));
    outputs(5372) <= not((layer0_outputs(281)) or (layer0_outputs(343)));
    outputs(5373) <= not(layer0_outputs(3437));
    outputs(5374) <= not((layer0_outputs(4168)) xor (layer0_outputs(3440)));
    outputs(5375) <= layer0_outputs(2639);
    outputs(5376) <= not(layer0_outputs(549)) or (layer0_outputs(4777));
    outputs(5377) <= not(layer0_outputs(6884)) or (layer0_outputs(3747));
    outputs(5378) <= layer0_outputs(4835);
    outputs(5379) <= layer0_outputs(1250);
    outputs(5380) <= (layer0_outputs(974)) xor (layer0_outputs(6503));
    outputs(5381) <= (layer0_outputs(1915)) or (layer0_outputs(6355));
    outputs(5382) <= (layer0_outputs(385)) and (layer0_outputs(878));
    outputs(5383) <= layer0_outputs(2403);
    outputs(5384) <= not(layer0_outputs(787));
    outputs(5385) <= not(layer0_outputs(6273));
    outputs(5386) <= (layer0_outputs(6525)) and not (layer0_outputs(2947));
    outputs(5387) <= layer0_outputs(2941);
    outputs(5388) <= not(layer0_outputs(1793));
    outputs(5389) <= not((layer0_outputs(6823)) or (layer0_outputs(4575)));
    outputs(5390) <= not((layer0_outputs(3781)) or (layer0_outputs(7145)));
    outputs(5391) <= not((layer0_outputs(3788)) or (layer0_outputs(387)));
    outputs(5392) <= layer0_outputs(4788);
    outputs(5393) <= not(layer0_outputs(2637));
    outputs(5394) <= not((layer0_outputs(2691)) or (layer0_outputs(2417)));
    outputs(5395) <= not(layer0_outputs(941));
    outputs(5396) <= not(layer0_outputs(6073));
    outputs(5397) <= not(layer0_outputs(6852));
    outputs(5398) <= (layer0_outputs(6034)) and not (layer0_outputs(880));
    outputs(5399) <= not((layer0_outputs(5899)) or (layer0_outputs(6337)));
    outputs(5400) <= layer0_outputs(7609);
    outputs(5401) <= (layer0_outputs(6670)) and not (layer0_outputs(6232));
    outputs(5402) <= not((layer0_outputs(6880)) xor (layer0_outputs(2325)));
    outputs(5403) <= layer0_outputs(654);
    outputs(5404) <= layer0_outputs(3208);
    outputs(5405) <= layer0_outputs(7306);
    outputs(5406) <= not((layer0_outputs(2374)) or (layer0_outputs(1021)));
    outputs(5407) <= not(layer0_outputs(4390));
    outputs(5408) <= (layer0_outputs(5406)) or (layer0_outputs(7128));
    outputs(5409) <= not(layer0_outputs(195));
    outputs(5410) <= layer0_outputs(4178);
    outputs(5411) <= layer0_outputs(2652);
    outputs(5412) <= not(layer0_outputs(1289));
    outputs(5413) <= not(layer0_outputs(2168));
    outputs(5414) <= not((layer0_outputs(1255)) or (layer0_outputs(2637)));
    outputs(5415) <= not((layer0_outputs(7376)) xor (layer0_outputs(4495)));
    outputs(5416) <= layer0_outputs(3744);
    outputs(5417) <= not(layer0_outputs(4355));
    outputs(5418) <= layer0_outputs(1317);
    outputs(5419) <= not(layer0_outputs(2958));
    outputs(5420) <= not(layer0_outputs(3116));
    outputs(5421) <= (layer0_outputs(3304)) and not (layer0_outputs(651));
    outputs(5422) <= not(layer0_outputs(4967));
    outputs(5423) <= layer0_outputs(7489);
    outputs(5424) <= (layer0_outputs(4115)) and not (layer0_outputs(5562));
    outputs(5425) <= not((layer0_outputs(6805)) xor (layer0_outputs(3996)));
    outputs(5426) <= not(layer0_outputs(5223)) or (layer0_outputs(5187));
    outputs(5427) <= layer0_outputs(5879);
    outputs(5428) <= not((layer0_outputs(1969)) xor (layer0_outputs(4185)));
    outputs(5429) <= not(layer0_outputs(1605));
    outputs(5430) <= (layer0_outputs(1559)) or (layer0_outputs(4033));
    outputs(5431) <= layer0_outputs(4952);
    outputs(5432) <= layer0_outputs(5526);
    outputs(5433) <= (layer0_outputs(6714)) and not (layer0_outputs(289));
    outputs(5434) <= not(layer0_outputs(5777));
    outputs(5435) <= layer0_outputs(3023);
    outputs(5436) <= not(layer0_outputs(483));
    outputs(5437) <= (layer0_outputs(2774)) and not (layer0_outputs(6412));
    outputs(5438) <= (layer0_outputs(1354)) and not (layer0_outputs(3275));
    outputs(5439) <= layer0_outputs(3892);
    outputs(5440) <= layer0_outputs(1552);
    outputs(5441) <= not(layer0_outputs(130));
    outputs(5442) <= layer0_outputs(4143);
    outputs(5443) <= (layer0_outputs(1160)) or (layer0_outputs(1026));
    outputs(5444) <= (layer0_outputs(2988)) and not (layer0_outputs(165));
    outputs(5445) <= layer0_outputs(1619);
    outputs(5446) <= not((layer0_outputs(6998)) or (layer0_outputs(1468)));
    outputs(5447) <= (layer0_outputs(3629)) and not (layer0_outputs(4698));
    outputs(5448) <= not(layer0_outputs(5033));
    outputs(5449) <= layer0_outputs(3670);
    outputs(5450) <= not(layer0_outputs(4455));
    outputs(5451) <= (layer0_outputs(6526)) and not (layer0_outputs(5542));
    outputs(5452) <= not(layer0_outputs(1515));
    outputs(5453) <= layer0_outputs(4940);
    outputs(5454) <= (layer0_outputs(2256)) and not (layer0_outputs(5447));
    outputs(5455) <= not(layer0_outputs(4048));
    outputs(5456) <= not(layer0_outputs(6807));
    outputs(5457) <= (layer0_outputs(7193)) xor (layer0_outputs(6684));
    outputs(5458) <= (layer0_outputs(4392)) and not (layer0_outputs(5967));
    outputs(5459) <= not(layer0_outputs(5520));
    outputs(5460) <= layer0_outputs(3872);
    outputs(5461) <= layer0_outputs(662);
    outputs(5462) <= (layer0_outputs(3264)) or (layer0_outputs(4332));
    outputs(5463) <= layer0_outputs(448);
    outputs(5464) <= not(layer0_outputs(3043));
    outputs(5465) <= not(layer0_outputs(6657)) or (layer0_outputs(6241));
    outputs(5466) <= not(layer0_outputs(2679)) or (layer0_outputs(4562));
    outputs(5467) <= (layer0_outputs(1098)) and (layer0_outputs(6302));
    outputs(5468) <= not((layer0_outputs(1352)) or (layer0_outputs(1312)));
    outputs(5469) <= not((layer0_outputs(556)) and (layer0_outputs(866)));
    outputs(5470) <= (layer0_outputs(4493)) and (layer0_outputs(1639));
    outputs(5471) <= not(layer0_outputs(2812));
    outputs(5472) <= not(layer0_outputs(5010));
    outputs(5473) <= layer0_outputs(6727);
    outputs(5474) <= not(layer0_outputs(4688));
    outputs(5475) <= not(layer0_outputs(6682));
    outputs(5476) <= not(layer0_outputs(1272));
    outputs(5477) <= not(layer0_outputs(1114)) or (layer0_outputs(6065));
    outputs(5478) <= not((layer0_outputs(522)) xor (layer0_outputs(7456)));
    outputs(5479) <= not(layer0_outputs(1984));
    outputs(5480) <= (layer0_outputs(2939)) xor (layer0_outputs(6516));
    outputs(5481) <= not(layer0_outputs(1616));
    outputs(5482) <= not(layer0_outputs(5660));
    outputs(5483) <= not(layer0_outputs(2676));
    outputs(5484) <= (layer0_outputs(4989)) and not (layer0_outputs(5052));
    outputs(5485) <= layer0_outputs(7198);
    outputs(5486) <= not(layer0_outputs(3199));
    outputs(5487) <= not((layer0_outputs(3553)) or (layer0_outputs(7440)));
    outputs(5488) <= (layer0_outputs(3226)) and not (layer0_outputs(5152));
    outputs(5489) <= not(layer0_outputs(1404));
    outputs(5490) <= (layer0_outputs(6133)) xor (layer0_outputs(2932));
    outputs(5491) <= (layer0_outputs(311)) and not (layer0_outputs(1676));
    outputs(5492) <= not(layer0_outputs(5530));
    outputs(5493) <= layer0_outputs(5068);
    outputs(5494) <= layer0_outputs(5149);
    outputs(5495) <= (layer0_outputs(3592)) xor (layer0_outputs(4171));
    outputs(5496) <= not(layer0_outputs(4402));
    outputs(5497) <= (layer0_outputs(4865)) and not (layer0_outputs(6609));
    outputs(5498) <= not((layer0_outputs(3705)) or (layer0_outputs(2257)));
    outputs(5499) <= layer0_outputs(5853);
    outputs(5500) <= (layer0_outputs(1699)) and not (layer0_outputs(849));
    outputs(5501) <= not(layer0_outputs(4667));
    outputs(5502) <= (layer0_outputs(4692)) and (layer0_outputs(1271));
    outputs(5503) <= not((layer0_outputs(2450)) or (layer0_outputs(3337)));
    outputs(5504) <= (layer0_outputs(3456)) and not (layer0_outputs(3984));
    outputs(5505) <= (layer0_outputs(3958)) or (layer0_outputs(476));
    outputs(5506) <= (layer0_outputs(215)) and not (layer0_outputs(369));
    outputs(5507) <= not((layer0_outputs(7059)) xor (layer0_outputs(631)));
    outputs(5508) <= (layer0_outputs(3323)) xor (layer0_outputs(2865));
    outputs(5509) <= layer0_outputs(1530);
    outputs(5510) <= (layer0_outputs(184)) and not (layer0_outputs(4231));
    outputs(5511) <= (layer0_outputs(2856)) and not (layer0_outputs(1233));
    outputs(5512) <= (layer0_outputs(4180)) xor (layer0_outputs(3446));
    outputs(5513) <= (layer0_outputs(382)) and not (layer0_outputs(5683));
    outputs(5514) <= layer0_outputs(4211);
    outputs(5515) <= layer0_outputs(6834);
    outputs(5516) <= (layer0_outputs(4217)) and not (layer0_outputs(3552));
    outputs(5517) <= layer0_outputs(1962);
    outputs(5518) <= (layer0_outputs(4145)) and not (layer0_outputs(7310));
    outputs(5519) <= layer0_outputs(5663);
    outputs(5520) <= not(layer0_outputs(3740));
    outputs(5521) <= not(layer0_outputs(4958)) or (layer0_outputs(642));
    outputs(5522) <= layer0_outputs(5782);
    outputs(5523) <= not((layer0_outputs(7421)) xor (layer0_outputs(224)));
    outputs(5524) <= not(layer0_outputs(6756));
    outputs(5525) <= layer0_outputs(420);
    outputs(5526) <= layer0_outputs(3835);
    outputs(5527) <= (layer0_outputs(804)) and (layer0_outputs(5131));
    outputs(5528) <= not(layer0_outputs(2805));
    outputs(5529) <= (layer0_outputs(6176)) and not (layer0_outputs(4721));
    outputs(5530) <= not(layer0_outputs(5666));
    outputs(5531) <= (layer0_outputs(5342)) and (layer0_outputs(1317));
    outputs(5532) <= not(layer0_outputs(3273));
    outputs(5533) <= (layer0_outputs(2420)) xor (layer0_outputs(4396));
    outputs(5534) <= (layer0_outputs(443)) and (layer0_outputs(2568));
    outputs(5535) <= (layer0_outputs(3543)) and (layer0_outputs(1412));
    outputs(5536) <= not(layer0_outputs(6358));
    outputs(5537) <= not((layer0_outputs(5413)) and (layer0_outputs(4103)));
    outputs(5538) <= not(layer0_outputs(6028));
    outputs(5539) <= layer0_outputs(7501);
    outputs(5540) <= (layer0_outputs(6681)) and (layer0_outputs(1976));
    outputs(5541) <= not(layer0_outputs(5072)) or (layer0_outputs(7327));
    outputs(5542) <= (layer0_outputs(4014)) xor (layer0_outputs(307));
    outputs(5543) <= layer0_outputs(4);
    outputs(5544) <= layer0_outputs(2056);
    outputs(5545) <= (layer0_outputs(5576)) and not (layer0_outputs(1094));
    outputs(5546) <= (layer0_outputs(2657)) xor (layer0_outputs(902));
    outputs(5547) <= layer0_outputs(7395);
    outputs(5548) <= (layer0_outputs(5831)) or (layer0_outputs(2796));
    outputs(5549) <= not(layer0_outputs(148));
    outputs(5550) <= not(layer0_outputs(36));
    outputs(5551) <= (layer0_outputs(1830)) xor (layer0_outputs(5836));
    outputs(5552) <= not(layer0_outputs(865));
    outputs(5553) <= (layer0_outputs(4195)) and not (layer0_outputs(7473));
    outputs(5554) <= (layer0_outputs(181)) and not (layer0_outputs(3879));
    outputs(5555) <= not((layer0_outputs(122)) xor (layer0_outputs(2716)));
    outputs(5556) <= (layer0_outputs(990)) and (layer0_outputs(7295));
    outputs(5557) <= not(layer0_outputs(5606));
    outputs(5558) <= (layer0_outputs(6291)) and not (layer0_outputs(6319));
    outputs(5559) <= not(layer0_outputs(959));
    outputs(5560) <= (layer0_outputs(3297)) and (layer0_outputs(3081));
    outputs(5561) <= not((layer0_outputs(327)) or (layer0_outputs(298)));
    outputs(5562) <= (layer0_outputs(5347)) and (layer0_outputs(6865));
    outputs(5563) <= (layer0_outputs(3574)) xor (layer0_outputs(4245));
    outputs(5564) <= layer0_outputs(3989);
    outputs(5565) <= (layer0_outputs(1569)) and (layer0_outputs(1133));
    outputs(5566) <= layer0_outputs(1162);
    outputs(5567) <= not((layer0_outputs(5875)) xor (layer0_outputs(5083)));
    outputs(5568) <= not(layer0_outputs(1848));
    outputs(5569) <= layer0_outputs(6690);
    outputs(5570) <= layer0_outputs(2915);
    outputs(5571) <= (layer0_outputs(5013)) xor (layer0_outputs(1737));
    outputs(5572) <= not((layer0_outputs(4495)) xor (layer0_outputs(1897)));
    outputs(5573) <= layer0_outputs(3256);
    outputs(5574) <= (layer0_outputs(1342)) and not (layer0_outputs(6635));
    outputs(5575) <= not((layer0_outputs(4902)) or (layer0_outputs(3025)));
    outputs(5576) <= not(layer0_outputs(879));
    outputs(5577) <= layer0_outputs(4557);
    outputs(5578) <= (layer0_outputs(4623)) and (layer0_outputs(948));
    outputs(5579) <= not(layer0_outputs(6869));
    outputs(5580) <= (layer0_outputs(7060)) and (layer0_outputs(6387));
    outputs(5581) <= (layer0_outputs(2301)) and not (layer0_outputs(6399));
    outputs(5582) <= layer0_outputs(338);
    outputs(5583) <= (layer0_outputs(3631)) and not (layer0_outputs(1531));
    outputs(5584) <= (layer0_outputs(7379)) and (layer0_outputs(6897));
    outputs(5585) <= (layer0_outputs(999)) xor (layer0_outputs(6148));
    outputs(5586) <= (layer0_outputs(6921)) and not (layer0_outputs(2951));
    outputs(5587) <= not(layer0_outputs(3234));
    outputs(5588) <= layer0_outputs(5093);
    outputs(5589) <= not((layer0_outputs(7057)) xor (layer0_outputs(2124)));
    outputs(5590) <= not((layer0_outputs(1909)) or (layer0_outputs(6648)));
    outputs(5591) <= (layer0_outputs(1246)) or (layer0_outputs(6194));
    outputs(5592) <= layer0_outputs(1824);
    outputs(5593) <= not((layer0_outputs(6014)) xor (layer0_outputs(4423)));
    outputs(5594) <= not(layer0_outputs(3737));
    outputs(5595) <= not(layer0_outputs(687));
    outputs(5596) <= (layer0_outputs(7309)) and not (layer0_outputs(4512));
    outputs(5597) <= not(layer0_outputs(6428));
    outputs(5598) <= not((layer0_outputs(2960)) and (layer0_outputs(3243)));
    outputs(5599) <= not((layer0_outputs(7406)) xor (layer0_outputs(4146)));
    outputs(5600) <= (layer0_outputs(362)) or (layer0_outputs(2645));
    outputs(5601) <= not(layer0_outputs(3904));
    outputs(5602) <= layer0_outputs(159);
    outputs(5603) <= not((layer0_outputs(161)) xor (layer0_outputs(3486)));
    outputs(5604) <= (layer0_outputs(4445)) xor (layer0_outputs(1759));
    outputs(5605) <= (layer0_outputs(3159)) and not (layer0_outputs(2970));
    outputs(5606) <= (layer0_outputs(7264)) and (layer0_outputs(7670));
    outputs(5607) <= not(layer0_outputs(5283));
    outputs(5608) <= not((layer0_outputs(18)) and (layer0_outputs(4550)));
    outputs(5609) <= layer0_outputs(1361);
    outputs(5610) <= layer0_outputs(6341);
    outputs(5611) <= not(layer0_outputs(1857)) or (layer0_outputs(3409));
    outputs(5612) <= not((layer0_outputs(279)) or (layer0_outputs(6620)));
    outputs(5613) <= not(layer0_outputs(39));
    outputs(5614) <= not(layer0_outputs(2713));
    outputs(5615) <= not(layer0_outputs(1297));
    outputs(5616) <= not(layer0_outputs(2055));
    outputs(5617) <= (layer0_outputs(838)) and not (layer0_outputs(4453));
    outputs(5618) <= layer0_outputs(2655);
    outputs(5619) <= not(layer0_outputs(541));
    outputs(5620) <= (layer0_outputs(576)) xor (layer0_outputs(4810));
    outputs(5621) <= not(layer0_outputs(6884));
    outputs(5622) <= not(layer0_outputs(2344));
    outputs(5623) <= not((layer0_outputs(24)) xor (layer0_outputs(1190)));
    outputs(5624) <= (layer0_outputs(2098)) and (layer0_outputs(5517));
    outputs(5625) <= layer0_outputs(3466);
    outputs(5626) <= layer0_outputs(5232);
    outputs(5627) <= layer0_outputs(180);
    outputs(5628) <= not((layer0_outputs(2756)) or (layer0_outputs(411)));
    outputs(5629) <= (layer0_outputs(1119)) and not (layer0_outputs(3981));
    outputs(5630) <= not(layer0_outputs(6494));
    outputs(5631) <= layer0_outputs(2035);
    outputs(5632) <= (layer0_outputs(5393)) and (layer0_outputs(1049));
    outputs(5633) <= not((layer0_outputs(3733)) or (layer0_outputs(2666)));
    outputs(5634) <= layer0_outputs(7021);
    outputs(5635) <= (layer0_outputs(4102)) or (layer0_outputs(4229));
    outputs(5636) <= layer0_outputs(1937);
    outputs(5637) <= layer0_outputs(903);
    outputs(5638) <= not((layer0_outputs(4558)) xor (layer0_outputs(5071)));
    outputs(5639) <= not(layer0_outputs(5682));
    outputs(5640) <= not(layer0_outputs(5562));
    outputs(5641) <= (layer0_outputs(3134)) and (layer0_outputs(1561));
    outputs(5642) <= (layer0_outputs(4884)) or (layer0_outputs(6847));
    outputs(5643) <= layer0_outputs(5932);
    outputs(5644) <= (layer0_outputs(2930)) and (layer0_outputs(6037));
    outputs(5645) <= (layer0_outputs(2967)) and (layer0_outputs(4789));
    outputs(5646) <= not(layer0_outputs(2898));
    outputs(5647) <= layer0_outputs(568);
    outputs(5648) <= layer0_outputs(6681);
    outputs(5649) <= layer0_outputs(3274);
    outputs(5650) <= (layer0_outputs(800)) and not (layer0_outputs(4009));
    outputs(5651) <= (layer0_outputs(3233)) or (layer0_outputs(4563));
    outputs(5652) <= (layer0_outputs(3898)) or (layer0_outputs(617));
    outputs(5653) <= not(layer0_outputs(3405));
    outputs(5654) <= (layer0_outputs(857)) or (layer0_outputs(6742));
    outputs(5655) <= not(layer0_outputs(4833));
    outputs(5656) <= layer0_outputs(1115);
    outputs(5657) <= layer0_outputs(384);
    outputs(5658) <= not(layer0_outputs(6988));
    outputs(5659) <= layer0_outputs(1769);
    outputs(5660) <= layer0_outputs(7280);
    outputs(5661) <= not(layer0_outputs(6994));
    outputs(5662) <= not(layer0_outputs(694)) or (layer0_outputs(6918));
    outputs(5663) <= not((layer0_outputs(2985)) or (layer0_outputs(2505)));
    outputs(5664) <= not((layer0_outputs(6733)) xor (layer0_outputs(5028)));
    outputs(5665) <= layer0_outputs(676);
    outputs(5666) <= not((layer0_outputs(7035)) or (layer0_outputs(2982)));
    outputs(5667) <= (layer0_outputs(2013)) and (layer0_outputs(2022));
    outputs(5668) <= layer0_outputs(2548);
    outputs(5669) <= (layer0_outputs(10)) or (layer0_outputs(6677));
    outputs(5670) <= not(layer0_outputs(2450));
    outputs(5671) <= not(layer0_outputs(6299));
    outputs(5672) <= layer0_outputs(2219);
    outputs(5673) <= (layer0_outputs(5346)) and not (layer0_outputs(629));
    outputs(5674) <= not((layer0_outputs(3296)) or (layer0_outputs(1709)));
    outputs(5675) <= (layer0_outputs(763)) and not (layer0_outputs(7416));
    outputs(5676) <= (layer0_outputs(2034)) xor (layer0_outputs(1330));
    outputs(5677) <= layer0_outputs(7444);
    outputs(5678) <= (layer0_outputs(6583)) and not (layer0_outputs(5017));
    outputs(5679) <= (layer0_outputs(6974)) and not (layer0_outputs(479));
    outputs(5680) <= layer0_outputs(4665);
    outputs(5681) <= not(layer0_outputs(2033));
    outputs(5682) <= layer0_outputs(5906);
    outputs(5683) <= layer0_outputs(7617);
    outputs(5684) <= layer0_outputs(1066);
    outputs(5685) <= (layer0_outputs(718)) and (layer0_outputs(4687));
    outputs(5686) <= layer0_outputs(6715);
    outputs(5687) <= not((layer0_outputs(5289)) or (layer0_outputs(4270)));
    outputs(5688) <= (layer0_outputs(4917)) xor (layer0_outputs(5602));
    outputs(5689) <= (layer0_outputs(4646)) and (layer0_outputs(4963));
    outputs(5690) <= (layer0_outputs(3653)) and not (layer0_outputs(7024));
    outputs(5691) <= not((layer0_outputs(2889)) xor (layer0_outputs(3521)));
    outputs(5692) <= layer0_outputs(4454);
    outputs(5693) <= (layer0_outputs(858)) and not (layer0_outputs(5258));
    outputs(5694) <= not(layer0_outputs(7351));
    outputs(5695) <= (layer0_outputs(7188)) and not (layer0_outputs(3763));
    outputs(5696) <= not(layer0_outputs(3661));
    outputs(5697) <= layer0_outputs(4367);
    outputs(5698) <= not(layer0_outputs(2805));
    outputs(5699) <= layer0_outputs(3180);
    outputs(5700) <= layer0_outputs(6290);
    outputs(5701) <= layer0_outputs(2354);
    outputs(5702) <= not(layer0_outputs(6811));
    outputs(5703) <= not((layer0_outputs(1131)) or (layer0_outputs(6624)));
    outputs(5704) <= layer0_outputs(41);
    outputs(5705) <= not((layer0_outputs(1348)) or (layer0_outputs(2467)));
    outputs(5706) <= (layer0_outputs(3547)) and not (layer0_outputs(3830));
    outputs(5707) <= not(layer0_outputs(6764));
    outputs(5708) <= layer0_outputs(6927);
    outputs(5709) <= not((layer0_outputs(3893)) or (layer0_outputs(1890)));
    outputs(5710) <= not(layer0_outputs(406));
    outputs(5711) <= (layer0_outputs(2358)) and (layer0_outputs(5208));
    outputs(5712) <= layer0_outputs(5438);
    outputs(5713) <= layer0_outputs(913);
    outputs(5714) <= layer0_outputs(4992);
    outputs(5715) <= not(layer0_outputs(894));
    outputs(5716) <= not((layer0_outputs(4615)) or (layer0_outputs(5821)));
    outputs(5717) <= layer0_outputs(3749);
    outputs(5718) <= not(layer0_outputs(2188)) or (layer0_outputs(7374));
    outputs(5719) <= not(layer0_outputs(3673));
    outputs(5720) <= layer0_outputs(6985);
    outputs(5721) <= layer0_outputs(3613);
    outputs(5722) <= (layer0_outputs(4172)) and not (layer0_outputs(6804));
    outputs(5723) <= (layer0_outputs(3314)) and not (layer0_outputs(2285));
    outputs(5724) <= layer0_outputs(3049);
    outputs(5725) <= (layer0_outputs(3369)) xor (layer0_outputs(1503));
    outputs(5726) <= not(layer0_outputs(327));
    outputs(5727) <= (layer0_outputs(5186)) or (layer0_outputs(1791));
    outputs(5728) <= (layer0_outputs(4127)) or (layer0_outputs(5355));
    outputs(5729) <= not((layer0_outputs(1798)) or (layer0_outputs(1302)));
    outputs(5730) <= layer0_outputs(3023);
    outputs(5731) <= (layer0_outputs(5521)) and not (layer0_outputs(2144));
    outputs(5732) <= (layer0_outputs(905)) and (layer0_outputs(537));
    outputs(5733) <= (layer0_outputs(5763)) and not (layer0_outputs(7540));
    outputs(5734) <= layer0_outputs(6567);
    outputs(5735) <= not(layer0_outputs(6425));
    outputs(5736) <= layer0_outputs(215);
    outputs(5737) <= (layer0_outputs(6531)) or (layer0_outputs(3581));
    outputs(5738) <= not(layer0_outputs(2344));
    outputs(5739) <= not(layer0_outputs(2426));
    outputs(5740) <= not(layer0_outputs(5979));
    outputs(5741) <= not(layer0_outputs(7043));
    outputs(5742) <= layer0_outputs(295);
    outputs(5743) <= not(layer0_outputs(2191));
    outputs(5744) <= layer0_outputs(5293);
    outputs(5745) <= layer0_outputs(3144);
    outputs(5746) <= (layer0_outputs(5269)) and not (layer0_outputs(6767));
    outputs(5747) <= not(layer0_outputs(4530));
    outputs(5748) <= layer0_outputs(2108);
    outputs(5749) <= not(layer0_outputs(115));
    outputs(5750) <= (layer0_outputs(6638)) and (layer0_outputs(3421));
    outputs(5751) <= not((layer0_outputs(4902)) or (layer0_outputs(2642)));
    outputs(5752) <= layer0_outputs(7471);
    outputs(5753) <= not((layer0_outputs(847)) and (layer0_outputs(545)));
    outputs(5754) <= not(layer0_outputs(6818)) or (layer0_outputs(3226));
    outputs(5755) <= not(layer0_outputs(901));
    outputs(5756) <= layer0_outputs(3622);
    outputs(5757) <= not(layer0_outputs(7624));
    outputs(5758) <= not((layer0_outputs(3881)) and (layer0_outputs(5129)));
    outputs(5759) <= layer0_outputs(6847);
    outputs(5760) <= not(layer0_outputs(2349)) or (layer0_outputs(5359));
    outputs(5761) <= (layer0_outputs(3726)) and (layer0_outputs(4611));
    outputs(5762) <= layer0_outputs(1962);
    outputs(5763) <= (layer0_outputs(6734)) and not (layer0_outputs(5477));
    outputs(5764) <= not((layer0_outputs(6089)) and (layer0_outputs(7409)));
    outputs(5765) <= not(layer0_outputs(4868));
    outputs(5766) <= layer0_outputs(785);
    outputs(5767) <= (layer0_outputs(5881)) xor (layer0_outputs(6617));
    outputs(5768) <= (layer0_outputs(4635)) and not (layer0_outputs(3024));
    outputs(5769) <= (layer0_outputs(2043)) and not (layer0_outputs(4130));
    outputs(5770) <= layer0_outputs(2155);
    outputs(5771) <= layer0_outputs(874);
    outputs(5772) <= (layer0_outputs(2138)) or (layer0_outputs(2278));
    outputs(5773) <= layer0_outputs(4768);
    outputs(5774) <= not(layer0_outputs(5288));
    outputs(5775) <= (layer0_outputs(1156)) and not (layer0_outputs(770));
    outputs(5776) <= (layer0_outputs(5834)) xor (layer0_outputs(3438));
    outputs(5777) <= not(layer0_outputs(7205));
    outputs(5778) <= not((layer0_outputs(5511)) or (layer0_outputs(3429)));
    outputs(5779) <= not(layer0_outputs(7629));
    outputs(5780) <= not(layer0_outputs(7212));
    outputs(5781) <= not((layer0_outputs(5270)) or (layer0_outputs(110)));
    outputs(5782) <= layer0_outputs(2352);
    outputs(5783) <= (layer0_outputs(6710)) and not (layer0_outputs(4521));
    outputs(5784) <= layer0_outputs(4927);
    outputs(5785) <= not(layer0_outputs(1320));
    outputs(5786) <= not(layer0_outputs(4072));
    outputs(5787) <= not(layer0_outputs(6202));
    outputs(5788) <= not((layer0_outputs(5762)) xor (layer0_outputs(278)));
    outputs(5789) <= not(layer0_outputs(1727));
    outputs(5790) <= not((layer0_outputs(3155)) or (layer0_outputs(5795)));
    outputs(5791) <= not(layer0_outputs(7290));
    outputs(5792) <= not(layer0_outputs(4394));
    outputs(5793) <= (layer0_outputs(3247)) xor (layer0_outputs(4321));
    outputs(5794) <= layer0_outputs(3770);
    outputs(5795) <= layer0_outputs(5060);
    outputs(5796) <= layer0_outputs(3471);
    outputs(5797) <= not(layer0_outputs(1608));
    outputs(5798) <= (layer0_outputs(2942)) and (layer0_outputs(627));
    outputs(5799) <= layer0_outputs(397);
    outputs(5800) <= (layer0_outputs(1036)) and not (layer0_outputs(6096));
    outputs(5801) <= not((layer0_outputs(4045)) xor (layer0_outputs(2769)));
    outputs(5802) <= not(layer0_outputs(3289));
    outputs(5803) <= (layer0_outputs(4220)) and (layer0_outputs(1439));
    outputs(5804) <= not(layer0_outputs(3490));
    outputs(5805) <= layer0_outputs(4686);
    outputs(5806) <= not((layer0_outputs(1894)) xor (layer0_outputs(3182)));
    outputs(5807) <= not(layer0_outputs(724));
    outputs(5808) <= not(layer0_outputs(5672));
    outputs(5809) <= not(layer0_outputs(2773));
    outputs(5810) <= not((layer0_outputs(452)) or (layer0_outputs(1059)));
    outputs(5811) <= layer0_outputs(6323);
    outputs(5812) <= (layer0_outputs(2458)) and (layer0_outputs(804));
    outputs(5813) <= not((layer0_outputs(2541)) xor (layer0_outputs(2134)));
    outputs(5814) <= not(layer0_outputs(7204));
    outputs(5815) <= (layer0_outputs(4913)) and (layer0_outputs(5081));
    outputs(5816) <= layer0_outputs(4641);
    outputs(5817) <= layer0_outputs(5522);
    outputs(5818) <= not(layer0_outputs(651));
    outputs(5819) <= (layer0_outputs(7410)) and (layer0_outputs(4814));
    outputs(5820) <= not(layer0_outputs(7441)) or (layer0_outputs(4763));
    outputs(5821) <= layer0_outputs(2235);
    outputs(5822) <= (layer0_outputs(4865)) and not (layer0_outputs(2337));
    outputs(5823) <= layer0_outputs(3280);
    outputs(5824) <= not((layer0_outputs(7645)) and (layer0_outputs(5551)));
    outputs(5825) <= not(layer0_outputs(2561));
    outputs(5826) <= not((layer0_outputs(1625)) and (layer0_outputs(6070)));
    outputs(5827) <= not(layer0_outputs(6940));
    outputs(5828) <= not(layer0_outputs(195)) or (layer0_outputs(4609));
    outputs(5829) <= not(layer0_outputs(6720));
    outputs(5830) <= layer0_outputs(2127);
    outputs(5831) <= not(layer0_outputs(6366));
    outputs(5832) <= layer0_outputs(7608);
    outputs(5833) <= layer0_outputs(3961);
    outputs(5834) <= (layer0_outputs(2556)) and (layer0_outputs(4336));
    outputs(5835) <= not(layer0_outputs(5237));
    outputs(5836) <= not((layer0_outputs(157)) xor (layer0_outputs(6577)));
    outputs(5837) <= (layer0_outputs(3990)) and (layer0_outputs(7045));
    outputs(5838) <= layer0_outputs(869);
    outputs(5839) <= layer0_outputs(6478);
    outputs(5840) <= not((layer0_outputs(3076)) or (layer0_outputs(261)));
    outputs(5841) <= layer0_outputs(6836);
    outputs(5842) <= (layer0_outputs(3172)) and not (layer0_outputs(3222));
    outputs(5843) <= (layer0_outputs(208)) and not (layer0_outputs(6524));
    outputs(5844) <= layer0_outputs(3711);
    outputs(5845) <= layer0_outputs(2220);
    outputs(5846) <= layer0_outputs(7102);
    outputs(5847) <= not(layer0_outputs(3235)) or (layer0_outputs(2943));
    outputs(5848) <= not((layer0_outputs(547)) or (layer0_outputs(6217)));
    outputs(5849) <= (layer0_outputs(5692)) and not (layer0_outputs(6110));
    outputs(5850) <= not((layer0_outputs(2552)) and (layer0_outputs(6189)));
    outputs(5851) <= (layer0_outputs(2640)) and not (layer0_outputs(842));
    outputs(5852) <= (layer0_outputs(7535)) and (layer0_outputs(3093));
    outputs(5853) <= not(layer0_outputs(5472));
    outputs(5854) <= (layer0_outputs(5072)) xor (layer0_outputs(69));
    outputs(5855) <= (layer0_outputs(1550)) and not (layer0_outputs(3266));
    outputs(5856) <= (layer0_outputs(6789)) and (layer0_outputs(6468));
    outputs(5857) <= layer0_outputs(3692);
    outputs(5858) <= not((layer0_outputs(2148)) or (layer0_outputs(6339)));
    outputs(5859) <= not((layer0_outputs(5310)) or (layer0_outputs(3864)));
    outputs(5860) <= (layer0_outputs(7337)) and (layer0_outputs(6885));
    outputs(5861) <= (layer0_outputs(1459)) or (layer0_outputs(1963));
    outputs(5862) <= (layer0_outputs(7164)) and not (layer0_outputs(2242));
    outputs(5863) <= not(layer0_outputs(1199));
    outputs(5864) <= (layer0_outputs(1095)) and not (layer0_outputs(3002));
    outputs(5865) <= layer0_outputs(6109);
    outputs(5866) <= not(layer0_outputs(6481));
    outputs(5867) <= not(layer0_outputs(5506));
    outputs(5868) <= not((layer0_outputs(3167)) xor (layer0_outputs(7419)));
    outputs(5869) <= not(layer0_outputs(610)) or (layer0_outputs(5978));
    outputs(5870) <= layer0_outputs(2987);
    outputs(5871) <= layer0_outputs(4055);
    outputs(5872) <= (layer0_outputs(382)) and not (layer0_outputs(4270));
    outputs(5873) <= not((layer0_outputs(3973)) xor (layer0_outputs(2112)));
    outputs(5874) <= layer0_outputs(7016);
    outputs(5875) <= layer0_outputs(5894);
    outputs(5876) <= layer0_outputs(4408);
    outputs(5877) <= (layer0_outputs(7584)) and not (layer0_outputs(1954));
    outputs(5878) <= not(layer0_outputs(5070));
    outputs(5879) <= layer0_outputs(4489);
    outputs(5880) <= (layer0_outputs(1160)) and not (layer0_outputs(5151));
    outputs(5881) <= not((layer0_outputs(563)) or (layer0_outputs(231)));
    outputs(5882) <= (layer0_outputs(5000)) or (layer0_outputs(7027));
    outputs(5883) <= layer0_outputs(1303);
    outputs(5884) <= not((layer0_outputs(4440)) or (layer0_outputs(7329)));
    outputs(5885) <= (layer0_outputs(2111)) and not (layer0_outputs(2956));
    outputs(5886) <= layer0_outputs(3903);
    outputs(5887) <= not((layer0_outputs(2474)) xor (layer0_outputs(7149)));
    outputs(5888) <= layer0_outputs(6835);
    outputs(5889) <= not(layer0_outputs(2334));
    outputs(5890) <= not(layer0_outputs(781));
    outputs(5891) <= not((layer0_outputs(967)) or (layer0_outputs(2807)));
    outputs(5892) <= layer0_outputs(1576);
    outputs(5893) <= not(layer0_outputs(406));
    outputs(5894) <= not((layer0_outputs(4885)) or (layer0_outputs(374)));
    outputs(5895) <= not(layer0_outputs(4428));
    outputs(5896) <= not(layer0_outputs(2192)) or (layer0_outputs(6512));
    outputs(5897) <= not(layer0_outputs(4450));
    outputs(5898) <= not((layer0_outputs(5164)) xor (layer0_outputs(5055)));
    outputs(5899) <= layer0_outputs(7380);
    outputs(5900) <= not(layer0_outputs(2703));
    outputs(5901) <= (layer0_outputs(1058)) and not (layer0_outputs(2153));
    outputs(5902) <= (layer0_outputs(6535)) and (layer0_outputs(747));
    outputs(5903) <= (layer0_outputs(3867)) and (layer0_outputs(5294));
    outputs(5904) <= (layer0_outputs(6025)) xor (layer0_outputs(3207));
    outputs(5905) <= layer0_outputs(6473);
    outputs(5906) <= layer0_outputs(5026);
    outputs(5907) <= layer0_outputs(106);
    outputs(5908) <= not((layer0_outputs(2709)) or (layer0_outputs(1623)));
    outputs(5909) <= layer0_outputs(3807);
    outputs(5910) <= not((layer0_outputs(6886)) and (layer0_outputs(5474)));
    outputs(5911) <= layer0_outputs(484);
    outputs(5912) <= layer0_outputs(226);
    outputs(5913) <= not(layer0_outputs(2092)) or (layer0_outputs(4403));
    outputs(5914) <= not(layer0_outputs(1549));
    outputs(5915) <= (layer0_outputs(3349)) and not (layer0_outputs(2446));
    outputs(5916) <= not((layer0_outputs(2613)) or (layer0_outputs(2338)));
    outputs(5917) <= not(layer0_outputs(2977));
    outputs(5918) <= layer0_outputs(4235);
    outputs(5919) <= (layer0_outputs(3336)) and not (layer0_outputs(3376));
    outputs(5920) <= (layer0_outputs(4064)) and not (layer0_outputs(1711));
    outputs(5921) <= not(layer0_outputs(603));
    outputs(5922) <= (layer0_outputs(7352)) or (layer0_outputs(5831));
    outputs(5923) <= not(layer0_outputs(893));
    outputs(5924) <= (layer0_outputs(1072)) and (layer0_outputs(4203));
    outputs(5925) <= (layer0_outputs(6297)) xor (layer0_outputs(1331));
    outputs(5926) <= not((layer0_outputs(1041)) and (layer0_outputs(960)));
    outputs(5927) <= layer0_outputs(6724);
    outputs(5928) <= not(layer0_outputs(7253)) or (layer0_outputs(5060));
    outputs(5929) <= (layer0_outputs(614)) and not (layer0_outputs(4381));
    outputs(5930) <= layer0_outputs(4717);
    outputs(5931) <= not((layer0_outputs(2193)) xor (layer0_outputs(2575)));
    outputs(5932) <= (layer0_outputs(6171)) and (layer0_outputs(4728));
    outputs(5933) <= not(layer0_outputs(5997));
    outputs(5934) <= not((layer0_outputs(5391)) xor (layer0_outputs(355)));
    outputs(5935) <= (layer0_outputs(6453)) and not (layer0_outputs(2897));
    outputs(5936) <= not((layer0_outputs(1229)) or (layer0_outputs(6446)));
    outputs(5937) <= not(layer0_outputs(4250)) or (layer0_outputs(1726));
    outputs(5938) <= (layer0_outputs(2412)) and not (layer0_outputs(2840));
    outputs(5939) <= layer0_outputs(3778);
    outputs(5940) <= (layer0_outputs(2274)) and not (layer0_outputs(4808));
    outputs(5941) <= not(layer0_outputs(1802));
    outputs(5942) <= not((layer0_outputs(3786)) xor (layer0_outputs(5868)));
    outputs(5943) <= layer0_outputs(7001);
    outputs(5944) <= (layer0_outputs(5449)) and (layer0_outputs(6538));
    outputs(5945) <= (layer0_outputs(5593)) and not (layer0_outputs(6611));
    outputs(5946) <= not((layer0_outputs(5563)) xor (layer0_outputs(2072)));
    outputs(5947) <= layer0_outputs(3174);
    outputs(5948) <= layer0_outputs(136);
    outputs(5949) <= layer0_outputs(3641);
    outputs(5950) <= not(layer0_outputs(1487));
    outputs(5951) <= (layer0_outputs(3438)) and (layer0_outputs(2065));
    outputs(5952) <= (layer0_outputs(6470)) and not (layer0_outputs(5165));
    outputs(5953) <= not((layer0_outputs(1086)) and (layer0_outputs(6906)));
    outputs(5954) <= layer0_outputs(5593);
    outputs(5955) <= (layer0_outputs(5538)) and not (layer0_outputs(481));
    outputs(5956) <= not(layer0_outputs(4046));
    outputs(5957) <= (layer0_outputs(5894)) and not (layer0_outputs(6313));
    outputs(5958) <= layer0_outputs(5624);
    outputs(5959) <= (layer0_outputs(3624)) and (layer0_outputs(3154));
    outputs(5960) <= not(layer0_outputs(2130));
    outputs(5961) <= not((layer0_outputs(3983)) or (layer0_outputs(1854)));
    outputs(5962) <= not(layer0_outputs(4100));
    outputs(5963) <= (layer0_outputs(3640)) and not (layer0_outputs(4355));
    outputs(5964) <= (layer0_outputs(7337)) and (layer0_outputs(4143));
    outputs(5965) <= layer0_outputs(6646);
    outputs(5966) <= (layer0_outputs(6220)) and not (layer0_outputs(5011));
    outputs(5967) <= not(layer0_outputs(3234));
    outputs(5968) <= (layer0_outputs(908)) or (layer0_outputs(5454));
    outputs(5969) <= not(layer0_outputs(1032));
    outputs(5970) <= (layer0_outputs(2733)) and not (layer0_outputs(1217));
    outputs(5971) <= layer0_outputs(568);
    outputs(5972) <= not((layer0_outputs(1236)) xor (layer0_outputs(6379)));
    outputs(5973) <= (layer0_outputs(5550)) xor (layer0_outputs(5747));
    outputs(5974) <= not((layer0_outputs(5675)) xor (layer0_outputs(2182)));
    outputs(5975) <= not((layer0_outputs(7477)) or (layer0_outputs(628)));
    outputs(5976) <= not((layer0_outputs(1445)) or (layer0_outputs(6956)));
    outputs(5977) <= (layer0_outputs(6361)) or (layer0_outputs(3585));
    outputs(5978) <= (layer0_outputs(2987)) and not (layer0_outputs(767));
    outputs(5979) <= (layer0_outputs(3078)) and not (layer0_outputs(3430));
    outputs(5980) <= layer0_outputs(6375);
    outputs(5981) <= not(layer0_outputs(2126));
    outputs(5982) <= (layer0_outputs(1063)) and not (layer0_outputs(5869));
    outputs(5983) <= layer0_outputs(2132);
    outputs(5984) <= (layer0_outputs(1588)) and (layer0_outputs(3815));
    outputs(5985) <= (layer0_outputs(7651)) and not (layer0_outputs(6609));
    outputs(5986) <= layer0_outputs(757);
    outputs(5987) <= not((layer0_outputs(4388)) or (layer0_outputs(6169)));
    outputs(5988) <= not(layer0_outputs(4561));
    outputs(5989) <= not(layer0_outputs(7627));
    outputs(5990) <= (layer0_outputs(3444)) and not (layer0_outputs(1416));
    outputs(5991) <= layer0_outputs(2935);
    outputs(5992) <= (layer0_outputs(6142)) and (layer0_outputs(7100));
    outputs(5993) <= not(layer0_outputs(1467));
    outputs(5994) <= not(layer0_outputs(4139));
    outputs(5995) <= not(layer0_outputs(5088));
    outputs(5996) <= layer0_outputs(1042);
    outputs(5997) <= layer0_outputs(2116);
    outputs(5998) <= (layer0_outputs(2086)) and not (layer0_outputs(7458));
    outputs(5999) <= (layer0_outputs(3706)) and (layer0_outputs(4720));
    outputs(6000) <= layer0_outputs(2744);
    outputs(6001) <= not((layer0_outputs(1934)) or (layer0_outputs(533)));
    outputs(6002) <= layer0_outputs(2967);
    outputs(6003) <= (layer0_outputs(4903)) and not (layer0_outputs(6597));
    outputs(6004) <= layer0_outputs(384);
    outputs(6005) <= (layer0_outputs(4674)) and (layer0_outputs(5767));
    outputs(6006) <= layer0_outputs(696);
    outputs(6007) <= (layer0_outputs(6113)) and not (layer0_outputs(5097));
    outputs(6008) <= (layer0_outputs(3145)) xor (layer0_outputs(3761));
    outputs(6009) <= not((layer0_outputs(3217)) or (layer0_outputs(3406)));
    outputs(6010) <= not(layer0_outputs(32));
    outputs(6011) <= not(layer0_outputs(1587));
    outputs(6012) <= not((layer0_outputs(6579)) or (layer0_outputs(5352)));
    outputs(6013) <= (layer0_outputs(3860)) and (layer0_outputs(7585));
    outputs(6014) <= not(layer0_outputs(3750));
    outputs(6015) <= layer0_outputs(4239);
    outputs(6016) <= not((layer0_outputs(7601)) xor (layer0_outputs(4498)));
    outputs(6017) <= (layer0_outputs(1212)) or (layer0_outputs(6830));
    outputs(6018) <= not(layer0_outputs(5753));
    outputs(6019) <= layer0_outputs(3008);
    outputs(6020) <= not(layer0_outputs(4114));
    outputs(6021) <= not((layer0_outputs(4292)) or (layer0_outputs(5031)));
    outputs(6022) <= not((layer0_outputs(5815)) xor (layer0_outputs(2764)));
    outputs(6023) <= (layer0_outputs(435)) and (layer0_outputs(4345));
    outputs(6024) <= not(layer0_outputs(981));
    outputs(6025) <= layer0_outputs(5056);
    outputs(6026) <= not(layer0_outputs(5511));
    outputs(6027) <= (layer0_outputs(6292)) xor (layer0_outputs(6966));
    outputs(6028) <= (layer0_outputs(591)) xor (layer0_outputs(861));
    outputs(6029) <= not(layer0_outputs(7587));
    outputs(6030) <= layer0_outputs(180);
    outputs(6031) <= (layer0_outputs(6402)) and not (layer0_outputs(2656));
    outputs(6032) <= not(layer0_outputs(7104));
    outputs(6033) <= (layer0_outputs(2777)) and not (layer0_outputs(7546));
    outputs(6034) <= not(layer0_outputs(4889));
    outputs(6035) <= (layer0_outputs(5756)) and not (layer0_outputs(580));
    outputs(6036) <= layer0_outputs(2845);
    outputs(6037) <= (layer0_outputs(7175)) or (layer0_outputs(6948));
    outputs(6038) <= not((layer0_outputs(1341)) and (layer0_outputs(7619)));
    outputs(6039) <= not(layer0_outputs(5733));
    outputs(6040) <= not(layer0_outputs(6564));
    outputs(6041) <= (layer0_outputs(3858)) and (layer0_outputs(1567));
    outputs(6042) <= (layer0_outputs(5228)) and (layer0_outputs(598));
    outputs(6043) <= not(layer0_outputs(5937));
    outputs(6044) <= not(layer0_outputs(3905));
    outputs(6045) <= (layer0_outputs(1126)) and (layer0_outputs(2355));
    outputs(6046) <= not(layer0_outputs(4278));
    outputs(6047) <= layer0_outputs(5046);
    outputs(6048) <= (layer0_outputs(2923)) xor (layer0_outputs(2008));
    outputs(6049) <= (layer0_outputs(6752)) and (layer0_outputs(3794));
    outputs(6050) <= (layer0_outputs(1195)) and (layer0_outputs(2232));
    outputs(6051) <= not(layer0_outputs(5778));
    outputs(6052) <= layer0_outputs(7114);
    outputs(6053) <= not(layer0_outputs(4142)) or (layer0_outputs(6621));
    outputs(6054) <= not(layer0_outputs(6193));
    outputs(6055) <= layer0_outputs(3503);
    outputs(6056) <= (layer0_outputs(6836)) and not (layer0_outputs(5597));
    outputs(6057) <= layer0_outputs(3244);
    outputs(6058) <= (layer0_outputs(7424)) and not (layer0_outputs(7080));
    outputs(6059) <= layer0_outputs(2296);
    outputs(6060) <= not(layer0_outputs(6426));
    outputs(6061) <= (layer0_outputs(4085)) xor (layer0_outputs(5867));
    outputs(6062) <= (layer0_outputs(5144)) and not (layer0_outputs(1587));
    outputs(6063) <= not(layer0_outputs(6344));
    outputs(6064) <= not(layer0_outputs(6657));
    outputs(6065) <= not((layer0_outputs(3714)) xor (layer0_outputs(3309)));
    outputs(6066) <= layer0_outputs(6977);
    outputs(6067) <= not((layer0_outputs(3231)) or (layer0_outputs(1468)));
    outputs(6068) <= (layer0_outputs(4828)) and not (layer0_outputs(3896));
    outputs(6069) <= not(layer0_outputs(4645));
    outputs(6070) <= layer0_outputs(674);
    outputs(6071) <= layer0_outputs(1359);
    outputs(6072) <= not((layer0_outputs(516)) xor (layer0_outputs(3736)));
    outputs(6073) <= (layer0_outputs(7197)) and (layer0_outputs(3689));
    outputs(6074) <= not(layer0_outputs(1113));
    outputs(6075) <= layer0_outputs(1427);
    outputs(6076) <= not((layer0_outputs(7267)) or (layer0_outputs(723)));
    outputs(6077) <= layer0_outputs(2532);
    outputs(6078) <= (layer0_outputs(1455)) and not (layer0_outputs(6110));
    outputs(6079) <= (layer0_outputs(4668)) and (layer0_outputs(7141));
    outputs(6080) <= (layer0_outputs(3410)) and (layer0_outputs(3564));
    outputs(6081) <= (layer0_outputs(1414)) and (layer0_outputs(4726));
    outputs(6082) <= layer0_outputs(3332);
    outputs(6083) <= not(layer0_outputs(1383));
    outputs(6084) <= layer0_outputs(2045);
    outputs(6085) <= not(layer0_outputs(2962));
    outputs(6086) <= layer0_outputs(4685);
    outputs(6087) <= (layer0_outputs(7332)) and not (layer0_outputs(6384));
    outputs(6088) <= not(layer0_outputs(1397));
    outputs(6089) <= not(layer0_outputs(7635));
    outputs(6090) <= layer0_outputs(6922);
    outputs(6091) <= not((layer0_outputs(4150)) xor (layer0_outputs(3312)));
    outputs(6092) <= (layer0_outputs(2318)) and (layer0_outputs(3684));
    outputs(6093) <= (layer0_outputs(4693)) and (layer0_outputs(5144));
    outputs(6094) <= not(layer0_outputs(689));
    outputs(6095) <= not(layer0_outputs(3028));
    outputs(6096) <= (layer0_outputs(3998)) and (layer0_outputs(5829));
    outputs(6097) <= not((layer0_outputs(3020)) or (layer0_outputs(3535)));
    outputs(6098) <= layer0_outputs(662);
    outputs(6099) <= not(layer0_outputs(2812));
    outputs(6100) <= layer0_outputs(232);
    outputs(6101) <= (layer0_outputs(7485)) and (layer0_outputs(1427));
    outputs(6102) <= layer0_outputs(712);
    outputs(6103) <= not(layer0_outputs(6555));
    outputs(6104) <= not((layer0_outputs(1175)) or (layer0_outputs(5048)));
    outputs(6105) <= layer0_outputs(5586);
    outputs(6106) <= (layer0_outputs(3796)) and not (layer0_outputs(3875));
    outputs(6107) <= layer0_outputs(5391);
    outputs(6108) <= not(layer0_outputs(6006));
    outputs(6109) <= (layer0_outputs(6910)) and not (layer0_outputs(4608));
    outputs(6110) <= (layer0_outputs(2243)) and not (layer0_outputs(1613));
    outputs(6111) <= (layer0_outputs(1161)) xor (layer0_outputs(4311));
    outputs(6112) <= not(layer0_outputs(796));
    outputs(6113) <= not((layer0_outputs(6371)) xor (layer0_outputs(4573)));
    outputs(6114) <= layer0_outputs(5171);
    outputs(6115) <= (layer0_outputs(3322)) and not (layer0_outputs(6273));
    outputs(6116) <= (layer0_outputs(7218)) and (layer0_outputs(2903));
    outputs(6117) <= (layer0_outputs(7194)) and not (layer0_outputs(561));
    outputs(6118) <= layer0_outputs(637);
    outputs(6119) <= not(layer0_outputs(6182));
    outputs(6120) <= not((layer0_outputs(1167)) and (layer0_outputs(4246)));
    outputs(6121) <= layer0_outputs(7388);
    outputs(6122) <= layer0_outputs(3625);
    outputs(6123) <= not((layer0_outputs(631)) or (layer0_outputs(4253)));
    outputs(6124) <= layer0_outputs(1239);
    outputs(6125) <= not((layer0_outputs(1326)) or (layer0_outputs(3183)));
    outputs(6126) <= (layer0_outputs(7288)) and not (layer0_outputs(5910));
    outputs(6127) <= not(layer0_outputs(2613));
    outputs(6128) <= layer0_outputs(5074);
    outputs(6129) <= layer0_outputs(1899);
    outputs(6130) <= (layer0_outputs(4467)) and (layer0_outputs(5205));
    outputs(6131) <= (layer0_outputs(6945)) and not (layer0_outputs(3691));
    outputs(6132) <= not(layer0_outputs(5403));
    outputs(6133) <= layer0_outputs(762);
    outputs(6134) <= not((layer0_outputs(5823)) xor (layer0_outputs(600)));
    outputs(6135) <= (layer0_outputs(3977)) xor (layer0_outputs(6309));
    outputs(6136) <= (layer0_outputs(1614)) and not (layer0_outputs(6943));
    outputs(6137) <= (layer0_outputs(1846)) xor (layer0_outputs(4036));
    outputs(6138) <= (layer0_outputs(1377)) and not (layer0_outputs(722));
    outputs(6139) <= not((layer0_outputs(7658)) or (layer0_outputs(1891)));
    outputs(6140) <= not(layer0_outputs(5486));
    outputs(6141) <= layer0_outputs(6566);
    outputs(6142) <= layer0_outputs(5718);
    outputs(6143) <= (layer0_outputs(4234)) or (layer0_outputs(3912));
    outputs(6144) <= not(layer0_outputs(6642));
    outputs(6145) <= (layer0_outputs(77)) xor (layer0_outputs(4884));
    outputs(6146) <= not(layer0_outputs(670));
    outputs(6147) <= layer0_outputs(3960);
    outputs(6148) <= not(layer0_outputs(4086));
    outputs(6149) <= (layer0_outputs(2277)) xor (layer0_outputs(4462));
    outputs(6150) <= (layer0_outputs(2185)) xor (layer0_outputs(7607));
    outputs(6151) <= not(layer0_outputs(2693));
    outputs(6152) <= not(layer0_outputs(6037));
    outputs(6153) <= not(layer0_outputs(5238)) or (layer0_outputs(4073));
    outputs(6154) <= layer0_outputs(2);
    outputs(6155) <= not(layer0_outputs(3844));
    outputs(6156) <= (layer0_outputs(5170)) and (layer0_outputs(2127));
    outputs(6157) <= layer0_outputs(7591);
    outputs(6158) <= (layer0_outputs(7675)) and (layer0_outputs(589));
    outputs(6159) <= not(layer0_outputs(7355)) or (layer0_outputs(5170));
    outputs(6160) <= not((layer0_outputs(939)) xor (layer0_outputs(6658)));
    outputs(6161) <= layer0_outputs(2712);
    outputs(6162) <= not((layer0_outputs(2140)) xor (layer0_outputs(169)));
    outputs(6163) <= not(layer0_outputs(293));
    outputs(6164) <= not(layer0_outputs(4776));
    outputs(6165) <= not(layer0_outputs(3546)) or (layer0_outputs(7640));
    outputs(6166) <= (layer0_outputs(6500)) xor (layer0_outputs(812));
    outputs(6167) <= layer0_outputs(6166);
    outputs(6168) <= not((layer0_outputs(2282)) xor (layer0_outputs(1980)));
    outputs(6169) <= (layer0_outputs(4515)) or (layer0_outputs(5123));
    outputs(6170) <= (layer0_outputs(1141)) xor (layer0_outputs(6213));
    outputs(6171) <= not(layer0_outputs(4968)) or (layer0_outputs(1957));
    outputs(6172) <= not(layer0_outputs(4912)) or (layer0_outputs(1576));
    outputs(6173) <= not((layer0_outputs(1105)) xor (layer0_outputs(3909)));
    outputs(6174) <= layer0_outputs(6342);
    outputs(6175) <= not((layer0_outputs(1235)) or (layer0_outputs(7555)));
    outputs(6176) <= (layer0_outputs(6295)) and not (layer0_outputs(5380));
    outputs(6177) <= (layer0_outputs(5343)) and not (layer0_outputs(4483));
    outputs(6178) <= (layer0_outputs(3988)) xor (layer0_outputs(1745));
    outputs(6179) <= not(layer0_outputs(2925));
    outputs(6180) <= (layer0_outputs(2472)) xor (layer0_outputs(223));
    outputs(6181) <= layer0_outputs(3803);
    outputs(6182) <= not((layer0_outputs(83)) xor (layer0_outputs(7)));
    outputs(6183) <= layer0_outputs(3476);
    outputs(6184) <= (layer0_outputs(1389)) xor (layer0_outputs(4549));
    outputs(6185) <= layer0_outputs(4833);
    outputs(6186) <= layer0_outputs(752);
    outputs(6187) <= not((layer0_outputs(2480)) and (layer0_outputs(6560)));
    outputs(6188) <= layer0_outputs(2763);
    outputs(6189) <= (layer0_outputs(823)) xor (layer0_outputs(6957));
    outputs(6190) <= (layer0_outputs(65)) xor (layer0_outputs(7438));
    outputs(6191) <= not((layer0_outputs(6728)) xor (layer0_outputs(5417)));
    outputs(6192) <= layer0_outputs(4363);
    outputs(6193) <= layer0_outputs(529);
    outputs(6194) <= layer0_outputs(59);
    outputs(6195) <= layer0_outputs(1754);
    outputs(6196) <= (layer0_outputs(3927)) and not (layer0_outputs(2152));
    outputs(6197) <= (layer0_outputs(4990)) xor (layer0_outputs(6863));
    outputs(6198) <= not((layer0_outputs(1437)) xor (layer0_outputs(5755)));
    outputs(6199) <= not(layer0_outputs(2010)) or (layer0_outputs(1101));
    outputs(6200) <= not(layer0_outputs(4474));
    outputs(6201) <= layer0_outputs(7363);
    outputs(6202) <= '1';
    outputs(6203) <= not(layer0_outputs(3402));
    outputs(6204) <= not((layer0_outputs(5890)) xor (layer0_outputs(870)));
    outputs(6205) <= layer0_outputs(308);
    outputs(6206) <= not((layer0_outputs(2636)) xor (layer0_outputs(5445)));
    outputs(6207) <= not((layer0_outputs(377)) and (layer0_outputs(7565)));
    outputs(6208) <= not(layer0_outputs(2705));
    outputs(6209) <= not((layer0_outputs(3324)) xor (layer0_outputs(7502)));
    outputs(6210) <= not(layer0_outputs(3241)) or (layer0_outputs(3053));
    outputs(6211) <= not(layer0_outputs(2653));
    outputs(6212) <= (layer0_outputs(7670)) or (layer0_outputs(928));
    outputs(6213) <= not((layer0_outputs(3492)) xor (layer0_outputs(2818)));
    outputs(6214) <= not(layer0_outputs(1373));
    outputs(6215) <= not(layer0_outputs(5042));
    outputs(6216) <= layer0_outputs(254);
    outputs(6217) <= '1';
    outputs(6218) <= layer0_outputs(7078);
    outputs(6219) <= not((layer0_outputs(2536)) and (layer0_outputs(5408)));
    outputs(6220) <= layer0_outputs(308);
    outputs(6221) <= (layer0_outputs(4480)) xor (layer0_outputs(2477));
    outputs(6222) <= not(layer0_outputs(2351));
    outputs(6223) <= not(layer0_outputs(2089));
    outputs(6224) <= (layer0_outputs(5183)) and (layer0_outputs(3966));
    outputs(6225) <= layer0_outputs(6269);
    outputs(6226) <= (layer0_outputs(6130)) and (layer0_outputs(161));
    outputs(6227) <= not(layer0_outputs(3293));
    outputs(6228) <= (layer0_outputs(5504)) and (layer0_outputs(5905));
    outputs(6229) <= (layer0_outputs(4967)) or (layer0_outputs(1189));
    outputs(6230) <= (layer0_outputs(3218)) and not (layer0_outputs(1447));
    outputs(6231) <= not(layer0_outputs(7094));
    outputs(6232) <= layer0_outputs(1630);
    outputs(6233) <= (layer0_outputs(335)) xor (layer0_outputs(4069));
    outputs(6234) <= not(layer0_outputs(4976));
    outputs(6235) <= (layer0_outputs(5220)) and not (layer0_outputs(3780));
    outputs(6236) <= (layer0_outputs(1184)) and not (layer0_outputs(5814));
    outputs(6237) <= not(layer0_outputs(5311));
    outputs(6238) <= not((layer0_outputs(2619)) or (layer0_outputs(6205)));
    outputs(6239) <= not(layer0_outputs(368));
    outputs(6240) <= (layer0_outputs(4753)) xor (layer0_outputs(5861));
    outputs(6241) <= not(layer0_outputs(2991));
    outputs(6242) <= layer0_outputs(3157);
    outputs(6243) <= not((layer0_outputs(4602)) xor (layer0_outputs(7410)));
    outputs(6244) <= (layer0_outputs(1012)) xor (layer0_outputs(854));
    outputs(6245) <= layer0_outputs(7372);
    outputs(6246) <= not(layer0_outputs(5763)) or (layer0_outputs(1652));
    outputs(6247) <= not((layer0_outputs(6941)) and (layer0_outputs(7495)));
    outputs(6248) <= not(layer0_outputs(4820));
    outputs(6249) <= not(layer0_outputs(5826)) or (layer0_outputs(7493));
    outputs(6250) <= not((layer0_outputs(4813)) or (layer0_outputs(2687)));
    outputs(6251) <= (layer0_outputs(1077)) and not (layer0_outputs(3776));
    outputs(6252) <= layer0_outputs(1287);
    outputs(6253) <= not((layer0_outputs(3698)) xor (layer0_outputs(4020)));
    outputs(6254) <= not(layer0_outputs(2935)) or (layer0_outputs(1489));
    outputs(6255) <= not((layer0_outputs(3980)) or (layer0_outputs(2079)));
    outputs(6256) <= not((layer0_outputs(7662)) xor (layer0_outputs(2137)));
    outputs(6257) <= (layer0_outputs(3299)) and not (layer0_outputs(6873));
    outputs(6258) <= not(layer0_outputs(3800));
    outputs(6259) <= (layer0_outputs(6237)) and (layer0_outputs(5851));
    outputs(6260) <= not(layer0_outputs(3194));
    outputs(6261) <= (layer0_outputs(2773)) and not (layer0_outputs(3563));
    outputs(6262) <= layer0_outputs(4366);
    outputs(6263) <= not(layer0_outputs(4291)) or (layer0_outputs(2352));
    outputs(6264) <= (layer0_outputs(6055)) xor (layer0_outputs(5878));
    outputs(6265) <= layer0_outputs(5492);
    outputs(6266) <= not((layer0_outputs(4157)) xor (layer0_outputs(915)));
    outputs(6267) <= (layer0_outputs(7434)) and (layer0_outputs(3486));
    outputs(6268) <= layer0_outputs(2422);
    outputs(6269) <= (layer0_outputs(5276)) and not (layer0_outputs(6159));
    outputs(6270) <= (layer0_outputs(163)) or (layer0_outputs(7432));
    outputs(6271) <= (layer0_outputs(4857)) and not (layer0_outputs(4999));
    outputs(6272) <= (layer0_outputs(6529)) xor (layer0_outputs(3475));
    outputs(6273) <= not(layer0_outputs(2761));
    outputs(6274) <= not(layer0_outputs(2688)) or (layer0_outputs(3114));
    outputs(6275) <= (layer0_outputs(1885)) xor (layer0_outputs(7002));
    outputs(6276) <= layer0_outputs(1222);
    outputs(6277) <= not((layer0_outputs(6963)) and (layer0_outputs(3596)));
    outputs(6278) <= not(layer0_outputs(1955));
    outputs(6279) <= not(layer0_outputs(203)) or (layer0_outputs(3557));
    outputs(6280) <= (layer0_outputs(2293)) xor (layer0_outputs(3989));
    outputs(6281) <= layer0_outputs(5636);
    outputs(6282) <= layer0_outputs(5219);
    outputs(6283) <= not(layer0_outputs(6220));
    outputs(6284) <= layer0_outputs(2955);
    outputs(6285) <= not(layer0_outputs(4883));
    outputs(6286) <= not(layer0_outputs(7270)) or (layer0_outputs(6178));
    outputs(6287) <= layer0_outputs(3117);
    outputs(6288) <= not((layer0_outputs(2522)) xor (layer0_outputs(2156)));
    outputs(6289) <= not((layer0_outputs(5281)) and (layer0_outputs(6522)));
    outputs(6290) <= layer0_outputs(7588);
    outputs(6291) <= layer0_outputs(185);
    outputs(6292) <= not(layer0_outputs(2628)) or (layer0_outputs(6209));
    outputs(6293) <= not(layer0_outputs(2558)) or (layer0_outputs(5013));
    outputs(6294) <= layer0_outputs(7254);
    outputs(6295) <= not((layer0_outputs(3544)) and (layer0_outputs(5638)));
    outputs(6296) <= not((layer0_outputs(2811)) and (layer0_outputs(6243)));
    outputs(6297) <= layer0_outputs(5926);
    outputs(6298) <= (layer0_outputs(1495)) xor (layer0_outputs(586));
    outputs(6299) <= layer0_outputs(5752);
    outputs(6300) <= (layer0_outputs(6101)) and not (layer0_outputs(1308));
    outputs(6301) <= not(layer0_outputs(379));
    outputs(6302) <= not(layer0_outputs(2934)) or (layer0_outputs(4872));
    outputs(6303) <= not(layer0_outputs(825));
    outputs(6304) <= not((layer0_outputs(1177)) xor (layer0_outputs(6717)));
    outputs(6305) <= not((layer0_outputs(5928)) and (layer0_outputs(7151)));
    outputs(6306) <= not(layer0_outputs(3980));
    outputs(6307) <= (layer0_outputs(1759)) and not (layer0_outputs(1323));
    outputs(6308) <= not(layer0_outputs(3916));
    outputs(6309) <= layer0_outputs(2004);
    outputs(6310) <= layer0_outputs(1815);
    outputs(6311) <= not(layer0_outputs(3224)) or (layer0_outputs(5505));
    outputs(6312) <= (layer0_outputs(2177)) xor (layer0_outputs(7469));
    outputs(6313) <= not((layer0_outputs(4137)) xor (layer0_outputs(6791)));
    outputs(6314) <= not(layer0_outputs(272));
    outputs(6315) <= layer0_outputs(5038);
    outputs(6316) <= not((layer0_outputs(4468)) xor (layer0_outputs(2934)));
    outputs(6317) <= (layer0_outputs(2601)) or (layer0_outputs(244));
    outputs(6318) <= not((layer0_outputs(341)) xor (layer0_outputs(6228)));
    outputs(6319) <= not(layer0_outputs(1481)) or (layer0_outputs(3046));
    outputs(6320) <= not((layer0_outputs(1975)) xor (layer0_outputs(6857)));
    outputs(6321) <= not(layer0_outputs(5008)) or (layer0_outputs(4614));
    outputs(6322) <= not(layer0_outputs(5214));
    outputs(6323) <= (layer0_outputs(599)) xor (layer0_outputs(3822));
    outputs(6324) <= layer0_outputs(3583);
    outputs(6325) <= (layer0_outputs(4296)) or (layer0_outputs(5891));
    outputs(6326) <= not(layer0_outputs(6418));
    outputs(6327) <= layer0_outputs(4014);
    outputs(6328) <= not(layer0_outputs(706));
    outputs(6329) <= not(layer0_outputs(2798));
    outputs(6330) <= not(layer0_outputs(1906));
    outputs(6331) <= not(layer0_outputs(3597));
    outputs(6332) <= not(layer0_outputs(5053));
    outputs(6333) <= not(layer0_outputs(2303)) or (layer0_outputs(4441));
    outputs(6334) <= (layer0_outputs(205)) and not (layer0_outputs(806));
    outputs(6335) <= not((layer0_outputs(7240)) xor (layer0_outputs(6709)));
    outputs(6336) <= (layer0_outputs(437)) and not (layer0_outputs(5225));
    outputs(6337) <= not((layer0_outputs(7253)) and (layer0_outputs(1472)));
    outputs(6338) <= not((layer0_outputs(6586)) xor (layer0_outputs(3689)));
    outputs(6339) <= (layer0_outputs(4063)) and (layer0_outputs(6822));
    outputs(6340) <= layer0_outputs(2057);
    outputs(6341) <= not((layer0_outputs(6118)) xor (layer0_outputs(874)));
    outputs(6342) <= (layer0_outputs(324)) xor (layer0_outputs(4627));
    outputs(6343) <= (layer0_outputs(4397)) and not (layer0_outputs(597));
    outputs(6344) <= not((layer0_outputs(4930)) xor (layer0_outputs(319)));
    outputs(6345) <= not((layer0_outputs(939)) xor (layer0_outputs(862)));
    outputs(6346) <= not(layer0_outputs(6141));
    outputs(6347) <= not(layer0_outputs(2175)) or (layer0_outputs(4226));
    outputs(6348) <= (layer0_outputs(7363)) and not (layer0_outputs(3877));
    outputs(6349) <= not(layer0_outputs(2611));
    outputs(6350) <= layer0_outputs(4950);
    outputs(6351) <= not(layer0_outputs(6814)) or (layer0_outputs(2071));
    outputs(6352) <= (layer0_outputs(6810)) and (layer0_outputs(7434));
    outputs(6353) <= layer0_outputs(5379);
    outputs(6354) <= layer0_outputs(2470);
    outputs(6355) <= not((layer0_outputs(4207)) and (layer0_outputs(3504)));
    outputs(6356) <= (layer0_outputs(7449)) or (layer0_outputs(3153));
    outputs(6357) <= not(layer0_outputs(2081));
    outputs(6358) <= layer0_outputs(3782);
    outputs(6359) <= not(layer0_outputs(6203));
    outputs(6360) <= not((layer0_outputs(4585)) or (layer0_outputs(5549)));
    outputs(6361) <= layer0_outputs(702);
    outputs(6362) <= not((layer0_outputs(2797)) xor (layer0_outputs(5439)));
    outputs(6363) <= layer0_outputs(5629);
    outputs(6364) <= not(layer0_outputs(1634));
    outputs(6365) <= not(layer0_outputs(4595));
    outputs(6366) <= not((layer0_outputs(1288)) xor (layer0_outputs(3399)));
    outputs(6367) <= not((layer0_outputs(6640)) xor (layer0_outputs(3449)));
    outputs(6368) <= not(layer0_outputs(5587));
    outputs(6369) <= (layer0_outputs(45)) xor (layer0_outputs(1820));
    outputs(6370) <= not(layer0_outputs(5746));
    outputs(6371) <= (layer0_outputs(5738)) xor (layer0_outputs(5945));
    outputs(6372) <= not(layer0_outputs(3568));
    outputs(6373) <= (layer0_outputs(4029)) or (layer0_outputs(2655));
    outputs(6374) <= not((layer0_outputs(5565)) xor (layer0_outputs(6146)));
    outputs(6375) <= (layer0_outputs(3984)) xor (layer0_outputs(1111));
    outputs(6376) <= not(layer0_outputs(2410)) or (layer0_outputs(6359));
    outputs(6377) <= not(layer0_outputs(3325));
    outputs(6378) <= not((layer0_outputs(2363)) and (layer0_outputs(3215)));
    outputs(6379) <= not(layer0_outputs(3485));
    outputs(6380) <= (layer0_outputs(5429)) or (layer0_outputs(6987));
    outputs(6381) <= layer0_outputs(7217);
    outputs(6382) <= layer0_outputs(7666);
    outputs(6383) <= not((layer0_outputs(2699)) and (layer0_outputs(897)));
    outputs(6384) <= layer0_outputs(2395);
    outputs(6385) <= (layer0_outputs(3148)) and not (layer0_outputs(4113));
    outputs(6386) <= not(layer0_outputs(7575));
    outputs(6387) <= not(layer0_outputs(1370));
    outputs(6388) <= not(layer0_outputs(6776));
    outputs(6389) <= (layer0_outputs(5512)) and (layer0_outputs(6055));
    outputs(6390) <= layer0_outputs(5922);
    outputs(6391) <= (layer0_outputs(1366)) xor (layer0_outputs(796));
    outputs(6392) <= layer0_outputs(7641);
    outputs(6393) <= not(layer0_outputs(4693));
    outputs(6394) <= (layer0_outputs(2815)) and (layer0_outputs(2128));
    outputs(6395) <= (layer0_outputs(4868)) xor (layer0_outputs(6013));
    outputs(6396) <= (layer0_outputs(996)) xor (layer0_outputs(2159));
    outputs(6397) <= layer0_outputs(4338);
    outputs(6398) <= not((layer0_outputs(3423)) xor (layer0_outputs(2870)));
    outputs(6399) <= not(layer0_outputs(1657));
    outputs(6400) <= (layer0_outputs(2831)) xor (layer0_outputs(4818));
    outputs(6401) <= (layer0_outputs(1563)) and not (layer0_outputs(7482));
    outputs(6402) <= not((layer0_outputs(7195)) and (layer0_outputs(7143)));
    outputs(6403) <= not(layer0_outputs(3938)) or (layer0_outputs(2526));
    outputs(6404) <= (layer0_outputs(5360)) or (layer0_outputs(4540));
    outputs(6405) <= not(layer0_outputs(6172));
    outputs(6406) <= layer0_outputs(2424);
    outputs(6407) <= not(layer0_outputs(4676)) or (layer0_outputs(2107));
    outputs(6408) <= layer0_outputs(1612);
    outputs(6409) <= (layer0_outputs(2077)) and not (layer0_outputs(4916));
    outputs(6410) <= not((layer0_outputs(1749)) and (layer0_outputs(4323)));
    outputs(6411) <= layer0_outputs(6580);
    outputs(6412) <= not((layer0_outputs(2266)) and (layer0_outputs(2829)));
    outputs(6413) <= not((layer0_outputs(4120)) and (layer0_outputs(2924)));
    outputs(6414) <= (layer0_outputs(2040)) or (layer0_outputs(2171));
    outputs(6415) <= (layer0_outputs(15)) and (layer0_outputs(7132));
    outputs(6416) <= not(layer0_outputs(4503));
    outputs(6417) <= (layer0_outputs(3269)) xor (layer0_outputs(334));
    outputs(6418) <= layer0_outputs(2621);
    outputs(6419) <= not((layer0_outputs(4675)) xor (layer0_outputs(5689)));
    outputs(6420) <= (layer0_outputs(6502)) xor (layer0_outputs(7567));
    outputs(6421) <= not((layer0_outputs(2360)) and (layer0_outputs(1914)));
    outputs(6422) <= (layer0_outputs(7231)) xor (layer0_outputs(6890));
    outputs(6423) <= not(layer0_outputs(133));
    outputs(6424) <= layer0_outputs(7190);
    outputs(6425) <= not((layer0_outputs(1104)) or (layer0_outputs(4628)));
    outputs(6426) <= layer0_outputs(881);
    outputs(6427) <= not((layer0_outputs(4528)) xor (layer0_outputs(7662)));
    outputs(6428) <= not(layer0_outputs(993)) or (layer0_outputs(3183));
    outputs(6429) <= not((layer0_outputs(6815)) and (layer0_outputs(2734)));
    outputs(6430) <= layer0_outputs(6545);
    outputs(6431) <= (layer0_outputs(5419)) or (layer0_outputs(1638));
    outputs(6432) <= not(layer0_outputs(4651)) or (layer0_outputs(839));
    outputs(6433) <= not(layer0_outputs(5871));
    outputs(6434) <= layer0_outputs(3871);
    outputs(6435) <= not(layer0_outputs(1067));
    outputs(6436) <= not((layer0_outputs(7291)) and (layer0_outputs(21)));
    outputs(6437) <= not(layer0_outputs(4207)) or (layer0_outputs(3997));
    outputs(6438) <= layer0_outputs(560);
    outputs(6439) <= not(layer0_outputs(5326));
    outputs(6440) <= (layer0_outputs(4706)) and not (layer0_outputs(1663));
    outputs(6441) <= not(layer0_outputs(5584));
    outputs(6442) <= (layer0_outputs(7481)) xor (layer0_outputs(2197));
    outputs(6443) <= not(layer0_outputs(3457));
    outputs(6444) <= layer0_outputs(3733);
    outputs(6445) <= layer0_outputs(6094);
    outputs(6446) <= (layer0_outputs(260)) xor (layer0_outputs(3940));
    outputs(6447) <= layer0_outputs(7267);
    outputs(6448) <= layer0_outputs(2044);
    outputs(6449) <= not(layer0_outputs(6541));
    outputs(6450) <= not((layer0_outputs(6391)) xor (layer0_outputs(5169)));
    outputs(6451) <= not((layer0_outputs(7266)) and (layer0_outputs(6583)));
    outputs(6452) <= not((layer0_outputs(5768)) xor (layer0_outputs(3360)));
    outputs(6453) <= (layer0_outputs(6819)) xor (layer0_outputs(6156));
    outputs(6454) <= not(layer0_outputs(4587));
    outputs(6455) <= layer0_outputs(4019);
    outputs(6456) <= layer0_outputs(2886);
    outputs(6457) <= layer0_outputs(2073);
    outputs(6458) <= (layer0_outputs(688)) or (layer0_outputs(4726));
    outputs(6459) <= not(layer0_outputs(1903));
    outputs(6460) <= layer0_outputs(1849);
    outputs(6461) <= not((layer0_outputs(911)) xor (layer0_outputs(2727)));
    outputs(6462) <= not(layer0_outputs(352));
    outputs(6463) <= (layer0_outputs(5732)) and (layer0_outputs(2270));
    outputs(6464) <= not(layer0_outputs(1256));
    outputs(6465) <= (layer0_outputs(5963)) xor (layer0_outputs(2733));
    outputs(6466) <= (layer0_outputs(6360)) xor (layer0_outputs(4658));
    outputs(6467) <= layer0_outputs(1505);
    outputs(6468) <= (layer0_outputs(3493)) xor (layer0_outputs(3821));
    outputs(6469) <= not((layer0_outputs(3418)) or (layer0_outputs(6277)));
    outputs(6470) <= not((layer0_outputs(5120)) and (layer0_outputs(7667)));
    outputs(6471) <= not((layer0_outputs(1494)) xor (layer0_outputs(707)));
    outputs(6472) <= (layer0_outputs(7050)) xor (layer0_outputs(6255));
    outputs(6473) <= (layer0_outputs(6917)) and (layer0_outputs(2403));
    outputs(6474) <= (layer0_outputs(693)) xor (layer0_outputs(6440));
    outputs(6475) <= not(layer0_outputs(5848));
    outputs(6476) <= layer0_outputs(5207);
    outputs(6477) <= not(layer0_outputs(5714));
    outputs(6478) <= layer0_outputs(5914);
    outputs(6479) <= layer0_outputs(2063);
    outputs(6480) <= (layer0_outputs(4405)) xor (layer0_outputs(5884));
    outputs(6481) <= layer0_outputs(837);
    outputs(6482) <= (layer0_outputs(1764)) xor (layer0_outputs(2146));
    outputs(6483) <= not((layer0_outputs(7181)) xor (layer0_outputs(1781)));
    outputs(6484) <= layer0_outputs(3852);
    outputs(6485) <= layer0_outputs(6931);
    outputs(6486) <= not((layer0_outputs(1660)) xor (layer0_outputs(7676)));
    outputs(6487) <= (layer0_outputs(1615)) or (layer0_outputs(5285));
    outputs(6488) <= layer0_outputs(969);
    outputs(6489) <= not(layer0_outputs(1274));
    outputs(6490) <= (layer0_outputs(4548)) and not (layer0_outputs(6784));
    outputs(6491) <= not((layer0_outputs(5224)) xor (layer0_outputs(544)));
    outputs(6492) <= not(layer0_outputs(5312));
    outputs(6493) <= not(layer0_outputs(3936));
    outputs(6494) <= layer0_outputs(5835);
    outputs(6495) <= layer0_outputs(2660);
    outputs(6496) <= (layer0_outputs(16)) or (layer0_outputs(3068));
    outputs(6497) <= not((layer0_outputs(3483)) and (layer0_outputs(1537)));
    outputs(6498) <= (layer0_outputs(6149)) and not (layer0_outputs(1772));
    outputs(6499) <= layer0_outputs(3843);
    outputs(6500) <= not(layer0_outputs(7388));
    outputs(6501) <= (layer0_outputs(468)) xor (layer0_outputs(6656));
    outputs(6502) <= not(layer0_outputs(6384)) or (layer0_outputs(530));
    outputs(6503) <= (layer0_outputs(1929)) xor (layer0_outputs(7399));
    outputs(6504) <= layer0_outputs(7524);
    outputs(6505) <= not(layer0_outputs(2028));
    outputs(6506) <= not(layer0_outputs(4129));
    outputs(6507) <= not((layer0_outputs(5001)) and (layer0_outputs(7349)));
    outputs(6508) <= not((layer0_outputs(182)) and (layer0_outputs(2370)));
    outputs(6509) <= (layer0_outputs(36)) xor (layer0_outputs(6340));
    outputs(6510) <= not((layer0_outputs(5252)) or (layer0_outputs(3380)));
    outputs(6511) <= layer0_outputs(7462);
    outputs(6512) <= (layer0_outputs(5496)) and not (layer0_outputs(2340));
    outputs(6513) <= (layer0_outputs(2298)) xor (layer0_outputs(847));
    outputs(6514) <= layer0_outputs(441);
    outputs(6515) <= not((layer0_outputs(3092)) and (layer0_outputs(6604)));
    outputs(6516) <= (layer0_outputs(613)) xor (layer0_outputs(5940));
    outputs(6517) <= layer0_outputs(6730);
    outputs(6518) <= not((layer0_outputs(7318)) or (layer0_outputs(2097)));
    outputs(6519) <= layer0_outputs(4230);
    outputs(6520) <= (layer0_outputs(227)) and not (layer0_outputs(3230));
    outputs(6521) <= (layer0_outputs(7647)) or (layer0_outputs(409));
    outputs(6522) <= not((layer0_outputs(4135)) xor (layer0_outputs(1042)));
    outputs(6523) <= not(layer0_outputs(5628));
    outputs(6524) <= (layer0_outputs(2063)) xor (layer0_outputs(7479));
    outputs(6525) <= not(layer0_outputs(6403)) or (layer0_outputs(4991));
    outputs(6526) <= not((layer0_outputs(2246)) xor (layer0_outputs(1202)));
    outputs(6527) <= not((layer0_outputs(7230)) xor (layer0_outputs(2206)));
    outputs(6528) <= (layer0_outputs(6019)) xor (layer0_outputs(459));
    outputs(6529) <= not(layer0_outputs(754)) or (layer0_outputs(5601));
    outputs(6530) <= not((layer0_outputs(1911)) xor (layer0_outputs(888)));
    outputs(6531) <= not(layer0_outputs(4486));
    outputs(6532) <= (layer0_outputs(5740)) xor (layer0_outputs(860));
    outputs(6533) <= not((layer0_outputs(991)) and (layer0_outputs(4838)));
    outputs(6534) <= not(layer0_outputs(1700));
    outputs(6535) <= not(layer0_outputs(4018)) or (layer0_outputs(7252));
    outputs(6536) <= layer0_outputs(2813);
    outputs(6537) <= not((layer0_outputs(4085)) and (layer0_outputs(7671)));
    outputs(6538) <= (layer0_outputs(1157)) and not (layer0_outputs(4568));
    outputs(6539) <= layer0_outputs(2039);
    outputs(6540) <= not(layer0_outputs(5416)) or (layer0_outputs(3898));
    outputs(6541) <= not(layer0_outputs(5212)) or (layer0_outputs(4202));
    outputs(6542) <= layer0_outputs(4172);
    outputs(6543) <= (layer0_outputs(2178)) and not (layer0_outputs(903));
    outputs(6544) <= not(layer0_outputs(3906)) or (layer0_outputs(1922));
    outputs(6545) <= not(layer0_outputs(4140));
    outputs(6546) <= (layer0_outputs(2535)) xor (layer0_outputs(4928));
    outputs(6547) <= not(layer0_outputs(753));
    outputs(6548) <= not(layer0_outputs(5426));
    outputs(6549) <= layer0_outputs(6655);
    outputs(6550) <= (layer0_outputs(5950)) and (layer0_outputs(2050));
    outputs(6551) <= not((layer0_outputs(4760)) and (layer0_outputs(6841)));
    outputs(6552) <= not(layer0_outputs(5431));
    outputs(6553) <= (layer0_outputs(1227)) and (layer0_outputs(3591));
    outputs(6554) <= not((layer0_outputs(5483)) xor (layer0_outputs(4938)));
    outputs(6555) <= (layer0_outputs(3525)) or (layer0_outputs(6206));
    outputs(6556) <= layer0_outputs(6261);
    outputs(6557) <= not((layer0_outputs(2067)) xor (layer0_outputs(6192)));
    outputs(6558) <= layer0_outputs(7392);
    outputs(6559) <= layer0_outputs(7420);
    outputs(6560) <= layer0_outputs(132);
    outputs(6561) <= (layer0_outputs(6686)) xor (layer0_outputs(2115));
    outputs(6562) <= layer0_outputs(2302);
    outputs(6563) <= (layer0_outputs(3061)) and not (layer0_outputs(4219));
    outputs(6564) <= (layer0_outputs(6682)) and not (layer0_outputs(5404));
    outputs(6565) <= not(layer0_outputs(2015)) or (layer0_outputs(6119));
    outputs(6566) <= not(layer0_outputs(6372));
    outputs(6567) <= (layer0_outputs(4228)) xor (layer0_outputs(6093));
    outputs(6568) <= (layer0_outputs(4821)) or (layer0_outputs(7472));
    outputs(6569) <= layer0_outputs(7549);
    outputs(6570) <= (layer0_outputs(5697)) xor (layer0_outputs(3124));
    outputs(6571) <= not((layer0_outputs(3209)) and (layer0_outputs(591)));
    outputs(6572) <= layer0_outputs(6624);
    outputs(6573) <= layer0_outputs(5137);
    outputs(6574) <= not(layer0_outputs(4978)) or (layer0_outputs(4764));
    outputs(6575) <= not(layer0_outputs(461)) or (layer0_outputs(1536));
    outputs(6576) <= layer0_outputs(1513);
    outputs(6577) <= not(layer0_outputs(7539)) or (layer0_outputs(4528));
    outputs(6578) <= not(layer0_outputs(2487));
    outputs(6579) <= layer0_outputs(994);
    outputs(6580) <= (layer0_outputs(2128)) and not (layer0_outputs(7316));
    outputs(6581) <= not((layer0_outputs(1909)) and (layer0_outputs(7628)));
    outputs(6582) <= (layer0_outputs(3245)) and not (layer0_outputs(4587));
    outputs(6583) <= layer0_outputs(3769);
    outputs(6584) <= layer0_outputs(1023);
    outputs(6585) <= not(layer0_outputs(6077));
    outputs(6586) <= not(layer0_outputs(444));
    outputs(6587) <= not(layer0_outputs(4701)) or (layer0_outputs(2959));
    outputs(6588) <= (layer0_outputs(294)) or (layer0_outputs(4029));
    outputs(6589) <= not(layer0_outputs(7563)) or (layer0_outputs(916));
    outputs(6590) <= not((layer0_outputs(2753)) xor (layer0_outputs(410)));
    outputs(6591) <= not((layer0_outputs(5503)) xor (layer0_outputs(6233)));
    outputs(6592) <= not(layer0_outputs(7644));
    outputs(6593) <= not((layer0_outputs(7140)) xor (layer0_outputs(3170)));
    outputs(6594) <= not(layer0_outputs(4949));
    outputs(6595) <= not(layer0_outputs(7480)) or (layer0_outputs(1520));
    outputs(6596) <= (layer0_outputs(7455)) xor (layer0_outputs(6486));
    outputs(6597) <= not(layer0_outputs(2583));
    outputs(6598) <= layer0_outputs(2737);
    outputs(6599) <= (layer0_outputs(7323)) or (layer0_outputs(2809));
    outputs(6600) <= (layer0_outputs(6346)) xor (layer0_outputs(6416));
    outputs(6601) <= layer0_outputs(1469);
    outputs(6602) <= (layer0_outputs(7478)) and not (layer0_outputs(3625));
    outputs(6603) <= (layer0_outputs(4562)) or (layer0_outputs(6195));
    outputs(6604) <= not(layer0_outputs(3649));
    outputs(6605) <= (layer0_outputs(4582)) xor (layer0_outputs(4325));
    outputs(6606) <= layer0_outputs(576);
    outputs(6607) <= layer0_outputs(4768);
    outputs(6608) <= not((layer0_outputs(779)) and (layer0_outputs(435)));
    outputs(6609) <= not((layer0_outputs(4696)) or (layer0_outputs(1051)));
    outputs(6610) <= not((layer0_outputs(5279)) and (layer0_outputs(2300)));
    outputs(6611) <= layer0_outputs(5633);
    outputs(6612) <= not(layer0_outputs(3495)) or (layer0_outputs(4187));
    outputs(6613) <= layer0_outputs(4023);
    outputs(6614) <= (layer0_outputs(1688)) and (layer0_outputs(1732));
    outputs(6615) <= layer0_outputs(6854);
    outputs(6616) <= layer0_outputs(3355);
    outputs(6617) <= (layer0_outputs(5234)) xor (layer0_outputs(2011));
    outputs(6618) <= layer0_outputs(6610);
    outputs(6619) <= not(layer0_outputs(5917));
    outputs(6620) <= not(layer0_outputs(2939)) or (layer0_outputs(1849));
    outputs(6621) <= (layer0_outputs(7378)) xor (layer0_outputs(6260));
    outputs(6622) <= not((layer0_outputs(5951)) xor (layer0_outputs(4133)));
    outputs(6623) <= layer0_outputs(5160);
    outputs(6624) <= layer0_outputs(6349);
    outputs(6625) <= (layer0_outputs(4017)) xor (layer0_outputs(6850));
    outputs(6626) <= not(layer0_outputs(1942));
    outputs(6627) <= (layer0_outputs(3645)) and not (layer0_outputs(5305));
    outputs(6628) <= (layer0_outputs(750)) and (layer0_outputs(1673));
    outputs(6629) <= layer0_outputs(1024);
    outputs(6630) <= (layer0_outputs(1270)) and not (layer0_outputs(964));
    outputs(6631) <= (layer0_outputs(4930)) xor (layer0_outputs(1602));
    outputs(6632) <= not(layer0_outputs(5690));
    outputs(6633) <= layer0_outputs(5379);
    outputs(6634) <= (layer0_outputs(3693)) and not (layer0_outputs(4305));
    outputs(6635) <= layer0_outputs(7098);
    outputs(6636) <= not(layer0_outputs(4750));
    outputs(6637) <= layer0_outputs(4388);
    outputs(6638) <= not(layer0_outputs(6433));
    outputs(6639) <= not(layer0_outputs(6072)) or (layer0_outputs(7277));
    outputs(6640) <= layer0_outputs(3383);
    outputs(6641) <= not((layer0_outputs(7483)) xor (layer0_outputs(1652)));
    outputs(6642) <= (layer0_outputs(3667)) xor (layer0_outputs(67));
    outputs(6643) <= not(layer0_outputs(5581)) or (layer0_outputs(7596));
    outputs(6644) <= layer0_outputs(966);
    outputs(6645) <= layer0_outputs(3684);
    outputs(6646) <= (layer0_outputs(4779)) xor (layer0_outputs(4022));
    outputs(6647) <= not((layer0_outputs(6021)) xor (layer0_outputs(5982)));
    outputs(6648) <= layer0_outputs(1021);
    outputs(6649) <= (layer0_outputs(3176)) and not (layer0_outputs(4129));
    outputs(6650) <= layer0_outputs(5306);
    outputs(6651) <= layer0_outputs(1030);
    outputs(6652) <= (layer0_outputs(4509)) xor (layer0_outputs(2765));
    outputs(6653) <= not(layer0_outputs(511)) or (layer0_outputs(7536));
    outputs(6654) <= not(layer0_outputs(1391));
    outputs(6655) <= not(layer0_outputs(7622));
    outputs(6656) <= not(layer0_outputs(4922));
    outputs(6657) <= not(layer0_outputs(5325));
    outputs(6658) <= layer0_outputs(4713);
    outputs(6659) <= (layer0_outputs(2007)) or (layer0_outputs(1175));
    outputs(6660) <= not(layer0_outputs(663));
    outputs(6661) <= layer0_outputs(148);
    outputs(6662) <= (layer0_outputs(4955)) or (layer0_outputs(7423));
    outputs(6663) <= layer0_outputs(6582);
    outputs(6664) <= (layer0_outputs(925)) and (layer0_outputs(927));
    outputs(6665) <= not(layer0_outputs(2804));
    outputs(6666) <= layer0_outputs(4201);
    outputs(6667) <= (layer0_outputs(471)) and (layer0_outputs(6280));
    outputs(6668) <= layer0_outputs(5834);
    outputs(6669) <= not((layer0_outputs(46)) and (layer0_outputs(2012)));
    outputs(6670) <= not(layer0_outputs(926)) or (layer0_outputs(5254));
    outputs(6671) <= not((layer0_outputs(4935)) xor (layer0_outputs(3027)));
    outputs(6672) <= not(layer0_outputs(749)) or (layer0_outputs(7633));
    outputs(6673) <= layer0_outputs(2404);
    outputs(6674) <= not(layer0_outputs(832)) or (layer0_outputs(1491));
    outputs(6675) <= not(layer0_outputs(6185)) or (layer0_outputs(5889));
    outputs(6676) <= not((layer0_outputs(5517)) xor (layer0_outputs(1881)));
    outputs(6677) <= not(layer0_outputs(3052));
    outputs(6678) <= layer0_outputs(6140);
    outputs(6679) <= layer0_outputs(240);
    outputs(6680) <= (layer0_outputs(5632)) and not (layer0_outputs(4458));
    outputs(6681) <= (layer0_outputs(6255)) and not (layer0_outputs(1445));
    outputs(6682) <= not(layer0_outputs(2012)) or (layer0_outputs(566));
    outputs(6683) <= layer0_outputs(3965);
    outputs(6684) <= (layer0_outputs(2323)) or (layer0_outputs(1673));
    outputs(6685) <= not((layer0_outputs(2058)) xor (layer0_outputs(2815)));
    outputs(6686) <= not((layer0_outputs(731)) or (layer0_outputs(5180)));
    outputs(6687) <= (layer0_outputs(5901)) xor (layer0_outputs(87));
    outputs(6688) <= not(layer0_outputs(2766)) or (layer0_outputs(1003));
    outputs(6689) <= not(layer0_outputs(4126));
    outputs(6690) <= layer0_outputs(2883);
    outputs(6691) <= layer0_outputs(607);
    outputs(6692) <= layer0_outputs(5863);
    outputs(6693) <= not(layer0_outputs(7634));
    outputs(6694) <= not(layer0_outputs(6373)) or (layer0_outputs(5892));
    outputs(6695) <= layer0_outputs(5377);
    outputs(6696) <= not((layer0_outputs(6690)) or (layer0_outputs(1883)));
    outputs(6697) <= layer0_outputs(4173);
    outputs(6698) <= layer0_outputs(7319);
    outputs(6699) <= layer0_outputs(6929);
    outputs(6700) <= (layer0_outputs(4419)) xor (layer0_outputs(3732));
    outputs(6701) <= not(layer0_outputs(2333)) or (layer0_outputs(2523));
    outputs(6702) <= not(layer0_outputs(7639));
    outputs(6703) <= not(layer0_outputs(1332));
    outputs(6704) <= not(layer0_outputs(7100));
    outputs(6705) <= layer0_outputs(6223);
    outputs(6706) <= (layer0_outputs(4519)) and not (layer0_outputs(4259));
    outputs(6707) <= layer0_outputs(1536);
    outputs(6708) <= not(layer0_outputs(2862));
    outputs(6709) <= (layer0_outputs(6396)) and not (layer0_outputs(7103));
    outputs(6710) <= (layer0_outputs(266)) xor (layer0_outputs(6726));
    outputs(6711) <= not((layer0_outputs(5199)) xor (layer0_outputs(1154)));
    outputs(6712) <= layer0_outputs(4636);
    outputs(6713) <= (layer0_outputs(4438)) xor (layer0_outputs(4273));
    outputs(6714) <= layer0_outputs(970);
    outputs(6715) <= not(layer0_outputs(5610));
    outputs(6716) <= not((layer0_outputs(2634)) xor (layer0_outputs(1084)));
    outputs(6717) <= not(layer0_outputs(7437));
    outputs(6718) <= layer0_outputs(1080);
    outputs(6719) <= not((layer0_outputs(7226)) xor (layer0_outputs(57)));
    outputs(6720) <= (layer0_outputs(1448)) or (layer0_outputs(6972));
    outputs(6721) <= not((layer0_outputs(4263)) xor (layer0_outputs(1675)));
    outputs(6722) <= (layer0_outputs(3647)) and not (layer0_outputs(374));
    outputs(6723) <= not(layer0_outputs(6108)) or (layer0_outputs(2514));
    outputs(6724) <= (layer0_outputs(2319)) xor (layer0_outputs(1871));
    outputs(6725) <= layer0_outputs(1630);
    outputs(6726) <= not(layer0_outputs(6327));
    outputs(6727) <= layer0_outputs(3634);
    outputs(6728) <= not(layer0_outputs(5626));
    outputs(6729) <= not((layer0_outputs(7344)) xor (layer0_outputs(1073)));
    outputs(6730) <= not((layer0_outputs(3049)) xor (layer0_outputs(4318)));
    outputs(6731) <= not(layer0_outputs(6623)) or (layer0_outputs(3327));
    outputs(6732) <= not(layer0_outputs(7039));
    outputs(6733) <= not((layer0_outputs(3974)) and (layer0_outputs(5319)));
    outputs(6734) <= layer0_outputs(2135);
    outputs(6735) <= (layer0_outputs(5235)) or (layer0_outputs(3162));
    outputs(6736) <= not(layer0_outputs(1339));
    outputs(6737) <= not(layer0_outputs(1522)) or (layer0_outputs(3617));
    outputs(6738) <= not(layer0_outputs(6522));
    outputs(6739) <= (layer0_outputs(6796)) or (layer0_outputs(6301));
    outputs(6740) <= not(layer0_outputs(6867));
    outputs(6741) <= not(layer0_outputs(691));
    outputs(6742) <= (layer0_outputs(754)) xor (layer0_outputs(2336));
    outputs(6743) <= not(layer0_outputs(6542));
    outputs(6744) <= not(layer0_outputs(5745)) or (layer0_outputs(4688));
    outputs(6745) <= layer0_outputs(4294);
    outputs(6746) <= layer0_outputs(3100);
    outputs(6747) <= not(layer0_outputs(1002));
    outputs(6748) <= (layer0_outputs(2305)) xor (layer0_outputs(6732));
    outputs(6749) <= layer0_outputs(1933);
    outputs(6750) <= not((layer0_outputs(234)) xor (layer0_outputs(6760)));
    outputs(6751) <= not(layer0_outputs(4784));
    outputs(6752) <= not(layer0_outputs(6544));
    outputs(6753) <= not((layer0_outputs(4518)) xor (layer0_outputs(1098)));
    outputs(6754) <= not((layer0_outputs(1151)) or (layer0_outputs(4506)));
    outputs(6755) <= layer0_outputs(2758);
    outputs(6756) <= not((layer0_outputs(5307)) xor (layer0_outputs(7421)));
    outputs(6757) <= layer0_outputs(5029);
    outputs(6758) <= layer0_outputs(6543);
    outputs(6759) <= (layer0_outputs(123)) xor (layer0_outputs(332));
    outputs(6760) <= not(layer0_outputs(1032)) or (layer0_outputs(1033));
    outputs(6761) <= not(layer0_outputs(3015));
    outputs(6762) <= (layer0_outputs(5740)) xor (layer0_outputs(3907));
    outputs(6763) <= not((layer0_outputs(5397)) or (layer0_outputs(2052)));
    outputs(6764) <= not((layer0_outputs(6267)) or (layer0_outputs(6984)));
    outputs(6765) <= layer0_outputs(5278);
    outputs(6766) <= not(layer0_outputs(735));
    outputs(6767) <= not(layer0_outputs(12)) or (layer0_outputs(4048));
    outputs(6768) <= (layer0_outputs(2717)) xor (layer0_outputs(7320));
    outputs(6769) <= (layer0_outputs(3637)) and not (layer0_outputs(2035));
    outputs(6770) <= (layer0_outputs(5505)) and not (layer0_outputs(7470));
    outputs(6771) <= not(layer0_outputs(5659));
    outputs(6772) <= layer0_outputs(404);
    outputs(6773) <= not(layer0_outputs(2964));
    outputs(6774) <= not(layer0_outputs(25));
    outputs(6775) <= layer0_outputs(5082);
    outputs(6776) <= not(layer0_outputs(5782));
    outputs(6777) <= (layer0_outputs(7458)) xor (layer0_outputs(5604));
    outputs(6778) <= not(layer0_outputs(7000));
    outputs(6779) <= not(layer0_outputs(5545)) or (layer0_outputs(2873));
    outputs(6780) <= layer0_outputs(3559);
    outputs(6781) <= not((layer0_outputs(1712)) and (layer0_outputs(4984)));
    outputs(6782) <= (layer0_outputs(4167)) xor (layer0_outputs(5583));
    outputs(6783) <= not((layer0_outputs(930)) and (layer0_outputs(1934)));
    outputs(6784) <= not(layer0_outputs(2788)) or (layer0_outputs(4734));
    outputs(6785) <= not((layer0_outputs(7081)) xor (layer0_outputs(6463)));
    outputs(6786) <= not((layer0_outputs(2350)) xor (layer0_outputs(5446)));
    outputs(6787) <= not((layer0_outputs(3808)) xor (layer0_outputs(394)));
    outputs(6788) <= layer0_outputs(2599);
    outputs(6789) <= not((layer0_outputs(7661)) xor (layer0_outputs(7673)));
    outputs(6790) <= not((layer0_outputs(3955)) xor (layer0_outputs(7237)));
    outputs(6791) <= (layer0_outputs(4764)) or (layer0_outputs(6034));
    outputs(6792) <= layer0_outputs(2489);
    outputs(6793) <= not(layer0_outputs(3502)) or (layer0_outputs(3804));
    outputs(6794) <= (layer0_outputs(2704)) xor (layer0_outputs(764));
    outputs(6795) <= (layer0_outputs(6227)) xor (layer0_outputs(6422));
    outputs(6796) <= (layer0_outputs(5556)) or (layer0_outputs(3705));
    outputs(6797) <= layer0_outputs(2372);
    outputs(6798) <= (layer0_outputs(5685)) xor (layer0_outputs(3102));
    outputs(6799) <= layer0_outputs(6436);
    outputs(6800) <= not(layer0_outputs(1738));
    outputs(6801) <= layer0_outputs(5033);
    outputs(6802) <= layer0_outputs(1891);
    outputs(6803) <= layer0_outputs(7212);
    outputs(6804) <= not(layer0_outputs(3994));
    outputs(6805) <= not(layer0_outputs(3725));
    outputs(6806) <= not(layer0_outputs(957));
    outputs(6807) <= not(layer0_outputs(381));
    outputs(6808) <= not(layer0_outputs(2440));
    outputs(6809) <= not(layer0_outputs(6920));
    outputs(6810) <= not((layer0_outputs(4654)) xor (layer0_outputs(3110)));
    outputs(6811) <= not(layer0_outputs(3862));
    outputs(6812) <= layer0_outputs(5360);
    outputs(6813) <= (layer0_outputs(3662)) xor (layer0_outputs(3575));
    outputs(6814) <= not((layer0_outputs(6353)) and (layer0_outputs(1609)));
    outputs(6815) <= layer0_outputs(3526);
    outputs(6816) <= (layer0_outputs(4669)) xor (layer0_outputs(7003));
    outputs(6817) <= not(layer0_outputs(4703));
    outputs(6818) <= layer0_outputs(424);
    outputs(6819) <= not(layer0_outputs(5096));
    outputs(6820) <= not(layer0_outputs(2113)) or (layer0_outputs(5898));
    outputs(6821) <= layer0_outputs(5681);
    outputs(6822) <= (layer0_outputs(1129)) xor (layer0_outputs(2237));
    outputs(6823) <= layer0_outputs(3481);
    outputs(6824) <= not(layer0_outputs(3058));
    outputs(6825) <= not(layer0_outputs(7650));
    outputs(6826) <= (layer0_outputs(6946)) and not (layer0_outputs(7020));
    outputs(6827) <= (layer0_outputs(7288)) or (layer0_outputs(1699));
    outputs(6828) <= layer0_outputs(1343);
    outputs(6829) <= (layer0_outputs(6103)) and not (layer0_outputs(463));
    outputs(6830) <= not((layer0_outputs(4167)) xor (layer0_outputs(5930)));
    outputs(6831) <= (layer0_outputs(243)) and not (layer0_outputs(3363));
    outputs(6832) <= layer0_outputs(2060);
    outputs(6833) <= layer0_outputs(186);
    outputs(6834) <= layer0_outputs(6552);
    outputs(6835) <= not((layer0_outputs(7261)) or (layer0_outputs(7007)));
    outputs(6836) <= not(layer0_outputs(6151));
    outputs(6837) <= (layer0_outputs(1002)) xor (layer0_outputs(4178));
    outputs(6838) <= not(layer0_outputs(1810));
    outputs(6839) <= not(layer0_outputs(3933)) or (layer0_outputs(1479));
    outputs(6840) <= not((layer0_outputs(4234)) or (layer0_outputs(150)));
    outputs(6841) <= layer0_outputs(5856);
    outputs(6842) <= layer0_outputs(4264);
    outputs(6843) <= layer0_outputs(3602);
    outputs(6844) <= not((layer0_outputs(5810)) xor (layer0_outputs(715)));
    outputs(6845) <= layer0_outputs(4434);
    outputs(6846) <= not((layer0_outputs(4624)) and (layer0_outputs(6827)));
    outputs(6847) <= not((layer0_outputs(1599)) xor (layer0_outputs(4963)));
    outputs(6848) <= not((layer0_outputs(944)) xor (layer0_outputs(6238)));
    outputs(6849) <= not(layer0_outputs(6667));
    outputs(6850) <= (layer0_outputs(4457)) xor (layer0_outputs(3798));
    outputs(6851) <= (layer0_outputs(1243)) and (layer0_outputs(2212));
    outputs(6852) <= not((layer0_outputs(3584)) or (layer0_outputs(4763)));
    outputs(6853) <= (layer0_outputs(3163)) and not (layer0_outputs(846));
    outputs(6854) <= layer0_outputs(6854);
    outputs(6855) <= not(layer0_outputs(4895)) or (layer0_outputs(4982));
    outputs(6856) <= (layer0_outputs(3091)) or (layer0_outputs(989));
    outputs(6857) <= not((layer0_outputs(7060)) and (layer0_outputs(5935)));
    outputs(6858) <= layer0_outputs(3012);
    outputs(6859) <= not((layer0_outputs(1344)) and (layer0_outputs(1819)));
    outputs(6860) <= (layer0_outputs(4301)) and (layer0_outputs(7255));
    outputs(6861) <= layer0_outputs(7625);
    outputs(6862) <= layer0_outputs(2441);
    outputs(6863) <= not(layer0_outputs(3720));
    outputs(6864) <= not(layer0_outputs(2756));
    outputs(6865) <= (layer0_outputs(1200)) or (layer0_outputs(5994));
    outputs(6866) <= (layer0_outputs(292)) and not (layer0_outputs(458));
    outputs(6867) <= not((layer0_outputs(7635)) xor (layer0_outputs(4378)));
    outputs(6868) <= not((layer0_outputs(6262)) xor (layer0_outputs(6515)));
    outputs(6869) <= not((layer0_outputs(3447)) xor (layer0_outputs(5021)));
    outputs(6870) <= not((layer0_outputs(5544)) xor (layer0_outputs(1478)));
    outputs(6871) <= layer0_outputs(2544);
    outputs(6872) <= not((layer0_outputs(3063)) xor (layer0_outputs(7107)));
    outputs(6873) <= layer0_outputs(345);
    outputs(6874) <= layer0_outputs(4986);
    outputs(6875) <= not((layer0_outputs(1684)) xor (layer0_outputs(4051)));
    outputs(6876) <= not(layer0_outputs(3597));
    outputs(6877) <= (layer0_outputs(2857)) or (layer0_outputs(5280));
    outputs(6878) <= not(layer0_outputs(7465));
    outputs(6879) <= layer0_outputs(7464);
    outputs(6880) <= layer0_outputs(3749);
    outputs(6881) <= (layer0_outputs(7017)) xor (layer0_outputs(7422));
    outputs(6882) <= not(layer0_outputs(4944));
    outputs(6883) <= layer0_outputs(1949);
    outputs(6884) <= not(layer0_outputs(1736));
    outputs(6885) <= not((layer0_outputs(1178)) and (layer0_outputs(3408)));
    outputs(6886) <= not(layer0_outputs(3428));
    outputs(6887) <= not((layer0_outputs(1840)) or (layer0_outputs(974)));
    outputs(6888) <= (layer0_outputs(5051)) xor (layer0_outputs(1883));
    outputs(6889) <= (layer0_outputs(321)) xor (layer0_outputs(469));
    outputs(6890) <= layer0_outputs(1845);
    outputs(6891) <= not((layer0_outputs(3264)) xor (layer0_outputs(1065)));
    outputs(6892) <= layer0_outputs(2928);
    outputs(6893) <= not(layer0_outputs(5686));
    outputs(6894) <= (layer0_outputs(1732)) or (layer0_outputs(3088));
    outputs(6895) <= not(layer0_outputs(3214));
    outputs(6896) <= layer0_outputs(119);
    outputs(6897) <= (layer0_outputs(7602)) xor (layer0_outputs(2649));
    outputs(6898) <= not(layer0_outputs(2895));
    outputs(6899) <= (layer0_outputs(5434)) or (layer0_outputs(7133));
    outputs(6900) <= layer0_outputs(3656);
    outputs(6901) <= not(layer0_outputs(3403)) or (layer0_outputs(3210));
    outputs(6902) <= not(layer0_outputs(1568));
    outputs(6903) <= not(layer0_outputs(2658)) or (layer0_outputs(3415));
    outputs(6904) <= layer0_outputs(2704);
    outputs(6905) <= not((layer0_outputs(4475)) xor (layer0_outputs(2730)));
    outputs(6906) <= layer0_outputs(4450);
    outputs(6907) <= not(layer0_outputs(6518));
    outputs(6908) <= (layer0_outputs(2260)) and (layer0_outputs(3128));
    outputs(6909) <= (layer0_outputs(7106)) and not (layer0_outputs(4409));
    outputs(6910) <= not(layer0_outputs(4439)) or (layer0_outputs(3374));
    outputs(6911) <= not((layer0_outputs(5907)) xor (layer0_outputs(1143)));
    outputs(6912) <= layer0_outputs(3599);
    outputs(6913) <= (layer0_outputs(3668)) xor (layer0_outputs(6442));
    outputs(6914) <= not(layer0_outputs(4443));
    outputs(6915) <= not(layer0_outputs(1105)) or (layer0_outputs(1493));
    outputs(6916) <= (layer0_outputs(2891)) and not (layer0_outputs(821));
    outputs(6917) <= not((layer0_outputs(236)) or (layer0_outputs(1916)));
    outputs(6918) <= not(layer0_outputs(6066));
    outputs(6919) <= not((layer0_outputs(2245)) and (layer0_outputs(5862)));
    outputs(6920) <= layer0_outputs(1632);
    outputs(6921) <= not(layer0_outputs(5655));
    outputs(6922) <= layer0_outputs(6550);
    outputs(6923) <= layer0_outputs(6235);
    outputs(6924) <= not(layer0_outputs(481));
    outputs(6925) <= layer0_outputs(797);
    outputs(6926) <= (layer0_outputs(532)) and not (layer0_outputs(212));
    outputs(6927) <= (layer0_outputs(1195)) xor (layer0_outputs(99));
    outputs(6928) <= (layer0_outputs(6476)) and not (layer0_outputs(7520));
    outputs(6929) <= not((layer0_outputs(4618)) or (layer0_outputs(2696)));
    outputs(6930) <= (layer0_outputs(1145)) xor (layer0_outputs(5981));
    outputs(6931) <= (layer0_outputs(2741)) xor (layer0_outputs(5598));
    outputs(6932) <= not((layer0_outputs(2940)) xor (layer0_outputs(5169)));
    outputs(6933) <= not(layer0_outputs(3187));
    outputs(6934) <= (layer0_outputs(4415)) xor (layer0_outputs(3994));
    outputs(6935) <= not(layer0_outputs(7545)) or (layer0_outputs(1659));
    outputs(6936) <= not((layer0_outputs(6887)) and (layer0_outputs(6127)));
    outputs(6937) <= not((layer0_outputs(3201)) or (layer0_outputs(28)));
    outputs(6938) <= (layer0_outputs(5209)) and not (layer0_outputs(5674));
    outputs(6939) <= not((layer0_outputs(467)) or (layer0_outputs(1321)));
    outputs(6940) <= layer0_outputs(2136);
    outputs(6941) <= (layer0_outputs(7169)) or (layer0_outputs(3869));
    outputs(6942) <= layer0_outputs(1061);
    outputs(6943) <= layer0_outputs(3034);
    outputs(6944) <= layer0_outputs(1539);
    outputs(6945) <= layer0_outputs(2361);
    outputs(6946) <= not(layer0_outputs(1689));
    outputs(6947) <= not(layer0_outputs(4530));
    outputs(6948) <= not(layer0_outputs(5394));
    outputs(6949) <= not(layer0_outputs(473));
    outputs(6950) <= not((layer0_outputs(2410)) xor (layer0_outputs(524)));
    outputs(6951) <= layer0_outputs(3594);
    outputs(6952) <= layer0_outputs(3607);
    outputs(6953) <= layer0_outputs(4462);
    outputs(6954) <= not((layer0_outputs(153)) xor (layer0_outputs(792)));
    outputs(6955) <= not(layer0_outputs(2780));
    outputs(6956) <= layer0_outputs(6957);
    outputs(6957) <= (layer0_outputs(5275)) xor (layer0_outputs(4850));
    outputs(6958) <= not(layer0_outputs(4773)) or (layer0_outputs(5742));
    outputs(6959) <= not((layer0_outputs(1626)) or (layer0_outputs(6458)));
    outputs(6960) <= not((layer0_outputs(7223)) or (layer0_outputs(6967)));
    outputs(6961) <= layer0_outputs(492);
    outputs(6962) <= not(layer0_outputs(354));
    outputs(6963) <= not(layer0_outputs(4449));
    outputs(6964) <= layer0_outputs(4160);
    outputs(6965) <= layer0_outputs(5242);
    outputs(6966) <= (layer0_outputs(1034)) and not (layer0_outputs(6643));
    outputs(6967) <= layer0_outputs(1957);
    outputs(6968) <= not((layer0_outputs(2261)) xor (layer0_outputs(5600)));
    outputs(6969) <= (layer0_outputs(1814)) and (layer0_outputs(3462));
    outputs(6970) <= not((layer0_outputs(738)) or (layer0_outputs(1735)));
    outputs(6971) <= (layer0_outputs(3892)) and not (layer0_outputs(852));
    outputs(6972) <= layer0_outputs(3139);
    outputs(6973) <= not(layer0_outputs(535));
    outputs(6974) <= not(layer0_outputs(4219));
    outputs(6975) <= layer0_outputs(3);
    outputs(6976) <= not(layer0_outputs(4529));
    outputs(6977) <= not((layer0_outputs(3677)) or (layer0_outputs(4452)));
    outputs(6978) <= layer0_outputs(7065);
    outputs(6979) <= not(layer0_outputs(6692));
    outputs(6980) <= not((layer0_outputs(6383)) and (layer0_outputs(3967)));
    outputs(6981) <= layer0_outputs(1555);
    outputs(6982) <= (layer0_outputs(1543)) and not (layer0_outputs(7325));
    outputs(6983) <= not(layer0_outputs(4347));
    outputs(6984) <= not((layer0_outputs(2161)) and (layer0_outputs(3554)));
    outputs(6985) <= (layer0_outputs(3558)) and not (layer0_outputs(4461));
    outputs(6986) <= not(layer0_outputs(7487));
    outputs(6987) <= not((layer0_outputs(7615)) or (layer0_outputs(3745)));
    outputs(6988) <= not(layer0_outputs(6395));
    outputs(6989) <= not((layer0_outputs(3686)) xor (layer0_outputs(3431)));
    outputs(6990) <= layer0_outputs(3182);
    outputs(6991) <= not(layer0_outputs(1851));
    outputs(6992) <= layer0_outputs(1688);
    outputs(6993) <= not(layer0_outputs(4502)) or (layer0_outputs(3583));
    outputs(6994) <= (layer0_outputs(3278)) and not (layer0_outputs(4299));
    outputs(6995) <= (layer0_outputs(5929)) or (layer0_outputs(6264));
    outputs(6996) <= not(layer0_outputs(1582));
    outputs(6997) <= (layer0_outputs(2838)) and not (layer0_outputs(7499));
    outputs(6998) <= (layer0_outputs(1209)) and not (layer0_outputs(5541));
    outputs(6999) <= not(layer0_outputs(5394));
    outputs(7000) <= (layer0_outputs(5428)) and not (layer0_outputs(7564));
    outputs(7001) <= not(layer0_outputs(5322)) or (layer0_outputs(3626));
    outputs(7002) <= layer0_outputs(3484);
    outputs(7003) <= (layer0_outputs(251)) and not (layer0_outputs(239));
    outputs(7004) <= (layer0_outputs(3361)) xor (layer0_outputs(2963));
    outputs(7005) <= (layer0_outputs(2081)) xor (layer0_outputs(1809));
    outputs(7006) <= layer0_outputs(3464);
    outputs(7007) <= not((layer0_outputs(5262)) xor (layer0_outputs(3012)));
    outputs(7008) <= (layer0_outputs(2700)) xor (layer0_outputs(1207));
    outputs(7009) <= layer0_outputs(5458);
    outputs(7010) <= (layer0_outputs(1031)) and (layer0_outputs(5448));
    outputs(7011) <= not(layer0_outputs(7019));
    outputs(7012) <= layer0_outputs(4053);
    outputs(7013) <= not(layer0_outputs(3115)) or (layer0_outputs(5234));
    outputs(7014) <= not((layer0_outputs(240)) xor (layer0_outputs(1231)));
    outputs(7015) <= not(layer0_outputs(6335));
    outputs(7016) <= not(layer0_outputs(2162));
    outputs(7017) <= not((layer0_outputs(986)) or (layer0_outputs(4000)));
    outputs(7018) <= not(layer0_outputs(7561));
    outputs(7019) <= not(layer0_outputs(1322));
    outputs(7020) <= layer0_outputs(3255);
    outputs(7021) <= layer0_outputs(1528);
    outputs(7022) <= (layer0_outputs(1411)) and not (layer0_outputs(1963));
    outputs(7023) <= (layer0_outputs(3253)) and not (layer0_outputs(187));
    outputs(7024) <= not((layer0_outputs(4321)) xor (layer0_outputs(1806)));
    outputs(7025) <= not((layer0_outputs(2064)) or (layer0_outputs(196)));
    outputs(7026) <= (layer0_outputs(877)) xor (layer0_outputs(6458));
    outputs(7027) <= not(layer0_outputs(4431));
    outputs(7028) <= not(layer0_outputs(6087));
    outputs(7029) <= not(layer0_outputs(7192));
    outputs(7030) <= not((layer0_outputs(7109)) or (layer0_outputs(645)));
    outputs(7031) <= not((layer0_outputs(1367)) or (layer0_outputs(7025)));
    outputs(7032) <= not(layer0_outputs(3737));
    outputs(7033) <= not(layer0_outputs(3569));
    outputs(7034) <= not((layer0_outputs(2910)) xor (layer0_outputs(5891)));
    outputs(7035) <= layer0_outputs(1767);
    outputs(7036) <= layer0_outputs(494);
    outputs(7037) <= (layer0_outputs(1418)) xor (layer0_outputs(6325));
    outputs(7038) <= layer0_outputs(3857);
    outputs(7039) <= not(layer0_outputs(4662));
    outputs(7040) <= not((layer0_outputs(7263)) xor (layer0_outputs(4831)));
    outputs(7041) <= not((layer0_outputs(3406)) or (layer0_outputs(771)));
    outputs(7042) <= not(layer0_outputs(5040)) or (layer0_outputs(1203));
    outputs(7043) <= not(layer0_outputs(6814));
    outputs(7044) <= layer0_outputs(2048);
    outputs(7045) <= (layer0_outputs(7548)) and not (layer0_outputs(6775));
    outputs(7046) <= layer0_outputs(1461);
    outputs(7047) <= layer0_outputs(2209);
    outputs(7048) <= layer0_outputs(3646);
    outputs(7049) <= (layer0_outputs(1737)) and (layer0_outputs(2169));
    outputs(7050) <= not(layer0_outputs(6514));
    outputs(7051) <= not((layer0_outputs(5461)) xor (layer0_outputs(5735)));
    outputs(7052) <= not(layer0_outputs(2571));
    outputs(7053) <= not(layer0_outputs(7048));
    outputs(7054) <= (layer0_outputs(3572)) and (layer0_outputs(4832));
    outputs(7055) <= not((layer0_outputs(2571)) or (layer0_outputs(4709)));
    outputs(7056) <= not((layer0_outputs(4929)) or (layer0_outputs(4949)));
    outputs(7057) <= layer0_outputs(5274);
    outputs(7058) <= not((layer0_outputs(1556)) or (layer0_outputs(585)));
    outputs(7059) <= layer0_outputs(674);
    outputs(7060) <= not(layer0_outputs(2195));
    outputs(7061) <= not(layer0_outputs(6876));
    outputs(7062) <= (layer0_outputs(122)) and not (layer0_outputs(5102));
    outputs(7063) <= not((layer0_outputs(4001)) xor (layer0_outputs(3880)));
    outputs(7064) <= not((layer0_outputs(5654)) xor (layer0_outputs(371)));
    outputs(7065) <= not(layer0_outputs(6623));
    outputs(7066) <= (layer0_outputs(4623)) xor (layer0_outputs(4306));
    outputs(7067) <= not(layer0_outputs(1369));
    outputs(7068) <= not(layer0_outputs(5349)) or (layer0_outputs(5007));
    outputs(7069) <= not(layer0_outputs(7602));
    outputs(7070) <= not(layer0_outputs(3836));
    outputs(7071) <= not(layer0_outputs(5631));
    outputs(7072) <= not((layer0_outputs(4845)) or (layer0_outputs(405)));
    outputs(7073) <= (layer0_outputs(3237)) and not (layer0_outputs(573));
    outputs(7074) <= layer0_outputs(2496);
    outputs(7075) <= layer0_outputs(417);
    outputs(7076) <= not(layer0_outputs(4439));
    outputs(7077) <= not((layer0_outputs(10)) or (layer0_outputs(2214)));
    outputs(7078) <= not(layer0_outputs(6820));
    outputs(7079) <= layer0_outputs(5413);
    outputs(7080) <= not((layer0_outputs(2028)) xor (layer0_outputs(7296)));
    outputs(7081) <= layer0_outputs(7519);
    outputs(7082) <= layer0_outputs(1635);
    outputs(7083) <= (layer0_outputs(5610)) xor (layer0_outputs(718));
    outputs(7084) <= not((layer0_outputs(3910)) xor (layer0_outputs(5985)));
    outputs(7085) <= not(layer0_outputs(3453));
    outputs(7086) <= not(layer0_outputs(988));
    outputs(7087) <= layer0_outputs(4053);
    outputs(7088) <= layer0_outputs(2421);
    outputs(7089) <= not((layer0_outputs(4093)) or (layer0_outputs(38)));
    outputs(7090) <= (layer0_outputs(6821)) and (layer0_outputs(1425));
    outputs(7091) <= not((layer0_outputs(2547)) or (layer0_outputs(5339)));
    outputs(7092) <= (layer0_outputs(6257)) and not (layer0_outputs(2029));
    outputs(7093) <= not(layer0_outputs(1739)) or (layer0_outputs(983));
    outputs(7094) <= not((layer0_outputs(7219)) and (layer0_outputs(4923)));
    outputs(7095) <= not((layer0_outputs(5749)) and (layer0_outputs(1679)));
    outputs(7096) <= not(layer0_outputs(954));
    outputs(7097) <= layer0_outputs(2108);
    outputs(7098) <= not(layer0_outputs(3452));
    outputs(7099) <= not(layer0_outputs(2720));
    outputs(7100) <= layer0_outputs(5468);
    outputs(7101) <= not(layer0_outputs(7430));
    outputs(7102) <= (layer0_outputs(5956)) and (layer0_outputs(2520));
    outputs(7103) <= layer0_outputs(1681);
    outputs(7104) <= (layer0_outputs(1879)) xor (layer0_outputs(6264));
    outputs(7105) <= not(layer0_outputs(4213)) or (layer0_outputs(7328));
    outputs(7106) <= not(layer0_outputs(6136));
    outputs(7107) <= layer0_outputs(3451);
    outputs(7108) <= not(layer0_outputs(3493));
    outputs(7109) <= (layer0_outputs(6921)) xor (layer0_outputs(4534));
    outputs(7110) <= layer0_outputs(6181);
    outputs(7111) <= layer0_outputs(199);
    outputs(7112) <= not(layer0_outputs(5620));
    outputs(7113) <= not(layer0_outputs(1078));
    outputs(7114) <= (layer0_outputs(3478)) and not (layer0_outputs(2069));
    outputs(7115) <= (layer0_outputs(3516)) and not (layer0_outputs(2612));
    outputs(7116) <= layer0_outputs(890);
    outputs(7117) <= (layer0_outputs(4154)) and not (layer0_outputs(6412));
    outputs(7118) <= not((layer0_outputs(3863)) xor (layer0_outputs(7070)));
    outputs(7119) <= (layer0_outputs(1642)) or (layer0_outputs(4004));
    outputs(7120) <= not(layer0_outputs(6120));
    outputs(7121) <= not(layer0_outputs(3470));
    outputs(7122) <= not(layer0_outputs(1524)) or (layer0_outputs(5105));
    outputs(7123) <= (layer0_outputs(6868)) or (layer0_outputs(5704));
    outputs(7124) <= not(layer0_outputs(3569));
    outputs(7125) <= (layer0_outputs(5487)) and not (layer0_outputs(6401));
    outputs(7126) <= layer0_outputs(6631);
    outputs(7127) <= (layer0_outputs(7151)) xor (layer0_outputs(3794));
    outputs(7128) <= (layer0_outputs(3105)) and not (layer0_outputs(317));
    outputs(7129) <= layer0_outputs(2625);
    outputs(7130) <= not(layer0_outputs(7266));
    outputs(7131) <= not((layer0_outputs(3615)) or (layer0_outputs(606)));
    outputs(7132) <= layer0_outputs(2908);
    outputs(7133) <= (layer0_outputs(1262)) and (layer0_outputs(5764));
    outputs(7134) <= not((layer0_outputs(7330)) or (layer0_outputs(608)));
    outputs(7135) <= layer0_outputs(621);
    outputs(7136) <= (layer0_outputs(339)) and not (layer0_outputs(6693));
    outputs(7137) <= not((layer0_outputs(5272)) xor (layer0_outputs(4364)));
    outputs(7138) <= (layer0_outputs(1704)) and not (layer0_outputs(6781));
    outputs(7139) <= (layer0_outputs(2027)) and not (layer0_outputs(1610));
    outputs(7140) <= (layer0_outputs(302)) and (layer0_outputs(7442));
    outputs(7141) <= not(layer0_outputs(3883));
    outputs(7142) <= (layer0_outputs(7463)) and (layer0_outputs(2719));
    outputs(7143) <= (layer0_outputs(3840)) and not (layer0_outputs(6493));
    outputs(7144) <= not(layer0_outputs(6093));
    outputs(7145) <= layer0_outputs(3823);
    outputs(7146) <= (layer0_outputs(7369)) and not (layer0_outputs(1159));
    outputs(7147) <= layer0_outputs(3407);
    outputs(7148) <= (layer0_outputs(4538)) xor (layer0_outputs(6627));
    outputs(7149) <= (layer0_outputs(7328)) and not (layer0_outputs(4809));
    outputs(7150) <= not(layer0_outputs(722));
    outputs(7151) <= layer0_outputs(2771);
    outputs(7152) <= layer0_outputs(307);
    outputs(7153) <= not(layer0_outputs(5267)) or (layer0_outputs(2570));
    outputs(7154) <= layer0_outputs(1575);
    outputs(7155) <= (layer0_outputs(3789)) and not (layer0_outputs(4473));
    outputs(7156) <= not(layer0_outputs(4259));
    outputs(7157) <= layer0_outputs(4420);
    outputs(7158) <= not(layer0_outputs(7569));
    outputs(7159) <= (layer0_outputs(2978)) and (layer0_outputs(534));
    outputs(7160) <= not((layer0_outputs(6789)) xor (layer0_outputs(7172)));
    outputs(7161) <= layer0_outputs(678);
    outputs(7162) <= not((layer0_outputs(6416)) xor (layer0_outputs(4900)));
    outputs(7163) <= layer0_outputs(5575);
    outputs(7164) <= layer0_outputs(1579);
    outputs(7165) <= not(layer0_outputs(1771));
    outputs(7166) <= layer0_outputs(2537);
    outputs(7167) <= layer0_outputs(2729);
    outputs(7168) <= not(layer0_outputs(4184));
    outputs(7169) <= not(layer0_outputs(6211));
    outputs(7170) <= (layer0_outputs(1882)) xor (layer0_outputs(2572));
    outputs(7171) <= (layer0_outputs(575)) and not (layer0_outputs(6155));
    outputs(7172) <= (layer0_outputs(3721)) and not (layer0_outputs(4542));
    outputs(7173) <= not((layer0_outputs(1054)) and (layer0_outputs(183)));
    outputs(7174) <= (layer0_outputs(7366)) and (layer0_outputs(4115));
    outputs(7175) <= not((layer0_outputs(4047)) and (layer0_outputs(4936)));
    outputs(7176) <= (layer0_outputs(2228)) and (layer0_outputs(5732));
    outputs(7177) <= not(layer0_outputs(4138)) or (layer0_outputs(2328));
    outputs(7178) <= (layer0_outputs(6332)) and (layer0_outputs(4752));
    outputs(7179) <= layer0_outputs(6945);
    outputs(7180) <= not((layer0_outputs(6622)) or (layer0_outputs(6381)));
    outputs(7181) <= layer0_outputs(6101);
    outputs(7182) <= (layer0_outputs(7440)) xor (layer0_outputs(6831));
    outputs(7183) <= not(layer0_outputs(7629));
    outputs(7184) <= (layer0_outputs(6477)) and not (layer0_outputs(7157));
    outputs(7185) <= (layer0_outputs(5095)) and not (layer0_outputs(6784));
    outputs(7186) <= (layer0_outputs(2850)) and not (layer0_outputs(7112));
    outputs(7187) <= layer0_outputs(2908);
    outputs(7188) <= (layer0_outputs(5128)) and not (layer0_outputs(4669));
    outputs(7189) <= layer0_outputs(1985);
    outputs(7190) <= not(layer0_outputs(5398));
    outputs(7191) <= not((layer0_outputs(5464)) and (layer0_outputs(789)));
    outputs(7192) <= not((layer0_outputs(1770)) or (layer0_outputs(1316)));
    outputs(7193) <= layer0_outputs(4012);
    outputs(7194) <= layer0_outputs(3711);
    outputs(7195) <= (layer0_outputs(4555)) and not (layer0_outputs(1426));
    outputs(7196) <= layer0_outputs(5195);
    outputs(7197) <= layer0_outputs(3809);
    outputs(7198) <= not(layer0_outputs(3231)) or (layer0_outputs(2739));
    outputs(7199) <= layer0_outputs(5146);
    outputs(7200) <= not(layer0_outputs(4647));
    outputs(7201) <= not((layer0_outputs(7082)) and (layer0_outputs(1496)));
    outputs(7202) <= not((layer0_outputs(325)) xor (layer0_outputs(3871)));
    outputs(7203) <= (layer0_outputs(296)) xor (layer0_outputs(3910));
    outputs(7204) <= not((layer0_outputs(3354)) xor (layer0_outputs(2790)));
    outputs(7205) <= not(layer0_outputs(7332));
    outputs(7206) <= not((layer0_outputs(1410)) or (layer0_outputs(2416)));
    outputs(7207) <= not(layer0_outputs(2936));
    outputs(7208) <= not(layer0_outputs(5883));
    outputs(7209) <= (layer0_outputs(6723)) and not (layer0_outputs(1306));
    outputs(7210) <= not((layer0_outputs(744)) or (layer0_outputs(4376)));
    outputs(7211) <= (layer0_outputs(6521)) xor (layer0_outputs(889));
    outputs(7212) <= (layer0_outputs(1364)) and (layer0_outputs(4841));
    outputs(7213) <= not(layer0_outputs(2701));
    outputs(7214) <= (layer0_outputs(3322)) and not (layer0_outputs(284));
    outputs(7215) <= layer0_outputs(6954);
    outputs(7216) <= not(layer0_outputs(3963));
    outputs(7217) <= not((layer0_outputs(5463)) xor (layer0_outputs(2383)));
    outputs(7218) <= not(layer0_outputs(7118));
    outputs(7219) <= not(layer0_outputs(1961));
    outputs(7220) <= not((layer0_outputs(7572)) or (layer0_outputs(2982)));
    outputs(7221) <= layer0_outputs(2921);
    outputs(7222) <= (layer0_outputs(1460)) xor (layer0_outputs(7343));
    outputs(7223) <= not(layer0_outputs(3793));
    outputs(7224) <= (layer0_outputs(2685)) and not (layer0_outputs(7254));
    outputs(7225) <= not((layer0_outputs(998)) and (layer0_outputs(3819)));
    outputs(7226) <= (layer0_outputs(3560)) xor (layer0_outputs(3482));
    outputs(7227) <= (layer0_outputs(5837)) and not (layer0_outputs(4711));
    outputs(7228) <= (layer0_outputs(5154)) and (layer0_outputs(995));
    outputs(7229) <= (layer0_outputs(6236)) and (layer0_outputs(6586));
    outputs(7230) <= not(layer0_outputs(7317));
    outputs(7231) <= (layer0_outputs(4397)) and not (layer0_outputs(3865));
    outputs(7232) <= not((layer0_outputs(4618)) xor (layer0_outputs(5056)));
    outputs(7233) <= '0';
    outputs(7234) <= layer0_outputs(4012);
    outputs(7235) <= layer0_outputs(6024);
    outputs(7236) <= (layer0_outputs(7654)) xor (layer0_outputs(291));
    outputs(7237) <= not(layer0_outputs(391));
    outputs(7238) <= (layer0_outputs(12)) and not (layer0_outputs(5919));
    outputs(7239) <= not(layer0_outputs(5790));
    outputs(7240) <= not((layer0_outputs(1089)) and (layer0_outputs(3399)));
    outputs(7241) <= not((layer0_outputs(5221)) or (layer0_outputs(2832)));
    outputs(7242) <= layer0_outputs(6525);
    outputs(7243) <= (layer0_outputs(2943)) and not (layer0_outputs(3249));
    outputs(7244) <= not((layer0_outputs(212)) or (layer0_outputs(4463)));
    outputs(7245) <= (layer0_outputs(1722)) and (layer0_outputs(1767));
    outputs(7246) <= layer0_outputs(2868);
    outputs(7247) <= not(layer0_outputs(7186));
    outputs(7248) <= (layer0_outputs(1354)) and not (layer0_outputs(542));
    outputs(7249) <= layer0_outputs(4177);
    outputs(7250) <= (layer0_outputs(1507)) and not (layer0_outputs(2095));
    outputs(7251) <= layer0_outputs(6407);
    outputs(7252) <= not((layer0_outputs(7056)) xor (layer0_outputs(2792)));
    outputs(7253) <= not(layer0_outputs(7447));
    outputs(7254) <= not((layer0_outputs(5371)) or (layer0_outputs(734)));
    outputs(7255) <= not((layer0_outputs(6621)) xor (layer0_outputs(868)));
    outputs(7256) <= not((layer0_outputs(861)) or (layer0_outputs(4694)));
    outputs(7257) <= not(layer0_outputs(7557));
    outputs(7258) <= layer0_outputs(3456);
    outputs(7259) <= not(layer0_outputs(3924));
    outputs(7260) <= layer0_outputs(3257);
    outputs(7261) <= layer0_outputs(5915);
    outputs(7262) <= not(layer0_outputs(4875));
    outputs(7263) <= not((layer0_outputs(3888)) or (layer0_outputs(4149)));
    outputs(7264) <= not((layer0_outputs(2749)) or (layer0_outputs(7568)));
    outputs(7265) <= not(layer0_outputs(813));
    outputs(7266) <= (layer0_outputs(6742)) and (layer0_outputs(1182));
    outputs(7267) <= (layer0_outputs(3609)) and not (layer0_outputs(2540));
    outputs(7268) <= (layer0_outputs(2996)) and not (layer0_outputs(5435));
    outputs(7269) <= not(layer0_outputs(5570));
    outputs(7270) <= not(layer0_outputs(3216));
    outputs(7271) <= layer0_outputs(397);
    outputs(7272) <= layer0_outputs(399);
    outputs(7273) <= not((layer0_outputs(5897)) xor (layer0_outputs(6426)));
    outputs(7274) <= layer0_outputs(2719);
    outputs(7275) <= layer0_outputs(49);
    outputs(7276) <= layer0_outputs(1661);
    outputs(7277) <= layer0_outputs(7519);
    outputs(7278) <= layer0_outputs(636);
    outputs(7279) <= layer0_outputs(6779);
    outputs(7280) <= (layer0_outputs(904)) xor (layer0_outputs(3839));
    outputs(7281) <= layer0_outputs(4464);
    outputs(7282) <= layer0_outputs(3952);
    outputs(7283) <= not(layer0_outputs(845));
    outputs(7284) <= not(layer0_outputs(7118));
    outputs(7285) <= (layer0_outputs(2744)) and not (layer0_outputs(4835));
    outputs(7286) <= not(layer0_outputs(7064));
    outputs(7287) <= not(layer0_outputs(5006)) or (layer0_outputs(26));
    outputs(7288) <= (layer0_outputs(4998)) xor (layer0_outputs(6674));
    outputs(7289) <= layer0_outputs(3498);
    outputs(7290) <= not(layer0_outputs(783));
    outputs(7291) <= (layer0_outputs(1856)) and (layer0_outputs(7174));
    outputs(7292) <= layer0_outputs(3419);
    outputs(7293) <= (layer0_outputs(5402)) and not (layer0_outputs(1309));
    outputs(7294) <= (layer0_outputs(7061)) and not (layer0_outputs(2701));
    outputs(7295) <= layer0_outputs(6821);
    outputs(7296) <= layer0_outputs(6051);
    outputs(7297) <= not(layer0_outputs(1449));
    outputs(7298) <= layer0_outputs(6338);
    outputs(7299) <= layer0_outputs(400);
    outputs(7300) <= (layer0_outputs(5451)) and not (layer0_outputs(5736));
    outputs(7301) <= layer0_outputs(3920);
    outputs(7302) <= (layer0_outputs(4580)) xor (layer0_outputs(1808));
    outputs(7303) <= (layer0_outputs(3790)) or (layer0_outputs(1844));
    outputs(7304) <= layer0_outputs(1748);
    outputs(7305) <= layer0_outputs(444);
    outputs(7306) <= (layer0_outputs(2755)) and not (layer0_outputs(2600));
    outputs(7307) <= not(layer0_outputs(1255));
    outputs(7308) <= not(layer0_outputs(4376));
    outputs(7309) <= not((layer0_outputs(4700)) xor (layer0_outputs(3385)));
    outputs(7310) <= layer0_outputs(5756);
    outputs(7311) <= not((layer0_outputs(1136)) xor (layer0_outputs(498)));
    outputs(7312) <= (layer0_outputs(2506)) and not (layer0_outputs(6759));
    outputs(7313) <= layer0_outputs(2262);
    outputs(7314) <= not(layer0_outputs(1430)) or (layer0_outputs(2609));
    outputs(7315) <= (layer0_outputs(2229)) and (layer0_outputs(3355));
    outputs(7316) <= not((layer0_outputs(175)) xor (layer0_outputs(6839)));
    outputs(7317) <= not(layer0_outputs(4300));
    outputs(7318) <= layer0_outputs(5731);
    outputs(7319) <= layer0_outputs(1668);
    outputs(7320) <= not((layer0_outputs(6160)) or (layer0_outputs(4003)));
    outputs(7321) <= (layer0_outputs(5012)) and not (layer0_outputs(4331));
    outputs(7322) <= layer0_outputs(217);
    outputs(7323) <= (layer0_outputs(4233)) xor (layer0_outputs(2339));
    outputs(7324) <= layer0_outputs(2803);
    outputs(7325) <= (layer0_outputs(2355)) and not (layer0_outputs(3876));
    outputs(7326) <= layer0_outputs(4257);
    outputs(7327) <= layer0_outputs(2149);
    outputs(7328) <= layer0_outputs(6959);
    outputs(7329) <= (layer0_outputs(7417)) and not (layer0_outputs(6860));
    outputs(7330) <= layer0_outputs(6713);
    outputs(7331) <= layer0_outputs(1928);
    outputs(7332) <= not((layer0_outputs(4567)) or (layer0_outputs(6106)));
    outputs(7333) <= layer0_outputs(933);
    outputs(7334) <= layer0_outputs(6578);
    outputs(7335) <= (layer0_outputs(4559)) and not (layer0_outputs(1676));
    outputs(7336) <= layer0_outputs(6201);
    outputs(7337) <= layer0_outputs(3362);
    outputs(7338) <= not((layer0_outputs(989)) or (layer0_outputs(1599)));
    outputs(7339) <= (layer0_outputs(3065)) and not (layer0_outputs(7300));
    outputs(7340) <= (layer0_outputs(6230)) and (layer0_outputs(1345));
    outputs(7341) <= (layer0_outputs(2916)) and (layer0_outputs(4481));
    outputs(7342) <= (layer0_outputs(2283)) and not (layer0_outputs(3672));
    outputs(7343) <= not(layer0_outputs(5747));
    outputs(7344) <= (layer0_outputs(1897)) xor (layer0_outputs(5609));
    outputs(7345) <= not(layer0_outputs(5707));
    outputs(7346) <= not((layer0_outputs(3240)) or (layer0_outputs(1146)));
    outputs(7347) <= not(layer0_outputs(5332));
    outputs(7348) <= not((layer0_outputs(2488)) xor (layer0_outputs(951)));
    outputs(7349) <= (layer0_outputs(623)) and not (layer0_outputs(1144));
    outputs(7350) <= not((layer0_outputs(1610)) xor (layer0_outputs(3039)));
    outputs(7351) <= layer0_outputs(2009);
    outputs(7352) <= not(layer0_outputs(4112));
    outputs(7353) <= not(layer0_outputs(6004));
    outputs(7354) <= not(layer0_outputs(1456));
    outputs(7355) <= not(layer0_outputs(2117));
    outputs(7356) <= (layer0_outputs(7238)) and not (layer0_outputs(2150));
    outputs(7357) <= (layer0_outputs(3262)) and not (layer0_outputs(4759));
    outputs(7358) <= not((layer0_outputs(3148)) xor (layer0_outputs(7615)));
    outputs(7359) <= not(layer0_outputs(7596));
    outputs(7360) <= not(layer0_outputs(2468));
    outputs(7361) <= not((layer0_outputs(5399)) xor (layer0_outputs(3145)));
    outputs(7362) <= not(layer0_outputs(4678));
    outputs(7363) <= not((layer0_outputs(1973)) and (layer0_outputs(1342)));
    outputs(7364) <= layer0_outputs(5751);
    outputs(7365) <= not(layer0_outputs(5691));
    outputs(7366) <= not(layer0_outputs(3077));
    outputs(7367) <= not(layer0_outputs(6448));
    outputs(7368) <= (layer0_outputs(3533)) and not (layer0_outputs(7460));
    outputs(7369) <= not((layer0_outputs(4760)) and (layer0_outputs(6770)));
    outputs(7370) <= not((layer0_outputs(231)) xor (layer0_outputs(2472)));
    outputs(7371) <= not((layer0_outputs(7606)) or (layer0_outputs(2090)));
    outputs(7372) <= (layer0_outputs(4769)) and not (layer0_outputs(2455));
    outputs(7373) <= layer0_outputs(4591);
    outputs(7374) <= (layer0_outputs(2927)) and (layer0_outputs(220));
    outputs(7375) <= (layer0_outputs(2010)) and not (layer0_outputs(279));
    outputs(7376) <= (layer0_outputs(3544)) and not (layer0_outputs(5282));
    outputs(7377) <= not(layer0_outputs(7595));
    outputs(7378) <= not((layer0_outputs(6320)) xor (layer0_outputs(2292)));
    outputs(7379) <= (layer0_outputs(3975)) xor (layer0_outputs(1010));
    outputs(7380) <= layer0_outputs(4630);
    outputs(7381) <= layer0_outputs(1069);
    outputs(7382) <= not(layer0_outputs(7040));
    outputs(7383) <= not(layer0_outputs(3177));
    outputs(7384) <= layer0_outputs(564);
    outputs(7385) <= (layer0_outputs(512)) and not (layer0_outputs(1107));
    outputs(7386) <= not(layer0_outputs(2749));
    outputs(7387) <= layer0_outputs(2575);
    outputs(7388) <= not((layer0_outputs(4775)) and (layer0_outputs(2662)));
    outputs(7389) <= layer0_outputs(7032);
    outputs(7390) <= (layer0_outputs(4092)) xor (layer0_outputs(5699));
    outputs(7391) <= not((layer0_outputs(3968)) or (layer0_outputs(5964)));
    outputs(7392) <= not((layer0_outputs(2881)) xor (layer0_outputs(6445)));
    outputs(7393) <= layer0_outputs(1776);
    outputs(7394) <= layer0_outputs(2315);
    outputs(7395) <= (layer0_outputs(5227)) and (layer0_outputs(5374));
    outputs(7396) <= not(layer0_outputs(5061));
    outputs(7397) <= not((layer0_outputs(2648)) and (layer0_outputs(3992)));
    outputs(7398) <= not(layer0_outputs(4508)) or (layer0_outputs(1578));
    outputs(7399) <= not(layer0_outputs(5705));
    outputs(7400) <= not(layer0_outputs(6510));
    outputs(7401) <= not((layer0_outputs(4333)) xor (layer0_outputs(6509)));
    outputs(7402) <= layer0_outputs(1852);
    outputs(7403) <= not((layer0_outputs(4015)) or (layer0_outputs(5649)));
    outputs(7404) <= not(layer0_outputs(900));
    outputs(7405) <= (layer0_outputs(2288)) and (layer0_outputs(4997));
    outputs(7406) <= layer0_outputs(5557);
    outputs(7407) <= not((layer0_outputs(2453)) xor (layer0_outputs(3732)));
    outputs(7408) <= layer0_outputs(6581);
    outputs(7409) <= not(layer0_outputs(4493));
    outputs(7410) <= not((layer0_outputs(2215)) or (layer0_outputs(6305)));
    outputs(7411) <= (layer0_outputs(2369)) and (layer0_outputs(4945));
    outputs(7412) <= layer0_outputs(2838);
    outputs(7413) <= (layer0_outputs(6632)) and not (layer0_outputs(1291));
    outputs(7414) <= (layer0_outputs(742)) and (layer0_outputs(2643));
    outputs(7415) <= (layer0_outputs(4867)) xor (layer0_outputs(559));
    outputs(7416) <= layer0_outputs(1391);
    outputs(7417) <= not((layer0_outputs(7004)) or (layer0_outputs(7177)));
    outputs(7418) <= not((layer0_outputs(3712)) and (layer0_outputs(4395)));
    outputs(7419) <= not(layer0_outputs(570)) or (layer0_outputs(4812));
    outputs(7420) <= layer0_outputs(4553);
    outputs(7421) <= not(layer0_outputs(4980));
    outputs(7422) <= not(layer0_outputs(4024));
    outputs(7423) <= not(layer0_outputs(7394));
    outputs(7424) <= not(layer0_outputs(228));
    outputs(7425) <= (layer0_outputs(243)) and (layer0_outputs(7353));
    outputs(7426) <= not((layer0_outputs(4782)) xor (layer0_outputs(5422)));
    outputs(7427) <= not(layer0_outputs(5847));
    outputs(7428) <= (layer0_outputs(4499)) and (layer0_outputs(3306));
    outputs(7429) <= not(layer0_outputs(6068));
    outputs(7430) <= not((layer0_outputs(316)) xor (layer0_outputs(7446)));
    outputs(7431) <= not(layer0_outputs(4007));
    outputs(7432) <= not(layer0_outputs(5225));
    outputs(7433) <= (layer0_outputs(5625)) and (layer0_outputs(6869));
    outputs(7434) <= not(layer0_outputs(7430));
    outputs(7435) <= not((layer0_outputs(872)) or (layer0_outputs(2555)));
    outputs(7436) <= not((layer0_outputs(6427)) xor (layer0_outputs(1004)));
    outputs(7437) <= (layer0_outputs(89)) or (layer0_outputs(424));
    outputs(7438) <= layer0_outputs(3542);
    outputs(7439) <= not(layer0_outputs(3411));
    outputs(7440) <= layer0_outputs(3188);
    outputs(7441) <= not(layer0_outputs(6651));
    outputs(7442) <= not(layer0_outputs(6792));
    outputs(7443) <= (layer0_outputs(3242)) and (layer0_outputs(6372));
    outputs(7444) <= not(layer0_outputs(1462));
    outputs(7445) <= (layer0_outputs(3307)) or (layer0_outputs(2633));
    outputs(7446) <= not(layer0_outputs(411));
    outputs(7447) <= layer0_outputs(4401);
    outputs(7448) <= (layer0_outputs(3787)) xor (layer0_outputs(1269));
    outputs(7449) <= not((layer0_outputs(7307)) and (layer0_outputs(5712)));
    outputs(7450) <= (layer0_outputs(5251)) xor (layer0_outputs(5806));
    outputs(7451) <= not(layer0_outputs(6191)) or (layer0_outputs(3461));
    outputs(7452) <= (layer0_outputs(2263)) xor (layer0_outputs(4399));
    outputs(7453) <= (layer0_outputs(5765)) and (layer0_outputs(7135));
    outputs(7454) <= not((layer0_outputs(652)) xor (layer0_outputs(4514)));
    outputs(7455) <= not(layer0_outputs(855));
    outputs(7456) <= (layer0_outputs(7334)) or (layer0_outputs(2275));
    outputs(7457) <= not(layer0_outputs(1228));
    outputs(7458) <= not((layer0_outputs(7011)) xor (layer0_outputs(1212)));
    outputs(7459) <= (layer0_outputs(6955)) and (layer0_outputs(2252));
    outputs(7460) <= (layer0_outputs(4344)) and (layer0_outputs(3959));
    outputs(7461) <= not(layer0_outputs(4047));
    outputs(7462) <= (layer0_outputs(6229)) and not (layer0_outputs(6234));
    outputs(7463) <= layer0_outputs(1376);
    outputs(7464) <= not((layer0_outputs(4442)) xor (layer0_outputs(633)));
    outputs(7465) <= (layer0_outputs(1101)) and not (layer0_outputs(6719));
    outputs(7466) <= not((layer0_outputs(2279)) xor (layer0_outputs(5373)));
    outputs(7467) <= not((layer0_outputs(4774)) or (layer0_outputs(1420)));
    outputs(7468) <= not(layer0_outputs(326));
    outputs(7469) <= (layer0_outputs(437)) and not (layer0_outputs(3672));
    outputs(7470) <= not((layer0_outputs(3978)) or (layer0_outputs(5529)));
    outputs(7471) <= layer0_outputs(2900);
    outputs(7472) <= not(layer0_outputs(345));
    outputs(7473) <= (layer0_outputs(1833)) and not (layer0_outputs(4170));
    outputs(7474) <= (layer0_outputs(5627)) or (layer0_outputs(4719));
    outputs(7475) <= not(layer0_outputs(5790));
    outputs(7476) <= (layer0_outputs(3744)) and not (layer0_outputs(3002));
    outputs(7477) <= (layer0_outputs(4043)) and not (layer0_outputs(3866));
    outputs(7478) <= (layer0_outputs(5974)) and not (layer0_outputs(1551));
    outputs(7479) <= (layer0_outputs(4948)) and not (layer0_outputs(7044));
    outputs(7480) <= not((layer0_outputs(2971)) xor (layer0_outputs(5506)));
    outputs(7481) <= not(layer0_outputs(7648));
    outputs(7482) <= (layer0_outputs(5431)) and not (layer0_outputs(2459));
    outputs(7483) <= (layer0_outputs(6550)) and not (layer0_outputs(810));
    outputs(7484) <= not(layer0_outputs(4964));
    outputs(7485) <= (layer0_outputs(1581)) xor (layer0_outputs(4413));
    outputs(7486) <= not(layer0_outputs(1734));
    outputs(7487) <= layer0_outputs(280);
    outputs(7488) <= not(layer0_outputs(6691));
    outputs(7489) <= not(layer0_outputs(1811));
    outputs(7490) <= not((layer0_outputs(5481)) xor (layer0_outputs(7015)));
    outputs(7491) <= not(layer0_outputs(1217));
    outputs(7492) <= not((layer0_outputs(7036)) or (layer0_outputs(5881)));
    outputs(7493) <= (layer0_outputs(4600)) and not (layer0_outputs(2411));
    outputs(7494) <= not(layer0_outputs(5537));
    outputs(7495) <= (layer0_outputs(1627)) and not (layer0_outputs(1959));
    outputs(7496) <= not((layer0_outputs(6358)) or (layer0_outputs(3072)));
    outputs(7497) <= not((layer0_outputs(1922)) xor (layer0_outputs(5811)));
    outputs(7498) <= layer0_outputs(6978);
    outputs(7499) <= (layer0_outputs(2726)) and (layer0_outputs(1507));
    outputs(7500) <= layer0_outputs(3205);
    outputs(7501) <= layer0_outputs(2395);
    outputs(7502) <= not(layer0_outputs(6798));
    outputs(7503) <= not(layer0_outputs(3070));
    outputs(7504) <= layer0_outputs(5822);
    outputs(7505) <= not(layer0_outputs(5554));
    outputs(7506) <= not(layer0_outputs(2272));
    outputs(7507) <= layer0_outputs(3650);
    outputs(7508) <= not(layer0_outputs(1422)) or (layer0_outputs(5016));
    outputs(7509) <= not((layer0_outputs(4971)) or (layer0_outputs(6431)));
    outputs(7510) <= not(layer0_outputs(299));
    outputs(7511) <= (layer0_outputs(1188)) or (layer0_outputs(245));
    outputs(7512) <= not(layer0_outputs(4679)) or (layer0_outputs(1510));
    outputs(7513) <= (layer0_outputs(3897)) and not (layer0_outputs(3138));
    outputs(7514) <= not(layer0_outputs(3576));
    outputs(7515) <= layer0_outputs(2444);
    outputs(7516) <= layer0_outputs(2868);
    outputs(7517) <= not(layer0_outputs(2937));
    outputs(7518) <= not(layer0_outputs(3576));
    outputs(7519) <= '0';
    outputs(7520) <= not(layer0_outputs(959));
    outputs(7521) <= not((layer0_outputs(3059)) or (layer0_outputs(5872)));
    outputs(7522) <= layer0_outputs(647);
    outputs(7523) <= layer0_outputs(3768);
    outputs(7524) <= (layer0_outputs(4560)) xor (layer0_outputs(5532));
    outputs(7525) <= layer0_outputs(4752);
    outputs(7526) <= not(layer0_outputs(7538));
    outputs(7527) <= (layer0_outputs(5851)) xor (layer0_outputs(6173));
    outputs(7528) <= (layer0_outputs(1103)) xor (layer0_outputs(1677));
    outputs(7529) <= (layer0_outputs(7454)) and (layer0_outputs(1061));
    outputs(7530) <= not(layer0_outputs(544));
    outputs(7531) <= not(layer0_outputs(1743));
    outputs(7532) <= not((layer0_outputs(3589)) xor (layer0_outputs(1017)));
    outputs(7533) <= not(layer0_outputs(5040)) or (layer0_outputs(6685));
    outputs(7534) <= layer0_outputs(7010);
    outputs(7535) <= (layer0_outputs(6904)) or (layer0_outputs(3986));
    outputs(7536) <= (layer0_outputs(5959)) and (layer0_outputs(1552));
    outputs(7537) <= not(layer0_outputs(4137)) or (layer0_outputs(2698));
    outputs(7538) <= not(layer0_outputs(5064)) or (layer0_outputs(4197));
    outputs(7539) <= not(layer0_outputs(811));
    outputs(7540) <= layer0_outputs(1506);
    outputs(7541) <= layer0_outputs(2402);
    outputs(7542) <= (layer0_outputs(5364)) and not (layer0_outputs(239));
    outputs(7543) <= not(layer0_outputs(323));
    outputs(7544) <= not(layer0_outputs(7092));
    outputs(7545) <= (layer0_outputs(512)) and not (layer0_outputs(4005));
    outputs(7546) <= not((layer0_outputs(958)) or (layer0_outputs(2974)));
    outputs(7547) <= not((layer0_outputs(6602)) xor (layer0_outputs(5421)));
    outputs(7548) <= not(layer0_outputs(3221));
    outputs(7549) <= layer0_outputs(7272);
    outputs(7550) <= not(layer0_outputs(679));
    outputs(7551) <= (layer0_outputs(2753)) and (layer0_outputs(3153));
    outputs(7552) <= not((layer0_outputs(7124)) or (layer0_outputs(2906)));
    outputs(7553) <= not(layer0_outputs(7146));
    outputs(7554) <= layer0_outputs(3704);
    outputs(7555) <= not(layer0_outputs(2282));
    outputs(7556) <= not(layer0_outputs(7610)) or (layer0_outputs(1490));
    outputs(7557) <= layer0_outputs(156);
    outputs(7558) <= layer0_outputs(3318);
    outputs(7559) <= layer0_outputs(4380);
    outputs(7560) <= not((layer0_outputs(3618)) and (layer0_outputs(7436)));
    outputs(7561) <= layer0_outputs(5779);
    outputs(7562) <= not((layer0_outputs(2255)) xor (layer0_outputs(5563)));
    outputs(7563) <= (layer0_outputs(465)) xor (layer0_outputs(6170));
    outputs(7564) <= not(layer0_outputs(2478));
    outputs(7565) <= not(layer0_outputs(3550));
    outputs(7566) <= (layer0_outputs(5534)) and not (layer0_outputs(4508));
    outputs(7567) <= not((layer0_outputs(7110)) xor (layer0_outputs(6036)));
    outputs(7568) <= layer0_outputs(4778);
    outputs(7569) <= (layer0_outputs(5218)) xor (layer0_outputs(4327));
    outputs(7570) <= not((layer0_outputs(913)) and (layer0_outputs(4406)));
    outputs(7571) <= (layer0_outputs(646)) xor (layer0_outputs(6651));
    outputs(7572) <= not((layer0_outputs(633)) xor (layer0_outputs(7403)));
    outputs(7573) <= layer0_outputs(5078);
    outputs(7574) <= not(layer0_outputs(873));
    outputs(7575) <= not(layer0_outputs(4049));
    outputs(7576) <= not((layer0_outputs(6874)) xor (layer0_outputs(2233)));
    outputs(7577) <= not(layer0_outputs(5730));
    outputs(7578) <= layer0_outputs(931);
    outputs(7579) <= not((layer0_outputs(4551)) xor (layer0_outputs(5200)));
    outputs(7580) <= layer0_outputs(1635);
    outputs(7581) <= not(layer0_outputs(5248));
    outputs(7582) <= layer0_outputs(1782);
    outputs(7583) <= (layer0_outputs(7618)) and not (layer0_outputs(5515));
    outputs(7584) <= not(layer0_outputs(3127));
    outputs(7585) <= (layer0_outputs(2489)) and not (layer0_outputs(3402));
    outputs(7586) <= (layer0_outputs(4583)) and not (layer0_outputs(1146));
    outputs(7587) <= not(layer0_outputs(6043));
    outputs(7588) <= not((layer0_outputs(2436)) or (layer0_outputs(3838)));
    outputs(7589) <= not(layer0_outputs(1319));
    outputs(7590) <= (layer0_outputs(6022)) and not (layer0_outputs(1701));
    outputs(7591) <= layer0_outputs(2597);
    outputs(7592) <= not((layer0_outputs(5773)) xor (layer0_outputs(1203)));
    outputs(7593) <= (layer0_outputs(760)) or (layer0_outputs(5030));
    outputs(7594) <= not((layer0_outputs(4161)) xor (layer0_outputs(386)));
    outputs(7595) <= not(layer0_outputs(3025));
    outputs(7596) <= not(layer0_outputs(4307));
    outputs(7597) <= layer0_outputs(210);
    outputs(7598) <= (layer0_outputs(5208)) and not (layer0_outputs(90));
    outputs(7599) <= not((layer0_outputs(2258)) or (layer0_outputs(2508)));
    outputs(7600) <= layer0_outputs(4819);
    outputs(7601) <= layer0_outputs(7273);
    outputs(7602) <= not((layer0_outputs(2455)) or (layer0_outputs(6488)));
    outputs(7603) <= layer0_outputs(862);
    outputs(7604) <= layer0_outputs(1405);
    outputs(7605) <= not((layer0_outputs(565)) or (layer0_outputs(6875)));
    outputs(7606) <= not(layer0_outputs(769));
    outputs(7607) <= (layer0_outputs(7461)) and not (layer0_outputs(3329));
    outputs(7608) <= layer0_outputs(4844);
    outputs(7609) <= (layer0_outputs(1987)) and not (layer0_outputs(190));
    outputs(7610) <= (layer0_outputs(1564)) and not (layer0_outputs(608));
    outputs(7611) <= not(layer0_outputs(1174));
    outputs(7612) <= not(layer0_outputs(6030)) or (layer0_outputs(7613));
    outputs(7613) <= not(layer0_outputs(7597));
    outputs(7614) <= layer0_outputs(7156);
    outputs(7615) <= (layer0_outputs(3571)) xor (layer0_outputs(1062));
    outputs(7616) <= layer0_outputs(5667);
    outputs(7617) <= (layer0_outputs(2032)) and not (layer0_outputs(5045));
    outputs(7618) <= (layer0_outputs(2995)) and not (layer0_outputs(5707));
    outputs(7619) <= layer0_outputs(23);
    outputs(7620) <= (layer0_outputs(3419)) and (layer0_outputs(4925));
    outputs(7621) <= not(layer0_outputs(6491)) or (layer0_outputs(6632));
    outputs(7622) <= layer0_outputs(2718);
    outputs(7623) <= (layer0_outputs(6371)) and not (layer0_outputs(7623));
    outputs(7624) <= (layer0_outputs(217)) and not (layer0_outputs(5417));
    outputs(7625) <= layer0_outputs(2247);
    outputs(7626) <= not((layer0_outputs(1754)) or (layer0_outputs(1351)));
    outputs(7627) <= (layer0_outputs(53)) xor (layer0_outputs(3057));
    outputs(7628) <= (layer0_outputs(7551)) and (layer0_outputs(2210));
    outputs(7629) <= not(layer0_outputs(87));
    outputs(7630) <= layer0_outputs(642);
    outputs(7631) <= layer0_outputs(5792);
    outputs(7632) <= not(layer0_outputs(4606));
    outputs(7633) <= (layer0_outputs(1276)) xor (layer0_outputs(5700));
    outputs(7634) <= not(layer0_outputs(6440));
    outputs(7635) <= layer0_outputs(5661);
    outputs(7636) <= (layer0_outputs(7506)) and not (layer0_outputs(1006));
    outputs(7637) <= layer0_outputs(2938);
    outputs(7638) <= not(layer0_outputs(3901));
    outputs(7639) <= not((layer0_outputs(4891)) or (layer0_outputs(6514)));
    outputs(7640) <= not(layer0_outputs(610)) or (layer0_outputs(4692));
    outputs(7641) <= layer0_outputs(6492);
    outputs(7642) <= layer0_outputs(2077);
    outputs(7643) <= layer0_outputs(423);
    outputs(7644) <= layer0_outputs(5625);
    outputs(7645) <= (layer0_outputs(4496)) and (layer0_outputs(6469));
    outputs(7646) <= (layer0_outputs(2456)) xor (layer0_outputs(1252));
    outputs(7647) <= not((layer0_outputs(6045)) xor (layer0_outputs(6717)));
    outputs(7648) <= (layer0_outputs(5743)) and not (layer0_outputs(3518));
    outputs(7649) <= layer0_outputs(1009);
    outputs(7650) <= layer0_outputs(6171);
    outputs(7651) <= not(layer0_outputs(2351));
    outputs(7652) <= not(layer0_outputs(1371)) or (layer0_outputs(1859));
    outputs(7653) <= not(layer0_outputs(3941));
    outputs(7654) <= not(layer0_outputs(2240));
    outputs(7655) <= (layer0_outputs(5402)) and not (layer0_outputs(455));
    outputs(7656) <= not(layer0_outputs(2090));
    outputs(7657) <= (layer0_outputs(3294)) and not (layer0_outputs(1328));
    outputs(7658) <= not(layer0_outputs(6572));
    outputs(7659) <= not(layer0_outputs(6696));
    outputs(7660) <= layer0_outputs(103);
    outputs(7661) <= (layer0_outputs(5885)) xor (layer0_outputs(5953));
    outputs(7662) <= not(layer0_outputs(2391));
    outputs(7663) <= not((layer0_outputs(6948)) xor (layer0_outputs(2170)));
    outputs(7664) <= layer0_outputs(6954);
    outputs(7665) <= (layer0_outputs(5298)) and not (layer0_outputs(3191));
    outputs(7666) <= (layer0_outputs(1245)) or (layer0_outputs(3176));
    outputs(7667) <= (layer0_outputs(4895)) and not (layer0_outputs(507));
    outputs(7668) <= (layer0_outputs(7313)) or (layer0_outputs(1368));
    outputs(7669) <= not((layer0_outputs(6981)) or (layer0_outputs(7568)));
    outputs(7670) <= (layer0_outputs(515)) and (layer0_outputs(5419));
    outputs(7671) <= not((layer0_outputs(5309)) or (layer0_outputs(901)));
    outputs(7672) <= not(layer0_outputs(6562));
    outputs(7673) <= not(layer0_outputs(5237));
    outputs(7674) <= (layer0_outputs(5142)) xor (layer0_outputs(6420));
    outputs(7675) <= layer0_outputs(3586);
    outputs(7676) <= (layer0_outputs(2519)) and (layer0_outputs(3436));
    outputs(7677) <= (layer0_outputs(7128)) and not (layer0_outputs(5127));
    outputs(7678) <= layer0_outputs(6415);
    outputs(7679) <= (layer0_outputs(4267)) and not (layer0_outputs(4534));

end Behavioral;
