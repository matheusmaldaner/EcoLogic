library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(2559 downto 0);
    signal layer1_outputs: std_logic_vector(2559 downto 0);
    signal layer2_outputs: std_logic_vector(2559 downto 0);
    signal layer3_outputs: std_logic_vector(2559 downto 0);
    signal layer4_outputs: std_logic_vector(2559 downto 0);

begin
    layer0_outputs(0) <= a or b;
    layer0_outputs(1) <= a and not b;
    layer0_outputs(2) <= a and not b;
    layer0_outputs(3) <= a and not b;
    layer0_outputs(4) <= a and not b;
    layer0_outputs(5) <= b;
    layer0_outputs(6) <= a or b;
    layer0_outputs(7) <= a xor b;
    layer0_outputs(8) <= not (a or b);
    layer0_outputs(9) <= a or b;
    layer0_outputs(10) <= a or b;
    layer0_outputs(11) <= not a;
    layer0_outputs(12) <= not a or b;
    layer0_outputs(13) <= a or b;
    layer0_outputs(14) <= 1'b1;
    layer0_outputs(15) <= not (a and b);
    layer0_outputs(16) <= 1'b0;
    layer0_outputs(17) <= not a;
    layer0_outputs(18) <= not b or a;
    layer0_outputs(19) <= not b or a;
    layer0_outputs(20) <= a or b;
    layer0_outputs(21) <= not (a or b);
    layer0_outputs(22) <= not b;
    layer0_outputs(23) <= not (a xor b);
    layer0_outputs(24) <= not a;
    layer0_outputs(25) <= not a or b;
    layer0_outputs(26) <= b and not a;
    layer0_outputs(27) <= a and not b;
    layer0_outputs(28) <= a and not b;
    layer0_outputs(29) <= a or b;
    layer0_outputs(30) <= 1'b1;
    layer0_outputs(31) <= not b or a;
    layer0_outputs(32) <= not a;
    layer0_outputs(33) <= not (a xor b);
    layer0_outputs(34) <= a or b;
    layer0_outputs(35) <= a and b;
    layer0_outputs(36) <= not a or b;
    layer0_outputs(37) <= not (a xor b);
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= a;
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= 1'b1;
    layer0_outputs(42) <= 1'b0;
    layer0_outputs(43) <= a and not b;
    layer0_outputs(44) <= a and not b;
    layer0_outputs(45) <= not a or b;
    layer0_outputs(46) <= 1'b1;
    layer0_outputs(47) <= a or b;
    layer0_outputs(48) <= b;
    layer0_outputs(49) <= a;
    layer0_outputs(50) <= a;
    layer0_outputs(51) <= not a;
    layer0_outputs(52) <= not a or b;
    layer0_outputs(53) <= not b or a;
    layer0_outputs(54) <= not (a or b);
    layer0_outputs(55) <= a or b;
    layer0_outputs(56) <= not b;
    layer0_outputs(57) <= 1'b1;
    layer0_outputs(58) <= 1'b0;
    layer0_outputs(59) <= not (a and b);
    layer0_outputs(60) <= not a;
    layer0_outputs(61) <= a or b;
    layer0_outputs(62) <= a and b;
    layer0_outputs(63) <= b and not a;
    layer0_outputs(64) <= not b or a;
    layer0_outputs(65) <= not b or a;
    layer0_outputs(66) <= 1'b1;
    layer0_outputs(67) <= b;
    layer0_outputs(68) <= not (a or b);
    layer0_outputs(69) <= not a or b;
    layer0_outputs(70) <= a and b;
    layer0_outputs(71) <= not b;
    layer0_outputs(72) <= b;
    layer0_outputs(73) <= not (a xor b);
    layer0_outputs(74) <= b and not a;
    layer0_outputs(75) <= a or b;
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= a and not b;
    layer0_outputs(78) <= a;
    layer0_outputs(79) <= a;
    layer0_outputs(80) <= not a or b;
    layer0_outputs(81) <= not (a or b);
    layer0_outputs(82) <= not (a xor b);
    layer0_outputs(83) <= not (a or b);
    layer0_outputs(84) <= not b;
    layer0_outputs(85) <= a;
    layer0_outputs(86) <= not (a xor b);
    layer0_outputs(87) <= not b;
    layer0_outputs(88) <= a or b;
    layer0_outputs(89) <= not (a or b);
    layer0_outputs(90) <= not a;
    layer0_outputs(91) <= a or b;
    layer0_outputs(92) <= 1'b1;
    layer0_outputs(93) <= not b or a;
    layer0_outputs(94) <= a and not b;
    layer0_outputs(95) <= not (a and b);
    layer0_outputs(96) <= b;
    layer0_outputs(97) <= 1'b1;
    layer0_outputs(98) <= a;
    layer0_outputs(99) <= 1'b1;
    layer0_outputs(100) <= not (a xor b);
    layer0_outputs(101) <= a and not b;
    layer0_outputs(102) <= not a;
    layer0_outputs(103) <= a xor b;
    layer0_outputs(104) <= not a or b;
    layer0_outputs(105) <= b;
    layer0_outputs(106) <= b and not a;
    layer0_outputs(107) <= not (a or b);
    layer0_outputs(108) <= a;
    layer0_outputs(109) <= b;
    layer0_outputs(110) <= a and b;
    layer0_outputs(111) <= a xor b;
    layer0_outputs(112) <= b and not a;
    layer0_outputs(113) <= 1'b1;
    layer0_outputs(114) <= not a;
    layer0_outputs(115) <= b and not a;
    layer0_outputs(116) <= not (a or b);
    layer0_outputs(117) <= not b;
    layer0_outputs(118) <= a;
    layer0_outputs(119) <= not (a or b);
    layer0_outputs(120) <= a xor b;
    layer0_outputs(121) <= b;
    layer0_outputs(122) <= not b or a;
    layer0_outputs(123) <= a;
    layer0_outputs(124) <= not b;
    layer0_outputs(125) <= not (a xor b);
    layer0_outputs(126) <= 1'b1;
    layer0_outputs(127) <= b and not a;
    layer0_outputs(128) <= a and b;
    layer0_outputs(129) <= 1'b0;
    layer0_outputs(130) <= not b;
    layer0_outputs(131) <= a and not b;
    layer0_outputs(132) <= a;
    layer0_outputs(133) <= b and not a;
    layer0_outputs(134) <= not b;
    layer0_outputs(135) <= b and not a;
    layer0_outputs(136) <= not (a or b);
    layer0_outputs(137) <= b and not a;
    layer0_outputs(138) <= not (a xor b);
    layer0_outputs(139) <= not b;
    layer0_outputs(140) <= not (a and b);
    layer0_outputs(141) <= b;
    layer0_outputs(142) <= a;
    layer0_outputs(143) <= a;
    layer0_outputs(144) <= a or b;
    layer0_outputs(145) <= not a or b;
    layer0_outputs(146) <= b and not a;
    layer0_outputs(147) <= not b or a;
    layer0_outputs(148) <= not b;
    layer0_outputs(149) <= not a;
    layer0_outputs(150) <= a;
    layer0_outputs(151) <= not a or b;
    layer0_outputs(152) <= not a;
    layer0_outputs(153) <= a;
    layer0_outputs(154) <= a xor b;
    layer0_outputs(155) <= a or b;
    layer0_outputs(156) <= a;
    layer0_outputs(157) <= a xor b;
    layer0_outputs(158) <= a or b;
    layer0_outputs(159) <= b;
    layer0_outputs(160) <= b and not a;
    layer0_outputs(161) <= not a;
    layer0_outputs(162) <= a;
    layer0_outputs(163) <= a or b;
    layer0_outputs(164) <= not a;
    layer0_outputs(165) <= 1'b1;
    layer0_outputs(166) <= a xor b;
    layer0_outputs(167) <= not b or a;
    layer0_outputs(168) <= 1'b1;
    layer0_outputs(169) <= not (a and b);
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= not a;
    layer0_outputs(172) <= not a;
    layer0_outputs(173) <= not (a or b);
    layer0_outputs(174) <= not (a and b);
    layer0_outputs(175) <= a;
    layer0_outputs(176) <= b and not a;
    layer0_outputs(177) <= 1'b0;
    layer0_outputs(178) <= not (a or b);
    layer0_outputs(179) <= a and b;
    layer0_outputs(180) <= b;
    layer0_outputs(181) <= b;
    layer0_outputs(182) <= 1'b0;
    layer0_outputs(183) <= not (a or b);
    layer0_outputs(184) <= a;
    layer0_outputs(185) <= a and not b;
    layer0_outputs(186) <= a and b;
    layer0_outputs(187) <= not (a or b);
    layer0_outputs(188) <= a or b;
    layer0_outputs(189) <= not (a xor b);
    layer0_outputs(190) <= a;
    layer0_outputs(191) <= not (a or b);
    layer0_outputs(192) <= not a;
    layer0_outputs(193) <= a or b;
    layer0_outputs(194) <= not b;
    layer0_outputs(195) <= not a;
    layer0_outputs(196) <= 1'b0;
    layer0_outputs(197) <= a and not b;
    layer0_outputs(198) <= 1'b1;
    layer0_outputs(199) <= a and b;
    layer0_outputs(200) <= not (a xor b);
    layer0_outputs(201) <= a or b;
    layer0_outputs(202) <= not (a or b);
    layer0_outputs(203) <= b;
    layer0_outputs(204) <= not b;
    layer0_outputs(205) <= not b or a;
    layer0_outputs(206) <= a;
    layer0_outputs(207) <= a and b;
    layer0_outputs(208) <= not a or b;
    layer0_outputs(209) <= a or b;
    layer0_outputs(210) <= 1'b1;
    layer0_outputs(211) <= not (a xor b);
    layer0_outputs(212) <= a or b;
    layer0_outputs(213) <= a or b;
    layer0_outputs(214) <= a or b;
    layer0_outputs(215) <= b;
    layer0_outputs(216) <= not a or b;
    layer0_outputs(217) <= a;
    layer0_outputs(218) <= not b or a;
    layer0_outputs(219) <= not (a or b);
    layer0_outputs(220) <= not (a xor b);
    layer0_outputs(221) <= not b;
    layer0_outputs(222) <= b;
    layer0_outputs(223) <= b and not a;
    layer0_outputs(224) <= not a or b;
    layer0_outputs(225) <= not b;
    layer0_outputs(226) <= not (a or b);
    layer0_outputs(227) <= not a;
    layer0_outputs(228) <= b and not a;
    layer0_outputs(229) <= a;
    layer0_outputs(230) <= not a;
    layer0_outputs(231) <= b;
    layer0_outputs(232) <= not b or a;
    layer0_outputs(233) <= not (a xor b);
    layer0_outputs(234) <= not b or a;
    layer0_outputs(235) <= 1'b0;
    layer0_outputs(236) <= not (a xor b);
    layer0_outputs(237) <= not (a or b);
    layer0_outputs(238) <= a;
    layer0_outputs(239) <= 1'b0;
    layer0_outputs(240) <= b;
    layer0_outputs(241) <= not a or b;
    layer0_outputs(242) <= 1'b1;
    layer0_outputs(243) <= a;
    layer0_outputs(244) <= b and not a;
    layer0_outputs(245) <= 1'b1;
    layer0_outputs(246) <= not b or a;
    layer0_outputs(247) <= b and not a;
    layer0_outputs(248) <= b;
    layer0_outputs(249) <= not b;
    layer0_outputs(250) <= b and not a;
    layer0_outputs(251) <= not (a or b);
    layer0_outputs(252) <= 1'b1;
    layer0_outputs(253) <= a and not b;
    layer0_outputs(254) <= not b;
    layer0_outputs(255) <= not (a and b);
    layer0_outputs(256) <= not (a or b);
    layer0_outputs(257) <= not (a or b);
    layer0_outputs(258) <= a xor b;
    layer0_outputs(259) <= not b or a;
    layer0_outputs(260) <= not (a or b);
    layer0_outputs(261) <= not (a or b);
    layer0_outputs(262) <= b;
    layer0_outputs(263) <= not a;
    layer0_outputs(264) <= not (a xor b);
    layer0_outputs(265) <= not (a xor b);
    layer0_outputs(266) <= 1'b1;
    layer0_outputs(267) <= not a;
    layer0_outputs(268) <= 1'b0;
    layer0_outputs(269) <= not a;
    layer0_outputs(270) <= a or b;
    layer0_outputs(271) <= 1'b1;
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= a xor b;
    layer0_outputs(274) <= b;
    layer0_outputs(275) <= not a;
    layer0_outputs(276) <= 1'b1;
    layer0_outputs(277) <= b;
    layer0_outputs(278) <= a or b;
    layer0_outputs(279) <= not (a or b);
    layer0_outputs(280) <= not b or a;
    layer0_outputs(281) <= a or b;
    layer0_outputs(282) <= not a or b;
    layer0_outputs(283) <= not b;
    layer0_outputs(284) <= a and b;
    layer0_outputs(285) <= b and not a;
    layer0_outputs(286) <= a and not b;
    layer0_outputs(287) <= a or b;
    layer0_outputs(288) <= a;
    layer0_outputs(289) <= not (a and b);
    layer0_outputs(290) <= 1'b1;
    layer0_outputs(291) <= not a or b;
    layer0_outputs(292) <= not a or b;
    layer0_outputs(293) <= a and not b;
    layer0_outputs(294) <= b;
    layer0_outputs(295) <= not a or b;
    layer0_outputs(296) <= a and not b;
    layer0_outputs(297) <= a and not b;
    layer0_outputs(298) <= a and not b;
    layer0_outputs(299) <= a and not b;
    layer0_outputs(300) <= not a or b;
    layer0_outputs(301) <= not a;
    layer0_outputs(302) <= a;
    layer0_outputs(303) <= 1'b1;
    layer0_outputs(304) <= a or b;
    layer0_outputs(305) <= a;
    layer0_outputs(306) <= a;
    layer0_outputs(307) <= a or b;
    layer0_outputs(308) <= b;
    layer0_outputs(309) <= not (a and b);
    layer0_outputs(310) <= not (a or b);
    layer0_outputs(311) <= a or b;
    layer0_outputs(312) <= a and b;
    layer0_outputs(313) <= a or b;
    layer0_outputs(314) <= not b or a;
    layer0_outputs(315) <= not b;
    layer0_outputs(316) <= b;
    layer0_outputs(317) <= not a;
    layer0_outputs(318) <= a or b;
    layer0_outputs(319) <= b;
    layer0_outputs(320) <= b;
    layer0_outputs(321) <= a;
    layer0_outputs(322) <= b;
    layer0_outputs(323) <= not a or b;
    layer0_outputs(324) <= not a;
    layer0_outputs(325) <= b;
    layer0_outputs(326) <= not b or a;
    layer0_outputs(327) <= not (a or b);
    layer0_outputs(328) <= a or b;
    layer0_outputs(329) <= not a or b;
    layer0_outputs(330) <= a;
    layer0_outputs(331) <= b;
    layer0_outputs(332) <= not b;
    layer0_outputs(333) <= not b;
    layer0_outputs(334) <= not b;
    layer0_outputs(335) <= a and b;
    layer0_outputs(336) <= not (a or b);
    layer0_outputs(337) <= a or b;
    layer0_outputs(338) <= b;
    layer0_outputs(339) <= 1'b1;
    layer0_outputs(340) <= not (a xor b);
    layer0_outputs(341) <= not a or b;
    layer0_outputs(342) <= b and not a;
    layer0_outputs(343) <= b and not a;
    layer0_outputs(344) <= a or b;
    layer0_outputs(345) <= b and not a;
    layer0_outputs(346) <= a and not b;
    layer0_outputs(347) <= a or b;
    layer0_outputs(348) <= not a;
    layer0_outputs(349) <= not (a and b);
    layer0_outputs(350) <= not (a or b);
    layer0_outputs(351) <= not b;
    layer0_outputs(352) <= not a or b;
    layer0_outputs(353) <= b;
    layer0_outputs(354) <= not (a or b);
    layer0_outputs(355) <= not a or b;
    layer0_outputs(356) <= not (a or b);
    layer0_outputs(357) <= a;
    layer0_outputs(358) <= not (a or b);
    layer0_outputs(359) <= not a;
    layer0_outputs(360) <= not (a or b);
    layer0_outputs(361) <= a or b;
    layer0_outputs(362) <= b;
    layer0_outputs(363) <= a or b;
    layer0_outputs(364) <= a or b;
    layer0_outputs(365) <= not a;
    layer0_outputs(366) <= a and b;
    layer0_outputs(367) <= not b;
    layer0_outputs(368) <= not a or b;
    layer0_outputs(369) <= not a;
    layer0_outputs(370) <= not (a or b);
    layer0_outputs(371) <= a and not b;
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= a or b;
    layer0_outputs(374) <= a and not b;
    layer0_outputs(375) <= not b;
    layer0_outputs(376) <= a;
    layer0_outputs(377) <= a or b;
    layer0_outputs(378) <= not b or a;
    layer0_outputs(379) <= not (a or b);
    layer0_outputs(380) <= a;
    layer0_outputs(381) <= a or b;
    layer0_outputs(382) <= a or b;
    layer0_outputs(383) <= not (a and b);
    layer0_outputs(384) <= not (a or b);
    layer0_outputs(385) <= not a;
    layer0_outputs(386) <= not (a xor b);
    layer0_outputs(387) <= 1'b1;
    layer0_outputs(388) <= b and not a;
    layer0_outputs(389) <= not b;
    layer0_outputs(390) <= not b;
    layer0_outputs(391) <= a or b;
    layer0_outputs(392) <= a or b;
    layer0_outputs(393) <= b and not a;
    layer0_outputs(394) <= a and not b;
    layer0_outputs(395) <= a or b;
    layer0_outputs(396) <= not (a xor b);
    layer0_outputs(397) <= a and not b;
    layer0_outputs(398) <= b and not a;
    layer0_outputs(399) <= not b;
    layer0_outputs(400) <= not (a or b);
    layer0_outputs(401) <= not (a and b);
    layer0_outputs(402) <= not b;
    layer0_outputs(403) <= not (a and b);
    layer0_outputs(404) <= b and not a;
    layer0_outputs(405) <= 1'b1;
    layer0_outputs(406) <= b and not a;
    layer0_outputs(407) <= a and b;
    layer0_outputs(408) <= not (a or b);
    layer0_outputs(409) <= 1'b1;
    layer0_outputs(410) <= b;
    layer0_outputs(411) <= b;
    layer0_outputs(412) <= a xor b;
    layer0_outputs(413) <= b;
    layer0_outputs(414) <= a and not b;
    layer0_outputs(415) <= not (a xor b);
    layer0_outputs(416) <= not a or b;
    layer0_outputs(417) <= not b;
    layer0_outputs(418) <= a and not b;
    layer0_outputs(419) <= a and b;
    layer0_outputs(420) <= not a or b;
    layer0_outputs(421) <= b;
    layer0_outputs(422) <= not b or a;
    layer0_outputs(423) <= not a or b;
    layer0_outputs(424) <= not (a xor b);
    layer0_outputs(425) <= a and not b;
    layer0_outputs(426) <= b and not a;
    layer0_outputs(427) <= a or b;
    layer0_outputs(428) <= not b or a;
    layer0_outputs(429) <= b and not a;
    layer0_outputs(430) <= a and not b;
    layer0_outputs(431) <= 1'b1;
    layer0_outputs(432) <= a and b;
    layer0_outputs(433) <= not b or a;
    layer0_outputs(434) <= not (a xor b);
    layer0_outputs(435) <= not b;
    layer0_outputs(436) <= a or b;
    layer0_outputs(437) <= a;
    layer0_outputs(438) <= a or b;
    layer0_outputs(439) <= a and not b;
    layer0_outputs(440) <= b and not a;
    layer0_outputs(441) <= not (a or b);
    layer0_outputs(442) <= a xor b;
    layer0_outputs(443) <= not b;
    layer0_outputs(444) <= a;
    layer0_outputs(445) <= 1'b1;
    layer0_outputs(446) <= not b;
    layer0_outputs(447) <= not a or b;
    layer0_outputs(448) <= a;
    layer0_outputs(449) <= 1'b1;
    layer0_outputs(450) <= not b;
    layer0_outputs(451) <= 1'b1;
    layer0_outputs(452) <= 1'b0;
    layer0_outputs(453) <= a;
    layer0_outputs(454) <= b;
    layer0_outputs(455) <= b and not a;
    layer0_outputs(456) <= not a or b;
    layer0_outputs(457) <= a xor b;
    layer0_outputs(458) <= not a;
    layer0_outputs(459) <= b;
    layer0_outputs(460) <= b;
    layer0_outputs(461) <= not a;
    layer0_outputs(462) <= not (a or b);
    layer0_outputs(463) <= 1'b1;
    layer0_outputs(464) <= not b;
    layer0_outputs(465) <= b;
    layer0_outputs(466) <= a xor b;
    layer0_outputs(467) <= a and not b;
    layer0_outputs(468) <= b and not a;
    layer0_outputs(469) <= 1'b0;
    layer0_outputs(470) <= b;
    layer0_outputs(471) <= 1'b0;
    layer0_outputs(472) <= not a;
    layer0_outputs(473) <= not (a or b);
    layer0_outputs(474) <= b and not a;
    layer0_outputs(475) <= a or b;
    layer0_outputs(476) <= not (a or b);
    layer0_outputs(477) <= not b;
    layer0_outputs(478) <= a xor b;
    layer0_outputs(479) <= not (a or b);
    layer0_outputs(480) <= 1'b1;
    layer0_outputs(481) <= not b;
    layer0_outputs(482) <= not b or a;
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= a;
    layer0_outputs(485) <= b;
    layer0_outputs(486) <= not (a or b);
    layer0_outputs(487) <= not (a or b);
    layer0_outputs(488) <= a or b;
    layer0_outputs(489) <= a and b;
    layer0_outputs(490) <= not (a or b);
    layer0_outputs(491) <= a and not b;
    layer0_outputs(492) <= not (a xor b);
    layer0_outputs(493) <= a or b;
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= not a;
    layer0_outputs(496) <= not (a or b);
    layer0_outputs(497) <= not (a and b);
    layer0_outputs(498) <= 1'b0;
    layer0_outputs(499) <= a and not b;
    layer0_outputs(500) <= b and not a;
    layer0_outputs(501) <= a or b;
    layer0_outputs(502) <= 1'b1;
    layer0_outputs(503) <= a and b;
    layer0_outputs(504) <= a;
    layer0_outputs(505) <= not a or b;
    layer0_outputs(506) <= a xor b;
    layer0_outputs(507) <= 1'b1;
    layer0_outputs(508) <= a xor b;
    layer0_outputs(509) <= not b or a;
    layer0_outputs(510) <= not a;
    layer0_outputs(511) <= not b;
    layer0_outputs(512) <= not a or b;
    layer0_outputs(513) <= b;
    layer0_outputs(514) <= a xor b;
    layer0_outputs(515) <= a xor b;
    layer0_outputs(516) <= not a or b;
    layer0_outputs(517) <= not a;
    layer0_outputs(518) <= 1'b0;
    layer0_outputs(519) <= a and not b;
    layer0_outputs(520) <= a xor b;
    layer0_outputs(521) <= not a;
    layer0_outputs(522) <= not (a xor b);
    layer0_outputs(523) <= not (a xor b);
    layer0_outputs(524) <= a and b;
    layer0_outputs(525) <= not (a or b);
    layer0_outputs(526) <= a and b;
    layer0_outputs(527) <= a;
    layer0_outputs(528) <= a and b;
    layer0_outputs(529) <= not b;
    layer0_outputs(530) <= a and b;
    layer0_outputs(531) <= not a;
    layer0_outputs(532) <= not a or b;
    layer0_outputs(533) <= 1'b1;
    layer0_outputs(534) <= a or b;
    layer0_outputs(535) <= b;
    layer0_outputs(536) <= 1'b0;
    layer0_outputs(537) <= a and not b;
    layer0_outputs(538) <= a and not b;
    layer0_outputs(539) <= not (a or b);
    layer0_outputs(540) <= a;
    layer0_outputs(541) <= not b or a;
    layer0_outputs(542) <= not (a or b);
    layer0_outputs(543) <= b;
    layer0_outputs(544) <= a;
    layer0_outputs(545) <= a xor b;
    layer0_outputs(546) <= a and b;
    layer0_outputs(547) <= not (a or b);
    layer0_outputs(548) <= b;
    layer0_outputs(549) <= not a;
    layer0_outputs(550) <= a or b;
    layer0_outputs(551) <= a;
    layer0_outputs(552) <= a;
    layer0_outputs(553) <= a and b;
    layer0_outputs(554) <= not b;
    layer0_outputs(555) <= not (a or b);
    layer0_outputs(556) <= not b;
    layer0_outputs(557) <= not a;
    layer0_outputs(558) <= a;
    layer0_outputs(559) <= not (a xor b);
    layer0_outputs(560) <= a and not b;
    layer0_outputs(561) <= a xor b;
    layer0_outputs(562) <= b and not a;
    layer0_outputs(563) <= b;
    layer0_outputs(564) <= not a or b;
    layer0_outputs(565) <= not b;
    layer0_outputs(566) <= not (a and b);
    layer0_outputs(567) <= not a;
    layer0_outputs(568) <= a and not b;
    layer0_outputs(569) <= 1'b0;
    layer0_outputs(570) <= not a;
    layer0_outputs(571) <= not a;
    layer0_outputs(572) <= not (a and b);
    layer0_outputs(573) <= a;
    layer0_outputs(574) <= not a or b;
    layer0_outputs(575) <= not a;
    layer0_outputs(576) <= not a or b;
    layer0_outputs(577) <= not a;
    layer0_outputs(578) <= not b;
    layer0_outputs(579) <= not (a xor b);
    layer0_outputs(580) <= a xor b;
    layer0_outputs(581) <= a or b;
    layer0_outputs(582) <= a and not b;
    layer0_outputs(583) <= not b or a;
    layer0_outputs(584) <= b and not a;
    layer0_outputs(585) <= a or b;
    layer0_outputs(586) <= a and not b;
    layer0_outputs(587) <= not b;
    layer0_outputs(588) <= 1'b0;
    layer0_outputs(589) <= a xor b;
    layer0_outputs(590) <= not (a xor b);
    layer0_outputs(591) <= not b;
    layer0_outputs(592) <= a;
    layer0_outputs(593) <= not (a xor b);
    layer0_outputs(594) <= not (a and b);
    layer0_outputs(595) <= not (a and b);
    layer0_outputs(596) <= not (a xor b);
    layer0_outputs(597) <= not a;
    layer0_outputs(598) <= 1'b0;
    layer0_outputs(599) <= a;
    layer0_outputs(600) <= a or b;
    layer0_outputs(601) <= not (a or b);
    layer0_outputs(602) <= not (a or b);
    layer0_outputs(603) <= b;
    layer0_outputs(604) <= a xor b;
    layer0_outputs(605) <= not a;
    layer0_outputs(606) <= not a or b;
    layer0_outputs(607) <= not b or a;
    layer0_outputs(608) <= not b;
    layer0_outputs(609) <= a and not b;
    layer0_outputs(610) <= a;
    layer0_outputs(611) <= not (a or b);
    layer0_outputs(612) <= not b;
    layer0_outputs(613) <= a;
    layer0_outputs(614) <= a and b;
    layer0_outputs(615) <= not b or a;
    layer0_outputs(616) <= a or b;
    layer0_outputs(617) <= not a;
    layer0_outputs(618) <= 1'b1;
    layer0_outputs(619) <= b and not a;
    layer0_outputs(620) <= a and not b;
    layer0_outputs(621) <= a;
    layer0_outputs(622) <= b;
    layer0_outputs(623) <= not (a or b);
    layer0_outputs(624) <= b and not a;
    layer0_outputs(625) <= not (a xor b);
    layer0_outputs(626) <= a or b;
    layer0_outputs(627) <= b;
    layer0_outputs(628) <= not a or b;
    layer0_outputs(629) <= 1'b0;
    layer0_outputs(630) <= b and not a;
    layer0_outputs(631) <= b;
    layer0_outputs(632) <= not b or a;
    layer0_outputs(633) <= not a;
    layer0_outputs(634) <= b and not a;
    layer0_outputs(635) <= 1'b1;
    layer0_outputs(636) <= not b;
    layer0_outputs(637) <= not b or a;
    layer0_outputs(638) <= not (a or b);
    layer0_outputs(639) <= a;
    layer0_outputs(640) <= b and not a;
    layer0_outputs(641) <= a and not b;
    layer0_outputs(642) <= not (a or b);
    layer0_outputs(643) <= a or b;
    layer0_outputs(644) <= not (a or b);
    layer0_outputs(645) <= not (a xor b);
    layer0_outputs(646) <= b;
    layer0_outputs(647) <= a and not b;
    layer0_outputs(648) <= not a or b;
    layer0_outputs(649) <= not (a or b);
    layer0_outputs(650) <= not a;
    layer0_outputs(651) <= a and not b;
    layer0_outputs(652) <= b and not a;
    layer0_outputs(653) <= not (a or b);
    layer0_outputs(654) <= not a or b;
    layer0_outputs(655) <= not b;
    layer0_outputs(656) <= not b;
    layer0_outputs(657) <= b and not a;
    layer0_outputs(658) <= not a or b;
    layer0_outputs(659) <= not a;
    layer0_outputs(660) <= not (a and b);
    layer0_outputs(661) <= a;
    layer0_outputs(662) <= not b;
    layer0_outputs(663) <= not b or a;
    layer0_outputs(664) <= not (a xor b);
    layer0_outputs(665) <= not (a xor b);
    layer0_outputs(666) <= not a;
    layer0_outputs(667) <= 1'b0;
    layer0_outputs(668) <= not (a or b);
    layer0_outputs(669) <= not (a or b);
    layer0_outputs(670) <= not (a and b);
    layer0_outputs(671) <= not b;
    layer0_outputs(672) <= not b;
    layer0_outputs(673) <= a and not b;
    layer0_outputs(674) <= b;
    layer0_outputs(675) <= a or b;
    layer0_outputs(676) <= a;
    layer0_outputs(677) <= not (a or b);
    layer0_outputs(678) <= a or b;
    layer0_outputs(679) <= a or b;
    layer0_outputs(680) <= a and b;
    layer0_outputs(681) <= not b;
    layer0_outputs(682) <= not (a xor b);
    layer0_outputs(683) <= not b or a;
    layer0_outputs(684) <= a or b;
    layer0_outputs(685) <= not a or b;
    layer0_outputs(686) <= not (a and b);
    layer0_outputs(687) <= not (a xor b);
    layer0_outputs(688) <= not b;
    layer0_outputs(689) <= a and b;
    layer0_outputs(690) <= not (a or b);
    layer0_outputs(691) <= not (a or b);
    layer0_outputs(692) <= not (a or b);
    layer0_outputs(693) <= a xor b;
    layer0_outputs(694) <= not a or b;
    layer0_outputs(695) <= not (a xor b);
    layer0_outputs(696) <= a xor b;
    layer0_outputs(697) <= a xor b;
    layer0_outputs(698) <= not a;
    layer0_outputs(699) <= b;
    layer0_outputs(700) <= not b;
    layer0_outputs(701) <= not a or b;
    layer0_outputs(702) <= not b or a;
    layer0_outputs(703) <= a;
    layer0_outputs(704) <= b;
    layer0_outputs(705) <= 1'b0;
    layer0_outputs(706) <= b;
    layer0_outputs(707) <= b;
    layer0_outputs(708) <= a and b;
    layer0_outputs(709) <= not (a or b);
    layer0_outputs(710) <= not (a or b);
    layer0_outputs(711) <= a xor b;
    layer0_outputs(712) <= not a;
    layer0_outputs(713) <= 1'b0;
    layer0_outputs(714) <= not (a xor b);
    layer0_outputs(715) <= b;
    layer0_outputs(716) <= a and b;
    layer0_outputs(717) <= not b or a;
    layer0_outputs(718) <= a;
    layer0_outputs(719) <= not (a xor b);
    layer0_outputs(720) <= 1'b1;
    layer0_outputs(721) <= not (a or b);
    layer0_outputs(722) <= a;
    layer0_outputs(723) <= not a or b;
    layer0_outputs(724) <= not a;
    layer0_outputs(725) <= b;
    layer0_outputs(726) <= not (a xor b);
    layer0_outputs(727) <= b and not a;
    layer0_outputs(728) <= not b or a;
    layer0_outputs(729) <= a and not b;
    layer0_outputs(730) <= not (a and b);
    layer0_outputs(731) <= not (a and b);
    layer0_outputs(732) <= not (a xor b);
    layer0_outputs(733) <= 1'b1;
    layer0_outputs(734) <= 1'b1;
    layer0_outputs(735) <= a;
    layer0_outputs(736) <= not b or a;
    layer0_outputs(737) <= not b or a;
    layer0_outputs(738) <= not (a xor b);
    layer0_outputs(739) <= a;
    layer0_outputs(740) <= not (a or b);
    layer0_outputs(741) <= a or b;
    layer0_outputs(742) <= not (a or b);
    layer0_outputs(743) <= a;
    layer0_outputs(744) <= 1'b1;
    layer0_outputs(745) <= not b;
    layer0_outputs(746) <= not a;
    layer0_outputs(747) <= a or b;
    layer0_outputs(748) <= a xor b;
    layer0_outputs(749) <= not a;
    layer0_outputs(750) <= not (a or b);
    layer0_outputs(751) <= not (a and b);
    layer0_outputs(752) <= a xor b;
    layer0_outputs(753) <= b;
    layer0_outputs(754) <= not (a or b);
    layer0_outputs(755) <= not (a and b);
    layer0_outputs(756) <= not (a xor b);
    layer0_outputs(757) <= not b;
    layer0_outputs(758) <= a and not b;
    layer0_outputs(759) <= not b;
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= a xor b;
    layer0_outputs(762) <= not b;
    layer0_outputs(763) <= not (a or b);
    layer0_outputs(764) <= 1'b0;
    layer0_outputs(765) <= not a or b;
    layer0_outputs(766) <= not (a or b);
    layer0_outputs(767) <= not b or a;
    layer0_outputs(768) <= a and b;
    layer0_outputs(769) <= not a or b;
    layer0_outputs(770) <= not b or a;
    layer0_outputs(771) <= not (a or b);
    layer0_outputs(772) <= a and not b;
    layer0_outputs(773) <= not a or b;
    layer0_outputs(774) <= not a or b;
    layer0_outputs(775) <= a or b;
    layer0_outputs(776) <= a;
    layer0_outputs(777) <= a or b;
    layer0_outputs(778) <= b and not a;
    layer0_outputs(779) <= not a or b;
    layer0_outputs(780) <= not b;
    layer0_outputs(781) <= not a;
    layer0_outputs(782) <= not b or a;
    layer0_outputs(783) <= a and b;
    layer0_outputs(784) <= a or b;
    layer0_outputs(785) <= a and not b;
    layer0_outputs(786) <= a;
    layer0_outputs(787) <= a;
    layer0_outputs(788) <= not a;
    layer0_outputs(789) <= not a;
    layer0_outputs(790) <= b and not a;
    layer0_outputs(791) <= b;
    layer0_outputs(792) <= not b;
    layer0_outputs(793) <= not b;
    layer0_outputs(794) <= not b or a;
    layer0_outputs(795) <= not a or b;
    layer0_outputs(796) <= a or b;
    layer0_outputs(797) <= not (a xor b);
    layer0_outputs(798) <= a xor b;
    layer0_outputs(799) <= not b;
    layer0_outputs(800) <= 1'b0;
    layer0_outputs(801) <= not a or b;
    layer0_outputs(802) <= a;
    layer0_outputs(803) <= b;
    layer0_outputs(804) <= a;
    layer0_outputs(805) <= a;
    layer0_outputs(806) <= a;
    layer0_outputs(807) <= a and b;
    layer0_outputs(808) <= not a;
    layer0_outputs(809) <= not a;
    layer0_outputs(810) <= not (a xor b);
    layer0_outputs(811) <= 1'b1;
    layer0_outputs(812) <= b and not a;
    layer0_outputs(813) <= not a;
    layer0_outputs(814) <= b and not a;
    layer0_outputs(815) <= a or b;
    layer0_outputs(816) <= 1'b0;
    layer0_outputs(817) <= a or b;
    layer0_outputs(818) <= not (a xor b);
    layer0_outputs(819) <= a or b;
    layer0_outputs(820) <= not b;
    layer0_outputs(821) <= not b or a;
    layer0_outputs(822) <= a and not b;
    layer0_outputs(823) <= not b or a;
    layer0_outputs(824) <= b;
    layer0_outputs(825) <= not (a or b);
    layer0_outputs(826) <= not (a xor b);
    layer0_outputs(827) <= b and not a;
    layer0_outputs(828) <= not b or a;
    layer0_outputs(829) <= a;
    layer0_outputs(830) <= not b;
    layer0_outputs(831) <= a;
    layer0_outputs(832) <= not b or a;
    layer0_outputs(833) <= not a;
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= b and not a;
    layer0_outputs(836) <= not a;
    layer0_outputs(837) <= not a;
    layer0_outputs(838) <= a or b;
    layer0_outputs(839) <= not a;
    layer0_outputs(840) <= not b;
    layer0_outputs(841) <= a or b;
    layer0_outputs(842) <= a or b;
    layer0_outputs(843) <= a;
    layer0_outputs(844) <= a or b;
    layer0_outputs(845) <= not (a or b);
    layer0_outputs(846) <= 1'b0;
    layer0_outputs(847) <= a and b;
    layer0_outputs(848) <= not (a or b);
    layer0_outputs(849) <= not b or a;
    layer0_outputs(850) <= not (a and b);
    layer0_outputs(851) <= a and b;
    layer0_outputs(852) <= a;
    layer0_outputs(853) <= not (a xor b);
    layer0_outputs(854) <= not b or a;
    layer0_outputs(855) <= a and not b;
    layer0_outputs(856) <= not a;
    layer0_outputs(857) <= not b or a;
    layer0_outputs(858) <= not a;
    layer0_outputs(859) <= not a;
    layer0_outputs(860) <= not a;
    layer0_outputs(861) <= not a or b;
    layer0_outputs(862) <= not (a xor b);
    layer0_outputs(863) <= 1'b0;
    layer0_outputs(864) <= a or b;
    layer0_outputs(865) <= a xor b;
    layer0_outputs(866) <= b;
    layer0_outputs(867) <= not (a xor b);
    layer0_outputs(868) <= a and not b;
    layer0_outputs(869) <= not (a or b);
    layer0_outputs(870) <= not b or a;
    layer0_outputs(871) <= not a;
    layer0_outputs(872) <= not (a xor b);
    layer0_outputs(873) <= not (a or b);
    layer0_outputs(874) <= not b;
    layer0_outputs(875) <= not (a or b);
    layer0_outputs(876) <= b;
    layer0_outputs(877) <= not (a xor b);
    layer0_outputs(878) <= not (a or b);
    layer0_outputs(879) <= not b or a;
    layer0_outputs(880) <= b and not a;
    layer0_outputs(881) <= a or b;
    layer0_outputs(882) <= not a or b;
    layer0_outputs(883) <= not a;
    layer0_outputs(884) <= a or b;
    layer0_outputs(885) <= not b;
    layer0_outputs(886) <= a xor b;
    layer0_outputs(887) <= not a or b;
    layer0_outputs(888) <= a or b;
    layer0_outputs(889) <= a xor b;
    layer0_outputs(890) <= 1'b1;
    layer0_outputs(891) <= a and not b;
    layer0_outputs(892) <= a or b;
    layer0_outputs(893) <= not a or b;
    layer0_outputs(894) <= a or b;
    layer0_outputs(895) <= not a or b;
    layer0_outputs(896) <= b and not a;
    layer0_outputs(897) <= not (a or b);
    layer0_outputs(898) <= not b;
    layer0_outputs(899) <= not b or a;
    layer0_outputs(900) <= not b;
    layer0_outputs(901) <= a or b;
    layer0_outputs(902) <= not (a or b);
    layer0_outputs(903) <= a or b;
    layer0_outputs(904) <= not a;
    layer0_outputs(905) <= not a;
    layer0_outputs(906) <= a and not b;
    layer0_outputs(907) <= a;
    layer0_outputs(908) <= not a or b;
    layer0_outputs(909) <= a;
    layer0_outputs(910) <= a or b;
    layer0_outputs(911) <= not (a xor b);
    layer0_outputs(912) <= a or b;
    layer0_outputs(913) <= a or b;
    layer0_outputs(914) <= a and not b;
    layer0_outputs(915) <= a;
    layer0_outputs(916) <= b and not a;
    layer0_outputs(917) <= not a or b;
    layer0_outputs(918) <= not b or a;
    layer0_outputs(919) <= a;
    layer0_outputs(920) <= not a or b;
    layer0_outputs(921) <= not (a or b);
    layer0_outputs(922) <= not (a or b);
    layer0_outputs(923) <= not a or b;
    layer0_outputs(924) <= b and not a;
    layer0_outputs(925) <= 1'b1;
    layer0_outputs(926) <= b;
    layer0_outputs(927) <= b;
    layer0_outputs(928) <= b;
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= b;
    layer0_outputs(931) <= a;
    layer0_outputs(932) <= a;
    layer0_outputs(933) <= not a or b;
    layer0_outputs(934) <= b;
    layer0_outputs(935) <= not b;
    layer0_outputs(936) <= a or b;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= b;
    layer0_outputs(939) <= not (a xor b);
    layer0_outputs(940) <= b;
    layer0_outputs(941) <= b and not a;
    layer0_outputs(942) <= a and not b;
    layer0_outputs(943) <= a;
    layer0_outputs(944) <= b and not a;
    layer0_outputs(945) <= b and not a;
    layer0_outputs(946) <= a and b;
    layer0_outputs(947) <= not (a or b);
    layer0_outputs(948) <= not b or a;
    layer0_outputs(949) <= a;
    layer0_outputs(950) <= a;
    layer0_outputs(951) <= not a or b;
    layer0_outputs(952) <= a or b;
    layer0_outputs(953) <= not (a or b);
    layer0_outputs(954) <= not (a xor b);
    layer0_outputs(955) <= not b or a;
    layer0_outputs(956) <= b and not a;
    layer0_outputs(957) <= not (a xor b);
    layer0_outputs(958) <= not b or a;
    layer0_outputs(959) <= not b;
    layer0_outputs(960) <= not b or a;
    layer0_outputs(961) <= not b;
    layer0_outputs(962) <= a xor b;
    layer0_outputs(963) <= not (a or b);
    layer0_outputs(964) <= 1'b1;
    layer0_outputs(965) <= not (a or b);
    layer0_outputs(966) <= not a;
    layer0_outputs(967) <= b and not a;
    layer0_outputs(968) <= a and b;
    layer0_outputs(969) <= b;
    layer0_outputs(970) <= a and b;
    layer0_outputs(971) <= not a;
    layer0_outputs(972) <= a and not b;
    layer0_outputs(973) <= not (a or b);
    layer0_outputs(974) <= not a;
    layer0_outputs(975) <= 1'b1;
    layer0_outputs(976) <= a or b;
    layer0_outputs(977) <= b;
    layer0_outputs(978) <= not a;
    layer0_outputs(979) <= 1'b1;
    layer0_outputs(980) <= not a;
    layer0_outputs(981) <= not (a xor b);
    layer0_outputs(982) <= a or b;
    layer0_outputs(983) <= not (a or b);
    layer0_outputs(984) <= a xor b;
    layer0_outputs(985) <= not (a xor b);
    layer0_outputs(986) <= not b or a;
    layer0_outputs(987) <= a;
    layer0_outputs(988) <= 1'b1;
    layer0_outputs(989) <= not (a and b);
    layer0_outputs(990) <= b;
    layer0_outputs(991) <= a and not b;
    layer0_outputs(992) <= a and not b;
    layer0_outputs(993) <= not (a or b);
    layer0_outputs(994) <= b;
    layer0_outputs(995) <= not b or a;
    layer0_outputs(996) <= a or b;
    layer0_outputs(997) <= b and not a;
    layer0_outputs(998) <= not b or a;
    layer0_outputs(999) <= not b or a;
    layer0_outputs(1000) <= a or b;
    layer0_outputs(1001) <= b;
    layer0_outputs(1002) <= not a;
    layer0_outputs(1003) <= b and not a;
    layer0_outputs(1004) <= a xor b;
    layer0_outputs(1005) <= not b;
    layer0_outputs(1006) <= a and not b;
    layer0_outputs(1007) <= a xor b;
    layer0_outputs(1008) <= b;
    layer0_outputs(1009) <= not (a xor b);
    layer0_outputs(1010) <= a xor b;
    layer0_outputs(1011) <= not a;
    layer0_outputs(1012) <= a or b;
    layer0_outputs(1013) <= a or b;
    layer0_outputs(1014) <= not (a or b);
    layer0_outputs(1015) <= not (a and b);
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= not a or b;
    layer0_outputs(1018) <= a xor b;
    layer0_outputs(1019) <= not b;
    layer0_outputs(1020) <= not a;
    layer0_outputs(1021) <= a and b;
    layer0_outputs(1022) <= 1'b0;
    layer0_outputs(1023) <= b;
    layer0_outputs(1024) <= a;
    layer0_outputs(1025) <= not (a xor b);
    layer0_outputs(1026) <= a or b;
    layer0_outputs(1027) <= not b;
    layer0_outputs(1028) <= a or b;
    layer0_outputs(1029) <= b and not a;
    layer0_outputs(1030) <= a;
    layer0_outputs(1031) <= b and not a;
    layer0_outputs(1032) <= a xor b;
    layer0_outputs(1033) <= not b or a;
    layer0_outputs(1034) <= not a;
    layer0_outputs(1035) <= a;
    layer0_outputs(1036) <= a xor b;
    layer0_outputs(1037) <= not b;
    layer0_outputs(1038) <= not a or b;
    layer0_outputs(1039) <= 1'b1;
    layer0_outputs(1040) <= a and b;
    layer0_outputs(1041) <= b;
    layer0_outputs(1042) <= b;
    layer0_outputs(1043) <= a or b;
    layer0_outputs(1044) <= 1'b0;
    layer0_outputs(1045) <= not (a or b);
    layer0_outputs(1046) <= a;
    layer0_outputs(1047) <= b;
    layer0_outputs(1048) <= b and not a;
    layer0_outputs(1049) <= 1'b1;
    layer0_outputs(1050) <= not (a and b);
    layer0_outputs(1051) <= b;
    layer0_outputs(1052) <= not a;
    layer0_outputs(1053) <= not a;
    layer0_outputs(1054) <= not b or a;
    layer0_outputs(1055) <= not a;
    layer0_outputs(1056) <= not a;
    layer0_outputs(1057) <= 1'b0;
    layer0_outputs(1058) <= not b;
    layer0_outputs(1059) <= not (a and b);
    layer0_outputs(1060) <= b;
    layer0_outputs(1061) <= 1'b1;
    layer0_outputs(1062) <= not (a xor b);
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= not a or b;
    layer0_outputs(1065) <= not a;
    layer0_outputs(1066) <= a or b;
    layer0_outputs(1067) <= not a;
    layer0_outputs(1068) <= not b or a;
    layer0_outputs(1069) <= not (a and b);
    layer0_outputs(1070) <= b;
    layer0_outputs(1071) <= not (a or b);
    layer0_outputs(1072) <= not a;
    layer0_outputs(1073) <= a or b;
    layer0_outputs(1074) <= b;
    layer0_outputs(1075) <= a and not b;
    layer0_outputs(1076) <= a xor b;
    layer0_outputs(1077) <= not (a xor b);
    layer0_outputs(1078) <= a;
    layer0_outputs(1079) <= not b;
    layer0_outputs(1080) <= not b;
    layer0_outputs(1081) <= a and not b;
    layer0_outputs(1082) <= 1'b0;
    layer0_outputs(1083) <= not (a or b);
    layer0_outputs(1084) <= not (a xor b);
    layer0_outputs(1085) <= not (a xor b);
    layer0_outputs(1086) <= not b or a;
    layer0_outputs(1087) <= not a;
    layer0_outputs(1088) <= not a or b;
    layer0_outputs(1089) <= a and not b;
    layer0_outputs(1090) <= not (a or b);
    layer0_outputs(1091) <= a;
    layer0_outputs(1092) <= a xor b;
    layer0_outputs(1093) <= a and b;
    layer0_outputs(1094) <= not b or a;
    layer0_outputs(1095) <= a;
    layer0_outputs(1096) <= not b;
    layer0_outputs(1097) <= not a;
    layer0_outputs(1098) <= 1'b0;
    layer0_outputs(1099) <= a and not b;
    layer0_outputs(1100) <= not b or a;
    layer0_outputs(1101) <= b;
    layer0_outputs(1102) <= b;
    layer0_outputs(1103) <= a or b;
    layer0_outputs(1104) <= not b;
    layer0_outputs(1105) <= not b;
    layer0_outputs(1106) <= a or b;
    layer0_outputs(1107) <= a or b;
    layer0_outputs(1108) <= 1'b0;
    layer0_outputs(1109) <= not (a or b);
    layer0_outputs(1110) <= not a;
    layer0_outputs(1111) <= not b;
    layer0_outputs(1112) <= a or b;
    layer0_outputs(1113) <= b;
    layer0_outputs(1114) <= not (a or b);
    layer0_outputs(1115) <= not b or a;
    layer0_outputs(1116) <= not (a or b);
    layer0_outputs(1117) <= not (a or b);
    layer0_outputs(1118) <= not a;
    layer0_outputs(1119) <= a and not b;
    layer0_outputs(1120) <= not (a or b);
    layer0_outputs(1121) <= a;
    layer0_outputs(1122) <= not (a xor b);
    layer0_outputs(1123) <= b;
    layer0_outputs(1124) <= not b or a;
    layer0_outputs(1125) <= not b;
    layer0_outputs(1126) <= b;
    layer0_outputs(1127) <= not (a or b);
    layer0_outputs(1128) <= a xor b;
    layer0_outputs(1129) <= b and not a;
    layer0_outputs(1130) <= 1'b0;
    layer0_outputs(1131) <= not (a xor b);
    layer0_outputs(1132) <= not b or a;
    layer0_outputs(1133) <= not (a or b);
    layer0_outputs(1134) <= not b or a;
    layer0_outputs(1135) <= a and b;
    layer0_outputs(1136) <= 1'b0;
    layer0_outputs(1137) <= not (a xor b);
    layer0_outputs(1138) <= 1'b0;
    layer0_outputs(1139) <= b and not a;
    layer0_outputs(1140) <= a or b;
    layer0_outputs(1141) <= not a;
    layer0_outputs(1142) <= b and not a;
    layer0_outputs(1143) <= a and b;
    layer0_outputs(1144) <= a or b;
    layer0_outputs(1145) <= not a or b;
    layer0_outputs(1146) <= not (a or b);
    layer0_outputs(1147) <= b;
    layer0_outputs(1148) <= a;
    layer0_outputs(1149) <= b;
    layer0_outputs(1150) <= not (a and b);
    layer0_outputs(1151) <= not (a and b);
    layer0_outputs(1152) <= not b or a;
    layer0_outputs(1153) <= not b or a;
    layer0_outputs(1154) <= a or b;
    layer0_outputs(1155) <= not (a and b);
    layer0_outputs(1156) <= not a or b;
    layer0_outputs(1157) <= not a or b;
    layer0_outputs(1158) <= not (a and b);
    layer0_outputs(1159) <= a or b;
    layer0_outputs(1160) <= not b or a;
    layer0_outputs(1161) <= not b or a;
    layer0_outputs(1162) <= not (a or b);
    layer0_outputs(1163) <= a and b;
    layer0_outputs(1164) <= not (a and b);
    layer0_outputs(1165) <= a xor b;
    layer0_outputs(1166) <= not (a xor b);
    layer0_outputs(1167) <= a xor b;
    layer0_outputs(1168) <= not (a and b);
    layer0_outputs(1169) <= a;
    layer0_outputs(1170) <= 1'b0;
    layer0_outputs(1171) <= not a or b;
    layer0_outputs(1172) <= not (a or b);
    layer0_outputs(1173) <= b;
    layer0_outputs(1174) <= b and not a;
    layer0_outputs(1175) <= not b;
    layer0_outputs(1176) <= b and not a;
    layer0_outputs(1177) <= a xor b;
    layer0_outputs(1178) <= not (a and b);
    layer0_outputs(1179) <= not b;
    layer0_outputs(1180) <= b;
    layer0_outputs(1181) <= not (a xor b);
    layer0_outputs(1182) <= a or b;
    layer0_outputs(1183) <= 1'b1;
    layer0_outputs(1184) <= not a or b;
    layer0_outputs(1185) <= 1'b0;
    layer0_outputs(1186) <= not (a and b);
    layer0_outputs(1187) <= a xor b;
    layer0_outputs(1188) <= not (a or b);
    layer0_outputs(1189) <= a or b;
    layer0_outputs(1190) <= a;
    layer0_outputs(1191) <= a;
    layer0_outputs(1192) <= a or b;
    layer0_outputs(1193) <= not (a or b);
    layer0_outputs(1194) <= not a or b;
    layer0_outputs(1195) <= 1'b0;
    layer0_outputs(1196) <= a xor b;
    layer0_outputs(1197) <= not a or b;
    layer0_outputs(1198) <= a xor b;
    layer0_outputs(1199) <= not (a xor b);
    layer0_outputs(1200) <= a;
    layer0_outputs(1201) <= not (a or b);
    layer0_outputs(1202) <= not a or b;
    layer0_outputs(1203) <= a xor b;
    layer0_outputs(1204) <= not a or b;
    layer0_outputs(1205) <= not b or a;
    layer0_outputs(1206) <= not b;
    layer0_outputs(1207) <= not (a or b);
    layer0_outputs(1208) <= not (a or b);
    layer0_outputs(1209) <= a;
    layer0_outputs(1210) <= not b or a;
    layer0_outputs(1211) <= a or b;
    layer0_outputs(1212) <= not (a and b);
    layer0_outputs(1213) <= not (a xor b);
    layer0_outputs(1214) <= not a;
    layer0_outputs(1215) <= not a;
    layer0_outputs(1216) <= a or b;
    layer0_outputs(1217) <= not (a or b);
    layer0_outputs(1218) <= a and not b;
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= not b;
    layer0_outputs(1221) <= not b or a;
    layer0_outputs(1222) <= a or b;
    layer0_outputs(1223) <= a xor b;
    layer0_outputs(1224) <= not (a or b);
    layer0_outputs(1225) <= not b or a;
    layer0_outputs(1226) <= a and not b;
    layer0_outputs(1227) <= not b;
    layer0_outputs(1228) <= a or b;
    layer0_outputs(1229) <= not b or a;
    layer0_outputs(1230) <= not b;
    layer0_outputs(1231) <= a xor b;
    layer0_outputs(1232) <= a xor b;
    layer0_outputs(1233) <= not (a and b);
    layer0_outputs(1234) <= a or b;
    layer0_outputs(1235) <= not (a and b);
    layer0_outputs(1236) <= not b or a;
    layer0_outputs(1237) <= a xor b;
    layer0_outputs(1238) <= not a or b;
    layer0_outputs(1239) <= b and not a;
    layer0_outputs(1240) <= a;
    layer0_outputs(1241) <= not a;
    layer0_outputs(1242) <= b and not a;
    layer0_outputs(1243) <= a or b;
    layer0_outputs(1244) <= not (a or b);
    layer0_outputs(1245) <= a;
    layer0_outputs(1246) <= 1'b1;
    layer0_outputs(1247) <= a or b;
    layer0_outputs(1248) <= a or b;
    layer0_outputs(1249) <= not b;
    layer0_outputs(1250) <= not a or b;
    layer0_outputs(1251) <= not (a or b);
    layer0_outputs(1252) <= b and not a;
    layer0_outputs(1253) <= not (a or b);
    layer0_outputs(1254) <= not a or b;
    layer0_outputs(1255) <= b;
    layer0_outputs(1256) <= not (a and b);
    layer0_outputs(1257) <= b;
    layer0_outputs(1258) <= not a;
    layer0_outputs(1259) <= b and not a;
    layer0_outputs(1260) <= not (a or b);
    layer0_outputs(1261) <= b;
    layer0_outputs(1262) <= b;
    layer0_outputs(1263) <= 1'b0;
    layer0_outputs(1264) <= not b;
    layer0_outputs(1265) <= a and b;
    layer0_outputs(1266) <= 1'b0;
    layer0_outputs(1267) <= not (a or b);
    layer0_outputs(1268) <= not (a xor b);
    layer0_outputs(1269) <= b and not a;
    layer0_outputs(1270) <= b;
    layer0_outputs(1271) <= not b or a;
    layer0_outputs(1272) <= a or b;
    layer0_outputs(1273) <= a or b;
    layer0_outputs(1274) <= a and b;
    layer0_outputs(1275) <= a and not b;
    layer0_outputs(1276) <= a and not b;
    layer0_outputs(1277) <= a xor b;
    layer0_outputs(1278) <= not (a or b);
    layer0_outputs(1279) <= not a or b;
    layer0_outputs(1280) <= 1'b0;
    layer0_outputs(1281) <= not a or b;
    layer0_outputs(1282) <= b;
    layer0_outputs(1283) <= not (a or b);
    layer0_outputs(1284) <= b and not a;
    layer0_outputs(1285) <= not (a and b);
    layer0_outputs(1286) <= not (a and b);
    layer0_outputs(1287) <= not a;
    layer0_outputs(1288) <= not b or a;
    layer0_outputs(1289) <= a and not b;
    layer0_outputs(1290) <= a or b;
    layer0_outputs(1291) <= 1'b1;
    layer0_outputs(1292) <= a;
    layer0_outputs(1293) <= b and not a;
    layer0_outputs(1294) <= a;
    layer0_outputs(1295) <= a;
    layer0_outputs(1296) <= 1'b1;
    layer0_outputs(1297) <= a xor b;
    layer0_outputs(1298) <= not (a or b);
    layer0_outputs(1299) <= not a;
    layer0_outputs(1300) <= a xor b;
    layer0_outputs(1301) <= 1'b0;
    layer0_outputs(1302) <= a and b;
    layer0_outputs(1303) <= not (a or b);
    layer0_outputs(1304) <= a or b;
    layer0_outputs(1305) <= not (a xor b);
    layer0_outputs(1306) <= not (a or b);
    layer0_outputs(1307) <= not (a xor b);
    layer0_outputs(1308) <= not (a or b);
    layer0_outputs(1309) <= not (a or b);
    layer0_outputs(1310) <= not (a xor b);
    layer0_outputs(1311) <= not b;
    layer0_outputs(1312) <= a or b;
    layer0_outputs(1313) <= a;
    layer0_outputs(1314) <= 1'b1;
    layer0_outputs(1315) <= a and b;
    layer0_outputs(1316) <= 1'b1;
    layer0_outputs(1317) <= not (a and b);
    layer0_outputs(1318) <= not a or b;
    layer0_outputs(1319) <= not a or b;
    layer0_outputs(1320) <= not b or a;
    layer0_outputs(1321) <= not (a and b);
    layer0_outputs(1322) <= a;
    layer0_outputs(1323) <= not b or a;
    layer0_outputs(1324) <= b;
    layer0_outputs(1325) <= not a;
    layer0_outputs(1326) <= not (a or b);
    layer0_outputs(1327) <= a;
    layer0_outputs(1328) <= not b;
    layer0_outputs(1329) <= not (a and b);
    layer0_outputs(1330) <= a and not b;
    layer0_outputs(1331) <= not (a and b);
    layer0_outputs(1332) <= 1'b1;
    layer0_outputs(1333) <= not b;
    layer0_outputs(1334) <= not (a or b);
    layer0_outputs(1335) <= not a;
    layer0_outputs(1336) <= b;
    layer0_outputs(1337) <= a;
    layer0_outputs(1338) <= a;
    layer0_outputs(1339) <= not (a or b);
    layer0_outputs(1340) <= a;
    layer0_outputs(1341) <= not b;
    layer0_outputs(1342) <= not (a or b);
    layer0_outputs(1343) <= a or b;
    layer0_outputs(1344) <= a or b;
    layer0_outputs(1345) <= a or b;
    layer0_outputs(1346) <= not a or b;
    layer0_outputs(1347) <= a xor b;
    layer0_outputs(1348) <= b and not a;
    layer0_outputs(1349) <= 1'b1;
    layer0_outputs(1350) <= b;
    layer0_outputs(1351) <= b and not a;
    layer0_outputs(1352) <= 1'b0;
    layer0_outputs(1353) <= 1'b0;
    layer0_outputs(1354) <= not a;
    layer0_outputs(1355) <= b;
    layer0_outputs(1356) <= a;
    layer0_outputs(1357) <= a and b;
    layer0_outputs(1358) <= 1'b0;
    layer0_outputs(1359) <= not a;
    layer0_outputs(1360) <= not b or a;
    layer0_outputs(1361) <= not (a or b);
    layer0_outputs(1362) <= b;
    layer0_outputs(1363) <= not b or a;
    layer0_outputs(1364) <= not (a xor b);
    layer0_outputs(1365) <= a;
    layer0_outputs(1366) <= not a or b;
    layer0_outputs(1367) <= not (a or b);
    layer0_outputs(1368) <= not (a or b);
    layer0_outputs(1369) <= a;
    layer0_outputs(1370) <= not (a or b);
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= not (a xor b);
    layer0_outputs(1373) <= not (a xor b);
    layer0_outputs(1374) <= not (a or b);
    layer0_outputs(1375) <= not (a and b);
    layer0_outputs(1376) <= not b or a;
    layer0_outputs(1377) <= not b;
    layer0_outputs(1378) <= not (a or b);
    layer0_outputs(1379) <= b and not a;
    layer0_outputs(1380) <= a and not b;
    layer0_outputs(1381) <= not (a and b);
    layer0_outputs(1382) <= a and not b;
    layer0_outputs(1383) <= b;
    layer0_outputs(1384) <= a or b;
    layer0_outputs(1385) <= a and not b;
    layer0_outputs(1386) <= a or b;
    layer0_outputs(1387) <= a or b;
    layer0_outputs(1388) <= not b or a;
    layer0_outputs(1389) <= not (a and b);
    layer0_outputs(1390) <= not (a or b);
    layer0_outputs(1391) <= not (a and b);
    layer0_outputs(1392) <= 1'b0;
    layer0_outputs(1393) <= not (a or b);
    layer0_outputs(1394) <= not b;
    layer0_outputs(1395) <= b;
    layer0_outputs(1396) <= b;
    layer0_outputs(1397) <= b and not a;
    layer0_outputs(1398) <= not b;
    layer0_outputs(1399) <= b and not a;
    layer0_outputs(1400) <= not b;
    layer0_outputs(1401) <= b;
    layer0_outputs(1402) <= not a;
    layer0_outputs(1403) <= not (a or b);
    layer0_outputs(1404) <= a xor b;
    layer0_outputs(1405) <= a or b;
    layer0_outputs(1406) <= 1'b0;
    layer0_outputs(1407) <= a;
    layer0_outputs(1408) <= not (a and b);
    layer0_outputs(1409) <= a xor b;
    layer0_outputs(1410) <= not a or b;
    layer0_outputs(1411) <= b;
    layer0_outputs(1412) <= a or b;
    layer0_outputs(1413) <= 1'b0;
    layer0_outputs(1414) <= not (a or b);
    layer0_outputs(1415) <= not a;
    layer0_outputs(1416) <= a;
    layer0_outputs(1417) <= b;
    layer0_outputs(1418) <= a and not b;
    layer0_outputs(1419) <= a and not b;
    layer0_outputs(1420) <= b;
    layer0_outputs(1421) <= not (a or b);
    layer0_outputs(1422) <= b and not a;
    layer0_outputs(1423) <= a;
    layer0_outputs(1424) <= a or b;
    layer0_outputs(1425) <= not a;
    layer0_outputs(1426) <= b and not a;
    layer0_outputs(1427) <= not (a or b);
    layer0_outputs(1428) <= 1'b1;
    layer0_outputs(1429) <= a or b;
    layer0_outputs(1430) <= not (a xor b);
    layer0_outputs(1431) <= not b;
    layer0_outputs(1432) <= not a or b;
    layer0_outputs(1433) <= 1'b1;
    layer0_outputs(1434) <= not a;
    layer0_outputs(1435) <= a and b;
    layer0_outputs(1436) <= a or b;
    layer0_outputs(1437) <= a;
    layer0_outputs(1438) <= a;
    layer0_outputs(1439) <= not (a or b);
    layer0_outputs(1440) <= not a or b;
    layer0_outputs(1441) <= not b;
    layer0_outputs(1442) <= a and b;
    layer0_outputs(1443) <= a xor b;
    layer0_outputs(1444) <= not (a or b);
    layer0_outputs(1445) <= a or b;
    layer0_outputs(1446) <= not (a xor b);
    layer0_outputs(1447) <= a and not b;
    layer0_outputs(1448) <= a and not b;
    layer0_outputs(1449) <= not b or a;
    layer0_outputs(1450) <= not (a and b);
    layer0_outputs(1451) <= a or b;
    layer0_outputs(1452) <= not a or b;
    layer0_outputs(1453) <= not (a or b);
    layer0_outputs(1454) <= b and not a;
    layer0_outputs(1455) <= not (a xor b);
    layer0_outputs(1456) <= a;
    layer0_outputs(1457) <= a;
    layer0_outputs(1458) <= b;
    layer0_outputs(1459) <= 1'b1;
    layer0_outputs(1460) <= b;
    layer0_outputs(1461) <= not a;
    layer0_outputs(1462) <= a and b;
    layer0_outputs(1463) <= a and not b;
    layer0_outputs(1464) <= a;
    layer0_outputs(1465) <= not b;
    layer0_outputs(1466) <= a xor b;
    layer0_outputs(1467) <= not a;
    layer0_outputs(1468) <= a xor b;
    layer0_outputs(1469) <= not (a or b);
    layer0_outputs(1470) <= a xor b;
    layer0_outputs(1471) <= a;
    layer0_outputs(1472) <= not b or a;
    layer0_outputs(1473) <= a or b;
    layer0_outputs(1474) <= b;
    layer0_outputs(1475) <= b and not a;
    layer0_outputs(1476) <= not (a or b);
    layer0_outputs(1477) <= not a;
    layer0_outputs(1478) <= b;
    layer0_outputs(1479) <= a;
    layer0_outputs(1480) <= a or b;
    layer0_outputs(1481) <= not (a or b);
    layer0_outputs(1482) <= not a;
    layer0_outputs(1483) <= a and not b;
    layer0_outputs(1484) <= a;
    layer0_outputs(1485) <= not a;
    layer0_outputs(1486) <= not a or b;
    layer0_outputs(1487) <= not (a xor b);
    layer0_outputs(1488) <= b;
    layer0_outputs(1489) <= not a;
    layer0_outputs(1490) <= not b;
    layer0_outputs(1491) <= a;
    layer0_outputs(1492) <= not (a xor b);
    layer0_outputs(1493) <= a or b;
    layer0_outputs(1494) <= not a or b;
    layer0_outputs(1495) <= not (a or b);
    layer0_outputs(1496) <= 1'b1;
    layer0_outputs(1497) <= 1'b1;
    layer0_outputs(1498) <= a or b;
    layer0_outputs(1499) <= b;
    layer0_outputs(1500) <= 1'b0;
    layer0_outputs(1501) <= b;
    layer0_outputs(1502) <= a and b;
    layer0_outputs(1503) <= a;
    layer0_outputs(1504) <= not (a or b);
    layer0_outputs(1505) <= a or b;
    layer0_outputs(1506) <= not b;
    layer0_outputs(1507) <= not (a xor b);
    layer0_outputs(1508) <= not a;
    layer0_outputs(1509) <= b and not a;
    layer0_outputs(1510) <= not a;
    layer0_outputs(1511) <= not a;
    layer0_outputs(1512) <= 1'b0;
    layer0_outputs(1513) <= not b or a;
    layer0_outputs(1514) <= a and not b;
    layer0_outputs(1515) <= a or b;
    layer0_outputs(1516) <= b and not a;
    layer0_outputs(1517) <= not (a and b);
    layer0_outputs(1518) <= not (a or b);
    layer0_outputs(1519) <= a or b;
    layer0_outputs(1520) <= a and b;
    layer0_outputs(1521) <= not b or a;
    layer0_outputs(1522) <= not (a xor b);
    layer0_outputs(1523) <= a xor b;
    layer0_outputs(1524) <= a xor b;
    layer0_outputs(1525) <= not b;
    layer0_outputs(1526) <= not b or a;
    layer0_outputs(1527) <= b;
    layer0_outputs(1528) <= not a or b;
    layer0_outputs(1529) <= b;
    layer0_outputs(1530) <= a and not b;
    layer0_outputs(1531) <= not (a xor b);
    layer0_outputs(1532) <= a and not b;
    layer0_outputs(1533) <= a and not b;
    layer0_outputs(1534) <= not a or b;
    layer0_outputs(1535) <= b and not a;
    layer0_outputs(1536) <= b;
    layer0_outputs(1537) <= not b;
    layer0_outputs(1538) <= not (a or b);
    layer0_outputs(1539) <= not a;
    layer0_outputs(1540) <= a or b;
    layer0_outputs(1541) <= a;
    layer0_outputs(1542) <= a or b;
    layer0_outputs(1543) <= a or b;
    layer0_outputs(1544) <= not b or a;
    layer0_outputs(1545) <= not a or b;
    layer0_outputs(1546) <= not a;
    layer0_outputs(1547) <= a or b;
    layer0_outputs(1548) <= not b or a;
    layer0_outputs(1549) <= b;
    layer0_outputs(1550) <= not b or a;
    layer0_outputs(1551) <= not b;
    layer0_outputs(1552) <= not a;
    layer0_outputs(1553) <= a;
    layer0_outputs(1554) <= a or b;
    layer0_outputs(1555) <= a and b;
    layer0_outputs(1556) <= not (a or b);
    layer0_outputs(1557) <= b;
    layer0_outputs(1558) <= a;
    layer0_outputs(1559) <= not (a xor b);
    layer0_outputs(1560) <= a;
    layer0_outputs(1561) <= b and not a;
    layer0_outputs(1562) <= not b;
    layer0_outputs(1563) <= 1'b0;
    layer0_outputs(1564) <= 1'b1;
    layer0_outputs(1565) <= a or b;
    layer0_outputs(1566) <= not b;
    layer0_outputs(1567) <= a xor b;
    layer0_outputs(1568) <= a;
    layer0_outputs(1569) <= not (a and b);
    layer0_outputs(1570) <= a xor b;
    layer0_outputs(1571) <= a;
    layer0_outputs(1572) <= not b;
    layer0_outputs(1573) <= not a;
    layer0_outputs(1574) <= 1'b1;
    layer0_outputs(1575) <= not b;
    layer0_outputs(1576) <= b;
    layer0_outputs(1577) <= not b;
    layer0_outputs(1578) <= 1'b0;
    layer0_outputs(1579) <= not b;
    layer0_outputs(1580) <= a and not b;
    layer0_outputs(1581) <= b;
    layer0_outputs(1582) <= not b;
    layer0_outputs(1583) <= a or b;
    layer0_outputs(1584) <= not (a or b);
    layer0_outputs(1585) <= not (a and b);
    layer0_outputs(1586) <= not a or b;
    layer0_outputs(1587) <= b;
    layer0_outputs(1588) <= a xor b;
    layer0_outputs(1589) <= not (a xor b);
    layer0_outputs(1590) <= not (a or b);
    layer0_outputs(1591) <= not b;
    layer0_outputs(1592) <= not a;
    layer0_outputs(1593) <= b;
    layer0_outputs(1594) <= not b or a;
    layer0_outputs(1595) <= not b or a;
    layer0_outputs(1596) <= not b;
    layer0_outputs(1597) <= a or b;
    layer0_outputs(1598) <= 1'b1;
    layer0_outputs(1599) <= 1'b1;
    layer0_outputs(1600) <= a xor b;
    layer0_outputs(1601) <= a xor b;
    layer0_outputs(1602) <= not a;
    layer0_outputs(1603) <= a and not b;
    layer0_outputs(1604) <= b;
    layer0_outputs(1605) <= not a;
    layer0_outputs(1606) <= 1'b1;
    layer0_outputs(1607) <= b and not a;
    layer0_outputs(1608) <= a or b;
    layer0_outputs(1609) <= not (a xor b);
    layer0_outputs(1610) <= not b or a;
    layer0_outputs(1611) <= b and not a;
    layer0_outputs(1612) <= not b or a;
    layer0_outputs(1613) <= a or b;
    layer0_outputs(1614) <= a or b;
    layer0_outputs(1615) <= a or b;
    layer0_outputs(1616) <= not a;
    layer0_outputs(1617) <= a or b;
    layer0_outputs(1618) <= not b;
    layer0_outputs(1619) <= not b;
    layer0_outputs(1620) <= not (a xor b);
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= b;
    layer0_outputs(1623) <= b;
    layer0_outputs(1624) <= a and b;
    layer0_outputs(1625) <= not b or a;
    layer0_outputs(1626) <= not (a xor b);
    layer0_outputs(1627) <= not (a xor b);
    layer0_outputs(1628) <= not (a and b);
    layer0_outputs(1629) <= a;
    layer0_outputs(1630) <= not (a xor b);
    layer0_outputs(1631) <= a or b;
    layer0_outputs(1632) <= a and not b;
    layer0_outputs(1633) <= not a or b;
    layer0_outputs(1634) <= a or b;
    layer0_outputs(1635) <= not (a xor b);
    layer0_outputs(1636) <= not a or b;
    layer0_outputs(1637) <= not (a or b);
    layer0_outputs(1638) <= not (a and b);
    layer0_outputs(1639) <= a or b;
    layer0_outputs(1640) <= 1'b0;
    layer0_outputs(1641) <= not b or a;
    layer0_outputs(1642) <= not a;
    layer0_outputs(1643) <= a xor b;
    layer0_outputs(1644) <= not a;
    layer0_outputs(1645) <= not a or b;
    layer0_outputs(1646) <= not (a xor b);
    layer0_outputs(1647) <= not (a or b);
    layer0_outputs(1648) <= a and not b;
    layer0_outputs(1649) <= a;
    layer0_outputs(1650) <= 1'b0;
    layer0_outputs(1651) <= a;
    layer0_outputs(1652) <= not b or a;
    layer0_outputs(1653) <= not (a xor b);
    layer0_outputs(1654) <= a or b;
    layer0_outputs(1655) <= a or b;
    layer0_outputs(1656) <= not b or a;
    layer0_outputs(1657) <= not (a and b);
    layer0_outputs(1658) <= not b;
    layer0_outputs(1659) <= not b;
    layer0_outputs(1660) <= not a or b;
    layer0_outputs(1661) <= a;
    layer0_outputs(1662) <= not b;
    layer0_outputs(1663) <= a and not b;
    layer0_outputs(1664) <= 1'b0;
    layer0_outputs(1665) <= 1'b1;
    layer0_outputs(1666) <= not b;
    layer0_outputs(1667) <= a;
    layer0_outputs(1668) <= 1'b0;
    layer0_outputs(1669) <= a;
    layer0_outputs(1670) <= a and not b;
    layer0_outputs(1671) <= not a;
    layer0_outputs(1672) <= a and not b;
    layer0_outputs(1673) <= not a;
    layer0_outputs(1674) <= not b;
    layer0_outputs(1675) <= a;
    layer0_outputs(1676) <= a and not b;
    layer0_outputs(1677) <= a and not b;
    layer0_outputs(1678) <= not (a xor b);
    layer0_outputs(1679) <= not a or b;
    layer0_outputs(1680) <= b and not a;
    layer0_outputs(1681) <= not (a xor b);
    layer0_outputs(1682) <= a and not b;
    layer0_outputs(1683) <= not a or b;
    layer0_outputs(1684) <= not (a and b);
    layer0_outputs(1685) <= a and b;
    layer0_outputs(1686) <= a or b;
    layer0_outputs(1687) <= not b or a;
    layer0_outputs(1688) <= b and not a;
    layer0_outputs(1689) <= not b or a;
    layer0_outputs(1690) <= a;
    layer0_outputs(1691) <= a or b;
    layer0_outputs(1692) <= a and b;
    layer0_outputs(1693) <= b;
    layer0_outputs(1694) <= not a;
    layer0_outputs(1695) <= b;
    layer0_outputs(1696) <= not b;
    layer0_outputs(1697) <= 1'b0;
    layer0_outputs(1698) <= a xor b;
    layer0_outputs(1699) <= not a;
    layer0_outputs(1700) <= not b or a;
    layer0_outputs(1701) <= a or b;
    layer0_outputs(1702) <= not (a or b);
    layer0_outputs(1703) <= not b;
    layer0_outputs(1704) <= not (a or b);
    layer0_outputs(1705) <= not a;
    layer0_outputs(1706) <= not (a or b);
    layer0_outputs(1707) <= not b or a;
    layer0_outputs(1708) <= a;
    layer0_outputs(1709) <= b;
    layer0_outputs(1710) <= not a;
    layer0_outputs(1711) <= not b or a;
    layer0_outputs(1712) <= not (a or b);
    layer0_outputs(1713) <= b and not a;
    layer0_outputs(1714) <= not (a or b);
    layer0_outputs(1715) <= not b or a;
    layer0_outputs(1716) <= a or b;
    layer0_outputs(1717) <= a and not b;
    layer0_outputs(1718) <= not (a xor b);
    layer0_outputs(1719) <= not a;
    layer0_outputs(1720) <= a or b;
    layer0_outputs(1721) <= b and not a;
    layer0_outputs(1722) <= a and not b;
    layer0_outputs(1723) <= a;
    layer0_outputs(1724) <= b;
    layer0_outputs(1725) <= 1'b1;
    layer0_outputs(1726) <= not (a xor b);
    layer0_outputs(1727) <= 1'b0;
    layer0_outputs(1728) <= not a or b;
    layer0_outputs(1729) <= a;
    layer0_outputs(1730) <= a and not b;
    layer0_outputs(1731) <= not (a or b);
    layer0_outputs(1732) <= b and not a;
    layer0_outputs(1733) <= 1'b0;
    layer0_outputs(1734) <= a and not b;
    layer0_outputs(1735) <= a or b;
    layer0_outputs(1736) <= not (a or b);
    layer0_outputs(1737) <= not (a xor b);
    layer0_outputs(1738) <= not (a xor b);
    layer0_outputs(1739) <= not b;
    layer0_outputs(1740) <= a xor b;
    layer0_outputs(1741) <= b;
    layer0_outputs(1742) <= not a;
    layer0_outputs(1743) <= a;
    layer0_outputs(1744) <= a;
    layer0_outputs(1745) <= not b;
    layer0_outputs(1746) <= b;
    layer0_outputs(1747) <= not (a xor b);
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= not (a or b);
    layer0_outputs(1750) <= a or b;
    layer0_outputs(1751) <= a and not b;
    layer0_outputs(1752) <= not (a xor b);
    layer0_outputs(1753) <= 1'b1;
    layer0_outputs(1754) <= not a;
    layer0_outputs(1755) <= a;
    layer0_outputs(1756) <= 1'b1;
    layer0_outputs(1757) <= not (a xor b);
    layer0_outputs(1758) <= 1'b1;
    layer0_outputs(1759) <= not b or a;
    layer0_outputs(1760) <= not (a xor b);
    layer0_outputs(1761) <= a xor b;
    layer0_outputs(1762) <= 1'b1;
    layer0_outputs(1763) <= not (a or b);
    layer0_outputs(1764) <= a;
    layer0_outputs(1765) <= a;
    layer0_outputs(1766) <= not (a or b);
    layer0_outputs(1767) <= not b or a;
    layer0_outputs(1768) <= not b;
    layer0_outputs(1769) <= a or b;
    layer0_outputs(1770) <= not a;
    layer0_outputs(1771) <= a and b;
    layer0_outputs(1772) <= a and b;
    layer0_outputs(1773) <= b;
    layer0_outputs(1774) <= not a;
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= a or b;
    layer0_outputs(1777) <= a or b;
    layer0_outputs(1778) <= not (a or b);
    layer0_outputs(1779) <= not (a xor b);
    layer0_outputs(1780) <= not b or a;
    layer0_outputs(1781) <= not b or a;
    layer0_outputs(1782) <= a;
    layer0_outputs(1783) <= a and b;
    layer0_outputs(1784) <= not b;
    layer0_outputs(1785) <= 1'b1;
    layer0_outputs(1786) <= not (a xor b);
    layer0_outputs(1787) <= b;
    layer0_outputs(1788) <= a or b;
    layer0_outputs(1789) <= b;
    layer0_outputs(1790) <= 1'b0;
    layer0_outputs(1791) <= 1'b0;
    layer0_outputs(1792) <= not a;
    layer0_outputs(1793) <= not a;
    layer0_outputs(1794) <= 1'b1;
    layer0_outputs(1795) <= 1'b0;
    layer0_outputs(1796) <= not b;
    layer0_outputs(1797) <= not (a or b);
    layer0_outputs(1798) <= b and not a;
    layer0_outputs(1799) <= a;
    layer0_outputs(1800) <= not (a or b);
    layer0_outputs(1801) <= b and not a;
    layer0_outputs(1802) <= not b or a;
    layer0_outputs(1803) <= b;
    layer0_outputs(1804) <= b;
    layer0_outputs(1805) <= a or b;
    layer0_outputs(1806) <= a xor b;
    layer0_outputs(1807) <= a and not b;
    layer0_outputs(1808) <= a;
    layer0_outputs(1809) <= not (a or b);
    layer0_outputs(1810) <= a and not b;
    layer0_outputs(1811) <= a and not b;
    layer0_outputs(1812) <= b;
    layer0_outputs(1813) <= a or b;
    layer0_outputs(1814) <= a or b;
    layer0_outputs(1815) <= a or b;
    layer0_outputs(1816) <= 1'b0;
    layer0_outputs(1817) <= not b;
    layer0_outputs(1818) <= a or b;
    layer0_outputs(1819) <= 1'b0;
    layer0_outputs(1820) <= not b or a;
    layer0_outputs(1821) <= a and not b;
    layer0_outputs(1822) <= b and not a;
    layer0_outputs(1823) <= not a;
    layer0_outputs(1824) <= a and b;
    layer0_outputs(1825) <= not b;
    layer0_outputs(1826) <= not (a xor b);
    layer0_outputs(1827) <= a xor b;
    layer0_outputs(1828) <= b;
    layer0_outputs(1829) <= not b;
    layer0_outputs(1830) <= not b;
    layer0_outputs(1831) <= a or b;
    layer0_outputs(1832) <= not a or b;
    layer0_outputs(1833) <= 1'b1;
    layer0_outputs(1834) <= not a or b;
    layer0_outputs(1835) <= b;
    layer0_outputs(1836) <= a or b;
    layer0_outputs(1837) <= not a or b;
    layer0_outputs(1838) <= b and not a;
    layer0_outputs(1839) <= a and not b;
    layer0_outputs(1840) <= not (a xor b);
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= b;
    layer0_outputs(1843) <= b;
    layer0_outputs(1844) <= not (a or b);
    layer0_outputs(1845) <= 1'b0;
    layer0_outputs(1846) <= not b;
    layer0_outputs(1847) <= a and b;
    layer0_outputs(1848) <= not a;
    layer0_outputs(1849) <= not (a or b);
    layer0_outputs(1850) <= 1'b0;
    layer0_outputs(1851) <= not b;
    layer0_outputs(1852) <= a or b;
    layer0_outputs(1853) <= a and not b;
    layer0_outputs(1854) <= not b or a;
    layer0_outputs(1855) <= not b or a;
    layer0_outputs(1856) <= not (a and b);
    layer0_outputs(1857) <= a or b;
    layer0_outputs(1858) <= a;
    layer0_outputs(1859) <= a or b;
    layer0_outputs(1860) <= not a;
    layer0_outputs(1861) <= b;
    layer0_outputs(1862) <= not a or b;
    layer0_outputs(1863) <= not b or a;
    layer0_outputs(1864) <= a or b;
    layer0_outputs(1865) <= not b;
    layer0_outputs(1866) <= a and not b;
    layer0_outputs(1867) <= not (a xor b);
    layer0_outputs(1868) <= 1'b1;
    layer0_outputs(1869) <= 1'b0;
    layer0_outputs(1870) <= b;
    layer0_outputs(1871) <= a and not b;
    layer0_outputs(1872) <= a or b;
    layer0_outputs(1873) <= b;
    layer0_outputs(1874) <= a;
    layer0_outputs(1875) <= not (a or b);
    layer0_outputs(1876) <= not (a or b);
    layer0_outputs(1877) <= a;
    layer0_outputs(1878) <= b and not a;
    layer0_outputs(1879) <= not b;
    layer0_outputs(1880) <= not (a and b);
    layer0_outputs(1881) <= b and not a;
    layer0_outputs(1882) <= not b or a;
    layer0_outputs(1883) <= not a or b;
    layer0_outputs(1884) <= a or b;
    layer0_outputs(1885) <= not (a xor b);
    layer0_outputs(1886) <= not a;
    layer0_outputs(1887) <= a or b;
    layer0_outputs(1888) <= a;
    layer0_outputs(1889) <= not b or a;
    layer0_outputs(1890) <= a and b;
    layer0_outputs(1891) <= a;
    layer0_outputs(1892) <= a or b;
    layer0_outputs(1893) <= not b;
    layer0_outputs(1894) <= 1'b0;
    layer0_outputs(1895) <= a and not b;
    layer0_outputs(1896) <= not (a and b);
    layer0_outputs(1897) <= not (a or b);
    layer0_outputs(1898) <= not (a xor b);
    layer0_outputs(1899) <= a;
    layer0_outputs(1900) <= a or b;
    layer0_outputs(1901) <= a and not b;
    layer0_outputs(1902) <= a or b;
    layer0_outputs(1903) <= a;
    layer0_outputs(1904) <= b and not a;
    layer0_outputs(1905) <= a;
    layer0_outputs(1906) <= a xor b;
    layer0_outputs(1907) <= 1'b1;
    layer0_outputs(1908) <= not (a xor b);
    layer0_outputs(1909) <= not (a xor b);
    layer0_outputs(1910) <= b;
    layer0_outputs(1911) <= not (a and b);
    layer0_outputs(1912) <= b and not a;
    layer0_outputs(1913) <= a or b;
    layer0_outputs(1914) <= a xor b;
    layer0_outputs(1915) <= b and not a;
    layer0_outputs(1916) <= 1'b1;
    layer0_outputs(1917) <= a;
    layer0_outputs(1918) <= b and not a;
    layer0_outputs(1919) <= b and not a;
    layer0_outputs(1920) <= a or b;
    layer0_outputs(1921) <= not b or a;
    layer0_outputs(1922) <= not (a xor b);
    layer0_outputs(1923) <= not (a xor b);
    layer0_outputs(1924) <= b;
    layer0_outputs(1925) <= not b or a;
    layer0_outputs(1926) <= a and not b;
    layer0_outputs(1927) <= not a or b;
    layer0_outputs(1928) <= a or b;
    layer0_outputs(1929) <= 1'b0;
    layer0_outputs(1930) <= a and b;
    layer0_outputs(1931) <= a xor b;
    layer0_outputs(1932) <= a xor b;
    layer0_outputs(1933) <= b;
    layer0_outputs(1934) <= a or b;
    layer0_outputs(1935) <= a xor b;
    layer0_outputs(1936) <= not (a xor b);
    layer0_outputs(1937) <= a;
    layer0_outputs(1938) <= a;
    layer0_outputs(1939) <= a;
    layer0_outputs(1940) <= a;
    layer0_outputs(1941) <= a;
    layer0_outputs(1942) <= a;
    layer0_outputs(1943) <= not (a xor b);
    layer0_outputs(1944) <= b;
    layer0_outputs(1945) <= a and not b;
    layer0_outputs(1946) <= a xor b;
    layer0_outputs(1947) <= not a or b;
    layer0_outputs(1948) <= not a;
    layer0_outputs(1949) <= a and not b;
    layer0_outputs(1950) <= not (a and b);
    layer0_outputs(1951) <= not (a or b);
    layer0_outputs(1952) <= not a;
    layer0_outputs(1953) <= a;
    layer0_outputs(1954) <= b and not a;
    layer0_outputs(1955) <= not a;
    layer0_outputs(1956) <= b;
    layer0_outputs(1957) <= a;
    layer0_outputs(1958) <= not (a and b);
    layer0_outputs(1959) <= b;
    layer0_outputs(1960) <= not (a and b);
    layer0_outputs(1961) <= not a;
    layer0_outputs(1962) <= not (a and b);
    layer0_outputs(1963) <= not a;
    layer0_outputs(1964) <= b;
    layer0_outputs(1965) <= a or b;
    layer0_outputs(1966) <= not a;
    layer0_outputs(1967) <= a;
    layer0_outputs(1968) <= not (a xor b);
    layer0_outputs(1969) <= not (a or b);
    layer0_outputs(1970) <= not a;
    layer0_outputs(1971) <= a xor b;
    layer0_outputs(1972) <= a;
    layer0_outputs(1973) <= not a or b;
    layer0_outputs(1974) <= a and not b;
    layer0_outputs(1975) <= not a;
    layer0_outputs(1976) <= b;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= not (a xor b);
    layer0_outputs(1979) <= a;
    layer0_outputs(1980) <= a and b;
    layer0_outputs(1981) <= not b or a;
    layer0_outputs(1982) <= b;
    layer0_outputs(1983) <= b and not a;
    layer0_outputs(1984) <= not b;
    layer0_outputs(1985) <= not (a or b);
    layer0_outputs(1986) <= 1'b0;
    layer0_outputs(1987) <= not b;
    layer0_outputs(1988) <= b;
    layer0_outputs(1989) <= 1'b1;
    layer0_outputs(1990) <= a;
    layer0_outputs(1991) <= a or b;
    layer0_outputs(1992) <= a and not b;
    layer0_outputs(1993) <= not a;
    layer0_outputs(1994) <= a and not b;
    layer0_outputs(1995) <= not (a and b);
    layer0_outputs(1996) <= not (a or b);
    layer0_outputs(1997) <= a and not b;
    layer0_outputs(1998) <= a;
    layer0_outputs(1999) <= not b or a;
    layer0_outputs(2000) <= 1'b0;
    layer0_outputs(2001) <= a or b;
    layer0_outputs(2002) <= not a;
    layer0_outputs(2003) <= a xor b;
    layer0_outputs(2004) <= not b or a;
    layer0_outputs(2005) <= b;
    layer0_outputs(2006) <= not (a xor b);
    layer0_outputs(2007) <= not (a and b);
    layer0_outputs(2008) <= not (a xor b);
    layer0_outputs(2009) <= not a or b;
    layer0_outputs(2010) <= a and b;
    layer0_outputs(2011) <= not (a or b);
    layer0_outputs(2012) <= not (a xor b);
    layer0_outputs(2013) <= not b;
    layer0_outputs(2014) <= 1'b1;
    layer0_outputs(2015) <= not (a xor b);
    layer0_outputs(2016) <= not (a xor b);
    layer0_outputs(2017) <= not b;
    layer0_outputs(2018) <= a or b;
    layer0_outputs(2019) <= 1'b0;
    layer0_outputs(2020) <= not (a xor b);
    layer0_outputs(2021) <= not (a or b);
    layer0_outputs(2022) <= not (a or b);
    layer0_outputs(2023) <= a and b;
    layer0_outputs(2024) <= not a;
    layer0_outputs(2025) <= a or b;
    layer0_outputs(2026) <= a or b;
    layer0_outputs(2027) <= not (a and b);
    layer0_outputs(2028) <= not a or b;
    layer0_outputs(2029) <= 1'b1;
    layer0_outputs(2030) <= b and not a;
    layer0_outputs(2031) <= a or b;
    layer0_outputs(2032) <= a or b;
    layer0_outputs(2033) <= b;
    layer0_outputs(2034) <= not (a xor b);
    layer0_outputs(2035) <= not (a xor b);
    layer0_outputs(2036) <= not (a or b);
    layer0_outputs(2037) <= not (a and b);
    layer0_outputs(2038) <= not b;
    layer0_outputs(2039) <= a xor b;
    layer0_outputs(2040) <= a and b;
    layer0_outputs(2041) <= not a;
    layer0_outputs(2042) <= b and not a;
    layer0_outputs(2043) <= a or b;
    layer0_outputs(2044) <= not (a and b);
    layer0_outputs(2045) <= b;
    layer0_outputs(2046) <= a;
    layer0_outputs(2047) <= not (a or b);
    layer0_outputs(2048) <= a and not b;
    layer0_outputs(2049) <= a and not b;
    layer0_outputs(2050) <= not (a or b);
    layer0_outputs(2051) <= 1'b0;
    layer0_outputs(2052) <= not (a or b);
    layer0_outputs(2053) <= not (a xor b);
    layer0_outputs(2054) <= not (a xor b);
    layer0_outputs(2055) <= not (a or b);
    layer0_outputs(2056) <= a;
    layer0_outputs(2057) <= not (a or b);
    layer0_outputs(2058) <= a or b;
    layer0_outputs(2059) <= not (a or b);
    layer0_outputs(2060) <= a and not b;
    layer0_outputs(2061) <= not a;
    layer0_outputs(2062) <= not a or b;
    layer0_outputs(2063) <= not b or a;
    layer0_outputs(2064) <= a xor b;
    layer0_outputs(2065) <= not (a xor b);
    layer0_outputs(2066) <= not b;
    layer0_outputs(2067) <= 1'b1;
    layer0_outputs(2068) <= 1'b1;
    layer0_outputs(2069) <= not (a or b);
    layer0_outputs(2070) <= not a or b;
    layer0_outputs(2071) <= 1'b1;
    layer0_outputs(2072) <= not b or a;
    layer0_outputs(2073) <= not b or a;
    layer0_outputs(2074) <= not (a and b);
    layer0_outputs(2075) <= not (a or b);
    layer0_outputs(2076) <= not b;
    layer0_outputs(2077) <= a and not b;
    layer0_outputs(2078) <= a xor b;
    layer0_outputs(2079) <= not (a or b);
    layer0_outputs(2080) <= not (a xor b);
    layer0_outputs(2081) <= a or b;
    layer0_outputs(2082) <= not a;
    layer0_outputs(2083) <= not (a or b);
    layer0_outputs(2084) <= not b;
    layer0_outputs(2085) <= a or b;
    layer0_outputs(2086) <= not b;
    layer0_outputs(2087) <= not a;
    layer0_outputs(2088) <= b and not a;
    layer0_outputs(2089) <= a or b;
    layer0_outputs(2090) <= not b;
    layer0_outputs(2091) <= b;
    layer0_outputs(2092) <= a xor b;
    layer0_outputs(2093) <= a;
    layer0_outputs(2094) <= a and not b;
    layer0_outputs(2095) <= not (a or b);
    layer0_outputs(2096) <= a;
    layer0_outputs(2097) <= a and not b;
    layer0_outputs(2098) <= not b;
    layer0_outputs(2099) <= 1'b0;
    layer0_outputs(2100) <= b and not a;
    layer0_outputs(2101) <= a and not b;
    layer0_outputs(2102) <= a and not b;
    layer0_outputs(2103) <= not (a xor b);
    layer0_outputs(2104) <= not a;
    layer0_outputs(2105) <= a or b;
    layer0_outputs(2106) <= not (a or b);
    layer0_outputs(2107) <= a and b;
    layer0_outputs(2108) <= a or b;
    layer0_outputs(2109) <= 1'b0;
    layer0_outputs(2110) <= not a;
    layer0_outputs(2111) <= not a or b;
    layer0_outputs(2112) <= 1'b1;
    layer0_outputs(2113) <= not (a and b);
    layer0_outputs(2114) <= not a or b;
    layer0_outputs(2115) <= not a;
    layer0_outputs(2116) <= not (a or b);
    layer0_outputs(2117) <= not b;
    layer0_outputs(2118) <= b and not a;
    layer0_outputs(2119) <= 1'b1;
    layer0_outputs(2120) <= not a;
    layer0_outputs(2121) <= a or b;
    layer0_outputs(2122) <= not a;
    layer0_outputs(2123) <= not (a xor b);
    layer0_outputs(2124) <= not b or a;
    layer0_outputs(2125) <= not (a or b);
    layer0_outputs(2126) <= not b or a;
    layer0_outputs(2127) <= not (a or b);
    layer0_outputs(2128) <= not (a and b);
    layer0_outputs(2129) <= a and not b;
    layer0_outputs(2130) <= not (a or b);
    layer0_outputs(2131) <= not (a and b);
    layer0_outputs(2132) <= b and not a;
    layer0_outputs(2133) <= not b;
    layer0_outputs(2134) <= a or b;
    layer0_outputs(2135) <= a and b;
    layer0_outputs(2136) <= not b;
    layer0_outputs(2137) <= not (a or b);
    layer0_outputs(2138) <= a and not b;
    layer0_outputs(2139) <= b and not a;
    layer0_outputs(2140) <= not a;
    layer0_outputs(2141) <= not (a or b);
    layer0_outputs(2142) <= not (a and b);
    layer0_outputs(2143) <= not b;
    layer0_outputs(2144) <= b and not a;
    layer0_outputs(2145) <= 1'b0;
    layer0_outputs(2146) <= a xor b;
    layer0_outputs(2147) <= not a;
    layer0_outputs(2148) <= a or b;
    layer0_outputs(2149) <= b and not a;
    layer0_outputs(2150) <= not (a or b);
    layer0_outputs(2151) <= not (a or b);
    layer0_outputs(2152) <= not a;
    layer0_outputs(2153) <= a or b;
    layer0_outputs(2154) <= b and not a;
    layer0_outputs(2155) <= b and not a;
    layer0_outputs(2156) <= 1'b1;
    layer0_outputs(2157) <= b and not a;
    layer0_outputs(2158) <= not b;
    layer0_outputs(2159) <= not a or b;
    layer0_outputs(2160) <= a or b;
    layer0_outputs(2161) <= not (a or b);
    layer0_outputs(2162) <= not a;
    layer0_outputs(2163) <= not b;
    layer0_outputs(2164) <= a and not b;
    layer0_outputs(2165) <= not (a xor b);
    layer0_outputs(2166) <= a and not b;
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= a;
    layer0_outputs(2169) <= b and not a;
    layer0_outputs(2170) <= not b;
    layer0_outputs(2171) <= not (a xor b);
    layer0_outputs(2172) <= 1'b1;
    layer0_outputs(2173) <= b;
    layer0_outputs(2174) <= b;
    layer0_outputs(2175) <= not (a or b);
    layer0_outputs(2176) <= not (a xor b);
    layer0_outputs(2177) <= b;
    layer0_outputs(2178) <= a or b;
    layer0_outputs(2179) <= not (a and b);
    layer0_outputs(2180) <= a or b;
    layer0_outputs(2181) <= a and b;
    layer0_outputs(2182) <= not b;
    layer0_outputs(2183) <= not a or b;
    layer0_outputs(2184) <= not (a or b);
    layer0_outputs(2185) <= not (a or b);
    layer0_outputs(2186) <= a and not b;
    layer0_outputs(2187) <= a and b;
    layer0_outputs(2188) <= not a or b;
    layer0_outputs(2189) <= a;
    layer0_outputs(2190) <= a;
    layer0_outputs(2191) <= b and not a;
    layer0_outputs(2192) <= b;
    layer0_outputs(2193) <= a and not b;
    layer0_outputs(2194) <= b;
    layer0_outputs(2195) <= not (a or b);
    layer0_outputs(2196) <= a or b;
    layer0_outputs(2197) <= not a;
    layer0_outputs(2198) <= a and b;
    layer0_outputs(2199) <= a;
    layer0_outputs(2200) <= not (a xor b);
    layer0_outputs(2201) <= a and b;
    layer0_outputs(2202) <= a and b;
    layer0_outputs(2203) <= not (a xor b);
    layer0_outputs(2204) <= a or b;
    layer0_outputs(2205) <= not (a or b);
    layer0_outputs(2206) <= a and not b;
    layer0_outputs(2207) <= not (a or b);
    layer0_outputs(2208) <= a or b;
    layer0_outputs(2209) <= b and not a;
    layer0_outputs(2210) <= a;
    layer0_outputs(2211) <= not a;
    layer0_outputs(2212) <= a or b;
    layer0_outputs(2213) <= b and not a;
    layer0_outputs(2214) <= a xor b;
    layer0_outputs(2215) <= 1'b1;
    layer0_outputs(2216) <= not (a or b);
    layer0_outputs(2217) <= b and not a;
    layer0_outputs(2218) <= not b or a;
    layer0_outputs(2219) <= not (a and b);
    layer0_outputs(2220) <= b;
    layer0_outputs(2221) <= a;
    layer0_outputs(2222) <= a;
    layer0_outputs(2223) <= a or b;
    layer0_outputs(2224) <= 1'b0;
    layer0_outputs(2225) <= a xor b;
    layer0_outputs(2226) <= b;
    layer0_outputs(2227) <= not a or b;
    layer0_outputs(2228) <= not (a xor b);
    layer0_outputs(2229) <= a and b;
    layer0_outputs(2230) <= not (a or b);
    layer0_outputs(2231) <= a and not b;
    layer0_outputs(2232) <= not b or a;
    layer0_outputs(2233) <= not a or b;
    layer0_outputs(2234) <= 1'b1;
    layer0_outputs(2235) <= a or b;
    layer0_outputs(2236) <= 1'b0;
    layer0_outputs(2237) <= a and b;
    layer0_outputs(2238) <= not b or a;
    layer0_outputs(2239) <= not (a xor b);
    layer0_outputs(2240) <= not a;
    layer0_outputs(2241) <= not (a or b);
    layer0_outputs(2242) <= 1'b1;
    layer0_outputs(2243) <= b;
    layer0_outputs(2244) <= a or b;
    layer0_outputs(2245) <= a or b;
    layer0_outputs(2246) <= not a or b;
    layer0_outputs(2247) <= not (a or b);
    layer0_outputs(2248) <= b;
    layer0_outputs(2249) <= not b;
    layer0_outputs(2250) <= a;
    layer0_outputs(2251) <= a or b;
    layer0_outputs(2252) <= not a;
    layer0_outputs(2253) <= not (a and b);
    layer0_outputs(2254) <= not a or b;
    layer0_outputs(2255) <= a xor b;
    layer0_outputs(2256) <= a or b;
    layer0_outputs(2257) <= not a or b;
    layer0_outputs(2258) <= not a;
    layer0_outputs(2259) <= not a or b;
    layer0_outputs(2260) <= a;
    layer0_outputs(2261) <= a and not b;
    layer0_outputs(2262) <= a or b;
    layer0_outputs(2263) <= a and not b;
    layer0_outputs(2264) <= a or b;
    layer0_outputs(2265) <= a xor b;
    layer0_outputs(2266) <= a;
    layer0_outputs(2267) <= b and not a;
    layer0_outputs(2268) <= not b or a;
    layer0_outputs(2269) <= 1'b0;
    layer0_outputs(2270) <= not (a xor b);
    layer0_outputs(2271) <= 1'b0;
    layer0_outputs(2272) <= a or b;
    layer0_outputs(2273) <= b;
    layer0_outputs(2274) <= not a;
    layer0_outputs(2275) <= a and not b;
    layer0_outputs(2276) <= a;
    layer0_outputs(2277) <= b;
    layer0_outputs(2278) <= not b or a;
    layer0_outputs(2279) <= a and b;
    layer0_outputs(2280) <= a or b;
    layer0_outputs(2281) <= not a;
    layer0_outputs(2282) <= a or b;
    layer0_outputs(2283) <= 1'b1;
    layer0_outputs(2284) <= not b;
    layer0_outputs(2285) <= a or b;
    layer0_outputs(2286) <= a;
    layer0_outputs(2287) <= not a;
    layer0_outputs(2288) <= 1'b1;
    layer0_outputs(2289) <= a and not b;
    layer0_outputs(2290) <= not a or b;
    layer0_outputs(2291) <= a;
    layer0_outputs(2292) <= a;
    layer0_outputs(2293) <= b;
    layer0_outputs(2294) <= not (a and b);
    layer0_outputs(2295) <= b and not a;
    layer0_outputs(2296) <= 1'b0;
    layer0_outputs(2297) <= not (a xor b);
    layer0_outputs(2298) <= a;
    layer0_outputs(2299) <= a;
    layer0_outputs(2300) <= not a or b;
    layer0_outputs(2301) <= a or b;
    layer0_outputs(2302) <= not a;
    layer0_outputs(2303) <= not a;
    layer0_outputs(2304) <= a and b;
    layer0_outputs(2305) <= not a or b;
    layer0_outputs(2306) <= b and not a;
    layer0_outputs(2307) <= a xor b;
    layer0_outputs(2308) <= a or b;
    layer0_outputs(2309) <= not b or a;
    layer0_outputs(2310) <= b and not a;
    layer0_outputs(2311) <= a or b;
    layer0_outputs(2312) <= b;
    layer0_outputs(2313) <= a or b;
    layer0_outputs(2314) <= not a or b;
    layer0_outputs(2315) <= not a;
    layer0_outputs(2316) <= not b;
    layer0_outputs(2317) <= not b or a;
    layer0_outputs(2318) <= not (a xor b);
    layer0_outputs(2319) <= a and not b;
    layer0_outputs(2320) <= b and not a;
    layer0_outputs(2321) <= 1'b0;
    layer0_outputs(2322) <= not b or a;
    layer0_outputs(2323) <= a and b;
    layer0_outputs(2324) <= not a or b;
    layer0_outputs(2325) <= a or b;
    layer0_outputs(2326) <= a and not b;
    layer0_outputs(2327) <= not (a or b);
    layer0_outputs(2328) <= not (a or b);
    layer0_outputs(2329) <= not b or a;
    layer0_outputs(2330) <= b;
    layer0_outputs(2331) <= 1'b1;
    layer0_outputs(2332) <= not a;
    layer0_outputs(2333) <= 1'b0;
    layer0_outputs(2334) <= b;
    layer0_outputs(2335) <= not b;
    layer0_outputs(2336) <= 1'b0;
    layer0_outputs(2337) <= not (a and b);
    layer0_outputs(2338) <= not a;
    layer0_outputs(2339) <= a and not b;
    layer0_outputs(2340) <= not a;
    layer0_outputs(2341) <= not (a and b);
    layer0_outputs(2342) <= a and not b;
    layer0_outputs(2343) <= a;
    layer0_outputs(2344) <= not a or b;
    layer0_outputs(2345) <= 1'b0;
    layer0_outputs(2346) <= not a;
    layer0_outputs(2347) <= a and b;
    layer0_outputs(2348) <= b;
    layer0_outputs(2349) <= not a;
    layer0_outputs(2350) <= not (a or b);
    layer0_outputs(2351) <= b;
    layer0_outputs(2352) <= b and not a;
    layer0_outputs(2353) <= a;
    layer0_outputs(2354) <= not (a xor b);
    layer0_outputs(2355) <= not (a and b);
    layer0_outputs(2356) <= a and not b;
    layer0_outputs(2357) <= a or b;
    layer0_outputs(2358) <= b;
    layer0_outputs(2359) <= b;
    layer0_outputs(2360) <= not (a or b);
    layer0_outputs(2361) <= not b or a;
    layer0_outputs(2362) <= not b or a;
    layer0_outputs(2363) <= a or b;
    layer0_outputs(2364) <= not (a xor b);
    layer0_outputs(2365) <= 1'b1;
    layer0_outputs(2366) <= a and b;
    layer0_outputs(2367) <= not a;
    layer0_outputs(2368) <= a;
    layer0_outputs(2369) <= a xor b;
    layer0_outputs(2370) <= a and b;
    layer0_outputs(2371) <= not (a xor b);
    layer0_outputs(2372) <= a;
    layer0_outputs(2373) <= not a;
    layer0_outputs(2374) <= not (a or b);
    layer0_outputs(2375) <= a and not b;
    layer0_outputs(2376) <= not b;
    layer0_outputs(2377) <= a xor b;
    layer0_outputs(2378) <= a xor b;
    layer0_outputs(2379) <= not a or b;
    layer0_outputs(2380) <= a and b;
    layer0_outputs(2381) <= not a;
    layer0_outputs(2382) <= a xor b;
    layer0_outputs(2383) <= b and not a;
    layer0_outputs(2384) <= a or b;
    layer0_outputs(2385) <= not b;
    layer0_outputs(2386) <= a;
    layer0_outputs(2387) <= a;
    layer0_outputs(2388) <= not b;
    layer0_outputs(2389) <= b and not a;
    layer0_outputs(2390) <= a or b;
    layer0_outputs(2391) <= not b or a;
    layer0_outputs(2392) <= not a;
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= not a or b;
    layer0_outputs(2395) <= a and not b;
    layer0_outputs(2396) <= a or b;
    layer0_outputs(2397) <= a and b;
    layer0_outputs(2398) <= a xor b;
    layer0_outputs(2399) <= a;
    layer0_outputs(2400) <= a and not b;
    layer0_outputs(2401) <= a or b;
    layer0_outputs(2402) <= b and not a;
    layer0_outputs(2403) <= not b or a;
    layer0_outputs(2404) <= not a;
    layer0_outputs(2405) <= 1'b0;
    layer0_outputs(2406) <= a or b;
    layer0_outputs(2407) <= b;
    layer0_outputs(2408) <= a and b;
    layer0_outputs(2409) <= a and not b;
    layer0_outputs(2410) <= a xor b;
    layer0_outputs(2411) <= not (a or b);
    layer0_outputs(2412) <= 1'b0;
    layer0_outputs(2413) <= a xor b;
    layer0_outputs(2414) <= a;
    layer0_outputs(2415) <= a and not b;
    layer0_outputs(2416) <= a xor b;
    layer0_outputs(2417) <= 1'b0;
    layer0_outputs(2418) <= a;
    layer0_outputs(2419) <= 1'b1;
    layer0_outputs(2420) <= a or b;
    layer0_outputs(2421) <= a;
    layer0_outputs(2422) <= not a;
    layer0_outputs(2423) <= not a;
    layer0_outputs(2424) <= not a or b;
    layer0_outputs(2425) <= a;
    layer0_outputs(2426) <= not (a or b);
    layer0_outputs(2427) <= a xor b;
    layer0_outputs(2428) <= a and not b;
    layer0_outputs(2429) <= a or b;
    layer0_outputs(2430) <= not a or b;
    layer0_outputs(2431) <= b;
    layer0_outputs(2432) <= 1'b0;
    layer0_outputs(2433) <= b and not a;
    layer0_outputs(2434) <= not b;
    layer0_outputs(2435) <= not a;
    layer0_outputs(2436) <= not a;
    layer0_outputs(2437) <= a;
    layer0_outputs(2438) <= not (a or b);
    layer0_outputs(2439) <= not a or b;
    layer0_outputs(2440) <= not (a or b);
    layer0_outputs(2441) <= not a;
    layer0_outputs(2442) <= not (a or b);
    layer0_outputs(2443) <= a and b;
    layer0_outputs(2444) <= a or b;
    layer0_outputs(2445) <= a xor b;
    layer0_outputs(2446) <= not a;
    layer0_outputs(2447) <= not (a and b);
    layer0_outputs(2448) <= a xor b;
    layer0_outputs(2449) <= a xor b;
    layer0_outputs(2450) <= a;
    layer0_outputs(2451) <= not (a xor b);
    layer0_outputs(2452) <= not a;
    layer0_outputs(2453) <= not (a or b);
    layer0_outputs(2454) <= a;
    layer0_outputs(2455) <= not (a and b);
    layer0_outputs(2456) <= not a;
    layer0_outputs(2457) <= not (a xor b);
    layer0_outputs(2458) <= not b;
    layer0_outputs(2459) <= not (a or b);
    layer0_outputs(2460) <= 1'b0;
    layer0_outputs(2461) <= not (a xor b);
    layer0_outputs(2462) <= b;
    layer0_outputs(2463) <= b;
    layer0_outputs(2464) <= a or b;
    layer0_outputs(2465) <= a and not b;
    layer0_outputs(2466) <= a;
    layer0_outputs(2467) <= not b;
    layer0_outputs(2468) <= a;
    layer0_outputs(2469) <= a or b;
    layer0_outputs(2470) <= not a or b;
    layer0_outputs(2471) <= b;
    layer0_outputs(2472) <= b and not a;
    layer0_outputs(2473) <= a;
    layer0_outputs(2474) <= not (a or b);
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= not (a or b);
    layer0_outputs(2477) <= a or b;
    layer0_outputs(2478) <= not (a or b);
    layer0_outputs(2479) <= not b;
    layer0_outputs(2480) <= b and not a;
    layer0_outputs(2481) <= not a or b;
    layer0_outputs(2482) <= a;
    layer0_outputs(2483) <= not b;
    layer0_outputs(2484) <= not (a and b);
    layer0_outputs(2485) <= not (a xor b);
    layer0_outputs(2486) <= not b;
    layer0_outputs(2487) <= not a or b;
    layer0_outputs(2488) <= a or b;
    layer0_outputs(2489) <= a;
    layer0_outputs(2490) <= not a or b;
    layer0_outputs(2491) <= b and not a;
    layer0_outputs(2492) <= b and not a;
    layer0_outputs(2493) <= a and b;
    layer0_outputs(2494) <= a;
    layer0_outputs(2495) <= a or b;
    layer0_outputs(2496) <= not (a or b);
    layer0_outputs(2497) <= not (a or b);
    layer0_outputs(2498) <= a xor b;
    layer0_outputs(2499) <= not b;
    layer0_outputs(2500) <= b and not a;
    layer0_outputs(2501) <= not a;
    layer0_outputs(2502) <= a or b;
    layer0_outputs(2503) <= a xor b;
    layer0_outputs(2504) <= a or b;
    layer0_outputs(2505) <= not b or a;
    layer0_outputs(2506) <= a and b;
    layer0_outputs(2507) <= not (a or b);
    layer0_outputs(2508) <= a and not b;
    layer0_outputs(2509) <= a and b;
    layer0_outputs(2510) <= not a;
    layer0_outputs(2511) <= b and not a;
    layer0_outputs(2512) <= not a;
    layer0_outputs(2513) <= a or b;
    layer0_outputs(2514) <= b;
    layer0_outputs(2515) <= not (a or b);
    layer0_outputs(2516) <= not b;
    layer0_outputs(2517) <= not b;
    layer0_outputs(2518) <= not (a xor b);
    layer0_outputs(2519) <= not a;
    layer0_outputs(2520) <= not (a xor b);
    layer0_outputs(2521) <= not b or a;
    layer0_outputs(2522) <= a and not b;
    layer0_outputs(2523) <= not b;
    layer0_outputs(2524) <= not (a xor b);
    layer0_outputs(2525) <= not (a or b);
    layer0_outputs(2526) <= 1'b1;
    layer0_outputs(2527) <= not b;
    layer0_outputs(2528) <= 1'b0;
    layer0_outputs(2529) <= not b;
    layer0_outputs(2530) <= not (a and b);
    layer0_outputs(2531) <= a;
    layer0_outputs(2532) <= not b;
    layer0_outputs(2533) <= not (a or b);
    layer0_outputs(2534) <= a;
    layer0_outputs(2535) <= a or b;
    layer0_outputs(2536) <= not a or b;
    layer0_outputs(2537) <= not (a or b);
    layer0_outputs(2538) <= not b or a;
    layer0_outputs(2539) <= a and not b;
    layer0_outputs(2540) <= b;
    layer0_outputs(2541) <= not (a or b);
    layer0_outputs(2542) <= not b;
    layer0_outputs(2543) <= a or b;
    layer0_outputs(2544) <= not b or a;
    layer0_outputs(2545) <= b and not a;
    layer0_outputs(2546) <= a;
    layer0_outputs(2547) <= a xor b;
    layer0_outputs(2548) <= not (a xor b);
    layer0_outputs(2549) <= a and b;
    layer0_outputs(2550) <= b;
    layer0_outputs(2551) <= b and not a;
    layer0_outputs(2552) <= not (a xor b);
    layer0_outputs(2553) <= a or b;
    layer0_outputs(2554) <= not a;
    layer0_outputs(2555) <= not (a or b);
    layer0_outputs(2556) <= a or b;
    layer0_outputs(2557) <= not (a or b);
    layer0_outputs(2558) <= not a or b;
    layer0_outputs(2559) <= a;
    layer1_outputs(0) <= not a;
    layer1_outputs(1) <= a or b;
    layer1_outputs(2) <= a and not b;
    layer1_outputs(3) <= a and b;
    layer1_outputs(4) <= a and not b;
    layer1_outputs(5) <= a and b;
    layer1_outputs(6) <= not (a and b);
    layer1_outputs(7) <= not b or a;
    layer1_outputs(8) <= not (a xor b);
    layer1_outputs(9) <= a and not b;
    layer1_outputs(10) <= not a;
    layer1_outputs(11) <= not a or b;
    layer1_outputs(12) <= not b or a;
    layer1_outputs(13) <= not a or b;
    layer1_outputs(14) <= b;
    layer1_outputs(15) <= b;
    layer1_outputs(16) <= not (a and b);
    layer1_outputs(17) <= not b or a;
    layer1_outputs(18) <= a and b;
    layer1_outputs(19) <= 1'b0;
    layer1_outputs(20) <= a and b;
    layer1_outputs(21) <= a and not b;
    layer1_outputs(22) <= a and not b;
    layer1_outputs(23) <= a and b;
    layer1_outputs(24) <= a xor b;
    layer1_outputs(25) <= a and b;
    layer1_outputs(26) <= a;
    layer1_outputs(27) <= not a;
    layer1_outputs(28) <= not b;
    layer1_outputs(29) <= b;
    layer1_outputs(30) <= not (a and b);
    layer1_outputs(31) <= not a or b;
    layer1_outputs(32) <= not (a or b);
    layer1_outputs(33) <= not a or b;
    layer1_outputs(34) <= not a or b;
    layer1_outputs(35) <= not a;
    layer1_outputs(36) <= not a;
    layer1_outputs(37) <= a;
    layer1_outputs(38) <= not a or b;
    layer1_outputs(39) <= not a or b;
    layer1_outputs(40) <= b and not a;
    layer1_outputs(41) <= a and b;
    layer1_outputs(42) <= not b;
    layer1_outputs(43) <= a and not b;
    layer1_outputs(44) <= a and b;
    layer1_outputs(45) <= b;
    layer1_outputs(46) <= 1'b1;
    layer1_outputs(47) <= not a or b;
    layer1_outputs(48) <= a or b;
    layer1_outputs(49) <= a and not b;
    layer1_outputs(50) <= not (a and b);
    layer1_outputs(51) <= b and not a;
    layer1_outputs(52) <= not b;
    layer1_outputs(53) <= b;
    layer1_outputs(54) <= not (a and b);
    layer1_outputs(55) <= 1'b1;
    layer1_outputs(56) <= a or b;
    layer1_outputs(57) <= not (a xor b);
    layer1_outputs(58) <= 1'b1;
    layer1_outputs(59) <= a or b;
    layer1_outputs(60) <= a xor b;
    layer1_outputs(61) <= 1'b1;
    layer1_outputs(62) <= b;
    layer1_outputs(63) <= not a or b;
    layer1_outputs(64) <= not b or a;
    layer1_outputs(65) <= a xor b;
    layer1_outputs(66) <= a or b;
    layer1_outputs(67) <= b and not a;
    layer1_outputs(68) <= not (a or b);
    layer1_outputs(69) <= not (a xor b);
    layer1_outputs(70) <= a;
    layer1_outputs(71) <= b;
    layer1_outputs(72) <= not b or a;
    layer1_outputs(73) <= b and not a;
    layer1_outputs(74) <= not (a and b);
    layer1_outputs(75) <= not a;
    layer1_outputs(76) <= a or b;
    layer1_outputs(77) <= not b or a;
    layer1_outputs(78) <= not (a or b);
    layer1_outputs(79) <= not b;
    layer1_outputs(80) <= a;
    layer1_outputs(81) <= not (a and b);
    layer1_outputs(82) <= not a;
    layer1_outputs(83) <= not (a or b);
    layer1_outputs(84) <= b and not a;
    layer1_outputs(85) <= a and not b;
    layer1_outputs(86) <= 1'b0;
    layer1_outputs(87) <= a;
    layer1_outputs(88) <= b and not a;
    layer1_outputs(89) <= a and not b;
    layer1_outputs(90) <= not (a xor b);
    layer1_outputs(91) <= b and not a;
    layer1_outputs(92) <= a xor b;
    layer1_outputs(93) <= not (a or b);
    layer1_outputs(94) <= a;
    layer1_outputs(95) <= not a or b;
    layer1_outputs(96) <= b and not a;
    layer1_outputs(97) <= a or b;
    layer1_outputs(98) <= not (a or b);
    layer1_outputs(99) <= a;
    layer1_outputs(100) <= not a or b;
    layer1_outputs(101) <= not (a or b);
    layer1_outputs(102) <= not b or a;
    layer1_outputs(103) <= not (a xor b);
    layer1_outputs(104) <= a and not b;
    layer1_outputs(105) <= a and not b;
    layer1_outputs(106) <= a or b;
    layer1_outputs(107) <= a;
    layer1_outputs(108) <= a or b;
    layer1_outputs(109) <= not a;
    layer1_outputs(110) <= not b;
    layer1_outputs(111) <= not (a and b);
    layer1_outputs(112) <= 1'b0;
    layer1_outputs(113) <= not b;
    layer1_outputs(114) <= not b or a;
    layer1_outputs(115) <= a and not b;
    layer1_outputs(116) <= b;
    layer1_outputs(117) <= a and b;
    layer1_outputs(118) <= a;
    layer1_outputs(119) <= b;
    layer1_outputs(120) <= a and not b;
    layer1_outputs(121) <= a;
    layer1_outputs(122) <= not a;
    layer1_outputs(123) <= b;
    layer1_outputs(124) <= not a;
    layer1_outputs(125) <= a xor b;
    layer1_outputs(126) <= not a;
    layer1_outputs(127) <= a and b;
    layer1_outputs(128) <= not (a or b);
    layer1_outputs(129) <= a or b;
    layer1_outputs(130) <= 1'b0;
    layer1_outputs(131) <= not b;
    layer1_outputs(132) <= not b or a;
    layer1_outputs(133) <= not a or b;
    layer1_outputs(134) <= not a or b;
    layer1_outputs(135) <= b and not a;
    layer1_outputs(136) <= not a;
    layer1_outputs(137) <= b;
    layer1_outputs(138) <= a or b;
    layer1_outputs(139) <= a and b;
    layer1_outputs(140) <= not (a or b);
    layer1_outputs(141) <= not a or b;
    layer1_outputs(142) <= not b;
    layer1_outputs(143) <= not (a and b);
    layer1_outputs(144) <= not (a and b);
    layer1_outputs(145) <= not (a and b);
    layer1_outputs(146) <= not (a and b);
    layer1_outputs(147) <= not (a or b);
    layer1_outputs(148) <= not b;
    layer1_outputs(149) <= not (a or b);
    layer1_outputs(150) <= a and not b;
    layer1_outputs(151) <= not a;
    layer1_outputs(152) <= b and not a;
    layer1_outputs(153) <= not (a xor b);
    layer1_outputs(154) <= not a or b;
    layer1_outputs(155) <= a and b;
    layer1_outputs(156) <= not a;
    layer1_outputs(157) <= b;
    layer1_outputs(158) <= not b or a;
    layer1_outputs(159) <= not a;
    layer1_outputs(160) <= not b;
    layer1_outputs(161) <= a or b;
    layer1_outputs(162) <= b;
    layer1_outputs(163) <= not (a or b);
    layer1_outputs(164) <= b;
    layer1_outputs(165) <= not (a xor b);
    layer1_outputs(166) <= not (a or b);
    layer1_outputs(167) <= 1'b1;
    layer1_outputs(168) <= not a;
    layer1_outputs(169) <= a and b;
    layer1_outputs(170) <= a and b;
    layer1_outputs(171) <= not a;
    layer1_outputs(172) <= a and not b;
    layer1_outputs(173) <= b and not a;
    layer1_outputs(174) <= 1'b1;
    layer1_outputs(175) <= a and not b;
    layer1_outputs(176) <= not (a and b);
    layer1_outputs(177) <= b;
    layer1_outputs(178) <= not (a and b);
    layer1_outputs(179) <= not b;
    layer1_outputs(180) <= a xor b;
    layer1_outputs(181) <= not a;
    layer1_outputs(182) <= not b or a;
    layer1_outputs(183) <= 1'b1;
    layer1_outputs(184) <= a or b;
    layer1_outputs(185) <= not b;
    layer1_outputs(186) <= a;
    layer1_outputs(187) <= a and not b;
    layer1_outputs(188) <= not (a or b);
    layer1_outputs(189) <= b;
    layer1_outputs(190) <= b and not a;
    layer1_outputs(191) <= a and not b;
    layer1_outputs(192) <= b;
    layer1_outputs(193) <= not b or a;
    layer1_outputs(194) <= b;
    layer1_outputs(195) <= not b;
    layer1_outputs(196) <= a and not b;
    layer1_outputs(197) <= 1'b0;
    layer1_outputs(198) <= b and not a;
    layer1_outputs(199) <= a;
    layer1_outputs(200) <= 1'b0;
    layer1_outputs(201) <= a and not b;
    layer1_outputs(202) <= 1'b1;
    layer1_outputs(203) <= 1'b0;
    layer1_outputs(204) <= not a or b;
    layer1_outputs(205) <= a and b;
    layer1_outputs(206) <= 1'b1;
    layer1_outputs(207) <= a or b;
    layer1_outputs(208) <= not b;
    layer1_outputs(209) <= not b or a;
    layer1_outputs(210) <= not a or b;
    layer1_outputs(211) <= a;
    layer1_outputs(212) <= a or b;
    layer1_outputs(213) <= a or b;
    layer1_outputs(214) <= 1'b1;
    layer1_outputs(215) <= not (a xor b);
    layer1_outputs(216) <= a or b;
    layer1_outputs(217) <= not a or b;
    layer1_outputs(218) <= not a or b;
    layer1_outputs(219) <= a and not b;
    layer1_outputs(220) <= not b;
    layer1_outputs(221) <= 1'b0;
    layer1_outputs(222) <= not (a or b);
    layer1_outputs(223) <= 1'b1;
    layer1_outputs(224) <= a and not b;
    layer1_outputs(225) <= a;
    layer1_outputs(226) <= a;
    layer1_outputs(227) <= a or b;
    layer1_outputs(228) <= a;
    layer1_outputs(229) <= not a or b;
    layer1_outputs(230) <= a xor b;
    layer1_outputs(231) <= not b;
    layer1_outputs(232) <= not (a or b);
    layer1_outputs(233) <= b;
    layer1_outputs(234) <= b;
    layer1_outputs(235) <= not b or a;
    layer1_outputs(236) <= b;
    layer1_outputs(237) <= a;
    layer1_outputs(238) <= not b;
    layer1_outputs(239) <= b and not a;
    layer1_outputs(240) <= 1'b1;
    layer1_outputs(241) <= a and not b;
    layer1_outputs(242) <= b;
    layer1_outputs(243) <= not b;
    layer1_outputs(244) <= not (a xor b);
    layer1_outputs(245) <= b;
    layer1_outputs(246) <= not (a and b);
    layer1_outputs(247) <= not a;
    layer1_outputs(248) <= not a or b;
    layer1_outputs(249) <= a;
    layer1_outputs(250) <= not a;
    layer1_outputs(251) <= a and b;
    layer1_outputs(252) <= not a or b;
    layer1_outputs(253) <= a;
    layer1_outputs(254) <= not b;
    layer1_outputs(255) <= not a;
    layer1_outputs(256) <= not b or a;
    layer1_outputs(257) <= a and not b;
    layer1_outputs(258) <= not b;
    layer1_outputs(259) <= not b or a;
    layer1_outputs(260) <= not (a and b);
    layer1_outputs(261) <= b and not a;
    layer1_outputs(262) <= a or b;
    layer1_outputs(263) <= not (a or b);
    layer1_outputs(264) <= a or b;
    layer1_outputs(265) <= a and not b;
    layer1_outputs(266) <= a or b;
    layer1_outputs(267) <= not a;
    layer1_outputs(268) <= not (a xor b);
    layer1_outputs(269) <= a and not b;
    layer1_outputs(270) <= b;
    layer1_outputs(271) <= not (a and b);
    layer1_outputs(272) <= b and not a;
    layer1_outputs(273) <= b;
    layer1_outputs(274) <= a;
    layer1_outputs(275) <= b;
    layer1_outputs(276) <= not a;
    layer1_outputs(277) <= not a or b;
    layer1_outputs(278) <= a and not b;
    layer1_outputs(279) <= not b or a;
    layer1_outputs(280) <= a;
    layer1_outputs(281) <= not (a xor b);
    layer1_outputs(282) <= b;
    layer1_outputs(283) <= b;
    layer1_outputs(284) <= not (a xor b);
    layer1_outputs(285) <= a;
    layer1_outputs(286) <= not a;
    layer1_outputs(287) <= b;
    layer1_outputs(288) <= not b or a;
    layer1_outputs(289) <= 1'b1;
    layer1_outputs(290) <= b;
    layer1_outputs(291) <= b and not a;
    layer1_outputs(292) <= a;
    layer1_outputs(293) <= b;
    layer1_outputs(294) <= not a or b;
    layer1_outputs(295) <= not a;
    layer1_outputs(296) <= a or b;
    layer1_outputs(297) <= a xor b;
    layer1_outputs(298) <= not b or a;
    layer1_outputs(299) <= not b;
    layer1_outputs(300) <= not a;
    layer1_outputs(301) <= b and not a;
    layer1_outputs(302) <= not (a and b);
    layer1_outputs(303) <= not b;
    layer1_outputs(304) <= 1'b0;
    layer1_outputs(305) <= not a;
    layer1_outputs(306) <= a;
    layer1_outputs(307) <= b and not a;
    layer1_outputs(308) <= not b or a;
    layer1_outputs(309) <= not a or b;
    layer1_outputs(310) <= not b or a;
    layer1_outputs(311) <= a or b;
    layer1_outputs(312) <= b and not a;
    layer1_outputs(313) <= not b or a;
    layer1_outputs(314) <= 1'b0;
    layer1_outputs(315) <= a and not b;
    layer1_outputs(316) <= not a or b;
    layer1_outputs(317) <= not (a or b);
    layer1_outputs(318) <= b and not a;
    layer1_outputs(319) <= a;
    layer1_outputs(320) <= a and b;
    layer1_outputs(321) <= a;
    layer1_outputs(322) <= not a;
    layer1_outputs(323) <= not (a or b);
    layer1_outputs(324) <= not b or a;
    layer1_outputs(325) <= a and b;
    layer1_outputs(326) <= a xor b;
    layer1_outputs(327) <= b and not a;
    layer1_outputs(328) <= b and not a;
    layer1_outputs(329) <= not b;
    layer1_outputs(330) <= a;
    layer1_outputs(331) <= 1'b1;
    layer1_outputs(332) <= b and not a;
    layer1_outputs(333) <= b and not a;
    layer1_outputs(334) <= not (a and b);
    layer1_outputs(335) <= a;
    layer1_outputs(336) <= 1'b0;
    layer1_outputs(337) <= not a;
    layer1_outputs(338) <= 1'b1;
    layer1_outputs(339) <= not (a and b);
    layer1_outputs(340) <= 1'b1;
    layer1_outputs(341) <= b and not a;
    layer1_outputs(342) <= b and not a;
    layer1_outputs(343) <= not b or a;
    layer1_outputs(344) <= a and b;
    layer1_outputs(345) <= a and not b;
    layer1_outputs(346) <= not a;
    layer1_outputs(347) <= a or b;
    layer1_outputs(348) <= a xor b;
    layer1_outputs(349) <= not a or b;
    layer1_outputs(350) <= b and not a;
    layer1_outputs(351) <= not a or b;
    layer1_outputs(352) <= not a or b;
    layer1_outputs(353) <= a;
    layer1_outputs(354) <= not b;
    layer1_outputs(355) <= a and b;
    layer1_outputs(356) <= a;
    layer1_outputs(357) <= not (a or b);
    layer1_outputs(358) <= a and not b;
    layer1_outputs(359) <= b and not a;
    layer1_outputs(360) <= 1'b0;
    layer1_outputs(361) <= 1'b1;
    layer1_outputs(362) <= 1'b1;
    layer1_outputs(363) <= not b or a;
    layer1_outputs(364) <= not (a and b);
    layer1_outputs(365) <= a xor b;
    layer1_outputs(366) <= a and b;
    layer1_outputs(367) <= not (a and b);
    layer1_outputs(368) <= not (a and b);
    layer1_outputs(369) <= not (a and b);
    layer1_outputs(370) <= not a or b;
    layer1_outputs(371) <= not b;
    layer1_outputs(372) <= a;
    layer1_outputs(373) <= b;
    layer1_outputs(374) <= not b;
    layer1_outputs(375) <= b;
    layer1_outputs(376) <= not a or b;
    layer1_outputs(377) <= a;
    layer1_outputs(378) <= not b;
    layer1_outputs(379) <= not (a and b);
    layer1_outputs(380) <= not (a and b);
    layer1_outputs(381) <= not (a and b);
    layer1_outputs(382) <= a;
    layer1_outputs(383) <= a and not b;
    layer1_outputs(384) <= not a or b;
    layer1_outputs(385) <= a;
    layer1_outputs(386) <= a and b;
    layer1_outputs(387) <= not b;
    layer1_outputs(388) <= a or b;
    layer1_outputs(389) <= a;
    layer1_outputs(390) <= a or b;
    layer1_outputs(391) <= 1'b1;
    layer1_outputs(392) <= a;
    layer1_outputs(393) <= a xor b;
    layer1_outputs(394) <= a and b;
    layer1_outputs(395) <= not a or b;
    layer1_outputs(396) <= not b or a;
    layer1_outputs(397) <= not a or b;
    layer1_outputs(398) <= b;
    layer1_outputs(399) <= not a;
    layer1_outputs(400) <= a;
    layer1_outputs(401) <= a;
    layer1_outputs(402) <= b and not a;
    layer1_outputs(403) <= b and not a;
    layer1_outputs(404) <= b;
    layer1_outputs(405) <= not (a or b);
    layer1_outputs(406) <= not a;
    layer1_outputs(407) <= b and not a;
    layer1_outputs(408) <= not b;
    layer1_outputs(409) <= not b or a;
    layer1_outputs(410) <= not b;
    layer1_outputs(411) <= a;
    layer1_outputs(412) <= a;
    layer1_outputs(413) <= not (a and b);
    layer1_outputs(414) <= b;
    layer1_outputs(415) <= a;
    layer1_outputs(416) <= not a or b;
    layer1_outputs(417) <= 1'b1;
    layer1_outputs(418) <= a;
    layer1_outputs(419) <= a and not b;
    layer1_outputs(420) <= b;
    layer1_outputs(421) <= not b;
    layer1_outputs(422) <= not (a and b);
    layer1_outputs(423) <= a and b;
    layer1_outputs(424) <= not (a xor b);
    layer1_outputs(425) <= not b or a;
    layer1_outputs(426) <= not (a or b);
    layer1_outputs(427) <= not (a or b);
    layer1_outputs(428) <= b;
    layer1_outputs(429) <= a;
    layer1_outputs(430) <= 1'b1;
    layer1_outputs(431) <= a and not b;
    layer1_outputs(432) <= not b;
    layer1_outputs(433) <= not b;
    layer1_outputs(434) <= not b;
    layer1_outputs(435) <= not b or a;
    layer1_outputs(436) <= not a or b;
    layer1_outputs(437) <= not a;
    layer1_outputs(438) <= a;
    layer1_outputs(439) <= a and b;
    layer1_outputs(440) <= b;
    layer1_outputs(441) <= not a;
    layer1_outputs(442) <= 1'b0;
    layer1_outputs(443) <= a or b;
    layer1_outputs(444) <= a xor b;
    layer1_outputs(445) <= a;
    layer1_outputs(446) <= a and not b;
    layer1_outputs(447) <= b;
    layer1_outputs(448) <= a xor b;
    layer1_outputs(449) <= 1'b1;
    layer1_outputs(450) <= 1'b1;
    layer1_outputs(451) <= b;
    layer1_outputs(452) <= 1'b0;
    layer1_outputs(453) <= a;
    layer1_outputs(454) <= not b;
    layer1_outputs(455) <= not (a or b);
    layer1_outputs(456) <= 1'b0;
    layer1_outputs(457) <= b and not a;
    layer1_outputs(458) <= not b;
    layer1_outputs(459) <= b and not a;
    layer1_outputs(460) <= not b;
    layer1_outputs(461) <= not (a or b);
    layer1_outputs(462) <= not b;
    layer1_outputs(463) <= 1'b1;
    layer1_outputs(464) <= a xor b;
    layer1_outputs(465) <= a or b;
    layer1_outputs(466) <= b and not a;
    layer1_outputs(467) <= not b or a;
    layer1_outputs(468) <= 1'b0;
    layer1_outputs(469) <= a xor b;
    layer1_outputs(470) <= b and not a;
    layer1_outputs(471) <= b and not a;
    layer1_outputs(472) <= b and not a;
    layer1_outputs(473) <= a xor b;
    layer1_outputs(474) <= 1'b1;
    layer1_outputs(475) <= not b;
    layer1_outputs(476) <= a or b;
    layer1_outputs(477) <= a and not b;
    layer1_outputs(478) <= not a;
    layer1_outputs(479) <= not b;
    layer1_outputs(480) <= not (a or b);
    layer1_outputs(481) <= not a or b;
    layer1_outputs(482) <= a;
    layer1_outputs(483) <= not a;
    layer1_outputs(484) <= a and not b;
    layer1_outputs(485) <= a and b;
    layer1_outputs(486) <= a;
    layer1_outputs(487) <= not (a or b);
    layer1_outputs(488) <= b and not a;
    layer1_outputs(489) <= not a;
    layer1_outputs(490) <= 1'b1;
    layer1_outputs(491) <= not b;
    layer1_outputs(492) <= not b or a;
    layer1_outputs(493) <= a;
    layer1_outputs(494) <= not (a or b);
    layer1_outputs(495) <= not a or b;
    layer1_outputs(496) <= a and b;
    layer1_outputs(497) <= 1'b1;
    layer1_outputs(498) <= b and not a;
    layer1_outputs(499) <= not a or b;
    layer1_outputs(500) <= not b;
    layer1_outputs(501) <= not b or a;
    layer1_outputs(502) <= not (a or b);
    layer1_outputs(503) <= a and not b;
    layer1_outputs(504) <= not (a or b);
    layer1_outputs(505) <= a or b;
    layer1_outputs(506) <= a and not b;
    layer1_outputs(507) <= not a;
    layer1_outputs(508) <= a;
    layer1_outputs(509) <= not a or b;
    layer1_outputs(510) <= a;
    layer1_outputs(511) <= not a or b;
    layer1_outputs(512) <= a or b;
    layer1_outputs(513) <= b and not a;
    layer1_outputs(514) <= a and not b;
    layer1_outputs(515) <= not (a xor b);
    layer1_outputs(516) <= a or b;
    layer1_outputs(517) <= not (a or b);
    layer1_outputs(518) <= a or b;
    layer1_outputs(519) <= 1'b1;
    layer1_outputs(520) <= not (a or b);
    layer1_outputs(521) <= not b;
    layer1_outputs(522) <= b;
    layer1_outputs(523) <= a or b;
    layer1_outputs(524) <= not b or a;
    layer1_outputs(525) <= not b;
    layer1_outputs(526) <= 1'b0;
    layer1_outputs(527) <= not (a and b);
    layer1_outputs(528) <= b and not a;
    layer1_outputs(529) <= a or b;
    layer1_outputs(530) <= a or b;
    layer1_outputs(531) <= b and not a;
    layer1_outputs(532) <= b and not a;
    layer1_outputs(533) <= b;
    layer1_outputs(534) <= not (a or b);
    layer1_outputs(535) <= not (a or b);
    layer1_outputs(536) <= not (a or b);
    layer1_outputs(537) <= not a or b;
    layer1_outputs(538) <= not a or b;
    layer1_outputs(539) <= a or b;
    layer1_outputs(540) <= not (a and b);
    layer1_outputs(541) <= a and b;
    layer1_outputs(542) <= a and not b;
    layer1_outputs(543) <= not a;
    layer1_outputs(544) <= a or b;
    layer1_outputs(545) <= b and not a;
    layer1_outputs(546) <= b;
    layer1_outputs(547) <= not (a and b);
    layer1_outputs(548) <= b;
    layer1_outputs(549) <= b and not a;
    layer1_outputs(550) <= b and not a;
    layer1_outputs(551) <= not (a and b);
    layer1_outputs(552) <= not a or b;
    layer1_outputs(553) <= not b or a;
    layer1_outputs(554) <= not b;
    layer1_outputs(555) <= not (a or b);
    layer1_outputs(556) <= a and not b;
    layer1_outputs(557) <= b;
    layer1_outputs(558) <= not a or b;
    layer1_outputs(559) <= not (a or b);
    layer1_outputs(560) <= a and not b;
    layer1_outputs(561) <= not (a or b);
    layer1_outputs(562) <= b;
    layer1_outputs(563) <= not (a or b);
    layer1_outputs(564) <= a or b;
    layer1_outputs(565) <= a;
    layer1_outputs(566) <= a;
    layer1_outputs(567) <= a or b;
    layer1_outputs(568) <= 1'b0;
    layer1_outputs(569) <= not (a or b);
    layer1_outputs(570) <= a and b;
    layer1_outputs(571) <= b and not a;
    layer1_outputs(572) <= not a or b;
    layer1_outputs(573) <= a or b;
    layer1_outputs(574) <= not b;
    layer1_outputs(575) <= not a;
    layer1_outputs(576) <= not (a and b);
    layer1_outputs(577) <= a and b;
    layer1_outputs(578) <= not b;
    layer1_outputs(579) <= not b;
    layer1_outputs(580) <= not (a and b);
    layer1_outputs(581) <= 1'b1;
    layer1_outputs(582) <= not (a and b);
    layer1_outputs(583) <= a;
    layer1_outputs(584) <= not a;
    layer1_outputs(585) <= not (a or b);
    layer1_outputs(586) <= b and not a;
    layer1_outputs(587) <= not (a and b);
    layer1_outputs(588) <= a or b;
    layer1_outputs(589) <= not a;
    layer1_outputs(590) <= not a or b;
    layer1_outputs(591) <= not a or b;
    layer1_outputs(592) <= 1'b0;
    layer1_outputs(593) <= a or b;
    layer1_outputs(594) <= 1'b1;
    layer1_outputs(595) <= 1'b0;
    layer1_outputs(596) <= not b;
    layer1_outputs(597) <= b and not a;
    layer1_outputs(598) <= not b;
    layer1_outputs(599) <= not (a and b);
    layer1_outputs(600) <= not b or a;
    layer1_outputs(601) <= not b;
    layer1_outputs(602) <= not b;
    layer1_outputs(603) <= not b or a;
    layer1_outputs(604) <= not (a or b);
    layer1_outputs(605) <= a and b;
    layer1_outputs(606) <= not b or a;
    layer1_outputs(607) <= not a;
    layer1_outputs(608) <= not b or a;
    layer1_outputs(609) <= b;
    layer1_outputs(610) <= not b or a;
    layer1_outputs(611) <= 1'b1;
    layer1_outputs(612) <= 1'b0;
    layer1_outputs(613) <= a and b;
    layer1_outputs(614) <= not b or a;
    layer1_outputs(615) <= not a;
    layer1_outputs(616) <= a;
    layer1_outputs(617) <= a and not b;
    layer1_outputs(618) <= 1'b0;
    layer1_outputs(619) <= not (a xor b);
    layer1_outputs(620) <= 1'b1;
    layer1_outputs(621) <= not a or b;
    layer1_outputs(622) <= a or b;
    layer1_outputs(623) <= not a or b;
    layer1_outputs(624) <= b;
    layer1_outputs(625) <= 1'b0;
    layer1_outputs(626) <= b;
    layer1_outputs(627) <= not a;
    layer1_outputs(628) <= b;
    layer1_outputs(629) <= b;
    layer1_outputs(630) <= b;
    layer1_outputs(631) <= not b;
    layer1_outputs(632) <= a and not b;
    layer1_outputs(633) <= b;
    layer1_outputs(634) <= a;
    layer1_outputs(635) <= 1'b1;
    layer1_outputs(636) <= a or b;
    layer1_outputs(637) <= not (a and b);
    layer1_outputs(638) <= a;
    layer1_outputs(639) <= a and not b;
    layer1_outputs(640) <= not a;
    layer1_outputs(641) <= b and not a;
    layer1_outputs(642) <= not a or b;
    layer1_outputs(643) <= a;
    layer1_outputs(644) <= not (a and b);
    layer1_outputs(645) <= not a or b;
    layer1_outputs(646) <= a and not b;
    layer1_outputs(647) <= not b;
    layer1_outputs(648) <= not a;
    layer1_outputs(649) <= not (a xor b);
    layer1_outputs(650) <= a;
    layer1_outputs(651) <= b and not a;
    layer1_outputs(652) <= a;
    layer1_outputs(653) <= a and b;
    layer1_outputs(654) <= not b or a;
    layer1_outputs(655) <= not b or a;
    layer1_outputs(656) <= not (a and b);
    layer1_outputs(657) <= not (a or b);
    layer1_outputs(658) <= 1'b1;
    layer1_outputs(659) <= a and not b;
    layer1_outputs(660) <= b and not a;
    layer1_outputs(661) <= 1'b1;
    layer1_outputs(662) <= not (a or b);
    layer1_outputs(663) <= a and not b;
    layer1_outputs(664) <= b;
    layer1_outputs(665) <= 1'b0;
    layer1_outputs(666) <= not b;
    layer1_outputs(667) <= a and b;
    layer1_outputs(668) <= a and b;
    layer1_outputs(669) <= a or b;
    layer1_outputs(670) <= a and b;
    layer1_outputs(671) <= b;
    layer1_outputs(672) <= b and not a;
    layer1_outputs(673) <= b and not a;
    layer1_outputs(674) <= not b or a;
    layer1_outputs(675) <= a xor b;
    layer1_outputs(676) <= a and not b;
    layer1_outputs(677) <= not a or b;
    layer1_outputs(678) <= not a or b;
    layer1_outputs(679) <= not b;
    layer1_outputs(680) <= a;
    layer1_outputs(681) <= not (a xor b);
    layer1_outputs(682) <= 1'b1;
    layer1_outputs(683) <= a;
    layer1_outputs(684) <= not a;
    layer1_outputs(685) <= not b or a;
    layer1_outputs(686) <= a and b;
    layer1_outputs(687) <= a and not b;
    layer1_outputs(688) <= b;
    layer1_outputs(689) <= a xor b;
    layer1_outputs(690) <= not b or a;
    layer1_outputs(691) <= 1'b0;
    layer1_outputs(692) <= a and not b;
    layer1_outputs(693) <= b and not a;
    layer1_outputs(694) <= not (a or b);
    layer1_outputs(695) <= b and not a;
    layer1_outputs(696) <= a and b;
    layer1_outputs(697) <= 1'b1;
    layer1_outputs(698) <= a xor b;
    layer1_outputs(699) <= 1'b1;
    layer1_outputs(700) <= b and not a;
    layer1_outputs(701) <= b and not a;
    layer1_outputs(702) <= 1'b0;
    layer1_outputs(703) <= b;
    layer1_outputs(704) <= a;
    layer1_outputs(705) <= not (a or b);
    layer1_outputs(706) <= a and not b;
    layer1_outputs(707) <= not b or a;
    layer1_outputs(708) <= not b;
    layer1_outputs(709) <= a;
    layer1_outputs(710) <= 1'b0;
    layer1_outputs(711) <= a and b;
    layer1_outputs(712) <= a;
    layer1_outputs(713) <= not b or a;
    layer1_outputs(714) <= 1'b0;
    layer1_outputs(715) <= a;
    layer1_outputs(716) <= not a or b;
    layer1_outputs(717) <= not b;
    layer1_outputs(718) <= b and not a;
    layer1_outputs(719) <= not b or a;
    layer1_outputs(720) <= not b;
    layer1_outputs(721) <= not a;
    layer1_outputs(722) <= b;
    layer1_outputs(723) <= a or b;
    layer1_outputs(724) <= a and not b;
    layer1_outputs(725) <= a and not b;
    layer1_outputs(726) <= not (a and b);
    layer1_outputs(727) <= not (a or b);
    layer1_outputs(728) <= not a or b;
    layer1_outputs(729) <= not a;
    layer1_outputs(730) <= b;
    layer1_outputs(731) <= not b;
    layer1_outputs(732) <= a and b;
    layer1_outputs(733) <= not (a or b);
    layer1_outputs(734) <= not (a xor b);
    layer1_outputs(735) <= 1'b1;
    layer1_outputs(736) <= not b;
    layer1_outputs(737) <= a;
    layer1_outputs(738) <= not b;
    layer1_outputs(739) <= a;
    layer1_outputs(740) <= 1'b0;
    layer1_outputs(741) <= a and not b;
    layer1_outputs(742) <= a xor b;
    layer1_outputs(743) <= 1'b0;
    layer1_outputs(744) <= not a;
    layer1_outputs(745) <= not b;
    layer1_outputs(746) <= b and not a;
    layer1_outputs(747) <= not a;
    layer1_outputs(748) <= 1'b0;
    layer1_outputs(749) <= not (a and b);
    layer1_outputs(750) <= a or b;
    layer1_outputs(751) <= b and not a;
    layer1_outputs(752) <= b and not a;
    layer1_outputs(753) <= not (a and b);
    layer1_outputs(754) <= not b;
    layer1_outputs(755) <= 1'b0;
    layer1_outputs(756) <= not (a or b);
    layer1_outputs(757) <= b and not a;
    layer1_outputs(758) <= not (a xor b);
    layer1_outputs(759) <= a and b;
    layer1_outputs(760) <= a or b;
    layer1_outputs(761) <= a xor b;
    layer1_outputs(762) <= not a;
    layer1_outputs(763) <= 1'b1;
    layer1_outputs(764) <= not a;
    layer1_outputs(765) <= not a or b;
    layer1_outputs(766) <= not a;
    layer1_outputs(767) <= a;
    layer1_outputs(768) <= not (a or b);
    layer1_outputs(769) <= a and not b;
    layer1_outputs(770) <= not a;
    layer1_outputs(771) <= not b or a;
    layer1_outputs(772) <= a or b;
    layer1_outputs(773) <= b;
    layer1_outputs(774) <= a or b;
    layer1_outputs(775) <= not b or a;
    layer1_outputs(776) <= not (a and b);
    layer1_outputs(777) <= not a or b;
    layer1_outputs(778) <= not a;
    layer1_outputs(779) <= a;
    layer1_outputs(780) <= not a or b;
    layer1_outputs(781) <= not b;
    layer1_outputs(782) <= a;
    layer1_outputs(783) <= 1'b0;
    layer1_outputs(784) <= not b or a;
    layer1_outputs(785) <= not a;
    layer1_outputs(786) <= a;
    layer1_outputs(787) <= not a;
    layer1_outputs(788) <= not a;
    layer1_outputs(789) <= a or b;
    layer1_outputs(790) <= not a;
    layer1_outputs(791) <= not a;
    layer1_outputs(792) <= not (a or b);
    layer1_outputs(793) <= a xor b;
    layer1_outputs(794) <= not (a and b);
    layer1_outputs(795) <= not a;
    layer1_outputs(796) <= not (a or b);
    layer1_outputs(797) <= not a or b;
    layer1_outputs(798) <= 1'b1;
    layer1_outputs(799) <= not b;
    layer1_outputs(800) <= 1'b1;
    layer1_outputs(801) <= b and not a;
    layer1_outputs(802) <= not b or a;
    layer1_outputs(803) <= a and b;
    layer1_outputs(804) <= a and b;
    layer1_outputs(805) <= a;
    layer1_outputs(806) <= not (a or b);
    layer1_outputs(807) <= a or b;
    layer1_outputs(808) <= not a;
    layer1_outputs(809) <= not b;
    layer1_outputs(810) <= a;
    layer1_outputs(811) <= not b;
    layer1_outputs(812) <= a;
    layer1_outputs(813) <= a or b;
    layer1_outputs(814) <= b;
    layer1_outputs(815) <= not a;
    layer1_outputs(816) <= b;
    layer1_outputs(817) <= not b;
    layer1_outputs(818) <= 1'b1;
    layer1_outputs(819) <= not (a or b);
    layer1_outputs(820) <= a or b;
    layer1_outputs(821) <= a xor b;
    layer1_outputs(822) <= 1'b0;
    layer1_outputs(823) <= not b or a;
    layer1_outputs(824) <= not b;
    layer1_outputs(825) <= a and b;
    layer1_outputs(826) <= a and b;
    layer1_outputs(827) <= a;
    layer1_outputs(828) <= a;
    layer1_outputs(829) <= a and b;
    layer1_outputs(830) <= not b;
    layer1_outputs(831) <= not (a and b);
    layer1_outputs(832) <= not b;
    layer1_outputs(833) <= 1'b0;
    layer1_outputs(834) <= a;
    layer1_outputs(835) <= not (a and b);
    layer1_outputs(836) <= not b;
    layer1_outputs(837) <= a and not b;
    layer1_outputs(838) <= not b or a;
    layer1_outputs(839) <= not a or b;
    layer1_outputs(840) <= not b or a;
    layer1_outputs(841) <= a and b;
    layer1_outputs(842) <= a and b;
    layer1_outputs(843) <= b;
    layer1_outputs(844) <= b and not a;
    layer1_outputs(845) <= a;
    layer1_outputs(846) <= not a;
    layer1_outputs(847) <= a;
    layer1_outputs(848) <= not a or b;
    layer1_outputs(849) <= a;
    layer1_outputs(850) <= 1'b0;
    layer1_outputs(851) <= a and not b;
    layer1_outputs(852) <= b and not a;
    layer1_outputs(853) <= b and not a;
    layer1_outputs(854) <= not a;
    layer1_outputs(855) <= b and not a;
    layer1_outputs(856) <= a xor b;
    layer1_outputs(857) <= a;
    layer1_outputs(858) <= not (a and b);
    layer1_outputs(859) <= b and not a;
    layer1_outputs(860) <= 1'b1;
    layer1_outputs(861) <= not a;
    layer1_outputs(862) <= a xor b;
    layer1_outputs(863) <= not (a or b);
    layer1_outputs(864) <= a;
    layer1_outputs(865) <= a;
    layer1_outputs(866) <= not a;
    layer1_outputs(867) <= not (a and b);
    layer1_outputs(868) <= not b;
    layer1_outputs(869) <= a;
    layer1_outputs(870) <= not (a or b);
    layer1_outputs(871) <= not b;
    layer1_outputs(872) <= a or b;
    layer1_outputs(873) <= not b;
    layer1_outputs(874) <= b and not a;
    layer1_outputs(875) <= not (a xor b);
    layer1_outputs(876) <= 1'b0;
    layer1_outputs(877) <= not (a or b);
    layer1_outputs(878) <= a and not b;
    layer1_outputs(879) <= not b or a;
    layer1_outputs(880) <= not (a and b);
    layer1_outputs(881) <= b;
    layer1_outputs(882) <= a xor b;
    layer1_outputs(883) <= a xor b;
    layer1_outputs(884) <= not a or b;
    layer1_outputs(885) <= not a or b;
    layer1_outputs(886) <= not (a xor b);
    layer1_outputs(887) <= a and not b;
    layer1_outputs(888) <= 1'b1;
    layer1_outputs(889) <= a and not b;
    layer1_outputs(890) <= b and not a;
    layer1_outputs(891) <= a and b;
    layer1_outputs(892) <= a;
    layer1_outputs(893) <= b;
    layer1_outputs(894) <= not b or a;
    layer1_outputs(895) <= not a or b;
    layer1_outputs(896) <= not b or a;
    layer1_outputs(897) <= a xor b;
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= a;
    layer1_outputs(900) <= not (a and b);
    layer1_outputs(901) <= not a or b;
    layer1_outputs(902) <= not b;
    layer1_outputs(903) <= not (a xor b);
    layer1_outputs(904) <= not (a or b);
    layer1_outputs(905) <= 1'b1;
    layer1_outputs(906) <= not b or a;
    layer1_outputs(907) <= b;
    layer1_outputs(908) <= not a or b;
    layer1_outputs(909) <= b;
    layer1_outputs(910) <= 1'b1;
    layer1_outputs(911) <= not a or b;
    layer1_outputs(912) <= b;
    layer1_outputs(913) <= not b or a;
    layer1_outputs(914) <= a and b;
    layer1_outputs(915) <= not (a xor b);
    layer1_outputs(916) <= b;
    layer1_outputs(917) <= a or b;
    layer1_outputs(918) <= b;
    layer1_outputs(919) <= not (a and b);
    layer1_outputs(920) <= a or b;
    layer1_outputs(921) <= 1'b0;
    layer1_outputs(922) <= not (a and b);
    layer1_outputs(923) <= b;
    layer1_outputs(924) <= not a;
    layer1_outputs(925) <= 1'b0;
    layer1_outputs(926) <= not b or a;
    layer1_outputs(927) <= not b;
    layer1_outputs(928) <= a or b;
    layer1_outputs(929) <= not a;
    layer1_outputs(930) <= a and b;
    layer1_outputs(931) <= a;
    layer1_outputs(932) <= not a or b;
    layer1_outputs(933) <= not b or a;
    layer1_outputs(934) <= not b or a;
    layer1_outputs(935) <= not (a and b);
    layer1_outputs(936) <= not (a and b);
    layer1_outputs(937) <= 1'b0;
    layer1_outputs(938) <= not b;
    layer1_outputs(939) <= 1'b1;
    layer1_outputs(940) <= not a;
    layer1_outputs(941) <= not (a and b);
    layer1_outputs(942) <= a;
    layer1_outputs(943) <= not (a and b);
    layer1_outputs(944) <= a;
    layer1_outputs(945) <= not a;
    layer1_outputs(946) <= a or b;
    layer1_outputs(947) <= not a or b;
    layer1_outputs(948) <= not (a and b);
    layer1_outputs(949) <= a and not b;
    layer1_outputs(950) <= a;
    layer1_outputs(951) <= a;
    layer1_outputs(952) <= not b or a;
    layer1_outputs(953) <= a and b;
    layer1_outputs(954) <= not (a xor b);
    layer1_outputs(955) <= not (a or b);
    layer1_outputs(956) <= not b;
    layer1_outputs(957) <= 1'b0;
    layer1_outputs(958) <= not a;
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= a;
    layer1_outputs(961) <= not (a and b);
    layer1_outputs(962) <= not b or a;
    layer1_outputs(963) <= not a or b;
    layer1_outputs(964) <= a and b;
    layer1_outputs(965) <= a and b;
    layer1_outputs(966) <= not b or a;
    layer1_outputs(967) <= not a;
    layer1_outputs(968) <= a and not b;
    layer1_outputs(969) <= a and not b;
    layer1_outputs(970) <= a xor b;
    layer1_outputs(971) <= not (a or b);
    layer1_outputs(972) <= a and b;
    layer1_outputs(973) <= 1'b1;
    layer1_outputs(974) <= a;
    layer1_outputs(975) <= not (a xor b);
    layer1_outputs(976) <= not b;
    layer1_outputs(977) <= a or b;
    layer1_outputs(978) <= a and not b;
    layer1_outputs(979) <= not a;
    layer1_outputs(980) <= 1'b1;
    layer1_outputs(981) <= a;
    layer1_outputs(982) <= a or b;
    layer1_outputs(983) <= not b;
    layer1_outputs(984) <= a;
    layer1_outputs(985) <= b;
    layer1_outputs(986) <= b;
    layer1_outputs(987) <= not b or a;
    layer1_outputs(988) <= not (a or b);
    layer1_outputs(989) <= not b or a;
    layer1_outputs(990) <= not (a xor b);
    layer1_outputs(991) <= not (a or b);
    layer1_outputs(992) <= a and b;
    layer1_outputs(993) <= a or b;
    layer1_outputs(994) <= not (a and b);
    layer1_outputs(995) <= not a;
    layer1_outputs(996) <= not b;
    layer1_outputs(997) <= not b or a;
    layer1_outputs(998) <= not b or a;
    layer1_outputs(999) <= 1'b0;
    layer1_outputs(1000) <= a and not b;
    layer1_outputs(1001) <= a xor b;
    layer1_outputs(1002) <= a and not b;
    layer1_outputs(1003) <= not (a xor b);
    layer1_outputs(1004) <= a and not b;
    layer1_outputs(1005) <= not b or a;
    layer1_outputs(1006) <= a or b;
    layer1_outputs(1007) <= not a;
    layer1_outputs(1008) <= not a;
    layer1_outputs(1009) <= 1'b0;
    layer1_outputs(1010) <= 1'b1;
    layer1_outputs(1011) <= b;
    layer1_outputs(1012) <= b;
    layer1_outputs(1013) <= a;
    layer1_outputs(1014) <= a and not b;
    layer1_outputs(1015) <= b;
    layer1_outputs(1016) <= not a or b;
    layer1_outputs(1017) <= not (a or b);
    layer1_outputs(1018) <= not a;
    layer1_outputs(1019) <= b and not a;
    layer1_outputs(1020) <= b;
    layer1_outputs(1021) <= not (a and b);
    layer1_outputs(1022) <= not a or b;
    layer1_outputs(1023) <= a;
    layer1_outputs(1024) <= b and not a;
    layer1_outputs(1025) <= a xor b;
    layer1_outputs(1026) <= b;
    layer1_outputs(1027) <= a;
    layer1_outputs(1028) <= not a;
    layer1_outputs(1029) <= not (a and b);
    layer1_outputs(1030) <= not (a or b);
    layer1_outputs(1031) <= not b;
    layer1_outputs(1032) <= not a;
    layer1_outputs(1033) <= not b;
    layer1_outputs(1034) <= not b;
    layer1_outputs(1035) <= not (a and b);
    layer1_outputs(1036) <= a and b;
    layer1_outputs(1037) <= a and b;
    layer1_outputs(1038) <= a and b;
    layer1_outputs(1039) <= a;
    layer1_outputs(1040) <= b;
    layer1_outputs(1041) <= a and b;
    layer1_outputs(1042) <= not a or b;
    layer1_outputs(1043) <= b;
    layer1_outputs(1044) <= not b or a;
    layer1_outputs(1045) <= not a;
    layer1_outputs(1046) <= b and not a;
    layer1_outputs(1047) <= not (a xor b);
    layer1_outputs(1048) <= b and not a;
    layer1_outputs(1049) <= b;
    layer1_outputs(1050) <= not (a or b);
    layer1_outputs(1051) <= a and b;
    layer1_outputs(1052) <= not b;
    layer1_outputs(1053) <= a and b;
    layer1_outputs(1054) <= not (a or b);
    layer1_outputs(1055) <= not b or a;
    layer1_outputs(1056) <= 1'b0;
    layer1_outputs(1057) <= not a;
    layer1_outputs(1058) <= 1'b0;
    layer1_outputs(1059) <= not a or b;
    layer1_outputs(1060) <= not b;
    layer1_outputs(1061) <= a;
    layer1_outputs(1062) <= not b or a;
    layer1_outputs(1063) <= not (a or b);
    layer1_outputs(1064) <= 1'b1;
    layer1_outputs(1065) <= not a;
    layer1_outputs(1066) <= not a or b;
    layer1_outputs(1067) <= not (a or b);
    layer1_outputs(1068) <= not a or b;
    layer1_outputs(1069) <= b;
    layer1_outputs(1070) <= a and not b;
    layer1_outputs(1071) <= not b;
    layer1_outputs(1072) <= 1'b1;
    layer1_outputs(1073) <= a and b;
    layer1_outputs(1074) <= b and not a;
    layer1_outputs(1075) <= a;
    layer1_outputs(1076) <= b;
    layer1_outputs(1077) <= b;
    layer1_outputs(1078) <= 1'b1;
    layer1_outputs(1079) <= not a;
    layer1_outputs(1080) <= not b or a;
    layer1_outputs(1081) <= not a;
    layer1_outputs(1082) <= not a;
    layer1_outputs(1083) <= b and not a;
    layer1_outputs(1084) <= a and b;
    layer1_outputs(1085) <= a and not b;
    layer1_outputs(1086) <= not a or b;
    layer1_outputs(1087) <= b and not a;
    layer1_outputs(1088) <= not a;
    layer1_outputs(1089) <= not (a and b);
    layer1_outputs(1090) <= a and b;
    layer1_outputs(1091) <= a xor b;
    layer1_outputs(1092) <= not (a or b);
    layer1_outputs(1093) <= a xor b;
    layer1_outputs(1094) <= a;
    layer1_outputs(1095) <= not (a xor b);
    layer1_outputs(1096) <= 1'b0;
    layer1_outputs(1097) <= 1'b1;
    layer1_outputs(1098) <= not (a or b);
    layer1_outputs(1099) <= not (a and b);
    layer1_outputs(1100) <= a or b;
    layer1_outputs(1101) <= 1'b1;
    layer1_outputs(1102) <= 1'b1;
    layer1_outputs(1103) <= b;
    layer1_outputs(1104) <= not b;
    layer1_outputs(1105) <= a;
    layer1_outputs(1106) <= not (a xor b);
    layer1_outputs(1107) <= 1'b0;
    layer1_outputs(1108) <= a or b;
    layer1_outputs(1109) <= not (a or b);
    layer1_outputs(1110) <= a and b;
    layer1_outputs(1111) <= not b or a;
    layer1_outputs(1112) <= a xor b;
    layer1_outputs(1113) <= not (a xor b);
    layer1_outputs(1114) <= not a;
    layer1_outputs(1115) <= not a or b;
    layer1_outputs(1116) <= not (a and b);
    layer1_outputs(1117) <= a;
    layer1_outputs(1118) <= a and b;
    layer1_outputs(1119) <= a and not b;
    layer1_outputs(1120) <= not b or a;
    layer1_outputs(1121) <= b;
    layer1_outputs(1122) <= b;
    layer1_outputs(1123) <= a;
    layer1_outputs(1124) <= 1'b1;
    layer1_outputs(1125) <= not (a or b);
    layer1_outputs(1126) <= not a;
    layer1_outputs(1127) <= 1'b1;
    layer1_outputs(1128) <= a or b;
    layer1_outputs(1129) <= b and not a;
    layer1_outputs(1130) <= a and b;
    layer1_outputs(1131) <= a or b;
    layer1_outputs(1132) <= a or b;
    layer1_outputs(1133) <= not (a or b);
    layer1_outputs(1134) <= a;
    layer1_outputs(1135) <= not a or b;
    layer1_outputs(1136) <= a;
    layer1_outputs(1137) <= not b;
    layer1_outputs(1138) <= 1'b1;
    layer1_outputs(1139) <= not a;
    layer1_outputs(1140) <= not (a or b);
    layer1_outputs(1141) <= a and b;
    layer1_outputs(1142) <= a xor b;
    layer1_outputs(1143) <= not a;
    layer1_outputs(1144) <= not a or b;
    layer1_outputs(1145) <= b;
    layer1_outputs(1146) <= not a;
    layer1_outputs(1147) <= a and not b;
    layer1_outputs(1148) <= not (a or b);
    layer1_outputs(1149) <= not b;
    layer1_outputs(1150) <= b and not a;
    layer1_outputs(1151) <= a and b;
    layer1_outputs(1152) <= not (a and b);
    layer1_outputs(1153) <= b;
    layer1_outputs(1154) <= not a;
    layer1_outputs(1155) <= not a or b;
    layer1_outputs(1156) <= a and b;
    layer1_outputs(1157) <= not a;
    layer1_outputs(1158) <= not a or b;
    layer1_outputs(1159) <= not a;
    layer1_outputs(1160) <= 1'b0;
    layer1_outputs(1161) <= a;
    layer1_outputs(1162) <= a and b;
    layer1_outputs(1163) <= b;
    layer1_outputs(1164) <= a;
    layer1_outputs(1165) <= not (a or b);
    layer1_outputs(1166) <= not a;
    layer1_outputs(1167) <= 1'b0;
    layer1_outputs(1168) <= a;
    layer1_outputs(1169) <= 1'b0;
    layer1_outputs(1170) <= not (a or b);
    layer1_outputs(1171) <= a or b;
    layer1_outputs(1172) <= not a;
    layer1_outputs(1173) <= a;
    layer1_outputs(1174) <= not (a or b);
    layer1_outputs(1175) <= a and b;
    layer1_outputs(1176) <= not (a and b);
    layer1_outputs(1177) <= not (a and b);
    layer1_outputs(1178) <= not a;
    layer1_outputs(1179) <= not b;
    layer1_outputs(1180) <= not a;
    layer1_outputs(1181) <= not b or a;
    layer1_outputs(1182) <= b and not a;
    layer1_outputs(1183) <= a or b;
    layer1_outputs(1184) <= a and b;
    layer1_outputs(1185) <= b;
    layer1_outputs(1186) <= not b;
    layer1_outputs(1187) <= b and not a;
    layer1_outputs(1188) <= not a;
    layer1_outputs(1189) <= not b or a;
    layer1_outputs(1190) <= not b or a;
    layer1_outputs(1191) <= b;
    layer1_outputs(1192) <= a or b;
    layer1_outputs(1193) <= not a;
    layer1_outputs(1194) <= b;
    layer1_outputs(1195) <= not (a or b);
    layer1_outputs(1196) <= not b;
    layer1_outputs(1197) <= not (a or b);
    layer1_outputs(1198) <= b;
    layer1_outputs(1199) <= a and not b;
    layer1_outputs(1200) <= not (a and b);
    layer1_outputs(1201) <= not (a and b);
    layer1_outputs(1202) <= a and not b;
    layer1_outputs(1203) <= a xor b;
    layer1_outputs(1204) <= not b;
    layer1_outputs(1205) <= b;
    layer1_outputs(1206) <= b;
    layer1_outputs(1207) <= not b or a;
    layer1_outputs(1208) <= a or b;
    layer1_outputs(1209) <= 1'b1;
    layer1_outputs(1210) <= not (a or b);
    layer1_outputs(1211) <= b;
    layer1_outputs(1212) <= a or b;
    layer1_outputs(1213) <= a and not b;
    layer1_outputs(1214) <= not (a or b);
    layer1_outputs(1215) <= a and b;
    layer1_outputs(1216) <= not b;
    layer1_outputs(1217) <= a and not b;
    layer1_outputs(1218) <= 1'b1;
    layer1_outputs(1219) <= b and not a;
    layer1_outputs(1220) <= not a or b;
    layer1_outputs(1221) <= not b;
    layer1_outputs(1222) <= b;
    layer1_outputs(1223) <= 1'b0;
    layer1_outputs(1224) <= not a or b;
    layer1_outputs(1225) <= a;
    layer1_outputs(1226) <= not (a or b);
    layer1_outputs(1227) <= not b or a;
    layer1_outputs(1228) <= a;
    layer1_outputs(1229) <= not a;
    layer1_outputs(1230) <= not (a and b);
    layer1_outputs(1231) <= not b or a;
    layer1_outputs(1232) <= not (a xor b);
    layer1_outputs(1233) <= b and not a;
    layer1_outputs(1234) <= not b;
    layer1_outputs(1235) <= not (a xor b);
    layer1_outputs(1236) <= a xor b;
    layer1_outputs(1237) <= a and not b;
    layer1_outputs(1238) <= not a;
    layer1_outputs(1239) <= a and b;
    layer1_outputs(1240) <= 1'b0;
    layer1_outputs(1241) <= b;
    layer1_outputs(1242) <= not a;
    layer1_outputs(1243) <= a xor b;
    layer1_outputs(1244) <= not (a and b);
    layer1_outputs(1245) <= not a;
    layer1_outputs(1246) <= a;
    layer1_outputs(1247) <= not b or a;
    layer1_outputs(1248) <= 1'b1;
    layer1_outputs(1249) <= not b;
    layer1_outputs(1250) <= not a or b;
    layer1_outputs(1251) <= not (a and b);
    layer1_outputs(1252) <= not a or b;
    layer1_outputs(1253) <= not (a and b);
    layer1_outputs(1254) <= not (a or b);
    layer1_outputs(1255) <= a and not b;
    layer1_outputs(1256) <= not (a and b);
    layer1_outputs(1257) <= not (a or b);
    layer1_outputs(1258) <= not a;
    layer1_outputs(1259) <= not (a and b);
    layer1_outputs(1260) <= a and b;
    layer1_outputs(1261) <= not (a and b);
    layer1_outputs(1262) <= not (a or b);
    layer1_outputs(1263) <= 1'b1;
    layer1_outputs(1264) <= a and b;
    layer1_outputs(1265) <= a and b;
    layer1_outputs(1266) <= a xor b;
    layer1_outputs(1267) <= a and b;
    layer1_outputs(1268) <= not (a xor b);
    layer1_outputs(1269) <= not b;
    layer1_outputs(1270) <= not a or b;
    layer1_outputs(1271) <= 1'b1;
    layer1_outputs(1272) <= not (a xor b);
    layer1_outputs(1273) <= b;
    layer1_outputs(1274) <= not a;
    layer1_outputs(1275) <= not b;
    layer1_outputs(1276) <= not b;
    layer1_outputs(1277) <= b;
    layer1_outputs(1278) <= b and not a;
    layer1_outputs(1279) <= not a;
    layer1_outputs(1280) <= not (a and b);
    layer1_outputs(1281) <= 1'b0;
    layer1_outputs(1282) <= not b;
    layer1_outputs(1283) <= a;
    layer1_outputs(1284) <= not a;
    layer1_outputs(1285) <= 1'b0;
    layer1_outputs(1286) <= not b;
    layer1_outputs(1287) <= not (a or b);
    layer1_outputs(1288) <= not (a or b);
    layer1_outputs(1289) <= not a;
    layer1_outputs(1290) <= 1'b0;
    layer1_outputs(1291) <= a or b;
    layer1_outputs(1292) <= not (a or b);
    layer1_outputs(1293) <= not (a or b);
    layer1_outputs(1294) <= not (a xor b);
    layer1_outputs(1295) <= b;
    layer1_outputs(1296) <= not b;
    layer1_outputs(1297) <= a and b;
    layer1_outputs(1298) <= a xor b;
    layer1_outputs(1299) <= not a or b;
    layer1_outputs(1300) <= not (a and b);
    layer1_outputs(1301) <= not (a and b);
    layer1_outputs(1302) <= a and b;
    layer1_outputs(1303) <= b and not a;
    layer1_outputs(1304) <= b and not a;
    layer1_outputs(1305) <= not (a or b);
    layer1_outputs(1306) <= a xor b;
    layer1_outputs(1307) <= b and not a;
    layer1_outputs(1308) <= not a or b;
    layer1_outputs(1309) <= b;
    layer1_outputs(1310) <= a;
    layer1_outputs(1311) <= not (a or b);
    layer1_outputs(1312) <= not a;
    layer1_outputs(1313) <= not a;
    layer1_outputs(1314) <= not a;
    layer1_outputs(1315) <= not b;
    layer1_outputs(1316) <= a;
    layer1_outputs(1317) <= not (a xor b);
    layer1_outputs(1318) <= not b or a;
    layer1_outputs(1319) <= not (a xor b);
    layer1_outputs(1320) <= not a;
    layer1_outputs(1321) <= not b;
    layer1_outputs(1322) <= not a;
    layer1_outputs(1323) <= a and not b;
    layer1_outputs(1324) <= not a or b;
    layer1_outputs(1325) <= a or b;
    layer1_outputs(1326) <= b;
    layer1_outputs(1327) <= not a;
    layer1_outputs(1328) <= not b;
    layer1_outputs(1329) <= a and not b;
    layer1_outputs(1330) <= a or b;
    layer1_outputs(1331) <= not (a and b);
    layer1_outputs(1332) <= not a;
    layer1_outputs(1333) <= not a;
    layer1_outputs(1334) <= a;
    layer1_outputs(1335) <= b and not a;
    layer1_outputs(1336) <= a;
    layer1_outputs(1337) <= not (a and b);
    layer1_outputs(1338) <= not b or a;
    layer1_outputs(1339) <= not a;
    layer1_outputs(1340) <= b and not a;
    layer1_outputs(1341) <= a and not b;
    layer1_outputs(1342) <= not (a or b);
    layer1_outputs(1343) <= b;
    layer1_outputs(1344) <= not b;
    layer1_outputs(1345) <= not b;
    layer1_outputs(1346) <= a;
    layer1_outputs(1347) <= a or b;
    layer1_outputs(1348) <= a and not b;
    layer1_outputs(1349) <= a;
    layer1_outputs(1350) <= a and b;
    layer1_outputs(1351) <= not (a and b);
    layer1_outputs(1352) <= not b;
    layer1_outputs(1353) <= not (a and b);
    layer1_outputs(1354) <= b;
    layer1_outputs(1355) <= a and b;
    layer1_outputs(1356) <= not b;
    layer1_outputs(1357) <= 1'b1;
    layer1_outputs(1358) <= not a or b;
    layer1_outputs(1359) <= not b or a;
    layer1_outputs(1360) <= a xor b;
    layer1_outputs(1361) <= not (a or b);
    layer1_outputs(1362) <= not (a and b);
    layer1_outputs(1363) <= a or b;
    layer1_outputs(1364) <= a and b;
    layer1_outputs(1365) <= not b;
    layer1_outputs(1366) <= b and not a;
    layer1_outputs(1367) <= not b or a;
    layer1_outputs(1368) <= a or b;
    layer1_outputs(1369) <= not b or a;
    layer1_outputs(1370) <= not b or a;
    layer1_outputs(1371) <= a and b;
    layer1_outputs(1372) <= not (a or b);
    layer1_outputs(1373) <= b and not a;
    layer1_outputs(1374) <= not (a or b);
    layer1_outputs(1375) <= 1'b0;
    layer1_outputs(1376) <= not (a and b);
    layer1_outputs(1377) <= not (a and b);
    layer1_outputs(1378) <= 1'b0;
    layer1_outputs(1379) <= 1'b0;
    layer1_outputs(1380) <= not a or b;
    layer1_outputs(1381) <= not b or a;
    layer1_outputs(1382) <= a and not b;
    layer1_outputs(1383) <= not (a xor b);
    layer1_outputs(1384) <= b;
    layer1_outputs(1385) <= not b;
    layer1_outputs(1386) <= not (a xor b);
    layer1_outputs(1387) <= a and not b;
    layer1_outputs(1388) <= not b;
    layer1_outputs(1389) <= b;
    layer1_outputs(1390) <= not (a and b);
    layer1_outputs(1391) <= not (a xor b);
    layer1_outputs(1392) <= not (a and b);
    layer1_outputs(1393) <= 1'b1;
    layer1_outputs(1394) <= not a;
    layer1_outputs(1395) <= not b or a;
    layer1_outputs(1396) <= b;
    layer1_outputs(1397) <= not (a and b);
    layer1_outputs(1398) <= not b;
    layer1_outputs(1399) <= 1'b0;
    layer1_outputs(1400) <= not b;
    layer1_outputs(1401) <= not b or a;
    layer1_outputs(1402) <= not a;
    layer1_outputs(1403) <= not b;
    layer1_outputs(1404) <= not a;
    layer1_outputs(1405) <= b;
    layer1_outputs(1406) <= a xor b;
    layer1_outputs(1407) <= b and not a;
    layer1_outputs(1408) <= a xor b;
    layer1_outputs(1409) <= not a;
    layer1_outputs(1410) <= b and not a;
    layer1_outputs(1411) <= 1'b0;
    layer1_outputs(1412) <= b;
    layer1_outputs(1413) <= not b;
    layer1_outputs(1414) <= b and not a;
    layer1_outputs(1415) <= not a or b;
    layer1_outputs(1416) <= a;
    layer1_outputs(1417) <= a;
    layer1_outputs(1418) <= not b;
    layer1_outputs(1419) <= not a or b;
    layer1_outputs(1420) <= b;
    layer1_outputs(1421) <= not a or b;
    layer1_outputs(1422) <= a;
    layer1_outputs(1423) <= not (a xor b);
    layer1_outputs(1424) <= a and b;
    layer1_outputs(1425) <= not a;
    layer1_outputs(1426) <= not a or b;
    layer1_outputs(1427) <= not (a and b);
    layer1_outputs(1428) <= a and not b;
    layer1_outputs(1429) <= a and b;
    layer1_outputs(1430) <= not b;
    layer1_outputs(1431) <= b and not a;
    layer1_outputs(1432) <= b and not a;
    layer1_outputs(1433) <= b and not a;
    layer1_outputs(1434) <= 1'b1;
    layer1_outputs(1435) <= b and not a;
    layer1_outputs(1436) <= b;
    layer1_outputs(1437) <= not a;
    layer1_outputs(1438) <= b and not a;
    layer1_outputs(1439) <= 1'b0;
    layer1_outputs(1440) <= 1'b0;
    layer1_outputs(1441) <= a and b;
    layer1_outputs(1442) <= not (a or b);
    layer1_outputs(1443) <= not b or a;
    layer1_outputs(1444) <= not a;
    layer1_outputs(1445) <= b and not a;
    layer1_outputs(1446) <= b;
    layer1_outputs(1447) <= not b or a;
    layer1_outputs(1448) <= not (a or b);
    layer1_outputs(1449) <= a;
    layer1_outputs(1450) <= not (a or b);
    layer1_outputs(1451) <= not b;
    layer1_outputs(1452) <= 1'b1;
    layer1_outputs(1453) <= a;
    layer1_outputs(1454) <= not b;
    layer1_outputs(1455) <= a and not b;
    layer1_outputs(1456) <= a and b;
    layer1_outputs(1457) <= b and not a;
    layer1_outputs(1458) <= not b;
    layer1_outputs(1459) <= not (a xor b);
    layer1_outputs(1460) <= a;
    layer1_outputs(1461) <= a;
    layer1_outputs(1462) <= a and not b;
    layer1_outputs(1463) <= not a;
    layer1_outputs(1464) <= not a or b;
    layer1_outputs(1465) <= a;
    layer1_outputs(1466) <= 1'b1;
    layer1_outputs(1467) <= a and b;
    layer1_outputs(1468) <= b and not a;
    layer1_outputs(1469) <= not (a and b);
    layer1_outputs(1470) <= not b or a;
    layer1_outputs(1471) <= not a;
    layer1_outputs(1472) <= a;
    layer1_outputs(1473) <= a;
    layer1_outputs(1474) <= a and not b;
    layer1_outputs(1475) <= not (a or b);
    layer1_outputs(1476) <= 1'b1;
    layer1_outputs(1477) <= a and b;
    layer1_outputs(1478) <= not (a or b);
    layer1_outputs(1479) <= not b or a;
    layer1_outputs(1480) <= a and not b;
    layer1_outputs(1481) <= not b;
    layer1_outputs(1482) <= not b;
    layer1_outputs(1483) <= a;
    layer1_outputs(1484) <= not a;
    layer1_outputs(1485) <= a or b;
    layer1_outputs(1486) <= not (a or b);
    layer1_outputs(1487) <= b and not a;
    layer1_outputs(1488) <= b;
    layer1_outputs(1489) <= b;
    layer1_outputs(1490) <= not a or b;
    layer1_outputs(1491) <= 1'b1;
    layer1_outputs(1492) <= 1'b1;
    layer1_outputs(1493) <= 1'b0;
    layer1_outputs(1494) <= b and not a;
    layer1_outputs(1495) <= b and not a;
    layer1_outputs(1496) <= 1'b0;
    layer1_outputs(1497) <= b and not a;
    layer1_outputs(1498) <= not a;
    layer1_outputs(1499) <= b;
    layer1_outputs(1500) <= 1'b0;
    layer1_outputs(1501) <= not b or a;
    layer1_outputs(1502) <= not b;
    layer1_outputs(1503) <= 1'b1;
    layer1_outputs(1504) <= b;
    layer1_outputs(1505) <= not b or a;
    layer1_outputs(1506) <= 1'b1;
    layer1_outputs(1507) <= not b;
    layer1_outputs(1508) <= a or b;
    layer1_outputs(1509) <= 1'b1;
    layer1_outputs(1510) <= a or b;
    layer1_outputs(1511) <= not b;
    layer1_outputs(1512) <= b;
    layer1_outputs(1513) <= b and not a;
    layer1_outputs(1514) <= a xor b;
    layer1_outputs(1515) <= a and b;
    layer1_outputs(1516) <= not (a and b);
    layer1_outputs(1517) <= not a;
    layer1_outputs(1518) <= 1'b1;
    layer1_outputs(1519) <= a xor b;
    layer1_outputs(1520) <= b;
    layer1_outputs(1521) <= b;
    layer1_outputs(1522) <= 1'b1;
    layer1_outputs(1523) <= not (a and b);
    layer1_outputs(1524) <= a and b;
    layer1_outputs(1525) <= 1'b1;
    layer1_outputs(1526) <= a;
    layer1_outputs(1527) <= a xor b;
    layer1_outputs(1528) <= not a or b;
    layer1_outputs(1529) <= not b;
    layer1_outputs(1530) <= 1'b0;
    layer1_outputs(1531) <= not a or b;
    layer1_outputs(1532) <= not a;
    layer1_outputs(1533) <= a and b;
    layer1_outputs(1534) <= b;
    layer1_outputs(1535) <= a or b;
    layer1_outputs(1536) <= not (a or b);
    layer1_outputs(1537) <= b;
    layer1_outputs(1538) <= not (a and b);
    layer1_outputs(1539) <= not b or a;
    layer1_outputs(1540) <= a and not b;
    layer1_outputs(1541) <= a or b;
    layer1_outputs(1542) <= a;
    layer1_outputs(1543) <= a and not b;
    layer1_outputs(1544) <= not a;
    layer1_outputs(1545) <= b;
    layer1_outputs(1546) <= 1'b0;
    layer1_outputs(1547) <= 1'b0;
    layer1_outputs(1548) <= a;
    layer1_outputs(1549) <= not a or b;
    layer1_outputs(1550) <= not a;
    layer1_outputs(1551) <= not b;
    layer1_outputs(1552) <= not (a xor b);
    layer1_outputs(1553) <= not b or a;
    layer1_outputs(1554) <= not (a or b);
    layer1_outputs(1555) <= not (a xor b);
    layer1_outputs(1556) <= a and b;
    layer1_outputs(1557) <= not b or a;
    layer1_outputs(1558) <= 1'b1;
    layer1_outputs(1559) <= b and not a;
    layer1_outputs(1560) <= a;
    layer1_outputs(1561) <= b;
    layer1_outputs(1562) <= not a;
    layer1_outputs(1563) <= a;
    layer1_outputs(1564) <= a and not b;
    layer1_outputs(1565) <= 1'b1;
    layer1_outputs(1566) <= a and not b;
    layer1_outputs(1567) <= a and not b;
    layer1_outputs(1568) <= a;
    layer1_outputs(1569) <= not (a or b);
    layer1_outputs(1570) <= 1'b0;
    layer1_outputs(1571) <= 1'b0;
    layer1_outputs(1572) <= b;
    layer1_outputs(1573) <= 1'b0;
    layer1_outputs(1574) <= not b;
    layer1_outputs(1575) <= not b;
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= 1'b1;
    layer1_outputs(1578) <= not b or a;
    layer1_outputs(1579) <= not b or a;
    layer1_outputs(1580) <= b and not a;
    layer1_outputs(1581) <= not (a or b);
    layer1_outputs(1582) <= not b;
    layer1_outputs(1583) <= b and not a;
    layer1_outputs(1584) <= not b;
    layer1_outputs(1585) <= not a;
    layer1_outputs(1586) <= a;
    layer1_outputs(1587) <= b;
    layer1_outputs(1588) <= a and not b;
    layer1_outputs(1589) <= b and not a;
    layer1_outputs(1590) <= not (a or b);
    layer1_outputs(1591) <= not b;
    layer1_outputs(1592) <= a and not b;
    layer1_outputs(1593) <= a;
    layer1_outputs(1594) <= not (a or b);
    layer1_outputs(1595) <= 1'b1;
    layer1_outputs(1596) <= not (a or b);
    layer1_outputs(1597) <= a;
    layer1_outputs(1598) <= not (a xor b);
    layer1_outputs(1599) <= b and not a;
    layer1_outputs(1600) <= not b or a;
    layer1_outputs(1601) <= not a;
    layer1_outputs(1602) <= not (a or b);
    layer1_outputs(1603) <= b;
    layer1_outputs(1604) <= a and not b;
    layer1_outputs(1605) <= not a or b;
    layer1_outputs(1606) <= a xor b;
    layer1_outputs(1607) <= not a;
    layer1_outputs(1608) <= 1'b0;
    layer1_outputs(1609) <= not b;
    layer1_outputs(1610) <= not b or a;
    layer1_outputs(1611) <= b and not a;
    layer1_outputs(1612) <= not (a and b);
    layer1_outputs(1613) <= 1'b1;
    layer1_outputs(1614) <= not (a or b);
    layer1_outputs(1615) <= a xor b;
    layer1_outputs(1616) <= not b or a;
    layer1_outputs(1617) <= b and not a;
    layer1_outputs(1618) <= not (a and b);
    layer1_outputs(1619) <= b;
    layer1_outputs(1620) <= not a;
    layer1_outputs(1621) <= not (a xor b);
    layer1_outputs(1622) <= not b;
    layer1_outputs(1623) <= not (a and b);
    layer1_outputs(1624) <= a;
    layer1_outputs(1625) <= a and not b;
    layer1_outputs(1626) <= not (a and b);
    layer1_outputs(1627) <= a;
    layer1_outputs(1628) <= not b;
    layer1_outputs(1629) <= 1'b1;
    layer1_outputs(1630) <= b;
    layer1_outputs(1631) <= not (a xor b);
    layer1_outputs(1632) <= a and not b;
    layer1_outputs(1633) <= a or b;
    layer1_outputs(1634) <= a and not b;
    layer1_outputs(1635) <= not (a and b);
    layer1_outputs(1636) <= a and not b;
    layer1_outputs(1637) <= not b;
    layer1_outputs(1638) <= not a or b;
    layer1_outputs(1639) <= not (a and b);
    layer1_outputs(1640) <= not (a and b);
    layer1_outputs(1641) <= a;
    layer1_outputs(1642) <= 1'b0;
    layer1_outputs(1643) <= b and not a;
    layer1_outputs(1644) <= not (a and b);
    layer1_outputs(1645) <= b and not a;
    layer1_outputs(1646) <= a xor b;
    layer1_outputs(1647) <= b;
    layer1_outputs(1648) <= not a or b;
    layer1_outputs(1649) <= not (a or b);
    layer1_outputs(1650) <= 1'b1;
    layer1_outputs(1651) <= not b or a;
    layer1_outputs(1652) <= a and b;
    layer1_outputs(1653) <= b and not a;
    layer1_outputs(1654) <= not b;
    layer1_outputs(1655) <= a or b;
    layer1_outputs(1656) <= a or b;
    layer1_outputs(1657) <= 1'b0;
    layer1_outputs(1658) <= not a or b;
    layer1_outputs(1659) <= not b or a;
    layer1_outputs(1660) <= not a;
    layer1_outputs(1661) <= b;
    layer1_outputs(1662) <= a;
    layer1_outputs(1663) <= b and not a;
    layer1_outputs(1664) <= a or b;
    layer1_outputs(1665) <= not a;
    layer1_outputs(1666) <= not (a and b);
    layer1_outputs(1667) <= a and b;
    layer1_outputs(1668) <= not a;
    layer1_outputs(1669) <= not b or a;
    layer1_outputs(1670) <= 1'b1;
    layer1_outputs(1671) <= not b or a;
    layer1_outputs(1672) <= not b;
    layer1_outputs(1673) <= b;
    layer1_outputs(1674) <= not a or b;
    layer1_outputs(1675) <= 1'b1;
    layer1_outputs(1676) <= not (a or b);
    layer1_outputs(1677) <= a and not b;
    layer1_outputs(1678) <= not a;
    layer1_outputs(1679) <= not b or a;
    layer1_outputs(1680) <= not (a and b);
    layer1_outputs(1681) <= not (a and b);
    layer1_outputs(1682) <= not a;
    layer1_outputs(1683) <= not b or a;
    layer1_outputs(1684) <= 1'b0;
    layer1_outputs(1685) <= not a or b;
    layer1_outputs(1686) <= a or b;
    layer1_outputs(1687) <= b;
    layer1_outputs(1688) <= not (a and b);
    layer1_outputs(1689) <= not (a and b);
    layer1_outputs(1690) <= not b or a;
    layer1_outputs(1691) <= b;
    layer1_outputs(1692) <= a and not b;
    layer1_outputs(1693) <= not b or a;
    layer1_outputs(1694) <= a or b;
    layer1_outputs(1695) <= b;
    layer1_outputs(1696) <= a or b;
    layer1_outputs(1697) <= b and not a;
    layer1_outputs(1698) <= not (a or b);
    layer1_outputs(1699) <= a;
    layer1_outputs(1700) <= a and not b;
    layer1_outputs(1701) <= a and b;
    layer1_outputs(1702) <= 1'b0;
    layer1_outputs(1703) <= b;
    layer1_outputs(1704) <= a and not b;
    layer1_outputs(1705) <= 1'b1;
    layer1_outputs(1706) <= b and not a;
    layer1_outputs(1707) <= not b;
    layer1_outputs(1708) <= b and not a;
    layer1_outputs(1709) <= a or b;
    layer1_outputs(1710) <= not (a or b);
    layer1_outputs(1711) <= not a;
    layer1_outputs(1712) <= not (a or b);
    layer1_outputs(1713) <= a and b;
    layer1_outputs(1714) <= a and b;
    layer1_outputs(1715) <= not b or a;
    layer1_outputs(1716) <= 1'b0;
    layer1_outputs(1717) <= a;
    layer1_outputs(1718) <= a xor b;
    layer1_outputs(1719) <= not (a or b);
    layer1_outputs(1720) <= not (a and b);
    layer1_outputs(1721) <= b and not a;
    layer1_outputs(1722) <= 1'b1;
    layer1_outputs(1723) <= not (a or b);
    layer1_outputs(1724) <= not b;
    layer1_outputs(1725) <= b;
    layer1_outputs(1726) <= b and not a;
    layer1_outputs(1727) <= b and not a;
    layer1_outputs(1728) <= not a or b;
    layer1_outputs(1729) <= a;
    layer1_outputs(1730) <= not a or b;
    layer1_outputs(1731) <= not a;
    layer1_outputs(1732) <= not b or a;
    layer1_outputs(1733) <= b;
    layer1_outputs(1734) <= a and b;
    layer1_outputs(1735) <= not a;
    layer1_outputs(1736) <= not b or a;
    layer1_outputs(1737) <= not a or b;
    layer1_outputs(1738) <= a and not b;
    layer1_outputs(1739) <= a and not b;
    layer1_outputs(1740) <= not (a and b);
    layer1_outputs(1741) <= not (a and b);
    layer1_outputs(1742) <= a or b;
    layer1_outputs(1743) <= not a or b;
    layer1_outputs(1744) <= a and not b;
    layer1_outputs(1745) <= not (a xor b);
    layer1_outputs(1746) <= not a;
    layer1_outputs(1747) <= a;
    layer1_outputs(1748) <= b;
    layer1_outputs(1749) <= a or b;
    layer1_outputs(1750) <= b;
    layer1_outputs(1751) <= b and not a;
    layer1_outputs(1752) <= not a;
    layer1_outputs(1753) <= not a or b;
    layer1_outputs(1754) <= not (a or b);
    layer1_outputs(1755) <= b and not a;
    layer1_outputs(1756) <= not (a and b);
    layer1_outputs(1757) <= not a or b;
    layer1_outputs(1758) <= not b;
    layer1_outputs(1759) <= a and b;
    layer1_outputs(1760) <= b and not a;
    layer1_outputs(1761) <= a and not b;
    layer1_outputs(1762) <= not b or a;
    layer1_outputs(1763) <= a xor b;
    layer1_outputs(1764) <= b and not a;
    layer1_outputs(1765) <= not a or b;
    layer1_outputs(1766) <= a and not b;
    layer1_outputs(1767) <= not a or b;
    layer1_outputs(1768) <= b;
    layer1_outputs(1769) <= a;
    layer1_outputs(1770) <= a and not b;
    layer1_outputs(1771) <= not a;
    layer1_outputs(1772) <= not b;
    layer1_outputs(1773) <= b;
    layer1_outputs(1774) <= b and not a;
    layer1_outputs(1775) <= a;
    layer1_outputs(1776) <= a;
    layer1_outputs(1777) <= 1'b1;
    layer1_outputs(1778) <= not a;
    layer1_outputs(1779) <= a and not b;
    layer1_outputs(1780) <= a;
    layer1_outputs(1781) <= not b;
    layer1_outputs(1782) <= not a or b;
    layer1_outputs(1783) <= a;
    layer1_outputs(1784) <= b and not a;
    layer1_outputs(1785) <= not (a or b);
    layer1_outputs(1786) <= b;
    layer1_outputs(1787) <= b and not a;
    layer1_outputs(1788) <= not b;
    layer1_outputs(1789) <= not b or a;
    layer1_outputs(1790) <= 1'b0;
    layer1_outputs(1791) <= 1'b1;
    layer1_outputs(1792) <= not (a xor b);
    layer1_outputs(1793) <= not a;
    layer1_outputs(1794) <= not b;
    layer1_outputs(1795) <= not (a and b);
    layer1_outputs(1796) <= not b;
    layer1_outputs(1797) <= 1'b0;
    layer1_outputs(1798) <= not b or a;
    layer1_outputs(1799) <= a and not b;
    layer1_outputs(1800) <= not b or a;
    layer1_outputs(1801) <= a or b;
    layer1_outputs(1802) <= not a or b;
    layer1_outputs(1803) <= a or b;
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= 1'b0;
    layer1_outputs(1806) <= not a;
    layer1_outputs(1807) <= a and not b;
    layer1_outputs(1808) <= 1'b0;
    layer1_outputs(1809) <= 1'b1;
    layer1_outputs(1810) <= not a;
    layer1_outputs(1811) <= not a;
    layer1_outputs(1812) <= a xor b;
    layer1_outputs(1813) <= a and b;
    layer1_outputs(1814) <= not (a or b);
    layer1_outputs(1815) <= not a;
    layer1_outputs(1816) <= a;
    layer1_outputs(1817) <= not (a xor b);
    layer1_outputs(1818) <= not a;
    layer1_outputs(1819) <= not (a xor b);
    layer1_outputs(1820) <= b and not a;
    layer1_outputs(1821) <= b;
    layer1_outputs(1822) <= not a;
    layer1_outputs(1823) <= not (a or b);
    layer1_outputs(1824) <= not a;
    layer1_outputs(1825) <= b;
    layer1_outputs(1826) <= a and not b;
    layer1_outputs(1827) <= a;
    layer1_outputs(1828) <= a;
    layer1_outputs(1829) <= not b or a;
    layer1_outputs(1830) <= not (a or b);
    layer1_outputs(1831) <= not a;
    layer1_outputs(1832) <= not (a or b);
    layer1_outputs(1833) <= not a or b;
    layer1_outputs(1834) <= not b;
    layer1_outputs(1835) <= not (a and b);
    layer1_outputs(1836) <= not b;
    layer1_outputs(1837) <= not a or b;
    layer1_outputs(1838) <= not b or a;
    layer1_outputs(1839) <= not (a and b);
    layer1_outputs(1840) <= not b;
    layer1_outputs(1841) <= not b;
    layer1_outputs(1842) <= a xor b;
    layer1_outputs(1843) <= not (a and b);
    layer1_outputs(1844) <= b and not a;
    layer1_outputs(1845) <= not a or b;
    layer1_outputs(1846) <= not (a or b);
    layer1_outputs(1847) <= not a or b;
    layer1_outputs(1848) <= not b or a;
    layer1_outputs(1849) <= not b;
    layer1_outputs(1850) <= b and not a;
    layer1_outputs(1851) <= not (a or b);
    layer1_outputs(1852) <= not (a and b);
    layer1_outputs(1853) <= not a or b;
    layer1_outputs(1854) <= a and b;
    layer1_outputs(1855) <= b;
    layer1_outputs(1856) <= not a;
    layer1_outputs(1857) <= 1'b1;
    layer1_outputs(1858) <= a and not b;
    layer1_outputs(1859) <= not b or a;
    layer1_outputs(1860) <= a and not b;
    layer1_outputs(1861) <= not a;
    layer1_outputs(1862) <= not b;
    layer1_outputs(1863) <= b;
    layer1_outputs(1864) <= b and not a;
    layer1_outputs(1865) <= not b;
    layer1_outputs(1866) <= b and not a;
    layer1_outputs(1867) <= not b or a;
    layer1_outputs(1868) <= a and not b;
    layer1_outputs(1869) <= not (a and b);
    layer1_outputs(1870) <= b;
    layer1_outputs(1871) <= a or b;
    layer1_outputs(1872) <= a;
    layer1_outputs(1873) <= not b;
    layer1_outputs(1874) <= 1'b0;
    layer1_outputs(1875) <= 1'b0;
    layer1_outputs(1876) <= b;
    layer1_outputs(1877) <= 1'b1;
    layer1_outputs(1878) <= a;
    layer1_outputs(1879) <= a or b;
    layer1_outputs(1880) <= a;
    layer1_outputs(1881) <= not a;
    layer1_outputs(1882) <= 1'b1;
    layer1_outputs(1883) <= not a;
    layer1_outputs(1884) <= not b;
    layer1_outputs(1885) <= not b;
    layer1_outputs(1886) <= b and not a;
    layer1_outputs(1887) <= a;
    layer1_outputs(1888) <= not (a and b);
    layer1_outputs(1889) <= not (a xor b);
    layer1_outputs(1890) <= not (a or b);
    layer1_outputs(1891) <= not a;
    layer1_outputs(1892) <= not (a and b);
    layer1_outputs(1893) <= b;
    layer1_outputs(1894) <= b;
    layer1_outputs(1895) <= a;
    layer1_outputs(1896) <= a xor b;
    layer1_outputs(1897) <= b and not a;
    layer1_outputs(1898) <= a and b;
    layer1_outputs(1899) <= not (a or b);
    layer1_outputs(1900) <= a;
    layer1_outputs(1901) <= b;
    layer1_outputs(1902) <= 1'b0;
    layer1_outputs(1903) <= not (a and b);
    layer1_outputs(1904) <= not (a and b);
    layer1_outputs(1905) <= not (a or b);
    layer1_outputs(1906) <= b;
    layer1_outputs(1907) <= 1'b1;
    layer1_outputs(1908) <= a;
    layer1_outputs(1909) <= not (a and b);
    layer1_outputs(1910) <= b;
    layer1_outputs(1911) <= a xor b;
    layer1_outputs(1912) <= a xor b;
    layer1_outputs(1913) <= not b;
    layer1_outputs(1914) <= b;
    layer1_outputs(1915) <= not b or a;
    layer1_outputs(1916) <= not b;
    layer1_outputs(1917) <= a and b;
    layer1_outputs(1918) <= not a;
    layer1_outputs(1919) <= a or b;
    layer1_outputs(1920) <= not (a and b);
    layer1_outputs(1921) <= not (a and b);
    layer1_outputs(1922) <= not b;
    layer1_outputs(1923) <= a;
    layer1_outputs(1924) <= a or b;
    layer1_outputs(1925) <= b and not a;
    layer1_outputs(1926) <= not (a xor b);
    layer1_outputs(1927) <= a or b;
    layer1_outputs(1928) <= not (a xor b);
    layer1_outputs(1929) <= a xor b;
    layer1_outputs(1930) <= not (a and b);
    layer1_outputs(1931) <= not a or b;
    layer1_outputs(1932) <= not b or a;
    layer1_outputs(1933) <= not (a or b);
    layer1_outputs(1934) <= not a;
    layer1_outputs(1935) <= not b;
    layer1_outputs(1936) <= a or b;
    layer1_outputs(1937) <= a and b;
    layer1_outputs(1938) <= a;
    layer1_outputs(1939) <= a or b;
    layer1_outputs(1940) <= not (a or b);
    layer1_outputs(1941) <= a and b;
    layer1_outputs(1942) <= a or b;
    layer1_outputs(1943) <= a and b;
    layer1_outputs(1944) <= not b;
    layer1_outputs(1945) <= a or b;
    layer1_outputs(1946) <= not a or b;
    layer1_outputs(1947) <= not a or b;
    layer1_outputs(1948) <= 1'b1;
    layer1_outputs(1949) <= a;
    layer1_outputs(1950) <= not a or b;
    layer1_outputs(1951) <= a;
    layer1_outputs(1952) <= not a;
    layer1_outputs(1953) <= 1'b0;
    layer1_outputs(1954) <= not a or b;
    layer1_outputs(1955) <= 1'b0;
    layer1_outputs(1956) <= not a or b;
    layer1_outputs(1957) <= not (a or b);
    layer1_outputs(1958) <= a xor b;
    layer1_outputs(1959) <= a and not b;
    layer1_outputs(1960) <= a or b;
    layer1_outputs(1961) <= not (a or b);
    layer1_outputs(1962) <= b and not a;
    layer1_outputs(1963) <= a xor b;
    layer1_outputs(1964) <= not b;
    layer1_outputs(1965) <= 1'b0;
    layer1_outputs(1966) <= 1'b0;
    layer1_outputs(1967) <= not b or a;
    layer1_outputs(1968) <= a or b;
    layer1_outputs(1969) <= a and b;
    layer1_outputs(1970) <= not a or b;
    layer1_outputs(1971) <= a or b;
    layer1_outputs(1972) <= not (a and b);
    layer1_outputs(1973) <= a or b;
    layer1_outputs(1974) <= b;
    layer1_outputs(1975) <= not (a and b);
    layer1_outputs(1976) <= a and b;
    layer1_outputs(1977) <= b and not a;
    layer1_outputs(1978) <= not b;
    layer1_outputs(1979) <= a or b;
    layer1_outputs(1980) <= not (a and b);
    layer1_outputs(1981) <= 1'b1;
    layer1_outputs(1982) <= not b or a;
    layer1_outputs(1983) <= not a or b;
    layer1_outputs(1984) <= a or b;
    layer1_outputs(1985) <= b and not a;
    layer1_outputs(1986) <= 1'b1;
    layer1_outputs(1987) <= not a or b;
    layer1_outputs(1988) <= not b or a;
    layer1_outputs(1989) <= not (a xor b);
    layer1_outputs(1990) <= a and not b;
    layer1_outputs(1991) <= not a or b;
    layer1_outputs(1992) <= b and not a;
    layer1_outputs(1993) <= a and not b;
    layer1_outputs(1994) <= b and not a;
    layer1_outputs(1995) <= b;
    layer1_outputs(1996) <= b and not a;
    layer1_outputs(1997) <= not a or b;
    layer1_outputs(1998) <= not b or a;
    layer1_outputs(1999) <= 1'b0;
    layer1_outputs(2000) <= a or b;
    layer1_outputs(2001) <= not a;
    layer1_outputs(2002) <= a or b;
    layer1_outputs(2003) <= not (a or b);
    layer1_outputs(2004) <= not a or b;
    layer1_outputs(2005) <= not b;
    layer1_outputs(2006) <= b;
    layer1_outputs(2007) <= not b or a;
    layer1_outputs(2008) <= a xor b;
    layer1_outputs(2009) <= not b or a;
    layer1_outputs(2010) <= not b;
    layer1_outputs(2011) <= b;
    layer1_outputs(2012) <= not b or a;
    layer1_outputs(2013) <= a xor b;
    layer1_outputs(2014) <= 1'b0;
    layer1_outputs(2015) <= not (a and b);
    layer1_outputs(2016) <= not a;
    layer1_outputs(2017) <= b and not a;
    layer1_outputs(2018) <= not (a and b);
    layer1_outputs(2019) <= a;
    layer1_outputs(2020) <= b;
    layer1_outputs(2021) <= 1'b0;
    layer1_outputs(2022) <= 1'b1;
    layer1_outputs(2023) <= not b or a;
    layer1_outputs(2024) <= a and not b;
    layer1_outputs(2025) <= not (a and b);
    layer1_outputs(2026) <= a;
    layer1_outputs(2027) <= not a;
    layer1_outputs(2028) <= not a or b;
    layer1_outputs(2029) <= 1'b0;
    layer1_outputs(2030) <= not b;
    layer1_outputs(2031) <= b;
    layer1_outputs(2032) <= not b;
    layer1_outputs(2033) <= not b or a;
    layer1_outputs(2034) <= not a or b;
    layer1_outputs(2035) <= not b;
    layer1_outputs(2036) <= not b or a;
    layer1_outputs(2037) <= not b or a;
    layer1_outputs(2038) <= a and not b;
    layer1_outputs(2039) <= b;
    layer1_outputs(2040) <= a xor b;
    layer1_outputs(2041) <= not b or a;
    layer1_outputs(2042) <= not b;
    layer1_outputs(2043) <= not a or b;
    layer1_outputs(2044) <= a and b;
    layer1_outputs(2045) <= a and b;
    layer1_outputs(2046) <= not (a xor b);
    layer1_outputs(2047) <= 1'b0;
    layer1_outputs(2048) <= not (a or b);
    layer1_outputs(2049) <= b;
    layer1_outputs(2050) <= not (a and b);
    layer1_outputs(2051) <= not a or b;
    layer1_outputs(2052) <= 1'b1;
    layer1_outputs(2053) <= not a;
    layer1_outputs(2054) <= a or b;
    layer1_outputs(2055) <= 1'b1;
    layer1_outputs(2056) <= a and b;
    layer1_outputs(2057) <= not b;
    layer1_outputs(2058) <= not (a or b);
    layer1_outputs(2059) <= not b;
    layer1_outputs(2060) <= b;
    layer1_outputs(2061) <= not a;
    layer1_outputs(2062) <= a or b;
    layer1_outputs(2063) <= not (a and b);
    layer1_outputs(2064) <= not a;
    layer1_outputs(2065) <= not b or a;
    layer1_outputs(2066) <= a and b;
    layer1_outputs(2067) <= a xor b;
    layer1_outputs(2068) <= a;
    layer1_outputs(2069) <= not a or b;
    layer1_outputs(2070) <= not a;
    layer1_outputs(2071) <= 1'b1;
    layer1_outputs(2072) <= a and not b;
    layer1_outputs(2073) <= not b or a;
    layer1_outputs(2074) <= a or b;
    layer1_outputs(2075) <= b;
    layer1_outputs(2076) <= not a or b;
    layer1_outputs(2077) <= b;
    layer1_outputs(2078) <= not (a and b);
    layer1_outputs(2079) <= 1'b1;
    layer1_outputs(2080) <= not a;
    layer1_outputs(2081) <= a or b;
    layer1_outputs(2082) <= a and not b;
    layer1_outputs(2083) <= not (a and b);
    layer1_outputs(2084) <= a and b;
    layer1_outputs(2085) <= a xor b;
    layer1_outputs(2086) <= not a;
    layer1_outputs(2087) <= 1'b0;
    layer1_outputs(2088) <= 1'b1;
    layer1_outputs(2089) <= not a or b;
    layer1_outputs(2090) <= not b;
    layer1_outputs(2091) <= a xor b;
    layer1_outputs(2092) <= not b or a;
    layer1_outputs(2093) <= b;
    layer1_outputs(2094) <= a;
    layer1_outputs(2095) <= 1'b0;
    layer1_outputs(2096) <= not (a or b);
    layer1_outputs(2097) <= a;
    layer1_outputs(2098) <= not a;
    layer1_outputs(2099) <= not b;
    layer1_outputs(2100) <= not (a or b);
    layer1_outputs(2101) <= not (a or b);
    layer1_outputs(2102) <= a and b;
    layer1_outputs(2103) <= not a;
    layer1_outputs(2104) <= b and not a;
    layer1_outputs(2105) <= a and b;
    layer1_outputs(2106) <= b and not a;
    layer1_outputs(2107) <= a;
    layer1_outputs(2108) <= a and b;
    layer1_outputs(2109) <= not a or b;
    layer1_outputs(2110) <= a and not b;
    layer1_outputs(2111) <= not a;
    layer1_outputs(2112) <= a and b;
    layer1_outputs(2113) <= a and b;
    layer1_outputs(2114) <= not (a xor b);
    layer1_outputs(2115) <= not a or b;
    layer1_outputs(2116) <= a and not b;
    layer1_outputs(2117) <= b;
    layer1_outputs(2118) <= 1'b1;
    layer1_outputs(2119) <= not (a and b);
    layer1_outputs(2120) <= not (a and b);
    layer1_outputs(2121) <= a and b;
    layer1_outputs(2122) <= b and not a;
    layer1_outputs(2123) <= not a or b;
    layer1_outputs(2124) <= a and b;
    layer1_outputs(2125) <= not a or b;
    layer1_outputs(2126) <= b;
    layer1_outputs(2127) <= a or b;
    layer1_outputs(2128) <= not b or a;
    layer1_outputs(2129) <= b;
    layer1_outputs(2130) <= not a or b;
    layer1_outputs(2131) <= a or b;
    layer1_outputs(2132) <= not (a and b);
    layer1_outputs(2133) <= not (a or b);
    layer1_outputs(2134) <= not (a or b);
    layer1_outputs(2135) <= 1'b1;
    layer1_outputs(2136) <= a;
    layer1_outputs(2137) <= 1'b0;
    layer1_outputs(2138) <= a;
    layer1_outputs(2139) <= not b or a;
    layer1_outputs(2140) <= b and not a;
    layer1_outputs(2141) <= not (a and b);
    layer1_outputs(2142) <= a or b;
    layer1_outputs(2143) <= not a or b;
    layer1_outputs(2144) <= a and not b;
    layer1_outputs(2145) <= b;
    layer1_outputs(2146) <= b and not a;
    layer1_outputs(2147) <= a xor b;
    layer1_outputs(2148) <= not (a and b);
    layer1_outputs(2149) <= 1'b1;
    layer1_outputs(2150) <= not a or b;
    layer1_outputs(2151) <= not a or b;
    layer1_outputs(2152) <= a xor b;
    layer1_outputs(2153) <= b;
    layer1_outputs(2154) <= b and not a;
    layer1_outputs(2155) <= a and not b;
    layer1_outputs(2156) <= not (a xor b);
    layer1_outputs(2157) <= b;
    layer1_outputs(2158) <= not a or b;
    layer1_outputs(2159) <= not a or b;
    layer1_outputs(2160) <= not b or a;
    layer1_outputs(2161) <= b;
    layer1_outputs(2162) <= not (a or b);
    layer1_outputs(2163) <= 1'b1;
    layer1_outputs(2164) <= 1'b0;
    layer1_outputs(2165) <= 1'b0;
    layer1_outputs(2166) <= a and not b;
    layer1_outputs(2167) <= not (a xor b);
    layer1_outputs(2168) <= not (a and b);
    layer1_outputs(2169) <= not a;
    layer1_outputs(2170) <= not (a or b);
    layer1_outputs(2171) <= b and not a;
    layer1_outputs(2172) <= not (a or b);
    layer1_outputs(2173) <= b;
    layer1_outputs(2174) <= b;
    layer1_outputs(2175) <= b;
    layer1_outputs(2176) <= not b or a;
    layer1_outputs(2177) <= not a or b;
    layer1_outputs(2178) <= a or b;
    layer1_outputs(2179) <= a and b;
    layer1_outputs(2180) <= not b;
    layer1_outputs(2181) <= a and b;
    layer1_outputs(2182) <= a xor b;
    layer1_outputs(2183) <= 1'b0;
    layer1_outputs(2184) <= b;
    layer1_outputs(2185) <= not b or a;
    layer1_outputs(2186) <= b;
    layer1_outputs(2187) <= not b;
    layer1_outputs(2188) <= a and b;
    layer1_outputs(2189) <= not a;
    layer1_outputs(2190) <= 1'b1;
    layer1_outputs(2191) <= not b or a;
    layer1_outputs(2192) <= not (a or b);
    layer1_outputs(2193) <= not b or a;
    layer1_outputs(2194) <= a;
    layer1_outputs(2195) <= not b;
    layer1_outputs(2196) <= not a or b;
    layer1_outputs(2197) <= a and not b;
    layer1_outputs(2198) <= a;
    layer1_outputs(2199) <= a xor b;
    layer1_outputs(2200) <= a or b;
    layer1_outputs(2201) <= not (a or b);
    layer1_outputs(2202) <= a;
    layer1_outputs(2203) <= b and not a;
    layer1_outputs(2204) <= b and not a;
    layer1_outputs(2205) <= not (a xor b);
    layer1_outputs(2206) <= a;
    layer1_outputs(2207) <= a or b;
    layer1_outputs(2208) <= not a or b;
    layer1_outputs(2209) <= not a or b;
    layer1_outputs(2210) <= not a;
    layer1_outputs(2211) <= not b;
    layer1_outputs(2212) <= not (a and b);
    layer1_outputs(2213) <= a and not b;
    layer1_outputs(2214) <= a;
    layer1_outputs(2215) <= a and b;
    layer1_outputs(2216) <= not b or a;
    layer1_outputs(2217) <= a and b;
    layer1_outputs(2218) <= b and not a;
    layer1_outputs(2219) <= a and not b;
    layer1_outputs(2220) <= a or b;
    layer1_outputs(2221) <= a or b;
    layer1_outputs(2222) <= a;
    layer1_outputs(2223) <= b;
    layer1_outputs(2224) <= 1'b1;
    layer1_outputs(2225) <= 1'b1;
    layer1_outputs(2226) <= a or b;
    layer1_outputs(2227) <= b;
    layer1_outputs(2228) <= not b;
    layer1_outputs(2229) <= not b or a;
    layer1_outputs(2230) <= a and not b;
    layer1_outputs(2231) <= not b;
    layer1_outputs(2232) <= not (a xor b);
    layer1_outputs(2233) <= 1'b0;
    layer1_outputs(2234) <= not (a and b);
    layer1_outputs(2235) <= a or b;
    layer1_outputs(2236) <= a or b;
    layer1_outputs(2237) <= b and not a;
    layer1_outputs(2238) <= a;
    layer1_outputs(2239) <= not a or b;
    layer1_outputs(2240) <= a xor b;
    layer1_outputs(2241) <= a and not b;
    layer1_outputs(2242) <= a xor b;
    layer1_outputs(2243) <= not (a and b);
    layer1_outputs(2244) <= not (a and b);
    layer1_outputs(2245) <= a;
    layer1_outputs(2246) <= a and not b;
    layer1_outputs(2247) <= 1'b1;
    layer1_outputs(2248) <= a and b;
    layer1_outputs(2249) <= not b or a;
    layer1_outputs(2250) <= 1'b0;
    layer1_outputs(2251) <= a or b;
    layer1_outputs(2252) <= not (a xor b);
    layer1_outputs(2253) <= 1'b0;
    layer1_outputs(2254) <= not (a and b);
    layer1_outputs(2255) <= b and not a;
    layer1_outputs(2256) <= b;
    layer1_outputs(2257) <= 1'b0;
    layer1_outputs(2258) <= not b or a;
    layer1_outputs(2259) <= not (a xor b);
    layer1_outputs(2260) <= not b or a;
    layer1_outputs(2261) <= 1'b0;
    layer1_outputs(2262) <= not (a and b);
    layer1_outputs(2263) <= not (a xor b);
    layer1_outputs(2264) <= a and b;
    layer1_outputs(2265) <= not a;
    layer1_outputs(2266) <= a and b;
    layer1_outputs(2267) <= not b;
    layer1_outputs(2268) <= not b or a;
    layer1_outputs(2269) <= b and not a;
    layer1_outputs(2270) <= b and not a;
    layer1_outputs(2271) <= 1'b0;
    layer1_outputs(2272) <= not (a xor b);
    layer1_outputs(2273) <= not a;
    layer1_outputs(2274) <= not b or a;
    layer1_outputs(2275) <= not b;
    layer1_outputs(2276) <= 1'b0;
    layer1_outputs(2277) <= 1'b0;
    layer1_outputs(2278) <= not (a and b);
    layer1_outputs(2279) <= not (a xor b);
    layer1_outputs(2280) <= a or b;
    layer1_outputs(2281) <= not a;
    layer1_outputs(2282) <= not a;
    layer1_outputs(2283) <= a;
    layer1_outputs(2284) <= b and not a;
    layer1_outputs(2285) <= 1'b0;
    layer1_outputs(2286) <= a and b;
    layer1_outputs(2287) <= b;
    layer1_outputs(2288) <= not b;
    layer1_outputs(2289) <= b and not a;
    layer1_outputs(2290) <= b and not a;
    layer1_outputs(2291) <= a or b;
    layer1_outputs(2292) <= b;
    layer1_outputs(2293) <= not (a or b);
    layer1_outputs(2294) <= not a or b;
    layer1_outputs(2295) <= a or b;
    layer1_outputs(2296) <= not (a and b);
    layer1_outputs(2297) <= a or b;
    layer1_outputs(2298) <= not (a or b);
    layer1_outputs(2299) <= b;
    layer1_outputs(2300) <= not a;
    layer1_outputs(2301) <= a and b;
    layer1_outputs(2302) <= not (a and b);
    layer1_outputs(2303) <= 1'b1;
    layer1_outputs(2304) <= a and b;
    layer1_outputs(2305) <= not a;
    layer1_outputs(2306) <= b and not a;
    layer1_outputs(2307) <= not (a or b);
    layer1_outputs(2308) <= not (a or b);
    layer1_outputs(2309) <= not b;
    layer1_outputs(2310) <= not b;
    layer1_outputs(2311) <= not (a or b);
    layer1_outputs(2312) <= not (a xor b);
    layer1_outputs(2313) <= not (a or b);
    layer1_outputs(2314) <= not (a or b);
    layer1_outputs(2315) <= not b or a;
    layer1_outputs(2316) <= not (a or b);
    layer1_outputs(2317) <= not a;
    layer1_outputs(2318) <= not a;
    layer1_outputs(2319) <= not a or b;
    layer1_outputs(2320) <= a or b;
    layer1_outputs(2321) <= not a;
    layer1_outputs(2322) <= not (a and b);
    layer1_outputs(2323) <= a;
    layer1_outputs(2324) <= not a;
    layer1_outputs(2325) <= not (a or b);
    layer1_outputs(2326) <= not b or a;
    layer1_outputs(2327) <= not b;
    layer1_outputs(2328) <= not (a or b);
    layer1_outputs(2329) <= not (a xor b);
    layer1_outputs(2330) <= not b;
    layer1_outputs(2331) <= a or b;
    layer1_outputs(2332) <= not (a or b);
    layer1_outputs(2333) <= not (a or b);
    layer1_outputs(2334) <= a or b;
    layer1_outputs(2335) <= not (a or b);
    layer1_outputs(2336) <= not (a and b);
    layer1_outputs(2337) <= not a;
    layer1_outputs(2338) <= not a;
    layer1_outputs(2339) <= a and not b;
    layer1_outputs(2340) <= a and not b;
    layer1_outputs(2341) <= not (a and b);
    layer1_outputs(2342) <= b and not a;
    layer1_outputs(2343) <= not b;
    layer1_outputs(2344) <= not a or b;
    layer1_outputs(2345) <= a;
    layer1_outputs(2346) <= a or b;
    layer1_outputs(2347) <= not a;
    layer1_outputs(2348) <= 1'b1;
    layer1_outputs(2349) <= not b;
    layer1_outputs(2350) <= not b;
    layer1_outputs(2351) <= not a or b;
    layer1_outputs(2352) <= a;
    layer1_outputs(2353) <= a;
    layer1_outputs(2354) <= not b;
    layer1_outputs(2355) <= a;
    layer1_outputs(2356) <= not (a xor b);
    layer1_outputs(2357) <= not (a or b);
    layer1_outputs(2358) <= not (a or b);
    layer1_outputs(2359) <= b;
    layer1_outputs(2360) <= not b or a;
    layer1_outputs(2361) <= not a or b;
    layer1_outputs(2362) <= not b;
    layer1_outputs(2363) <= a and b;
    layer1_outputs(2364) <= not a;
    layer1_outputs(2365) <= a or b;
    layer1_outputs(2366) <= 1'b0;
    layer1_outputs(2367) <= not b;
    layer1_outputs(2368) <= a;
    layer1_outputs(2369) <= b;
    layer1_outputs(2370) <= not a or b;
    layer1_outputs(2371) <= a;
    layer1_outputs(2372) <= not a;
    layer1_outputs(2373) <= not a;
    layer1_outputs(2374) <= a;
    layer1_outputs(2375) <= a or b;
    layer1_outputs(2376) <= a;
    layer1_outputs(2377) <= 1'b1;
    layer1_outputs(2378) <= b;
    layer1_outputs(2379) <= not a;
    layer1_outputs(2380) <= not a or b;
    layer1_outputs(2381) <= 1'b0;
    layer1_outputs(2382) <= not a;
    layer1_outputs(2383) <= a and b;
    layer1_outputs(2384) <= not a or b;
    layer1_outputs(2385) <= not a or b;
    layer1_outputs(2386) <= 1'b0;
    layer1_outputs(2387) <= not a;
    layer1_outputs(2388) <= not a;
    layer1_outputs(2389) <= a and not b;
    layer1_outputs(2390) <= 1'b0;
    layer1_outputs(2391) <= not a;
    layer1_outputs(2392) <= a xor b;
    layer1_outputs(2393) <= a;
    layer1_outputs(2394) <= a;
    layer1_outputs(2395) <= not b or a;
    layer1_outputs(2396) <= not a;
    layer1_outputs(2397) <= not b;
    layer1_outputs(2398) <= a and b;
    layer1_outputs(2399) <= not a;
    layer1_outputs(2400) <= a;
    layer1_outputs(2401) <= a and b;
    layer1_outputs(2402) <= not b or a;
    layer1_outputs(2403) <= not b;
    layer1_outputs(2404) <= not b or a;
    layer1_outputs(2405) <= not b or a;
    layer1_outputs(2406) <= 1'b1;
    layer1_outputs(2407) <= b;
    layer1_outputs(2408) <= a and not b;
    layer1_outputs(2409) <= 1'b0;
    layer1_outputs(2410) <= not b or a;
    layer1_outputs(2411) <= 1'b1;
    layer1_outputs(2412) <= b and not a;
    layer1_outputs(2413) <= a;
    layer1_outputs(2414) <= not (a or b);
    layer1_outputs(2415) <= a;
    layer1_outputs(2416) <= not (a or b);
    layer1_outputs(2417) <= a and not b;
    layer1_outputs(2418) <= a and not b;
    layer1_outputs(2419) <= b;
    layer1_outputs(2420) <= a;
    layer1_outputs(2421) <= b;
    layer1_outputs(2422) <= a and not b;
    layer1_outputs(2423) <= not (a and b);
    layer1_outputs(2424) <= 1'b0;
    layer1_outputs(2425) <= a or b;
    layer1_outputs(2426) <= not a;
    layer1_outputs(2427) <= b;
    layer1_outputs(2428) <= b and not a;
    layer1_outputs(2429) <= not (a xor b);
    layer1_outputs(2430) <= not (a and b);
    layer1_outputs(2431) <= not a;
    layer1_outputs(2432) <= not b or a;
    layer1_outputs(2433) <= not (a or b);
    layer1_outputs(2434) <= not (a or b);
    layer1_outputs(2435) <= b and not a;
    layer1_outputs(2436) <= a or b;
    layer1_outputs(2437) <= not (a and b);
    layer1_outputs(2438) <= not (a and b);
    layer1_outputs(2439) <= 1'b1;
    layer1_outputs(2440) <= b;
    layer1_outputs(2441) <= a and b;
    layer1_outputs(2442) <= a and b;
    layer1_outputs(2443) <= not a;
    layer1_outputs(2444) <= 1'b0;
    layer1_outputs(2445) <= not (a or b);
    layer1_outputs(2446) <= a;
    layer1_outputs(2447) <= b;
    layer1_outputs(2448) <= not b;
    layer1_outputs(2449) <= a and not b;
    layer1_outputs(2450) <= not b or a;
    layer1_outputs(2451) <= not b or a;
    layer1_outputs(2452) <= not (a or b);
    layer1_outputs(2453) <= b and not a;
    layer1_outputs(2454) <= not (a or b);
    layer1_outputs(2455) <= not b;
    layer1_outputs(2456) <= not (a and b);
    layer1_outputs(2457) <= not b;
    layer1_outputs(2458) <= not b;
    layer1_outputs(2459) <= a;
    layer1_outputs(2460) <= b;
    layer1_outputs(2461) <= not a;
    layer1_outputs(2462) <= not (a xor b);
    layer1_outputs(2463) <= not b;
    layer1_outputs(2464) <= not (a or b);
    layer1_outputs(2465) <= not a;
    layer1_outputs(2466) <= a and not b;
    layer1_outputs(2467) <= not a or b;
    layer1_outputs(2468) <= a xor b;
    layer1_outputs(2469) <= 1'b1;
    layer1_outputs(2470) <= not b;
    layer1_outputs(2471) <= a xor b;
    layer1_outputs(2472) <= b and not a;
    layer1_outputs(2473) <= not (a or b);
    layer1_outputs(2474) <= not b;
    layer1_outputs(2475) <= a;
    layer1_outputs(2476) <= a;
    layer1_outputs(2477) <= a;
    layer1_outputs(2478) <= a or b;
    layer1_outputs(2479) <= not a;
    layer1_outputs(2480) <= not b;
    layer1_outputs(2481) <= not (a xor b);
    layer1_outputs(2482) <= not a;
    layer1_outputs(2483) <= not b;
    layer1_outputs(2484) <= not b or a;
    layer1_outputs(2485) <= a and b;
    layer1_outputs(2486) <= a and b;
    layer1_outputs(2487) <= b;
    layer1_outputs(2488) <= not a or b;
    layer1_outputs(2489) <= not (a and b);
    layer1_outputs(2490) <= a;
    layer1_outputs(2491) <= a;
    layer1_outputs(2492) <= b and not a;
    layer1_outputs(2493) <= a or b;
    layer1_outputs(2494) <= 1'b1;
    layer1_outputs(2495) <= a and not b;
    layer1_outputs(2496) <= b and not a;
    layer1_outputs(2497) <= not (a and b);
    layer1_outputs(2498) <= a and not b;
    layer1_outputs(2499) <= 1'b1;
    layer1_outputs(2500) <= not a;
    layer1_outputs(2501) <= not a or b;
    layer1_outputs(2502) <= not b;
    layer1_outputs(2503) <= not b or a;
    layer1_outputs(2504) <= not a;
    layer1_outputs(2505) <= not b;
    layer1_outputs(2506) <= not b or a;
    layer1_outputs(2507) <= not (a and b);
    layer1_outputs(2508) <= a xor b;
    layer1_outputs(2509) <= not a;
    layer1_outputs(2510) <= not (a and b);
    layer1_outputs(2511) <= not a or b;
    layer1_outputs(2512) <= b;
    layer1_outputs(2513) <= b;
    layer1_outputs(2514) <= a and b;
    layer1_outputs(2515) <= a and not b;
    layer1_outputs(2516) <= not (a or b);
    layer1_outputs(2517) <= not (a or b);
    layer1_outputs(2518) <= b and not a;
    layer1_outputs(2519) <= a and not b;
    layer1_outputs(2520) <= not b;
    layer1_outputs(2521) <= b;
    layer1_outputs(2522) <= a and not b;
    layer1_outputs(2523) <= a or b;
    layer1_outputs(2524) <= not b;
    layer1_outputs(2525) <= b and not a;
    layer1_outputs(2526) <= 1'b1;
    layer1_outputs(2527) <= a and b;
    layer1_outputs(2528) <= not a or b;
    layer1_outputs(2529) <= not a or b;
    layer1_outputs(2530) <= not (a xor b);
    layer1_outputs(2531) <= not a;
    layer1_outputs(2532) <= not (a xor b);
    layer1_outputs(2533) <= not (a or b);
    layer1_outputs(2534) <= not a;
    layer1_outputs(2535) <= a and not b;
    layer1_outputs(2536) <= not b or a;
    layer1_outputs(2537) <= a;
    layer1_outputs(2538) <= not a or b;
    layer1_outputs(2539) <= a or b;
    layer1_outputs(2540) <= not a or b;
    layer1_outputs(2541) <= b;
    layer1_outputs(2542) <= a and b;
    layer1_outputs(2543) <= not (a xor b);
    layer1_outputs(2544) <= not (a and b);
    layer1_outputs(2545) <= not b;
    layer1_outputs(2546) <= a;
    layer1_outputs(2547) <= not (a and b);
    layer1_outputs(2548) <= not b or a;
    layer1_outputs(2549) <= not b or a;
    layer1_outputs(2550) <= a and b;
    layer1_outputs(2551) <= a;
    layer1_outputs(2552) <= not a or b;
    layer1_outputs(2553) <= 1'b1;
    layer1_outputs(2554) <= 1'b1;
    layer1_outputs(2555) <= a;
    layer1_outputs(2556) <= a;
    layer1_outputs(2557) <= not a;
    layer1_outputs(2558) <= a and b;
    layer1_outputs(2559) <= a and b;
    layer2_outputs(0) <= 1'b0;
    layer2_outputs(1) <= b;
    layer2_outputs(2) <= not a or b;
    layer2_outputs(3) <= not b or a;
    layer2_outputs(4) <= not b;
    layer2_outputs(5) <= not a or b;
    layer2_outputs(6) <= a;
    layer2_outputs(7) <= not a;
    layer2_outputs(8) <= b;
    layer2_outputs(9) <= not b;
    layer2_outputs(10) <= not (a xor b);
    layer2_outputs(11) <= not (a or b);
    layer2_outputs(12) <= not a or b;
    layer2_outputs(13) <= not a;
    layer2_outputs(14) <= 1'b1;
    layer2_outputs(15) <= not a or b;
    layer2_outputs(16) <= 1'b1;
    layer2_outputs(17) <= not b;
    layer2_outputs(18) <= a and not b;
    layer2_outputs(19) <= b;
    layer2_outputs(20) <= not b;
    layer2_outputs(21) <= b and not a;
    layer2_outputs(22) <= not (a and b);
    layer2_outputs(23) <= not a;
    layer2_outputs(24) <= not b;
    layer2_outputs(25) <= not (a and b);
    layer2_outputs(26) <= 1'b0;
    layer2_outputs(27) <= a or b;
    layer2_outputs(28) <= not (a or b);
    layer2_outputs(29) <= a or b;
    layer2_outputs(30) <= not (a or b);
    layer2_outputs(31) <= b and not a;
    layer2_outputs(32) <= a and not b;
    layer2_outputs(33) <= not b;
    layer2_outputs(34) <= b;
    layer2_outputs(35) <= not b;
    layer2_outputs(36) <= not b or a;
    layer2_outputs(37) <= 1'b1;
    layer2_outputs(38) <= not b or a;
    layer2_outputs(39) <= b;
    layer2_outputs(40) <= 1'b0;
    layer2_outputs(41) <= not a or b;
    layer2_outputs(42) <= not a;
    layer2_outputs(43) <= b;
    layer2_outputs(44) <= not b or a;
    layer2_outputs(45) <= not a;
    layer2_outputs(46) <= b and not a;
    layer2_outputs(47) <= not b;
    layer2_outputs(48) <= not a;
    layer2_outputs(49) <= a or b;
    layer2_outputs(50) <= a;
    layer2_outputs(51) <= b;
    layer2_outputs(52) <= a;
    layer2_outputs(53) <= b and not a;
    layer2_outputs(54) <= a and not b;
    layer2_outputs(55) <= not b;
    layer2_outputs(56) <= b;
    layer2_outputs(57) <= not b or a;
    layer2_outputs(58) <= b;
    layer2_outputs(59) <= not (a or b);
    layer2_outputs(60) <= b and not a;
    layer2_outputs(61) <= not (a and b);
    layer2_outputs(62) <= a and b;
    layer2_outputs(63) <= not b;
    layer2_outputs(64) <= not (a and b);
    layer2_outputs(65) <= b and not a;
    layer2_outputs(66) <= b and not a;
    layer2_outputs(67) <= 1'b1;
    layer2_outputs(68) <= 1'b0;
    layer2_outputs(69) <= not b;
    layer2_outputs(70) <= b and not a;
    layer2_outputs(71) <= 1'b1;
    layer2_outputs(72) <= not a or b;
    layer2_outputs(73) <= a and b;
    layer2_outputs(74) <= not a;
    layer2_outputs(75) <= a xor b;
    layer2_outputs(76) <= a;
    layer2_outputs(77) <= a and not b;
    layer2_outputs(78) <= a xor b;
    layer2_outputs(79) <= not b or a;
    layer2_outputs(80) <= a;
    layer2_outputs(81) <= b and not a;
    layer2_outputs(82) <= a and b;
    layer2_outputs(83) <= a;
    layer2_outputs(84) <= b;
    layer2_outputs(85) <= a and b;
    layer2_outputs(86) <= b and not a;
    layer2_outputs(87) <= not b;
    layer2_outputs(88) <= a and b;
    layer2_outputs(89) <= b;
    layer2_outputs(90) <= not a or b;
    layer2_outputs(91) <= not a;
    layer2_outputs(92) <= b and not a;
    layer2_outputs(93) <= a or b;
    layer2_outputs(94) <= 1'b0;
    layer2_outputs(95) <= a and b;
    layer2_outputs(96) <= not a or b;
    layer2_outputs(97) <= not a or b;
    layer2_outputs(98) <= not (a and b);
    layer2_outputs(99) <= not (a xor b);
    layer2_outputs(100) <= not (a xor b);
    layer2_outputs(101) <= b;
    layer2_outputs(102) <= b;
    layer2_outputs(103) <= a;
    layer2_outputs(104) <= a and not b;
    layer2_outputs(105) <= not a;
    layer2_outputs(106) <= a or b;
    layer2_outputs(107) <= not (a and b);
    layer2_outputs(108) <= not (a or b);
    layer2_outputs(109) <= a and not b;
    layer2_outputs(110) <= not b;
    layer2_outputs(111) <= a xor b;
    layer2_outputs(112) <= 1'b1;
    layer2_outputs(113) <= a;
    layer2_outputs(114) <= b and not a;
    layer2_outputs(115) <= b and not a;
    layer2_outputs(116) <= b and not a;
    layer2_outputs(117) <= a or b;
    layer2_outputs(118) <= not (a xor b);
    layer2_outputs(119) <= a and b;
    layer2_outputs(120) <= a and not b;
    layer2_outputs(121) <= not a;
    layer2_outputs(122) <= not (a and b);
    layer2_outputs(123) <= a and b;
    layer2_outputs(124) <= 1'b0;
    layer2_outputs(125) <= b;
    layer2_outputs(126) <= not b or a;
    layer2_outputs(127) <= a and not b;
    layer2_outputs(128) <= b;
    layer2_outputs(129) <= not (a or b);
    layer2_outputs(130) <= 1'b0;
    layer2_outputs(131) <= not (a and b);
    layer2_outputs(132) <= not a;
    layer2_outputs(133) <= not (a or b);
    layer2_outputs(134) <= 1'b1;
    layer2_outputs(135) <= not (a and b);
    layer2_outputs(136) <= 1'b1;
    layer2_outputs(137) <= not a or b;
    layer2_outputs(138) <= a and not b;
    layer2_outputs(139) <= not (a and b);
    layer2_outputs(140) <= not a;
    layer2_outputs(141) <= not a;
    layer2_outputs(142) <= a;
    layer2_outputs(143) <= a and not b;
    layer2_outputs(144) <= not a;
    layer2_outputs(145) <= a and not b;
    layer2_outputs(146) <= a or b;
    layer2_outputs(147) <= a and b;
    layer2_outputs(148) <= a or b;
    layer2_outputs(149) <= b;
    layer2_outputs(150) <= a;
    layer2_outputs(151) <= a xor b;
    layer2_outputs(152) <= a and b;
    layer2_outputs(153) <= not (a or b);
    layer2_outputs(154) <= a;
    layer2_outputs(155) <= not b;
    layer2_outputs(156) <= not (a or b);
    layer2_outputs(157) <= b;
    layer2_outputs(158) <= a or b;
    layer2_outputs(159) <= not (a or b);
    layer2_outputs(160) <= not b or a;
    layer2_outputs(161) <= not b;
    layer2_outputs(162) <= not (a or b);
    layer2_outputs(163) <= b;
    layer2_outputs(164) <= b;
    layer2_outputs(165) <= not a or b;
    layer2_outputs(166) <= b and not a;
    layer2_outputs(167) <= b and not a;
    layer2_outputs(168) <= a;
    layer2_outputs(169) <= not b or a;
    layer2_outputs(170) <= 1'b1;
    layer2_outputs(171) <= not a or b;
    layer2_outputs(172) <= a xor b;
    layer2_outputs(173) <= b;
    layer2_outputs(174) <= 1'b1;
    layer2_outputs(175) <= not a or b;
    layer2_outputs(176) <= a and not b;
    layer2_outputs(177) <= not b or a;
    layer2_outputs(178) <= a and b;
    layer2_outputs(179) <= b;
    layer2_outputs(180) <= not a or b;
    layer2_outputs(181) <= not a or b;
    layer2_outputs(182) <= a xor b;
    layer2_outputs(183) <= b and not a;
    layer2_outputs(184) <= a;
    layer2_outputs(185) <= not b or a;
    layer2_outputs(186) <= not (a or b);
    layer2_outputs(187) <= not (a and b);
    layer2_outputs(188) <= 1'b0;
    layer2_outputs(189) <= b and not a;
    layer2_outputs(190) <= a and b;
    layer2_outputs(191) <= 1'b0;
    layer2_outputs(192) <= 1'b0;
    layer2_outputs(193) <= a;
    layer2_outputs(194) <= a or b;
    layer2_outputs(195) <= not (a and b);
    layer2_outputs(196) <= a;
    layer2_outputs(197) <= not a or b;
    layer2_outputs(198) <= not (a and b);
    layer2_outputs(199) <= 1'b1;
    layer2_outputs(200) <= not (a or b);
    layer2_outputs(201) <= a or b;
    layer2_outputs(202) <= a and b;
    layer2_outputs(203) <= not (a and b);
    layer2_outputs(204) <= not a;
    layer2_outputs(205) <= b and not a;
    layer2_outputs(206) <= not b;
    layer2_outputs(207) <= b and not a;
    layer2_outputs(208) <= not a or b;
    layer2_outputs(209) <= a xor b;
    layer2_outputs(210) <= b;
    layer2_outputs(211) <= not b or a;
    layer2_outputs(212) <= not b;
    layer2_outputs(213) <= a;
    layer2_outputs(214) <= b and not a;
    layer2_outputs(215) <= a;
    layer2_outputs(216) <= not b;
    layer2_outputs(217) <= a or b;
    layer2_outputs(218) <= b;
    layer2_outputs(219) <= a;
    layer2_outputs(220) <= a;
    layer2_outputs(221) <= 1'b0;
    layer2_outputs(222) <= a;
    layer2_outputs(223) <= a;
    layer2_outputs(224) <= a and not b;
    layer2_outputs(225) <= b;
    layer2_outputs(226) <= not a or b;
    layer2_outputs(227) <= a and not b;
    layer2_outputs(228) <= a or b;
    layer2_outputs(229) <= b and not a;
    layer2_outputs(230) <= a and b;
    layer2_outputs(231) <= not b;
    layer2_outputs(232) <= not a;
    layer2_outputs(233) <= b and not a;
    layer2_outputs(234) <= b;
    layer2_outputs(235) <= not b or a;
    layer2_outputs(236) <= not (a and b);
    layer2_outputs(237) <= not b;
    layer2_outputs(238) <= b and not a;
    layer2_outputs(239) <= a and not b;
    layer2_outputs(240) <= not (a or b);
    layer2_outputs(241) <= not a;
    layer2_outputs(242) <= not (a and b);
    layer2_outputs(243) <= not b;
    layer2_outputs(244) <= a and b;
    layer2_outputs(245) <= a;
    layer2_outputs(246) <= not a;
    layer2_outputs(247) <= a and not b;
    layer2_outputs(248) <= 1'b1;
    layer2_outputs(249) <= a or b;
    layer2_outputs(250) <= not a;
    layer2_outputs(251) <= not a;
    layer2_outputs(252) <= a;
    layer2_outputs(253) <= not a;
    layer2_outputs(254) <= a and not b;
    layer2_outputs(255) <= a or b;
    layer2_outputs(256) <= not a or b;
    layer2_outputs(257) <= a xor b;
    layer2_outputs(258) <= a;
    layer2_outputs(259) <= not (a or b);
    layer2_outputs(260) <= a;
    layer2_outputs(261) <= not b;
    layer2_outputs(262) <= 1'b0;
    layer2_outputs(263) <= not (a or b);
    layer2_outputs(264) <= not b or a;
    layer2_outputs(265) <= a and not b;
    layer2_outputs(266) <= not (a and b);
    layer2_outputs(267) <= a or b;
    layer2_outputs(268) <= a and b;
    layer2_outputs(269) <= a and b;
    layer2_outputs(270) <= not b;
    layer2_outputs(271) <= 1'b0;
    layer2_outputs(272) <= not b;
    layer2_outputs(273) <= 1'b1;
    layer2_outputs(274) <= a xor b;
    layer2_outputs(275) <= a;
    layer2_outputs(276) <= not (a and b);
    layer2_outputs(277) <= 1'b1;
    layer2_outputs(278) <= a;
    layer2_outputs(279) <= b;
    layer2_outputs(280) <= b and not a;
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= a or b;
    layer2_outputs(283) <= a and not b;
    layer2_outputs(284) <= not b or a;
    layer2_outputs(285) <= b;
    layer2_outputs(286) <= a and b;
    layer2_outputs(287) <= not a;
    layer2_outputs(288) <= not a;
    layer2_outputs(289) <= a;
    layer2_outputs(290) <= not b or a;
    layer2_outputs(291) <= a;
    layer2_outputs(292) <= a and not b;
    layer2_outputs(293) <= not b;
    layer2_outputs(294) <= not (a and b);
    layer2_outputs(295) <= b and not a;
    layer2_outputs(296) <= b and not a;
    layer2_outputs(297) <= 1'b0;
    layer2_outputs(298) <= not a or b;
    layer2_outputs(299) <= b;
    layer2_outputs(300) <= not b or a;
    layer2_outputs(301) <= a or b;
    layer2_outputs(302) <= not b;
    layer2_outputs(303) <= b and not a;
    layer2_outputs(304) <= b;
    layer2_outputs(305) <= not b;
    layer2_outputs(306) <= not b or a;
    layer2_outputs(307) <= a;
    layer2_outputs(308) <= not b or a;
    layer2_outputs(309) <= not a;
    layer2_outputs(310) <= 1'b1;
    layer2_outputs(311) <= not a;
    layer2_outputs(312) <= a and b;
    layer2_outputs(313) <= not a;
    layer2_outputs(314) <= not a;
    layer2_outputs(315) <= not (a and b);
    layer2_outputs(316) <= not a;
    layer2_outputs(317) <= not b or a;
    layer2_outputs(318) <= a and b;
    layer2_outputs(319) <= not b;
    layer2_outputs(320) <= a or b;
    layer2_outputs(321) <= a or b;
    layer2_outputs(322) <= 1'b1;
    layer2_outputs(323) <= not b;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= a xor b;
    layer2_outputs(326) <= a;
    layer2_outputs(327) <= not (a and b);
    layer2_outputs(328) <= not b or a;
    layer2_outputs(329) <= not (a and b);
    layer2_outputs(330) <= not a or b;
    layer2_outputs(331) <= b and not a;
    layer2_outputs(332) <= b and not a;
    layer2_outputs(333) <= 1'b0;
    layer2_outputs(334) <= b;
    layer2_outputs(335) <= a and not b;
    layer2_outputs(336) <= a and b;
    layer2_outputs(337) <= a;
    layer2_outputs(338) <= a or b;
    layer2_outputs(339) <= 1'b0;
    layer2_outputs(340) <= b and not a;
    layer2_outputs(341) <= 1'b0;
    layer2_outputs(342) <= not a;
    layer2_outputs(343) <= 1'b0;
    layer2_outputs(344) <= a;
    layer2_outputs(345) <= not a or b;
    layer2_outputs(346) <= not b;
    layer2_outputs(347) <= b and not a;
    layer2_outputs(348) <= not b or a;
    layer2_outputs(349) <= not a;
    layer2_outputs(350) <= not (a and b);
    layer2_outputs(351) <= not b;
    layer2_outputs(352) <= a and b;
    layer2_outputs(353) <= not b or a;
    layer2_outputs(354) <= b;
    layer2_outputs(355) <= a;
    layer2_outputs(356) <= not b;
    layer2_outputs(357) <= not b;
    layer2_outputs(358) <= a or b;
    layer2_outputs(359) <= a;
    layer2_outputs(360) <= b and not a;
    layer2_outputs(361) <= a;
    layer2_outputs(362) <= b;
    layer2_outputs(363) <= not (a or b);
    layer2_outputs(364) <= not (a and b);
    layer2_outputs(365) <= b and not a;
    layer2_outputs(366) <= a and not b;
    layer2_outputs(367) <= b;
    layer2_outputs(368) <= b and not a;
    layer2_outputs(369) <= a and b;
    layer2_outputs(370) <= a or b;
    layer2_outputs(371) <= not a or b;
    layer2_outputs(372) <= a and b;
    layer2_outputs(373) <= not a;
    layer2_outputs(374) <= a;
    layer2_outputs(375) <= a;
    layer2_outputs(376) <= 1'b0;
    layer2_outputs(377) <= not b;
    layer2_outputs(378) <= a and b;
    layer2_outputs(379) <= not b;
    layer2_outputs(380) <= a;
    layer2_outputs(381) <= not b or a;
    layer2_outputs(382) <= b and not a;
    layer2_outputs(383) <= not a;
    layer2_outputs(384) <= not b;
    layer2_outputs(385) <= b and not a;
    layer2_outputs(386) <= a and b;
    layer2_outputs(387) <= a or b;
    layer2_outputs(388) <= a and not b;
    layer2_outputs(389) <= not b or a;
    layer2_outputs(390) <= not b;
    layer2_outputs(391) <= not (a or b);
    layer2_outputs(392) <= not a or b;
    layer2_outputs(393) <= b and not a;
    layer2_outputs(394) <= a;
    layer2_outputs(395) <= not (a or b);
    layer2_outputs(396) <= 1'b1;
    layer2_outputs(397) <= a and b;
    layer2_outputs(398) <= b and not a;
    layer2_outputs(399) <= 1'b0;
    layer2_outputs(400) <= not (a or b);
    layer2_outputs(401) <= b and not a;
    layer2_outputs(402) <= not b;
    layer2_outputs(403) <= not (a and b);
    layer2_outputs(404) <= b;
    layer2_outputs(405) <= not a or b;
    layer2_outputs(406) <= not b or a;
    layer2_outputs(407) <= a and b;
    layer2_outputs(408) <= a xor b;
    layer2_outputs(409) <= b;
    layer2_outputs(410) <= a and b;
    layer2_outputs(411) <= 1'b1;
    layer2_outputs(412) <= not (a and b);
    layer2_outputs(413) <= a;
    layer2_outputs(414) <= not (a or b);
    layer2_outputs(415) <= not (a xor b);
    layer2_outputs(416) <= b;
    layer2_outputs(417) <= b;
    layer2_outputs(418) <= a and not b;
    layer2_outputs(419) <= not b;
    layer2_outputs(420) <= not a;
    layer2_outputs(421) <= b and not a;
    layer2_outputs(422) <= not a or b;
    layer2_outputs(423) <= not (a xor b);
    layer2_outputs(424) <= not (a or b);
    layer2_outputs(425) <= a xor b;
    layer2_outputs(426) <= not (a or b);
    layer2_outputs(427) <= b and not a;
    layer2_outputs(428) <= not (a and b);
    layer2_outputs(429) <= 1'b0;
    layer2_outputs(430) <= not (a or b);
    layer2_outputs(431) <= b and not a;
    layer2_outputs(432) <= not (a xor b);
    layer2_outputs(433) <= b;
    layer2_outputs(434) <= not b or a;
    layer2_outputs(435) <= not (a or b);
    layer2_outputs(436) <= 1'b1;
    layer2_outputs(437) <= not b or a;
    layer2_outputs(438) <= b;
    layer2_outputs(439) <= a or b;
    layer2_outputs(440) <= not b or a;
    layer2_outputs(441) <= a or b;
    layer2_outputs(442) <= not (a or b);
    layer2_outputs(443) <= a;
    layer2_outputs(444) <= not a or b;
    layer2_outputs(445) <= a xor b;
    layer2_outputs(446) <= not b;
    layer2_outputs(447) <= 1'b1;
    layer2_outputs(448) <= not a or b;
    layer2_outputs(449) <= a or b;
    layer2_outputs(450) <= not b;
    layer2_outputs(451) <= b and not a;
    layer2_outputs(452) <= not b;
    layer2_outputs(453) <= a or b;
    layer2_outputs(454) <= not b;
    layer2_outputs(455) <= not b;
    layer2_outputs(456) <= not (a and b);
    layer2_outputs(457) <= not (a or b);
    layer2_outputs(458) <= a;
    layer2_outputs(459) <= not (a or b);
    layer2_outputs(460) <= not b or a;
    layer2_outputs(461) <= a or b;
    layer2_outputs(462) <= not b;
    layer2_outputs(463) <= a and not b;
    layer2_outputs(464) <= not (a and b);
    layer2_outputs(465) <= not (a xor b);
    layer2_outputs(466) <= not (a and b);
    layer2_outputs(467) <= a and not b;
    layer2_outputs(468) <= not (a or b);
    layer2_outputs(469) <= not a;
    layer2_outputs(470) <= a or b;
    layer2_outputs(471) <= a;
    layer2_outputs(472) <= b and not a;
    layer2_outputs(473) <= 1'b1;
    layer2_outputs(474) <= not a;
    layer2_outputs(475) <= 1'b0;
    layer2_outputs(476) <= b and not a;
    layer2_outputs(477) <= not a;
    layer2_outputs(478) <= not a or b;
    layer2_outputs(479) <= b and not a;
    layer2_outputs(480) <= not b;
    layer2_outputs(481) <= not a;
    layer2_outputs(482) <= not b;
    layer2_outputs(483) <= not b;
    layer2_outputs(484) <= b;
    layer2_outputs(485) <= b;
    layer2_outputs(486) <= not b;
    layer2_outputs(487) <= not a;
    layer2_outputs(488) <= a or b;
    layer2_outputs(489) <= not a;
    layer2_outputs(490) <= not (a or b);
    layer2_outputs(491) <= not a;
    layer2_outputs(492) <= not b or a;
    layer2_outputs(493) <= b;
    layer2_outputs(494) <= not (a and b);
    layer2_outputs(495) <= a or b;
    layer2_outputs(496) <= not (a and b);
    layer2_outputs(497) <= b;
    layer2_outputs(498) <= not a;
    layer2_outputs(499) <= not b;
    layer2_outputs(500) <= a or b;
    layer2_outputs(501) <= not a;
    layer2_outputs(502) <= b and not a;
    layer2_outputs(503) <= not b;
    layer2_outputs(504) <= not (a and b);
    layer2_outputs(505) <= b;
    layer2_outputs(506) <= not b;
    layer2_outputs(507) <= not (a and b);
    layer2_outputs(508) <= not b or a;
    layer2_outputs(509) <= not b or a;
    layer2_outputs(510) <= a or b;
    layer2_outputs(511) <= b and not a;
    layer2_outputs(512) <= not (a and b);
    layer2_outputs(513) <= not (a and b);
    layer2_outputs(514) <= b;
    layer2_outputs(515) <= b;
    layer2_outputs(516) <= not a;
    layer2_outputs(517) <= not a;
    layer2_outputs(518) <= not (a or b);
    layer2_outputs(519) <= b;
    layer2_outputs(520) <= a;
    layer2_outputs(521) <= 1'b1;
    layer2_outputs(522) <= a and not b;
    layer2_outputs(523) <= not (a xor b);
    layer2_outputs(524) <= not b or a;
    layer2_outputs(525) <= not (a and b);
    layer2_outputs(526) <= 1'b1;
    layer2_outputs(527) <= not b or a;
    layer2_outputs(528) <= not b or a;
    layer2_outputs(529) <= not (a xor b);
    layer2_outputs(530) <= not a or b;
    layer2_outputs(531) <= not b;
    layer2_outputs(532) <= not (a or b);
    layer2_outputs(533) <= not a or b;
    layer2_outputs(534) <= not (a or b);
    layer2_outputs(535) <= not a or b;
    layer2_outputs(536) <= not (a or b);
    layer2_outputs(537) <= b and not a;
    layer2_outputs(538) <= a;
    layer2_outputs(539) <= not a or b;
    layer2_outputs(540) <= 1'b1;
    layer2_outputs(541) <= not (a xor b);
    layer2_outputs(542) <= 1'b0;
    layer2_outputs(543) <= a;
    layer2_outputs(544) <= a and not b;
    layer2_outputs(545) <= a or b;
    layer2_outputs(546) <= a and not b;
    layer2_outputs(547) <= a and b;
    layer2_outputs(548) <= a or b;
    layer2_outputs(549) <= b;
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= a and b;
    layer2_outputs(552) <= a;
    layer2_outputs(553) <= not a or b;
    layer2_outputs(554) <= not a;
    layer2_outputs(555) <= not b;
    layer2_outputs(556) <= a and not b;
    layer2_outputs(557) <= b and not a;
    layer2_outputs(558) <= not (a and b);
    layer2_outputs(559) <= b;
    layer2_outputs(560) <= not b;
    layer2_outputs(561) <= a or b;
    layer2_outputs(562) <= a xor b;
    layer2_outputs(563) <= a and b;
    layer2_outputs(564) <= a xor b;
    layer2_outputs(565) <= not a or b;
    layer2_outputs(566) <= not b;
    layer2_outputs(567) <= not (a xor b);
    layer2_outputs(568) <= a or b;
    layer2_outputs(569) <= not (a or b);
    layer2_outputs(570) <= a;
    layer2_outputs(571) <= b and not a;
    layer2_outputs(572) <= a or b;
    layer2_outputs(573) <= a xor b;
    layer2_outputs(574) <= a and b;
    layer2_outputs(575) <= not a;
    layer2_outputs(576) <= not (a xor b);
    layer2_outputs(577) <= not (a and b);
    layer2_outputs(578) <= not a;
    layer2_outputs(579) <= not (a and b);
    layer2_outputs(580) <= a and not b;
    layer2_outputs(581) <= a;
    layer2_outputs(582) <= a and b;
    layer2_outputs(583) <= not (a or b);
    layer2_outputs(584) <= a;
    layer2_outputs(585) <= a;
    layer2_outputs(586) <= not a;
    layer2_outputs(587) <= not b;
    layer2_outputs(588) <= a and not b;
    layer2_outputs(589) <= not (a and b);
    layer2_outputs(590) <= not (a and b);
    layer2_outputs(591) <= not b;
    layer2_outputs(592) <= not b or a;
    layer2_outputs(593) <= b and not a;
    layer2_outputs(594) <= a;
    layer2_outputs(595) <= a and b;
    layer2_outputs(596) <= a and b;
    layer2_outputs(597) <= a;
    layer2_outputs(598) <= a and b;
    layer2_outputs(599) <= not b;
    layer2_outputs(600) <= not b;
    layer2_outputs(601) <= not (a and b);
    layer2_outputs(602) <= b and not a;
    layer2_outputs(603) <= b and not a;
    layer2_outputs(604) <= 1'b0;
    layer2_outputs(605) <= a and b;
    layer2_outputs(606) <= b;
    layer2_outputs(607) <= b;
    layer2_outputs(608) <= not b;
    layer2_outputs(609) <= not b;
    layer2_outputs(610) <= a;
    layer2_outputs(611) <= not (a xor b);
    layer2_outputs(612) <= a or b;
    layer2_outputs(613) <= not b;
    layer2_outputs(614) <= a;
    layer2_outputs(615) <= not (a xor b);
    layer2_outputs(616) <= not b;
    layer2_outputs(617) <= not b or a;
    layer2_outputs(618) <= not a or b;
    layer2_outputs(619) <= not b;
    layer2_outputs(620) <= not a or b;
    layer2_outputs(621) <= b;
    layer2_outputs(622) <= b;
    layer2_outputs(623) <= not b or a;
    layer2_outputs(624) <= not a;
    layer2_outputs(625) <= a;
    layer2_outputs(626) <= not b;
    layer2_outputs(627) <= not b;
    layer2_outputs(628) <= not b;
    layer2_outputs(629) <= b;
    layer2_outputs(630) <= a or b;
    layer2_outputs(631) <= a;
    layer2_outputs(632) <= not (a or b);
    layer2_outputs(633) <= a;
    layer2_outputs(634) <= a or b;
    layer2_outputs(635) <= b and not a;
    layer2_outputs(636) <= not b;
    layer2_outputs(637) <= not (a and b);
    layer2_outputs(638) <= a;
    layer2_outputs(639) <= a and b;
    layer2_outputs(640) <= not (a or b);
    layer2_outputs(641) <= 1'b1;
    layer2_outputs(642) <= not b;
    layer2_outputs(643) <= a and not b;
    layer2_outputs(644) <= not b;
    layer2_outputs(645) <= b;
    layer2_outputs(646) <= b;
    layer2_outputs(647) <= not a or b;
    layer2_outputs(648) <= not (a xor b);
    layer2_outputs(649) <= a and b;
    layer2_outputs(650) <= b;
    layer2_outputs(651) <= a and b;
    layer2_outputs(652) <= b;
    layer2_outputs(653) <= not b;
    layer2_outputs(654) <= a and b;
    layer2_outputs(655) <= not a;
    layer2_outputs(656) <= a or b;
    layer2_outputs(657) <= not a;
    layer2_outputs(658) <= not a or b;
    layer2_outputs(659) <= not (a and b);
    layer2_outputs(660) <= not a;
    layer2_outputs(661) <= not a;
    layer2_outputs(662) <= not b or a;
    layer2_outputs(663) <= not a;
    layer2_outputs(664) <= not (a xor b);
    layer2_outputs(665) <= b and not a;
    layer2_outputs(666) <= 1'b1;
    layer2_outputs(667) <= b;
    layer2_outputs(668) <= a and not b;
    layer2_outputs(669) <= not (a or b);
    layer2_outputs(670) <= not a;
    layer2_outputs(671) <= not (a and b);
    layer2_outputs(672) <= b and not a;
    layer2_outputs(673) <= not a or b;
    layer2_outputs(674) <= a;
    layer2_outputs(675) <= b and not a;
    layer2_outputs(676) <= a;
    layer2_outputs(677) <= not b;
    layer2_outputs(678) <= not b or a;
    layer2_outputs(679) <= a;
    layer2_outputs(680) <= a;
    layer2_outputs(681) <= a;
    layer2_outputs(682) <= a and not b;
    layer2_outputs(683) <= not (a or b);
    layer2_outputs(684) <= b;
    layer2_outputs(685) <= a;
    layer2_outputs(686) <= not a;
    layer2_outputs(687) <= 1'b0;
    layer2_outputs(688) <= b;
    layer2_outputs(689) <= a or b;
    layer2_outputs(690) <= not b;
    layer2_outputs(691) <= a;
    layer2_outputs(692) <= not (a and b);
    layer2_outputs(693) <= not (a and b);
    layer2_outputs(694) <= not b or a;
    layer2_outputs(695) <= not a or b;
    layer2_outputs(696) <= not a or b;
    layer2_outputs(697) <= a and b;
    layer2_outputs(698) <= a;
    layer2_outputs(699) <= b;
    layer2_outputs(700) <= not b;
    layer2_outputs(701) <= not a;
    layer2_outputs(702) <= a;
    layer2_outputs(703) <= not (a or b);
    layer2_outputs(704) <= a xor b;
    layer2_outputs(705) <= not (a and b);
    layer2_outputs(706) <= b;
    layer2_outputs(707) <= a;
    layer2_outputs(708) <= not a;
    layer2_outputs(709) <= a and b;
    layer2_outputs(710) <= not (a or b);
    layer2_outputs(711) <= a and not b;
    layer2_outputs(712) <= a and not b;
    layer2_outputs(713) <= b;
    layer2_outputs(714) <= a xor b;
    layer2_outputs(715) <= b;
    layer2_outputs(716) <= a;
    layer2_outputs(717) <= not b or a;
    layer2_outputs(718) <= not a or b;
    layer2_outputs(719) <= a and b;
    layer2_outputs(720) <= a and not b;
    layer2_outputs(721) <= not (a or b);
    layer2_outputs(722) <= not a or b;
    layer2_outputs(723) <= not (a or b);
    layer2_outputs(724) <= b and not a;
    layer2_outputs(725) <= b;
    layer2_outputs(726) <= not a;
    layer2_outputs(727) <= b;
    layer2_outputs(728) <= b;
    layer2_outputs(729) <= not (a or b);
    layer2_outputs(730) <= a and b;
    layer2_outputs(731) <= not (a and b);
    layer2_outputs(732) <= not a;
    layer2_outputs(733) <= 1'b1;
    layer2_outputs(734) <= b and not a;
    layer2_outputs(735) <= a and b;
    layer2_outputs(736) <= a or b;
    layer2_outputs(737) <= not (a and b);
    layer2_outputs(738) <= a and not b;
    layer2_outputs(739) <= b and not a;
    layer2_outputs(740) <= not (a or b);
    layer2_outputs(741) <= not a or b;
    layer2_outputs(742) <= b;
    layer2_outputs(743) <= not a or b;
    layer2_outputs(744) <= not (a xor b);
    layer2_outputs(745) <= not (a or b);
    layer2_outputs(746) <= a and not b;
    layer2_outputs(747) <= not (a or b);
    layer2_outputs(748) <= a and not b;
    layer2_outputs(749) <= 1'b1;
    layer2_outputs(750) <= b;
    layer2_outputs(751) <= not a or b;
    layer2_outputs(752) <= not b or a;
    layer2_outputs(753) <= 1'b0;
    layer2_outputs(754) <= not a or b;
    layer2_outputs(755) <= not a or b;
    layer2_outputs(756) <= not (a and b);
    layer2_outputs(757) <= a xor b;
    layer2_outputs(758) <= a or b;
    layer2_outputs(759) <= not (a and b);
    layer2_outputs(760) <= not (a or b);
    layer2_outputs(761) <= not a;
    layer2_outputs(762) <= a and b;
    layer2_outputs(763) <= not a;
    layer2_outputs(764) <= not b;
    layer2_outputs(765) <= a;
    layer2_outputs(766) <= a;
    layer2_outputs(767) <= not (a or b);
    layer2_outputs(768) <= not a;
    layer2_outputs(769) <= b;
    layer2_outputs(770) <= not (a or b);
    layer2_outputs(771) <= not a or b;
    layer2_outputs(772) <= a or b;
    layer2_outputs(773) <= a or b;
    layer2_outputs(774) <= a and b;
    layer2_outputs(775) <= not b or a;
    layer2_outputs(776) <= b and not a;
    layer2_outputs(777) <= a and not b;
    layer2_outputs(778) <= not b;
    layer2_outputs(779) <= not b;
    layer2_outputs(780) <= not b or a;
    layer2_outputs(781) <= not b;
    layer2_outputs(782) <= a or b;
    layer2_outputs(783) <= not b;
    layer2_outputs(784) <= b and not a;
    layer2_outputs(785) <= not a or b;
    layer2_outputs(786) <= a;
    layer2_outputs(787) <= not (a xor b);
    layer2_outputs(788) <= a or b;
    layer2_outputs(789) <= not a or b;
    layer2_outputs(790) <= a;
    layer2_outputs(791) <= not a;
    layer2_outputs(792) <= a and b;
    layer2_outputs(793) <= a or b;
    layer2_outputs(794) <= not b or a;
    layer2_outputs(795) <= b and not a;
    layer2_outputs(796) <= not a;
    layer2_outputs(797) <= not (a or b);
    layer2_outputs(798) <= b and not a;
    layer2_outputs(799) <= not b;
    layer2_outputs(800) <= a and b;
    layer2_outputs(801) <= not a;
    layer2_outputs(802) <= not b;
    layer2_outputs(803) <= not b;
    layer2_outputs(804) <= not (a or b);
    layer2_outputs(805) <= not (a xor b);
    layer2_outputs(806) <= not b;
    layer2_outputs(807) <= not b or a;
    layer2_outputs(808) <= a;
    layer2_outputs(809) <= not b;
    layer2_outputs(810) <= a or b;
    layer2_outputs(811) <= 1'b0;
    layer2_outputs(812) <= a;
    layer2_outputs(813) <= a or b;
    layer2_outputs(814) <= not a;
    layer2_outputs(815) <= a and b;
    layer2_outputs(816) <= not b;
    layer2_outputs(817) <= not a;
    layer2_outputs(818) <= 1'b1;
    layer2_outputs(819) <= not b;
    layer2_outputs(820) <= a and b;
    layer2_outputs(821) <= not a;
    layer2_outputs(822) <= a and b;
    layer2_outputs(823) <= a xor b;
    layer2_outputs(824) <= 1'b0;
    layer2_outputs(825) <= not b;
    layer2_outputs(826) <= a or b;
    layer2_outputs(827) <= a xor b;
    layer2_outputs(828) <= not b or a;
    layer2_outputs(829) <= b and not a;
    layer2_outputs(830) <= not b;
    layer2_outputs(831) <= not (a or b);
    layer2_outputs(832) <= not a;
    layer2_outputs(833) <= a and not b;
    layer2_outputs(834) <= a and b;
    layer2_outputs(835) <= b;
    layer2_outputs(836) <= not (a or b);
    layer2_outputs(837) <= a;
    layer2_outputs(838) <= not a;
    layer2_outputs(839) <= not b;
    layer2_outputs(840) <= not a;
    layer2_outputs(841) <= a and b;
    layer2_outputs(842) <= a;
    layer2_outputs(843) <= b;
    layer2_outputs(844) <= not b or a;
    layer2_outputs(845) <= 1'b1;
    layer2_outputs(846) <= a;
    layer2_outputs(847) <= not (a and b);
    layer2_outputs(848) <= a and not b;
    layer2_outputs(849) <= b;
    layer2_outputs(850) <= not (a or b);
    layer2_outputs(851) <= 1'b1;
    layer2_outputs(852) <= a xor b;
    layer2_outputs(853) <= a or b;
    layer2_outputs(854) <= a and not b;
    layer2_outputs(855) <= a or b;
    layer2_outputs(856) <= not b or a;
    layer2_outputs(857) <= 1'b1;
    layer2_outputs(858) <= b;
    layer2_outputs(859) <= a xor b;
    layer2_outputs(860) <= not a;
    layer2_outputs(861) <= a and b;
    layer2_outputs(862) <= a or b;
    layer2_outputs(863) <= a;
    layer2_outputs(864) <= not b;
    layer2_outputs(865) <= b;
    layer2_outputs(866) <= not b;
    layer2_outputs(867) <= not b;
    layer2_outputs(868) <= not (a and b);
    layer2_outputs(869) <= b;
    layer2_outputs(870) <= not (a or b);
    layer2_outputs(871) <= a;
    layer2_outputs(872) <= a or b;
    layer2_outputs(873) <= not (a or b);
    layer2_outputs(874) <= a;
    layer2_outputs(875) <= a;
    layer2_outputs(876) <= not a or b;
    layer2_outputs(877) <= not (a and b);
    layer2_outputs(878) <= not (a and b);
    layer2_outputs(879) <= a xor b;
    layer2_outputs(880) <= a or b;
    layer2_outputs(881) <= a or b;
    layer2_outputs(882) <= not a;
    layer2_outputs(883) <= not b or a;
    layer2_outputs(884) <= not a;
    layer2_outputs(885) <= not a or b;
    layer2_outputs(886) <= not a or b;
    layer2_outputs(887) <= not a or b;
    layer2_outputs(888) <= not a or b;
    layer2_outputs(889) <= a xor b;
    layer2_outputs(890) <= 1'b1;
    layer2_outputs(891) <= a;
    layer2_outputs(892) <= not (a or b);
    layer2_outputs(893) <= not (a and b);
    layer2_outputs(894) <= not b or a;
    layer2_outputs(895) <= b;
    layer2_outputs(896) <= not a;
    layer2_outputs(897) <= a or b;
    layer2_outputs(898) <= not b;
    layer2_outputs(899) <= not b;
    layer2_outputs(900) <= b;
    layer2_outputs(901) <= 1'b0;
    layer2_outputs(902) <= not (a and b);
    layer2_outputs(903) <= a and not b;
    layer2_outputs(904) <= a and b;
    layer2_outputs(905) <= 1'b0;
    layer2_outputs(906) <= not a;
    layer2_outputs(907) <= a;
    layer2_outputs(908) <= b;
    layer2_outputs(909) <= b;
    layer2_outputs(910) <= a;
    layer2_outputs(911) <= not b;
    layer2_outputs(912) <= not a or b;
    layer2_outputs(913) <= not a;
    layer2_outputs(914) <= not (a or b);
    layer2_outputs(915) <= a and not b;
    layer2_outputs(916) <= not b or a;
    layer2_outputs(917) <= not b;
    layer2_outputs(918) <= a or b;
    layer2_outputs(919) <= 1'b0;
    layer2_outputs(920) <= not (a or b);
    layer2_outputs(921) <= b and not a;
    layer2_outputs(922) <= b and not a;
    layer2_outputs(923) <= not a or b;
    layer2_outputs(924) <= a and b;
    layer2_outputs(925) <= not (a and b);
    layer2_outputs(926) <= a or b;
    layer2_outputs(927) <= 1'b0;
    layer2_outputs(928) <= not (a or b);
    layer2_outputs(929) <= not (a xor b);
    layer2_outputs(930) <= not a or b;
    layer2_outputs(931) <= 1'b1;
    layer2_outputs(932) <= a and not b;
    layer2_outputs(933) <= not (a or b);
    layer2_outputs(934) <= a and b;
    layer2_outputs(935) <= not b or a;
    layer2_outputs(936) <= b and not a;
    layer2_outputs(937) <= not a;
    layer2_outputs(938) <= b;
    layer2_outputs(939) <= b;
    layer2_outputs(940) <= not a;
    layer2_outputs(941) <= not (a xor b);
    layer2_outputs(942) <= not a or b;
    layer2_outputs(943) <= b;
    layer2_outputs(944) <= a;
    layer2_outputs(945) <= not (a or b);
    layer2_outputs(946) <= b;
    layer2_outputs(947) <= a or b;
    layer2_outputs(948) <= not a;
    layer2_outputs(949) <= not a or b;
    layer2_outputs(950) <= b and not a;
    layer2_outputs(951) <= b;
    layer2_outputs(952) <= not (a xor b);
    layer2_outputs(953) <= a and not b;
    layer2_outputs(954) <= not b;
    layer2_outputs(955) <= a and b;
    layer2_outputs(956) <= a and not b;
    layer2_outputs(957) <= not (a and b);
    layer2_outputs(958) <= 1'b0;
    layer2_outputs(959) <= a and not b;
    layer2_outputs(960) <= not b or a;
    layer2_outputs(961) <= b and not a;
    layer2_outputs(962) <= not (a and b);
    layer2_outputs(963) <= not b or a;
    layer2_outputs(964) <= b and not a;
    layer2_outputs(965) <= a and b;
    layer2_outputs(966) <= not (a or b);
    layer2_outputs(967) <= not (a or b);
    layer2_outputs(968) <= not (a or b);
    layer2_outputs(969) <= b;
    layer2_outputs(970) <= b;
    layer2_outputs(971) <= not a;
    layer2_outputs(972) <= a;
    layer2_outputs(973) <= 1'b0;
    layer2_outputs(974) <= not a;
    layer2_outputs(975) <= a or b;
    layer2_outputs(976) <= not a or b;
    layer2_outputs(977) <= not a or b;
    layer2_outputs(978) <= b and not a;
    layer2_outputs(979) <= 1'b1;
    layer2_outputs(980) <= a xor b;
    layer2_outputs(981) <= a;
    layer2_outputs(982) <= not b or a;
    layer2_outputs(983) <= a and not b;
    layer2_outputs(984) <= a or b;
    layer2_outputs(985) <= b;
    layer2_outputs(986) <= a and b;
    layer2_outputs(987) <= 1'b0;
    layer2_outputs(988) <= not a;
    layer2_outputs(989) <= a;
    layer2_outputs(990) <= not a;
    layer2_outputs(991) <= not a;
    layer2_outputs(992) <= not b;
    layer2_outputs(993) <= not b or a;
    layer2_outputs(994) <= a and b;
    layer2_outputs(995) <= not b or a;
    layer2_outputs(996) <= a xor b;
    layer2_outputs(997) <= b and not a;
    layer2_outputs(998) <= a;
    layer2_outputs(999) <= a;
    layer2_outputs(1000) <= not a;
    layer2_outputs(1001) <= not (a and b);
    layer2_outputs(1002) <= not (a xor b);
    layer2_outputs(1003) <= b;
    layer2_outputs(1004) <= a;
    layer2_outputs(1005) <= a and not b;
    layer2_outputs(1006) <= not b;
    layer2_outputs(1007) <= not b or a;
    layer2_outputs(1008) <= b;
    layer2_outputs(1009) <= a;
    layer2_outputs(1010) <= not a or b;
    layer2_outputs(1011) <= not b;
    layer2_outputs(1012) <= not b or a;
    layer2_outputs(1013) <= not a;
    layer2_outputs(1014) <= not a;
    layer2_outputs(1015) <= b and not a;
    layer2_outputs(1016) <= not a or b;
    layer2_outputs(1017) <= not b or a;
    layer2_outputs(1018) <= a and not b;
    layer2_outputs(1019) <= a or b;
    layer2_outputs(1020) <= not a;
    layer2_outputs(1021) <= b and not a;
    layer2_outputs(1022) <= b;
    layer2_outputs(1023) <= a or b;
    layer2_outputs(1024) <= 1'b0;
    layer2_outputs(1025) <= a and b;
    layer2_outputs(1026) <= not (a and b);
    layer2_outputs(1027) <= 1'b1;
    layer2_outputs(1028) <= not (a or b);
    layer2_outputs(1029) <= a or b;
    layer2_outputs(1030) <= a;
    layer2_outputs(1031) <= not a or b;
    layer2_outputs(1032) <= b;
    layer2_outputs(1033) <= not b;
    layer2_outputs(1034) <= not a;
    layer2_outputs(1035) <= a and b;
    layer2_outputs(1036) <= not b or a;
    layer2_outputs(1037) <= a and not b;
    layer2_outputs(1038) <= not (a or b);
    layer2_outputs(1039) <= not a or b;
    layer2_outputs(1040) <= a;
    layer2_outputs(1041) <= 1'b0;
    layer2_outputs(1042) <= a or b;
    layer2_outputs(1043) <= not b or a;
    layer2_outputs(1044) <= not a;
    layer2_outputs(1045) <= not a;
    layer2_outputs(1046) <= a and not b;
    layer2_outputs(1047) <= a or b;
    layer2_outputs(1048) <= a or b;
    layer2_outputs(1049) <= not a or b;
    layer2_outputs(1050) <= a and not b;
    layer2_outputs(1051) <= not a or b;
    layer2_outputs(1052) <= not a or b;
    layer2_outputs(1053) <= not a;
    layer2_outputs(1054) <= not a;
    layer2_outputs(1055) <= b;
    layer2_outputs(1056) <= not a;
    layer2_outputs(1057) <= a;
    layer2_outputs(1058) <= b;
    layer2_outputs(1059) <= not (a or b);
    layer2_outputs(1060) <= not b or a;
    layer2_outputs(1061) <= not (a and b);
    layer2_outputs(1062) <= 1'b0;
    layer2_outputs(1063) <= a;
    layer2_outputs(1064) <= not (a and b);
    layer2_outputs(1065) <= b and not a;
    layer2_outputs(1066) <= not (a and b);
    layer2_outputs(1067) <= not (a or b);
    layer2_outputs(1068) <= a and b;
    layer2_outputs(1069) <= a and b;
    layer2_outputs(1070) <= 1'b1;
    layer2_outputs(1071) <= not (a xor b);
    layer2_outputs(1072) <= not (a and b);
    layer2_outputs(1073) <= not b or a;
    layer2_outputs(1074) <= not b;
    layer2_outputs(1075) <= a and not b;
    layer2_outputs(1076) <= not b or a;
    layer2_outputs(1077) <= a or b;
    layer2_outputs(1078) <= not a;
    layer2_outputs(1079) <= not a;
    layer2_outputs(1080) <= not a;
    layer2_outputs(1081) <= 1'b0;
    layer2_outputs(1082) <= a;
    layer2_outputs(1083) <= not b;
    layer2_outputs(1084) <= not b;
    layer2_outputs(1085) <= not (a or b);
    layer2_outputs(1086) <= not (a xor b);
    layer2_outputs(1087) <= not b;
    layer2_outputs(1088) <= not a;
    layer2_outputs(1089) <= a and b;
    layer2_outputs(1090) <= a xor b;
    layer2_outputs(1091) <= not b or a;
    layer2_outputs(1092) <= 1'b0;
    layer2_outputs(1093) <= not a;
    layer2_outputs(1094) <= not (a or b);
    layer2_outputs(1095) <= b;
    layer2_outputs(1096) <= b and not a;
    layer2_outputs(1097) <= not a;
    layer2_outputs(1098) <= not a or b;
    layer2_outputs(1099) <= b;
    layer2_outputs(1100) <= not (a or b);
    layer2_outputs(1101) <= not a;
    layer2_outputs(1102) <= not a;
    layer2_outputs(1103) <= a and b;
    layer2_outputs(1104) <= not a;
    layer2_outputs(1105) <= b;
    layer2_outputs(1106) <= not (a and b);
    layer2_outputs(1107) <= a and not b;
    layer2_outputs(1108) <= a;
    layer2_outputs(1109) <= not b;
    layer2_outputs(1110) <= not a;
    layer2_outputs(1111) <= not a or b;
    layer2_outputs(1112) <= not a;
    layer2_outputs(1113) <= not b or a;
    layer2_outputs(1114) <= b and not a;
    layer2_outputs(1115) <= not (a and b);
    layer2_outputs(1116) <= not a or b;
    layer2_outputs(1117) <= b;
    layer2_outputs(1118) <= b and not a;
    layer2_outputs(1119) <= not b;
    layer2_outputs(1120) <= 1'b1;
    layer2_outputs(1121) <= a or b;
    layer2_outputs(1122) <= a;
    layer2_outputs(1123) <= b;
    layer2_outputs(1124) <= a;
    layer2_outputs(1125) <= b;
    layer2_outputs(1126) <= b;
    layer2_outputs(1127) <= b;
    layer2_outputs(1128) <= not (a xor b);
    layer2_outputs(1129) <= a;
    layer2_outputs(1130) <= a or b;
    layer2_outputs(1131) <= a or b;
    layer2_outputs(1132) <= not (a xor b);
    layer2_outputs(1133) <= not (a or b);
    layer2_outputs(1134) <= a;
    layer2_outputs(1135) <= not a;
    layer2_outputs(1136) <= 1'b1;
    layer2_outputs(1137) <= not (a and b);
    layer2_outputs(1138) <= not a or b;
    layer2_outputs(1139) <= not b;
    layer2_outputs(1140) <= b and not a;
    layer2_outputs(1141) <= not b;
    layer2_outputs(1142) <= a and b;
    layer2_outputs(1143) <= not b or a;
    layer2_outputs(1144) <= not (a and b);
    layer2_outputs(1145) <= not a;
    layer2_outputs(1146) <= not (a xor b);
    layer2_outputs(1147) <= a and not b;
    layer2_outputs(1148) <= a xor b;
    layer2_outputs(1149) <= a and b;
    layer2_outputs(1150) <= 1'b1;
    layer2_outputs(1151) <= a;
    layer2_outputs(1152) <= not b;
    layer2_outputs(1153) <= b;
    layer2_outputs(1154) <= not (a or b);
    layer2_outputs(1155) <= not (a xor b);
    layer2_outputs(1156) <= 1'b0;
    layer2_outputs(1157) <= b;
    layer2_outputs(1158) <= not b;
    layer2_outputs(1159) <= b;
    layer2_outputs(1160) <= not (a and b);
    layer2_outputs(1161) <= a xor b;
    layer2_outputs(1162) <= a and not b;
    layer2_outputs(1163) <= a xor b;
    layer2_outputs(1164) <= b;
    layer2_outputs(1165) <= not a or b;
    layer2_outputs(1166) <= b and not a;
    layer2_outputs(1167) <= not a;
    layer2_outputs(1168) <= b;
    layer2_outputs(1169) <= a or b;
    layer2_outputs(1170) <= not (a and b);
    layer2_outputs(1171) <= a xor b;
    layer2_outputs(1172) <= 1'b0;
    layer2_outputs(1173) <= not b or a;
    layer2_outputs(1174) <= a or b;
    layer2_outputs(1175) <= not (a and b);
    layer2_outputs(1176) <= b;
    layer2_outputs(1177) <= a;
    layer2_outputs(1178) <= not (a and b);
    layer2_outputs(1179) <= not (a and b);
    layer2_outputs(1180) <= not b;
    layer2_outputs(1181) <= b and not a;
    layer2_outputs(1182) <= not (a xor b);
    layer2_outputs(1183) <= a;
    layer2_outputs(1184) <= not (a or b);
    layer2_outputs(1185) <= a;
    layer2_outputs(1186) <= b and not a;
    layer2_outputs(1187) <= not (a or b);
    layer2_outputs(1188) <= a and not b;
    layer2_outputs(1189) <= not a;
    layer2_outputs(1190) <= not (a or b);
    layer2_outputs(1191) <= b;
    layer2_outputs(1192) <= a;
    layer2_outputs(1193) <= not (a and b);
    layer2_outputs(1194) <= not b or a;
    layer2_outputs(1195) <= not a;
    layer2_outputs(1196) <= b;
    layer2_outputs(1197) <= not (a or b);
    layer2_outputs(1198) <= a;
    layer2_outputs(1199) <= b;
    layer2_outputs(1200) <= a and not b;
    layer2_outputs(1201) <= a and b;
    layer2_outputs(1202) <= b;
    layer2_outputs(1203) <= not a;
    layer2_outputs(1204) <= a and not b;
    layer2_outputs(1205) <= b;
    layer2_outputs(1206) <= b;
    layer2_outputs(1207) <= not b;
    layer2_outputs(1208) <= not b or a;
    layer2_outputs(1209) <= b and not a;
    layer2_outputs(1210) <= a and not b;
    layer2_outputs(1211) <= a or b;
    layer2_outputs(1212) <= not (a and b);
    layer2_outputs(1213) <= b;
    layer2_outputs(1214) <= not b or a;
    layer2_outputs(1215) <= a and b;
    layer2_outputs(1216) <= a and b;
    layer2_outputs(1217) <= not a or b;
    layer2_outputs(1218) <= not a or b;
    layer2_outputs(1219) <= a and not b;
    layer2_outputs(1220) <= not a;
    layer2_outputs(1221) <= not a or b;
    layer2_outputs(1222) <= 1'b1;
    layer2_outputs(1223) <= not a or b;
    layer2_outputs(1224) <= not b or a;
    layer2_outputs(1225) <= a xor b;
    layer2_outputs(1226) <= b;
    layer2_outputs(1227) <= not a or b;
    layer2_outputs(1228) <= not b;
    layer2_outputs(1229) <= not b or a;
    layer2_outputs(1230) <= a;
    layer2_outputs(1231) <= not b or a;
    layer2_outputs(1232) <= b and not a;
    layer2_outputs(1233) <= not (a or b);
    layer2_outputs(1234) <= 1'b0;
    layer2_outputs(1235) <= b;
    layer2_outputs(1236) <= 1'b0;
    layer2_outputs(1237) <= not b;
    layer2_outputs(1238) <= not b;
    layer2_outputs(1239) <= not a;
    layer2_outputs(1240) <= a and b;
    layer2_outputs(1241) <= not a;
    layer2_outputs(1242) <= not (a or b);
    layer2_outputs(1243) <= a xor b;
    layer2_outputs(1244) <= not b;
    layer2_outputs(1245) <= b;
    layer2_outputs(1246) <= a or b;
    layer2_outputs(1247) <= not b or a;
    layer2_outputs(1248) <= not b or a;
    layer2_outputs(1249) <= a and not b;
    layer2_outputs(1250) <= a or b;
    layer2_outputs(1251) <= not b or a;
    layer2_outputs(1252) <= not (a or b);
    layer2_outputs(1253) <= a and b;
    layer2_outputs(1254) <= a and not b;
    layer2_outputs(1255) <= 1'b1;
    layer2_outputs(1256) <= not a;
    layer2_outputs(1257) <= not (a or b);
    layer2_outputs(1258) <= not b or a;
    layer2_outputs(1259) <= a and not b;
    layer2_outputs(1260) <= not a;
    layer2_outputs(1261) <= a and b;
    layer2_outputs(1262) <= a and not b;
    layer2_outputs(1263) <= b;
    layer2_outputs(1264) <= 1'b1;
    layer2_outputs(1265) <= not a;
    layer2_outputs(1266) <= not b;
    layer2_outputs(1267) <= b;
    layer2_outputs(1268) <= a or b;
    layer2_outputs(1269) <= b;
    layer2_outputs(1270) <= not (a or b);
    layer2_outputs(1271) <= not b;
    layer2_outputs(1272) <= not a or b;
    layer2_outputs(1273) <= not (a or b);
    layer2_outputs(1274) <= 1'b1;
    layer2_outputs(1275) <= a;
    layer2_outputs(1276) <= a or b;
    layer2_outputs(1277) <= 1'b1;
    layer2_outputs(1278) <= a and b;
    layer2_outputs(1279) <= b;
    layer2_outputs(1280) <= not a or b;
    layer2_outputs(1281) <= a;
    layer2_outputs(1282) <= not b;
    layer2_outputs(1283) <= b and not a;
    layer2_outputs(1284) <= a and not b;
    layer2_outputs(1285) <= not b;
    layer2_outputs(1286) <= b and not a;
    layer2_outputs(1287) <= a and b;
    layer2_outputs(1288) <= not (a or b);
    layer2_outputs(1289) <= a;
    layer2_outputs(1290) <= not a;
    layer2_outputs(1291) <= a and b;
    layer2_outputs(1292) <= a xor b;
    layer2_outputs(1293) <= b;
    layer2_outputs(1294) <= b;
    layer2_outputs(1295) <= not (a or b);
    layer2_outputs(1296) <= a and b;
    layer2_outputs(1297) <= b and not a;
    layer2_outputs(1298) <= not a;
    layer2_outputs(1299) <= b;
    layer2_outputs(1300) <= a and b;
    layer2_outputs(1301) <= not (a and b);
    layer2_outputs(1302) <= a and not b;
    layer2_outputs(1303) <= not (a or b);
    layer2_outputs(1304) <= b and not a;
    layer2_outputs(1305) <= a;
    layer2_outputs(1306) <= a;
    layer2_outputs(1307) <= a xor b;
    layer2_outputs(1308) <= not (a and b);
    layer2_outputs(1309) <= a and b;
    layer2_outputs(1310) <= not a;
    layer2_outputs(1311) <= a and b;
    layer2_outputs(1312) <= not a;
    layer2_outputs(1313) <= a or b;
    layer2_outputs(1314) <= not (a and b);
    layer2_outputs(1315) <= not a;
    layer2_outputs(1316) <= a or b;
    layer2_outputs(1317) <= not b;
    layer2_outputs(1318) <= a or b;
    layer2_outputs(1319) <= not a or b;
    layer2_outputs(1320) <= b;
    layer2_outputs(1321) <= a xor b;
    layer2_outputs(1322) <= b;
    layer2_outputs(1323) <= not (a and b);
    layer2_outputs(1324) <= 1'b0;
    layer2_outputs(1325) <= not (a or b);
    layer2_outputs(1326) <= not (a and b);
    layer2_outputs(1327) <= not (a and b);
    layer2_outputs(1328) <= a and not b;
    layer2_outputs(1329) <= b and not a;
    layer2_outputs(1330) <= a and b;
    layer2_outputs(1331) <= not (a xor b);
    layer2_outputs(1332) <= not b;
    layer2_outputs(1333) <= a;
    layer2_outputs(1334) <= a and not b;
    layer2_outputs(1335) <= not b or a;
    layer2_outputs(1336) <= a and not b;
    layer2_outputs(1337) <= not b;
    layer2_outputs(1338) <= not a;
    layer2_outputs(1339) <= b and not a;
    layer2_outputs(1340) <= not (a and b);
    layer2_outputs(1341) <= a xor b;
    layer2_outputs(1342) <= not b;
    layer2_outputs(1343) <= not a;
    layer2_outputs(1344) <= not (a and b);
    layer2_outputs(1345) <= not b;
    layer2_outputs(1346) <= a;
    layer2_outputs(1347) <= a or b;
    layer2_outputs(1348) <= a;
    layer2_outputs(1349) <= not (a and b);
    layer2_outputs(1350) <= not (a or b);
    layer2_outputs(1351) <= not a;
    layer2_outputs(1352) <= a and not b;
    layer2_outputs(1353) <= a and b;
    layer2_outputs(1354) <= not a;
    layer2_outputs(1355) <= a;
    layer2_outputs(1356) <= b;
    layer2_outputs(1357) <= a or b;
    layer2_outputs(1358) <= a;
    layer2_outputs(1359) <= not (a or b);
    layer2_outputs(1360) <= not b;
    layer2_outputs(1361) <= a and b;
    layer2_outputs(1362) <= not a;
    layer2_outputs(1363) <= not (a or b);
    layer2_outputs(1364) <= not (a or b);
    layer2_outputs(1365) <= a;
    layer2_outputs(1366) <= not b or a;
    layer2_outputs(1367) <= b;
    layer2_outputs(1368) <= a or b;
    layer2_outputs(1369) <= not (a and b);
    layer2_outputs(1370) <= not a or b;
    layer2_outputs(1371) <= 1'b0;
    layer2_outputs(1372) <= not a;
    layer2_outputs(1373) <= 1'b0;
    layer2_outputs(1374) <= a and not b;
    layer2_outputs(1375) <= 1'b0;
    layer2_outputs(1376) <= not (a or b);
    layer2_outputs(1377) <= a or b;
    layer2_outputs(1378) <= b;
    layer2_outputs(1379) <= not a;
    layer2_outputs(1380) <= 1'b1;
    layer2_outputs(1381) <= b and not a;
    layer2_outputs(1382) <= a;
    layer2_outputs(1383) <= not b;
    layer2_outputs(1384) <= b;
    layer2_outputs(1385) <= not b or a;
    layer2_outputs(1386) <= not (a or b);
    layer2_outputs(1387) <= b;
    layer2_outputs(1388) <= b;
    layer2_outputs(1389) <= b;
    layer2_outputs(1390) <= not (a or b);
    layer2_outputs(1391) <= a and b;
    layer2_outputs(1392) <= not a;
    layer2_outputs(1393) <= 1'b1;
    layer2_outputs(1394) <= 1'b0;
    layer2_outputs(1395) <= a xor b;
    layer2_outputs(1396) <= not b;
    layer2_outputs(1397) <= b;
    layer2_outputs(1398) <= not a;
    layer2_outputs(1399) <= b and not a;
    layer2_outputs(1400) <= a and b;
    layer2_outputs(1401) <= not (a or b);
    layer2_outputs(1402) <= a and not b;
    layer2_outputs(1403) <= not a;
    layer2_outputs(1404) <= not (a or b);
    layer2_outputs(1405) <= not a or b;
    layer2_outputs(1406) <= not (a or b);
    layer2_outputs(1407) <= not b or a;
    layer2_outputs(1408) <= not a;
    layer2_outputs(1409) <= a and not b;
    layer2_outputs(1410) <= not (a xor b);
    layer2_outputs(1411) <= not b;
    layer2_outputs(1412) <= a and not b;
    layer2_outputs(1413) <= b;
    layer2_outputs(1414) <= not (a or b);
    layer2_outputs(1415) <= not a;
    layer2_outputs(1416) <= not b;
    layer2_outputs(1417) <= a;
    layer2_outputs(1418) <= not b;
    layer2_outputs(1419) <= a and not b;
    layer2_outputs(1420) <= not b;
    layer2_outputs(1421) <= not a;
    layer2_outputs(1422) <= a;
    layer2_outputs(1423) <= not a or b;
    layer2_outputs(1424) <= a or b;
    layer2_outputs(1425) <= a or b;
    layer2_outputs(1426) <= not (a and b);
    layer2_outputs(1427) <= a;
    layer2_outputs(1428) <= not a or b;
    layer2_outputs(1429) <= a;
    layer2_outputs(1430) <= not (a and b);
    layer2_outputs(1431) <= not b or a;
    layer2_outputs(1432) <= not b;
    layer2_outputs(1433) <= a and not b;
    layer2_outputs(1434) <= b and not a;
    layer2_outputs(1435) <= not b or a;
    layer2_outputs(1436) <= a and not b;
    layer2_outputs(1437) <= a and not b;
    layer2_outputs(1438) <= not (a xor b);
    layer2_outputs(1439) <= a and not b;
    layer2_outputs(1440) <= b and not a;
    layer2_outputs(1441) <= a and b;
    layer2_outputs(1442) <= b;
    layer2_outputs(1443) <= not b or a;
    layer2_outputs(1444) <= 1'b1;
    layer2_outputs(1445) <= a and not b;
    layer2_outputs(1446) <= a or b;
    layer2_outputs(1447) <= not b;
    layer2_outputs(1448) <= a and not b;
    layer2_outputs(1449) <= a and not b;
    layer2_outputs(1450) <= a;
    layer2_outputs(1451) <= a;
    layer2_outputs(1452) <= a;
    layer2_outputs(1453) <= b;
    layer2_outputs(1454) <= not (a xor b);
    layer2_outputs(1455) <= not b;
    layer2_outputs(1456) <= a xor b;
    layer2_outputs(1457) <= a and b;
    layer2_outputs(1458) <= a and b;
    layer2_outputs(1459) <= a and not b;
    layer2_outputs(1460) <= a and b;
    layer2_outputs(1461) <= not (a and b);
    layer2_outputs(1462) <= b;
    layer2_outputs(1463) <= not a or b;
    layer2_outputs(1464) <= not (a and b);
    layer2_outputs(1465) <= b;
    layer2_outputs(1466) <= not a;
    layer2_outputs(1467) <= a;
    layer2_outputs(1468) <= a;
    layer2_outputs(1469) <= b and not a;
    layer2_outputs(1470) <= not (a xor b);
    layer2_outputs(1471) <= not a or b;
    layer2_outputs(1472) <= not b;
    layer2_outputs(1473) <= a;
    layer2_outputs(1474) <= a or b;
    layer2_outputs(1475) <= a xor b;
    layer2_outputs(1476) <= a;
    layer2_outputs(1477) <= not a;
    layer2_outputs(1478) <= not a or b;
    layer2_outputs(1479) <= a;
    layer2_outputs(1480) <= not b;
    layer2_outputs(1481) <= not b or a;
    layer2_outputs(1482) <= not (a and b);
    layer2_outputs(1483) <= not a;
    layer2_outputs(1484) <= a or b;
    layer2_outputs(1485) <= a;
    layer2_outputs(1486) <= a and b;
    layer2_outputs(1487) <= not b;
    layer2_outputs(1488) <= not (a or b);
    layer2_outputs(1489) <= a;
    layer2_outputs(1490) <= not a;
    layer2_outputs(1491) <= a or b;
    layer2_outputs(1492) <= a and not b;
    layer2_outputs(1493) <= not b or a;
    layer2_outputs(1494) <= not b;
    layer2_outputs(1495) <= a and b;
    layer2_outputs(1496) <= a and b;
    layer2_outputs(1497) <= not (a and b);
    layer2_outputs(1498) <= a;
    layer2_outputs(1499) <= 1'b1;
    layer2_outputs(1500) <= not a;
    layer2_outputs(1501) <= not (a xor b);
    layer2_outputs(1502) <= not a;
    layer2_outputs(1503) <= a and b;
    layer2_outputs(1504) <= not a;
    layer2_outputs(1505) <= 1'b0;
    layer2_outputs(1506) <= not b or a;
    layer2_outputs(1507) <= a;
    layer2_outputs(1508) <= 1'b0;
    layer2_outputs(1509) <= a and b;
    layer2_outputs(1510) <= a;
    layer2_outputs(1511) <= not (a or b);
    layer2_outputs(1512) <= a;
    layer2_outputs(1513) <= a;
    layer2_outputs(1514) <= 1'b0;
    layer2_outputs(1515) <= a xor b;
    layer2_outputs(1516) <= not b;
    layer2_outputs(1517) <= 1'b1;
    layer2_outputs(1518) <= b and not a;
    layer2_outputs(1519) <= not a;
    layer2_outputs(1520) <= not a;
    layer2_outputs(1521) <= 1'b1;
    layer2_outputs(1522) <= not (a and b);
    layer2_outputs(1523) <= b;
    layer2_outputs(1524) <= a;
    layer2_outputs(1525) <= b;
    layer2_outputs(1526) <= a;
    layer2_outputs(1527) <= not (a or b);
    layer2_outputs(1528) <= not (a and b);
    layer2_outputs(1529) <= b and not a;
    layer2_outputs(1530) <= not (a or b);
    layer2_outputs(1531) <= b and not a;
    layer2_outputs(1532) <= not a;
    layer2_outputs(1533) <= 1'b0;
    layer2_outputs(1534) <= not a or b;
    layer2_outputs(1535) <= a;
    layer2_outputs(1536) <= not (a and b);
    layer2_outputs(1537) <= 1'b1;
    layer2_outputs(1538) <= b and not a;
    layer2_outputs(1539) <= a and b;
    layer2_outputs(1540) <= not (a or b);
    layer2_outputs(1541) <= not b;
    layer2_outputs(1542) <= b;
    layer2_outputs(1543) <= 1'b0;
    layer2_outputs(1544) <= a and b;
    layer2_outputs(1545) <= not a;
    layer2_outputs(1546) <= a and b;
    layer2_outputs(1547) <= not a;
    layer2_outputs(1548) <= not b;
    layer2_outputs(1549) <= not (a and b);
    layer2_outputs(1550) <= a or b;
    layer2_outputs(1551) <= b;
    layer2_outputs(1552) <= a and not b;
    layer2_outputs(1553) <= a xor b;
    layer2_outputs(1554) <= not b or a;
    layer2_outputs(1555) <= not a;
    layer2_outputs(1556) <= not (a and b);
    layer2_outputs(1557) <= not (a and b);
    layer2_outputs(1558) <= a and not b;
    layer2_outputs(1559) <= b;
    layer2_outputs(1560) <= not b;
    layer2_outputs(1561) <= a and b;
    layer2_outputs(1562) <= not a;
    layer2_outputs(1563) <= not b;
    layer2_outputs(1564) <= not b or a;
    layer2_outputs(1565) <= 1'b0;
    layer2_outputs(1566) <= not a;
    layer2_outputs(1567) <= not a;
    layer2_outputs(1568) <= b;
    layer2_outputs(1569) <= a xor b;
    layer2_outputs(1570) <= b;
    layer2_outputs(1571) <= not (a and b);
    layer2_outputs(1572) <= a and b;
    layer2_outputs(1573) <= 1'b1;
    layer2_outputs(1574) <= not a;
    layer2_outputs(1575) <= not (a xor b);
    layer2_outputs(1576) <= not a or b;
    layer2_outputs(1577) <= a xor b;
    layer2_outputs(1578) <= not (a and b);
    layer2_outputs(1579) <= not a;
    layer2_outputs(1580) <= 1'b0;
    layer2_outputs(1581) <= not (a and b);
    layer2_outputs(1582) <= b;
    layer2_outputs(1583) <= a xor b;
    layer2_outputs(1584) <= not (a xor b);
    layer2_outputs(1585) <= a or b;
    layer2_outputs(1586) <= not b;
    layer2_outputs(1587) <= a or b;
    layer2_outputs(1588) <= not (a or b);
    layer2_outputs(1589) <= a;
    layer2_outputs(1590) <= a;
    layer2_outputs(1591) <= not (a and b);
    layer2_outputs(1592) <= a and b;
    layer2_outputs(1593) <= not b;
    layer2_outputs(1594) <= b;
    layer2_outputs(1595) <= not (a or b);
    layer2_outputs(1596) <= not b;
    layer2_outputs(1597) <= a or b;
    layer2_outputs(1598) <= not b;
    layer2_outputs(1599) <= not (a and b);
    layer2_outputs(1600) <= not (a or b);
    layer2_outputs(1601) <= not a;
    layer2_outputs(1602) <= a and not b;
    layer2_outputs(1603) <= b;
    layer2_outputs(1604) <= not b;
    layer2_outputs(1605) <= a and not b;
    layer2_outputs(1606) <= b and not a;
    layer2_outputs(1607) <= a and b;
    layer2_outputs(1608) <= not b;
    layer2_outputs(1609) <= not b;
    layer2_outputs(1610) <= a;
    layer2_outputs(1611) <= 1'b0;
    layer2_outputs(1612) <= a and not b;
    layer2_outputs(1613) <= not a;
    layer2_outputs(1614) <= a and b;
    layer2_outputs(1615) <= a;
    layer2_outputs(1616) <= not b or a;
    layer2_outputs(1617) <= a or b;
    layer2_outputs(1618) <= a or b;
    layer2_outputs(1619) <= a and b;
    layer2_outputs(1620) <= not b;
    layer2_outputs(1621) <= 1'b0;
    layer2_outputs(1622) <= a and b;
    layer2_outputs(1623) <= not a;
    layer2_outputs(1624) <= not b or a;
    layer2_outputs(1625) <= 1'b0;
    layer2_outputs(1626) <= not a;
    layer2_outputs(1627) <= b and not a;
    layer2_outputs(1628) <= b;
    layer2_outputs(1629) <= not a;
    layer2_outputs(1630) <= a;
    layer2_outputs(1631) <= not a;
    layer2_outputs(1632) <= not a;
    layer2_outputs(1633) <= not (a and b);
    layer2_outputs(1634) <= a or b;
    layer2_outputs(1635) <= a;
    layer2_outputs(1636) <= a;
    layer2_outputs(1637) <= a and b;
    layer2_outputs(1638) <= a and b;
    layer2_outputs(1639) <= not (a xor b);
    layer2_outputs(1640) <= a and not b;
    layer2_outputs(1641) <= not b;
    layer2_outputs(1642) <= 1'b1;
    layer2_outputs(1643) <= b and not a;
    layer2_outputs(1644) <= b and not a;
    layer2_outputs(1645) <= a and not b;
    layer2_outputs(1646) <= a or b;
    layer2_outputs(1647) <= not b or a;
    layer2_outputs(1648) <= not (a or b);
    layer2_outputs(1649) <= a;
    layer2_outputs(1650) <= a and not b;
    layer2_outputs(1651) <= not (a or b);
    layer2_outputs(1652) <= not a or b;
    layer2_outputs(1653) <= a xor b;
    layer2_outputs(1654) <= not b or a;
    layer2_outputs(1655) <= not (a or b);
    layer2_outputs(1656) <= not (a and b);
    layer2_outputs(1657) <= a and b;
    layer2_outputs(1658) <= not (a or b);
    layer2_outputs(1659) <= not (a or b);
    layer2_outputs(1660) <= not a or b;
    layer2_outputs(1661) <= a;
    layer2_outputs(1662) <= b and not a;
    layer2_outputs(1663) <= a or b;
    layer2_outputs(1664) <= not (a or b);
    layer2_outputs(1665) <= b and not a;
    layer2_outputs(1666) <= a;
    layer2_outputs(1667) <= not a or b;
    layer2_outputs(1668) <= a or b;
    layer2_outputs(1669) <= not b;
    layer2_outputs(1670) <= not a or b;
    layer2_outputs(1671) <= a and b;
    layer2_outputs(1672) <= 1'b1;
    layer2_outputs(1673) <= not b;
    layer2_outputs(1674) <= 1'b1;
    layer2_outputs(1675) <= not (a and b);
    layer2_outputs(1676) <= not (a or b);
    layer2_outputs(1677) <= b and not a;
    layer2_outputs(1678) <= a or b;
    layer2_outputs(1679) <= not (a and b);
    layer2_outputs(1680) <= not b or a;
    layer2_outputs(1681) <= not b;
    layer2_outputs(1682) <= a and b;
    layer2_outputs(1683) <= not a;
    layer2_outputs(1684) <= 1'b0;
    layer2_outputs(1685) <= not (a and b);
    layer2_outputs(1686) <= a;
    layer2_outputs(1687) <= not b or a;
    layer2_outputs(1688) <= b and not a;
    layer2_outputs(1689) <= 1'b1;
    layer2_outputs(1690) <= not a;
    layer2_outputs(1691) <= 1'b0;
    layer2_outputs(1692) <= b and not a;
    layer2_outputs(1693) <= not a;
    layer2_outputs(1694) <= not b;
    layer2_outputs(1695) <= a or b;
    layer2_outputs(1696) <= a and not b;
    layer2_outputs(1697) <= not (a or b);
    layer2_outputs(1698) <= b and not a;
    layer2_outputs(1699) <= not (a and b);
    layer2_outputs(1700) <= 1'b1;
    layer2_outputs(1701) <= not b;
    layer2_outputs(1702) <= b;
    layer2_outputs(1703) <= not a or b;
    layer2_outputs(1704) <= not a or b;
    layer2_outputs(1705) <= a;
    layer2_outputs(1706) <= b;
    layer2_outputs(1707) <= a and not b;
    layer2_outputs(1708) <= not b or a;
    layer2_outputs(1709) <= not b;
    layer2_outputs(1710) <= b;
    layer2_outputs(1711) <= not a;
    layer2_outputs(1712) <= a or b;
    layer2_outputs(1713) <= not (a or b);
    layer2_outputs(1714) <= not b;
    layer2_outputs(1715) <= not b;
    layer2_outputs(1716) <= not a;
    layer2_outputs(1717) <= not (a and b);
    layer2_outputs(1718) <= not a;
    layer2_outputs(1719) <= b;
    layer2_outputs(1720) <= a or b;
    layer2_outputs(1721) <= b;
    layer2_outputs(1722) <= not b or a;
    layer2_outputs(1723) <= not a;
    layer2_outputs(1724) <= a and b;
    layer2_outputs(1725) <= not a;
    layer2_outputs(1726) <= b;
    layer2_outputs(1727) <= b and not a;
    layer2_outputs(1728) <= b and not a;
    layer2_outputs(1729) <= not a or b;
    layer2_outputs(1730) <= not b;
    layer2_outputs(1731) <= b and not a;
    layer2_outputs(1732) <= a;
    layer2_outputs(1733) <= not (a and b);
    layer2_outputs(1734) <= a or b;
    layer2_outputs(1735) <= not (a or b);
    layer2_outputs(1736) <= not a;
    layer2_outputs(1737) <= 1'b1;
    layer2_outputs(1738) <= a;
    layer2_outputs(1739) <= b;
    layer2_outputs(1740) <= a;
    layer2_outputs(1741) <= a and b;
    layer2_outputs(1742) <= not (a and b);
    layer2_outputs(1743) <= not b or a;
    layer2_outputs(1744) <= not b;
    layer2_outputs(1745) <= a and not b;
    layer2_outputs(1746) <= b and not a;
    layer2_outputs(1747) <= a and not b;
    layer2_outputs(1748) <= a and b;
    layer2_outputs(1749) <= a and b;
    layer2_outputs(1750) <= a and b;
    layer2_outputs(1751) <= not a or b;
    layer2_outputs(1752) <= b;
    layer2_outputs(1753) <= not b;
    layer2_outputs(1754) <= not (a xor b);
    layer2_outputs(1755) <= not b or a;
    layer2_outputs(1756) <= not a or b;
    layer2_outputs(1757) <= not (a and b);
    layer2_outputs(1758) <= not b;
    layer2_outputs(1759) <= not a;
    layer2_outputs(1760) <= not a or b;
    layer2_outputs(1761) <= a and not b;
    layer2_outputs(1762) <= not (a and b);
    layer2_outputs(1763) <= a;
    layer2_outputs(1764) <= a or b;
    layer2_outputs(1765) <= not b;
    layer2_outputs(1766) <= a and not b;
    layer2_outputs(1767) <= not (a and b);
    layer2_outputs(1768) <= not b or a;
    layer2_outputs(1769) <= not (a and b);
    layer2_outputs(1770) <= not b or a;
    layer2_outputs(1771) <= b;
    layer2_outputs(1772) <= not b or a;
    layer2_outputs(1773) <= not b;
    layer2_outputs(1774) <= b and not a;
    layer2_outputs(1775) <= a or b;
    layer2_outputs(1776) <= not a or b;
    layer2_outputs(1777) <= a xor b;
    layer2_outputs(1778) <= 1'b0;
    layer2_outputs(1779) <= b and not a;
    layer2_outputs(1780) <= b;
    layer2_outputs(1781) <= not (a and b);
    layer2_outputs(1782) <= not a;
    layer2_outputs(1783) <= b and not a;
    layer2_outputs(1784) <= a;
    layer2_outputs(1785) <= not a;
    layer2_outputs(1786) <= a or b;
    layer2_outputs(1787) <= a;
    layer2_outputs(1788) <= not (a and b);
    layer2_outputs(1789) <= not b or a;
    layer2_outputs(1790) <= a;
    layer2_outputs(1791) <= b;
    layer2_outputs(1792) <= not a or b;
    layer2_outputs(1793) <= not a or b;
    layer2_outputs(1794) <= not b or a;
    layer2_outputs(1795) <= not a or b;
    layer2_outputs(1796) <= 1'b0;
    layer2_outputs(1797) <= a;
    layer2_outputs(1798) <= not (a and b);
    layer2_outputs(1799) <= a;
    layer2_outputs(1800) <= not b;
    layer2_outputs(1801) <= a;
    layer2_outputs(1802) <= not a;
    layer2_outputs(1803) <= a xor b;
    layer2_outputs(1804) <= b;
    layer2_outputs(1805) <= a and b;
    layer2_outputs(1806) <= b and not a;
    layer2_outputs(1807) <= not a;
    layer2_outputs(1808) <= b;
    layer2_outputs(1809) <= b and not a;
    layer2_outputs(1810) <= not a or b;
    layer2_outputs(1811) <= b and not a;
    layer2_outputs(1812) <= not (a or b);
    layer2_outputs(1813) <= not b;
    layer2_outputs(1814) <= not (a and b);
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= not a or b;
    layer2_outputs(1817) <= a or b;
    layer2_outputs(1818) <= a and b;
    layer2_outputs(1819) <= b;
    layer2_outputs(1820) <= b;
    layer2_outputs(1821) <= not b or a;
    layer2_outputs(1822) <= a;
    layer2_outputs(1823) <= not (a or b);
    layer2_outputs(1824) <= not a;
    layer2_outputs(1825) <= not a or b;
    layer2_outputs(1826) <= not a or b;
    layer2_outputs(1827) <= not a;
    layer2_outputs(1828) <= not (a and b);
    layer2_outputs(1829) <= b and not a;
    layer2_outputs(1830) <= a and b;
    layer2_outputs(1831) <= b;
    layer2_outputs(1832) <= a;
    layer2_outputs(1833) <= not b;
    layer2_outputs(1834) <= not b;
    layer2_outputs(1835) <= b;
    layer2_outputs(1836) <= b and not a;
    layer2_outputs(1837) <= a;
    layer2_outputs(1838) <= not a or b;
    layer2_outputs(1839) <= a or b;
    layer2_outputs(1840) <= a or b;
    layer2_outputs(1841) <= a;
    layer2_outputs(1842) <= a and b;
    layer2_outputs(1843) <= a and not b;
    layer2_outputs(1844) <= not (a or b);
    layer2_outputs(1845) <= a;
    layer2_outputs(1846) <= not a or b;
    layer2_outputs(1847) <= not (a and b);
    layer2_outputs(1848) <= not (a and b);
    layer2_outputs(1849) <= not a;
    layer2_outputs(1850) <= b;
    layer2_outputs(1851) <= b;
    layer2_outputs(1852) <= not (a or b);
    layer2_outputs(1853) <= not a or b;
    layer2_outputs(1854) <= a or b;
    layer2_outputs(1855) <= 1'b0;
    layer2_outputs(1856) <= a and b;
    layer2_outputs(1857) <= b;
    layer2_outputs(1858) <= a;
    layer2_outputs(1859) <= not (a or b);
    layer2_outputs(1860) <= not b or a;
    layer2_outputs(1861) <= not (a and b);
    layer2_outputs(1862) <= a;
    layer2_outputs(1863) <= a or b;
    layer2_outputs(1864) <= not (a or b);
    layer2_outputs(1865) <= a or b;
    layer2_outputs(1866) <= not (a or b);
    layer2_outputs(1867) <= b;
    layer2_outputs(1868) <= a xor b;
    layer2_outputs(1869) <= b;
    layer2_outputs(1870) <= a or b;
    layer2_outputs(1871) <= b;
    layer2_outputs(1872) <= not (a xor b);
    layer2_outputs(1873) <= not a;
    layer2_outputs(1874) <= a and b;
    layer2_outputs(1875) <= not (a xor b);
    layer2_outputs(1876) <= b;
    layer2_outputs(1877) <= not b or a;
    layer2_outputs(1878) <= a;
    layer2_outputs(1879) <= not (a and b);
    layer2_outputs(1880) <= not (a xor b);
    layer2_outputs(1881) <= a;
    layer2_outputs(1882) <= not b;
    layer2_outputs(1883) <= not (a or b);
    layer2_outputs(1884) <= not (a or b);
    layer2_outputs(1885) <= a and not b;
    layer2_outputs(1886) <= not a;
    layer2_outputs(1887) <= a and b;
    layer2_outputs(1888) <= a;
    layer2_outputs(1889) <= not a or b;
    layer2_outputs(1890) <= not a or b;
    layer2_outputs(1891) <= a and b;
    layer2_outputs(1892) <= a and not b;
    layer2_outputs(1893) <= a and b;
    layer2_outputs(1894) <= 1'b0;
    layer2_outputs(1895) <= b and not a;
    layer2_outputs(1896) <= b;
    layer2_outputs(1897) <= not a;
    layer2_outputs(1898) <= b;
    layer2_outputs(1899) <= not b;
    layer2_outputs(1900) <= 1'b0;
    layer2_outputs(1901) <= not b or a;
    layer2_outputs(1902) <= a xor b;
    layer2_outputs(1903) <= a xor b;
    layer2_outputs(1904) <= a and b;
    layer2_outputs(1905) <= not (a and b);
    layer2_outputs(1906) <= b;
    layer2_outputs(1907) <= not (a xor b);
    layer2_outputs(1908) <= not a;
    layer2_outputs(1909) <= not a;
    layer2_outputs(1910) <= 1'b0;
    layer2_outputs(1911) <= a and not b;
    layer2_outputs(1912) <= b;
    layer2_outputs(1913) <= b and not a;
    layer2_outputs(1914) <= not (a xor b);
    layer2_outputs(1915) <= not (a or b);
    layer2_outputs(1916) <= not b;
    layer2_outputs(1917) <= not b or a;
    layer2_outputs(1918) <= a and b;
    layer2_outputs(1919) <= b;
    layer2_outputs(1920) <= b and not a;
    layer2_outputs(1921) <= a and b;
    layer2_outputs(1922) <= a and not b;
    layer2_outputs(1923) <= b and not a;
    layer2_outputs(1924) <= b;
    layer2_outputs(1925) <= b;
    layer2_outputs(1926) <= not a or b;
    layer2_outputs(1927) <= b and not a;
    layer2_outputs(1928) <= b;
    layer2_outputs(1929) <= a or b;
    layer2_outputs(1930) <= b;
    layer2_outputs(1931) <= not a or b;
    layer2_outputs(1932) <= b and not a;
    layer2_outputs(1933) <= not b;
    layer2_outputs(1934) <= not (a or b);
    layer2_outputs(1935) <= not b or a;
    layer2_outputs(1936) <= a and b;
    layer2_outputs(1937) <= not a or b;
    layer2_outputs(1938) <= a and b;
    layer2_outputs(1939) <= a and b;
    layer2_outputs(1940) <= not b;
    layer2_outputs(1941) <= a and not b;
    layer2_outputs(1942) <= not b;
    layer2_outputs(1943) <= b;
    layer2_outputs(1944) <= not (a or b);
    layer2_outputs(1945) <= not b or a;
    layer2_outputs(1946) <= not b or a;
    layer2_outputs(1947) <= not a;
    layer2_outputs(1948) <= a;
    layer2_outputs(1949) <= not a or b;
    layer2_outputs(1950) <= not b;
    layer2_outputs(1951) <= not a;
    layer2_outputs(1952) <= a;
    layer2_outputs(1953) <= not (a and b);
    layer2_outputs(1954) <= a;
    layer2_outputs(1955) <= not a or b;
    layer2_outputs(1956) <= a;
    layer2_outputs(1957) <= not (a or b);
    layer2_outputs(1958) <= not b or a;
    layer2_outputs(1959) <= not (a and b);
    layer2_outputs(1960) <= not a;
    layer2_outputs(1961) <= not (a and b);
    layer2_outputs(1962) <= a and not b;
    layer2_outputs(1963) <= b and not a;
    layer2_outputs(1964) <= not b;
    layer2_outputs(1965) <= a and b;
    layer2_outputs(1966) <= a;
    layer2_outputs(1967) <= not b;
    layer2_outputs(1968) <= not b or a;
    layer2_outputs(1969) <= 1'b0;
    layer2_outputs(1970) <= not a;
    layer2_outputs(1971) <= a;
    layer2_outputs(1972) <= b and not a;
    layer2_outputs(1973) <= not (a or b);
    layer2_outputs(1974) <= not b or a;
    layer2_outputs(1975) <= b;
    layer2_outputs(1976) <= a and b;
    layer2_outputs(1977) <= b and not a;
    layer2_outputs(1978) <= not a or b;
    layer2_outputs(1979) <= not b or a;
    layer2_outputs(1980) <= not b or a;
    layer2_outputs(1981) <= b;
    layer2_outputs(1982) <= 1'b1;
    layer2_outputs(1983) <= not (a or b);
    layer2_outputs(1984) <= not b;
    layer2_outputs(1985) <= not a;
    layer2_outputs(1986) <= not a;
    layer2_outputs(1987) <= a xor b;
    layer2_outputs(1988) <= not b;
    layer2_outputs(1989) <= not b;
    layer2_outputs(1990) <= 1'b1;
    layer2_outputs(1991) <= a or b;
    layer2_outputs(1992) <= b;
    layer2_outputs(1993) <= not a;
    layer2_outputs(1994) <= not b or a;
    layer2_outputs(1995) <= 1'b0;
    layer2_outputs(1996) <= a xor b;
    layer2_outputs(1997) <= b and not a;
    layer2_outputs(1998) <= a and b;
    layer2_outputs(1999) <= a and not b;
    layer2_outputs(2000) <= not a;
    layer2_outputs(2001) <= not (a or b);
    layer2_outputs(2002) <= not b;
    layer2_outputs(2003) <= 1'b1;
    layer2_outputs(2004) <= not (a or b);
    layer2_outputs(2005) <= not (a and b);
    layer2_outputs(2006) <= not b or a;
    layer2_outputs(2007) <= not a or b;
    layer2_outputs(2008) <= a or b;
    layer2_outputs(2009) <= not a;
    layer2_outputs(2010) <= not a;
    layer2_outputs(2011) <= a and b;
    layer2_outputs(2012) <= not b or a;
    layer2_outputs(2013) <= b and not a;
    layer2_outputs(2014) <= a;
    layer2_outputs(2015) <= a or b;
    layer2_outputs(2016) <= not b;
    layer2_outputs(2017) <= not b;
    layer2_outputs(2018) <= not a;
    layer2_outputs(2019) <= 1'b0;
    layer2_outputs(2020) <= not b;
    layer2_outputs(2021) <= a or b;
    layer2_outputs(2022) <= not (a and b);
    layer2_outputs(2023) <= not b;
    layer2_outputs(2024) <= a or b;
    layer2_outputs(2025) <= a;
    layer2_outputs(2026) <= not b or a;
    layer2_outputs(2027) <= a;
    layer2_outputs(2028) <= b;
    layer2_outputs(2029) <= not (a xor b);
    layer2_outputs(2030) <= 1'b0;
    layer2_outputs(2031) <= not a or b;
    layer2_outputs(2032) <= not b;
    layer2_outputs(2033) <= a and not b;
    layer2_outputs(2034) <= a xor b;
    layer2_outputs(2035) <= 1'b1;
    layer2_outputs(2036) <= a and not b;
    layer2_outputs(2037) <= a;
    layer2_outputs(2038) <= a or b;
    layer2_outputs(2039) <= not (a and b);
    layer2_outputs(2040) <= a;
    layer2_outputs(2041) <= not a or b;
    layer2_outputs(2042) <= a and not b;
    layer2_outputs(2043) <= not a or b;
    layer2_outputs(2044) <= not b or a;
    layer2_outputs(2045) <= a;
    layer2_outputs(2046) <= not a;
    layer2_outputs(2047) <= a and not b;
    layer2_outputs(2048) <= not a;
    layer2_outputs(2049) <= a and not b;
    layer2_outputs(2050) <= not a;
    layer2_outputs(2051) <= not b;
    layer2_outputs(2052) <= not a or b;
    layer2_outputs(2053) <= not a or b;
    layer2_outputs(2054) <= not a;
    layer2_outputs(2055) <= a;
    layer2_outputs(2056) <= 1'b0;
    layer2_outputs(2057) <= not (a or b);
    layer2_outputs(2058) <= not b or a;
    layer2_outputs(2059) <= not a;
    layer2_outputs(2060) <= not (a or b);
    layer2_outputs(2061) <= b and not a;
    layer2_outputs(2062) <= b;
    layer2_outputs(2063) <= a or b;
    layer2_outputs(2064) <= not b;
    layer2_outputs(2065) <= 1'b1;
    layer2_outputs(2066) <= not (a and b);
    layer2_outputs(2067) <= a xor b;
    layer2_outputs(2068) <= 1'b0;
    layer2_outputs(2069) <= a;
    layer2_outputs(2070) <= a and not b;
    layer2_outputs(2071) <= a xor b;
    layer2_outputs(2072) <= not a;
    layer2_outputs(2073) <= a;
    layer2_outputs(2074) <= a or b;
    layer2_outputs(2075) <= a;
    layer2_outputs(2076) <= not (a or b);
    layer2_outputs(2077) <= a xor b;
    layer2_outputs(2078) <= a and b;
    layer2_outputs(2079) <= a xor b;
    layer2_outputs(2080) <= a;
    layer2_outputs(2081) <= not b;
    layer2_outputs(2082) <= not a or b;
    layer2_outputs(2083) <= a xor b;
    layer2_outputs(2084) <= a and b;
    layer2_outputs(2085) <= a;
    layer2_outputs(2086) <= not (a or b);
    layer2_outputs(2087) <= a xor b;
    layer2_outputs(2088) <= not a;
    layer2_outputs(2089) <= not (a or b);
    layer2_outputs(2090) <= a;
    layer2_outputs(2091) <= a and b;
    layer2_outputs(2092) <= a;
    layer2_outputs(2093) <= not (a and b);
    layer2_outputs(2094) <= b;
    layer2_outputs(2095) <= not a;
    layer2_outputs(2096) <= not (a or b);
    layer2_outputs(2097) <= 1'b0;
    layer2_outputs(2098) <= not (a and b);
    layer2_outputs(2099) <= not a or b;
    layer2_outputs(2100) <= a;
    layer2_outputs(2101) <= not (a or b);
    layer2_outputs(2102) <= a and not b;
    layer2_outputs(2103) <= a and b;
    layer2_outputs(2104) <= b and not a;
    layer2_outputs(2105) <= b;
    layer2_outputs(2106) <= a;
    layer2_outputs(2107) <= a;
    layer2_outputs(2108) <= b and not a;
    layer2_outputs(2109) <= not a or b;
    layer2_outputs(2110) <= not (a and b);
    layer2_outputs(2111) <= not b;
    layer2_outputs(2112) <= b;
    layer2_outputs(2113) <= not (a and b);
    layer2_outputs(2114) <= not a;
    layer2_outputs(2115) <= a xor b;
    layer2_outputs(2116) <= not (a or b);
    layer2_outputs(2117) <= not a;
    layer2_outputs(2118) <= b;
    layer2_outputs(2119) <= not a;
    layer2_outputs(2120) <= 1'b1;
    layer2_outputs(2121) <= not a;
    layer2_outputs(2122) <= b and not a;
    layer2_outputs(2123) <= a;
    layer2_outputs(2124) <= b;
    layer2_outputs(2125) <= not a;
    layer2_outputs(2126) <= not a or b;
    layer2_outputs(2127) <= a;
    layer2_outputs(2128) <= not a;
    layer2_outputs(2129) <= a;
    layer2_outputs(2130) <= a or b;
    layer2_outputs(2131) <= not (a and b);
    layer2_outputs(2132) <= not b;
    layer2_outputs(2133) <= b;
    layer2_outputs(2134) <= a or b;
    layer2_outputs(2135) <= a and not b;
    layer2_outputs(2136) <= 1'b0;
    layer2_outputs(2137) <= not b or a;
    layer2_outputs(2138) <= a and b;
    layer2_outputs(2139) <= b;
    layer2_outputs(2140) <= not (a and b);
    layer2_outputs(2141) <= not b or a;
    layer2_outputs(2142) <= b;
    layer2_outputs(2143) <= not a;
    layer2_outputs(2144) <= a;
    layer2_outputs(2145) <= 1'b1;
    layer2_outputs(2146) <= a or b;
    layer2_outputs(2147) <= not a;
    layer2_outputs(2148) <= not a;
    layer2_outputs(2149) <= not b or a;
    layer2_outputs(2150) <= not b;
    layer2_outputs(2151) <= a;
    layer2_outputs(2152) <= a and not b;
    layer2_outputs(2153) <= not a or b;
    layer2_outputs(2154) <= not b;
    layer2_outputs(2155) <= not (a or b);
    layer2_outputs(2156) <= b and not a;
    layer2_outputs(2157) <= not b or a;
    layer2_outputs(2158) <= 1'b1;
    layer2_outputs(2159) <= not a or b;
    layer2_outputs(2160) <= a;
    layer2_outputs(2161) <= not a;
    layer2_outputs(2162) <= a or b;
    layer2_outputs(2163) <= not a or b;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= b and not a;
    layer2_outputs(2166) <= not a;
    layer2_outputs(2167) <= not (a or b);
    layer2_outputs(2168) <= not a;
    layer2_outputs(2169) <= not b;
    layer2_outputs(2170) <= b;
    layer2_outputs(2171) <= not (a xor b);
    layer2_outputs(2172) <= a and not b;
    layer2_outputs(2173) <= not b;
    layer2_outputs(2174) <= not (a or b);
    layer2_outputs(2175) <= 1'b1;
    layer2_outputs(2176) <= not a;
    layer2_outputs(2177) <= not b;
    layer2_outputs(2178) <= not b;
    layer2_outputs(2179) <= a;
    layer2_outputs(2180) <= a and b;
    layer2_outputs(2181) <= not a or b;
    layer2_outputs(2182) <= b;
    layer2_outputs(2183) <= 1'b1;
    layer2_outputs(2184) <= not a;
    layer2_outputs(2185) <= not (a or b);
    layer2_outputs(2186) <= not b or a;
    layer2_outputs(2187) <= a and not b;
    layer2_outputs(2188) <= a and not b;
    layer2_outputs(2189) <= a xor b;
    layer2_outputs(2190) <= a and not b;
    layer2_outputs(2191) <= not b;
    layer2_outputs(2192) <= 1'b1;
    layer2_outputs(2193) <= not a;
    layer2_outputs(2194) <= not a or b;
    layer2_outputs(2195) <= not (a or b);
    layer2_outputs(2196) <= not (a and b);
    layer2_outputs(2197) <= a and not b;
    layer2_outputs(2198) <= not (a xor b);
    layer2_outputs(2199) <= not b or a;
    layer2_outputs(2200) <= not (a or b);
    layer2_outputs(2201) <= a xor b;
    layer2_outputs(2202) <= not a or b;
    layer2_outputs(2203) <= not b;
    layer2_outputs(2204) <= a;
    layer2_outputs(2205) <= not (a and b);
    layer2_outputs(2206) <= a;
    layer2_outputs(2207) <= not b or a;
    layer2_outputs(2208) <= not b;
    layer2_outputs(2209) <= not (a or b);
    layer2_outputs(2210) <= a or b;
    layer2_outputs(2211) <= a and not b;
    layer2_outputs(2212) <= b;
    layer2_outputs(2213) <= not a or b;
    layer2_outputs(2214) <= a;
    layer2_outputs(2215) <= not b or a;
    layer2_outputs(2216) <= not a;
    layer2_outputs(2217) <= not (a and b);
    layer2_outputs(2218) <= not (a and b);
    layer2_outputs(2219) <= not a;
    layer2_outputs(2220) <= not b;
    layer2_outputs(2221) <= a or b;
    layer2_outputs(2222) <= a xor b;
    layer2_outputs(2223) <= not b or a;
    layer2_outputs(2224) <= a;
    layer2_outputs(2225) <= not (a and b);
    layer2_outputs(2226) <= a or b;
    layer2_outputs(2227) <= a;
    layer2_outputs(2228) <= not b;
    layer2_outputs(2229) <= not b or a;
    layer2_outputs(2230) <= a and not b;
    layer2_outputs(2231) <= not a;
    layer2_outputs(2232) <= not (a or b);
    layer2_outputs(2233) <= not a or b;
    layer2_outputs(2234) <= not a or b;
    layer2_outputs(2235) <= a and not b;
    layer2_outputs(2236) <= not b or a;
    layer2_outputs(2237) <= b and not a;
    layer2_outputs(2238) <= b;
    layer2_outputs(2239) <= b;
    layer2_outputs(2240) <= not (a and b);
    layer2_outputs(2241) <= a and b;
    layer2_outputs(2242) <= a;
    layer2_outputs(2243) <= not b or a;
    layer2_outputs(2244) <= not a or b;
    layer2_outputs(2245) <= a or b;
    layer2_outputs(2246) <= not b;
    layer2_outputs(2247) <= not b;
    layer2_outputs(2248) <= not a;
    layer2_outputs(2249) <= 1'b0;
    layer2_outputs(2250) <= a;
    layer2_outputs(2251) <= b;
    layer2_outputs(2252) <= not a;
    layer2_outputs(2253) <= b;
    layer2_outputs(2254) <= not a or b;
    layer2_outputs(2255) <= not (a xor b);
    layer2_outputs(2256) <= b and not a;
    layer2_outputs(2257) <= a and b;
    layer2_outputs(2258) <= a or b;
    layer2_outputs(2259) <= b;
    layer2_outputs(2260) <= a and b;
    layer2_outputs(2261) <= b;
    layer2_outputs(2262) <= not (a xor b);
    layer2_outputs(2263) <= not (a and b);
    layer2_outputs(2264) <= not (a or b);
    layer2_outputs(2265) <= not (a or b);
    layer2_outputs(2266) <= not (a or b);
    layer2_outputs(2267) <= a or b;
    layer2_outputs(2268) <= not (a or b);
    layer2_outputs(2269) <= a and b;
    layer2_outputs(2270) <= not (a and b);
    layer2_outputs(2271) <= b;
    layer2_outputs(2272) <= b;
    layer2_outputs(2273) <= not b or a;
    layer2_outputs(2274) <= not b;
    layer2_outputs(2275) <= b;
    layer2_outputs(2276) <= not b;
    layer2_outputs(2277) <= 1'b0;
    layer2_outputs(2278) <= a or b;
    layer2_outputs(2279) <= a xor b;
    layer2_outputs(2280) <= a or b;
    layer2_outputs(2281) <= a or b;
    layer2_outputs(2282) <= b;
    layer2_outputs(2283) <= not b;
    layer2_outputs(2284) <= not (a and b);
    layer2_outputs(2285) <= not a;
    layer2_outputs(2286) <= a;
    layer2_outputs(2287) <= b and not a;
    layer2_outputs(2288) <= not b;
    layer2_outputs(2289) <= not a;
    layer2_outputs(2290) <= b;
    layer2_outputs(2291) <= not b or a;
    layer2_outputs(2292) <= a and not b;
    layer2_outputs(2293) <= a or b;
    layer2_outputs(2294) <= not b or a;
    layer2_outputs(2295) <= 1'b1;
    layer2_outputs(2296) <= a and b;
    layer2_outputs(2297) <= not (a and b);
    layer2_outputs(2298) <= a;
    layer2_outputs(2299) <= not (a or b);
    layer2_outputs(2300) <= a or b;
    layer2_outputs(2301) <= 1'b0;
    layer2_outputs(2302) <= a;
    layer2_outputs(2303) <= not b;
    layer2_outputs(2304) <= not (a or b);
    layer2_outputs(2305) <= not a;
    layer2_outputs(2306) <= 1'b1;
    layer2_outputs(2307) <= a and b;
    layer2_outputs(2308) <= not (a xor b);
    layer2_outputs(2309) <= not b or a;
    layer2_outputs(2310) <= not a;
    layer2_outputs(2311) <= not (a and b);
    layer2_outputs(2312) <= not (a and b);
    layer2_outputs(2313) <= not (a and b);
    layer2_outputs(2314) <= not a;
    layer2_outputs(2315) <= not (a or b);
    layer2_outputs(2316) <= a;
    layer2_outputs(2317) <= b and not a;
    layer2_outputs(2318) <= not a;
    layer2_outputs(2319) <= a;
    layer2_outputs(2320) <= not (a and b);
    layer2_outputs(2321) <= 1'b0;
    layer2_outputs(2322) <= 1'b1;
    layer2_outputs(2323) <= not (a or b);
    layer2_outputs(2324) <= a or b;
    layer2_outputs(2325) <= b and not a;
    layer2_outputs(2326) <= not a;
    layer2_outputs(2327) <= not b;
    layer2_outputs(2328) <= not a;
    layer2_outputs(2329) <= not a;
    layer2_outputs(2330) <= a and b;
    layer2_outputs(2331) <= not b;
    layer2_outputs(2332) <= a xor b;
    layer2_outputs(2333) <= not a;
    layer2_outputs(2334) <= not (a or b);
    layer2_outputs(2335) <= not a;
    layer2_outputs(2336) <= not a;
    layer2_outputs(2337) <= b and not a;
    layer2_outputs(2338) <= a and b;
    layer2_outputs(2339) <= a and not b;
    layer2_outputs(2340) <= b and not a;
    layer2_outputs(2341) <= 1'b0;
    layer2_outputs(2342) <= a and b;
    layer2_outputs(2343) <= a and b;
    layer2_outputs(2344) <= a and b;
    layer2_outputs(2345) <= a;
    layer2_outputs(2346) <= b;
    layer2_outputs(2347) <= not b or a;
    layer2_outputs(2348) <= b;
    layer2_outputs(2349) <= a;
    layer2_outputs(2350) <= a;
    layer2_outputs(2351) <= not b or a;
    layer2_outputs(2352) <= not (a xor b);
    layer2_outputs(2353) <= a;
    layer2_outputs(2354) <= not (a and b);
    layer2_outputs(2355) <= a and b;
    layer2_outputs(2356) <= not b or a;
    layer2_outputs(2357) <= a and b;
    layer2_outputs(2358) <= a or b;
    layer2_outputs(2359) <= not b;
    layer2_outputs(2360) <= a and b;
    layer2_outputs(2361) <= not b;
    layer2_outputs(2362) <= b and not a;
    layer2_outputs(2363) <= not b;
    layer2_outputs(2364) <= b;
    layer2_outputs(2365) <= not b or a;
    layer2_outputs(2366) <= not b;
    layer2_outputs(2367) <= not a;
    layer2_outputs(2368) <= a and b;
    layer2_outputs(2369) <= a;
    layer2_outputs(2370) <= a or b;
    layer2_outputs(2371) <= a xor b;
    layer2_outputs(2372) <= b and not a;
    layer2_outputs(2373) <= b;
    layer2_outputs(2374) <= a;
    layer2_outputs(2375) <= not b;
    layer2_outputs(2376) <= not a or b;
    layer2_outputs(2377) <= not a or b;
    layer2_outputs(2378) <= a;
    layer2_outputs(2379) <= b;
    layer2_outputs(2380) <= a;
    layer2_outputs(2381) <= a or b;
    layer2_outputs(2382) <= a and not b;
    layer2_outputs(2383) <= not b or a;
    layer2_outputs(2384) <= not a;
    layer2_outputs(2385) <= b and not a;
    layer2_outputs(2386) <= a or b;
    layer2_outputs(2387) <= not b;
    layer2_outputs(2388) <= a or b;
    layer2_outputs(2389) <= not a or b;
    layer2_outputs(2390) <= not (a and b);
    layer2_outputs(2391) <= a or b;
    layer2_outputs(2392) <= not a;
    layer2_outputs(2393) <= not (a xor b);
    layer2_outputs(2394) <= not a or b;
    layer2_outputs(2395) <= a and b;
    layer2_outputs(2396) <= not (a and b);
    layer2_outputs(2397) <= not (a and b);
    layer2_outputs(2398) <= a and b;
    layer2_outputs(2399) <= b and not a;
    layer2_outputs(2400) <= a;
    layer2_outputs(2401) <= a and b;
    layer2_outputs(2402) <= 1'b0;
    layer2_outputs(2403) <= not a or b;
    layer2_outputs(2404) <= not b or a;
    layer2_outputs(2405) <= a and b;
    layer2_outputs(2406) <= not (a and b);
    layer2_outputs(2407) <= 1'b1;
    layer2_outputs(2408) <= 1'b1;
    layer2_outputs(2409) <= a or b;
    layer2_outputs(2410) <= not (a and b);
    layer2_outputs(2411) <= a and b;
    layer2_outputs(2412) <= a and not b;
    layer2_outputs(2413) <= a and b;
    layer2_outputs(2414) <= not b;
    layer2_outputs(2415) <= b and not a;
    layer2_outputs(2416) <= a and not b;
    layer2_outputs(2417) <= not a or b;
    layer2_outputs(2418) <= a and b;
    layer2_outputs(2419) <= a xor b;
    layer2_outputs(2420) <= not a;
    layer2_outputs(2421) <= a or b;
    layer2_outputs(2422) <= not (a xor b);
    layer2_outputs(2423) <= a or b;
    layer2_outputs(2424) <= not (a and b);
    layer2_outputs(2425) <= not a or b;
    layer2_outputs(2426) <= a and b;
    layer2_outputs(2427) <= not (a xor b);
    layer2_outputs(2428) <= b;
    layer2_outputs(2429) <= a;
    layer2_outputs(2430) <= not a;
    layer2_outputs(2431) <= not (a and b);
    layer2_outputs(2432) <= b;
    layer2_outputs(2433) <= a and not b;
    layer2_outputs(2434) <= a;
    layer2_outputs(2435) <= not b or a;
    layer2_outputs(2436) <= not (a or b);
    layer2_outputs(2437) <= b and not a;
    layer2_outputs(2438) <= not (a or b);
    layer2_outputs(2439) <= not (a and b);
    layer2_outputs(2440) <= not b;
    layer2_outputs(2441) <= not a;
    layer2_outputs(2442) <= not b;
    layer2_outputs(2443) <= a or b;
    layer2_outputs(2444) <= not a or b;
    layer2_outputs(2445) <= not b;
    layer2_outputs(2446) <= a and not b;
    layer2_outputs(2447) <= not b;
    layer2_outputs(2448) <= not (a and b);
    layer2_outputs(2449) <= b;
    layer2_outputs(2450) <= not a;
    layer2_outputs(2451) <= 1'b0;
    layer2_outputs(2452) <= not b or a;
    layer2_outputs(2453) <= not b;
    layer2_outputs(2454) <= a and not b;
    layer2_outputs(2455) <= not b;
    layer2_outputs(2456) <= not a or b;
    layer2_outputs(2457) <= not b or a;
    layer2_outputs(2458) <= not (a xor b);
    layer2_outputs(2459) <= b;
    layer2_outputs(2460) <= not b or a;
    layer2_outputs(2461) <= not b;
    layer2_outputs(2462) <= not (a or b);
    layer2_outputs(2463) <= a;
    layer2_outputs(2464) <= not b;
    layer2_outputs(2465) <= not b;
    layer2_outputs(2466) <= a and b;
    layer2_outputs(2467) <= not b;
    layer2_outputs(2468) <= a;
    layer2_outputs(2469) <= not b or a;
    layer2_outputs(2470) <= a or b;
    layer2_outputs(2471) <= a and b;
    layer2_outputs(2472) <= not a;
    layer2_outputs(2473) <= not a or b;
    layer2_outputs(2474) <= a;
    layer2_outputs(2475) <= not b;
    layer2_outputs(2476) <= b;
    layer2_outputs(2477) <= a;
    layer2_outputs(2478) <= a or b;
    layer2_outputs(2479) <= a or b;
    layer2_outputs(2480) <= a;
    layer2_outputs(2481) <= a and b;
    layer2_outputs(2482) <= a;
    layer2_outputs(2483) <= not (a and b);
    layer2_outputs(2484) <= a;
    layer2_outputs(2485) <= not b;
    layer2_outputs(2486) <= b;
    layer2_outputs(2487) <= not a or b;
    layer2_outputs(2488) <= not (a or b);
    layer2_outputs(2489) <= not (a xor b);
    layer2_outputs(2490) <= not b or a;
    layer2_outputs(2491) <= not a;
    layer2_outputs(2492) <= 1'b1;
    layer2_outputs(2493) <= not a or b;
    layer2_outputs(2494) <= b;
    layer2_outputs(2495) <= a or b;
    layer2_outputs(2496) <= a and b;
    layer2_outputs(2497) <= not b or a;
    layer2_outputs(2498) <= not b;
    layer2_outputs(2499) <= not (a xor b);
    layer2_outputs(2500) <= 1'b1;
    layer2_outputs(2501) <= not a;
    layer2_outputs(2502) <= b;
    layer2_outputs(2503) <= b;
    layer2_outputs(2504) <= not a or b;
    layer2_outputs(2505) <= not a or b;
    layer2_outputs(2506) <= b;
    layer2_outputs(2507) <= b and not a;
    layer2_outputs(2508) <= not (a or b);
    layer2_outputs(2509) <= a or b;
    layer2_outputs(2510) <= a and not b;
    layer2_outputs(2511) <= a or b;
    layer2_outputs(2512) <= not b or a;
    layer2_outputs(2513) <= b and not a;
    layer2_outputs(2514) <= not (a or b);
    layer2_outputs(2515) <= not b;
    layer2_outputs(2516) <= not (a xor b);
    layer2_outputs(2517) <= not a;
    layer2_outputs(2518) <= not (a and b);
    layer2_outputs(2519) <= b and not a;
    layer2_outputs(2520) <= b and not a;
    layer2_outputs(2521) <= b and not a;
    layer2_outputs(2522) <= not (a and b);
    layer2_outputs(2523) <= not a;
    layer2_outputs(2524) <= not a;
    layer2_outputs(2525) <= not b;
    layer2_outputs(2526) <= a and not b;
    layer2_outputs(2527) <= a and not b;
    layer2_outputs(2528) <= a and not b;
    layer2_outputs(2529) <= not b;
    layer2_outputs(2530) <= not (a xor b);
    layer2_outputs(2531) <= not (a and b);
    layer2_outputs(2532) <= not a;
    layer2_outputs(2533) <= a and b;
    layer2_outputs(2534) <= not b;
    layer2_outputs(2535) <= a and b;
    layer2_outputs(2536) <= a and b;
    layer2_outputs(2537) <= a or b;
    layer2_outputs(2538) <= not a or b;
    layer2_outputs(2539) <= not (a or b);
    layer2_outputs(2540) <= b and not a;
    layer2_outputs(2541) <= a;
    layer2_outputs(2542) <= 1'b1;
    layer2_outputs(2543) <= a;
    layer2_outputs(2544) <= a and b;
    layer2_outputs(2545) <= not (a xor b);
    layer2_outputs(2546) <= not b or a;
    layer2_outputs(2547) <= not b;
    layer2_outputs(2548) <= not b;
    layer2_outputs(2549) <= 1'b0;
    layer2_outputs(2550) <= a xor b;
    layer2_outputs(2551) <= not (a or b);
    layer2_outputs(2552) <= b and not a;
    layer2_outputs(2553) <= not a or b;
    layer2_outputs(2554) <= not (a or b);
    layer2_outputs(2555) <= not a;
    layer2_outputs(2556) <= not a or b;
    layer2_outputs(2557) <= a and b;
    layer2_outputs(2558) <= not b;
    layer2_outputs(2559) <= b;
    layer3_outputs(0) <= not b or a;
    layer3_outputs(1) <= a;
    layer3_outputs(2) <= a xor b;
    layer3_outputs(3) <= b and not a;
    layer3_outputs(4) <= b;
    layer3_outputs(5) <= not b;
    layer3_outputs(6) <= a and b;
    layer3_outputs(7) <= not b or a;
    layer3_outputs(8) <= not (a or b);
    layer3_outputs(9) <= b and not a;
    layer3_outputs(10) <= not a or b;
    layer3_outputs(11) <= b and not a;
    layer3_outputs(12) <= b and not a;
    layer3_outputs(13) <= not a;
    layer3_outputs(14) <= not a;
    layer3_outputs(15) <= not a;
    layer3_outputs(16) <= a;
    layer3_outputs(17) <= a or b;
    layer3_outputs(18) <= a and b;
    layer3_outputs(19) <= b;
    layer3_outputs(20) <= not b;
    layer3_outputs(21) <= not b;
    layer3_outputs(22) <= not a;
    layer3_outputs(23) <= not (a or b);
    layer3_outputs(24) <= b;
    layer3_outputs(25) <= b;
    layer3_outputs(26) <= not a or b;
    layer3_outputs(27) <= a or b;
    layer3_outputs(28) <= not (a and b);
    layer3_outputs(29) <= a;
    layer3_outputs(30) <= b;
    layer3_outputs(31) <= a and b;
    layer3_outputs(32) <= not (a and b);
    layer3_outputs(33) <= not (a or b);
    layer3_outputs(34) <= b;
    layer3_outputs(35) <= b;
    layer3_outputs(36) <= b and not a;
    layer3_outputs(37) <= not b;
    layer3_outputs(38) <= a;
    layer3_outputs(39) <= not (a and b);
    layer3_outputs(40) <= not a;
    layer3_outputs(41) <= not (a or b);
    layer3_outputs(42) <= a;
    layer3_outputs(43) <= a and b;
    layer3_outputs(44) <= b and not a;
    layer3_outputs(45) <= b;
    layer3_outputs(46) <= b;
    layer3_outputs(47) <= b;
    layer3_outputs(48) <= b;
    layer3_outputs(49) <= not b;
    layer3_outputs(50) <= not a or b;
    layer3_outputs(51) <= not b;
    layer3_outputs(52) <= not a or b;
    layer3_outputs(53) <= a;
    layer3_outputs(54) <= a;
    layer3_outputs(55) <= a;
    layer3_outputs(56) <= not a;
    layer3_outputs(57) <= b;
    layer3_outputs(58) <= not a;
    layer3_outputs(59) <= a and not b;
    layer3_outputs(60) <= b;
    layer3_outputs(61) <= a and not b;
    layer3_outputs(62) <= a and not b;
    layer3_outputs(63) <= not b;
    layer3_outputs(64) <= b and not a;
    layer3_outputs(65) <= not a or b;
    layer3_outputs(66) <= a and not b;
    layer3_outputs(67) <= a or b;
    layer3_outputs(68) <= not a;
    layer3_outputs(69) <= not a;
    layer3_outputs(70) <= 1'b0;
    layer3_outputs(71) <= not b or a;
    layer3_outputs(72) <= b and not a;
    layer3_outputs(73) <= b;
    layer3_outputs(74) <= a and not b;
    layer3_outputs(75) <= b;
    layer3_outputs(76) <= a;
    layer3_outputs(77) <= a;
    layer3_outputs(78) <= a;
    layer3_outputs(79) <= a;
    layer3_outputs(80) <= b and not a;
    layer3_outputs(81) <= a or b;
    layer3_outputs(82) <= not b or a;
    layer3_outputs(83) <= not a or b;
    layer3_outputs(84) <= not b;
    layer3_outputs(85) <= not a or b;
    layer3_outputs(86) <= not (a and b);
    layer3_outputs(87) <= b;
    layer3_outputs(88) <= not b;
    layer3_outputs(89) <= not (a or b);
    layer3_outputs(90) <= b;
    layer3_outputs(91) <= b and not a;
    layer3_outputs(92) <= b;
    layer3_outputs(93) <= a and not b;
    layer3_outputs(94) <= a;
    layer3_outputs(95) <= not (a or b);
    layer3_outputs(96) <= not a;
    layer3_outputs(97) <= not b or a;
    layer3_outputs(98) <= a;
    layer3_outputs(99) <= not b or a;
    layer3_outputs(100) <= not b or a;
    layer3_outputs(101) <= a;
    layer3_outputs(102) <= not (a and b);
    layer3_outputs(103) <= not (a and b);
    layer3_outputs(104) <= not b or a;
    layer3_outputs(105) <= a or b;
    layer3_outputs(106) <= not a or b;
    layer3_outputs(107) <= not (a and b);
    layer3_outputs(108) <= b and not a;
    layer3_outputs(109) <= b;
    layer3_outputs(110) <= not b;
    layer3_outputs(111) <= b and not a;
    layer3_outputs(112) <= a;
    layer3_outputs(113) <= b;
    layer3_outputs(114) <= 1'b0;
    layer3_outputs(115) <= a and b;
    layer3_outputs(116) <= a or b;
    layer3_outputs(117) <= not a;
    layer3_outputs(118) <= not b;
    layer3_outputs(119) <= a and not b;
    layer3_outputs(120) <= a or b;
    layer3_outputs(121) <= a;
    layer3_outputs(122) <= not b;
    layer3_outputs(123) <= not b or a;
    layer3_outputs(124) <= b and not a;
    layer3_outputs(125) <= b;
    layer3_outputs(126) <= not a or b;
    layer3_outputs(127) <= not a;
    layer3_outputs(128) <= not a or b;
    layer3_outputs(129) <= 1'b1;
    layer3_outputs(130) <= not a;
    layer3_outputs(131) <= b;
    layer3_outputs(132) <= a and not b;
    layer3_outputs(133) <= a;
    layer3_outputs(134) <= not a;
    layer3_outputs(135) <= not b;
    layer3_outputs(136) <= b;
    layer3_outputs(137) <= not (a or b);
    layer3_outputs(138) <= b;
    layer3_outputs(139) <= a and not b;
    layer3_outputs(140) <= a or b;
    layer3_outputs(141) <= 1'b1;
    layer3_outputs(142) <= b and not a;
    layer3_outputs(143) <= not (a or b);
    layer3_outputs(144) <= 1'b0;
    layer3_outputs(145) <= a;
    layer3_outputs(146) <= not (a and b);
    layer3_outputs(147) <= not b;
    layer3_outputs(148) <= not (a and b);
    layer3_outputs(149) <= a and b;
    layer3_outputs(150) <= not (a or b);
    layer3_outputs(151) <= not (a or b);
    layer3_outputs(152) <= b and not a;
    layer3_outputs(153) <= not (a and b);
    layer3_outputs(154) <= 1'b0;
    layer3_outputs(155) <= a;
    layer3_outputs(156) <= a;
    layer3_outputs(157) <= not a;
    layer3_outputs(158) <= not a;
    layer3_outputs(159) <= b;
    layer3_outputs(160) <= not b;
    layer3_outputs(161) <= 1'b0;
    layer3_outputs(162) <= not b;
    layer3_outputs(163) <= not a;
    layer3_outputs(164) <= a and not b;
    layer3_outputs(165) <= not (a and b);
    layer3_outputs(166) <= not b;
    layer3_outputs(167) <= 1'b1;
    layer3_outputs(168) <= not b;
    layer3_outputs(169) <= not a;
    layer3_outputs(170) <= not (a or b);
    layer3_outputs(171) <= not b;
    layer3_outputs(172) <= b;
    layer3_outputs(173) <= a;
    layer3_outputs(174) <= 1'b0;
    layer3_outputs(175) <= 1'b0;
    layer3_outputs(176) <= a and b;
    layer3_outputs(177) <= a;
    layer3_outputs(178) <= b;
    layer3_outputs(179) <= not (a or b);
    layer3_outputs(180) <= not (a or b);
    layer3_outputs(181) <= b and not a;
    layer3_outputs(182) <= a and b;
    layer3_outputs(183) <= a;
    layer3_outputs(184) <= not b;
    layer3_outputs(185) <= not (a and b);
    layer3_outputs(186) <= b and not a;
    layer3_outputs(187) <= a or b;
    layer3_outputs(188) <= not a or b;
    layer3_outputs(189) <= a and b;
    layer3_outputs(190) <= a;
    layer3_outputs(191) <= a;
    layer3_outputs(192) <= not b or a;
    layer3_outputs(193) <= a and not b;
    layer3_outputs(194) <= 1'b1;
    layer3_outputs(195) <= not (a and b);
    layer3_outputs(196) <= b and not a;
    layer3_outputs(197) <= a xor b;
    layer3_outputs(198) <= b;
    layer3_outputs(199) <= a;
    layer3_outputs(200) <= not (a or b);
    layer3_outputs(201) <= not a or b;
    layer3_outputs(202) <= a and b;
    layer3_outputs(203) <= not (a and b);
    layer3_outputs(204) <= not (a xor b);
    layer3_outputs(205) <= a or b;
    layer3_outputs(206) <= a and b;
    layer3_outputs(207) <= a or b;
    layer3_outputs(208) <= a;
    layer3_outputs(209) <= not (a or b);
    layer3_outputs(210) <= 1'b0;
    layer3_outputs(211) <= not b;
    layer3_outputs(212) <= b and not a;
    layer3_outputs(213) <= b;
    layer3_outputs(214) <= not (a and b);
    layer3_outputs(215) <= not b or a;
    layer3_outputs(216) <= a or b;
    layer3_outputs(217) <= b;
    layer3_outputs(218) <= b and not a;
    layer3_outputs(219) <= not a;
    layer3_outputs(220) <= a and b;
    layer3_outputs(221) <= not (a and b);
    layer3_outputs(222) <= not a;
    layer3_outputs(223) <= not a;
    layer3_outputs(224) <= not (a or b);
    layer3_outputs(225) <= not (a or b);
    layer3_outputs(226) <= not a or b;
    layer3_outputs(227) <= a or b;
    layer3_outputs(228) <= b and not a;
    layer3_outputs(229) <= not (a or b);
    layer3_outputs(230) <= a;
    layer3_outputs(231) <= not a or b;
    layer3_outputs(232) <= b;
    layer3_outputs(233) <= 1'b1;
    layer3_outputs(234) <= not a;
    layer3_outputs(235) <= not b;
    layer3_outputs(236) <= not a;
    layer3_outputs(237) <= a or b;
    layer3_outputs(238) <= b;
    layer3_outputs(239) <= not b;
    layer3_outputs(240) <= not a;
    layer3_outputs(241) <= a and not b;
    layer3_outputs(242) <= a and not b;
    layer3_outputs(243) <= a;
    layer3_outputs(244) <= not a or b;
    layer3_outputs(245) <= not (a xor b);
    layer3_outputs(246) <= b and not a;
    layer3_outputs(247) <= not (a xor b);
    layer3_outputs(248) <= b and not a;
    layer3_outputs(249) <= a and b;
    layer3_outputs(250) <= not (a and b);
    layer3_outputs(251) <= a or b;
    layer3_outputs(252) <= not b;
    layer3_outputs(253) <= not b;
    layer3_outputs(254) <= a;
    layer3_outputs(255) <= a or b;
    layer3_outputs(256) <= a and not b;
    layer3_outputs(257) <= not (a and b);
    layer3_outputs(258) <= a and b;
    layer3_outputs(259) <= a or b;
    layer3_outputs(260) <= not a;
    layer3_outputs(261) <= 1'b0;
    layer3_outputs(262) <= not b;
    layer3_outputs(263) <= a;
    layer3_outputs(264) <= not (a and b);
    layer3_outputs(265) <= not (a and b);
    layer3_outputs(266) <= a and b;
    layer3_outputs(267) <= b and not a;
    layer3_outputs(268) <= a;
    layer3_outputs(269) <= a;
    layer3_outputs(270) <= 1'b0;
    layer3_outputs(271) <= not (a or b);
    layer3_outputs(272) <= not (a and b);
    layer3_outputs(273) <= not a;
    layer3_outputs(274) <= not (a or b);
    layer3_outputs(275) <= not (a xor b);
    layer3_outputs(276) <= not b;
    layer3_outputs(277) <= a and not b;
    layer3_outputs(278) <= a and not b;
    layer3_outputs(279) <= not b;
    layer3_outputs(280) <= b and not a;
    layer3_outputs(281) <= not a;
    layer3_outputs(282) <= not a or b;
    layer3_outputs(283) <= a;
    layer3_outputs(284) <= a and b;
    layer3_outputs(285) <= not b or a;
    layer3_outputs(286) <= not a;
    layer3_outputs(287) <= not (a or b);
    layer3_outputs(288) <= a and not b;
    layer3_outputs(289) <= not (a xor b);
    layer3_outputs(290) <= a and not b;
    layer3_outputs(291) <= not b;
    layer3_outputs(292) <= a and not b;
    layer3_outputs(293) <= a;
    layer3_outputs(294) <= not a;
    layer3_outputs(295) <= not a or b;
    layer3_outputs(296) <= not a;
    layer3_outputs(297) <= b and not a;
    layer3_outputs(298) <= not (a and b);
    layer3_outputs(299) <= not a;
    layer3_outputs(300) <= not a;
    layer3_outputs(301) <= not (a and b);
    layer3_outputs(302) <= 1'b0;
    layer3_outputs(303) <= b and not a;
    layer3_outputs(304) <= a;
    layer3_outputs(305) <= not b;
    layer3_outputs(306) <= not a;
    layer3_outputs(307) <= a;
    layer3_outputs(308) <= not a;
    layer3_outputs(309) <= not (a or b);
    layer3_outputs(310) <= not a or b;
    layer3_outputs(311) <= not a;
    layer3_outputs(312) <= a;
    layer3_outputs(313) <= not a or b;
    layer3_outputs(314) <= b;
    layer3_outputs(315) <= a and b;
    layer3_outputs(316) <= b;
    layer3_outputs(317) <= not a;
    layer3_outputs(318) <= not a or b;
    layer3_outputs(319) <= b;
    layer3_outputs(320) <= not (a or b);
    layer3_outputs(321) <= not a;
    layer3_outputs(322) <= a and not b;
    layer3_outputs(323) <= not b or a;
    layer3_outputs(324) <= not (a and b);
    layer3_outputs(325) <= not b;
    layer3_outputs(326) <= a;
    layer3_outputs(327) <= not (a and b);
    layer3_outputs(328) <= not (a or b);
    layer3_outputs(329) <= b;
    layer3_outputs(330) <= b;
    layer3_outputs(331) <= not a;
    layer3_outputs(332) <= a;
    layer3_outputs(333) <= 1'b1;
    layer3_outputs(334) <= not b;
    layer3_outputs(335) <= a and b;
    layer3_outputs(336) <= 1'b0;
    layer3_outputs(337) <= a or b;
    layer3_outputs(338) <= not b;
    layer3_outputs(339) <= not b;
    layer3_outputs(340) <= not a or b;
    layer3_outputs(341) <= not (a and b);
    layer3_outputs(342) <= a;
    layer3_outputs(343) <= b and not a;
    layer3_outputs(344) <= not a;
    layer3_outputs(345) <= not b;
    layer3_outputs(346) <= a or b;
    layer3_outputs(347) <= not b;
    layer3_outputs(348) <= a or b;
    layer3_outputs(349) <= not a;
    layer3_outputs(350) <= not (a or b);
    layer3_outputs(351) <= not (a or b);
    layer3_outputs(352) <= a xor b;
    layer3_outputs(353) <= b;
    layer3_outputs(354) <= not (a xor b);
    layer3_outputs(355) <= b and not a;
    layer3_outputs(356) <= not b or a;
    layer3_outputs(357) <= not a or b;
    layer3_outputs(358) <= not b;
    layer3_outputs(359) <= 1'b1;
    layer3_outputs(360) <= b;
    layer3_outputs(361) <= a and not b;
    layer3_outputs(362) <= 1'b1;
    layer3_outputs(363) <= not a;
    layer3_outputs(364) <= not a;
    layer3_outputs(365) <= not (a and b);
    layer3_outputs(366) <= not a or b;
    layer3_outputs(367) <= not (a or b);
    layer3_outputs(368) <= a;
    layer3_outputs(369) <= not (a or b);
    layer3_outputs(370) <= not b;
    layer3_outputs(371) <= not a;
    layer3_outputs(372) <= b;
    layer3_outputs(373) <= not a;
    layer3_outputs(374) <= a;
    layer3_outputs(375) <= not (a xor b);
    layer3_outputs(376) <= not a;
    layer3_outputs(377) <= not a or b;
    layer3_outputs(378) <= not (a or b);
    layer3_outputs(379) <= not a;
    layer3_outputs(380) <= not (a and b);
    layer3_outputs(381) <= a and b;
    layer3_outputs(382) <= b;
    layer3_outputs(383) <= not a or b;
    layer3_outputs(384) <= a or b;
    layer3_outputs(385) <= not (a or b);
    layer3_outputs(386) <= not (a or b);
    layer3_outputs(387) <= not b or a;
    layer3_outputs(388) <= a;
    layer3_outputs(389) <= a;
    layer3_outputs(390) <= not b or a;
    layer3_outputs(391) <= not a or b;
    layer3_outputs(392) <= a or b;
    layer3_outputs(393) <= not (a xor b);
    layer3_outputs(394) <= not b;
    layer3_outputs(395) <= b;
    layer3_outputs(396) <= not b or a;
    layer3_outputs(397) <= a and b;
    layer3_outputs(398) <= not b or a;
    layer3_outputs(399) <= not b;
    layer3_outputs(400) <= 1'b1;
    layer3_outputs(401) <= b and not a;
    layer3_outputs(402) <= b and not a;
    layer3_outputs(403) <= b;
    layer3_outputs(404) <= a and b;
    layer3_outputs(405) <= a and not b;
    layer3_outputs(406) <= a or b;
    layer3_outputs(407) <= b and not a;
    layer3_outputs(408) <= not a or b;
    layer3_outputs(409) <= b and not a;
    layer3_outputs(410) <= b;
    layer3_outputs(411) <= not b;
    layer3_outputs(412) <= a or b;
    layer3_outputs(413) <= not (a and b);
    layer3_outputs(414) <= a;
    layer3_outputs(415) <= a and not b;
    layer3_outputs(416) <= not (a xor b);
    layer3_outputs(417) <= not b;
    layer3_outputs(418) <= b;
    layer3_outputs(419) <= a xor b;
    layer3_outputs(420) <= not b;
    layer3_outputs(421) <= not (a and b);
    layer3_outputs(422) <= a or b;
    layer3_outputs(423) <= a and not b;
    layer3_outputs(424) <= a or b;
    layer3_outputs(425) <= 1'b1;
    layer3_outputs(426) <= 1'b1;
    layer3_outputs(427) <= b and not a;
    layer3_outputs(428) <= not a;
    layer3_outputs(429) <= not b;
    layer3_outputs(430) <= a or b;
    layer3_outputs(431) <= b and not a;
    layer3_outputs(432) <= not (a and b);
    layer3_outputs(433) <= a and not b;
    layer3_outputs(434) <= not (a xor b);
    layer3_outputs(435) <= a and not b;
    layer3_outputs(436) <= not (a or b);
    layer3_outputs(437) <= not (a or b);
    layer3_outputs(438) <= not (a and b);
    layer3_outputs(439) <= b and not a;
    layer3_outputs(440) <= b;
    layer3_outputs(441) <= a and b;
    layer3_outputs(442) <= not b or a;
    layer3_outputs(443) <= not (a and b);
    layer3_outputs(444) <= not a;
    layer3_outputs(445) <= b;
    layer3_outputs(446) <= not b or a;
    layer3_outputs(447) <= b;
    layer3_outputs(448) <= not (a and b);
    layer3_outputs(449) <= not (a or b);
    layer3_outputs(450) <= not b or a;
    layer3_outputs(451) <= not a;
    layer3_outputs(452) <= 1'b1;
    layer3_outputs(453) <= not a;
    layer3_outputs(454) <= not b;
    layer3_outputs(455) <= not b;
    layer3_outputs(456) <= a xor b;
    layer3_outputs(457) <= b and not a;
    layer3_outputs(458) <= b;
    layer3_outputs(459) <= a;
    layer3_outputs(460) <= b and not a;
    layer3_outputs(461) <= b;
    layer3_outputs(462) <= not a;
    layer3_outputs(463) <= not b;
    layer3_outputs(464) <= not (a or b);
    layer3_outputs(465) <= a and not b;
    layer3_outputs(466) <= not (a or b);
    layer3_outputs(467) <= b;
    layer3_outputs(468) <= not a;
    layer3_outputs(469) <= not b;
    layer3_outputs(470) <= not a;
    layer3_outputs(471) <= not (a or b);
    layer3_outputs(472) <= b and not a;
    layer3_outputs(473) <= a or b;
    layer3_outputs(474) <= a;
    layer3_outputs(475) <= not a or b;
    layer3_outputs(476) <= a and not b;
    layer3_outputs(477) <= a;
    layer3_outputs(478) <= not b or a;
    layer3_outputs(479) <= not (a and b);
    layer3_outputs(480) <= b and not a;
    layer3_outputs(481) <= b;
    layer3_outputs(482) <= b and not a;
    layer3_outputs(483) <= not (a or b);
    layer3_outputs(484) <= not b;
    layer3_outputs(485) <= b;
    layer3_outputs(486) <= not b;
    layer3_outputs(487) <= a or b;
    layer3_outputs(488) <= not b;
    layer3_outputs(489) <= a or b;
    layer3_outputs(490) <= b;
    layer3_outputs(491) <= b;
    layer3_outputs(492) <= not a;
    layer3_outputs(493) <= not b or a;
    layer3_outputs(494) <= not a;
    layer3_outputs(495) <= not a;
    layer3_outputs(496) <= 1'b1;
    layer3_outputs(497) <= a;
    layer3_outputs(498) <= not a;
    layer3_outputs(499) <= not a or b;
    layer3_outputs(500) <= not a;
    layer3_outputs(501) <= not a;
    layer3_outputs(502) <= 1'b0;
    layer3_outputs(503) <= not a;
    layer3_outputs(504) <= b and not a;
    layer3_outputs(505) <= 1'b1;
    layer3_outputs(506) <= b;
    layer3_outputs(507) <= not b or a;
    layer3_outputs(508) <= not (a or b);
    layer3_outputs(509) <= not (a xor b);
    layer3_outputs(510) <= a or b;
    layer3_outputs(511) <= 1'b1;
    layer3_outputs(512) <= not a or b;
    layer3_outputs(513) <= not a or b;
    layer3_outputs(514) <= a;
    layer3_outputs(515) <= a and b;
    layer3_outputs(516) <= a;
    layer3_outputs(517) <= a and b;
    layer3_outputs(518) <= b and not a;
    layer3_outputs(519) <= 1'b1;
    layer3_outputs(520) <= not (a and b);
    layer3_outputs(521) <= 1'b1;
    layer3_outputs(522) <= a;
    layer3_outputs(523) <= 1'b0;
    layer3_outputs(524) <= a xor b;
    layer3_outputs(525) <= not b or a;
    layer3_outputs(526) <= not (a or b);
    layer3_outputs(527) <= a and not b;
    layer3_outputs(528) <= a or b;
    layer3_outputs(529) <= not a or b;
    layer3_outputs(530) <= not (a or b);
    layer3_outputs(531) <= b and not a;
    layer3_outputs(532) <= not (a or b);
    layer3_outputs(533) <= b;
    layer3_outputs(534) <= a and b;
    layer3_outputs(535) <= not b or a;
    layer3_outputs(536) <= not b or a;
    layer3_outputs(537) <= a xor b;
    layer3_outputs(538) <= not a or b;
    layer3_outputs(539) <= b and not a;
    layer3_outputs(540) <= a;
    layer3_outputs(541) <= a and b;
    layer3_outputs(542) <= a and not b;
    layer3_outputs(543) <= not (a or b);
    layer3_outputs(544) <= a;
    layer3_outputs(545) <= a and not b;
    layer3_outputs(546) <= not b or a;
    layer3_outputs(547) <= b and not a;
    layer3_outputs(548) <= a or b;
    layer3_outputs(549) <= not a;
    layer3_outputs(550) <= a and b;
    layer3_outputs(551) <= not (a or b);
    layer3_outputs(552) <= not (a or b);
    layer3_outputs(553) <= not (a and b);
    layer3_outputs(554) <= not b or a;
    layer3_outputs(555) <= b and not a;
    layer3_outputs(556) <= b and not a;
    layer3_outputs(557) <= a or b;
    layer3_outputs(558) <= a xor b;
    layer3_outputs(559) <= not (a and b);
    layer3_outputs(560) <= not a or b;
    layer3_outputs(561) <= not a or b;
    layer3_outputs(562) <= not (a or b);
    layer3_outputs(563) <= 1'b0;
    layer3_outputs(564) <= not b;
    layer3_outputs(565) <= not a or b;
    layer3_outputs(566) <= a;
    layer3_outputs(567) <= 1'b1;
    layer3_outputs(568) <= not b or a;
    layer3_outputs(569) <= not b or a;
    layer3_outputs(570) <= a or b;
    layer3_outputs(571) <= not (a or b);
    layer3_outputs(572) <= 1'b1;
    layer3_outputs(573) <= 1'b1;
    layer3_outputs(574) <= not (a and b);
    layer3_outputs(575) <= a and b;
    layer3_outputs(576) <= b;
    layer3_outputs(577) <= not b;
    layer3_outputs(578) <= b;
    layer3_outputs(579) <= a and not b;
    layer3_outputs(580) <= not a;
    layer3_outputs(581) <= 1'b1;
    layer3_outputs(582) <= not a;
    layer3_outputs(583) <= not a;
    layer3_outputs(584) <= not b or a;
    layer3_outputs(585) <= not a;
    layer3_outputs(586) <= b and not a;
    layer3_outputs(587) <= not a or b;
    layer3_outputs(588) <= not (a and b);
    layer3_outputs(589) <= not b or a;
    layer3_outputs(590) <= not b or a;
    layer3_outputs(591) <= b;
    layer3_outputs(592) <= not (a and b);
    layer3_outputs(593) <= a;
    layer3_outputs(594) <= not (a and b);
    layer3_outputs(595) <= a xor b;
    layer3_outputs(596) <= not b;
    layer3_outputs(597) <= 1'b0;
    layer3_outputs(598) <= not b or a;
    layer3_outputs(599) <= a and not b;
    layer3_outputs(600) <= not a;
    layer3_outputs(601) <= not b;
    layer3_outputs(602) <= not a;
    layer3_outputs(603) <= not (a or b);
    layer3_outputs(604) <= b;
    layer3_outputs(605) <= not b or a;
    layer3_outputs(606) <= b;
    layer3_outputs(607) <= 1'b0;
    layer3_outputs(608) <= 1'b0;
    layer3_outputs(609) <= not a;
    layer3_outputs(610) <= a and not b;
    layer3_outputs(611) <= a;
    layer3_outputs(612) <= 1'b1;
    layer3_outputs(613) <= a;
    layer3_outputs(614) <= not (a and b);
    layer3_outputs(615) <= a and b;
    layer3_outputs(616) <= not (a or b);
    layer3_outputs(617) <= not b;
    layer3_outputs(618) <= not a;
    layer3_outputs(619) <= not a;
    layer3_outputs(620) <= b;
    layer3_outputs(621) <= a and b;
    layer3_outputs(622) <= a and not b;
    layer3_outputs(623) <= a;
    layer3_outputs(624) <= not a;
    layer3_outputs(625) <= not b or a;
    layer3_outputs(626) <= not a or b;
    layer3_outputs(627) <= a and b;
    layer3_outputs(628) <= a or b;
    layer3_outputs(629) <= not b;
    layer3_outputs(630) <= not a;
    layer3_outputs(631) <= a;
    layer3_outputs(632) <= not (a xor b);
    layer3_outputs(633) <= 1'b1;
    layer3_outputs(634) <= b;
    layer3_outputs(635) <= not a or b;
    layer3_outputs(636) <= a and b;
    layer3_outputs(637) <= a and b;
    layer3_outputs(638) <= not a;
    layer3_outputs(639) <= not (a or b);
    layer3_outputs(640) <= not a;
    layer3_outputs(641) <= a or b;
    layer3_outputs(642) <= not b or a;
    layer3_outputs(643) <= b;
    layer3_outputs(644) <= a and not b;
    layer3_outputs(645) <= b;
    layer3_outputs(646) <= not a;
    layer3_outputs(647) <= a and not b;
    layer3_outputs(648) <= a;
    layer3_outputs(649) <= a and not b;
    layer3_outputs(650) <= not a;
    layer3_outputs(651) <= not (a or b);
    layer3_outputs(652) <= not a;
    layer3_outputs(653) <= not b or a;
    layer3_outputs(654) <= not b;
    layer3_outputs(655) <= not (a and b);
    layer3_outputs(656) <= b;
    layer3_outputs(657) <= 1'b0;
    layer3_outputs(658) <= not a;
    layer3_outputs(659) <= not a;
    layer3_outputs(660) <= b and not a;
    layer3_outputs(661) <= a and not b;
    layer3_outputs(662) <= b;
    layer3_outputs(663) <= a and b;
    layer3_outputs(664) <= a or b;
    layer3_outputs(665) <= 1'b1;
    layer3_outputs(666) <= a and b;
    layer3_outputs(667) <= 1'b1;
    layer3_outputs(668) <= a;
    layer3_outputs(669) <= not a;
    layer3_outputs(670) <= not (a and b);
    layer3_outputs(671) <= not b;
    layer3_outputs(672) <= a;
    layer3_outputs(673) <= a and b;
    layer3_outputs(674) <= not a;
    layer3_outputs(675) <= not (a and b);
    layer3_outputs(676) <= b;
    layer3_outputs(677) <= not b;
    layer3_outputs(678) <= not (a xor b);
    layer3_outputs(679) <= not b;
    layer3_outputs(680) <= not (a and b);
    layer3_outputs(681) <= not a;
    layer3_outputs(682) <= not b;
    layer3_outputs(683) <= a and not b;
    layer3_outputs(684) <= not a or b;
    layer3_outputs(685) <= b and not a;
    layer3_outputs(686) <= not a;
    layer3_outputs(687) <= 1'b0;
    layer3_outputs(688) <= a and b;
    layer3_outputs(689) <= b;
    layer3_outputs(690) <= b;
    layer3_outputs(691) <= b and not a;
    layer3_outputs(692) <= not (a and b);
    layer3_outputs(693) <= not a;
    layer3_outputs(694) <= a and b;
    layer3_outputs(695) <= not a or b;
    layer3_outputs(696) <= a xor b;
    layer3_outputs(697) <= a xor b;
    layer3_outputs(698) <= not b;
    layer3_outputs(699) <= a and b;
    layer3_outputs(700) <= b and not a;
    layer3_outputs(701) <= a and b;
    layer3_outputs(702) <= a and not b;
    layer3_outputs(703) <= b;
    layer3_outputs(704) <= a and not b;
    layer3_outputs(705) <= a xor b;
    layer3_outputs(706) <= not b;
    layer3_outputs(707) <= a and b;
    layer3_outputs(708) <= b and not a;
    layer3_outputs(709) <= a;
    layer3_outputs(710) <= not b;
    layer3_outputs(711) <= b and not a;
    layer3_outputs(712) <= a or b;
    layer3_outputs(713) <= not a or b;
    layer3_outputs(714) <= not b;
    layer3_outputs(715) <= a;
    layer3_outputs(716) <= a and b;
    layer3_outputs(717) <= not (a and b);
    layer3_outputs(718) <= a xor b;
    layer3_outputs(719) <= not b or a;
    layer3_outputs(720) <= not (a xor b);
    layer3_outputs(721) <= a or b;
    layer3_outputs(722) <= a xor b;
    layer3_outputs(723) <= b and not a;
    layer3_outputs(724) <= not a or b;
    layer3_outputs(725) <= not b or a;
    layer3_outputs(726) <= a xor b;
    layer3_outputs(727) <= not (a and b);
    layer3_outputs(728) <= a or b;
    layer3_outputs(729) <= a and b;
    layer3_outputs(730) <= a;
    layer3_outputs(731) <= not (a xor b);
    layer3_outputs(732) <= a;
    layer3_outputs(733) <= b and not a;
    layer3_outputs(734) <= not a or b;
    layer3_outputs(735) <= not b or a;
    layer3_outputs(736) <= not b or a;
    layer3_outputs(737) <= not a;
    layer3_outputs(738) <= not (a and b);
    layer3_outputs(739) <= a or b;
    layer3_outputs(740) <= b and not a;
    layer3_outputs(741) <= not b;
    layer3_outputs(742) <= not a;
    layer3_outputs(743) <= b;
    layer3_outputs(744) <= not a;
    layer3_outputs(745) <= not (a or b);
    layer3_outputs(746) <= not (a or b);
    layer3_outputs(747) <= not b;
    layer3_outputs(748) <= not (a xor b);
    layer3_outputs(749) <= a xor b;
    layer3_outputs(750) <= a xor b;
    layer3_outputs(751) <= not b;
    layer3_outputs(752) <= a or b;
    layer3_outputs(753) <= not a;
    layer3_outputs(754) <= b;
    layer3_outputs(755) <= a and not b;
    layer3_outputs(756) <= 1'b0;
    layer3_outputs(757) <= not b or a;
    layer3_outputs(758) <= not a or b;
    layer3_outputs(759) <= a or b;
    layer3_outputs(760) <= not (a and b);
    layer3_outputs(761) <= a and b;
    layer3_outputs(762) <= not b;
    layer3_outputs(763) <= b and not a;
    layer3_outputs(764) <= b;
    layer3_outputs(765) <= not a;
    layer3_outputs(766) <= b;
    layer3_outputs(767) <= not b or a;
    layer3_outputs(768) <= b and not a;
    layer3_outputs(769) <= a;
    layer3_outputs(770) <= a;
    layer3_outputs(771) <= b;
    layer3_outputs(772) <= a and not b;
    layer3_outputs(773) <= b;
    layer3_outputs(774) <= b;
    layer3_outputs(775) <= not a;
    layer3_outputs(776) <= 1'b1;
    layer3_outputs(777) <= a xor b;
    layer3_outputs(778) <= b and not a;
    layer3_outputs(779) <= not a;
    layer3_outputs(780) <= not (a and b);
    layer3_outputs(781) <= a and not b;
    layer3_outputs(782) <= a or b;
    layer3_outputs(783) <= b and not a;
    layer3_outputs(784) <= not b;
    layer3_outputs(785) <= a or b;
    layer3_outputs(786) <= 1'b1;
    layer3_outputs(787) <= not b;
    layer3_outputs(788) <= 1'b1;
    layer3_outputs(789) <= b and not a;
    layer3_outputs(790) <= a and b;
    layer3_outputs(791) <= b and not a;
    layer3_outputs(792) <= 1'b0;
    layer3_outputs(793) <= not (a or b);
    layer3_outputs(794) <= a;
    layer3_outputs(795) <= not (a and b);
    layer3_outputs(796) <= a and b;
    layer3_outputs(797) <= b and not a;
    layer3_outputs(798) <= not b;
    layer3_outputs(799) <= not a or b;
    layer3_outputs(800) <= not (a and b);
    layer3_outputs(801) <= a or b;
    layer3_outputs(802) <= a;
    layer3_outputs(803) <= b;
    layer3_outputs(804) <= not b or a;
    layer3_outputs(805) <= not b;
    layer3_outputs(806) <= a;
    layer3_outputs(807) <= b and not a;
    layer3_outputs(808) <= a or b;
    layer3_outputs(809) <= a and not b;
    layer3_outputs(810) <= not a;
    layer3_outputs(811) <= not a;
    layer3_outputs(812) <= a;
    layer3_outputs(813) <= 1'b1;
    layer3_outputs(814) <= not (a or b);
    layer3_outputs(815) <= a and not b;
    layer3_outputs(816) <= not b;
    layer3_outputs(817) <= a;
    layer3_outputs(818) <= not (a xor b);
    layer3_outputs(819) <= not b or a;
    layer3_outputs(820) <= a;
    layer3_outputs(821) <= b;
    layer3_outputs(822) <= a;
    layer3_outputs(823) <= 1'b1;
    layer3_outputs(824) <= not a or b;
    layer3_outputs(825) <= not b;
    layer3_outputs(826) <= a and b;
    layer3_outputs(827) <= a and b;
    layer3_outputs(828) <= a and b;
    layer3_outputs(829) <= not (a and b);
    layer3_outputs(830) <= b;
    layer3_outputs(831) <= not (a and b);
    layer3_outputs(832) <= not b or a;
    layer3_outputs(833) <= not a or b;
    layer3_outputs(834) <= a xor b;
    layer3_outputs(835) <= 1'b1;
    layer3_outputs(836) <= not b or a;
    layer3_outputs(837) <= not a;
    layer3_outputs(838) <= not b;
    layer3_outputs(839) <= not a or b;
    layer3_outputs(840) <= not b;
    layer3_outputs(841) <= not b or a;
    layer3_outputs(842) <= b;
    layer3_outputs(843) <= a or b;
    layer3_outputs(844) <= not a;
    layer3_outputs(845) <= a;
    layer3_outputs(846) <= not a;
    layer3_outputs(847) <= not (a and b);
    layer3_outputs(848) <= not (a and b);
    layer3_outputs(849) <= not b or a;
    layer3_outputs(850) <= b;
    layer3_outputs(851) <= not a;
    layer3_outputs(852) <= not a;
    layer3_outputs(853) <= not b or a;
    layer3_outputs(854) <= not a;
    layer3_outputs(855) <= not a;
    layer3_outputs(856) <= not b or a;
    layer3_outputs(857) <= not b;
    layer3_outputs(858) <= a xor b;
    layer3_outputs(859) <= a or b;
    layer3_outputs(860) <= a;
    layer3_outputs(861) <= a;
    layer3_outputs(862) <= a;
    layer3_outputs(863) <= b;
    layer3_outputs(864) <= a and not b;
    layer3_outputs(865) <= a;
    layer3_outputs(866) <= a or b;
    layer3_outputs(867) <= b and not a;
    layer3_outputs(868) <= b and not a;
    layer3_outputs(869) <= a and not b;
    layer3_outputs(870) <= b and not a;
    layer3_outputs(871) <= b;
    layer3_outputs(872) <= not a;
    layer3_outputs(873) <= not (a or b);
    layer3_outputs(874) <= b;
    layer3_outputs(875) <= not a;
    layer3_outputs(876) <= not a;
    layer3_outputs(877) <= b;
    layer3_outputs(878) <= b;
    layer3_outputs(879) <= not (a and b);
    layer3_outputs(880) <= not a or b;
    layer3_outputs(881) <= not a or b;
    layer3_outputs(882) <= not (a or b);
    layer3_outputs(883) <= a xor b;
    layer3_outputs(884) <= a and not b;
    layer3_outputs(885) <= not (a or b);
    layer3_outputs(886) <= not (a xor b);
    layer3_outputs(887) <= 1'b1;
    layer3_outputs(888) <= a and not b;
    layer3_outputs(889) <= not a or b;
    layer3_outputs(890) <= not a or b;
    layer3_outputs(891) <= a and not b;
    layer3_outputs(892) <= a;
    layer3_outputs(893) <= not (a xor b);
    layer3_outputs(894) <= a;
    layer3_outputs(895) <= not (a and b);
    layer3_outputs(896) <= a or b;
    layer3_outputs(897) <= not (a and b);
    layer3_outputs(898) <= a and not b;
    layer3_outputs(899) <= not (a or b);
    layer3_outputs(900) <= not b;
    layer3_outputs(901) <= not a or b;
    layer3_outputs(902) <= a;
    layer3_outputs(903) <= a;
    layer3_outputs(904) <= a xor b;
    layer3_outputs(905) <= b;
    layer3_outputs(906) <= a;
    layer3_outputs(907) <= b and not a;
    layer3_outputs(908) <= not b or a;
    layer3_outputs(909) <= not a;
    layer3_outputs(910) <= not (a and b);
    layer3_outputs(911) <= not a or b;
    layer3_outputs(912) <= b and not a;
    layer3_outputs(913) <= a and not b;
    layer3_outputs(914) <= not b;
    layer3_outputs(915) <= not (a or b);
    layer3_outputs(916) <= b;
    layer3_outputs(917) <= a;
    layer3_outputs(918) <= a;
    layer3_outputs(919) <= not a or b;
    layer3_outputs(920) <= not a;
    layer3_outputs(921) <= a and not b;
    layer3_outputs(922) <= 1'b0;
    layer3_outputs(923) <= a;
    layer3_outputs(924) <= 1'b1;
    layer3_outputs(925) <= not (a or b);
    layer3_outputs(926) <= b and not a;
    layer3_outputs(927) <= 1'b1;
    layer3_outputs(928) <= b;
    layer3_outputs(929) <= a;
    layer3_outputs(930) <= a;
    layer3_outputs(931) <= a xor b;
    layer3_outputs(932) <= b;
    layer3_outputs(933) <= a and b;
    layer3_outputs(934) <= a and not b;
    layer3_outputs(935) <= a;
    layer3_outputs(936) <= a;
    layer3_outputs(937) <= not a;
    layer3_outputs(938) <= not a or b;
    layer3_outputs(939) <= not (a and b);
    layer3_outputs(940) <= a;
    layer3_outputs(941) <= not a;
    layer3_outputs(942) <= a and not b;
    layer3_outputs(943) <= not (a and b);
    layer3_outputs(944) <= a and b;
    layer3_outputs(945) <= not b;
    layer3_outputs(946) <= b;
    layer3_outputs(947) <= a;
    layer3_outputs(948) <= a xor b;
    layer3_outputs(949) <= not b;
    layer3_outputs(950) <= not a or b;
    layer3_outputs(951) <= a and not b;
    layer3_outputs(952) <= not (a or b);
    layer3_outputs(953) <= a or b;
    layer3_outputs(954) <= a and b;
    layer3_outputs(955) <= a or b;
    layer3_outputs(956) <= not b or a;
    layer3_outputs(957) <= not a;
    layer3_outputs(958) <= a;
    layer3_outputs(959) <= b and not a;
    layer3_outputs(960) <= b and not a;
    layer3_outputs(961) <= not a or b;
    layer3_outputs(962) <= a or b;
    layer3_outputs(963) <= a and not b;
    layer3_outputs(964) <= not (a or b);
    layer3_outputs(965) <= a and not b;
    layer3_outputs(966) <= not (a and b);
    layer3_outputs(967) <= a;
    layer3_outputs(968) <= not (a xor b);
    layer3_outputs(969) <= 1'b1;
    layer3_outputs(970) <= a;
    layer3_outputs(971) <= not (a and b);
    layer3_outputs(972) <= not b or a;
    layer3_outputs(973) <= b;
    layer3_outputs(974) <= a and not b;
    layer3_outputs(975) <= not a;
    layer3_outputs(976) <= a and not b;
    layer3_outputs(977) <= not b or a;
    layer3_outputs(978) <= not (a and b);
    layer3_outputs(979) <= not b;
    layer3_outputs(980) <= not a;
    layer3_outputs(981) <= a or b;
    layer3_outputs(982) <= b;
    layer3_outputs(983) <= not b;
    layer3_outputs(984) <= 1'b1;
    layer3_outputs(985) <= not b;
    layer3_outputs(986) <= b and not a;
    layer3_outputs(987) <= not b;
    layer3_outputs(988) <= not (a and b);
    layer3_outputs(989) <= not b;
    layer3_outputs(990) <= not b;
    layer3_outputs(991) <= 1'b0;
    layer3_outputs(992) <= a and not b;
    layer3_outputs(993) <= a and b;
    layer3_outputs(994) <= b;
    layer3_outputs(995) <= a;
    layer3_outputs(996) <= a or b;
    layer3_outputs(997) <= a and not b;
    layer3_outputs(998) <= not a;
    layer3_outputs(999) <= not a or b;
    layer3_outputs(1000) <= not (a and b);
    layer3_outputs(1001) <= a;
    layer3_outputs(1002) <= a xor b;
    layer3_outputs(1003) <= b;
    layer3_outputs(1004) <= a and b;
    layer3_outputs(1005) <= b and not a;
    layer3_outputs(1006) <= a or b;
    layer3_outputs(1007) <= a and not b;
    layer3_outputs(1008) <= not (a xor b);
    layer3_outputs(1009) <= 1'b1;
    layer3_outputs(1010) <= b;
    layer3_outputs(1011) <= not b;
    layer3_outputs(1012) <= a;
    layer3_outputs(1013) <= not a;
    layer3_outputs(1014) <= not a;
    layer3_outputs(1015) <= a or b;
    layer3_outputs(1016) <= a;
    layer3_outputs(1017) <= not (a xor b);
    layer3_outputs(1018) <= not a;
    layer3_outputs(1019) <= a;
    layer3_outputs(1020) <= a;
    layer3_outputs(1021) <= not a or b;
    layer3_outputs(1022) <= not a or b;
    layer3_outputs(1023) <= not a;
    layer3_outputs(1024) <= not b;
    layer3_outputs(1025) <= 1'b1;
    layer3_outputs(1026) <= not b;
    layer3_outputs(1027) <= b;
    layer3_outputs(1028) <= not b or a;
    layer3_outputs(1029) <= not a;
    layer3_outputs(1030) <= not (a and b);
    layer3_outputs(1031) <= not a or b;
    layer3_outputs(1032) <= a;
    layer3_outputs(1033) <= not a;
    layer3_outputs(1034) <= not b;
    layer3_outputs(1035) <= not b or a;
    layer3_outputs(1036) <= a or b;
    layer3_outputs(1037) <= not a;
    layer3_outputs(1038) <= not (a xor b);
    layer3_outputs(1039) <= 1'b1;
    layer3_outputs(1040) <= b and not a;
    layer3_outputs(1041) <= 1'b1;
    layer3_outputs(1042) <= not a;
    layer3_outputs(1043) <= b and not a;
    layer3_outputs(1044) <= b;
    layer3_outputs(1045) <= 1'b1;
    layer3_outputs(1046) <= b;
    layer3_outputs(1047) <= a and not b;
    layer3_outputs(1048) <= b;
    layer3_outputs(1049) <= not (a or b);
    layer3_outputs(1050) <= a;
    layer3_outputs(1051) <= not b;
    layer3_outputs(1052) <= not a or b;
    layer3_outputs(1053) <= a and b;
    layer3_outputs(1054) <= a and not b;
    layer3_outputs(1055) <= not (a and b);
    layer3_outputs(1056) <= a or b;
    layer3_outputs(1057) <= 1'b0;
    layer3_outputs(1058) <= b and not a;
    layer3_outputs(1059) <= not (a and b);
    layer3_outputs(1060) <= not (a xor b);
    layer3_outputs(1061) <= not a;
    layer3_outputs(1062) <= not b or a;
    layer3_outputs(1063) <= a and not b;
    layer3_outputs(1064) <= a and b;
    layer3_outputs(1065) <= not a;
    layer3_outputs(1066) <= a and b;
    layer3_outputs(1067) <= not a;
    layer3_outputs(1068) <= a xor b;
    layer3_outputs(1069) <= b and not a;
    layer3_outputs(1070) <= b;
    layer3_outputs(1071) <= a;
    layer3_outputs(1072) <= a xor b;
    layer3_outputs(1073) <= b;
    layer3_outputs(1074) <= not (a and b);
    layer3_outputs(1075) <= not a;
    layer3_outputs(1076) <= a and not b;
    layer3_outputs(1077) <= not a or b;
    layer3_outputs(1078) <= 1'b0;
    layer3_outputs(1079) <= b and not a;
    layer3_outputs(1080) <= not (a and b);
    layer3_outputs(1081) <= not b;
    layer3_outputs(1082) <= not a;
    layer3_outputs(1083) <= a and b;
    layer3_outputs(1084) <= not a;
    layer3_outputs(1085) <= not (a or b);
    layer3_outputs(1086) <= 1'b1;
    layer3_outputs(1087) <= not b or a;
    layer3_outputs(1088) <= not a;
    layer3_outputs(1089) <= a and not b;
    layer3_outputs(1090) <= not b or a;
    layer3_outputs(1091) <= not (a or b);
    layer3_outputs(1092) <= not a;
    layer3_outputs(1093) <= not a or b;
    layer3_outputs(1094) <= 1'b0;
    layer3_outputs(1095) <= not a;
    layer3_outputs(1096) <= 1'b0;
    layer3_outputs(1097) <= not (a xor b);
    layer3_outputs(1098) <= not a;
    layer3_outputs(1099) <= not b or a;
    layer3_outputs(1100) <= not (a xor b);
    layer3_outputs(1101) <= not a or b;
    layer3_outputs(1102) <= not a or b;
    layer3_outputs(1103) <= b;
    layer3_outputs(1104) <= a or b;
    layer3_outputs(1105) <= not a or b;
    layer3_outputs(1106) <= b;
    layer3_outputs(1107) <= not a;
    layer3_outputs(1108) <= not (a and b);
    layer3_outputs(1109) <= b and not a;
    layer3_outputs(1110) <= not a;
    layer3_outputs(1111) <= 1'b1;
    layer3_outputs(1112) <= not b;
    layer3_outputs(1113) <= a or b;
    layer3_outputs(1114) <= not (a or b);
    layer3_outputs(1115) <= a and b;
    layer3_outputs(1116) <= a or b;
    layer3_outputs(1117) <= a;
    layer3_outputs(1118) <= not a or b;
    layer3_outputs(1119) <= a and not b;
    layer3_outputs(1120) <= not (a or b);
    layer3_outputs(1121) <= not (a or b);
    layer3_outputs(1122) <= a xor b;
    layer3_outputs(1123) <= not (a and b);
    layer3_outputs(1124) <= b and not a;
    layer3_outputs(1125) <= not (a and b);
    layer3_outputs(1126) <= a or b;
    layer3_outputs(1127) <= not a;
    layer3_outputs(1128) <= 1'b1;
    layer3_outputs(1129) <= not b or a;
    layer3_outputs(1130) <= b;
    layer3_outputs(1131) <= not a or b;
    layer3_outputs(1132) <= a and not b;
    layer3_outputs(1133) <= a and b;
    layer3_outputs(1134) <= a and not b;
    layer3_outputs(1135) <= a and not b;
    layer3_outputs(1136) <= b;
    layer3_outputs(1137) <= b;
    layer3_outputs(1138) <= not b;
    layer3_outputs(1139) <= not b;
    layer3_outputs(1140) <= not (a and b);
    layer3_outputs(1141) <= not (a xor b);
    layer3_outputs(1142) <= 1'b0;
    layer3_outputs(1143) <= b;
    layer3_outputs(1144) <= not a or b;
    layer3_outputs(1145) <= a and b;
    layer3_outputs(1146) <= a;
    layer3_outputs(1147) <= a xor b;
    layer3_outputs(1148) <= not (a or b);
    layer3_outputs(1149) <= a and not b;
    layer3_outputs(1150) <= a;
    layer3_outputs(1151) <= b;
    layer3_outputs(1152) <= a and not b;
    layer3_outputs(1153) <= b;
    layer3_outputs(1154) <= not (a and b);
    layer3_outputs(1155) <= not (a or b);
    layer3_outputs(1156) <= b;
    layer3_outputs(1157) <= b;
    layer3_outputs(1158) <= not (a and b);
    layer3_outputs(1159) <= a;
    layer3_outputs(1160) <= b and not a;
    layer3_outputs(1161) <= b;
    layer3_outputs(1162) <= not a or b;
    layer3_outputs(1163) <= a and not b;
    layer3_outputs(1164) <= 1'b0;
    layer3_outputs(1165) <= not (a xor b);
    layer3_outputs(1166) <= not a or b;
    layer3_outputs(1167) <= not (a and b);
    layer3_outputs(1168) <= not b or a;
    layer3_outputs(1169) <= not a;
    layer3_outputs(1170) <= a and b;
    layer3_outputs(1171) <= not a or b;
    layer3_outputs(1172) <= not (a or b);
    layer3_outputs(1173) <= a;
    layer3_outputs(1174) <= b and not a;
    layer3_outputs(1175) <= not b or a;
    layer3_outputs(1176) <= a or b;
    layer3_outputs(1177) <= not b;
    layer3_outputs(1178) <= a or b;
    layer3_outputs(1179) <= b;
    layer3_outputs(1180) <= not (a and b);
    layer3_outputs(1181) <= a;
    layer3_outputs(1182) <= a or b;
    layer3_outputs(1183) <= a or b;
    layer3_outputs(1184) <= 1'b0;
    layer3_outputs(1185) <= a and b;
    layer3_outputs(1186) <= not b;
    layer3_outputs(1187) <= not b;
    layer3_outputs(1188) <= not (a and b);
    layer3_outputs(1189) <= b;
    layer3_outputs(1190) <= a or b;
    layer3_outputs(1191) <= a xor b;
    layer3_outputs(1192) <= b and not a;
    layer3_outputs(1193) <= not (a and b);
    layer3_outputs(1194) <= 1'b1;
    layer3_outputs(1195) <= 1'b1;
    layer3_outputs(1196) <= b;
    layer3_outputs(1197) <= b;
    layer3_outputs(1198) <= a xor b;
    layer3_outputs(1199) <= not (a or b);
    layer3_outputs(1200) <= not (a xor b);
    layer3_outputs(1201) <= not (a and b);
    layer3_outputs(1202) <= a and not b;
    layer3_outputs(1203) <= not b;
    layer3_outputs(1204) <= a xor b;
    layer3_outputs(1205) <= a and b;
    layer3_outputs(1206) <= not a or b;
    layer3_outputs(1207) <= not (a or b);
    layer3_outputs(1208) <= a or b;
    layer3_outputs(1209) <= a and not b;
    layer3_outputs(1210) <= not (a or b);
    layer3_outputs(1211) <= b and not a;
    layer3_outputs(1212) <= 1'b1;
    layer3_outputs(1213) <= a;
    layer3_outputs(1214) <= not a;
    layer3_outputs(1215) <= a or b;
    layer3_outputs(1216) <= not b;
    layer3_outputs(1217) <= a;
    layer3_outputs(1218) <= a;
    layer3_outputs(1219) <= b;
    layer3_outputs(1220) <= not b or a;
    layer3_outputs(1221) <= not (a xor b);
    layer3_outputs(1222) <= not a;
    layer3_outputs(1223) <= not b;
    layer3_outputs(1224) <= b and not a;
    layer3_outputs(1225) <= not (a and b);
    layer3_outputs(1226) <= not (a or b);
    layer3_outputs(1227) <= not a;
    layer3_outputs(1228) <= a or b;
    layer3_outputs(1229) <= not (a xor b);
    layer3_outputs(1230) <= not b or a;
    layer3_outputs(1231) <= not (a or b);
    layer3_outputs(1232) <= not b or a;
    layer3_outputs(1233) <= a;
    layer3_outputs(1234) <= a or b;
    layer3_outputs(1235) <= a and not b;
    layer3_outputs(1236) <= 1'b1;
    layer3_outputs(1237) <= not b;
    layer3_outputs(1238) <= not (a xor b);
    layer3_outputs(1239) <= 1'b0;
    layer3_outputs(1240) <= b;
    layer3_outputs(1241) <= not (a or b);
    layer3_outputs(1242) <= not (a or b);
    layer3_outputs(1243) <= b and not a;
    layer3_outputs(1244) <= b and not a;
    layer3_outputs(1245) <= not a or b;
    layer3_outputs(1246) <= not a or b;
    layer3_outputs(1247) <= not b;
    layer3_outputs(1248) <= not a or b;
    layer3_outputs(1249) <= not b or a;
    layer3_outputs(1250) <= a and not b;
    layer3_outputs(1251) <= not a;
    layer3_outputs(1252) <= not a;
    layer3_outputs(1253) <= a and not b;
    layer3_outputs(1254) <= b;
    layer3_outputs(1255) <= b;
    layer3_outputs(1256) <= not b or a;
    layer3_outputs(1257) <= a;
    layer3_outputs(1258) <= not b or a;
    layer3_outputs(1259) <= b and not a;
    layer3_outputs(1260) <= a and not b;
    layer3_outputs(1261) <= a and not b;
    layer3_outputs(1262) <= not a;
    layer3_outputs(1263) <= a;
    layer3_outputs(1264) <= a and not b;
    layer3_outputs(1265) <= not (a or b);
    layer3_outputs(1266) <= b;
    layer3_outputs(1267) <= not a;
    layer3_outputs(1268) <= a and b;
    layer3_outputs(1269) <= a or b;
    layer3_outputs(1270) <= a;
    layer3_outputs(1271) <= not a or b;
    layer3_outputs(1272) <= not a or b;
    layer3_outputs(1273) <= not (a and b);
    layer3_outputs(1274) <= not a;
    layer3_outputs(1275) <= not b or a;
    layer3_outputs(1276) <= not b;
    layer3_outputs(1277) <= not (a and b);
    layer3_outputs(1278) <= not (a xor b);
    layer3_outputs(1279) <= not (a and b);
    layer3_outputs(1280) <= not a;
    layer3_outputs(1281) <= not b;
    layer3_outputs(1282) <= not (a and b);
    layer3_outputs(1283) <= not b or a;
    layer3_outputs(1284) <= not a or b;
    layer3_outputs(1285) <= not a;
    layer3_outputs(1286) <= b and not a;
    layer3_outputs(1287) <= not a;
    layer3_outputs(1288) <= a and not b;
    layer3_outputs(1289) <= b and not a;
    layer3_outputs(1290) <= not a;
    layer3_outputs(1291) <= a or b;
    layer3_outputs(1292) <= not a;
    layer3_outputs(1293) <= a;
    layer3_outputs(1294) <= b and not a;
    layer3_outputs(1295) <= 1'b0;
    layer3_outputs(1296) <= not (a xor b);
    layer3_outputs(1297) <= b and not a;
    layer3_outputs(1298) <= a xor b;
    layer3_outputs(1299) <= not a;
    layer3_outputs(1300) <= not a;
    layer3_outputs(1301) <= not a;
    layer3_outputs(1302) <= not (a xor b);
    layer3_outputs(1303) <= not (a or b);
    layer3_outputs(1304) <= not b;
    layer3_outputs(1305) <= not (a or b);
    layer3_outputs(1306) <= not b or a;
    layer3_outputs(1307) <= a and b;
    layer3_outputs(1308) <= a and not b;
    layer3_outputs(1309) <= a;
    layer3_outputs(1310) <= a and b;
    layer3_outputs(1311) <= a;
    layer3_outputs(1312) <= b;
    layer3_outputs(1313) <= b and not a;
    layer3_outputs(1314) <= not (a and b);
    layer3_outputs(1315) <= not b or a;
    layer3_outputs(1316) <= not a;
    layer3_outputs(1317) <= not a or b;
    layer3_outputs(1318) <= b;
    layer3_outputs(1319) <= not b;
    layer3_outputs(1320) <= a xor b;
    layer3_outputs(1321) <= not b;
    layer3_outputs(1322) <= not a;
    layer3_outputs(1323) <= not b or a;
    layer3_outputs(1324) <= not a or b;
    layer3_outputs(1325) <= not (a or b);
    layer3_outputs(1326) <= not (a xor b);
    layer3_outputs(1327) <= a and b;
    layer3_outputs(1328) <= not (a and b);
    layer3_outputs(1329) <= a and b;
    layer3_outputs(1330) <= a;
    layer3_outputs(1331) <= not (a or b);
    layer3_outputs(1332) <= a and not b;
    layer3_outputs(1333) <= not (a xor b);
    layer3_outputs(1334) <= a;
    layer3_outputs(1335) <= a;
    layer3_outputs(1336) <= not a;
    layer3_outputs(1337) <= not a or b;
    layer3_outputs(1338) <= a and b;
    layer3_outputs(1339) <= b;
    layer3_outputs(1340) <= 1'b0;
    layer3_outputs(1341) <= not a or b;
    layer3_outputs(1342) <= a xor b;
    layer3_outputs(1343) <= not (a or b);
    layer3_outputs(1344) <= not b;
    layer3_outputs(1345) <= a and not b;
    layer3_outputs(1346) <= a;
    layer3_outputs(1347) <= b;
    layer3_outputs(1348) <= a;
    layer3_outputs(1349) <= a and b;
    layer3_outputs(1350) <= not (a and b);
    layer3_outputs(1351) <= b and not a;
    layer3_outputs(1352) <= not b;
    layer3_outputs(1353) <= a;
    layer3_outputs(1354) <= not a;
    layer3_outputs(1355) <= not a or b;
    layer3_outputs(1356) <= not b;
    layer3_outputs(1357) <= not a;
    layer3_outputs(1358) <= a and not b;
    layer3_outputs(1359) <= not b;
    layer3_outputs(1360) <= not b;
    layer3_outputs(1361) <= a and b;
    layer3_outputs(1362) <= a and b;
    layer3_outputs(1363) <= not (a and b);
    layer3_outputs(1364) <= b;
    layer3_outputs(1365) <= not b or a;
    layer3_outputs(1366) <= not a;
    layer3_outputs(1367) <= not a or b;
    layer3_outputs(1368) <= a and b;
    layer3_outputs(1369) <= a;
    layer3_outputs(1370) <= not (a xor b);
    layer3_outputs(1371) <= a;
    layer3_outputs(1372) <= not a;
    layer3_outputs(1373) <= b;
    layer3_outputs(1374) <= a;
    layer3_outputs(1375) <= a;
    layer3_outputs(1376) <= a and b;
    layer3_outputs(1377) <= not b or a;
    layer3_outputs(1378) <= not a;
    layer3_outputs(1379) <= b;
    layer3_outputs(1380) <= a and b;
    layer3_outputs(1381) <= a or b;
    layer3_outputs(1382) <= not a;
    layer3_outputs(1383) <= not a;
    layer3_outputs(1384) <= not (a and b);
    layer3_outputs(1385) <= not a or b;
    layer3_outputs(1386) <= not a or b;
    layer3_outputs(1387) <= a;
    layer3_outputs(1388) <= b;
    layer3_outputs(1389) <= a;
    layer3_outputs(1390) <= b;
    layer3_outputs(1391) <= not (a or b);
    layer3_outputs(1392) <= b;
    layer3_outputs(1393) <= not b or a;
    layer3_outputs(1394) <= not (a or b);
    layer3_outputs(1395) <= not a or b;
    layer3_outputs(1396) <= not b;
    layer3_outputs(1397) <= not b or a;
    layer3_outputs(1398) <= not b;
    layer3_outputs(1399) <= not (a and b);
    layer3_outputs(1400) <= not a;
    layer3_outputs(1401) <= a or b;
    layer3_outputs(1402) <= not b or a;
    layer3_outputs(1403) <= not b or a;
    layer3_outputs(1404) <= a and not b;
    layer3_outputs(1405) <= a and not b;
    layer3_outputs(1406) <= not a or b;
    layer3_outputs(1407) <= not a;
    layer3_outputs(1408) <= 1'b1;
    layer3_outputs(1409) <= not b or a;
    layer3_outputs(1410) <= not b;
    layer3_outputs(1411) <= b;
    layer3_outputs(1412) <= not a or b;
    layer3_outputs(1413) <= a and not b;
    layer3_outputs(1414) <= not a;
    layer3_outputs(1415) <= 1'b1;
    layer3_outputs(1416) <= a;
    layer3_outputs(1417) <= a or b;
    layer3_outputs(1418) <= not b or a;
    layer3_outputs(1419) <= not (a or b);
    layer3_outputs(1420) <= a or b;
    layer3_outputs(1421) <= not a;
    layer3_outputs(1422) <= not (a or b);
    layer3_outputs(1423) <= not a or b;
    layer3_outputs(1424) <= not (a and b);
    layer3_outputs(1425) <= not b;
    layer3_outputs(1426) <= a;
    layer3_outputs(1427) <= not b;
    layer3_outputs(1428) <= a and not b;
    layer3_outputs(1429) <= a xor b;
    layer3_outputs(1430) <= a and not b;
    layer3_outputs(1431) <= not (a or b);
    layer3_outputs(1432) <= a and b;
    layer3_outputs(1433) <= b and not a;
    layer3_outputs(1434) <= not (a and b);
    layer3_outputs(1435) <= b and not a;
    layer3_outputs(1436) <= not a or b;
    layer3_outputs(1437) <= not (a and b);
    layer3_outputs(1438) <= a;
    layer3_outputs(1439) <= b and not a;
    layer3_outputs(1440) <= not (a xor b);
    layer3_outputs(1441) <= b and not a;
    layer3_outputs(1442) <= not b or a;
    layer3_outputs(1443) <= not (a xor b);
    layer3_outputs(1444) <= a and b;
    layer3_outputs(1445) <= not a;
    layer3_outputs(1446) <= a or b;
    layer3_outputs(1447) <= b;
    layer3_outputs(1448) <= not a;
    layer3_outputs(1449) <= a;
    layer3_outputs(1450) <= not a;
    layer3_outputs(1451) <= b;
    layer3_outputs(1452) <= not a or b;
    layer3_outputs(1453) <= b and not a;
    layer3_outputs(1454) <= not (a xor b);
    layer3_outputs(1455) <= not b;
    layer3_outputs(1456) <= b;
    layer3_outputs(1457) <= not b;
    layer3_outputs(1458) <= a and b;
    layer3_outputs(1459) <= not (a xor b);
    layer3_outputs(1460) <= b;
    layer3_outputs(1461) <= a;
    layer3_outputs(1462) <= not (a xor b);
    layer3_outputs(1463) <= not b;
    layer3_outputs(1464) <= a and not b;
    layer3_outputs(1465) <= not (a xor b);
    layer3_outputs(1466) <= not a;
    layer3_outputs(1467) <= not (a and b);
    layer3_outputs(1468) <= not a;
    layer3_outputs(1469) <= b and not a;
    layer3_outputs(1470) <= a and b;
    layer3_outputs(1471) <= not (a or b);
    layer3_outputs(1472) <= not (a and b);
    layer3_outputs(1473) <= 1'b1;
    layer3_outputs(1474) <= a and not b;
    layer3_outputs(1475) <= a and not b;
    layer3_outputs(1476) <= b;
    layer3_outputs(1477) <= not a;
    layer3_outputs(1478) <= 1'b0;
    layer3_outputs(1479) <= b;
    layer3_outputs(1480) <= b and not a;
    layer3_outputs(1481) <= a;
    layer3_outputs(1482) <= not a;
    layer3_outputs(1483) <= not (a or b);
    layer3_outputs(1484) <= b;
    layer3_outputs(1485) <= not a or b;
    layer3_outputs(1486) <= not (a xor b);
    layer3_outputs(1487) <= b;
    layer3_outputs(1488) <= a or b;
    layer3_outputs(1489) <= b;
    layer3_outputs(1490) <= a xor b;
    layer3_outputs(1491) <= not b;
    layer3_outputs(1492) <= b and not a;
    layer3_outputs(1493) <= not (a and b);
    layer3_outputs(1494) <= not b;
    layer3_outputs(1495) <= b;
    layer3_outputs(1496) <= b and not a;
    layer3_outputs(1497) <= a and b;
    layer3_outputs(1498) <= a and not b;
    layer3_outputs(1499) <= not b or a;
    layer3_outputs(1500) <= not a or b;
    layer3_outputs(1501) <= not b;
    layer3_outputs(1502) <= not (a and b);
    layer3_outputs(1503) <= a or b;
    layer3_outputs(1504) <= a and b;
    layer3_outputs(1505) <= not (a and b);
    layer3_outputs(1506) <= not b;
    layer3_outputs(1507) <= a xor b;
    layer3_outputs(1508) <= not b;
    layer3_outputs(1509) <= not (a or b);
    layer3_outputs(1510) <= not b;
    layer3_outputs(1511) <= a and b;
    layer3_outputs(1512) <= not (a and b);
    layer3_outputs(1513) <= a and b;
    layer3_outputs(1514) <= not b;
    layer3_outputs(1515) <= a or b;
    layer3_outputs(1516) <= 1'b0;
    layer3_outputs(1517) <= 1'b0;
    layer3_outputs(1518) <= not b or a;
    layer3_outputs(1519) <= b;
    layer3_outputs(1520) <= 1'b0;
    layer3_outputs(1521) <= not b;
    layer3_outputs(1522) <= b and not a;
    layer3_outputs(1523) <= not a or b;
    layer3_outputs(1524) <= 1'b0;
    layer3_outputs(1525) <= not a or b;
    layer3_outputs(1526) <= a or b;
    layer3_outputs(1527) <= not b;
    layer3_outputs(1528) <= not a or b;
    layer3_outputs(1529) <= not (a and b);
    layer3_outputs(1530) <= not b;
    layer3_outputs(1531) <= a or b;
    layer3_outputs(1532) <= not a;
    layer3_outputs(1533) <= not (a or b);
    layer3_outputs(1534) <= not a;
    layer3_outputs(1535) <= a xor b;
    layer3_outputs(1536) <= 1'b0;
    layer3_outputs(1537) <= a or b;
    layer3_outputs(1538) <= not (a or b);
    layer3_outputs(1539) <= not b;
    layer3_outputs(1540) <= not (a or b);
    layer3_outputs(1541) <= b;
    layer3_outputs(1542) <= a xor b;
    layer3_outputs(1543) <= b and not a;
    layer3_outputs(1544) <= a or b;
    layer3_outputs(1545) <= a;
    layer3_outputs(1546) <= 1'b0;
    layer3_outputs(1547) <= a and not b;
    layer3_outputs(1548) <= a;
    layer3_outputs(1549) <= not b;
    layer3_outputs(1550) <= not a or b;
    layer3_outputs(1551) <= not b;
    layer3_outputs(1552) <= a or b;
    layer3_outputs(1553) <= a and b;
    layer3_outputs(1554) <= a and not b;
    layer3_outputs(1555) <= b;
    layer3_outputs(1556) <= not b or a;
    layer3_outputs(1557) <= not b;
    layer3_outputs(1558) <= not a or b;
    layer3_outputs(1559) <= a and not b;
    layer3_outputs(1560) <= not (a or b);
    layer3_outputs(1561) <= a;
    layer3_outputs(1562) <= not a or b;
    layer3_outputs(1563) <= not b or a;
    layer3_outputs(1564) <= not a;
    layer3_outputs(1565) <= a;
    layer3_outputs(1566) <= b and not a;
    layer3_outputs(1567) <= not b or a;
    layer3_outputs(1568) <= not b;
    layer3_outputs(1569) <= not (a xor b);
    layer3_outputs(1570) <= b;
    layer3_outputs(1571) <= a and b;
    layer3_outputs(1572) <= not a;
    layer3_outputs(1573) <= b and not a;
    layer3_outputs(1574) <= a and b;
    layer3_outputs(1575) <= not a;
    layer3_outputs(1576) <= a or b;
    layer3_outputs(1577) <= not a;
    layer3_outputs(1578) <= not (a and b);
    layer3_outputs(1579) <= not a;
    layer3_outputs(1580) <= not b;
    layer3_outputs(1581) <= not b;
    layer3_outputs(1582) <= b;
    layer3_outputs(1583) <= not b;
    layer3_outputs(1584) <= b;
    layer3_outputs(1585) <= b and not a;
    layer3_outputs(1586) <= not b;
    layer3_outputs(1587) <= b and not a;
    layer3_outputs(1588) <= not a;
    layer3_outputs(1589) <= a or b;
    layer3_outputs(1590) <= b and not a;
    layer3_outputs(1591) <= 1'b1;
    layer3_outputs(1592) <= a and not b;
    layer3_outputs(1593) <= b;
    layer3_outputs(1594) <= not b or a;
    layer3_outputs(1595) <= b;
    layer3_outputs(1596) <= not b;
    layer3_outputs(1597) <= not (a xor b);
    layer3_outputs(1598) <= b;
    layer3_outputs(1599) <= not a;
    layer3_outputs(1600) <= not b;
    layer3_outputs(1601) <= not b;
    layer3_outputs(1602) <= not a;
    layer3_outputs(1603) <= not (a or b);
    layer3_outputs(1604) <= not b or a;
    layer3_outputs(1605) <= a xor b;
    layer3_outputs(1606) <= b;
    layer3_outputs(1607) <= a and not b;
    layer3_outputs(1608) <= not b;
    layer3_outputs(1609) <= a or b;
    layer3_outputs(1610) <= a and not b;
    layer3_outputs(1611) <= not a;
    layer3_outputs(1612) <= a or b;
    layer3_outputs(1613) <= not (a or b);
    layer3_outputs(1614) <= not b or a;
    layer3_outputs(1615) <= a or b;
    layer3_outputs(1616) <= a and b;
    layer3_outputs(1617) <= a and not b;
    layer3_outputs(1618) <= not b;
    layer3_outputs(1619) <= a;
    layer3_outputs(1620) <= not b;
    layer3_outputs(1621) <= not (a and b);
    layer3_outputs(1622) <= b;
    layer3_outputs(1623) <= 1'b0;
    layer3_outputs(1624) <= not b;
    layer3_outputs(1625) <= not a;
    layer3_outputs(1626) <= a and not b;
    layer3_outputs(1627) <= not a;
    layer3_outputs(1628) <= 1'b1;
    layer3_outputs(1629) <= a or b;
    layer3_outputs(1630) <= not b;
    layer3_outputs(1631) <= not a or b;
    layer3_outputs(1632) <= b;
    layer3_outputs(1633) <= not a or b;
    layer3_outputs(1634) <= not (a or b);
    layer3_outputs(1635) <= a and b;
    layer3_outputs(1636) <= a;
    layer3_outputs(1637) <= a and not b;
    layer3_outputs(1638) <= a or b;
    layer3_outputs(1639) <= b and not a;
    layer3_outputs(1640) <= a and b;
    layer3_outputs(1641) <= not (a or b);
    layer3_outputs(1642) <= a;
    layer3_outputs(1643) <= not (a and b);
    layer3_outputs(1644) <= not b;
    layer3_outputs(1645) <= a and not b;
    layer3_outputs(1646) <= a;
    layer3_outputs(1647) <= b;
    layer3_outputs(1648) <= not a;
    layer3_outputs(1649) <= not b;
    layer3_outputs(1650) <= b;
    layer3_outputs(1651) <= a or b;
    layer3_outputs(1652) <= not b;
    layer3_outputs(1653) <= a or b;
    layer3_outputs(1654) <= not (a and b);
    layer3_outputs(1655) <= not (a or b);
    layer3_outputs(1656) <= not b or a;
    layer3_outputs(1657) <= not (a or b);
    layer3_outputs(1658) <= not a or b;
    layer3_outputs(1659) <= not a;
    layer3_outputs(1660) <= not b or a;
    layer3_outputs(1661) <= not a;
    layer3_outputs(1662) <= a and not b;
    layer3_outputs(1663) <= a and not b;
    layer3_outputs(1664) <= not a;
    layer3_outputs(1665) <= a and b;
    layer3_outputs(1666) <= not b or a;
    layer3_outputs(1667) <= not a;
    layer3_outputs(1668) <= not a;
    layer3_outputs(1669) <= a and b;
    layer3_outputs(1670) <= a;
    layer3_outputs(1671) <= not (a or b);
    layer3_outputs(1672) <= not b;
    layer3_outputs(1673) <= not b or a;
    layer3_outputs(1674) <= not (a or b);
    layer3_outputs(1675) <= not a or b;
    layer3_outputs(1676) <= not b or a;
    layer3_outputs(1677) <= 1'b0;
    layer3_outputs(1678) <= a or b;
    layer3_outputs(1679) <= b and not a;
    layer3_outputs(1680) <= not a or b;
    layer3_outputs(1681) <= a;
    layer3_outputs(1682) <= a and not b;
    layer3_outputs(1683) <= a;
    layer3_outputs(1684) <= not b or a;
    layer3_outputs(1685) <= not b or a;
    layer3_outputs(1686) <= a;
    layer3_outputs(1687) <= a xor b;
    layer3_outputs(1688) <= not a or b;
    layer3_outputs(1689) <= a or b;
    layer3_outputs(1690) <= not b;
    layer3_outputs(1691) <= b and not a;
    layer3_outputs(1692) <= not (a or b);
    layer3_outputs(1693) <= a and b;
    layer3_outputs(1694) <= a or b;
    layer3_outputs(1695) <= not a;
    layer3_outputs(1696) <= not b or a;
    layer3_outputs(1697) <= 1'b0;
    layer3_outputs(1698) <= not (a xor b);
    layer3_outputs(1699) <= not a;
    layer3_outputs(1700) <= a and b;
    layer3_outputs(1701) <= a;
    layer3_outputs(1702) <= not b;
    layer3_outputs(1703) <= not (a or b);
    layer3_outputs(1704) <= a and not b;
    layer3_outputs(1705) <= not (a xor b);
    layer3_outputs(1706) <= not b;
    layer3_outputs(1707) <= a and b;
    layer3_outputs(1708) <= 1'b1;
    layer3_outputs(1709) <= a and not b;
    layer3_outputs(1710) <= b and not a;
    layer3_outputs(1711) <= not (a or b);
    layer3_outputs(1712) <= a;
    layer3_outputs(1713) <= not b or a;
    layer3_outputs(1714) <= b and not a;
    layer3_outputs(1715) <= b and not a;
    layer3_outputs(1716) <= 1'b0;
    layer3_outputs(1717) <= a or b;
    layer3_outputs(1718) <= not a;
    layer3_outputs(1719) <= not b or a;
    layer3_outputs(1720) <= b;
    layer3_outputs(1721) <= b;
    layer3_outputs(1722) <= a and b;
    layer3_outputs(1723) <= a;
    layer3_outputs(1724) <= not a or b;
    layer3_outputs(1725) <= b;
    layer3_outputs(1726) <= not b;
    layer3_outputs(1727) <= b and not a;
    layer3_outputs(1728) <= a and b;
    layer3_outputs(1729) <= not b;
    layer3_outputs(1730) <= a;
    layer3_outputs(1731) <= b;
    layer3_outputs(1732) <= not a;
    layer3_outputs(1733) <= not (a and b);
    layer3_outputs(1734) <= a;
    layer3_outputs(1735) <= not b or a;
    layer3_outputs(1736) <= not b;
    layer3_outputs(1737) <= not b;
    layer3_outputs(1738) <= not a;
    layer3_outputs(1739) <= a and not b;
    layer3_outputs(1740) <= a or b;
    layer3_outputs(1741) <= a and not b;
    layer3_outputs(1742) <= not b;
    layer3_outputs(1743) <= not b or a;
    layer3_outputs(1744) <= not a;
    layer3_outputs(1745) <= a or b;
    layer3_outputs(1746) <= not b;
    layer3_outputs(1747) <= not a or b;
    layer3_outputs(1748) <= a and b;
    layer3_outputs(1749) <= b;
    layer3_outputs(1750) <= b and not a;
    layer3_outputs(1751) <= not b;
    layer3_outputs(1752) <= a;
    layer3_outputs(1753) <= not a or b;
    layer3_outputs(1754) <= b;
    layer3_outputs(1755) <= not a;
    layer3_outputs(1756) <= a and b;
    layer3_outputs(1757) <= b;
    layer3_outputs(1758) <= 1'b1;
    layer3_outputs(1759) <= not (a or b);
    layer3_outputs(1760) <= not a or b;
    layer3_outputs(1761) <= not a or b;
    layer3_outputs(1762) <= not b;
    layer3_outputs(1763) <= not a or b;
    layer3_outputs(1764) <= not a or b;
    layer3_outputs(1765) <= not a;
    layer3_outputs(1766) <= a and not b;
    layer3_outputs(1767) <= 1'b1;
    layer3_outputs(1768) <= a or b;
    layer3_outputs(1769) <= a and not b;
    layer3_outputs(1770) <= a and not b;
    layer3_outputs(1771) <= a or b;
    layer3_outputs(1772) <= 1'b1;
    layer3_outputs(1773) <= not b or a;
    layer3_outputs(1774) <= not a;
    layer3_outputs(1775) <= b;
    layer3_outputs(1776) <= not (a xor b);
    layer3_outputs(1777) <= b;
    layer3_outputs(1778) <= a and not b;
    layer3_outputs(1779) <= a or b;
    layer3_outputs(1780) <= not (a or b);
    layer3_outputs(1781) <= a;
    layer3_outputs(1782) <= a or b;
    layer3_outputs(1783) <= not a or b;
    layer3_outputs(1784) <= not (a and b);
    layer3_outputs(1785) <= b;
    layer3_outputs(1786) <= not a;
    layer3_outputs(1787) <= a or b;
    layer3_outputs(1788) <= not (a or b);
    layer3_outputs(1789) <= not b;
    layer3_outputs(1790) <= b;
    layer3_outputs(1791) <= not b or a;
    layer3_outputs(1792) <= not (a or b);
    layer3_outputs(1793) <= a and not b;
    layer3_outputs(1794) <= not b;
    layer3_outputs(1795) <= 1'b0;
    layer3_outputs(1796) <= a or b;
    layer3_outputs(1797) <= a or b;
    layer3_outputs(1798) <= not (a or b);
    layer3_outputs(1799) <= b;
    layer3_outputs(1800) <= not a;
    layer3_outputs(1801) <= not (a xor b);
    layer3_outputs(1802) <= not a;
    layer3_outputs(1803) <= b;
    layer3_outputs(1804) <= a;
    layer3_outputs(1805) <= not (a or b);
    layer3_outputs(1806) <= not a;
    layer3_outputs(1807) <= not b or a;
    layer3_outputs(1808) <= b;
    layer3_outputs(1809) <= b;
    layer3_outputs(1810) <= b;
    layer3_outputs(1811) <= not a or b;
    layer3_outputs(1812) <= b;
    layer3_outputs(1813) <= not b;
    layer3_outputs(1814) <= not (a or b);
    layer3_outputs(1815) <= a;
    layer3_outputs(1816) <= b;
    layer3_outputs(1817) <= a and b;
    layer3_outputs(1818) <= a or b;
    layer3_outputs(1819) <= not (a or b);
    layer3_outputs(1820) <= not a;
    layer3_outputs(1821) <= 1'b0;
    layer3_outputs(1822) <= not a or b;
    layer3_outputs(1823) <= not (a or b);
    layer3_outputs(1824) <= b;
    layer3_outputs(1825) <= not a;
    layer3_outputs(1826) <= not (a and b);
    layer3_outputs(1827) <= a and b;
    layer3_outputs(1828) <= not b;
    layer3_outputs(1829) <= a;
    layer3_outputs(1830) <= a or b;
    layer3_outputs(1831) <= not a;
    layer3_outputs(1832) <= not b;
    layer3_outputs(1833) <= a;
    layer3_outputs(1834) <= not a;
    layer3_outputs(1835) <= not (a or b);
    layer3_outputs(1836) <= a and b;
    layer3_outputs(1837) <= b;
    layer3_outputs(1838) <= b;
    layer3_outputs(1839) <= not b or a;
    layer3_outputs(1840) <= a and not b;
    layer3_outputs(1841) <= not b;
    layer3_outputs(1842) <= not (a and b);
    layer3_outputs(1843) <= not b;
    layer3_outputs(1844) <= not a or b;
    layer3_outputs(1845) <= 1'b0;
    layer3_outputs(1846) <= not b;
    layer3_outputs(1847) <= not b;
    layer3_outputs(1848) <= a and not b;
    layer3_outputs(1849) <= not b;
    layer3_outputs(1850) <= a or b;
    layer3_outputs(1851) <= not (a or b);
    layer3_outputs(1852) <= b and not a;
    layer3_outputs(1853) <= not (a and b);
    layer3_outputs(1854) <= a or b;
    layer3_outputs(1855) <= not a;
    layer3_outputs(1856) <= b;
    layer3_outputs(1857) <= not a or b;
    layer3_outputs(1858) <= a;
    layer3_outputs(1859) <= a or b;
    layer3_outputs(1860) <= a;
    layer3_outputs(1861) <= not (a xor b);
    layer3_outputs(1862) <= a;
    layer3_outputs(1863) <= not a;
    layer3_outputs(1864) <= a xor b;
    layer3_outputs(1865) <= b;
    layer3_outputs(1866) <= a;
    layer3_outputs(1867) <= not a;
    layer3_outputs(1868) <= not (a or b);
    layer3_outputs(1869) <= not (a or b);
    layer3_outputs(1870) <= a;
    layer3_outputs(1871) <= not (a or b);
    layer3_outputs(1872) <= not a or b;
    layer3_outputs(1873) <= not (a xor b);
    layer3_outputs(1874) <= not a;
    layer3_outputs(1875) <= not a;
    layer3_outputs(1876) <= not b or a;
    layer3_outputs(1877) <= a or b;
    layer3_outputs(1878) <= a or b;
    layer3_outputs(1879) <= b;
    layer3_outputs(1880) <= a;
    layer3_outputs(1881) <= b and not a;
    layer3_outputs(1882) <= not (a or b);
    layer3_outputs(1883) <= a xor b;
    layer3_outputs(1884) <= a;
    layer3_outputs(1885) <= not a or b;
    layer3_outputs(1886) <= not b;
    layer3_outputs(1887) <= not b or a;
    layer3_outputs(1888) <= not a;
    layer3_outputs(1889) <= a;
    layer3_outputs(1890) <= not b;
    layer3_outputs(1891) <= a and not b;
    layer3_outputs(1892) <= a and b;
    layer3_outputs(1893) <= not a or b;
    layer3_outputs(1894) <= b;
    layer3_outputs(1895) <= not b;
    layer3_outputs(1896) <= b and not a;
    layer3_outputs(1897) <= not (a and b);
    layer3_outputs(1898) <= 1'b1;
    layer3_outputs(1899) <= b;
    layer3_outputs(1900) <= b;
    layer3_outputs(1901) <= b;
    layer3_outputs(1902) <= a;
    layer3_outputs(1903) <= not (a and b);
    layer3_outputs(1904) <= not b;
    layer3_outputs(1905) <= not (a or b);
    layer3_outputs(1906) <= b;
    layer3_outputs(1907) <= a;
    layer3_outputs(1908) <= a or b;
    layer3_outputs(1909) <= a or b;
    layer3_outputs(1910) <= b;
    layer3_outputs(1911) <= a xor b;
    layer3_outputs(1912) <= 1'b1;
    layer3_outputs(1913) <= not a or b;
    layer3_outputs(1914) <= a;
    layer3_outputs(1915) <= a;
    layer3_outputs(1916) <= a and b;
    layer3_outputs(1917) <= not a or b;
    layer3_outputs(1918) <= b and not a;
    layer3_outputs(1919) <= not a;
    layer3_outputs(1920) <= not (a or b);
    layer3_outputs(1921) <= a and b;
    layer3_outputs(1922) <= b and not a;
    layer3_outputs(1923) <= not (a and b);
    layer3_outputs(1924) <= not a;
    layer3_outputs(1925) <= b;
    layer3_outputs(1926) <= a;
    layer3_outputs(1927) <= not a;
    layer3_outputs(1928) <= a and not b;
    layer3_outputs(1929) <= b;
    layer3_outputs(1930) <= b and not a;
    layer3_outputs(1931) <= not (a or b);
    layer3_outputs(1932) <= not (a or b);
    layer3_outputs(1933) <= not (a and b);
    layer3_outputs(1934) <= not a;
    layer3_outputs(1935) <= not a;
    layer3_outputs(1936) <= b;
    layer3_outputs(1937) <= not b;
    layer3_outputs(1938) <= a;
    layer3_outputs(1939) <= not (a or b);
    layer3_outputs(1940) <= not (a or b);
    layer3_outputs(1941) <= not (a xor b);
    layer3_outputs(1942) <= a and not b;
    layer3_outputs(1943) <= a or b;
    layer3_outputs(1944) <= 1'b1;
    layer3_outputs(1945) <= b and not a;
    layer3_outputs(1946) <= a;
    layer3_outputs(1947) <= a xor b;
    layer3_outputs(1948) <= not a or b;
    layer3_outputs(1949) <= a or b;
    layer3_outputs(1950) <= not b or a;
    layer3_outputs(1951) <= a or b;
    layer3_outputs(1952) <= a;
    layer3_outputs(1953) <= not b;
    layer3_outputs(1954) <= b;
    layer3_outputs(1955) <= not a or b;
    layer3_outputs(1956) <= a and b;
    layer3_outputs(1957) <= not b or a;
    layer3_outputs(1958) <= a;
    layer3_outputs(1959) <= b;
    layer3_outputs(1960) <= not (a and b);
    layer3_outputs(1961) <= not b;
    layer3_outputs(1962) <= not b or a;
    layer3_outputs(1963) <= not b;
    layer3_outputs(1964) <= b;
    layer3_outputs(1965) <= b;
    layer3_outputs(1966) <= not b;
    layer3_outputs(1967) <= b and not a;
    layer3_outputs(1968) <= a or b;
    layer3_outputs(1969) <= a and not b;
    layer3_outputs(1970) <= b and not a;
    layer3_outputs(1971) <= a and b;
    layer3_outputs(1972) <= a;
    layer3_outputs(1973) <= not a;
    layer3_outputs(1974) <= not b;
    layer3_outputs(1975) <= a;
    layer3_outputs(1976) <= a and not b;
    layer3_outputs(1977) <= a and not b;
    layer3_outputs(1978) <= not b or a;
    layer3_outputs(1979) <= b;
    layer3_outputs(1980) <= a and b;
    layer3_outputs(1981) <= a and not b;
    layer3_outputs(1982) <= 1'b1;
    layer3_outputs(1983) <= not b or a;
    layer3_outputs(1984) <= b;
    layer3_outputs(1985) <= a;
    layer3_outputs(1986) <= a or b;
    layer3_outputs(1987) <= a;
    layer3_outputs(1988) <= not a;
    layer3_outputs(1989) <= not (a and b);
    layer3_outputs(1990) <= not b;
    layer3_outputs(1991) <= not (a and b);
    layer3_outputs(1992) <= not a;
    layer3_outputs(1993) <= b and not a;
    layer3_outputs(1994) <= not (a or b);
    layer3_outputs(1995) <= b;
    layer3_outputs(1996) <= 1'b0;
    layer3_outputs(1997) <= 1'b0;
    layer3_outputs(1998) <= not (a and b);
    layer3_outputs(1999) <= not b;
    layer3_outputs(2000) <= a and not b;
    layer3_outputs(2001) <= a and b;
    layer3_outputs(2002) <= b and not a;
    layer3_outputs(2003) <= b;
    layer3_outputs(2004) <= a or b;
    layer3_outputs(2005) <= b and not a;
    layer3_outputs(2006) <= not b or a;
    layer3_outputs(2007) <= not a or b;
    layer3_outputs(2008) <= a and not b;
    layer3_outputs(2009) <= a xor b;
    layer3_outputs(2010) <= not b;
    layer3_outputs(2011) <= a;
    layer3_outputs(2012) <= not (a and b);
    layer3_outputs(2013) <= not a;
    layer3_outputs(2014) <= 1'b1;
    layer3_outputs(2015) <= not (a and b);
    layer3_outputs(2016) <= not b;
    layer3_outputs(2017) <= b;
    layer3_outputs(2018) <= not b;
    layer3_outputs(2019) <= not a or b;
    layer3_outputs(2020) <= not a;
    layer3_outputs(2021) <= not b or a;
    layer3_outputs(2022) <= b;
    layer3_outputs(2023) <= a and not b;
    layer3_outputs(2024) <= not (a and b);
    layer3_outputs(2025) <= a;
    layer3_outputs(2026) <= a;
    layer3_outputs(2027) <= b;
    layer3_outputs(2028) <= b and not a;
    layer3_outputs(2029) <= not a or b;
    layer3_outputs(2030) <= a and b;
    layer3_outputs(2031) <= not (a and b);
    layer3_outputs(2032) <= not a;
    layer3_outputs(2033) <= not a;
    layer3_outputs(2034) <= b;
    layer3_outputs(2035) <= a or b;
    layer3_outputs(2036) <= not a;
    layer3_outputs(2037) <= not b or a;
    layer3_outputs(2038) <= a and not b;
    layer3_outputs(2039) <= 1'b0;
    layer3_outputs(2040) <= a and b;
    layer3_outputs(2041) <= not a or b;
    layer3_outputs(2042) <= a;
    layer3_outputs(2043) <= b;
    layer3_outputs(2044) <= a and not b;
    layer3_outputs(2045) <= b;
    layer3_outputs(2046) <= a and b;
    layer3_outputs(2047) <= not (a or b);
    layer3_outputs(2048) <= a or b;
    layer3_outputs(2049) <= not (a or b);
    layer3_outputs(2050) <= a or b;
    layer3_outputs(2051) <= a and not b;
    layer3_outputs(2052) <= not (a or b);
    layer3_outputs(2053) <= not a or b;
    layer3_outputs(2054) <= a;
    layer3_outputs(2055) <= a and not b;
    layer3_outputs(2056) <= not a or b;
    layer3_outputs(2057) <= not b or a;
    layer3_outputs(2058) <= not b;
    layer3_outputs(2059) <= a;
    layer3_outputs(2060) <= b and not a;
    layer3_outputs(2061) <= not b;
    layer3_outputs(2062) <= a and b;
    layer3_outputs(2063) <= 1'b0;
    layer3_outputs(2064) <= not (a and b);
    layer3_outputs(2065) <= a and b;
    layer3_outputs(2066) <= not b;
    layer3_outputs(2067) <= b and not a;
    layer3_outputs(2068) <= not (a xor b);
    layer3_outputs(2069) <= not b;
    layer3_outputs(2070) <= 1'b0;
    layer3_outputs(2071) <= b;
    layer3_outputs(2072) <= not (a xor b);
    layer3_outputs(2073) <= 1'b0;
    layer3_outputs(2074) <= not b or a;
    layer3_outputs(2075) <= not b or a;
    layer3_outputs(2076) <= a and not b;
    layer3_outputs(2077) <= b and not a;
    layer3_outputs(2078) <= 1'b0;
    layer3_outputs(2079) <= not a or b;
    layer3_outputs(2080) <= a and not b;
    layer3_outputs(2081) <= not (a or b);
    layer3_outputs(2082) <= not b;
    layer3_outputs(2083) <= a and not b;
    layer3_outputs(2084) <= 1'b0;
    layer3_outputs(2085) <= not (a or b);
    layer3_outputs(2086) <= 1'b1;
    layer3_outputs(2087) <= not a;
    layer3_outputs(2088) <= a and not b;
    layer3_outputs(2089) <= a and not b;
    layer3_outputs(2090) <= not b;
    layer3_outputs(2091) <= b and not a;
    layer3_outputs(2092) <= a and not b;
    layer3_outputs(2093) <= a or b;
    layer3_outputs(2094) <= a or b;
    layer3_outputs(2095) <= a and not b;
    layer3_outputs(2096) <= not (a and b);
    layer3_outputs(2097) <= a;
    layer3_outputs(2098) <= not (a and b);
    layer3_outputs(2099) <= not (a or b);
    layer3_outputs(2100) <= not b;
    layer3_outputs(2101) <= not b or a;
    layer3_outputs(2102) <= a;
    layer3_outputs(2103) <= not b;
    layer3_outputs(2104) <= not (a xor b);
    layer3_outputs(2105) <= b;
    layer3_outputs(2106) <= b;
    layer3_outputs(2107) <= not (a and b);
    layer3_outputs(2108) <= 1'b0;
    layer3_outputs(2109) <= not b;
    layer3_outputs(2110) <= a;
    layer3_outputs(2111) <= not b or a;
    layer3_outputs(2112) <= a or b;
    layer3_outputs(2113) <= not a or b;
    layer3_outputs(2114) <= not a or b;
    layer3_outputs(2115) <= not (a and b);
    layer3_outputs(2116) <= a;
    layer3_outputs(2117) <= not b or a;
    layer3_outputs(2118) <= b;
    layer3_outputs(2119) <= not a;
    layer3_outputs(2120) <= a and not b;
    layer3_outputs(2121) <= not b;
    layer3_outputs(2122) <= a and not b;
    layer3_outputs(2123) <= not b;
    layer3_outputs(2124) <= a;
    layer3_outputs(2125) <= not b;
    layer3_outputs(2126) <= not a or b;
    layer3_outputs(2127) <= not (a or b);
    layer3_outputs(2128) <= a and not b;
    layer3_outputs(2129) <= not b or a;
    layer3_outputs(2130) <= not b or a;
    layer3_outputs(2131) <= not b or a;
    layer3_outputs(2132) <= not (a xor b);
    layer3_outputs(2133) <= not (a xor b);
    layer3_outputs(2134) <= not a or b;
    layer3_outputs(2135) <= b;
    layer3_outputs(2136) <= a;
    layer3_outputs(2137) <= b and not a;
    layer3_outputs(2138) <= 1'b1;
    layer3_outputs(2139) <= a or b;
    layer3_outputs(2140) <= 1'b1;
    layer3_outputs(2141) <= a and b;
    layer3_outputs(2142) <= a or b;
    layer3_outputs(2143) <= a;
    layer3_outputs(2144) <= b;
    layer3_outputs(2145) <= not a;
    layer3_outputs(2146) <= b;
    layer3_outputs(2147) <= not (a or b);
    layer3_outputs(2148) <= a and b;
    layer3_outputs(2149) <= not a;
    layer3_outputs(2150) <= not b or a;
    layer3_outputs(2151) <= not (a and b);
    layer3_outputs(2152) <= not a;
    layer3_outputs(2153) <= not a or b;
    layer3_outputs(2154) <= b;
    layer3_outputs(2155) <= b and not a;
    layer3_outputs(2156) <= a;
    layer3_outputs(2157) <= a;
    layer3_outputs(2158) <= a and not b;
    layer3_outputs(2159) <= a;
    layer3_outputs(2160) <= b and not a;
    layer3_outputs(2161) <= not (a or b);
    layer3_outputs(2162) <= not a;
    layer3_outputs(2163) <= a xor b;
    layer3_outputs(2164) <= b and not a;
    layer3_outputs(2165) <= a and b;
    layer3_outputs(2166) <= not b;
    layer3_outputs(2167) <= not b or a;
    layer3_outputs(2168) <= not (a and b);
    layer3_outputs(2169) <= not (a or b);
    layer3_outputs(2170) <= a and b;
    layer3_outputs(2171) <= a and b;
    layer3_outputs(2172) <= b;
    layer3_outputs(2173) <= not b;
    layer3_outputs(2174) <= a and b;
    layer3_outputs(2175) <= not b;
    layer3_outputs(2176) <= a;
    layer3_outputs(2177) <= not b or a;
    layer3_outputs(2178) <= b;
    layer3_outputs(2179) <= not a or b;
    layer3_outputs(2180) <= not b;
    layer3_outputs(2181) <= a;
    layer3_outputs(2182) <= b;
    layer3_outputs(2183) <= not b;
    layer3_outputs(2184) <= not (a and b);
    layer3_outputs(2185) <= not (a xor b);
    layer3_outputs(2186) <= b;
    layer3_outputs(2187) <= not b or a;
    layer3_outputs(2188) <= a or b;
    layer3_outputs(2189) <= b;
    layer3_outputs(2190) <= not (a xor b);
    layer3_outputs(2191) <= not b;
    layer3_outputs(2192) <= b and not a;
    layer3_outputs(2193) <= not b;
    layer3_outputs(2194) <= a and b;
    layer3_outputs(2195) <= not b;
    layer3_outputs(2196) <= a;
    layer3_outputs(2197) <= a or b;
    layer3_outputs(2198) <= b;
    layer3_outputs(2199) <= not (a xor b);
    layer3_outputs(2200) <= 1'b0;
    layer3_outputs(2201) <= a or b;
    layer3_outputs(2202) <= a;
    layer3_outputs(2203) <= not (a or b);
    layer3_outputs(2204) <= a;
    layer3_outputs(2205) <= not a or b;
    layer3_outputs(2206) <= not a;
    layer3_outputs(2207) <= b and not a;
    layer3_outputs(2208) <= not (a xor b);
    layer3_outputs(2209) <= not a;
    layer3_outputs(2210) <= not (a and b);
    layer3_outputs(2211) <= not a;
    layer3_outputs(2212) <= not b;
    layer3_outputs(2213) <= not b;
    layer3_outputs(2214) <= b and not a;
    layer3_outputs(2215) <= a and not b;
    layer3_outputs(2216) <= b;
    layer3_outputs(2217) <= a;
    layer3_outputs(2218) <= a;
    layer3_outputs(2219) <= not b or a;
    layer3_outputs(2220) <= a;
    layer3_outputs(2221) <= not a;
    layer3_outputs(2222) <= not b;
    layer3_outputs(2223) <= b and not a;
    layer3_outputs(2224) <= a and not b;
    layer3_outputs(2225) <= not b;
    layer3_outputs(2226) <= a xor b;
    layer3_outputs(2227) <= not (a or b);
    layer3_outputs(2228) <= b;
    layer3_outputs(2229) <= not b;
    layer3_outputs(2230) <= b;
    layer3_outputs(2231) <= not (a and b);
    layer3_outputs(2232) <= a xor b;
    layer3_outputs(2233) <= 1'b1;
    layer3_outputs(2234) <= b and not a;
    layer3_outputs(2235) <= not a;
    layer3_outputs(2236) <= not b;
    layer3_outputs(2237) <= b and not a;
    layer3_outputs(2238) <= b;
    layer3_outputs(2239) <= not a;
    layer3_outputs(2240) <= b;
    layer3_outputs(2241) <= b;
    layer3_outputs(2242) <= a and b;
    layer3_outputs(2243) <= not b;
    layer3_outputs(2244) <= not a or b;
    layer3_outputs(2245) <= a or b;
    layer3_outputs(2246) <= a and b;
    layer3_outputs(2247) <= b and not a;
    layer3_outputs(2248) <= a;
    layer3_outputs(2249) <= a xor b;
    layer3_outputs(2250) <= not (a and b);
    layer3_outputs(2251) <= not b;
    layer3_outputs(2252) <= a;
    layer3_outputs(2253) <= not (a xor b);
    layer3_outputs(2254) <= b and not a;
    layer3_outputs(2255) <= not b;
    layer3_outputs(2256) <= not (a xor b);
    layer3_outputs(2257) <= not b or a;
    layer3_outputs(2258) <= not b or a;
    layer3_outputs(2259) <= not (a and b);
    layer3_outputs(2260) <= not (a and b);
    layer3_outputs(2261) <= a and not b;
    layer3_outputs(2262) <= a and not b;
    layer3_outputs(2263) <= 1'b1;
    layer3_outputs(2264) <= a;
    layer3_outputs(2265) <= not (a and b);
    layer3_outputs(2266) <= b and not a;
    layer3_outputs(2267) <= a;
    layer3_outputs(2268) <= a xor b;
    layer3_outputs(2269) <= not (a or b);
    layer3_outputs(2270) <= not b or a;
    layer3_outputs(2271) <= a;
    layer3_outputs(2272) <= not a;
    layer3_outputs(2273) <= not b;
    layer3_outputs(2274) <= a;
    layer3_outputs(2275) <= not a or b;
    layer3_outputs(2276) <= a;
    layer3_outputs(2277) <= a;
    layer3_outputs(2278) <= not (a xor b);
    layer3_outputs(2279) <= b;
    layer3_outputs(2280) <= a;
    layer3_outputs(2281) <= 1'b1;
    layer3_outputs(2282) <= not a;
    layer3_outputs(2283) <= not (a xor b);
    layer3_outputs(2284) <= 1'b0;
    layer3_outputs(2285) <= a;
    layer3_outputs(2286) <= a and not b;
    layer3_outputs(2287) <= a;
    layer3_outputs(2288) <= not a;
    layer3_outputs(2289) <= not a;
    layer3_outputs(2290) <= 1'b0;
    layer3_outputs(2291) <= 1'b0;
    layer3_outputs(2292) <= not b;
    layer3_outputs(2293) <= a;
    layer3_outputs(2294) <= a and not b;
    layer3_outputs(2295) <= a;
    layer3_outputs(2296) <= b;
    layer3_outputs(2297) <= not b or a;
    layer3_outputs(2298) <= not b or a;
    layer3_outputs(2299) <= not (a and b);
    layer3_outputs(2300) <= not b;
    layer3_outputs(2301) <= not b or a;
    layer3_outputs(2302) <= not b or a;
    layer3_outputs(2303) <= b;
    layer3_outputs(2304) <= not b or a;
    layer3_outputs(2305) <= a and b;
    layer3_outputs(2306) <= not (a and b);
    layer3_outputs(2307) <= not a or b;
    layer3_outputs(2308) <= not a;
    layer3_outputs(2309) <= not a;
    layer3_outputs(2310) <= not a or b;
    layer3_outputs(2311) <= a or b;
    layer3_outputs(2312) <= a and not b;
    layer3_outputs(2313) <= a and b;
    layer3_outputs(2314) <= not a;
    layer3_outputs(2315) <= not a;
    layer3_outputs(2316) <= b;
    layer3_outputs(2317) <= b;
    layer3_outputs(2318) <= a xor b;
    layer3_outputs(2319) <= not a or b;
    layer3_outputs(2320) <= not a;
    layer3_outputs(2321) <= a;
    layer3_outputs(2322) <= not b or a;
    layer3_outputs(2323) <= b and not a;
    layer3_outputs(2324) <= not b;
    layer3_outputs(2325) <= b;
    layer3_outputs(2326) <= 1'b0;
    layer3_outputs(2327) <= not a;
    layer3_outputs(2328) <= not (a or b);
    layer3_outputs(2329) <= b;
    layer3_outputs(2330) <= a;
    layer3_outputs(2331) <= not b;
    layer3_outputs(2332) <= 1'b1;
    layer3_outputs(2333) <= a;
    layer3_outputs(2334) <= b;
    layer3_outputs(2335) <= a;
    layer3_outputs(2336) <= not a or b;
    layer3_outputs(2337) <= not a;
    layer3_outputs(2338) <= not b;
    layer3_outputs(2339) <= not a;
    layer3_outputs(2340) <= a;
    layer3_outputs(2341) <= not (a or b);
    layer3_outputs(2342) <= a or b;
    layer3_outputs(2343) <= a and b;
    layer3_outputs(2344) <= not a;
    layer3_outputs(2345) <= not (a and b);
    layer3_outputs(2346) <= b and not a;
    layer3_outputs(2347) <= not a;
    layer3_outputs(2348) <= not b;
    layer3_outputs(2349) <= a and b;
    layer3_outputs(2350) <= b and not a;
    layer3_outputs(2351) <= a;
    layer3_outputs(2352) <= b and not a;
    layer3_outputs(2353) <= not a;
    layer3_outputs(2354) <= a and b;
    layer3_outputs(2355) <= 1'b1;
    layer3_outputs(2356) <= not a;
    layer3_outputs(2357) <= a or b;
    layer3_outputs(2358) <= b and not a;
    layer3_outputs(2359) <= b;
    layer3_outputs(2360) <= not a or b;
    layer3_outputs(2361) <= not (a xor b);
    layer3_outputs(2362) <= not (a and b);
    layer3_outputs(2363) <= b and not a;
    layer3_outputs(2364) <= not b;
    layer3_outputs(2365) <= b;
    layer3_outputs(2366) <= not a;
    layer3_outputs(2367) <= not a;
    layer3_outputs(2368) <= not b;
    layer3_outputs(2369) <= b;
    layer3_outputs(2370) <= not b or a;
    layer3_outputs(2371) <= not b;
    layer3_outputs(2372) <= not a;
    layer3_outputs(2373) <= not b;
    layer3_outputs(2374) <= a and b;
    layer3_outputs(2375) <= b;
    layer3_outputs(2376) <= a;
    layer3_outputs(2377) <= b;
    layer3_outputs(2378) <= a or b;
    layer3_outputs(2379) <= a or b;
    layer3_outputs(2380) <= not a;
    layer3_outputs(2381) <= 1'b1;
    layer3_outputs(2382) <= not a or b;
    layer3_outputs(2383) <= a and b;
    layer3_outputs(2384) <= b;
    layer3_outputs(2385) <= not a;
    layer3_outputs(2386) <= not a or b;
    layer3_outputs(2387) <= b;
    layer3_outputs(2388) <= not (a xor b);
    layer3_outputs(2389) <= not (a and b);
    layer3_outputs(2390) <= b;
    layer3_outputs(2391) <= b;
    layer3_outputs(2392) <= a xor b;
    layer3_outputs(2393) <= a or b;
    layer3_outputs(2394) <= a and not b;
    layer3_outputs(2395) <= not b;
    layer3_outputs(2396) <= a and b;
    layer3_outputs(2397) <= not b;
    layer3_outputs(2398) <= not b;
    layer3_outputs(2399) <= a;
    layer3_outputs(2400) <= a and not b;
    layer3_outputs(2401) <= b;
    layer3_outputs(2402) <= a and not b;
    layer3_outputs(2403) <= a;
    layer3_outputs(2404) <= not a;
    layer3_outputs(2405) <= a;
    layer3_outputs(2406) <= a xor b;
    layer3_outputs(2407) <= a and not b;
    layer3_outputs(2408) <= not (a or b);
    layer3_outputs(2409) <= not (a and b);
    layer3_outputs(2410) <= a;
    layer3_outputs(2411) <= a and b;
    layer3_outputs(2412) <= b;
    layer3_outputs(2413) <= not a or b;
    layer3_outputs(2414) <= not (a and b);
    layer3_outputs(2415) <= not (a or b);
    layer3_outputs(2416) <= not b;
    layer3_outputs(2417) <= 1'b1;
    layer3_outputs(2418) <= not b;
    layer3_outputs(2419) <= a and b;
    layer3_outputs(2420) <= not a;
    layer3_outputs(2421) <= a xor b;
    layer3_outputs(2422) <= not a;
    layer3_outputs(2423) <= a and not b;
    layer3_outputs(2424) <= not a;
    layer3_outputs(2425) <= a and not b;
    layer3_outputs(2426) <= b;
    layer3_outputs(2427) <= not b;
    layer3_outputs(2428) <= a;
    layer3_outputs(2429) <= not a;
    layer3_outputs(2430) <= b;
    layer3_outputs(2431) <= not b or a;
    layer3_outputs(2432) <= not b;
    layer3_outputs(2433) <= not b;
    layer3_outputs(2434) <= a and not b;
    layer3_outputs(2435) <= a or b;
    layer3_outputs(2436) <= not a or b;
    layer3_outputs(2437) <= b;
    layer3_outputs(2438) <= not (a or b);
    layer3_outputs(2439) <= not a;
    layer3_outputs(2440) <= a xor b;
    layer3_outputs(2441) <= not b or a;
    layer3_outputs(2442) <= not a;
    layer3_outputs(2443) <= a;
    layer3_outputs(2444) <= not (a or b);
    layer3_outputs(2445) <= b;
    layer3_outputs(2446) <= not (a xor b);
    layer3_outputs(2447) <= a or b;
    layer3_outputs(2448) <= a xor b;
    layer3_outputs(2449) <= not b;
    layer3_outputs(2450) <= a and b;
    layer3_outputs(2451) <= b;
    layer3_outputs(2452) <= not (a and b);
    layer3_outputs(2453) <= b and not a;
    layer3_outputs(2454) <= b;
    layer3_outputs(2455) <= not (a or b);
    layer3_outputs(2456) <= a;
    layer3_outputs(2457) <= a;
    layer3_outputs(2458) <= a;
    layer3_outputs(2459) <= not a;
    layer3_outputs(2460) <= not a;
    layer3_outputs(2461) <= b;
    layer3_outputs(2462) <= a and not b;
    layer3_outputs(2463) <= a;
    layer3_outputs(2464) <= not b or a;
    layer3_outputs(2465) <= a;
    layer3_outputs(2466) <= not a;
    layer3_outputs(2467) <= 1'b0;
    layer3_outputs(2468) <= a xor b;
    layer3_outputs(2469) <= not a;
    layer3_outputs(2470) <= not a;
    layer3_outputs(2471) <= a xor b;
    layer3_outputs(2472) <= not b or a;
    layer3_outputs(2473) <= not a or b;
    layer3_outputs(2474) <= not (a and b);
    layer3_outputs(2475) <= not b;
    layer3_outputs(2476) <= not b or a;
    layer3_outputs(2477) <= 1'b1;
    layer3_outputs(2478) <= not b;
    layer3_outputs(2479) <= a and not b;
    layer3_outputs(2480) <= not (a or b);
    layer3_outputs(2481) <= not (a or b);
    layer3_outputs(2482) <= not b;
    layer3_outputs(2483) <= not (a and b);
    layer3_outputs(2484) <= not a or b;
    layer3_outputs(2485) <= not (a and b);
    layer3_outputs(2486) <= not (a and b);
    layer3_outputs(2487) <= not (a or b);
    layer3_outputs(2488) <= a and not b;
    layer3_outputs(2489) <= a xor b;
    layer3_outputs(2490) <= b and not a;
    layer3_outputs(2491) <= not (a and b);
    layer3_outputs(2492) <= not (a and b);
    layer3_outputs(2493) <= not b;
    layer3_outputs(2494) <= a;
    layer3_outputs(2495) <= not b or a;
    layer3_outputs(2496) <= a;
    layer3_outputs(2497) <= a and not b;
    layer3_outputs(2498) <= not a or b;
    layer3_outputs(2499) <= a and not b;
    layer3_outputs(2500) <= not b or a;
    layer3_outputs(2501) <= not b;
    layer3_outputs(2502) <= not a or b;
    layer3_outputs(2503) <= a and not b;
    layer3_outputs(2504) <= not (a xor b);
    layer3_outputs(2505) <= not a;
    layer3_outputs(2506) <= not a or b;
    layer3_outputs(2507) <= not (a or b);
    layer3_outputs(2508) <= b and not a;
    layer3_outputs(2509) <= not a;
    layer3_outputs(2510) <= a and b;
    layer3_outputs(2511) <= a and not b;
    layer3_outputs(2512) <= not (a and b);
    layer3_outputs(2513) <= a and b;
    layer3_outputs(2514) <= a and b;
    layer3_outputs(2515) <= not b;
    layer3_outputs(2516) <= not b or a;
    layer3_outputs(2517) <= not (a or b);
    layer3_outputs(2518) <= not a;
    layer3_outputs(2519) <= b and not a;
    layer3_outputs(2520) <= not b;
    layer3_outputs(2521) <= b;
    layer3_outputs(2522) <= a and b;
    layer3_outputs(2523) <= a;
    layer3_outputs(2524) <= a;
    layer3_outputs(2525) <= a;
    layer3_outputs(2526) <= not a or b;
    layer3_outputs(2527) <= not (a xor b);
    layer3_outputs(2528) <= not (a or b);
    layer3_outputs(2529) <= not b or a;
    layer3_outputs(2530) <= a and b;
    layer3_outputs(2531) <= not a;
    layer3_outputs(2532) <= b and not a;
    layer3_outputs(2533) <= not b;
    layer3_outputs(2534) <= a;
    layer3_outputs(2535) <= a or b;
    layer3_outputs(2536) <= not a;
    layer3_outputs(2537) <= not b or a;
    layer3_outputs(2538) <= not (a and b);
    layer3_outputs(2539) <= b and not a;
    layer3_outputs(2540) <= a;
    layer3_outputs(2541) <= not (a or b);
    layer3_outputs(2542) <= not b;
    layer3_outputs(2543) <= not a;
    layer3_outputs(2544) <= b;
    layer3_outputs(2545) <= not b or a;
    layer3_outputs(2546) <= b and not a;
    layer3_outputs(2547) <= not b or a;
    layer3_outputs(2548) <= not a or b;
    layer3_outputs(2549) <= not b or a;
    layer3_outputs(2550) <= not b or a;
    layer3_outputs(2551) <= b;
    layer3_outputs(2552) <= not a or b;
    layer3_outputs(2553) <= not b or a;
    layer3_outputs(2554) <= a;
    layer3_outputs(2555) <= b and not a;
    layer3_outputs(2556) <= a or b;
    layer3_outputs(2557) <= not (a xor b);
    layer3_outputs(2558) <= not a;
    layer3_outputs(2559) <= not a;
    layer4_outputs(0) <= not b;
    layer4_outputs(1) <= not a or b;
    layer4_outputs(2) <= not b;
    layer4_outputs(3) <= not (a or b);
    layer4_outputs(4) <= a and not b;
    layer4_outputs(5) <= b and not a;
    layer4_outputs(6) <= 1'b1;
    layer4_outputs(7) <= a or b;
    layer4_outputs(8) <= not (a or b);
    layer4_outputs(9) <= b and not a;
    layer4_outputs(10) <= a and b;
    layer4_outputs(11) <= a;
    layer4_outputs(12) <= a or b;
    layer4_outputs(13) <= not a;
    layer4_outputs(14) <= not b;
    layer4_outputs(15) <= a or b;
    layer4_outputs(16) <= not a;
    layer4_outputs(17) <= not b;
    layer4_outputs(18) <= a or b;
    layer4_outputs(19) <= a xor b;
    layer4_outputs(20) <= not b;
    layer4_outputs(21) <= b and not a;
    layer4_outputs(22) <= not (a and b);
    layer4_outputs(23) <= not b;
    layer4_outputs(24) <= not (a and b);
    layer4_outputs(25) <= a;
    layer4_outputs(26) <= not (a and b);
    layer4_outputs(27) <= not a or b;
    layer4_outputs(28) <= a and not b;
    layer4_outputs(29) <= not b;
    layer4_outputs(30) <= not b;
    layer4_outputs(31) <= b and not a;
    layer4_outputs(32) <= not (a xor b);
    layer4_outputs(33) <= not (a or b);
    layer4_outputs(34) <= not b or a;
    layer4_outputs(35) <= not a;
    layer4_outputs(36) <= not b;
    layer4_outputs(37) <= not a or b;
    layer4_outputs(38) <= not a;
    layer4_outputs(39) <= b;
    layer4_outputs(40) <= not (a or b);
    layer4_outputs(41) <= not b;
    layer4_outputs(42) <= a and b;
    layer4_outputs(43) <= not (a or b);
    layer4_outputs(44) <= a;
    layer4_outputs(45) <= a xor b;
    layer4_outputs(46) <= not a;
    layer4_outputs(47) <= a;
    layer4_outputs(48) <= a and b;
    layer4_outputs(49) <= not b or a;
    layer4_outputs(50) <= b and not a;
    layer4_outputs(51) <= a and b;
    layer4_outputs(52) <= not b;
    layer4_outputs(53) <= b;
    layer4_outputs(54) <= not (a xor b);
    layer4_outputs(55) <= 1'b1;
    layer4_outputs(56) <= not (a or b);
    layer4_outputs(57) <= a or b;
    layer4_outputs(58) <= b;
    layer4_outputs(59) <= b;
    layer4_outputs(60) <= b;
    layer4_outputs(61) <= a;
    layer4_outputs(62) <= a and not b;
    layer4_outputs(63) <= b;
    layer4_outputs(64) <= not a;
    layer4_outputs(65) <= not a or b;
    layer4_outputs(66) <= a;
    layer4_outputs(67) <= not (a and b);
    layer4_outputs(68) <= not b;
    layer4_outputs(69) <= b and not a;
    layer4_outputs(70) <= a;
    layer4_outputs(71) <= not (a xor b);
    layer4_outputs(72) <= not b;
    layer4_outputs(73) <= not b;
    layer4_outputs(74) <= not a;
    layer4_outputs(75) <= not a;
    layer4_outputs(76) <= not (a xor b);
    layer4_outputs(77) <= b and not a;
    layer4_outputs(78) <= not b;
    layer4_outputs(79) <= not (a or b);
    layer4_outputs(80) <= a;
    layer4_outputs(81) <= a and not b;
    layer4_outputs(82) <= not (a or b);
    layer4_outputs(83) <= not b;
    layer4_outputs(84) <= a;
    layer4_outputs(85) <= a;
    layer4_outputs(86) <= a or b;
    layer4_outputs(87) <= not (a xor b);
    layer4_outputs(88) <= not a;
    layer4_outputs(89) <= b and not a;
    layer4_outputs(90) <= not b or a;
    layer4_outputs(91) <= b;
    layer4_outputs(92) <= not (a and b);
    layer4_outputs(93) <= not (a xor b);
    layer4_outputs(94) <= not (a or b);
    layer4_outputs(95) <= not b;
    layer4_outputs(96) <= not b or a;
    layer4_outputs(97) <= not b or a;
    layer4_outputs(98) <= a;
    layer4_outputs(99) <= b;
    layer4_outputs(100) <= not b;
    layer4_outputs(101) <= not a;
    layer4_outputs(102) <= a;
    layer4_outputs(103) <= a and not b;
    layer4_outputs(104) <= not b;
    layer4_outputs(105) <= a xor b;
    layer4_outputs(106) <= not (a xor b);
    layer4_outputs(107) <= a;
    layer4_outputs(108) <= b;
    layer4_outputs(109) <= a;
    layer4_outputs(110) <= a;
    layer4_outputs(111) <= a and b;
    layer4_outputs(112) <= b;
    layer4_outputs(113) <= not b;
    layer4_outputs(114) <= a;
    layer4_outputs(115) <= b;
    layer4_outputs(116) <= b;
    layer4_outputs(117) <= a xor b;
    layer4_outputs(118) <= not a;
    layer4_outputs(119) <= a;
    layer4_outputs(120) <= not (a xor b);
    layer4_outputs(121) <= a or b;
    layer4_outputs(122) <= b;
    layer4_outputs(123) <= not b;
    layer4_outputs(124) <= not (a and b);
    layer4_outputs(125) <= a;
    layer4_outputs(126) <= a and not b;
    layer4_outputs(127) <= not a or b;
    layer4_outputs(128) <= b;
    layer4_outputs(129) <= a;
    layer4_outputs(130) <= a and not b;
    layer4_outputs(131) <= a and b;
    layer4_outputs(132) <= a xor b;
    layer4_outputs(133) <= a xor b;
    layer4_outputs(134) <= a;
    layer4_outputs(135) <= not (a or b);
    layer4_outputs(136) <= not (a or b);
    layer4_outputs(137) <= a or b;
    layer4_outputs(138) <= not a;
    layer4_outputs(139) <= not (a and b);
    layer4_outputs(140) <= b;
    layer4_outputs(141) <= b and not a;
    layer4_outputs(142) <= not b;
    layer4_outputs(143) <= b;
    layer4_outputs(144) <= not a;
    layer4_outputs(145) <= a or b;
    layer4_outputs(146) <= not a or b;
    layer4_outputs(147) <= a;
    layer4_outputs(148) <= b;
    layer4_outputs(149) <= not a or b;
    layer4_outputs(150) <= b and not a;
    layer4_outputs(151) <= not (a or b);
    layer4_outputs(152) <= a and not b;
    layer4_outputs(153) <= b;
    layer4_outputs(154) <= not (a or b);
    layer4_outputs(155) <= a and b;
    layer4_outputs(156) <= not a;
    layer4_outputs(157) <= not (a or b);
    layer4_outputs(158) <= a and b;
    layer4_outputs(159) <= a and b;
    layer4_outputs(160) <= not (a and b);
    layer4_outputs(161) <= not b;
    layer4_outputs(162) <= a and not b;
    layer4_outputs(163) <= not b;
    layer4_outputs(164) <= a;
    layer4_outputs(165) <= not (a xor b);
    layer4_outputs(166) <= b;
    layer4_outputs(167) <= not a;
    layer4_outputs(168) <= a and b;
    layer4_outputs(169) <= not a;
    layer4_outputs(170) <= not (a or b);
    layer4_outputs(171) <= not b or a;
    layer4_outputs(172) <= a or b;
    layer4_outputs(173) <= a and b;
    layer4_outputs(174) <= not b or a;
    layer4_outputs(175) <= not b or a;
    layer4_outputs(176) <= a xor b;
    layer4_outputs(177) <= b;
    layer4_outputs(178) <= a or b;
    layer4_outputs(179) <= b;
    layer4_outputs(180) <= not a;
    layer4_outputs(181) <= b;
    layer4_outputs(182) <= not b;
    layer4_outputs(183) <= a and b;
    layer4_outputs(184) <= a;
    layer4_outputs(185) <= b;
    layer4_outputs(186) <= a xor b;
    layer4_outputs(187) <= not (a or b);
    layer4_outputs(188) <= b and not a;
    layer4_outputs(189) <= not (a xor b);
    layer4_outputs(190) <= b and not a;
    layer4_outputs(191) <= not (a and b);
    layer4_outputs(192) <= b;
    layer4_outputs(193) <= b;
    layer4_outputs(194) <= not a;
    layer4_outputs(195) <= a and b;
    layer4_outputs(196) <= not (a and b);
    layer4_outputs(197) <= b;
    layer4_outputs(198) <= a or b;
    layer4_outputs(199) <= a and b;
    layer4_outputs(200) <= not (a or b);
    layer4_outputs(201) <= a or b;
    layer4_outputs(202) <= a;
    layer4_outputs(203) <= b;
    layer4_outputs(204) <= not a;
    layer4_outputs(205) <= not (a and b);
    layer4_outputs(206) <= a and b;
    layer4_outputs(207) <= b;
    layer4_outputs(208) <= b and not a;
    layer4_outputs(209) <= not (a and b);
    layer4_outputs(210) <= b;
    layer4_outputs(211) <= not (a or b);
    layer4_outputs(212) <= b;
    layer4_outputs(213) <= not (a xor b);
    layer4_outputs(214) <= b;
    layer4_outputs(215) <= not b;
    layer4_outputs(216) <= b and not a;
    layer4_outputs(217) <= a;
    layer4_outputs(218) <= a and not b;
    layer4_outputs(219) <= a or b;
    layer4_outputs(220) <= a;
    layer4_outputs(221) <= a xor b;
    layer4_outputs(222) <= not (a or b);
    layer4_outputs(223) <= a and not b;
    layer4_outputs(224) <= not a;
    layer4_outputs(225) <= not b;
    layer4_outputs(226) <= not a or b;
    layer4_outputs(227) <= not a or b;
    layer4_outputs(228) <= a xor b;
    layer4_outputs(229) <= not b;
    layer4_outputs(230) <= not b or a;
    layer4_outputs(231) <= not (a and b);
    layer4_outputs(232) <= a and b;
    layer4_outputs(233) <= b;
    layer4_outputs(234) <= a;
    layer4_outputs(235) <= a or b;
    layer4_outputs(236) <= not a;
    layer4_outputs(237) <= a;
    layer4_outputs(238) <= not (a xor b);
    layer4_outputs(239) <= not (a and b);
    layer4_outputs(240) <= a;
    layer4_outputs(241) <= not (a xor b);
    layer4_outputs(242) <= not a or b;
    layer4_outputs(243) <= not b or a;
    layer4_outputs(244) <= not a;
    layer4_outputs(245) <= not b or a;
    layer4_outputs(246) <= not (a or b);
    layer4_outputs(247) <= a xor b;
    layer4_outputs(248) <= a and not b;
    layer4_outputs(249) <= not b or a;
    layer4_outputs(250) <= not (a xor b);
    layer4_outputs(251) <= a and b;
    layer4_outputs(252) <= 1'b1;
    layer4_outputs(253) <= a xor b;
    layer4_outputs(254) <= b and not a;
    layer4_outputs(255) <= a and b;
    layer4_outputs(256) <= a;
    layer4_outputs(257) <= b;
    layer4_outputs(258) <= a and b;
    layer4_outputs(259) <= a;
    layer4_outputs(260) <= 1'b1;
    layer4_outputs(261) <= not a;
    layer4_outputs(262) <= not b;
    layer4_outputs(263) <= a;
    layer4_outputs(264) <= a and b;
    layer4_outputs(265) <= b;
    layer4_outputs(266) <= a and not b;
    layer4_outputs(267) <= not b;
    layer4_outputs(268) <= b;
    layer4_outputs(269) <= b;
    layer4_outputs(270) <= not a;
    layer4_outputs(271) <= not a or b;
    layer4_outputs(272) <= 1'b1;
    layer4_outputs(273) <= not (a or b);
    layer4_outputs(274) <= not a;
    layer4_outputs(275) <= not a or b;
    layer4_outputs(276) <= a;
    layer4_outputs(277) <= 1'b1;
    layer4_outputs(278) <= a and b;
    layer4_outputs(279) <= not (a xor b);
    layer4_outputs(280) <= not a;
    layer4_outputs(281) <= not b or a;
    layer4_outputs(282) <= not a or b;
    layer4_outputs(283) <= not (a or b);
    layer4_outputs(284) <= a or b;
    layer4_outputs(285) <= not b;
    layer4_outputs(286) <= a xor b;
    layer4_outputs(287) <= a and not b;
    layer4_outputs(288) <= a and b;
    layer4_outputs(289) <= 1'b0;
    layer4_outputs(290) <= a;
    layer4_outputs(291) <= not b or a;
    layer4_outputs(292) <= a;
    layer4_outputs(293) <= not (a xor b);
    layer4_outputs(294) <= not b;
    layer4_outputs(295) <= not b;
    layer4_outputs(296) <= not b or a;
    layer4_outputs(297) <= a or b;
    layer4_outputs(298) <= not a;
    layer4_outputs(299) <= not (a xor b);
    layer4_outputs(300) <= a;
    layer4_outputs(301) <= a;
    layer4_outputs(302) <= not a;
    layer4_outputs(303) <= a;
    layer4_outputs(304) <= not (a or b);
    layer4_outputs(305) <= not b or a;
    layer4_outputs(306) <= a and not b;
    layer4_outputs(307) <= a and b;
    layer4_outputs(308) <= not b;
    layer4_outputs(309) <= not a or b;
    layer4_outputs(310) <= a;
    layer4_outputs(311) <= not (a xor b);
    layer4_outputs(312) <= not a or b;
    layer4_outputs(313) <= not (a and b);
    layer4_outputs(314) <= not a;
    layer4_outputs(315) <= not b or a;
    layer4_outputs(316) <= not a or b;
    layer4_outputs(317) <= a or b;
    layer4_outputs(318) <= a and b;
    layer4_outputs(319) <= a and b;
    layer4_outputs(320) <= not (a xor b);
    layer4_outputs(321) <= not (a and b);
    layer4_outputs(322) <= not a or b;
    layer4_outputs(323) <= a and b;
    layer4_outputs(324) <= not (a and b);
    layer4_outputs(325) <= b;
    layer4_outputs(326) <= not a;
    layer4_outputs(327) <= not (a or b);
    layer4_outputs(328) <= a and not b;
    layer4_outputs(329) <= not a or b;
    layer4_outputs(330) <= not b;
    layer4_outputs(331) <= not a;
    layer4_outputs(332) <= a;
    layer4_outputs(333) <= b;
    layer4_outputs(334) <= a and not b;
    layer4_outputs(335) <= b;
    layer4_outputs(336) <= not (a or b);
    layer4_outputs(337) <= a;
    layer4_outputs(338) <= a xor b;
    layer4_outputs(339) <= b and not a;
    layer4_outputs(340) <= not a or b;
    layer4_outputs(341) <= b and not a;
    layer4_outputs(342) <= a and not b;
    layer4_outputs(343) <= not a;
    layer4_outputs(344) <= not (a xor b);
    layer4_outputs(345) <= a xor b;
    layer4_outputs(346) <= a and b;
    layer4_outputs(347) <= not (a and b);
    layer4_outputs(348) <= b;
    layer4_outputs(349) <= not (a or b);
    layer4_outputs(350) <= a;
    layer4_outputs(351) <= b and not a;
    layer4_outputs(352) <= not b;
    layer4_outputs(353) <= b;
    layer4_outputs(354) <= b and not a;
    layer4_outputs(355) <= not a;
    layer4_outputs(356) <= a or b;
    layer4_outputs(357) <= b and not a;
    layer4_outputs(358) <= not a;
    layer4_outputs(359) <= not b;
    layer4_outputs(360) <= not (a xor b);
    layer4_outputs(361) <= not a or b;
    layer4_outputs(362) <= a and b;
    layer4_outputs(363) <= a xor b;
    layer4_outputs(364) <= not a or b;
    layer4_outputs(365) <= a and not b;
    layer4_outputs(366) <= a and not b;
    layer4_outputs(367) <= not (a and b);
    layer4_outputs(368) <= not (a or b);
    layer4_outputs(369) <= b;
    layer4_outputs(370) <= b;
    layer4_outputs(371) <= not a or b;
    layer4_outputs(372) <= 1'b0;
    layer4_outputs(373) <= not b;
    layer4_outputs(374) <= a;
    layer4_outputs(375) <= not (a or b);
    layer4_outputs(376) <= not (a and b);
    layer4_outputs(377) <= a and not b;
    layer4_outputs(378) <= not b;
    layer4_outputs(379) <= not b or a;
    layer4_outputs(380) <= not (a and b);
    layer4_outputs(381) <= not (a or b);
    layer4_outputs(382) <= b;
    layer4_outputs(383) <= not (a xor b);
    layer4_outputs(384) <= not (a or b);
    layer4_outputs(385) <= not (a xor b);
    layer4_outputs(386) <= b;
    layer4_outputs(387) <= a;
    layer4_outputs(388) <= not b or a;
    layer4_outputs(389) <= a or b;
    layer4_outputs(390) <= not (a or b);
    layer4_outputs(391) <= a or b;
    layer4_outputs(392) <= a;
    layer4_outputs(393) <= a or b;
    layer4_outputs(394) <= a;
    layer4_outputs(395) <= a or b;
    layer4_outputs(396) <= a;
    layer4_outputs(397) <= not b or a;
    layer4_outputs(398) <= not b or a;
    layer4_outputs(399) <= a;
    layer4_outputs(400) <= a;
    layer4_outputs(401) <= not b;
    layer4_outputs(402) <= not b;
    layer4_outputs(403) <= not a or b;
    layer4_outputs(404) <= not a or b;
    layer4_outputs(405) <= not b;
    layer4_outputs(406) <= not a or b;
    layer4_outputs(407) <= a and b;
    layer4_outputs(408) <= a and b;
    layer4_outputs(409) <= a;
    layer4_outputs(410) <= b and not a;
    layer4_outputs(411) <= not b;
    layer4_outputs(412) <= a and b;
    layer4_outputs(413) <= not b;
    layer4_outputs(414) <= not b;
    layer4_outputs(415) <= not b or a;
    layer4_outputs(416) <= not b;
    layer4_outputs(417) <= not b or a;
    layer4_outputs(418) <= not a;
    layer4_outputs(419) <= not a or b;
    layer4_outputs(420) <= 1'b0;
    layer4_outputs(421) <= a and not b;
    layer4_outputs(422) <= not a or b;
    layer4_outputs(423) <= not b or a;
    layer4_outputs(424) <= not (a or b);
    layer4_outputs(425) <= a xor b;
    layer4_outputs(426) <= not (a or b);
    layer4_outputs(427) <= a or b;
    layer4_outputs(428) <= b;
    layer4_outputs(429) <= not b;
    layer4_outputs(430) <= not b;
    layer4_outputs(431) <= not b;
    layer4_outputs(432) <= a and b;
    layer4_outputs(433) <= not (a xor b);
    layer4_outputs(434) <= not b or a;
    layer4_outputs(435) <= a;
    layer4_outputs(436) <= a or b;
    layer4_outputs(437) <= a or b;
    layer4_outputs(438) <= not (a and b);
    layer4_outputs(439) <= not b;
    layer4_outputs(440) <= not (a or b);
    layer4_outputs(441) <= a;
    layer4_outputs(442) <= not b;
    layer4_outputs(443) <= a and not b;
    layer4_outputs(444) <= not a or b;
    layer4_outputs(445) <= not a or b;
    layer4_outputs(446) <= not (a xor b);
    layer4_outputs(447) <= a;
    layer4_outputs(448) <= a;
    layer4_outputs(449) <= not (a and b);
    layer4_outputs(450) <= not a;
    layer4_outputs(451) <= a xor b;
    layer4_outputs(452) <= not a;
    layer4_outputs(453) <= not a;
    layer4_outputs(454) <= not b or a;
    layer4_outputs(455) <= not b;
    layer4_outputs(456) <= not a;
    layer4_outputs(457) <= not a;
    layer4_outputs(458) <= not (a and b);
    layer4_outputs(459) <= b;
    layer4_outputs(460) <= not a or b;
    layer4_outputs(461) <= not a;
    layer4_outputs(462) <= a or b;
    layer4_outputs(463) <= not (a or b);
    layer4_outputs(464) <= a and b;
    layer4_outputs(465) <= not (a and b);
    layer4_outputs(466) <= not b;
    layer4_outputs(467) <= not (a xor b);
    layer4_outputs(468) <= not b;
    layer4_outputs(469) <= a;
    layer4_outputs(470) <= not a;
    layer4_outputs(471) <= b and not a;
    layer4_outputs(472) <= a;
    layer4_outputs(473) <= a;
    layer4_outputs(474) <= a and b;
    layer4_outputs(475) <= not (a or b);
    layer4_outputs(476) <= a xor b;
    layer4_outputs(477) <= not (a or b);
    layer4_outputs(478) <= b;
    layer4_outputs(479) <= 1'b1;
    layer4_outputs(480) <= b and not a;
    layer4_outputs(481) <= a or b;
    layer4_outputs(482) <= a xor b;
    layer4_outputs(483) <= not a or b;
    layer4_outputs(484) <= a;
    layer4_outputs(485) <= not a;
    layer4_outputs(486) <= a;
    layer4_outputs(487) <= not b;
    layer4_outputs(488) <= not (a xor b);
    layer4_outputs(489) <= a and not b;
    layer4_outputs(490) <= not (a and b);
    layer4_outputs(491) <= b;
    layer4_outputs(492) <= a and b;
    layer4_outputs(493) <= a;
    layer4_outputs(494) <= b;
    layer4_outputs(495) <= not b;
    layer4_outputs(496) <= b;
    layer4_outputs(497) <= not (a and b);
    layer4_outputs(498) <= not b or a;
    layer4_outputs(499) <= a;
    layer4_outputs(500) <= not a;
    layer4_outputs(501) <= b;
    layer4_outputs(502) <= not b or a;
    layer4_outputs(503) <= not b;
    layer4_outputs(504) <= not (a xor b);
    layer4_outputs(505) <= a or b;
    layer4_outputs(506) <= a;
    layer4_outputs(507) <= a and b;
    layer4_outputs(508) <= not a;
    layer4_outputs(509) <= a xor b;
    layer4_outputs(510) <= not a;
    layer4_outputs(511) <= not (a and b);
    layer4_outputs(512) <= not b or a;
    layer4_outputs(513) <= a xor b;
    layer4_outputs(514) <= not a or b;
    layer4_outputs(515) <= not a or b;
    layer4_outputs(516) <= not b;
    layer4_outputs(517) <= b;
    layer4_outputs(518) <= b;
    layer4_outputs(519) <= not a or b;
    layer4_outputs(520) <= not (a or b);
    layer4_outputs(521) <= not (a or b);
    layer4_outputs(522) <= b and not a;
    layer4_outputs(523) <= not (a or b);
    layer4_outputs(524) <= a and b;
    layer4_outputs(525) <= not a or b;
    layer4_outputs(526) <= not (a and b);
    layer4_outputs(527) <= not b;
    layer4_outputs(528) <= a and b;
    layer4_outputs(529) <= b and not a;
    layer4_outputs(530) <= not a;
    layer4_outputs(531) <= not (a and b);
    layer4_outputs(532) <= a;
    layer4_outputs(533) <= not b or a;
    layer4_outputs(534) <= not b;
    layer4_outputs(535) <= not (a and b);
    layer4_outputs(536) <= a or b;
    layer4_outputs(537) <= b;
    layer4_outputs(538) <= not b;
    layer4_outputs(539) <= a and not b;
    layer4_outputs(540) <= b;
    layer4_outputs(541) <= not (a and b);
    layer4_outputs(542) <= a or b;
    layer4_outputs(543) <= not a or b;
    layer4_outputs(544) <= b and not a;
    layer4_outputs(545) <= a;
    layer4_outputs(546) <= not a or b;
    layer4_outputs(547) <= not (a and b);
    layer4_outputs(548) <= not (a or b);
    layer4_outputs(549) <= a and not b;
    layer4_outputs(550) <= not (a or b);
    layer4_outputs(551) <= not (a and b);
    layer4_outputs(552) <= a;
    layer4_outputs(553) <= 1'b1;
    layer4_outputs(554) <= b and not a;
    layer4_outputs(555) <= a;
    layer4_outputs(556) <= b;
    layer4_outputs(557) <= a and b;
    layer4_outputs(558) <= not b;
    layer4_outputs(559) <= not a;
    layer4_outputs(560) <= b;
    layer4_outputs(561) <= a;
    layer4_outputs(562) <= a;
    layer4_outputs(563) <= not (a and b);
    layer4_outputs(564) <= not b;
    layer4_outputs(565) <= not b;
    layer4_outputs(566) <= not b;
    layer4_outputs(567) <= not b or a;
    layer4_outputs(568) <= a;
    layer4_outputs(569) <= b and not a;
    layer4_outputs(570) <= not a or b;
    layer4_outputs(571) <= not b or a;
    layer4_outputs(572) <= b;
    layer4_outputs(573) <= not a or b;
    layer4_outputs(574) <= a;
    layer4_outputs(575) <= not a;
    layer4_outputs(576) <= not a;
    layer4_outputs(577) <= not (a xor b);
    layer4_outputs(578) <= not b or a;
    layer4_outputs(579) <= b;
    layer4_outputs(580) <= b;
    layer4_outputs(581) <= a;
    layer4_outputs(582) <= not b;
    layer4_outputs(583) <= not b or a;
    layer4_outputs(584) <= not a or b;
    layer4_outputs(585) <= not b or a;
    layer4_outputs(586) <= a;
    layer4_outputs(587) <= not a or b;
    layer4_outputs(588) <= a or b;
    layer4_outputs(589) <= a or b;
    layer4_outputs(590) <= a or b;
    layer4_outputs(591) <= b and not a;
    layer4_outputs(592) <= not a;
    layer4_outputs(593) <= b;
    layer4_outputs(594) <= b;
    layer4_outputs(595) <= not (a or b);
    layer4_outputs(596) <= b;
    layer4_outputs(597) <= a;
    layer4_outputs(598) <= not b or a;
    layer4_outputs(599) <= not (a and b);
    layer4_outputs(600) <= a and not b;
    layer4_outputs(601) <= not b;
    layer4_outputs(602) <= b;
    layer4_outputs(603) <= not a or b;
    layer4_outputs(604) <= not b or a;
    layer4_outputs(605) <= b;
    layer4_outputs(606) <= not a;
    layer4_outputs(607) <= not a or b;
    layer4_outputs(608) <= b;
    layer4_outputs(609) <= a xor b;
    layer4_outputs(610) <= a xor b;
    layer4_outputs(611) <= a;
    layer4_outputs(612) <= not b;
    layer4_outputs(613) <= a;
    layer4_outputs(614) <= not (a or b);
    layer4_outputs(615) <= a and not b;
    layer4_outputs(616) <= not a;
    layer4_outputs(617) <= not (a xor b);
    layer4_outputs(618) <= not a;
    layer4_outputs(619) <= not b;
    layer4_outputs(620) <= a;
    layer4_outputs(621) <= b;
    layer4_outputs(622) <= a;
    layer4_outputs(623) <= not b;
    layer4_outputs(624) <= a and not b;
    layer4_outputs(625) <= a or b;
    layer4_outputs(626) <= a or b;
    layer4_outputs(627) <= not (a or b);
    layer4_outputs(628) <= not (a xor b);
    layer4_outputs(629) <= not b or a;
    layer4_outputs(630) <= b and not a;
    layer4_outputs(631) <= not (a or b);
    layer4_outputs(632) <= b;
    layer4_outputs(633) <= not b;
    layer4_outputs(634) <= b and not a;
    layer4_outputs(635) <= not a;
    layer4_outputs(636) <= not b;
    layer4_outputs(637) <= a or b;
    layer4_outputs(638) <= not b or a;
    layer4_outputs(639) <= not b or a;
    layer4_outputs(640) <= not a;
    layer4_outputs(641) <= not a;
    layer4_outputs(642) <= not a or b;
    layer4_outputs(643) <= b and not a;
    layer4_outputs(644) <= not b;
    layer4_outputs(645) <= not b;
    layer4_outputs(646) <= b;
    layer4_outputs(647) <= b;
    layer4_outputs(648) <= not (a and b);
    layer4_outputs(649) <= b;
    layer4_outputs(650) <= not b;
    layer4_outputs(651) <= a xor b;
    layer4_outputs(652) <= not a;
    layer4_outputs(653) <= not b;
    layer4_outputs(654) <= not b or a;
    layer4_outputs(655) <= not (a or b);
    layer4_outputs(656) <= a or b;
    layer4_outputs(657) <= not (a xor b);
    layer4_outputs(658) <= not b;
    layer4_outputs(659) <= 1'b1;
    layer4_outputs(660) <= not (a xor b);
    layer4_outputs(661) <= not (a and b);
    layer4_outputs(662) <= a and not b;
    layer4_outputs(663) <= not b or a;
    layer4_outputs(664) <= not b;
    layer4_outputs(665) <= not a;
    layer4_outputs(666) <= a xor b;
    layer4_outputs(667) <= not b;
    layer4_outputs(668) <= a xor b;
    layer4_outputs(669) <= not b;
    layer4_outputs(670) <= a or b;
    layer4_outputs(671) <= not a or b;
    layer4_outputs(672) <= not (a or b);
    layer4_outputs(673) <= not b or a;
    layer4_outputs(674) <= not a or b;
    layer4_outputs(675) <= not a;
    layer4_outputs(676) <= a and b;
    layer4_outputs(677) <= not a;
    layer4_outputs(678) <= a and not b;
    layer4_outputs(679) <= b and not a;
    layer4_outputs(680) <= b;
    layer4_outputs(681) <= not (a or b);
    layer4_outputs(682) <= not b;
    layer4_outputs(683) <= not b or a;
    layer4_outputs(684) <= a or b;
    layer4_outputs(685) <= not b or a;
    layer4_outputs(686) <= b and not a;
    layer4_outputs(687) <= not (a and b);
    layer4_outputs(688) <= a;
    layer4_outputs(689) <= a or b;
    layer4_outputs(690) <= a or b;
    layer4_outputs(691) <= a;
    layer4_outputs(692) <= b;
    layer4_outputs(693) <= not a;
    layer4_outputs(694) <= not a;
    layer4_outputs(695) <= a;
    layer4_outputs(696) <= a or b;
    layer4_outputs(697) <= not a or b;
    layer4_outputs(698) <= a and b;
    layer4_outputs(699) <= a;
    layer4_outputs(700) <= not (a and b);
    layer4_outputs(701) <= not a;
    layer4_outputs(702) <= a and b;
    layer4_outputs(703) <= a;
    layer4_outputs(704) <= not (a or b);
    layer4_outputs(705) <= a xor b;
    layer4_outputs(706) <= a and not b;
    layer4_outputs(707) <= not b;
    layer4_outputs(708) <= b and not a;
    layer4_outputs(709) <= not a;
    layer4_outputs(710) <= b;
    layer4_outputs(711) <= not b;
    layer4_outputs(712) <= a or b;
    layer4_outputs(713) <= a or b;
    layer4_outputs(714) <= a and b;
    layer4_outputs(715) <= a or b;
    layer4_outputs(716) <= a;
    layer4_outputs(717) <= 1'b1;
    layer4_outputs(718) <= b;
    layer4_outputs(719) <= b;
    layer4_outputs(720) <= not (a and b);
    layer4_outputs(721) <= not a or b;
    layer4_outputs(722) <= not (a or b);
    layer4_outputs(723) <= a and b;
    layer4_outputs(724) <= a;
    layer4_outputs(725) <= not b or a;
    layer4_outputs(726) <= a;
    layer4_outputs(727) <= a or b;
    layer4_outputs(728) <= not a or b;
    layer4_outputs(729) <= not b or a;
    layer4_outputs(730) <= not a or b;
    layer4_outputs(731) <= not (a xor b);
    layer4_outputs(732) <= not (a and b);
    layer4_outputs(733) <= not a or b;
    layer4_outputs(734) <= 1'b1;
    layer4_outputs(735) <= a or b;
    layer4_outputs(736) <= a or b;
    layer4_outputs(737) <= not (a and b);
    layer4_outputs(738) <= not a;
    layer4_outputs(739) <= not a;
    layer4_outputs(740) <= not a;
    layer4_outputs(741) <= not a;
    layer4_outputs(742) <= a xor b;
    layer4_outputs(743) <= a and b;
    layer4_outputs(744) <= not a;
    layer4_outputs(745) <= a;
    layer4_outputs(746) <= 1'b1;
    layer4_outputs(747) <= a xor b;
    layer4_outputs(748) <= a xor b;
    layer4_outputs(749) <= b;
    layer4_outputs(750) <= a;
    layer4_outputs(751) <= not a;
    layer4_outputs(752) <= not b;
    layer4_outputs(753) <= b;
    layer4_outputs(754) <= not b;
    layer4_outputs(755) <= a and b;
    layer4_outputs(756) <= a and not b;
    layer4_outputs(757) <= b;
    layer4_outputs(758) <= not b;
    layer4_outputs(759) <= a and b;
    layer4_outputs(760) <= not a;
    layer4_outputs(761) <= b;
    layer4_outputs(762) <= a and b;
    layer4_outputs(763) <= not a or b;
    layer4_outputs(764) <= a;
    layer4_outputs(765) <= not b;
    layer4_outputs(766) <= not b or a;
    layer4_outputs(767) <= not b;
    layer4_outputs(768) <= not b;
    layer4_outputs(769) <= 1'b0;
    layer4_outputs(770) <= not b or a;
    layer4_outputs(771) <= a and not b;
    layer4_outputs(772) <= not b;
    layer4_outputs(773) <= not b or a;
    layer4_outputs(774) <= not a;
    layer4_outputs(775) <= not (a and b);
    layer4_outputs(776) <= a and b;
    layer4_outputs(777) <= a xor b;
    layer4_outputs(778) <= b and not a;
    layer4_outputs(779) <= b;
    layer4_outputs(780) <= not a;
    layer4_outputs(781) <= not (a or b);
    layer4_outputs(782) <= not a or b;
    layer4_outputs(783) <= a;
    layer4_outputs(784) <= not (a and b);
    layer4_outputs(785) <= a;
    layer4_outputs(786) <= b and not a;
    layer4_outputs(787) <= not b or a;
    layer4_outputs(788) <= not a;
    layer4_outputs(789) <= not (a or b);
    layer4_outputs(790) <= a and b;
    layer4_outputs(791) <= a xor b;
    layer4_outputs(792) <= b;
    layer4_outputs(793) <= a and b;
    layer4_outputs(794) <= not (a xor b);
    layer4_outputs(795) <= not (a and b);
    layer4_outputs(796) <= not (a and b);
    layer4_outputs(797) <= b and not a;
    layer4_outputs(798) <= not b;
    layer4_outputs(799) <= b;
    layer4_outputs(800) <= not (a xor b);
    layer4_outputs(801) <= b and not a;
    layer4_outputs(802) <= b;
    layer4_outputs(803) <= not a;
    layer4_outputs(804) <= not a or b;
    layer4_outputs(805) <= a and b;
    layer4_outputs(806) <= not (a xor b);
    layer4_outputs(807) <= not b or a;
    layer4_outputs(808) <= a and not b;
    layer4_outputs(809) <= not a or b;
    layer4_outputs(810) <= b and not a;
    layer4_outputs(811) <= not a or b;
    layer4_outputs(812) <= not b;
    layer4_outputs(813) <= not (a or b);
    layer4_outputs(814) <= not (a or b);
    layer4_outputs(815) <= not a;
    layer4_outputs(816) <= a;
    layer4_outputs(817) <= a and not b;
    layer4_outputs(818) <= a;
    layer4_outputs(819) <= a;
    layer4_outputs(820) <= a;
    layer4_outputs(821) <= a;
    layer4_outputs(822) <= not a;
    layer4_outputs(823) <= not (a and b);
    layer4_outputs(824) <= a and b;
    layer4_outputs(825) <= not b;
    layer4_outputs(826) <= b and not a;
    layer4_outputs(827) <= a and not b;
    layer4_outputs(828) <= a;
    layer4_outputs(829) <= a and not b;
    layer4_outputs(830) <= a or b;
    layer4_outputs(831) <= b;
    layer4_outputs(832) <= not b or a;
    layer4_outputs(833) <= b;
    layer4_outputs(834) <= a or b;
    layer4_outputs(835) <= a xor b;
    layer4_outputs(836) <= not (a or b);
    layer4_outputs(837) <= b and not a;
    layer4_outputs(838) <= not b or a;
    layer4_outputs(839) <= not (a or b);
    layer4_outputs(840) <= a or b;
    layer4_outputs(841) <= b;
    layer4_outputs(842) <= a;
    layer4_outputs(843) <= not (a or b);
    layer4_outputs(844) <= a and b;
    layer4_outputs(845) <= a and not b;
    layer4_outputs(846) <= b;
    layer4_outputs(847) <= not b;
    layer4_outputs(848) <= b;
    layer4_outputs(849) <= b;
    layer4_outputs(850) <= not a or b;
    layer4_outputs(851) <= a;
    layer4_outputs(852) <= b;
    layer4_outputs(853) <= not b;
    layer4_outputs(854) <= not a;
    layer4_outputs(855) <= a;
    layer4_outputs(856) <= not (a and b);
    layer4_outputs(857) <= b and not a;
    layer4_outputs(858) <= a and b;
    layer4_outputs(859) <= b;
    layer4_outputs(860) <= a;
    layer4_outputs(861) <= not (a or b);
    layer4_outputs(862) <= a and not b;
    layer4_outputs(863) <= a and b;
    layer4_outputs(864) <= not a;
    layer4_outputs(865) <= b;
    layer4_outputs(866) <= not (a or b);
    layer4_outputs(867) <= not b or a;
    layer4_outputs(868) <= not (a or b);
    layer4_outputs(869) <= not (a and b);
    layer4_outputs(870) <= 1'b0;
    layer4_outputs(871) <= not a;
    layer4_outputs(872) <= not a;
    layer4_outputs(873) <= a;
    layer4_outputs(874) <= a or b;
    layer4_outputs(875) <= a xor b;
    layer4_outputs(876) <= not b;
    layer4_outputs(877) <= not a or b;
    layer4_outputs(878) <= not a or b;
    layer4_outputs(879) <= not b or a;
    layer4_outputs(880) <= b;
    layer4_outputs(881) <= a xor b;
    layer4_outputs(882) <= not (a or b);
    layer4_outputs(883) <= b;
    layer4_outputs(884) <= not b;
    layer4_outputs(885) <= b;
    layer4_outputs(886) <= b;
    layer4_outputs(887) <= not (a or b);
    layer4_outputs(888) <= a;
    layer4_outputs(889) <= not (a or b);
    layer4_outputs(890) <= not a;
    layer4_outputs(891) <= not (a or b);
    layer4_outputs(892) <= a and not b;
    layer4_outputs(893) <= a xor b;
    layer4_outputs(894) <= not a;
    layer4_outputs(895) <= not b or a;
    layer4_outputs(896) <= not a or b;
    layer4_outputs(897) <= a;
    layer4_outputs(898) <= not a or b;
    layer4_outputs(899) <= not a;
    layer4_outputs(900) <= a;
    layer4_outputs(901) <= a;
    layer4_outputs(902) <= not a;
    layer4_outputs(903) <= a;
    layer4_outputs(904) <= not a;
    layer4_outputs(905) <= a;
    layer4_outputs(906) <= not (a xor b);
    layer4_outputs(907) <= not (a or b);
    layer4_outputs(908) <= not a or b;
    layer4_outputs(909) <= a;
    layer4_outputs(910) <= not a or b;
    layer4_outputs(911) <= a or b;
    layer4_outputs(912) <= not a or b;
    layer4_outputs(913) <= not b;
    layer4_outputs(914) <= not b or a;
    layer4_outputs(915) <= not a;
    layer4_outputs(916) <= not (a xor b);
    layer4_outputs(917) <= a;
    layer4_outputs(918) <= not a or b;
    layer4_outputs(919) <= 1'b0;
    layer4_outputs(920) <= a and b;
    layer4_outputs(921) <= b;
    layer4_outputs(922) <= a;
    layer4_outputs(923) <= a and not b;
    layer4_outputs(924) <= not b or a;
    layer4_outputs(925) <= a and b;
    layer4_outputs(926) <= not b;
    layer4_outputs(927) <= not b;
    layer4_outputs(928) <= not a;
    layer4_outputs(929) <= not (a or b);
    layer4_outputs(930) <= not b;
    layer4_outputs(931) <= not (a or b);
    layer4_outputs(932) <= a and not b;
    layer4_outputs(933) <= not b;
    layer4_outputs(934) <= a;
    layer4_outputs(935) <= a or b;
    layer4_outputs(936) <= not b or a;
    layer4_outputs(937) <= not (a and b);
    layer4_outputs(938) <= not a or b;
    layer4_outputs(939) <= a;
    layer4_outputs(940) <= not a or b;
    layer4_outputs(941) <= not (a or b);
    layer4_outputs(942) <= a and not b;
    layer4_outputs(943) <= not (a xor b);
    layer4_outputs(944) <= not (a or b);
    layer4_outputs(945) <= a;
    layer4_outputs(946) <= a and not b;
    layer4_outputs(947) <= a;
    layer4_outputs(948) <= b;
    layer4_outputs(949) <= a or b;
    layer4_outputs(950) <= not a or b;
    layer4_outputs(951) <= b and not a;
    layer4_outputs(952) <= a and not b;
    layer4_outputs(953) <= not (a xor b);
    layer4_outputs(954) <= not (a or b);
    layer4_outputs(955) <= b;
    layer4_outputs(956) <= not (a and b);
    layer4_outputs(957) <= a and b;
    layer4_outputs(958) <= a;
    layer4_outputs(959) <= a and not b;
    layer4_outputs(960) <= b and not a;
    layer4_outputs(961) <= b and not a;
    layer4_outputs(962) <= not b;
    layer4_outputs(963) <= 1'b1;
    layer4_outputs(964) <= b and not a;
    layer4_outputs(965) <= a or b;
    layer4_outputs(966) <= not a;
    layer4_outputs(967) <= a and b;
    layer4_outputs(968) <= not (a and b);
    layer4_outputs(969) <= a or b;
    layer4_outputs(970) <= not a;
    layer4_outputs(971) <= not b or a;
    layer4_outputs(972) <= not (a xor b);
    layer4_outputs(973) <= not b;
    layer4_outputs(974) <= b;
    layer4_outputs(975) <= not b;
    layer4_outputs(976) <= a;
    layer4_outputs(977) <= not a;
    layer4_outputs(978) <= b and not a;
    layer4_outputs(979) <= not (a and b);
    layer4_outputs(980) <= not (a or b);
    layer4_outputs(981) <= not b or a;
    layer4_outputs(982) <= not a or b;
    layer4_outputs(983) <= not (a xor b);
    layer4_outputs(984) <= a and b;
    layer4_outputs(985) <= 1'b0;
    layer4_outputs(986) <= a and b;
    layer4_outputs(987) <= a;
    layer4_outputs(988) <= not a;
    layer4_outputs(989) <= a and not b;
    layer4_outputs(990) <= not a;
    layer4_outputs(991) <= a and b;
    layer4_outputs(992) <= a;
    layer4_outputs(993) <= b;
    layer4_outputs(994) <= b;
    layer4_outputs(995) <= not a;
    layer4_outputs(996) <= a xor b;
    layer4_outputs(997) <= a and not b;
    layer4_outputs(998) <= not a or b;
    layer4_outputs(999) <= not a or b;
    layer4_outputs(1000) <= not b;
    layer4_outputs(1001) <= a;
    layer4_outputs(1002) <= not (a or b);
    layer4_outputs(1003) <= b;
    layer4_outputs(1004) <= not (a and b);
    layer4_outputs(1005) <= b and not a;
    layer4_outputs(1006) <= a or b;
    layer4_outputs(1007) <= b and not a;
    layer4_outputs(1008) <= not a;
    layer4_outputs(1009) <= not b or a;
    layer4_outputs(1010) <= not b;
    layer4_outputs(1011) <= not a or b;
    layer4_outputs(1012) <= not a;
    layer4_outputs(1013) <= b and not a;
    layer4_outputs(1014) <= not a or b;
    layer4_outputs(1015) <= b;
    layer4_outputs(1016) <= not (a xor b);
    layer4_outputs(1017) <= a or b;
    layer4_outputs(1018) <= b;
    layer4_outputs(1019) <= b;
    layer4_outputs(1020) <= 1'b0;
    layer4_outputs(1021) <= a xor b;
    layer4_outputs(1022) <= a;
    layer4_outputs(1023) <= a xor b;
    layer4_outputs(1024) <= not b or a;
    layer4_outputs(1025) <= b and not a;
    layer4_outputs(1026) <= not b or a;
    layer4_outputs(1027) <= not (a and b);
    layer4_outputs(1028) <= b;
    layer4_outputs(1029) <= a or b;
    layer4_outputs(1030) <= b and not a;
    layer4_outputs(1031) <= a and b;
    layer4_outputs(1032) <= a and b;
    layer4_outputs(1033) <= a and b;
    layer4_outputs(1034) <= not a;
    layer4_outputs(1035) <= not b;
    layer4_outputs(1036) <= not (a or b);
    layer4_outputs(1037) <= not (a or b);
    layer4_outputs(1038) <= not a or b;
    layer4_outputs(1039) <= a xor b;
    layer4_outputs(1040) <= not (a and b);
    layer4_outputs(1041) <= b;
    layer4_outputs(1042) <= not a;
    layer4_outputs(1043) <= not (a and b);
    layer4_outputs(1044) <= b;
    layer4_outputs(1045) <= b;
    layer4_outputs(1046) <= b and not a;
    layer4_outputs(1047) <= not b or a;
    layer4_outputs(1048) <= not (a xor b);
    layer4_outputs(1049) <= not a or b;
    layer4_outputs(1050) <= not b;
    layer4_outputs(1051) <= a;
    layer4_outputs(1052) <= a;
    layer4_outputs(1053) <= not a or b;
    layer4_outputs(1054) <= b;
    layer4_outputs(1055) <= a;
    layer4_outputs(1056) <= a;
    layer4_outputs(1057) <= b and not a;
    layer4_outputs(1058) <= 1'b0;
    layer4_outputs(1059) <= a;
    layer4_outputs(1060) <= a or b;
    layer4_outputs(1061) <= b and not a;
    layer4_outputs(1062) <= not a;
    layer4_outputs(1063) <= a or b;
    layer4_outputs(1064) <= not a or b;
    layer4_outputs(1065) <= not a or b;
    layer4_outputs(1066) <= not a;
    layer4_outputs(1067) <= not (a or b);
    layer4_outputs(1068) <= not (a or b);
    layer4_outputs(1069) <= not a;
    layer4_outputs(1070) <= a;
    layer4_outputs(1071) <= not b or a;
    layer4_outputs(1072) <= b;
    layer4_outputs(1073) <= not (a xor b);
    layer4_outputs(1074) <= not a or b;
    layer4_outputs(1075) <= b;
    layer4_outputs(1076) <= not (a or b);
    layer4_outputs(1077) <= b and not a;
    layer4_outputs(1078) <= b;
    layer4_outputs(1079) <= b;
    layer4_outputs(1080) <= b;
    layer4_outputs(1081) <= a xor b;
    layer4_outputs(1082) <= not (a xor b);
    layer4_outputs(1083) <= a and b;
    layer4_outputs(1084) <= not b or a;
    layer4_outputs(1085) <= not b or a;
    layer4_outputs(1086) <= 1'b1;
    layer4_outputs(1087) <= b;
    layer4_outputs(1088) <= b;
    layer4_outputs(1089) <= b;
    layer4_outputs(1090) <= not (a and b);
    layer4_outputs(1091) <= b;
    layer4_outputs(1092) <= a;
    layer4_outputs(1093) <= not a or b;
    layer4_outputs(1094) <= not b;
    layer4_outputs(1095) <= not a;
    layer4_outputs(1096) <= not a;
    layer4_outputs(1097) <= not a or b;
    layer4_outputs(1098) <= not (a or b);
    layer4_outputs(1099) <= a and not b;
    layer4_outputs(1100) <= not a;
    layer4_outputs(1101) <= not b;
    layer4_outputs(1102) <= not a;
    layer4_outputs(1103) <= not (a or b);
    layer4_outputs(1104) <= not (a xor b);
    layer4_outputs(1105) <= a or b;
    layer4_outputs(1106) <= a and b;
    layer4_outputs(1107) <= a and b;
    layer4_outputs(1108) <= not b or a;
    layer4_outputs(1109) <= a or b;
    layer4_outputs(1110) <= not (a and b);
    layer4_outputs(1111) <= not a;
    layer4_outputs(1112) <= a;
    layer4_outputs(1113) <= not a;
    layer4_outputs(1114) <= b and not a;
    layer4_outputs(1115) <= not b;
    layer4_outputs(1116) <= not a or b;
    layer4_outputs(1117) <= a;
    layer4_outputs(1118) <= not b;
    layer4_outputs(1119) <= b;
    layer4_outputs(1120) <= b;
    layer4_outputs(1121) <= not a;
    layer4_outputs(1122) <= b;
    layer4_outputs(1123) <= a and not b;
    layer4_outputs(1124) <= not b;
    layer4_outputs(1125) <= not b;
    layer4_outputs(1126) <= b;
    layer4_outputs(1127) <= a and b;
    layer4_outputs(1128) <= b and not a;
    layer4_outputs(1129) <= not a;
    layer4_outputs(1130) <= b and not a;
    layer4_outputs(1131) <= not a;
    layer4_outputs(1132) <= b;
    layer4_outputs(1133) <= b;
    layer4_outputs(1134) <= b;
    layer4_outputs(1135) <= 1'b1;
    layer4_outputs(1136) <= a;
    layer4_outputs(1137) <= a or b;
    layer4_outputs(1138) <= not b;
    layer4_outputs(1139) <= not a;
    layer4_outputs(1140) <= 1'b0;
    layer4_outputs(1141) <= not (a or b);
    layer4_outputs(1142) <= not (a and b);
    layer4_outputs(1143) <= a;
    layer4_outputs(1144) <= a;
    layer4_outputs(1145) <= b;
    layer4_outputs(1146) <= a and b;
    layer4_outputs(1147) <= b and not a;
    layer4_outputs(1148) <= not a;
    layer4_outputs(1149) <= not (a and b);
    layer4_outputs(1150) <= not b;
    layer4_outputs(1151) <= a;
    layer4_outputs(1152) <= not b or a;
    layer4_outputs(1153) <= not (a and b);
    layer4_outputs(1154) <= b and not a;
    layer4_outputs(1155) <= a and not b;
    layer4_outputs(1156) <= not a;
    layer4_outputs(1157) <= b and not a;
    layer4_outputs(1158) <= a xor b;
    layer4_outputs(1159) <= a;
    layer4_outputs(1160) <= not b;
    layer4_outputs(1161) <= not b;
    layer4_outputs(1162) <= a xor b;
    layer4_outputs(1163) <= not b or a;
    layer4_outputs(1164) <= not a;
    layer4_outputs(1165) <= not a or b;
    layer4_outputs(1166) <= a xor b;
    layer4_outputs(1167) <= not (a or b);
    layer4_outputs(1168) <= a;
    layer4_outputs(1169) <= a;
    layer4_outputs(1170) <= not (a and b);
    layer4_outputs(1171) <= not a;
    layer4_outputs(1172) <= not (a or b);
    layer4_outputs(1173) <= a or b;
    layer4_outputs(1174) <= a and b;
    layer4_outputs(1175) <= a;
    layer4_outputs(1176) <= a xor b;
    layer4_outputs(1177) <= not (a or b);
    layer4_outputs(1178) <= not a or b;
    layer4_outputs(1179) <= not (a xor b);
    layer4_outputs(1180) <= not a;
    layer4_outputs(1181) <= not b or a;
    layer4_outputs(1182) <= not b;
    layer4_outputs(1183) <= not a or b;
    layer4_outputs(1184) <= not b;
    layer4_outputs(1185) <= a and not b;
    layer4_outputs(1186) <= not b;
    layer4_outputs(1187) <= not b;
    layer4_outputs(1188) <= not b;
    layer4_outputs(1189) <= a;
    layer4_outputs(1190) <= b;
    layer4_outputs(1191) <= not b;
    layer4_outputs(1192) <= not (a and b);
    layer4_outputs(1193) <= not a;
    layer4_outputs(1194) <= not a or b;
    layer4_outputs(1195) <= a and not b;
    layer4_outputs(1196) <= not a;
    layer4_outputs(1197) <= a or b;
    layer4_outputs(1198) <= not b;
    layer4_outputs(1199) <= a xor b;
    layer4_outputs(1200) <= a and not b;
    layer4_outputs(1201) <= a and b;
    layer4_outputs(1202) <= not a;
    layer4_outputs(1203) <= a and b;
    layer4_outputs(1204) <= a;
    layer4_outputs(1205) <= not b or a;
    layer4_outputs(1206) <= not a;
    layer4_outputs(1207) <= b;
    layer4_outputs(1208) <= not (a xor b);
    layer4_outputs(1209) <= a and b;
    layer4_outputs(1210) <= a or b;
    layer4_outputs(1211) <= b and not a;
    layer4_outputs(1212) <= not (a xor b);
    layer4_outputs(1213) <= a;
    layer4_outputs(1214) <= not b or a;
    layer4_outputs(1215) <= b;
    layer4_outputs(1216) <= not (a or b);
    layer4_outputs(1217) <= a or b;
    layer4_outputs(1218) <= 1'b1;
    layer4_outputs(1219) <= b and not a;
    layer4_outputs(1220) <= a and not b;
    layer4_outputs(1221) <= b and not a;
    layer4_outputs(1222) <= not (a xor b);
    layer4_outputs(1223) <= a and b;
    layer4_outputs(1224) <= not (a and b);
    layer4_outputs(1225) <= a and b;
    layer4_outputs(1226) <= not b or a;
    layer4_outputs(1227) <= not (a and b);
    layer4_outputs(1228) <= a xor b;
    layer4_outputs(1229) <= a;
    layer4_outputs(1230) <= a;
    layer4_outputs(1231) <= not (a or b);
    layer4_outputs(1232) <= b and not a;
    layer4_outputs(1233) <= a and not b;
    layer4_outputs(1234) <= a or b;
    layer4_outputs(1235) <= not a;
    layer4_outputs(1236) <= b;
    layer4_outputs(1237) <= not (a or b);
    layer4_outputs(1238) <= a and b;
    layer4_outputs(1239) <= a or b;
    layer4_outputs(1240) <= a;
    layer4_outputs(1241) <= b and not a;
    layer4_outputs(1242) <= not b;
    layer4_outputs(1243) <= a and b;
    layer4_outputs(1244) <= not a;
    layer4_outputs(1245) <= not (a xor b);
    layer4_outputs(1246) <= not a;
    layer4_outputs(1247) <= not b;
    layer4_outputs(1248) <= not a or b;
    layer4_outputs(1249) <= not (a and b);
    layer4_outputs(1250) <= a and b;
    layer4_outputs(1251) <= not a or b;
    layer4_outputs(1252) <= not a or b;
    layer4_outputs(1253) <= not b or a;
    layer4_outputs(1254) <= a;
    layer4_outputs(1255) <= b and not a;
    layer4_outputs(1256) <= not a;
    layer4_outputs(1257) <= not a or b;
    layer4_outputs(1258) <= not b;
    layer4_outputs(1259) <= not b;
    layer4_outputs(1260) <= a xor b;
    layer4_outputs(1261) <= not b;
    layer4_outputs(1262) <= b;
    layer4_outputs(1263) <= a and not b;
    layer4_outputs(1264) <= not (a and b);
    layer4_outputs(1265) <= not a or b;
    layer4_outputs(1266) <= b and not a;
    layer4_outputs(1267) <= not b or a;
    layer4_outputs(1268) <= not a;
    layer4_outputs(1269) <= not a;
    layer4_outputs(1270) <= not b or a;
    layer4_outputs(1271) <= not a;
    layer4_outputs(1272) <= not b;
    layer4_outputs(1273) <= b;
    layer4_outputs(1274) <= a or b;
    layer4_outputs(1275) <= not a;
    layer4_outputs(1276) <= a or b;
    layer4_outputs(1277) <= a and b;
    layer4_outputs(1278) <= not (a and b);
    layer4_outputs(1279) <= not a or b;
    layer4_outputs(1280) <= not a or b;
    layer4_outputs(1281) <= a and not b;
    layer4_outputs(1282) <= not a or b;
    layer4_outputs(1283) <= a and not b;
    layer4_outputs(1284) <= not b;
    layer4_outputs(1285) <= not b;
    layer4_outputs(1286) <= b;
    layer4_outputs(1287) <= a or b;
    layer4_outputs(1288) <= b and not a;
    layer4_outputs(1289) <= not (a and b);
    layer4_outputs(1290) <= a and b;
    layer4_outputs(1291) <= b;
    layer4_outputs(1292) <= a and not b;
    layer4_outputs(1293) <= a and not b;
    layer4_outputs(1294) <= a or b;
    layer4_outputs(1295) <= not (a xor b);
    layer4_outputs(1296) <= not a;
    layer4_outputs(1297) <= not a;
    layer4_outputs(1298) <= not a;
    layer4_outputs(1299) <= not a;
    layer4_outputs(1300) <= b;
    layer4_outputs(1301) <= a and b;
    layer4_outputs(1302) <= 1'b1;
    layer4_outputs(1303) <= b;
    layer4_outputs(1304) <= a and not b;
    layer4_outputs(1305) <= b;
    layer4_outputs(1306) <= not (a and b);
    layer4_outputs(1307) <= a and b;
    layer4_outputs(1308) <= a;
    layer4_outputs(1309) <= a or b;
    layer4_outputs(1310) <= not b;
    layer4_outputs(1311) <= not b or a;
    layer4_outputs(1312) <= not b or a;
    layer4_outputs(1313) <= not a;
    layer4_outputs(1314) <= not (a and b);
    layer4_outputs(1315) <= a;
    layer4_outputs(1316) <= not b;
    layer4_outputs(1317) <= not (a xor b);
    layer4_outputs(1318) <= a;
    layer4_outputs(1319) <= 1'b1;
    layer4_outputs(1320) <= a and not b;
    layer4_outputs(1321) <= not b;
    layer4_outputs(1322) <= not b or a;
    layer4_outputs(1323) <= not a;
    layer4_outputs(1324) <= not (a and b);
    layer4_outputs(1325) <= a;
    layer4_outputs(1326) <= not b or a;
    layer4_outputs(1327) <= not (a xor b);
    layer4_outputs(1328) <= a and b;
    layer4_outputs(1329) <= a;
    layer4_outputs(1330) <= a;
    layer4_outputs(1331) <= not (a and b);
    layer4_outputs(1332) <= not a;
    layer4_outputs(1333) <= not b;
    layer4_outputs(1334) <= a or b;
    layer4_outputs(1335) <= a;
    layer4_outputs(1336) <= not (a xor b);
    layer4_outputs(1337) <= a and b;
    layer4_outputs(1338) <= not b;
    layer4_outputs(1339) <= not b or a;
    layer4_outputs(1340) <= not b;
    layer4_outputs(1341) <= b and not a;
    layer4_outputs(1342) <= not (a and b);
    layer4_outputs(1343) <= a;
    layer4_outputs(1344) <= a;
    layer4_outputs(1345) <= not a or b;
    layer4_outputs(1346) <= not b or a;
    layer4_outputs(1347) <= not a;
    layer4_outputs(1348) <= b;
    layer4_outputs(1349) <= a;
    layer4_outputs(1350) <= not b;
    layer4_outputs(1351) <= b;
    layer4_outputs(1352) <= not (a or b);
    layer4_outputs(1353) <= a or b;
    layer4_outputs(1354) <= not (a and b);
    layer4_outputs(1355) <= not a;
    layer4_outputs(1356) <= a or b;
    layer4_outputs(1357) <= a or b;
    layer4_outputs(1358) <= b and not a;
    layer4_outputs(1359) <= a or b;
    layer4_outputs(1360) <= b and not a;
    layer4_outputs(1361) <= not a or b;
    layer4_outputs(1362) <= not (a and b);
    layer4_outputs(1363) <= b;
    layer4_outputs(1364) <= a xor b;
    layer4_outputs(1365) <= not a or b;
    layer4_outputs(1366) <= a;
    layer4_outputs(1367) <= not b;
    layer4_outputs(1368) <= a and b;
    layer4_outputs(1369) <= not a;
    layer4_outputs(1370) <= not a;
    layer4_outputs(1371) <= not (a or b);
    layer4_outputs(1372) <= a;
    layer4_outputs(1373) <= not (a or b);
    layer4_outputs(1374) <= not a or b;
    layer4_outputs(1375) <= a xor b;
    layer4_outputs(1376) <= not b;
    layer4_outputs(1377) <= a or b;
    layer4_outputs(1378) <= not (a xor b);
    layer4_outputs(1379) <= not b;
    layer4_outputs(1380) <= a;
    layer4_outputs(1381) <= not (a and b);
    layer4_outputs(1382) <= a;
    layer4_outputs(1383) <= a xor b;
    layer4_outputs(1384) <= not b;
    layer4_outputs(1385) <= 1'b0;
    layer4_outputs(1386) <= b and not a;
    layer4_outputs(1387) <= not a or b;
    layer4_outputs(1388) <= not a;
    layer4_outputs(1389) <= a;
    layer4_outputs(1390) <= not a;
    layer4_outputs(1391) <= a and not b;
    layer4_outputs(1392) <= not (a or b);
    layer4_outputs(1393) <= not a or b;
    layer4_outputs(1394) <= not (a and b);
    layer4_outputs(1395) <= not (a xor b);
    layer4_outputs(1396) <= not a;
    layer4_outputs(1397) <= not a;
    layer4_outputs(1398) <= not b or a;
    layer4_outputs(1399) <= not b;
    layer4_outputs(1400) <= a and not b;
    layer4_outputs(1401) <= a;
    layer4_outputs(1402) <= not b;
    layer4_outputs(1403) <= b;
    layer4_outputs(1404) <= not (a xor b);
    layer4_outputs(1405) <= not a;
    layer4_outputs(1406) <= not a;
    layer4_outputs(1407) <= a;
    layer4_outputs(1408) <= 1'b1;
    layer4_outputs(1409) <= not (a and b);
    layer4_outputs(1410) <= a and not b;
    layer4_outputs(1411) <= a;
    layer4_outputs(1412) <= not a;
    layer4_outputs(1413) <= b and not a;
    layer4_outputs(1414) <= not (a and b);
    layer4_outputs(1415) <= a;
    layer4_outputs(1416) <= a and not b;
    layer4_outputs(1417) <= not b;
    layer4_outputs(1418) <= not b;
    layer4_outputs(1419) <= not b;
    layer4_outputs(1420) <= a xor b;
    layer4_outputs(1421) <= not (a or b);
    layer4_outputs(1422) <= not (a and b);
    layer4_outputs(1423) <= not (a and b);
    layer4_outputs(1424) <= 1'b0;
    layer4_outputs(1425) <= not b;
    layer4_outputs(1426) <= a and b;
    layer4_outputs(1427) <= not a;
    layer4_outputs(1428) <= b and not a;
    layer4_outputs(1429) <= a or b;
    layer4_outputs(1430) <= not b;
    layer4_outputs(1431) <= a xor b;
    layer4_outputs(1432) <= b and not a;
    layer4_outputs(1433) <= a;
    layer4_outputs(1434) <= a xor b;
    layer4_outputs(1435) <= a and b;
    layer4_outputs(1436) <= not b;
    layer4_outputs(1437) <= a xor b;
    layer4_outputs(1438) <= a and not b;
    layer4_outputs(1439) <= not (a or b);
    layer4_outputs(1440) <= not (a or b);
    layer4_outputs(1441) <= a;
    layer4_outputs(1442) <= not (a xor b);
    layer4_outputs(1443) <= not b;
    layer4_outputs(1444) <= not (a or b);
    layer4_outputs(1445) <= not (a and b);
    layer4_outputs(1446) <= b and not a;
    layer4_outputs(1447) <= a;
    layer4_outputs(1448) <= b and not a;
    layer4_outputs(1449) <= a or b;
    layer4_outputs(1450) <= not (a and b);
    layer4_outputs(1451) <= a and not b;
    layer4_outputs(1452) <= not (a and b);
    layer4_outputs(1453) <= not b;
    layer4_outputs(1454) <= not (a and b);
    layer4_outputs(1455) <= a and b;
    layer4_outputs(1456) <= a and not b;
    layer4_outputs(1457) <= not a;
    layer4_outputs(1458) <= a;
    layer4_outputs(1459) <= a and b;
    layer4_outputs(1460) <= not a;
    layer4_outputs(1461) <= a;
    layer4_outputs(1462) <= b;
    layer4_outputs(1463) <= not a;
    layer4_outputs(1464) <= a and b;
    layer4_outputs(1465) <= not b or a;
    layer4_outputs(1466) <= b;
    layer4_outputs(1467) <= not b;
    layer4_outputs(1468) <= b;
    layer4_outputs(1469) <= not a;
    layer4_outputs(1470) <= not (a and b);
    layer4_outputs(1471) <= b and not a;
    layer4_outputs(1472) <= not (a xor b);
    layer4_outputs(1473) <= not a;
    layer4_outputs(1474) <= not a or b;
    layer4_outputs(1475) <= a or b;
    layer4_outputs(1476) <= not a;
    layer4_outputs(1477) <= 1'b0;
    layer4_outputs(1478) <= not a;
    layer4_outputs(1479) <= not b;
    layer4_outputs(1480) <= a or b;
    layer4_outputs(1481) <= not a;
    layer4_outputs(1482) <= b;
    layer4_outputs(1483) <= not a;
    layer4_outputs(1484) <= not b or a;
    layer4_outputs(1485) <= not a;
    layer4_outputs(1486) <= 1'b0;
    layer4_outputs(1487) <= not (a and b);
    layer4_outputs(1488) <= a and b;
    layer4_outputs(1489) <= not a or b;
    layer4_outputs(1490) <= b and not a;
    layer4_outputs(1491) <= not a or b;
    layer4_outputs(1492) <= a and b;
    layer4_outputs(1493) <= not a;
    layer4_outputs(1494) <= not b;
    layer4_outputs(1495) <= not b or a;
    layer4_outputs(1496) <= not a or b;
    layer4_outputs(1497) <= not a;
    layer4_outputs(1498) <= b;
    layer4_outputs(1499) <= not b;
    layer4_outputs(1500) <= b;
    layer4_outputs(1501) <= a;
    layer4_outputs(1502) <= b;
    layer4_outputs(1503) <= b;
    layer4_outputs(1504) <= a;
    layer4_outputs(1505) <= a or b;
    layer4_outputs(1506) <= not a or b;
    layer4_outputs(1507) <= not (a or b);
    layer4_outputs(1508) <= not (a or b);
    layer4_outputs(1509) <= a xor b;
    layer4_outputs(1510) <= b;
    layer4_outputs(1511) <= a and not b;
    layer4_outputs(1512) <= not b or a;
    layer4_outputs(1513) <= a;
    layer4_outputs(1514) <= b;
    layer4_outputs(1515) <= not a or b;
    layer4_outputs(1516) <= a;
    layer4_outputs(1517) <= a or b;
    layer4_outputs(1518) <= a;
    layer4_outputs(1519) <= a and not b;
    layer4_outputs(1520) <= a;
    layer4_outputs(1521) <= not a;
    layer4_outputs(1522) <= not b;
    layer4_outputs(1523) <= not a;
    layer4_outputs(1524) <= b and not a;
    layer4_outputs(1525) <= a and b;
    layer4_outputs(1526) <= not (a or b);
    layer4_outputs(1527) <= not a or b;
    layer4_outputs(1528) <= not b or a;
    layer4_outputs(1529) <= not (a and b);
    layer4_outputs(1530) <= b;
    layer4_outputs(1531) <= 1'b0;
    layer4_outputs(1532) <= not (a and b);
    layer4_outputs(1533) <= not b;
    layer4_outputs(1534) <= b;
    layer4_outputs(1535) <= not b;
    layer4_outputs(1536) <= a and not b;
    layer4_outputs(1537) <= not (a xor b);
    layer4_outputs(1538) <= b and not a;
    layer4_outputs(1539) <= not (a xor b);
    layer4_outputs(1540) <= not (a or b);
    layer4_outputs(1541) <= b and not a;
    layer4_outputs(1542) <= a and not b;
    layer4_outputs(1543) <= a or b;
    layer4_outputs(1544) <= not (a and b);
    layer4_outputs(1545) <= a and b;
    layer4_outputs(1546) <= b;
    layer4_outputs(1547) <= not b;
    layer4_outputs(1548) <= b;
    layer4_outputs(1549) <= a;
    layer4_outputs(1550) <= not a or b;
    layer4_outputs(1551) <= b and not a;
    layer4_outputs(1552) <= not b;
    layer4_outputs(1553) <= b and not a;
    layer4_outputs(1554) <= not a;
    layer4_outputs(1555) <= not a;
    layer4_outputs(1556) <= not a;
    layer4_outputs(1557) <= b and not a;
    layer4_outputs(1558) <= a;
    layer4_outputs(1559) <= a or b;
    layer4_outputs(1560) <= a and b;
    layer4_outputs(1561) <= not (a and b);
    layer4_outputs(1562) <= a and b;
    layer4_outputs(1563) <= not b or a;
    layer4_outputs(1564) <= not a or b;
    layer4_outputs(1565) <= not (a and b);
    layer4_outputs(1566) <= not b;
    layer4_outputs(1567) <= a xor b;
    layer4_outputs(1568) <= a and not b;
    layer4_outputs(1569) <= b;
    layer4_outputs(1570) <= a and not b;
    layer4_outputs(1571) <= a or b;
    layer4_outputs(1572) <= not (a or b);
    layer4_outputs(1573) <= not a;
    layer4_outputs(1574) <= b;
    layer4_outputs(1575) <= b;
    layer4_outputs(1576) <= a;
    layer4_outputs(1577) <= a xor b;
    layer4_outputs(1578) <= 1'b0;
    layer4_outputs(1579) <= b;
    layer4_outputs(1580) <= a xor b;
    layer4_outputs(1581) <= a and b;
    layer4_outputs(1582) <= not b;
    layer4_outputs(1583) <= a;
    layer4_outputs(1584) <= not a or b;
    layer4_outputs(1585) <= not b or a;
    layer4_outputs(1586) <= not a or b;
    layer4_outputs(1587) <= b and not a;
    layer4_outputs(1588) <= not a or b;
    layer4_outputs(1589) <= a and b;
    layer4_outputs(1590) <= b;
    layer4_outputs(1591) <= not (a and b);
    layer4_outputs(1592) <= a and not b;
    layer4_outputs(1593) <= not a or b;
    layer4_outputs(1594) <= not b or a;
    layer4_outputs(1595) <= a;
    layer4_outputs(1596) <= b and not a;
    layer4_outputs(1597) <= not b or a;
    layer4_outputs(1598) <= b and not a;
    layer4_outputs(1599) <= a;
    layer4_outputs(1600) <= b and not a;
    layer4_outputs(1601) <= a;
    layer4_outputs(1602) <= a;
    layer4_outputs(1603) <= not b or a;
    layer4_outputs(1604) <= not b;
    layer4_outputs(1605) <= not b;
    layer4_outputs(1606) <= not (a and b);
    layer4_outputs(1607) <= not a;
    layer4_outputs(1608) <= a or b;
    layer4_outputs(1609) <= not b;
    layer4_outputs(1610) <= a and b;
    layer4_outputs(1611) <= b and not a;
    layer4_outputs(1612) <= b;
    layer4_outputs(1613) <= not a or b;
    layer4_outputs(1614) <= a or b;
    layer4_outputs(1615) <= not b or a;
    layer4_outputs(1616) <= not b;
    layer4_outputs(1617) <= a;
    layer4_outputs(1618) <= a;
    layer4_outputs(1619) <= b and not a;
    layer4_outputs(1620) <= a xor b;
    layer4_outputs(1621) <= not (a or b);
    layer4_outputs(1622) <= a xor b;
    layer4_outputs(1623) <= b;
    layer4_outputs(1624) <= b;
    layer4_outputs(1625) <= not a;
    layer4_outputs(1626) <= not (a and b);
    layer4_outputs(1627) <= a or b;
    layer4_outputs(1628) <= not (a or b);
    layer4_outputs(1629) <= b and not a;
    layer4_outputs(1630) <= not (a and b);
    layer4_outputs(1631) <= b and not a;
    layer4_outputs(1632) <= a;
    layer4_outputs(1633) <= b;
    layer4_outputs(1634) <= not (a xor b);
    layer4_outputs(1635) <= not b;
    layer4_outputs(1636) <= not (a or b);
    layer4_outputs(1637) <= a or b;
    layer4_outputs(1638) <= b and not a;
    layer4_outputs(1639) <= not (a and b);
    layer4_outputs(1640) <= a and b;
    layer4_outputs(1641) <= b;
    layer4_outputs(1642) <= not a;
    layer4_outputs(1643) <= a or b;
    layer4_outputs(1644) <= not b;
    layer4_outputs(1645) <= not a or b;
    layer4_outputs(1646) <= not a;
    layer4_outputs(1647) <= a;
    layer4_outputs(1648) <= b;
    layer4_outputs(1649) <= not (a and b);
    layer4_outputs(1650) <= 1'b0;
    layer4_outputs(1651) <= a;
    layer4_outputs(1652) <= b;
    layer4_outputs(1653) <= b;
    layer4_outputs(1654) <= not a or b;
    layer4_outputs(1655) <= not (a and b);
    layer4_outputs(1656) <= not (a and b);
    layer4_outputs(1657) <= b and not a;
    layer4_outputs(1658) <= b and not a;
    layer4_outputs(1659) <= not a;
    layer4_outputs(1660) <= a;
    layer4_outputs(1661) <= a and not b;
    layer4_outputs(1662) <= not b;
    layer4_outputs(1663) <= not (a and b);
    layer4_outputs(1664) <= not (a xor b);
    layer4_outputs(1665) <= not b;
    layer4_outputs(1666) <= b and not a;
    layer4_outputs(1667) <= 1'b0;
    layer4_outputs(1668) <= not b;
    layer4_outputs(1669) <= b;
    layer4_outputs(1670) <= not b;
    layer4_outputs(1671) <= b and not a;
    layer4_outputs(1672) <= not a;
    layer4_outputs(1673) <= not b;
    layer4_outputs(1674) <= a xor b;
    layer4_outputs(1675) <= not b or a;
    layer4_outputs(1676) <= a or b;
    layer4_outputs(1677) <= not b;
    layer4_outputs(1678) <= not (a or b);
    layer4_outputs(1679) <= b;
    layer4_outputs(1680) <= not a or b;
    layer4_outputs(1681) <= a or b;
    layer4_outputs(1682) <= not a;
    layer4_outputs(1683) <= a and not b;
    layer4_outputs(1684) <= a or b;
    layer4_outputs(1685) <= not a;
    layer4_outputs(1686) <= a;
    layer4_outputs(1687) <= a and not b;
    layer4_outputs(1688) <= b and not a;
    layer4_outputs(1689) <= not (a or b);
    layer4_outputs(1690) <= not a;
    layer4_outputs(1691) <= not (a or b);
    layer4_outputs(1692) <= not a;
    layer4_outputs(1693) <= a xor b;
    layer4_outputs(1694) <= a;
    layer4_outputs(1695) <= not b;
    layer4_outputs(1696) <= not b;
    layer4_outputs(1697) <= b;
    layer4_outputs(1698) <= 1'b0;
    layer4_outputs(1699) <= not b;
    layer4_outputs(1700) <= a;
    layer4_outputs(1701) <= b;
    layer4_outputs(1702) <= a;
    layer4_outputs(1703) <= b;
    layer4_outputs(1704) <= not a;
    layer4_outputs(1705) <= not a;
    layer4_outputs(1706) <= not a;
    layer4_outputs(1707) <= not b or a;
    layer4_outputs(1708) <= not a or b;
    layer4_outputs(1709) <= 1'b0;
    layer4_outputs(1710) <= not (a and b);
    layer4_outputs(1711) <= not b;
    layer4_outputs(1712) <= not b;
    layer4_outputs(1713) <= not (a and b);
    layer4_outputs(1714) <= not a or b;
    layer4_outputs(1715) <= not b;
    layer4_outputs(1716) <= not a or b;
    layer4_outputs(1717) <= a and b;
    layer4_outputs(1718) <= a and b;
    layer4_outputs(1719) <= a or b;
    layer4_outputs(1720) <= a;
    layer4_outputs(1721) <= b;
    layer4_outputs(1722) <= a;
    layer4_outputs(1723) <= b;
    layer4_outputs(1724) <= not b;
    layer4_outputs(1725) <= not b;
    layer4_outputs(1726) <= 1'b1;
    layer4_outputs(1727) <= 1'b0;
    layer4_outputs(1728) <= a;
    layer4_outputs(1729) <= b and not a;
    layer4_outputs(1730) <= b;
    layer4_outputs(1731) <= not b;
    layer4_outputs(1732) <= not b or a;
    layer4_outputs(1733) <= a and not b;
    layer4_outputs(1734) <= not (a or b);
    layer4_outputs(1735) <= not (a or b);
    layer4_outputs(1736) <= not (a xor b);
    layer4_outputs(1737) <= not (a and b);
    layer4_outputs(1738) <= b and not a;
    layer4_outputs(1739) <= not b;
    layer4_outputs(1740) <= not (a or b);
    layer4_outputs(1741) <= not b or a;
    layer4_outputs(1742) <= b;
    layer4_outputs(1743) <= not a;
    layer4_outputs(1744) <= not b;
    layer4_outputs(1745) <= a;
    layer4_outputs(1746) <= not b;
    layer4_outputs(1747) <= not (a xor b);
    layer4_outputs(1748) <= not b or a;
    layer4_outputs(1749) <= b and not a;
    layer4_outputs(1750) <= a;
    layer4_outputs(1751) <= not b;
    layer4_outputs(1752) <= not b or a;
    layer4_outputs(1753) <= a;
    layer4_outputs(1754) <= a;
    layer4_outputs(1755) <= b and not a;
    layer4_outputs(1756) <= not a;
    layer4_outputs(1757) <= a and b;
    layer4_outputs(1758) <= not (a or b);
    layer4_outputs(1759) <= not b or a;
    layer4_outputs(1760) <= not (a and b);
    layer4_outputs(1761) <= not a;
    layer4_outputs(1762) <= not a or b;
    layer4_outputs(1763) <= b;
    layer4_outputs(1764) <= a;
    layer4_outputs(1765) <= b;
    layer4_outputs(1766) <= not a;
    layer4_outputs(1767) <= not b or a;
    layer4_outputs(1768) <= b;
    layer4_outputs(1769) <= not (a and b);
    layer4_outputs(1770) <= b;
    layer4_outputs(1771) <= a;
    layer4_outputs(1772) <= not b or a;
    layer4_outputs(1773) <= not b;
    layer4_outputs(1774) <= not b;
    layer4_outputs(1775) <= 1'b0;
    layer4_outputs(1776) <= a and not b;
    layer4_outputs(1777) <= not a or b;
    layer4_outputs(1778) <= not (a xor b);
    layer4_outputs(1779) <= not b or a;
    layer4_outputs(1780) <= not (a or b);
    layer4_outputs(1781) <= a and b;
    layer4_outputs(1782) <= not b;
    layer4_outputs(1783) <= not a or b;
    layer4_outputs(1784) <= not a or b;
    layer4_outputs(1785) <= not a;
    layer4_outputs(1786) <= a xor b;
    layer4_outputs(1787) <= not b;
    layer4_outputs(1788) <= a;
    layer4_outputs(1789) <= not b;
    layer4_outputs(1790) <= a;
    layer4_outputs(1791) <= not b;
    layer4_outputs(1792) <= a and not b;
    layer4_outputs(1793) <= b and not a;
    layer4_outputs(1794) <= not b;
    layer4_outputs(1795) <= not b;
    layer4_outputs(1796) <= not a;
    layer4_outputs(1797) <= 1'b1;
    layer4_outputs(1798) <= b and not a;
    layer4_outputs(1799) <= b;
    layer4_outputs(1800) <= b;
    layer4_outputs(1801) <= b and not a;
    layer4_outputs(1802) <= not b;
    layer4_outputs(1803) <= a or b;
    layer4_outputs(1804) <= a;
    layer4_outputs(1805) <= not a;
    layer4_outputs(1806) <= b and not a;
    layer4_outputs(1807) <= not (a or b);
    layer4_outputs(1808) <= a and not b;
    layer4_outputs(1809) <= not b or a;
    layer4_outputs(1810) <= not b;
    layer4_outputs(1811) <= a;
    layer4_outputs(1812) <= a or b;
    layer4_outputs(1813) <= not b or a;
    layer4_outputs(1814) <= b;
    layer4_outputs(1815) <= not (a and b);
    layer4_outputs(1816) <= not a or b;
    layer4_outputs(1817) <= not a;
    layer4_outputs(1818) <= a or b;
    layer4_outputs(1819) <= b;
    layer4_outputs(1820) <= a or b;
    layer4_outputs(1821) <= not a;
    layer4_outputs(1822) <= a;
    layer4_outputs(1823) <= not (a xor b);
    layer4_outputs(1824) <= b;
    layer4_outputs(1825) <= not (a xor b);
    layer4_outputs(1826) <= not a;
    layer4_outputs(1827) <= b and not a;
    layer4_outputs(1828) <= b;
    layer4_outputs(1829) <= b and not a;
    layer4_outputs(1830) <= not a;
    layer4_outputs(1831) <= not a;
    layer4_outputs(1832) <= a;
    layer4_outputs(1833) <= b;
    layer4_outputs(1834) <= not (a or b);
    layer4_outputs(1835) <= not a or b;
    layer4_outputs(1836) <= not a;
    layer4_outputs(1837) <= not (a and b);
    layer4_outputs(1838) <= not b or a;
    layer4_outputs(1839) <= b;
    layer4_outputs(1840) <= 1'b1;
    layer4_outputs(1841) <= a and not b;
    layer4_outputs(1842) <= a and b;
    layer4_outputs(1843) <= b;
    layer4_outputs(1844) <= not b;
    layer4_outputs(1845) <= a and not b;
    layer4_outputs(1846) <= a xor b;
    layer4_outputs(1847) <= a xor b;
    layer4_outputs(1848) <= b;
    layer4_outputs(1849) <= not b;
    layer4_outputs(1850) <= a and b;
    layer4_outputs(1851) <= not b or a;
    layer4_outputs(1852) <= not (a xor b);
    layer4_outputs(1853) <= a;
    layer4_outputs(1854) <= not (a and b);
    layer4_outputs(1855) <= not b or a;
    layer4_outputs(1856) <= b and not a;
    layer4_outputs(1857) <= a;
    layer4_outputs(1858) <= not b or a;
    layer4_outputs(1859) <= a and not b;
    layer4_outputs(1860) <= not a;
    layer4_outputs(1861) <= not a or b;
    layer4_outputs(1862) <= a;
    layer4_outputs(1863) <= not b;
    layer4_outputs(1864) <= not b;
    layer4_outputs(1865) <= a and not b;
    layer4_outputs(1866) <= not b;
    layer4_outputs(1867) <= a or b;
    layer4_outputs(1868) <= a and b;
    layer4_outputs(1869) <= not b;
    layer4_outputs(1870) <= not a;
    layer4_outputs(1871) <= not (a or b);
    layer4_outputs(1872) <= not (a or b);
    layer4_outputs(1873) <= a;
    layer4_outputs(1874) <= b and not a;
    layer4_outputs(1875) <= b;
    layer4_outputs(1876) <= not (a and b);
    layer4_outputs(1877) <= not a;
    layer4_outputs(1878) <= a xor b;
    layer4_outputs(1879) <= not (a xor b);
    layer4_outputs(1880) <= not (a or b);
    layer4_outputs(1881) <= a;
    layer4_outputs(1882) <= not b;
    layer4_outputs(1883) <= b and not a;
    layer4_outputs(1884) <= b and not a;
    layer4_outputs(1885) <= not (a and b);
    layer4_outputs(1886) <= a;
    layer4_outputs(1887) <= not a or b;
    layer4_outputs(1888) <= a;
    layer4_outputs(1889) <= not b or a;
    layer4_outputs(1890) <= b;
    layer4_outputs(1891) <= not b or a;
    layer4_outputs(1892) <= not a;
    layer4_outputs(1893) <= not a;
    layer4_outputs(1894) <= not a;
    layer4_outputs(1895) <= not (a or b);
    layer4_outputs(1896) <= a and b;
    layer4_outputs(1897) <= not b;
    layer4_outputs(1898) <= a;
    layer4_outputs(1899) <= not a;
    layer4_outputs(1900) <= not a;
    layer4_outputs(1901) <= not b or a;
    layer4_outputs(1902) <= 1'b1;
    layer4_outputs(1903) <= not (a xor b);
    layer4_outputs(1904) <= a and not b;
    layer4_outputs(1905) <= not b or a;
    layer4_outputs(1906) <= a xor b;
    layer4_outputs(1907) <= not b or a;
    layer4_outputs(1908) <= not (a or b);
    layer4_outputs(1909) <= not (a and b);
    layer4_outputs(1910) <= a xor b;
    layer4_outputs(1911) <= not (a xor b);
    layer4_outputs(1912) <= a xor b;
    layer4_outputs(1913) <= a;
    layer4_outputs(1914) <= not (a xor b);
    layer4_outputs(1915) <= b and not a;
    layer4_outputs(1916) <= a or b;
    layer4_outputs(1917) <= not a;
    layer4_outputs(1918) <= b and not a;
    layer4_outputs(1919) <= b;
    layer4_outputs(1920) <= not b;
    layer4_outputs(1921) <= a xor b;
    layer4_outputs(1922) <= not b;
    layer4_outputs(1923) <= a xor b;
    layer4_outputs(1924) <= not (a and b);
    layer4_outputs(1925) <= not b or a;
    layer4_outputs(1926) <= not b or a;
    layer4_outputs(1927) <= b and not a;
    layer4_outputs(1928) <= b;
    layer4_outputs(1929) <= not b;
    layer4_outputs(1930) <= not a or b;
    layer4_outputs(1931) <= a;
    layer4_outputs(1932) <= not a or b;
    layer4_outputs(1933) <= not (a and b);
    layer4_outputs(1934) <= not a;
    layer4_outputs(1935) <= not (a and b);
    layer4_outputs(1936) <= b and not a;
    layer4_outputs(1937) <= not a;
    layer4_outputs(1938) <= a or b;
    layer4_outputs(1939) <= not a or b;
    layer4_outputs(1940) <= not b;
    layer4_outputs(1941) <= a;
    layer4_outputs(1942) <= a;
    layer4_outputs(1943) <= not (a xor b);
    layer4_outputs(1944) <= not (a or b);
    layer4_outputs(1945) <= not a or b;
    layer4_outputs(1946) <= not (a or b);
    layer4_outputs(1947) <= not a;
    layer4_outputs(1948) <= a xor b;
    layer4_outputs(1949) <= not a;
    layer4_outputs(1950) <= not (a and b);
    layer4_outputs(1951) <= a xor b;
    layer4_outputs(1952) <= a and b;
    layer4_outputs(1953) <= not b or a;
    layer4_outputs(1954) <= a and b;
    layer4_outputs(1955) <= not a;
    layer4_outputs(1956) <= not a;
    layer4_outputs(1957) <= a or b;
    layer4_outputs(1958) <= a xor b;
    layer4_outputs(1959) <= not b or a;
    layer4_outputs(1960) <= not b;
    layer4_outputs(1961) <= not a;
    layer4_outputs(1962) <= b and not a;
    layer4_outputs(1963) <= not b;
    layer4_outputs(1964) <= not a or b;
    layer4_outputs(1965) <= a;
    layer4_outputs(1966) <= not (a and b);
    layer4_outputs(1967) <= not (a xor b);
    layer4_outputs(1968) <= a or b;
    layer4_outputs(1969) <= not b or a;
    layer4_outputs(1970) <= not b;
    layer4_outputs(1971) <= b and not a;
    layer4_outputs(1972) <= b;
    layer4_outputs(1973) <= not b;
    layer4_outputs(1974) <= b;
    layer4_outputs(1975) <= not a;
    layer4_outputs(1976) <= a and b;
    layer4_outputs(1977) <= a;
    layer4_outputs(1978) <= not b;
    layer4_outputs(1979) <= not a;
    layer4_outputs(1980) <= not a or b;
    layer4_outputs(1981) <= not (a xor b);
    layer4_outputs(1982) <= not b or a;
    layer4_outputs(1983) <= 1'b1;
    layer4_outputs(1984) <= a;
    layer4_outputs(1985) <= not (a xor b);
    layer4_outputs(1986) <= a and b;
    layer4_outputs(1987) <= not (a xor b);
    layer4_outputs(1988) <= not a;
    layer4_outputs(1989) <= not (a or b);
    layer4_outputs(1990) <= not (a and b);
    layer4_outputs(1991) <= not a;
    layer4_outputs(1992) <= not b;
    layer4_outputs(1993) <= not a;
    layer4_outputs(1994) <= not (a or b);
    layer4_outputs(1995) <= not (a and b);
    layer4_outputs(1996) <= b;
    layer4_outputs(1997) <= not (a and b);
    layer4_outputs(1998) <= not a or b;
    layer4_outputs(1999) <= a or b;
    layer4_outputs(2000) <= not b;
    layer4_outputs(2001) <= b and not a;
    layer4_outputs(2002) <= a and not b;
    layer4_outputs(2003) <= b;
    layer4_outputs(2004) <= b;
    layer4_outputs(2005) <= a;
    layer4_outputs(2006) <= a or b;
    layer4_outputs(2007) <= not a;
    layer4_outputs(2008) <= not (a xor b);
    layer4_outputs(2009) <= not (a or b);
    layer4_outputs(2010) <= a and b;
    layer4_outputs(2011) <= not a;
    layer4_outputs(2012) <= not a;
    layer4_outputs(2013) <= a and b;
    layer4_outputs(2014) <= b and not a;
    layer4_outputs(2015) <= b and not a;
    layer4_outputs(2016) <= a and b;
    layer4_outputs(2017) <= not a;
    layer4_outputs(2018) <= not a or b;
    layer4_outputs(2019) <= not (a and b);
    layer4_outputs(2020) <= a xor b;
    layer4_outputs(2021) <= not (a or b);
    layer4_outputs(2022) <= a;
    layer4_outputs(2023) <= a;
    layer4_outputs(2024) <= b;
    layer4_outputs(2025) <= a;
    layer4_outputs(2026) <= a xor b;
    layer4_outputs(2027) <= a and b;
    layer4_outputs(2028) <= not (a xor b);
    layer4_outputs(2029) <= not b;
    layer4_outputs(2030) <= b and not a;
    layer4_outputs(2031) <= a;
    layer4_outputs(2032) <= not a;
    layer4_outputs(2033) <= a and not b;
    layer4_outputs(2034) <= b;
    layer4_outputs(2035) <= not (a or b);
    layer4_outputs(2036) <= b and not a;
    layer4_outputs(2037) <= a and b;
    layer4_outputs(2038) <= a and b;
    layer4_outputs(2039) <= not a;
    layer4_outputs(2040) <= not (a xor b);
    layer4_outputs(2041) <= a;
    layer4_outputs(2042) <= b;
    layer4_outputs(2043) <= not (a or b);
    layer4_outputs(2044) <= not b;
    layer4_outputs(2045) <= a xor b;
    layer4_outputs(2046) <= b and not a;
    layer4_outputs(2047) <= a;
    layer4_outputs(2048) <= a and b;
    layer4_outputs(2049) <= not (a and b);
    layer4_outputs(2050) <= not (a or b);
    layer4_outputs(2051) <= not a or b;
    layer4_outputs(2052) <= not a;
    layer4_outputs(2053) <= not a or b;
    layer4_outputs(2054) <= a;
    layer4_outputs(2055) <= not (a and b);
    layer4_outputs(2056) <= not b or a;
    layer4_outputs(2057) <= a and b;
    layer4_outputs(2058) <= a;
    layer4_outputs(2059) <= not a or b;
    layer4_outputs(2060) <= b;
    layer4_outputs(2061) <= a or b;
    layer4_outputs(2062) <= not a;
    layer4_outputs(2063) <= a;
    layer4_outputs(2064) <= a and b;
    layer4_outputs(2065) <= not b;
    layer4_outputs(2066) <= not (a xor b);
    layer4_outputs(2067) <= not b;
    layer4_outputs(2068) <= not a;
    layer4_outputs(2069) <= a;
    layer4_outputs(2070) <= not b;
    layer4_outputs(2071) <= b;
    layer4_outputs(2072) <= a;
    layer4_outputs(2073) <= a;
    layer4_outputs(2074) <= not (a xor b);
    layer4_outputs(2075) <= not b or a;
    layer4_outputs(2076) <= b;
    layer4_outputs(2077) <= a or b;
    layer4_outputs(2078) <= not (a and b);
    layer4_outputs(2079) <= a and b;
    layer4_outputs(2080) <= a;
    layer4_outputs(2081) <= not b or a;
    layer4_outputs(2082) <= a;
    layer4_outputs(2083) <= b;
    layer4_outputs(2084) <= not b;
    layer4_outputs(2085) <= not a;
    layer4_outputs(2086) <= a or b;
    layer4_outputs(2087) <= not b;
    layer4_outputs(2088) <= a or b;
    layer4_outputs(2089) <= a;
    layer4_outputs(2090) <= not a or b;
    layer4_outputs(2091) <= not b;
    layer4_outputs(2092) <= a xor b;
    layer4_outputs(2093) <= b and not a;
    layer4_outputs(2094) <= a and b;
    layer4_outputs(2095) <= not b or a;
    layer4_outputs(2096) <= a;
    layer4_outputs(2097) <= not (a xor b);
    layer4_outputs(2098) <= a;
    layer4_outputs(2099) <= a and not b;
    layer4_outputs(2100) <= a or b;
    layer4_outputs(2101) <= not b;
    layer4_outputs(2102) <= not a;
    layer4_outputs(2103) <= not (a and b);
    layer4_outputs(2104) <= a and not b;
    layer4_outputs(2105) <= not (a xor b);
    layer4_outputs(2106) <= not (a or b);
    layer4_outputs(2107) <= a xor b;
    layer4_outputs(2108) <= not (a and b);
    layer4_outputs(2109) <= not (a or b);
    layer4_outputs(2110) <= b and not a;
    layer4_outputs(2111) <= b and not a;
    layer4_outputs(2112) <= not b;
    layer4_outputs(2113) <= not (a and b);
    layer4_outputs(2114) <= not b;
    layer4_outputs(2115) <= not (a or b);
    layer4_outputs(2116) <= b and not a;
    layer4_outputs(2117) <= not b or a;
    layer4_outputs(2118) <= a and not b;
    layer4_outputs(2119) <= a;
    layer4_outputs(2120) <= b;
    layer4_outputs(2121) <= a and not b;
    layer4_outputs(2122) <= not b or a;
    layer4_outputs(2123) <= not (a xor b);
    layer4_outputs(2124) <= not (a xor b);
    layer4_outputs(2125) <= b;
    layer4_outputs(2126) <= not (a xor b);
    layer4_outputs(2127) <= a or b;
    layer4_outputs(2128) <= a;
    layer4_outputs(2129) <= a or b;
    layer4_outputs(2130) <= a;
    layer4_outputs(2131) <= a;
    layer4_outputs(2132) <= not b;
    layer4_outputs(2133) <= a or b;
    layer4_outputs(2134) <= not a or b;
    layer4_outputs(2135) <= not a or b;
    layer4_outputs(2136) <= a and b;
    layer4_outputs(2137) <= a or b;
    layer4_outputs(2138) <= b;
    layer4_outputs(2139) <= a or b;
    layer4_outputs(2140) <= b;
    layer4_outputs(2141) <= a and b;
    layer4_outputs(2142) <= a or b;
    layer4_outputs(2143) <= not (a and b);
    layer4_outputs(2144) <= not (a or b);
    layer4_outputs(2145) <= a;
    layer4_outputs(2146) <= not (a or b);
    layer4_outputs(2147) <= a;
    layer4_outputs(2148) <= b;
    layer4_outputs(2149) <= not (a xor b);
    layer4_outputs(2150) <= a and b;
    layer4_outputs(2151) <= b;
    layer4_outputs(2152) <= not a or b;
    layer4_outputs(2153) <= a and b;
    layer4_outputs(2154) <= a;
    layer4_outputs(2155) <= not a;
    layer4_outputs(2156) <= not a;
    layer4_outputs(2157) <= a;
    layer4_outputs(2158) <= b;
    layer4_outputs(2159) <= not a or b;
    layer4_outputs(2160) <= not b;
    layer4_outputs(2161) <= a or b;
    layer4_outputs(2162) <= b;
    layer4_outputs(2163) <= not b;
    layer4_outputs(2164) <= a;
    layer4_outputs(2165) <= a and b;
    layer4_outputs(2166) <= b;
    layer4_outputs(2167) <= not b or a;
    layer4_outputs(2168) <= a;
    layer4_outputs(2169) <= not a or b;
    layer4_outputs(2170) <= a or b;
    layer4_outputs(2171) <= not b or a;
    layer4_outputs(2172) <= b;
    layer4_outputs(2173) <= b;
    layer4_outputs(2174) <= not a;
    layer4_outputs(2175) <= not (a and b);
    layer4_outputs(2176) <= not b;
    layer4_outputs(2177) <= not a or b;
    layer4_outputs(2178) <= 1'b1;
    layer4_outputs(2179) <= not (a and b);
    layer4_outputs(2180) <= a;
    layer4_outputs(2181) <= not b or a;
    layer4_outputs(2182) <= a;
    layer4_outputs(2183) <= a;
    layer4_outputs(2184) <= b and not a;
    layer4_outputs(2185) <= a;
    layer4_outputs(2186) <= 1'b0;
    layer4_outputs(2187) <= b;
    layer4_outputs(2188) <= a and not b;
    layer4_outputs(2189) <= not a or b;
    layer4_outputs(2190) <= not b or a;
    layer4_outputs(2191) <= a or b;
    layer4_outputs(2192) <= not a;
    layer4_outputs(2193) <= a;
    layer4_outputs(2194) <= a;
    layer4_outputs(2195) <= not b or a;
    layer4_outputs(2196) <= not a;
    layer4_outputs(2197) <= not b;
    layer4_outputs(2198) <= not b;
    layer4_outputs(2199) <= a and not b;
    layer4_outputs(2200) <= a;
    layer4_outputs(2201) <= not (a and b);
    layer4_outputs(2202) <= not a or b;
    layer4_outputs(2203) <= a xor b;
    layer4_outputs(2204) <= a;
    layer4_outputs(2205) <= not a or b;
    layer4_outputs(2206) <= not (a and b);
    layer4_outputs(2207) <= a xor b;
    layer4_outputs(2208) <= a and b;
    layer4_outputs(2209) <= a or b;
    layer4_outputs(2210) <= not a or b;
    layer4_outputs(2211) <= not a;
    layer4_outputs(2212) <= not b or a;
    layer4_outputs(2213) <= a and b;
    layer4_outputs(2214) <= not b or a;
    layer4_outputs(2215) <= b and not a;
    layer4_outputs(2216) <= a or b;
    layer4_outputs(2217) <= not a or b;
    layer4_outputs(2218) <= a and not b;
    layer4_outputs(2219) <= not a;
    layer4_outputs(2220) <= not a or b;
    layer4_outputs(2221) <= b;
    layer4_outputs(2222) <= a;
    layer4_outputs(2223) <= a or b;
    layer4_outputs(2224) <= b;
    layer4_outputs(2225) <= not b;
    layer4_outputs(2226) <= not (a and b);
    layer4_outputs(2227) <= not b;
    layer4_outputs(2228) <= not (a and b);
    layer4_outputs(2229) <= a;
    layer4_outputs(2230) <= a;
    layer4_outputs(2231) <= a and not b;
    layer4_outputs(2232) <= not b;
    layer4_outputs(2233) <= a;
    layer4_outputs(2234) <= not a;
    layer4_outputs(2235) <= b;
    layer4_outputs(2236) <= a and b;
    layer4_outputs(2237) <= a or b;
    layer4_outputs(2238) <= not a or b;
    layer4_outputs(2239) <= b;
    layer4_outputs(2240) <= b and not a;
    layer4_outputs(2241) <= a or b;
    layer4_outputs(2242) <= a;
    layer4_outputs(2243) <= b and not a;
    layer4_outputs(2244) <= b;
    layer4_outputs(2245) <= not (a or b);
    layer4_outputs(2246) <= not a or b;
    layer4_outputs(2247) <= a and not b;
    layer4_outputs(2248) <= b and not a;
    layer4_outputs(2249) <= not a or b;
    layer4_outputs(2250) <= not b;
    layer4_outputs(2251) <= not a or b;
    layer4_outputs(2252) <= not (a or b);
    layer4_outputs(2253) <= not b;
    layer4_outputs(2254) <= a and not b;
    layer4_outputs(2255) <= not b;
    layer4_outputs(2256) <= a and not b;
    layer4_outputs(2257) <= not b;
    layer4_outputs(2258) <= b;
    layer4_outputs(2259) <= not (a or b);
    layer4_outputs(2260) <= not a;
    layer4_outputs(2261) <= a or b;
    layer4_outputs(2262) <= not b;
    layer4_outputs(2263) <= b;
    layer4_outputs(2264) <= not a;
    layer4_outputs(2265) <= a xor b;
    layer4_outputs(2266) <= not a or b;
    layer4_outputs(2267) <= b and not a;
    layer4_outputs(2268) <= not b;
    layer4_outputs(2269) <= b;
    layer4_outputs(2270) <= not a;
    layer4_outputs(2271) <= b;
    layer4_outputs(2272) <= a;
    layer4_outputs(2273) <= not b;
    layer4_outputs(2274) <= a or b;
    layer4_outputs(2275) <= 1'b0;
    layer4_outputs(2276) <= not b or a;
    layer4_outputs(2277) <= a or b;
    layer4_outputs(2278) <= not (a or b);
    layer4_outputs(2279) <= not (a or b);
    layer4_outputs(2280) <= 1'b1;
    layer4_outputs(2281) <= not (a or b);
    layer4_outputs(2282) <= b;
    layer4_outputs(2283) <= not a or b;
    layer4_outputs(2284) <= not b or a;
    layer4_outputs(2285) <= a or b;
    layer4_outputs(2286) <= b;
    layer4_outputs(2287) <= a xor b;
    layer4_outputs(2288) <= not b or a;
    layer4_outputs(2289) <= a or b;
    layer4_outputs(2290) <= a and not b;
    layer4_outputs(2291) <= a and not b;
    layer4_outputs(2292) <= a;
    layer4_outputs(2293) <= not a;
    layer4_outputs(2294) <= b and not a;
    layer4_outputs(2295) <= not (a xor b);
    layer4_outputs(2296) <= a;
    layer4_outputs(2297) <= not (a or b);
    layer4_outputs(2298) <= not (a or b);
    layer4_outputs(2299) <= not (a and b);
    layer4_outputs(2300) <= a and b;
    layer4_outputs(2301) <= a;
    layer4_outputs(2302) <= not b;
    layer4_outputs(2303) <= not a;
    layer4_outputs(2304) <= not b or a;
    layer4_outputs(2305) <= not a;
    layer4_outputs(2306) <= not (a or b);
    layer4_outputs(2307) <= b;
    layer4_outputs(2308) <= a and not b;
    layer4_outputs(2309) <= not (a and b);
    layer4_outputs(2310) <= a xor b;
    layer4_outputs(2311) <= not b or a;
    layer4_outputs(2312) <= not (a or b);
    layer4_outputs(2313) <= a and b;
    layer4_outputs(2314) <= a or b;
    layer4_outputs(2315) <= a or b;
    layer4_outputs(2316) <= not b;
    layer4_outputs(2317) <= b;
    layer4_outputs(2318) <= a or b;
    layer4_outputs(2319) <= b;
    layer4_outputs(2320) <= not a;
    layer4_outputs(2321) <= a xor b;
    layer4_outputs(2322) <= b;
    layer4_outputs(2323) <= not b;
    layer4_outputs(2324) <= b;
    layer4_outputs(2325) <= 1'b0;
    layer4_outputs(2326) <= a or b;
    layer4_outputs(2327) <= b and not a;
    layer4_outputs(2328) <= not b;
    layer4_outputs(2329) <= not (a and b);
    layer4_outputs(2330) <= b;
    layer4_outputs(2331) <= not b;
    layer4_outputs(2332) <= b;
    layer4_outputs(2333) <= a;
    layer4_outputs(2334) <= not a;
    layer4_outputs(2335) <= not b or a;
    layer4_outputs(2336) <= not a;
    layer4_outputs(2337) <= not b;
    layer4_outputs(2338) <= a;
    layer4_outputs(2339) <= not b;
    layer4_outputs(2340) <= a;
    layer4_outputs(2341) <= b and not a;
    layer4_outputs(2342) <= a and not b;
    layer4_outputs(2343) <= b;
    layer4_outputs(2344) <= a and b;
    layer4_outputs(2345) <= not a or b;
    layer4_outputs(2346) <= b;
    layer4_outputs(2347) <= b;
    layer4_outputs(2348) <= not (a or b);
    layer4_outputs(2349) <= not a or b;
    layer4_outputs(2350) <= not a or b;
    layer4_outputs(2351) <= a;
    layer4_outputs(2352) <= a xor b;
    layer4_outputs(2353) <= not (a and b);
    layer4_outputs(2354) <= a;
    layer4_outputs(2355) <= a and b;
    layer4_outputs(2356) <= not b or a;
    layer4_outputs(2357) <= not (a xor b);
    layer4_outputs(2358) <= b;
    layer4_outputs(2359) <= not b;
    layer4_outputs(2360) <= not b;
    layer4_outputs(2361) <= not a;
    layer4_outputs(2362) <= b and not a;
    layer4_outputs(2363) <= not b or a;
    layer4_outputs(2364) <= not b;
    layer4_outputs(2365) <= not a or b;
    layer4_outputs(2366) <= not (a and b);
    layer4_outputs(2367) <= a and not b;
    layer4_outputs(2368) <= a and b;
    layer4_outputs(2369) <= not a;
    layer4_outputs(2370) <= a;
    layer4_outputs(2371) <= not b or a;
    layer4_outputs(2372) <= not (a or b);
    layer4_outputs(2373) <= not (a xor b);
    layer4_outputs(2374) <= not (a and b);
    layer4_outputs(2375) <= not (a and b);
    layer4_outputs(2376) <= not (a or b);
    layer4_outputs(2377) <= b;
    layer4_outputs(2378) <= not b or a;
    layer4_outputs(2379) <= a or b;
    layer4_outputs(2380) <= a and b;
    layer4_outputs(2381) <= not a;
    layer4_outputs(2382) <= a and not b;
    layer4_outputs(2383) <= b and not a;
    layer4_outputs(2384) <= a and b;
    layer4_outputs(2385) <= not b or a;
    layer4_outputs(2386) <= a;
    layer4_outputs(2387) <= not b;
    layer4_outputs(2388) <= not b;
    layer4_outputs(2389) <= not a or b;
    layer4_outputs(2390) <= not b;
    layer4_outputs(2391) <= b and not a;
    layer4_outputs(2392) <= not b;
    layer4_outputs(2393) <= not b;
    layer4_outputs(2394) <= a or b;
    layer4_outputs(2395) <= a and not b;
    layer4_outputs(2396) <= not b;
    layer4_outputs(2397) <= not a;
    layer4_outputs(2398) <= a and b;
    layer4_outputs(2399) <= a xor b;
    layer4_outputs(2400) <= not (a xor b);
    layer4_outputs(2401) <= not (a xor b);
    layer4_outputs(2402) <= not (a xor b);
    layer4_outputs(2403) <= not (a and b);
    layer4_outputs(2404) <= b;
    layer4_outputs(2405) <= not a;
    layer4_outputs(2406) <= a and b;
    layer4_outputs(2407) <= a and b;
    layer4_outputs(2408) <= b and not a;
    layer4_outputs(2409) <= a and b;
    layer4_outputs(2410) <= not a;
    layer4_outputs(2411) <= not b;
    layer4_outputs(2412) <= not b;
    layer4_outputs(2413) <= not b or a;
    layer4_outputs(2414) <= a and not b;
    layer4_outputs(2415) <= not b;
    layer4_outputs(2416) <= a and not b;
    layer4_outputs(2417) <= not b or a;
    layer4_outputs(2418) <= a and not b;
    layer4_outputs(2419) <= a xor b;
    layer4_outputs(2420) <= a;
    layer4_outputs(2421) <= a or b;
    layer4_outputs(2422) <= a;
    layer4_outputs(2423) <= not (a or b);
    layer4_outputs(2424) <= b and not a;
    layer4_outputs(2425) <= a;
    layer4_outputs(2426) <= a or b;
    layer4_outputs(2427) <= not a;
    layer4_outputs(2428) <= a and b;
    layer4_outputs(2429) <= not a;
    layer4_outputs(2430) <= a xor b;
    layer4_outputs(2431) <= a and not b;
    layer4_outputs(2432) <= not b or a;
    layer4_outputs(2433) <= not (a and b);
    layer4_outputs(2434) <= a or b;
    layer4_outputs(2435) <= a and not b;
    layer4_outputs(2436) <= not (a and b);
    layer4_outputs(2437) <= b;
    layer4_outputs(2438) <= 1'b1;
    layer4_outputs(2439) <= not b or a;
    layer4_outputs(2440) <= a xor b;
    layer4_outputs(2441) <= a;
    layer4_outputs(2442) <= not b or a;
    layer4_outputs(2443) <= not a or b;
    layer4_outputs(2444) <= a and b;
    layer4_outputs(2445) <= a and not b;
    layer4_outputs(2446) <= a and not b;
    layer4_outputs(2447) <= a or b;
    layer4_outputs(2448) <= not b;
    layer4_outputs(2449) <= not (a xor b);
    layer4_outputs(2450) <= not a or b;
    layer4_outputs(2451) <= a xor b;
    layer4_outputs(2452) <= not a;
    layer4_outputs(2453) <= not a or b;
    layer4_outputs(2454) <= a and b;
    layer4_outputs(2455) <= not (a xor b);
    layer4_outputs(2456) <= not a;
    layer4_outputs(2457) <= a;
    layer4_outputs(2458) <= 1'b0;
    layer4_outputs(2459) <= a and b;
    layer4_outputs(2460) <= not (a xor b);
    layer4_outputs(2461) <= not (a or b);
    layer4_outputs(2462) <= not a;
    layer4_outputs(2463) <= not (a and b);
    layer4_outputs(2464) <= not b;
    layer4_outputs(2465) <= a;
    layer4_outputs(2466) <= b;
    layer4_outputs(2467) <= b and not a;
    layer4_outputs(2468) <= a;
    layer4_outputs(2469) <= not a;
    layer4_outputs(2470) <= a and b;
    layer4_outputs(2471) <= not b;
    layer4_outputs(2472) <= not a or b;
    layer4_outputs(2473) <= b and not a;
    layer4_outputs(2474) <= a;
    layer4_outputs(2475) <= not b;
    layer4_outputs(2476) <= not b or a;
    layer4_outputs(2477) <= a or b;
    layer4_outputs(2478) <= not a or b;
    layer4_outputs(2479) <= b;
    layer4_outputs(2480) <= a xor b;
    layer4_outputs(2481) <= a;
    layer4_outputs(2482) <= not (a and b);
    layer4_outputs(2483) <= not a or b;
    layer4_outputs(2484) <= a or b;
    layer4_outputs(2485) <= a and b;
    layer4_outputs(2486) <= a;
    layer4_outputs(2487) <= not a or b;
    layer4_outputs(2488) <= a xor b;
    layer4_outputs(2489) <= a or b;
    layer4_outputs(2490) <= not a or b;
    layer4_outputs(2491) <= not a;
    layer4_outputs(2492) <= b;
    layer4_outputs(2493) <= not a or b;
    layer4_outputs(2494) <= a and not b;
    layer4_outputs(2495) <= b;
    layer4_outputs(2496) <= not b or a;
    layer4_outputs(2497) <= a xor b;
    layer4_outputs(2498) <= a or b;
    layer4_outputs(2499) <= not b or a;
    layer4_outputs(2500) <= b;
    layer4_outputs(2501) <= not b;
    layer4_outputs(2502) <= not (a xor b);
    layer4_outputs(2503) <= a or b;
    layer4_outputs(2504) <= 1'b1;
    layer4_outputs(2505) <= b;
    layer4_outputs(2506) <= not (a xor b);
    layer4_outputs(2507) <= a or b;
    layer4_outputs(2508) <= not a or b;
    layer4_outputs(2509) <= not (a xor b);
    layer4_outputs(2510) <= not a or b;
    layer4_outputs(2511) <= not (a or b);
    layer4_outputs(2512) <= not a;
    layer4_outputs(2513) <= not b;
    layer4_outputs(2514) <= not a;
    layer4_outputs(2515) <= not a;
    layer4_outputs(2516) <= not b;
    layer4_outputs(2517) <= a;
    layer4_outputs(2518) <= a and b;
    layer4_outputs(2519) <= not b;
    layer4_outputs(2520) <= b;
    layer4_outputs(2521) <= a;
    layer4_outputs(2522) <= not (a and b);
    layer4_outputs(2523) <= not b;
    layer4_outputs(2524) <= b and not a;
    layer4_outputs(2525) <= not a;
    layer4_outputs(2526) <= b and not a;
    layer4_outputs(2527) <= b;
    layer4_outputs(2528) <= b;
    layer4_outputs(2529) <= a and not b;
    layer4_outputs(2530) <= not a;
    layer4_outputs(2531) <= a and b;
    layer4_outputs(2532) <= a and not b;
    layer4_outputs(2533) <= 1'b0;
    layer4_outputs(2534) <= b;
    layer4_outputs(2535) <= not (a xor b);
    layer4_outputs(2536) <= b and not a;
    layer4_outputs(2537) <= not a;
    layer4_outputs(2538) <= a;
    layer4_outputs(2539) <= not (a xor b);
    layer4_outputs(2540) <= not (a and b);
    layer4_outputs(2541) <= a and b;
    layer4_outputs(2542) <= not a;
    layer4_outputs(2543) <= not a;
    layer4_outputs(2544) <= b;
    layer4_outputs(2545) <= b;
    layer4_outputs(2546) <= not b or a;
    layer4_outputs(2547) <= b and not a;
    layer4_outputs(2548) <= a and b;
    layer4_outputs(2549) <= not a or b;
    layer4_outputs(2550) <= not a;
    layer4_outputs(2551) <= not (a xor b);
    layer4_outputs(2552) <= not (a or b);
    layer4_outputs(2553) <= not (a or b);
    layer4_outputs(2554) <= not b;
    layer4_outputs(2555) <= not (a xor b);
    layer4_outputs(2556) <= not (a or b);
    layer4_outputs(2557) <= b;
    layer4_outputs(2558) <= a or b;
    layer4_outputs(2559) <= b and not a;
    outputs(0) <= a;
    outputs(1) <= a and b;
    outputs(2) <= a or b;
    outputs(3) <= a and b;
    outputs(4) <= not b;
    outputs(5) <= a and b;
    outputs(6) <= b;
    outputs(7) <= not b;
    outputs(8) <= b;
    outputs(9) <= a and b;
    outputs(10) <= a;
    outputs(11) <= not b;
    outputs(12) <= a and b;
    outputs(13) <= not (a or b);
    outputs(14) <= a;
    outputs(15) <= not a;
    outputs(16) <= not (a or b);
    outputs(17) <= not a;
    outputs(18) <= b and not a;
    outputs(19) <= not (a and b);
    outputs(20) <= b and not a;
    outputs(21) <= a and b;
    outputs(22) <= a and not b;
    outputs(23) <= b;
    outputs(24) <= not b;
    outputs(25) <= b and not a;
    outputs(26) <= not a;
    outputs(27) <= not a;
    outputs(28) <= a and not b;
    outputs(29) <= not b;
    outputs(30) <= not a or b;
    outputs(31) <= a and not b;
    outputs(32) <= not b or a;
    outputs(33) <= a and not b;
    outputs(34) <= b and not a;
    outputs(35) <= b and not a;
    outputs(36) <= a;
    outputs(37) <= not (a xor b);
    outputs(38) <= not (a and b);
    outputs(39) <= not a;
    outputs(40) <= not (a or b);
    outputs(41) <= not b;
    outputs(42) <= not (a or b);
    outputs(43) <= not (a xor b);
    outputs(44) <= not b or a;
    outputs(45) <= a;
    outputs(46) <= not b;
    outputs(47) <= a or b;
    outputs(48) <= not a;
    outputs(49) <= not b;
    outputs(50) <= a and b;
    outputs(51) <= a;
    outputs(52) <= not a;
    outputs(53) <= a and b;
    outputs(54) <= b;
    outputs(55) <= not (a or b);
    outputs(56) <= not b or a;
    outputs(57) <= not b;
    outputs(58) <= a and not b;
    outputs(59) <= not (a or b);
    outputs(60) <= a;
    outputs(61) <= not a;
    outputs(62) <= b;
    outputs(63) <= not (a or b);
    outputs(64) <= a xor b;
    outputs(65) <= b;
    outputs(66) <= not b;
    outputs(67) <= a;
    outputs(68) <= not b or a;
    outputs(69) <= not a;
    outputs(70) <= not b;
    outputs(71) <= b;
    outputs(72) <= not (a or b);
    outputs(73) <= not b;
    outputs(74) <= b and not a;
    outputs(75) <= b and not a;
    outputs(76) <= not (a or b);
    outputs(77) <= a or b;
    outputs(78) <= b;
    outputs(79) <= not a or b;
    outputs(80) <= a;
    outputs(81) <= b;
    outputs(82) <= b and not a;
    outputs(83) <= not a or b;
    outputs(84) <= a;
    outputs(85) <= b;
    outputs(86) <= a or b;
    outputs(87) <= not (a or b);
    outputs(88) <= not b;
    outputs(89) <= b and not a;
    outputs(90) <= a or b;
    outputs(91) <= not (a or b);
    outputs(92) <= b and not a;
    outputs(93) <= b;
    outputs(94) <= not a;
    outputs(95) <= not a;
    outputs(96) <= a and b;
    outputs(97) <= not b;
    outputs(98) <= a;
    outputs(99) <= not b;
    outputs(100) <= b;
    outputs(101) <= a;
    outputs(102) <= a and b;
    outputs(103) <= not b;
    outputs(104) <= b and not a;
    outputs(105) <= not a;
    outputs(106) <= b and not a;
    outputs(107) <= not a;
    outputs(108) <= not b;
    outputs(109) <= a and b;
    outputs(110) <= not b;
    outputs(111) <= b;
    outputs(112) <= not (a and b);
    outputs(113) <= not b;
    outputs(114) <= a and not b;
    outputs(115) <= a;
    outputs(116) <= b and not a;
    outputs(117) <= not a;
    outputs(118) <= b and not a;
    outputs(119) <= a;
    outputs(120) <= a;
    outputs(121) <= b and not a;
    outputs(122) <= a and not b;
    outputs(123) <= not a;
    outputs(124) <= a and not b;
    outputs(125) <= a and not b;
    outputs(126) <= a and b;
    outputs(127) <= a and b;
    outputs(128) <= not b;
    outputs(129) <= b;
    outputs(130) <= a and b;
    outputs(131) <= b and not a;
    outputs(132) <= a xor b;
    outputs(133) <= not a;
    outputs(134) <= a and b;
    outputs(135) <= not b;
    outputs(136) <= a and b;
    outputs(137) <= a;
    outputs(138) <= b;
    outputs(139) <= not a;
    outputs(140) <= a;
    outputs(141) <= b;
    outputs(142) <= not (a xor b);
    outputs(143) <= not (a or b);
    outputs(144) <= not (a or b);
    outputs(145) <= a;
    outputs(146) <= a and not b;
    outputs(147) <= b;
    outputs(148) <= a and not b;
    outputs(149) <= not b;
    outputs(150) <= a;
    outputs(151) <= not (a or b);
    outputs(152) <= not a;
    outputs(153) <= a and b;
    outputs(154) <= a xor b;
    outputs(155) <= not (a or b);
    outputs(156) <= a xor b;
    outputs(157) <= not a;
    outputs(158) <= b;
    outputs(159) <= a and b;
    outputs(160) <= b and not a;
    outputs(161) <= a xor b;
    outputs(162) <= a xor b;
    outputs(163) <= b;
    outputs(164) <= not (a or b);
    outputs(165) <= b;
    outputs(166) <= a and b;
    outputs(167) <= not a;
    outputs(168) <= a and b;
    outputs(169) <= not b;
    outputs(170) <= not b;
    outputs(171) <= not a;
    outputs(172) <= a;
    outputs(173) <= a and not b;
    outputs(174) <= b and not a;
    outputs(175) <= not a or b;
    outputs(176) <= a;
    outputs(177) <= a and not b;
    outputs(178) <= not a;
    outputs(179) <= not b or a;
    outputs(180) <= not (a or b);
    outputs(181) <= not b;
    outputs(182) <= a and b;
    outputs(183) <= b and not a;
    outputs(184) <= a and b;
    outputs(185) <= a and not b;
    outputs(186) <= not b;
    outputs(187) <= b and not a;
    outputs(188) <= b and not a;
    outputs(189) <= a and b;
    outputs(190) <= a and not b;
    outputs(191) <= a;
    outputs(192) <= not b;
    outputs(193) <= a;
    outputs(194) <= b and not a;
    outputs(195) <= not a;
    outputs(196) <= a and not b;
    outputs(197) <= a;
    outputs(198) <= a;
    outputs(199) <= not b;
    outputs(200) <= b and not a;
    outputs(201) <= a and not b;
    outputs(202) <= not a;
    outputs(203) <= a or b;
    outputs(204) <= not a;
    outputs(205) <= not a;
    outputs(206) <= not (a or b);
    outputs(207) <= b;
    outputs(208) <= a and b;
    outputs(209) <= not b;
    outputs(210) <= a xor b;
    outputs(211) <= not a;
    outputs(212) <= b and not a;
    outputs(213) <= a;
    outputs(214) <= a and not b;
    outputs(215) <= not a;
    outputs(216) <= not a or b;
    outputs(217) <= b;
    outputs(218) <= not b;
    outputs(219) <= a and b;
    outputs(220) <= not (a or b);
    outputs(221) <= a and not b;
    outputs(222) <= not a;
    outputs(223) <= a xor b;
    outputs(224) <= not b;
    outputs(225) <= b and not a;
    outputs(226) <= not a;
    outputs(227) <= not b or a;
    outputs(228) <= not a;
    outputs(229) <= not a;
    outputs(230) <= not a;
    outputs(231) <= a;
    outputs(232) <= a xor b;
    outputs(233) <= not b or a;
    outputs(234) <= a;
    outputs(235) <= not a;
    outputs(236) <= not b;
    outputs(237) <= not (a or b);
    outputs(238) <= b;
    outputs(239) <= a or b;
    outputs(240) <= a and b;
    outputs(241) <= not b;
    outputs(242) <= a;
    outputs(243) <= a;
    outputs(244) <= b;
    outputs(245) <= b and not a;
    outputs(246) <= a and b;
    outputs(247) <= a and b;
    outputs(248) <= not a;
    outputs(249) <= not b;
    outputs(250) <= b and not a;
    outputs(251) <= not b;
    outputs(252) <= not (a or b);
    outputs(253) <= not (a and b);
    outputs(254) <= a and not b;
    outputs(255) <= not a;
    outputs(256) <= not a;
    outputs(257) <= not (a or b);
    outputs(258) <= b and not a;
    outputs(259) <= a and b;
    outputs(260) <= not (a or b);
    outputs(261) <= not a;
    outputs(262) <= a and not b;
    outputs(263) <= a and b;
    outputs(264) <= not b;
    outputs(265) <= not b;
    outputs(266) <= a and b;
    outputs(267) <= a and not b;
    outputs(268) <= a;
    outputs(269) <= a and b;
    outputs(270) <= a and b;
    outputs(271) <= not (a or b);
    outputs(272) <= a;
    outputs(273) <= a;
    outputs(274) <= not a;
    outputs(275) <= not (a or b);
    outputs(276) <= not (a or b);
    outputs(277) <= not a;
    outputs(278) <= not a;
    outputs(279) <= a and b;
    outputs(280) <= not (a xor b);
    outputs(281) <= not (a or b);
    outputs(282) <= a and not b;
    outputs(283) <= a xor b;
    outputs(284) <= a;
    outputs(285) <= a and not b;
    outputs(286) <= b and not a;
    outputs(287) <= b and not a;
    outputs(288) <= a and not b;
    outputs(289) <= b;
    outputs(290) <= not a;
    outputs(291) <= not (a or b);
    outputs(292) <= not (a or b);
    outputs(293) <= b and not a;
    outputs(294) <= b;
    outputs(295) <= b and not a;
    outputs(296) <= not b;
    outputs(297) <= a and not b;
    outputs(298) <= a and b;
    outputs(299) <= not (a or b);
    outputs(300) <= a and b;
    outputs(301) <= a and b;
    outputs(302) <= b and not a;
    outputs(303) <= a;
    outputs(304) <= not b;
    outputs(305) <= not b;
    outputs(306) <= a and b;
    outputs(307) <= not b;
    outputs(308) <= not b;
    outputs(309) <= a and not b;
    outputs(310) <= a and not b;
    outputs(311) <= not (a xor b);
    outputs(312) <= b and not a;
    outputs(313) <= a and b;
    outputs(314) <= a and not b;
    outputs(315) <= a or b;
    outputs(316) <= not b;
    outputs(317) <= b and not a;
    outputs(318) <= b;
    outputs(319) <= b and not a;
    outputs(320) <= a xor b;
    outputs(321) <= a and b;
    outputs(322) <= not b;
    outputs(323) <= a and b;
    outputs(324) <= a and not b;
    outputs(325) <= a and b;
    outputs(326) <= not (a or b);
    outputs(327) <= b;
    outputs(328) <= not (a or b);
    outputs(329) <= not b;
    outputs(330) <= a and b;
    outputs(331) <= a and not b;
    outputs(332) <= not (a or b);
    outputs(333) <= not (a xor b);
    outputs(334) <= b and not a;
    outputs(335) <= b and not a;
    outputs(336) <= a and not b;
    outputs(337) <= a;
    outputs(338) <= a and not b;
    outputs(339) <= a;
    outputs(340) <= not (a or b);
    outputs(341) <= a and not b;
    outputs(342) <= a and not b;
    outputs(343) <= a;
    outputs(344) <= not (a or b);
    outputs(345) <= a and not b;
    outputs(346) <= b and not a;
    outputs(347) <= not b;
    outputs(348) <= b and not a;
    outputs(349) <= not a;
    outputs(350) <= a and b;
    outputs(351) <= not b;
    outputs(352) <= a;
    outputs(353) <= b;
    outputs(354) <= a and not b;
    outputs(355) <= b and not a;
    outputs(356) <= a and b;
    outputs(357) <= a and not b;
    outputs(358) <= a;
    outputs(359) <= b;
    outputs(360) <= a and not b;
    outputs(361) <= not a;
    outputs(362) <= b and not a;
    outputs(363) <= a and not b;
    outputs(364) <= b;
    outputs(365) <= b;
    outputs(366) <= b and not a;
    outputs(367) <= a and not b;
    outputs(368) <= not a;
    outputs(369) <= b and not a;
    outputs(370) <= not (a or b);
    outputs(371) <= not b;
    outputs(372) <= a and not b;
    outputs(373) <= b and not a;
    outputs(374) <= a;
    outputs(375) <= b;
    outputs(376) <= a and b;
    outputs(377) <= b and not a;
    outputs(378) <= b and not a;
    outputs(379) <= b and not a;
    outputs(380) <= not b;
    outputs(381) <= not (a or b);
    outputs(382) <= a and b;
    outputs(383) <= a and b;
    outputs(384) <= not (a or b);
    outputs(385) <= a;
    outputs(386) <= b and not a;
    outputs(387) <= not (a or b);
    outputs(388) <= a;
    outputs(389) <= not (a and b);
    outputs(390) <= not (a xor b);
    outputs(391) <= a xor b;
    outputs(392) <= a and not b;
    outputs(393) <= not a;
    outputs(394) <= not (a or b);
    outputs(395) <= not a;
    outputs(396) <= a and not b;
    outputs(397) <= a xor b;
    outputs(398) <= not (a or b);
    outputs(399) <= a and not b;
    outputs(400) <= b and not a;
    outputs(401) <= not (a xor b);
    outputs(402) <= b and not a;
    outputs(403) <= a and not b;
    outputs(404) <= not (a or b);
    outputs(405) <= a and b;
    outputs(406) <= a xor b;
    outputs(407) <= not (a or b);
    outputs(408) <= b and not a;
    outputs(409) <= a and not b;
    outputs(410) <= a and b;
    outputs(411) <= a and not b;
    outputs(412) <= b;
    outputs(413) <= a;
    outputs(414) <= a;
    outputs(415) <= not a;
    outputs(416) <= a xor b;
    outputs(417) <= a and not b;
    outputs(418) <= b and not a;
    outputs(419) <= not (a or b);
    outputs(420) <= not (a or b);
    outputs(421) <= a and b;
    outputs(422) <= not a;
    outputs(423) <= a and b;
    outputs(424) <= b and not a;
    outputs(425) <= a and b;
    outputs(426) <= not (a or b);
    outputs(427) <= a and not b;
    outputs(428) <= b;
    outputs(429) <= a;
    outputs(430) <= a and not b;
    outputs(431) <= b and not a;
    outputs(432) <= a;
    outputs(433) <= b and not a;
    outputs(434) <= a and b;
    outputs(435) <= not a;
    outputs(436) <= not a;
    outputs(437) <= not (a or b);
    outputs(438) <= a and not b;
    outputs(439) <= a and b;
    outputs(440) <= not (a or b);
    outputs(441) <= a and b;
    outputs(442) <= not (a xor b);
    outputs(443) <= not b or a;
    outputs(444) <= a and b;
    outputs(445) <= not (a xor b);
    outputs(446) <= b and not a;
    outputs(447) <= not (a or b);
    outputs(448) <= b;
    outputs(449) <= not (a or b);
    outputs(450) <= a xor b;
    outputs(451) <= b;
    outputs(452) <= a and not b;
    outputs(453) <= not (a or b);
    outputs(454) <= a and b;
    outputs(455) <= not b;
    outputs(456) <= a and not b;
    outputs(457) <= b and not a;
    outputs(458) <= a;
    outputs(459) <= b and not a;
    outputs(460) <= a and b;
    outputs(461) <= a and not b;
    outputs(462) <= b and not a;
    outputs(463) <= not (a or b);
    outputs(464) <= b and not a;
    outputs(465) <= b and not a;
    outputs(466) <= not (a or b);
    outputs(467) <= not (a or b);
    outputs(468) <= a;
    outputs(469) <= not a;
    outputs(470) <= b and not a;
    outputs(471) <= not b;
    outputs(472) <= a and not b;
    outputs(473) <= a xor b;
    outputs(474) <= a and b;
    outputs(475) <= not a;
    outputs(476) <= not a;
    outputs(477) <= a and b;
    outputs(478) <= not (a or b);
    outputs(479) <= not a;
    outputs(480) <= not (a or b);
    outputs(481) <= not a;
    outputs(482) <= not b;
    outputs(483) <= a and not b;
    outputs(484) <= b;
    outputs(485) <= a and b;
    outputs(486) <= a;
    outputs(487) <= not b;
    outputs(488) <= not (a and b);
    outputs(489) <= a and not b;
    outputs(490) <= a xor b;
    outputs(491) <= a and b;
    outputs(492) <= not (a xor b);
    outputs(493) <= not (a or b);
    outputs(494) <= not a;
    outputs(495) <= b and not a;
    outputs(496) <= a and b;
    outputs(497) <= a and b;
    outputs(498) <= a and b;
    outputs(499) <= b;
    outputs(500) <= b and not a;
    outputs(501) <= a;
    outputs(502) <= not a;
    outputs(503) <= not (a or b);
    outputs(504) <= not b or a;
    outputs(505) <= a and b;
    outputs(506) <= a and b;
    outputs(507) <= a and b;
    outputs(508) <= a and not b;
    outputs(509) <= not (a xor b);
    outputs(510) <= a;
    outputs(511) <= a and b;
    outputs(512) <= a xor b;
    outputs(513) <= a xor b;
    outputs(514) <= not b;
    outputs(515) <= not (a or b);
    outputs(516) <= not (a or b);
    outputs(517) <= a or b;
    outputs(518) <= a and not b;
    outputs(519) <= not (a xor b);
    outputs(520) <= not b;
    outputs(521) <= a xor b;
    outputs(522) <= not a;
    outputs(523) <= a xor b;
    outputs(524) <= a and not b;
    outputs(525) <= a;
    outputs(526) <= b;
    outputs(527) <= a and b;
    outputs(528) <= a;
    outputs(529) <= not (a or b);
    outputs(530) <= b;
    outputs(531) <= not b;
    outputs(532) <= not (a or b);
    outputs(533) <= not b;
    outputs(534) <= a;
    outputs(535) <= a and not b;
    outputs(536) <= a;
    outputs(537) <= a and b;
    outputs(538) <= a;
    outputs(539) <= b;
    outputs(540) <= not a or b;
    outputs(541) <= b;
    outputs(542) <= a or b;
    outputs(543) <= b and not a;
    outputs(544) <= b;
    outputs(545) <= b and not a;
    outputs(546) <= not b;
    outputs(547) <= not a;
    outputs(548) <= a;
    outputs(549) <= a;
    outputs(550) <= a and b;
    outputs(551) <= b;
    outputs(552) <= not a;
    outputs(553) <= a and not b;
    outputs(554) <= not (a or b);
    outputs(555) <= b;
    outputs(556) <= b;
    outputs(557) <= not a;
    outputs(558) <= not (a or b);
    outputs(559) <= a;
    outputs(560) <= not a;
    outputs(561) <= a or b;
    outputs(562) <= a and b;
    outputs(563) <= a;
    outputs(564) <= not b;
    outputs(565) <= b and not a;
    outputs(566) <= a xor b;
    outputs(567) <= not b;
    outputs(568) <= a and b;
    outputs(569) <= b;
    outputs(570) <= a;
    outputs(571) <= not b;
    outputs(572) <= b;
    outputs(573) <= not b;
    outputs(574) <= not a;
    outputs(575) <= b and not a;
    outputs(576) <= not b;
    outputs(577) <= a;
    outputs(578) <= not (a xor b);
    outputs(579) <= a;
    outputs(580) <= b;
    outputs(581) <= b;
    outputs(582) <= a and not b;
    outputs(583) <= a and b;
    outputs(584) <= a and not b;
    outputs(585) <= not a or b;
    outputs(586) <= not b;
    outputs(587) <= a and b;
    outputs(588) <= not a;
    outputs(589) <= b and not a;
    outputs(590) <= b;
    outputs(591) <= a xor b;
    outputs(592) <= not a;
    outputs(593) <= a and b;
    outputs(594) <= a and b;
    outputs(595) <= not a;
    outputs(596) <= not (a or b);
    outputs(597) <= a;
    outputs(598) <= a or b;
    outputs(599) <= b;
    outputs(600) <= a and not b;
    outputs(601) <= not (a and b);
    outputs(602) <= not b;
    outputs(603) <= not a;
    outputs(604) <= a and b;
    outputs(605) <= a xor b;
    outputs(606) <= not (a or b);
    outputs(607) <= not a or b;
    outputs(608) <= a and not b;
    outputs(609) <= a and not b;
    outputs(610) <= b;
    outputs(611) <= a;
    outputs(612) <= not b or a;
    outputs(613) <= a and not b;
    outputs(614) <= not b;
    outputs(615) <= not a;
    outputs(616) <= not (a or b);
    outputs(617) <= a;
    outputs(618) <= b;
    outputs(619) <= a and b;
    outputs(620) <= not a;
    outputs(621) <= not b;
    outputs(622) <= not a;
    outputs(623) <= not a;
    outputs(624) <= not a or b;
    outputs(625) <= a and b;
    outputs(626) <= a and b;
    outputs(627) <= a and b;
    outputs(628) <= not a;
    outputs(629) <= a;
    outputs(630) <= b;
    outputs(631) <= b and not a;
    outputs(632) <= b and not a;
    outputs(633) <= b;
    outputs(634) <= not b;
    outputs(635) <= not b;
    outputs(636) <= not b;
    outputs(637) <= a;
    outputs(638) <= not b;
    outputs(639) <= a and not b;
    outputs(640) <= a xor b;
    outputs(641) <= not b;
    outputs(642) <= a;
    outputs(643) <= not (a and b);
    outputs(644) <= b and not a;
    outputs(645) <= not a or b;
    outputs(646) <= not (a or b);
    outputs(647) <= a;
    outputs(648) <= b and not a;
    outputs(649) <= a xor b;
    outputs(650) <= not b;
    outputs(651) <= a and not b;
    outputs(652) <= a xor b;
    outputs(653) <= not (a or b);
    outputs(654) <= not b;
    outputs(655) <= not b;
    outputs(656) <= a;
    outputs(657) <= a and b;
    outputs(658) <= not a or b;
    outputs(659) <= not b or a;
    outputs(660) <= a;
    outputs(661) <= a or b;
    outputs(662) <= b;
    outputs(663) <= a;
    outputs(664) <= not a;
    outputs(665) <= not a;
    outputs(666) <= not b;
    outputs(667) <= not b or a;
    outputs(668) <= b and not a;
    outputs(669) <= b and not a;
    outputs(670) <= b;
    outputs(671) <= not a;
    outputs(672) <= not b;
    outputs(673) <= a xor b;
    outputs(674) <= a;
    outputs(675) <= not b;
    outputs(676) <= b and not a;
    outputs(677) <= a;
    outputs(678) <= a;
    outputs(679) <= not b or a;
    outputs(680) <= b and not a;
    outputs(681) <= not a;
    outputs(682) <= not (a xor b);
    outputs(683) <= b and not a;
    outputs(684) <= not (a or b);
    outputs(685) <= a;
    outputs(686) <= a xor b;
    outputs(687) <= not a;
    outputs(688) <= a or b;
    outputs(689) <= a;
    outputs(690) <= b and not a;
    outputs(691) <= not b;
    outputs(692) <= b;
    outputs(693) <= a and b;
    outputs(694) <= a and not b;
    outputs(695) <= a xor b;
    outputs(696) <= a;
    outputs(697) <= b and not a;
    outputs(698) <= a xor b;
    outputs(699) <= not a;
    outputs(700) <= a;
    outputs(701) <= not b or a;
    outputs(702) <= a and b;
    outputs(703) <= a xor b;
    outputs(704) <= a;
    outputs(705) <= a and b;
    outputs(706) <= not b or a;
    outputs(707) <= b;
    outputs(708) <= not a;
    outputs(709) <= not (a xor b);
    outputs(710) <= b and not a;
    outputs(711) <= not (a xor b);
    outputs(712) <= a and not b;
    outputs(713) <= not a;
    outputs(714) <= a;
    outputs(715) <= not b;
    outputs(716) <= b;
    outputs(717) <= a xor b;
    outputs(718) <= not a;
    outputs(719) <= not b;
    outputs(720) <= not (a or b);
    outputs(721) <= a;
    outputs(722) <= a;
    outputs(723) <= not a;
    outputs(724) <= a;
    outputs(725) <= not b;
    outputs(726) <= not (a xor b);
    outputs(727) <= a and b;
    outputs(728) <= not b or a;
    outputs(729) <= a and not b;
    outputs(730) <= not b or a;
    outputs(731) <= not a;
    outputs(732) <= not b;
    outputs(733) <= a and not b;
    outputs(734) <= a and not b;
    outputs(735) <= a and not b;
    outputs(736) <= not (a and b);
    outputs(737) <= not a;
    outputs(738) <= a and not b;
    outputs(739) <= a and not b;
    outputs(740) <= not (a xor b);
    outputs(741) <= not a or b;
    outputs(742) <= not a or b;
    outputs(743) <= not a;
    outputs(744) <= a and b;
    outputs(745) <= a and b;
    outputs(746) <= not b or a;
    outputs(747) <= a and not b;
    outputs(748) <= not a;
    outputs(749) <= not a;
    outputs(750) <= not b;
    outputs(751) <= not b or a;
    outputs(752) <= not (a or b);
    outputs(753) <= not (a or b);
    outputs(754) <= a xor b;
    outputs(755) <= a;
    outputs(756) <= a;
    outputs(757) <= a xor b;
    outputs(758) <= not (a xor b);
    outputs(759) <= b and not a;
    outputs(760) <= not a;
    outputs(761) <= b and not a;
    outputs(762) <= not b;
    outputs(763) <= not (a or b);
    outputs(764) <= a xor b;
    outputs(765) <= not (a and b);
    outputs(766) <= b and not a;
    outputs(767) <= not b;
    outputs(768) <= not (a xor b);
    outputs(769) <= b;
    outputs(770) <= not a;
    outputs(771) <= not b or a;
    outputs(772) <= not (a xor b);
    outputs(773) <= a and not b;
    outputs(774) <= not (a or b);
    outputs(775) <= a;
    outputs(776) <= b;
    outputs(777) <= b;
    outputs(778) <= not b;
    outputs(779) <= not b;
    outputs(780) <= not b;
    outputs(781) <= a and not b;
    outputs(782) <= not b;
    outputs(783) <= not b;
    outputs(784) <= a or b;
    outputs(785) <= a and b;
    outputs(786) <= a xor b;
    outputs(787) <= a and not b;
    outputs(788) <= not (a or b);
    outputs(789) <= a;
    outputs(790) <= not a;
    outputs(791) <= not (a and b);
    outputs(792) <= not b;
    outputs(793) <= not (a xor b);
    outputs(794) <= not (a or b);
    outputs(795) <= a and b;
    outputs(796) <= not a or b;
    outputs(797) <= not a;
    outputs(798) <= b and not a;
    outputs(799) <= not b;
    outputs(800) <= not (a and b);
    outputs(801) <= a and b;
    outputs(802) <= not a;
    outputs(803) <= not a;
    outputs(804) <= not a;
    outputs(805) <= not b;
    outputs(806) <= a and b;
    outputs(807) <= not a;
    outputs(808) <= not a or b;
    outputs(809) <= not a;
    outputs(810) <= not a;
    outputs(811) <= a or b;
    outputs(812) <= b;
    outputs(813) <= a and b;
    outputs(814) <= not a;
    outputs(815) <= a and b;
    outputs(816) <= not (a and b);
    outputs(817) <= a;
    outputs(818) <= not b;
    outputs(819) <= b;
    outputs(820) <= not a;
    outputs(821) <= b;
    outputs(822) <= b and not a;
    outputs(823) <= a and not b;
    outputs(824) <= a and not b;
    outputs(825) <= b;
    outputs(826) <= a and b;
    outputs(827) <= a and b;
    outputs(828) <= not a or b;
    outputs(829) <= b;
    outputs(830) <= b;
    outputs(831) <= not b;
    outputs(832) <= not b;
    outputs(833) <= a xor b;
    outputs(834) <= a;
    outputs(835) <= a;
    outputs(836) <= a xor b;
    outputs(837) <= not b;
    outputs(838) <= not a;
    outputs(839) <= b and not a;
    outputs(840) <= b and not a;
    outputs(841) <= not a;
    outputs(842) <= a;
    outputs(843) <= not a;
    outputs(844) <= not a;
    outputs(845) <= a and not b;
    outputs(846) <= b and not a;
    outputs(847) <= not b or a;
    outputs(848) <= a;
    outputs(849) <= b and not a;
    outputs(850) <= not (a xor b);
    outputs(851) <= a and not b;
    outputs(852) <= b;
    outputs(853) <= b and not a;
    outputs(854) <= b and not a;
    outputs(855) <= b;
    outputs(856) <= not (a or b);
    outputs(857) <= not b;
    outputs(858) <= a and b;
    outputs(859) <= a;
    outputs(860) <= b and not a;
    outputs(861) <= not a;
    outputs(862) <= not a or b;
    outputs(863) <= a;
    outputs(864) <= a and b;
    outputs(865) <= a xor b;
    outputs(866) <= a and b;
    outputs(867) <= a;
    outputs(868) <= b and not a;
    outputs(869) <= a xor b;
    outputs(870) <= b;
    outputs(871) <= not a;
    outputs(872) <= not b or a;
    outputs(873) <= a;
    outputs(874) <= not b;
    outputs(875) <= not a or b;
    outputs(876) <= a xor b;
    outputs(877) <= a and b;
    outputs(878) <= not b;
    outputs(879) <= not (a or b);
    outputs(880) <= a;
    outputs(881) <= not (a or b);
    outputs(882) <= b and not a;
    outputs(883) <= a;
    outputs(884) <= b;
    outputs(885) <= not (a xor b);
    outputs(886) <= a and b;
    outputs(887) <= not (a xor b);
    outputs(888) <= b;
    outputs(889) <= a;
    outputs(890) <= not a;
    outputs(891) <= a xor b;
    outputs(892) <= a xor b;
    outputs(893) <= a and b;
    outputs(894) <= b and not a;
    outputs(895) <= a;
    outputs(896) <= b;
    outputs(897) <= not b;
    outputs(898) <= a and b;
    outputs(899) <= not b;
    outputs(900) <= a and b;
    outputs(901) <= b;
    outputs(902) <= a;
    outputs(903) <= not a;
    outputs(904) <= not (a and b);
    outputs(905) <= b and not a;
    outputs(906) <= b;
    outputs(907) <= b and not a;
    outputs(908) <= a and not b;
    outputs(909) <= not a;
    outputs(910) <= b;
    outputs(911) <= b;
    outputs(912) <= a;
    outputs(913) <= b;
    outputs(914) <= a;
    outputs(915) <= b and not a;
    outputs(916) <= a xor b;
    outputs(917) <= a;
    outputs(918) <= b;
    outputs(919) <= b;
    outputs(920) <= a;
    outputs(921) <= a and not b;
    outputs(922) <= not a;
    outputs(923) <= a and not b;
    outputs(924) <= a;
    outputs(925) <= not (a or b);
    outputs(926) <= not b;
    outputs(927) <= b;
    outputs(928) <= not b or a;
    outputs(929) <= b and not a;
    outputs(930) <= not (a xor b);
    outputs(931) <= not (a or b);
    outputs(932) <= not a;
    outputs(933) <= not (a xor b);
    outputs(934) <= not a;
    outputs(935) <= a and not b;
    outputs(936) <= a or b;
    outputs(937) <= a and b;
    outputs(938) <= a;
    outputs(939) <= a xor b;
    outputs(940) <= b;
    outputs(941) <= b and not a;
    outputs(942) <= a;
    outputs(943) <= a;
    outputs(944) <= b and not a;
    outputs(945) <= a xor b;
    outputs(946) <= a xor b;
    outputs(947) <= b;
    outputs(948) <= not b;
    outputs(949) <= a and b;
    outputs(950) <= not (a or b);
    outputs(951) <= not b;
    outputs(952) <= a;
    outputs(953) <= b and not a;
    outputs(954) <= a;
    outputs(955) <= not b;
    outputs(956) <= a;
    outputs(957) <= a and not b;
    outputs(958) <= not (a and b);
    outputs(959) <= not a;
    outputs(960) <= b;
    outputs(961) <= not a or b;
    outputs(962) <= not b;
    outputs(963) <= not (a xor b);
    outputs(964) <= b and not a;
    outputs(965) <= a;
    outputs(966) <= not (a or b);
    outputs(967) <= not (a or b);
    outputs(968) <= not (a or b);
    outputs(969) <= not a;
    outputs(970) <= not b;
    outputs(971) <= b;
    outputs(972) <= b and not a;
    outputs(973) <= not b or a;
    outputs(974) <= not a or b;
    outputs(975) <= not (a xor b);
    outputs(976) <= a and not b;
    outputs(977) <= a;
    outputs(978) <= a;
    outputs(979) <= not b or a;
    outputs(980) <= not b;
    outputs(981) <= a and b;
    outputs(982) <= b;
    outputs(983) <= a and not b;
    outputs(984) <= b;
    outputs(985) <= b and not a;
    outputs(986) <= a and not b;
    outputs(987) <= b;
    outputs(988) <= not b;
    outputs(989) <= a xor b;
    outputs(990) <= a;
    outputs(991) <= not a;
    outputs(992) <= not (a or b);
    outputs(993) <= a and b;
    outputs(994) <= a and b;
    outputs(995) <= not b;
    outputs(996) <= not a;
    outputs(997) <= b;
    outputs(998) <= b;
    outputs(999) <= a;
    outputs(1000) <= b and not a;
    outputs(1001) <= not (a and b);
    outputs(1002) <= a and b;
    outputs(1003) <= a;
    outputs(1004) <= not b;
    outputs(1005) <= b and not a;
    outputs(1006) <= not a;
    outputs(1007) <= a;
    outputs(1008) <= a or b;
    outputs(1009) <= not b;
    outputs(1010) <= not a;
    outputs(1011) <= not a or b;
    outputs(1012) <= a and b;
    outputs(1013) <= not a;
    outputs(1014) <= not (a and b);
    outputs(1015) <= not (a or b);
    outputs(1016) <= not (a or b);
    outputs(1017) <= a and b;
    outputs(1018) <= a xor b;
    outputs(1019) <= a or b;
    outputs(1020) <= a;
    outputs(1021) <= a and not b;
    outputs(1022) <= not b;
    outputs(1023) <= not a;
    outputs(1024) <= not (a or b);
    outputs(1025) <= not b;
    outputs(1026) <= a and not b;
    outputs(1027) <= not a;
    outputs(1028) <= b and not a;
    outputs(1029) <= not b;
    outputs(1030) <= not b;
    outputs(1031) <= b;
    outputs(1032) <= not b;
    outputs(1033) <= b and not a;
    outputs(1034) <= not b;
    outputs(1035) <= not b;
    outputs(1036) <= not a;
    outputs(1037) <= not a;
    outputs(1038) <= a or b;
    outputs(1039) <= a;
    outputs(1040) <= a and not b;
    outputs(1041) <= not (a or b);
    outputs(1042) <= b and not a;
    outputs(1043) <= a;
    outputs(1044) <= b and not a;
    outputs(1045) <= a;
    outputs(1046) <= not b or a;
    outputs(1047) <= not a or b;
    outputs(1048) <= not (a xor b);
    outputs(1049) <= a and b;
    outputs(1050) <= b;
    outputs(1051) <= not a or b;
    outputs(1052) <= a and b;
    outputs(1053) <= b and not a;
    outputs(1054) <= not b;
    outputs(1055) <= not (a xor b);
    outputs(1056) <= not a or b;
    outputs(1057) <= b and not a;
    outputs(1058) <= a and not b;
    outputs(1059) <= b and not a;
    outputs(1060) <= not a;
    outputs(1061) <= a;
    outputs(1062) <= not a;
    outputs(1063) <= not a;
    outputs(1064) <= a;
    outputs(1065) <= b;
    outputs(1066) <= a and not b;
    outputs(1067) <= a xor b;
    outputs(1068) <= not (a or b);
    outputs(1069) <= not b;
    outputs(1070) <= not (a xor b);
    outputs(1071) <= a;
    outputs(1072) <= not b;
    outputs(1073) <= b and not a;
    outputs(1074) <= a;
    outputs(1075) <= not (a and b);
    outputs(1076) <= a and b;
    outputs(1077) <= b and not a;
    outputs(1078) <= b and not a;
    outputs(1079) <= not (a or b);
    outputs(1080) <= b and not a;
    outputs(1081) <= b and not a;
    outputs(1082) <= a;
    outputs(1083) <= b;
    outputs(1084) <= a and b;
    outputs(1085) <= a and b;
    outputs(1086) <= not (a or b);
    outputs(1087) <= b and not a;
    outputs(1088) <= not a;
    outputs(1089) <= b and not a;
    outputs(1090) <= a and b;
    outputs(1091) <= a;
    outputs(1092) <= not a;
    outputs(1093) <= a;
    outputs(1094) <= not b;
    outputs(1095) <= a;
    outputs(1096) <= not (a and b);
    outputs(1097) <= not b;
    outputs(1098) <= not b;
    outputs(1099) <= not (a or b);
    outputs(1100) <= not (a and b);
    outputs(1101) <= a and b;
    outputs(1102) <= b and not a;
    outputs(1103) <= not (a xor b);
    outputs(1104) <= b and not a;
    outputs(1105) <= b;
    outputs(1106) <= not (a or b);
    outputs(1107) <= not a;
    outputs(1108) <= not a;
    outputs(1109) <= not (a and b);
    outputs(1110) <= a and not b;
    outputs(1111) <= a;
    outputs(1112) <= not a;
    outputs(1113) <= a and b;
    outputs(1114) <= b and not a;
    outputs(1115) <= a and not b;
    outputs(1116) <= b and not a;
    outputs(1117) <= not (a xor b);
    outputs(1118) <= a and b;
    outputs(1119) <= not b;
    outputs(1120) <= a xor b;
    outputs(1121) <= not (a and b);
    outputs(1122) <= b and not a;
    outputs(1123) <= a and not b;
    outputs(1124) <= not b or a;
    outputs(1125) <= a;
    outputs(1126) <= a;
    outputs(1127) <= not b;
    outputs(1128) <= not (a or b);
    outputs(1129) <= a and b;
    outputs(1130) <= b;
    outputs(1131) <= b and not a;
    outputs(1132) <= not (a or b);
    outputs(1133) <= a xor b;
    outputs(1134) <= a and not b;
    outputs(1135) <= not (a or b);
    outputs(1136) <= not (a or b);
    outputs(1137) <= not (a or b);
    outputs(1138) <= not b;
    outputs(1139) <= a;
    outputs(1140) <= not (a or b);
    outputs(1141) <= not (a or b);
    outputs(1142) <= b;
    outputs(1143) <= b and not a;
    outputs(1144) <= not b;
    outputs(1145) <= not (a xor b);
    outputs(1146) <= b;
    outputs(1147) <= not (a or b);
    outputs(1148) <= not b;
    outputs(1149) <= a;
    outputs(1150) <= a;
    outputs(1151) <= a and b;
    outputs(1152) <= b;
    outputs(1153) <= not b;
    outputs(1154) <= b;
    outputs(1155) <= b;
    outputs(1156) <= b;
    outputs(1157) <= a;
    outputs(1158) <= not (a or b);
    outputs(1159) <= b;
    outputs(1160) <= b and not a;
    outputs(1161) <= a;
    outputs(1162) <= not a;
    outputs(1163) <= not (a xor b);
    outputs(1164) <= b;
    outputs(1165) <= a;
    outputs(1166) <= b;
    outputs(1167) <= not b;
    outputs(1168) <= a;
    outputs(1169) <= not a;
    outputs(1170) <= not (a or b);
    outputs(1171) <= not (a or b);
    outputs(1172) <= a;
    outputs(1173) <= not (a xor b);
    outputs(1174) <= b;
    outputs(1175) <= a;
    outputs(1176) <= not (a or b);
    outputs(1177) <= a and not b;
    outputs(1178) <= b and not a;
    outputs(1179) <= b;
    outputs(1180) <= not (a or b);
    outputs(1181) <= not a;
    outputs(1182) <= b;
    outputs(1183) <= not a or b;
    outputs(1184) <= b and not a;
    outputs(1185) <= not a or b;
    outputs(1186) <= not (a or b);
    outputs(1187) <= not b;
    outputs(1188) <= a and not b;
    outputs(1189) <= a and b;
    outputs(1190) <= not b;
    outputs(1191) <= not (a or b);
    outputs(1192) <= a and b;
    outputs(1193) <= a xor b;
    outputs(1194) <= not (a xor b);
    outputs(1195) <= not b;
    outputs(1196) <= a or b;
    outputs(1197) <= not (a or b);
    outputs(1198) <= not a;
    outputs(1199) <= b;
    outputs(1200) <= b;
    outputs(1201) <= not a;
    outputs(1202) <= not b or a;
    outputs(1203) <= not a;
    outputs(1204) <= a;
    outputs(1205) <= not b;
    outputs(1206) <= b;
    outputs(1207) <= not b or a;
    outputs(1208) <= a;
    outputs(1209) <= not b;
    outputs(1210) <= not a;
    outputs(1211) <= b and not a;
    outputs(1212) <= not (a xor b);
    outputs(1213) <= not (a or b);
    outputs(1214) <= b;
    outputs(1215) <= a or b;
    outputs(1216) <= a and b;
    outputs(1217) <= b;
    outputs(1218) <= b;
    outputs(1219) <= a;
    outputs(1220) <= a and not b;
    outputs(1221) <= a and b;
    outputs(1222) <= b;
    outputs(1223) <= a;
    outputs(1224) <= a;
    outputs(1225) <= not b;
    outputs(1226) <= not (a xor b);
    outputs(1227) <= a;
    outputs(1228) <= a;
    outputs(1229) <= a xor b;
    outputs(1230) <= b and not a;
    outputs(1231) <= not a;
    outputs(1232) <= not (a or b);
    outputs(1233) <= not (a or b);
    outputs(1234) <= a;
    outputs(1235) <= a and b;
    outputs(1236) <= a;
    outputs(1237) <= not a;
    outputs(1238) <= a and not b;
    outputs(1239) <= not (a or b);
    outputs(1240) <= a xor b;
    outputs(1241) <= b;
    outputs(1242) <= not (a or b);
    outputs(1243) <= not a;
    outputs(1244) <= a and b;
    outputs(1245) <= not b;
    outputs(1246) <= b and not a;
    outputs(1247) <= b;
    outputs(1248) <= a and not b;
    outputs(1249) <= a and not b;
    outputs(1250) <= not a;
    outputs(1251) <= not a or b;
    outputs(1252) <= not a or b;
    outputs(1253) <= not (a and b);
    outputs(1254) <= not (a xor b);
    outputs(1255) <= not (a or b);
    outputs(1256) <= a and not b;
    outputs(1257) <= not b;
    outputs(1258) <= not a or b;
    outputs(1259) <= not b;
    outputs(1260) <= b;
    outputs(1261) <= not b;
    outputs(1262) <= b and not a;
    outputs(1263) <= b;
    outputs(1264) <= not a;
    outputs(1265) <= a and not b;
    outputs(1266) <= b and not a;
    outputs(1267) <= a and b;
    outputs(1268) <= a and b;
    outputs(1269) <= b;
    outputs(1270) <= not a;
    outputs(1271) <= not a;
    outputs(1272) <= not b;
    outputs(1273) <= a and b;
    outputs(1274) <= a and not b;
    outputs(1275) <= not (a xor b);
    outputs(1276) <= a;
    outputs(1277) <= b;
    outputs(1278) <= a and not b;
    outputs(1279) <= b;
    outputs(1280) <= a or b;
    outputs(1281) <= not b;
    outputs(1282) <= not b;
    outputs(1283) <= a and not b;
    outputs(1284) <= b;
    outputs(1285) <= not b;
    outputs(1286) <= not b;
    outputs(1287) <= not (a or b);
    outputs(1288) <= a and not b;
    outputs(1289) <= a or b;
    outputs(1290) <= a xor b;
    outputs(1291) <= b;
    outputs(1292) <= b and not a;
    outputs(1293) <= not (a and b);
    outputs(1294) <= not b;
    outputs(1295) <= a xor b;
    outputs(1296) <= b;
    outputs(1297) <= not (a xor b);
    outputs(1298) <= not (a or b);
    outputs(1299) <= a or b;
    outputs(1300) <= a and b;
    outputs(1301) <= b;
    outputs(1302) <= not b;
    outputs(1303) <= not b;
    outputs(1304) <= a xor b;
    outputs(1305) <= a and not b;
    outputs(1306) <= b;
    outputs(1307) <= not b;
    outputs(1308) <= b and not a;
    outputs(1309) <= not b;
    outputs(1310) <= not a;
    outputs(1311) <= not a;
    outputs(1312) <= a xor b;
    outputs(1313) <= not b;
    outputs(1314) <= not a;
    outputs(1315) <= not a;
    outputs(1316) <= not b;
    outputs(1317) <= not b;
    outputs(1318) <= a;
    outputs(1319) <= b;
    outputs(1320) <= b and not a;
    outputs(1321) <= a xor b;
    outputs(1322) <= not (a or b);
    outputs(1323) <= not b;
    outputs(1324) <= not a;
    outputs(1325) <= not (a and b);
    outputs(1326) <= b;
    outputs(1327) <= b and not a;
    outputs(1328) <= not a or b;
    outputs(1329) <= not a;
    outputs(1330) <= a;
    outputs(1331) <= not a or b;
    outputs(1332) <= not b;
    outputs(1333) <= not (a xor b);
    outputs(1334) <= b;
    outputs(1335) <= b;
    outputs(1336) <= not (a and b);
    outputs(1337) <= not (a xor b);
    outputs(1338) <= b;
    outputs(1339) <= not a;
    outputs(1340) <= a xor b;
    outputs(1341) <= a xor b;
    outputs(1342) <= a and b;
    outputs(1343) <= b;
    outputs(1344) <= a xor b;
    outputs(1345) <= b;
    outputs(1346) <= not a or b;
    outputs(1347) <= a;
    outputs(1348) <= a;
    outputs(1349) <= not b;
    outputs(1350) <= not b;
    outputs(1351) <= a;
    outputs(1352) <= a xor b;
    outputs(1353) <= a xor b;
    outputs(1354) <= b;
    outputs(1355) <= b and not a;
    outputs(1356) <= not a;
    outputs(1357) <= not a;
    outputs(1358) <= b;
    outputs(1359) <= not a;
    outputs(1360) <= not b;
    outputs(1361) <= not (a or b);
    outputs(1362) <= not (a or b);
    outputs(1363) <= a or b;
    outputs(1364) <= b;
    outputs(1365) <= a;
    outputs(1366) <= a;
    outputs(1367) <= a;
    outputs(1368) <= not (a xor b);
    outputs(1369) <= not b;
    outputs(1370) <= not a;
    outputs(1371) <= not b;
    outputs(1372) <= not a;
    outputs(1373) <= not (a or b);
    outputs(1374) <= not (a xor b);
    outputs(1375) <= b and not a;
    outputs(1376) <= a xor b;
    outputs(1377) <= not (a xor b);
    outputs(1378) <= a xor b;
    outputs(1379) <= b;
    outputs(1380) <= b and not a;
    outputs(1381) <= b and not a;
    outputs(1382) <= not b or a;
    outputs(1383) <= a and b;
    outputs(1384) <= not (a xor b);
    outputs(1385) <= a and not b;
    outputs(1386) <= not b;
    outputs(1387) <= b;
    outputs(1388) <= not a;
    outputs(1389) <= b;
    outputs(1390) <= not (a or b);
    outputs(1391) <= not (a xor b);
    outputs(1392) <= b;
    outputs(1393) <= a;
    outputs(1394) <= a xor b;
    outputs(1395) <= a;
    outputs(1396) <= not b;
    outputs(1397) <= not b;
    outputs(1398) <= a;
    outputs(1399) <= not b or a;
    outputs(1400) <= not b;
    outputs(1401) <= not b;
    outputs(1402) <= b;
    outputs(1403) <= a or b;
    outputs(1404) <= a;
    outputs(1405) <= not b or a;
    outputs(1406) <= not a;
    outputs(1407) <= not (a xor b);
    outputs(1408) <= a and b;
    outputs(1409) <= a;
    outputs(1410) <= a xor b;
    outputs(1411) <= b;
    outputs(1412) <= not b or a;
    outputs(1413) <= b and not a;
    outputs(1414) <= not b;
    outputs(1415) <= a and not b;
    outputs(1416) <= not (a xor b);
    outputs(1417) <= not b;
    outputs(1418) <= a;
    outputs(1419) <= b and not a;
    outputs(1420) <= not a or b;
    outputs(1421) <= b and not a;
    outputs(1422) <= b;
    outputs(1423) <= b;
    outputs(1424) <= a and b;
    outputs(1425) <= b and not a;
    outputs(1426) <= b;
    outputs(1427) <= a and b;
    outputs(1428) <= b;
    outputs(1429) <= a or b;
    outputs(1430) <= a and b;
    outputs(1431) <= not a or b;
    outputs(1432) <= not a;
    outputs(1433) <= b and not a;
    outputs(1434) <= a xor b;
    outputs(1435) <= not a;
    outputs(1436) <= a and not b;
    outputs(1437) <= not a or b;
    outputs(1438) <= not b or a;
    outputs(1439) <= not (a and b);
    outputs(1440) <= a;
    outputs(1441) <= not (a xor b);
    outputs(1442) <= not (a and b);
    outputs(1443) <= a xor b;
    outputs(1444) <= a;
    outputs(1445) <= not (a xor b);
    outputs(1446) <= not a;
    outputs(1447) <= a and b;
    outputs(1448) <= a and not b;
    outputs(1449) <= b and not a;
    outputs(1450) <= a and b;
    outputs(1451) <= b and not a;
    outputs(1452) <= b and not a;
    outputs(1453) <= a and b;
    outputs(1454) <= a;
    outputs(1455) <= a;
    outputs(1456) <= not (a or b);
    outputs(1457) <= a and b;
    outputs(1458) <= not a;
    outputs(1459) <= a;
    outputs(1460) <= not (a or b);
    outputs(1461) <= a;
    outputs(1462) <= not a;
    outputs(1463) <= b and not a;
    outputs(1464) <= not (a or b);
    outputs(1465) <= a and not b;
    outputs(1466) <= b and not a;
    outputs(1467) <= not (a xor b);
    outputs(1468) <= b and not a;
    outputs(1469) <= b;
    outputs(1470) <= not a;
    outputs(1471) <= not (a or b);
    outputs(1472) <= not a;
    outputs(1473) <= b and not a;
    outputs(1474) <= a xor b;
    outputs(1475) <= a xor b;
    outputs(1476) <= b;
    outputs(1477) <= a;
    outputs(1478) <= not a or b;
    outputs(1479) <= not (a xor b);
    outputs(1480) <= not (a xor b);
    outputs(1481) <= a;
    outputs(1482) <= not b;
    outputs(1483) <= a or b;
    outputs(1484) <= not b;
    outputs(1485) <= not a;
    outputs(1486) <= b;
    outputs(1487) <= b and not a;
    outputs(1488) <= not (a xor b);
    outputs(1489) <= not (a and b);
    outputs(1490) <= not (a or b);
    outputs(1491) <= b;
    outputs(1492) <= not b;
    outputs(1493) <= b and not a;
    outputs(1494) <= not (a xor b);
    outputs(1495) <= not b;
    outputs(1496) <= a xor b;
    outputs(1497) <= not (a or b);
    outputs(1498) <= b;
    outputs(1499) <= not (a xor b);
    outputs(1500) <= b;
    outputs(1501) <= a;
    outputs(1502) <= not (a or b);
    outputs(1503) <= a;
    outputs(1504) <= b;
    outputs(1505) <= not (a and b);
    outputs(1506) <= a and not b;
    outputs(1507) <= a xor b;
    outputs(1508) <= not (a and b);
    outputs(1509) <= a and not b;
    outputs(1510) <= a and not b;
    outputs(1511) <= b;
    outputs(1512) <= not (a or b);
    outputs(1513) <= a and b;
    outputs(1514) <= not b or a;
    outputs(1515) <= not b;
    outputs(1516) <= b and not a;
    outputs(1517) <= not a;
    outputs(1518) <= not (a and b);
    outputs(1519) <= b;
    outputs(1520) <= not b;
    outputs(1521) <= not a;
    outputs(1522) <= b and not a;
    outputs(1523) <= not b;
    outputs(1524) <= not (a or b);
    outputs(1525) <= a;
    outputs(1526) <= not b;
    outputs(1527) <= not b;
    outputs(1528) <= a and not b;
    outputs(1529) <= a and not b;
    outputs(1530) <= not b;
    outputs(1531) <= not b;
    outputs(1532) <= b and not a;
    outputs(1533) <= not a or b;
    outputs(1534) <= a xor b;
    outputs(1535) <= b;
    outputs(1536) <= a;
    outputs(1537) <= b;
    outputs(1538) <= a and b;
    outputs(1539) <= not a;
    outputs(1540) <= a and b;
    outputs(1541) <= not a;
    outputs(1542) <= a and not b;
    outputs(1543) <= a xor b;
    outputs(1544) <= not a or b;
    outputs(1545) <= a xor b;
    outputs(1546) <= b and not a;
    outputs(1547) <= a xor b;
    outputs(1548) <= not b;
    outputs(1549) <= not b;
    outputs(1550) <= a and not b;
    outputs(1551) <= a and b;
    outputs(1552) <= a;
    outputs(1553) <= not b;
    outputs(1554) <= not (a xor b);
    outputs(1555) <= a;
    outputs(1556) <= not a;
    outputs(1557) <= a and not b;
    outputs(1558) <= b and not a;
    outputs(1559) <= a and b;
    outputs(1560) <= not (a or b);
    outputs(1561) <= not (a xor b);
    outputs(1562) <= not (a xor b);
    outputs(1563) <= b;
    outputs(1564) <= a;
    outputs(1565) <= not b;
    outputs(1566) <= b;
    outputs(1567) <= b;
    outputs(1568) <= not a;
    outputs(1569) <= not (a xor b);
    outputs(1570) <= a and not b;
    outputs(1571) <= a and b;
    outputs(1572) <= not b;
    outputs(1573) <= not a or b;
    outputs(1574) <= not a;
    outputs(1575) <= not a;
    outputs(1576) <= not b or a;
    outputs(1577) <= b;
    outputs(1578) <= b;
    outputs(1579) <= not b;
    outputs(1580) <= b;
    outputs(1581) <= a and b;
    outputs(1582) <= b;
    outputs(1583) <= a;
    outputs(1584) <= b and not a;
    outputs(1585) <= a;
    outputs(1586) <= not (a xor b);
    outputs(1587) <= not (a or b);
    outputs(1588) <= a xor b;
    outputs(1589) <= not (a or b);
    outputs(1590) <= not a;
    outputs(1591) <= not (a or b);
    outputs(1592) <= not (a and b);
    outputs(1593) <= b;
    outputs(1594) <= not b;
    outputs(1595) <= a;
    outputs(1596) <= b and not a;
    outputs(1597) <= not a;
    outputs(1598) <= a xor b;
    outputs(1599) <= not a or b;
    outputs(1600) <= not a;
    outputs(1601) <= not a or b;
    outputs(1602) <= not b;
    outputs(1603) <= a;
    outputs(1604) <= not b;
    outputs(1605) <= b and not a;
    outputs(1606) <= a;
    outputs(1607) <= a and b;
    outputs(1608) <= not a or b;
    outputs(1609) <= a;
    outputs(1610) <= not (a or b);
    outputs(1611) <= a and b;
    outputs(1612) <= b;
    outputs(1613) <= not b;
    outputs(1614) <= not b;
    outputs(1615) <= b;
    outputs(1616) <= a and not b;
    outputs(1617) <= not b;
    outputs(1618) <= a xor b;
    outputs(1619) <= a and b;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= a and b;
    outputs(1622) <= b;
    outputs(1623) <= b;
    outputs(1624) <= a and not b;
    outputs(1625) <= a xor b;
    outputs(1626) <= not (a xor b);
    outputs(1627) <= b;
    outputs(1628) <= b;
    outputs(1629) <= a and b;
    outputs(1630) <= not (a or b);
    outputs(1631) <= not (a or b);
    outputs(1632) <= not (a xor b);
    outputs(1633) <= not b;
    outputs(1634) <= b;
    outputs(1635) <= a and b;
    outputs(1636) <= a xor b;
    outputs(1637) <= not (a xor b);
    outputs(1638) <= a and b;
    outputs(1639) <= b and not a;
    outputs(1640) <= a;
    outputs(1641) <= a and b;
    outputs(1642) <= b;
    outputs(1643) <= not b;
    outputs(1644) <= a;
    outputs(1645) <= a and b;
    outputs(1646) <= a and not b;
    outputs(1647) <= a and not b;
    outputs(1648) <= a;
    outputs(1649) <= not b;
    outputs(1650) <= a;
    outputs(1651) <= b and not a;
    outputs(1652) <= not (a xor b);
    outputs(1653) <= not b;
    outputs(1654) <= b and not a;
    outputs(1655) <= a;
    outputs(1656) <= not a or b;
    outputs(1657) <= a and b;
    outputs(1658) <= a and b;
    outputs(1659) <= a and b;
    outputs(1660) <= a;
    outputs(1661) <= a and b;
    outputs(1662) <= a xor b;
    outputs(1663) <= a and b;
    outputs(1664) <= not a or b;
    outputs(1665) <= not b;
    outputs(1666) <= not b;
    outputs(1667) <= not b;
    outputs(1668) <= b;
    outputs(1669) <= a and not b;
    outputs(1670) <= b;
    outputs(1671) <= not b;
    outputs(1672) <= not b;
    outputs(1673) <= a and not b;
    outputs(1674) <= not a;
    outputs(1675) <= not (a and b);
    outputs(1676) <= b;
    outputs(1677) <= not a;
    outputs(1678) <= not a;
    outputs(1679) <= a;
    outputs(1680) <= not (a and b);
    outputs(1681) <= b;
    outputs(1682) <= a and not b;
    outputs(1683) <= not a;
    outputs(1684) <= b;
    outputs(1685) <= a;
    outputs(1686) <= a;
    outputs(1687) <= a;
    outputs(1688) <= b and not a;
    outputs(1689) <= a;
    outputs(1690) <= a and b;
    outputs(1691) <= a;
    outputs(1692) <= a;
    outputs(1693) <= a xor b;
    outputs(1694) <= not (a xor b);
    outputs(1695) <= not (a xor b);
    outputs(1696) <= b and not a;
    outputs(1697) <= not b;
    outputs(1698) <= b and not a;
    outputs(1699) <= a and not b;
    outputs(1700) <= not b;
    outputs(1701) <= not b;
    outputs(1702) <= not a or b;
    outputs(1703) <= not (a or b);
    outputs(1704) <= b and not a;
    outputs(1705) <= not (a xor b);
    outputs(1706) <= a and b;
    outputs(1707) <= not b;
    outputs(1708) <= a and not b;
    outputs(1709) <= not b;
    outputs(1710) <= not (a xor b);
    outputs(1711) <= a;
    outputs(1712) <= a xor b;
    outputs(1713) <= a and b;
    outputs(1714) <= not b;
    outputs(1715) <= a xor b;
    outputs(1716) <= not b;
    outputs(1717) <= not (a and b);
    outputs(1718) <= a;
    outputs(1719) <= not a;
    outputs(1720) <= not a;
    outputs(1721) <= not b;
    outputs(1722) <= not (a xor b);
    outputs(1723) <= not a;
    outputs(1724) <= not a;
    outputs(1725) <= b and not a;
    outputs(1726) <= not b;
    outputs(1727) <= not (a and b);
    outputs(1728) <= a and b;
    outputs(1729) <= b;
    outputs(1730) <= a and not b;
    outputs(1731) <= b;
    outputs(1732) <= b;
    outputs(1733) <= a xor b;
    outputs(1734) <= a and not b;
    outputs(1735) <= a and b;
    outputs(1736) <= a or b;
    outputs(1737) <= b;
    outputs(1738) <= not a;
    outputs(1739) <= not (a or b);
    outputs(1740) <= not b;
    outputs(1741) <= a and b;
    outputs(1742) <= not (a xor b);
    outputs(1743) <= a xor b;
    outputs(1744) <= a;
    outputs(1745) <= not b;
    outputs(1746) <= not (a xor b);
    outputs(1747) <= not (a or b);
    outputs(1748) <= a and b;
    outputs(1749) <= not a or b;
    outputs(1750) <= b;
    outputs(1751) <= b and not a;
    outputs(1752) <= not b;
    outputs(1753) <= b;
    outputs(1754) <= a;
    outputs(1755) <= not (a or b);
    outputs(1756) <= a xor b;
    outputs(1757) <= not b or a;
    outputs(1758) <= not (a xor b);
    outputs(1759) <= a and b;
    outputs(1760) <= not b;
    outputs(1761) <= not b;
    outputs(1762) <= not b or a;
    outputs(1763) <= not a or b;
    outputs(1764) <= b;
    outputs(1765) <= not b or a;
    outputs(1766) <= a or b;
    outputs(1767) <= a;
    outputs(1768) <= not b;
    outputs(1769) <= b and not a;
    outputs(1770) <= not b;
    outputs(1771) <= b and not a;
    outputs(1772) <= not b;
    outputs(1773) <= b;
    outputs(1774) <= a and not b;
    outputs(1775) <= not b;
    outputs(1776) <= b;
    outputs(1777) <= not b;
    outputs(1778) <= not b;
    outputs(1779) <= not a;
    outputs(1780) <= a and not b;
    outputs(1781) <= not a;
    outputs(1782) <= not a;
    outputs(1783) <= b;
    outputs(1784) <= b;
    outputs(1785) <= a;
    outputs(1786) <= b;
    outputs(1787) <= not b;
    outputs(1788) <= b and not a;
    outputs(1789) <= a;
    outputs(1790) <= b;
    outputs(1791) <= a and not b;
    outputs(1792) <= b;
    outputs(1793) <= not (a or b);
    outputs(1794) <= not (a or b);
    outputs(1795) <= b and not a;
    outputs(1796) <= b;
    outputs(1797) <= not b;
    outputs(1798) <= b;
    outputs(1799) <= a;
    outputs(1800) <= a and not b;
    outputs(1801) <= a and b;
    outputs(1802) <= a and b;
    outputs(1803) <= b;
    outputs(1804) <= b;
    outputs(1805) <= a and b;
    outputs(1806) <= not a;
    outputs(1807) <= a and b;
    outputs(1808) <= not (a or b);
    outputs(1809) <= a and b;
    outputs(1810) <= a and b;
    outputs(1811) <= b and not a;
    outputs(1812) <= not (a xor b);
    outputs(1813) <= a and b;
    outputs(1814) <= not a;
    outputs(1815) <= a and not b;
    outputs(1816) <= a and not b;
    outputs(1817) <= a and b;
    outputs(1818) <= not b;
    outputs(1819) <= b;
    outputs(1820) <= a and not b;
    outputs(1821) <= not a or b;
    outputs(1822) <= a;
    outputs(1823) <= b;
    outputs(1824) <= b and not a;
    outputs(1825) <= a;
    outputs(1826) <= not b;
    outputs(1827) <= a and not b;
    outputs(1828) <= a;
    outputs(1829) <= not (a and b);
    outputs(1830) <= b;
    outputs(1831) <= a;
    outputs(1832) <= a;
    outputs(1833) <= a xor b;
    outputs(1834) <= a and not b;
    outputs(1835) <= a and not b;
    outputs(1836) <= not (a or b);
    outputs(1837) <= a and not b;
    outputs(1838) <= not a or b;
    outputs(1839) <= not (a or b);
    outputs(1840) <= not (a and b);
    outputs(1841) <= a or b;
    outputs(1842) <= not a;
    outputs(1843) <= b and not a;
    outputs(1844) <= a or b;
    outputs(1845) <= b and not a;
    outputs(1846) <= b and not a;
    outputs(1847) <= a;
    outputs(1848) <= not a;
    outputs(1849) <= a;
    outputs(1850) <= not b;
    outputs(1851) <= not (a or b);
    outputs(1852) <= a and b;
    outputs(1853) <= b;
    outputs(1854) <= not a;
    outputs(1855) <= b and not a;
    outputs(1856) <= b and not a;
    outputs(1857) <= not b;
    outputs(1858) <= not (a or b);
    outputs(1859) <= not (a or b);
    outputs(1860) <= b and not a;
    outputs(1861) <= not a;
    outputs(1862) <= a;
    outputs(1863) <= a and not b;
    outputs(1864) <= not (a or b);
    outputs(1865) <= a and b;
    outputs(1866) <= a and not b;
    outputs(1867) <= not a;
    outputs(1868) <= not b;
    outputs(1869) <= b;
    outputs(1870) <= not (a xor b);
    outputs(1871) <= not (a or b);
    outputs(1872) <= a and not b;
    outputs(1873) <= a and not b;
    outputs(1874) <= a or b;
    outputs(1875) <= not (a xor b);
    outputs(1876) <= a and not b;
    outputs(1877) <= not (a xor b);
    outputs(1878) <= a;
    outputs(1879) <= a;
    outputs(1880) <= a and b;
    outputs(1881) <= a;
    outputs(1882) <= b and not a;
    outputs(1883) <= b;
    outputs(1884) <= a and not b;
    outputs(1885) <= b;
    outputs(1886) <= a xor b;
    outputs(1887) <= a and b;
    outputs(1888) <= not (a or b);
    outputs(1889) <= b;
    outputs(1890) <= a;
    outputs(1891) <= b;
    outputs(1892) <= not a;
    outputs(1893) <= a and not b;
    outputs(1894) <= b;
    outputs(1895) <= a and b;
    outputs(1896) <= b;
    outputs(1897) <= not (a xor b);
    outputs(1898) <= a and not b;
    outputs(1899) <= a and b;
    outputs(1900) <= b and not a;
    outputs(1901) <= a xor b;
    outputs(1902) <= not b;
    outputs(1903) <= b and not a;
    outputs(1904) <= not a;
    outputs(1905) <= a;
    outputs(1906) <= b and not a;
    outputs(1907) <= a and not b;
    outputs(1908) <= not a;
    outputs(1909) <= not (a or b);
    outputs(1910) <= not a;
    outputs(1911) <= a and b;
    outputs(1912) <= a and b;
    outputs(1913) <= a;
    outputs(1914) <= a and not b;
    outputs(1915) <= b and not a;
    outputs(1916) <= a;
    outputs(1917) <= not (a xor b);
    outputs(1918) <= a xor b;
    outputs(1919) <= a and not b;
    outputs(1920) <= a and b;
    outputs(1921) <= a and b;
    outputs(1922) <= b and not a;
    outputs(1923) <= b and not a;
    outputs(1924) <= a and not b;
    outputs(1925) <= a and not b;
    outputs(1926) <= a and b;
    outputs(1927) <= b and not a;
    outputs(1928) <= b;
    outputs(1929) <= a xor b;
    outputs(1930) <= not b;
    outputs(1931) <= a and not b;
    outputs(1932) <= not (a xor b);
    outputs(1933) <= not (a or b);
    outputs(1934) <= a and not b;
    outputs(1935) <= b and not a;
    outputs(1936) <= b and not a;
    outputs(1937) <= a and b;
    outputs(1938) <= a and not b;
    outputs(1939) <= a and b;
    outputs(1940) <= b and not a;
    outputs(1941) <= a;
    outputs(1942) <= not a;
    outputs(1943) <= b;
    outputs(1944) <= a and not b;
    outputs(1945) <= b and not a;
    outputs(1946) <= not a;
    outputs(1947) <= not a;
    outputs(1948) <= not (a or b);
    outputs(1949) <= a and b;
    outputs(1950) <= b;
    outputs(1951) <= not a or b;
    outputs(1952) <= not b;
    outputs(1953) <= b and not a;
    outputs(1954) <= a;
    outputs(1955) <= a and not b;
    outputs(1956) <= a;
    outputs(1957) <= a and b;
    outputs(1958) <= a and not b;
    outputs(1959) <= b and not a;
    outputs(1960) <= a and not b;
    outputs(1961) <= not (a xor b);
    outputs(1962) <= not b;
    outputs(1963) <= not b;
    outputs(1964) <= a;
    outputs(1965) <= not a;
    outputs(1966) <= a xor b;
    outputs(1967) <= not b;
    outputs(1968) <= not a;
    outputs(1969) <= not (a or b);
    outputs(1970) <= a and not b;
    outputs(1971) <= a and b;
    outputs(1972) <= not a;
    outputs(1973) <= a and b;
    outputs(1974) <= a and not b;
    outputs(1975) <= a and not b;
    outputs(1976) <= a;
    outputs(1977) <= a;
    outputs(1978) <= a and not b;
    outputs(1979) <= a;
    outputs(1980) <= not (a or b);
    outputs(1981) <= a and b;
    outputs(1982) <= b and not a;
    outputs(1983) <= b and not a;
    outputs(1984) <= b;
    outputs(1985) <= a xor b;
    outputs(1986) <= not a;
    outputs(1987) <= not (a or b);
    outputs(1988) <= a and b;
    outputs(1989) <= not a;
    outputs(1990) <= b;
    outputs(1991) <= a and b;
    outputs(1992) <= a and b;
    outputs(1993) <= b and not a;
    outputs(1994) <= a and not b;
    outputs(1995) <= not a;
    outputs(1996) <= a and b;
    outputs(1997) <= a;
    outputs(1998) <= not (a or b);
    outputs(1999) <= b;
    outputs(2000) <= a;
    outputs(2001) <= a;
    outputs(2002) <= not (a or b);
    outputs(2003) <= a and not b;
    outputs(2004) <= a and not b;
    outputs(2005) <= a and b;
    outputs(2006) <= not a or b;
    outputs(2007) <= a;
    outputs(2008) <= not a;
    outputs(2009) <= a and b;
    outputs(2010) <= a;
    outputs(2011) <= not a;
    outputs(2012) <= a;
    outputs(2013) <= not (a xor b);
    outputs(2014) <= a and not b;
    outputs(2015) <= not a;
    outputs(2016) <= not (a xor b);
    outputs(2017) <= a and not b;
    outputs(2018) <= a and b;
    outputs(2019) <= not (a or b);
    outputs(2020) <= a and b;
    outputs(2021) <= a;
    outputs(2022) <= a;
    outputs(2023) <= a;
    outputs(2024) <= a and b;
    outputs(2025) <= a and not b;
    outputs(2026) <= b and not a;
    outputs(2027) <= a xor b;
    outputs(2028) <= a and b;
    outputs(2029) <= not a;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= not (a xor b);
    outputs(2032) <= a and b;
    outputs(2033) <= not (a or b);
    outputs(2034) <= b and not a;
    outputs(2035) <= a;
    outputs(2036) <= a;
    outputs(2037) <= a;
    outputs(2038) <= not a;
    outputs(2039) <= not a;
    outputs(2040) <= not b;
    outputs(2041) <= not a;
    outputs(2042) <= not (a xor b);
    outputs(2043) <= b and not a;
    outputs(2044) <= not b;
    outputs(2045) <= a and b;
    outputs(2046) <= a;
    outputs(2047) <= not (a xor b);
    outputs(2048) <= a;
    outputs(2049) <= a xor b;
    outputs(2050) <= not (a and b);
    outputs(2051) <= a;
    outputs(2052) <= a;
    outputs(2053) <= not b;
    outputs(2054) <= a xor b;
    outputs(2055) <= not (a xor b);
    outputs(2056) <= a;
    outputs(2057) <= not (a and b);
    outputs(2058) <= a xor b;
    outputs(2059) <= not b or a;
    outputs(2060) <= b;
    outputs(2061) <= b;
    outputs(2062) <= a;
    outputs(2063) <= a xor b;
    outputs(2064) <= not (a xor b);
    outputs(2065) <= a;
    outputs(2066) <= not a or b;
    outputs(2067) <= b and not a;
    outputs(2068) <= not (a and b);
    outputs(2069) <= not b;
    outputs(2070) <= b;
    outputs(2071) <= not a;
    outputs(2072) <= b;
    outputs(2073) <= a xor b;
    outputs(2074) <= not a;
    outputs(2075) <= not b;
    outputs(2076) <= not a;
    outputs(2077) <= not (a and b);
    outputs(2078) <= b;
    outputs(2079) <= not (a and b);
    outputs(2080) <= a;
    outputs(2081) <= not a;
    outputs(2082) <= b and not a;
    outputs(2083) <= a or b;
    outputs(2084) <= not a;
    outputs(2085) <= a or b;
    outputs(2086) <= not (a or b);
    outputs(2087) <= not b;
    outputs(2088) <= not (a xor b);
    outputs(2089) <= a or b;
    outputs(2090) <= not (a or b);
    outputs(2091) <= a and b;
    outputs(2092) <= a;
    outputs(2093) <= a and b;
    outputs(2094) <= a xor b;
    outputs(2095) <= a and b;
    outputs(2096) <= not (a or b);
    outputs(2097) <= not a;
    outputs(2098) <= b and not a;
    outputs(2099) <= b;
    outputs(2100) <= a and b;
    outputs(2101) <= not (a or b);
    outputs(2102) <= a;
    outputs(2103) <= not b;
    outputs(2104) <= not b or a;
    outputs(2105) <= a;
    outputs(2106) <= a;
    outputs(2107) <= not (a xor b);
    outputs(2108) <= a and not b;
    outputs(2109) <= b and not a;
    outputs(2110) <= a and b;
    outputs(2111) <= a and not b;
    outputs(2112) <= not a;
    outputs(2113) <= not (a or b);
    outputs(2114) <= not b;
    outputs(2115) <= not (a or b);
    outputs(2116) <= b and not a;
    outputs(2117) <= not (a or b);
    outputs(2118) <= a or b;
    outputs(2119) <= not a;
    outputs(2120) <= not b;
    outputs(2121) <= not a;
    outputs(2122) <= a;
    outputs(2123) <= not b;
    outputs(2124) <= not a;
    outputs(2125) <= not (a or b);
    outputs(2126) <= b;
    outputs(2127) <= a;
    outputs(2128) <= a;
    outputs(2129) <= a and b;
    outputs(2130) <= a xor b;
    outputs(2131) <= not b;
    outputs(2132) <= not (a xor b);
    outputs(2133) <= not b or a;
    outputs(2134) <= a or b;
    outputs(2135) <= a;
    outputs(2136) <= not b;
    outputs(2137) <= b;
    outputs(2138) <= not (a xor b);
    outputs(2139) <= a xor b;
    outputs(2140) <= not (a or b);
    outputs(2141) <= not (a xor b);
    outputs(2142) <= not (a and b);
    outputs(2143) <= a xor b;
    outputs(2144) <= not (a or b);
    outputs(2145) <= not a;
    outputs(2146) <= not (a or b);
    outputs(2147) <= not a;
    outputs(2148) <= not (a and b);
    outputs(2149) <= b;
    outputs(2150) <= b;
    outputs(2151) <= b;
    outputs(2152) <= a or b;
    outputs(2153) <= a;
    outputs(2154) <= not a;
    outputs(2155) <= not (a xor b);
    outputs(2156) <= not a;
    outputs(2157) <= b and not a;
    outputs(2158) <= b;
    outputs(2159) <= not (a xor b);
    outputs(2160) <= a;
    outputs(2161) <= a and not b;
    outputs(2162) <= not (a xor b);
    outputs(2163) <= not b;
    outputs(2164) <= not b;
    outputs(2165) <= not (a xor b);
    outputs(2166) <= a xor b;
    outputs(2167) <= a;
    outputs(2168) <= b;
    outputs(2169) <= a xor b;
    outputs(2170) <= not b;
    outputs(2171) <= a;
    outputs(2172) <= a and b;
    outputs(2173) <= b;
    outputs(2174) <= b and not a;
    outputs(2175) <= not (a xor b);
    outputs(2176) <= not (a xor b);
    outputs(2177) <= not (a xor b);
    outputs(2178) <= b;
    outputs(2179) <= b and not a;
    outputs(2180) <= a xor b;
    outputs(2181) <= not a;
    outputs(2182) <= a and b;
    outputs(2183) <= not b;
    outputs(2184) <= not (a and b);
    outputs(2185) <= b;
    outputs(2186) <= not b;
    outputs(2187) <= not (a or b);
    outputs(2188) <= not (a and b);
    outputs(2189) <= a;
    outputs(2190) <= a and b;
    outputs(2191) <= not a;
    outputs(2192) <= b;
    outputs(2193) <= not b;
    outputs(2194) <= a xor b;
    outputs(2195) <= b;
    outputs(2196) <= not b;
    outputs(2197) <= a;
    outputs(2198) <= not (a or b);
    outputs(2199) <= not b;
    outputs(2200) <= a xor b;
    outputs(2201) <= a;
    outputs(2202) <= not a;
    outputs(2203) <= not b;
    outputs(2204) <= a;
    outputs(2205) <= a;
    outputs(2206) <= a and not b;
    outputs(2207) <= a;
    outputs(2208) <= b;
    outputs(2209) <= not a or b;
    outputs(2210) <= not a;
    outputs(2211) <= not a;
    outputs(2212) <= not (a or b);
    outputs(2213) <= not a;
    outputs(2214) <= not b or a;
    outputs(2215) <= not b or a;
    outputs(2216) <= not (a or b);
    outputs(2217) <= a and not b;
    outputs(2218) <= b;
    outputs(2219) <= not a;
    outputs(2220) <= a;
    outputs(2221) <= not (a xor b);
    outputs(2222) <= not (a xor b);
    outputs(2223) <= a and not b;
    outputs(2224) <= a;
    outputs(2225) <= a xor b;
    outputs(2226) <= b;
    outputs(2227) <= not (a xor b);
    outputs(2228) <= b;
    outputs(2229) <= b;
    outputs(2230) <= not (a xor b);
    outputs(2231) <= not (a and b);
    outputs(2232) <= a and not b;
    outputs(2233) <= a and b;
    outputs(2234) <= not (a xor b);
    outputs(2235) <= a and b;
    outputs(2236) <= b;
    outputs(2237) <= not a or b;
    outputs(2238) <= a or b;
    outputs(2239) <= a xor b;
    outputs(2240) <= not (a and b);
    outputs(2241) <= b and not a;
    outputs(2242) <= b;
    outputs(2243) <= not a;
    outputs(2244) <= a xor b;
    outputs(2245) <= a and not b;
    outputs(2246) <= not a;
    outputs(2247) <= a and not b;
    outputs(2248) <= not b or a;
    outputs(2249) <= not b or a;
    outputs(2250) <= b and not a;
    outputs(2251) <= not a;
    outputs(2252) <= a;
    outputs(2253) <= a and b;
    outputs(2254) <= a;
    outputs(2255) <= not b;
    outputs(2256) <= b and not a;
    outputs(2257) <= not a;
    outputs(2258) <= b and not a;
    outputs(2259) <= b;
    outputs(2260) <= a and not b;
    outputs(2261) <= b and not a;
    outputs(2262) <= b;
    outputs(2263) <= not a or b;
    outputs(2264) <= not (a or b);
    outputs(2265) <= not a or b;
    outputs(2266) <= a;
    outputs(2267) <= a and b;
    outputs(2268) <= b;
    outputs(2269) <= not b;
    outputs(2270) <= not b or a;
    outputs(2271) <= a;
    outputs(2272) <= not a or b;
    outputs(2273) <= b;
    outputs(2274) <= a;
    outputs(2275) <= a;
    outputs(2276) <= b;
    outputs(2277) <= not a;
    outputs(2278) <= not a;
    outputs(2279) <= not a or b;
    outputs(2280) <= a and b;
    outputs(2281) <= not a;
    outputs(2282) <= a xor b;
    outputs(2283) <= not (a and b);
    outputs(2284) <= not b;
    outputs(2285) <= b;
    outputs(2286) <= not (a or b);
    outputs(2287) <= not a;
    outputs(2288) <= not a;
    outputs(2289) <= a and not b;
    outputs(2290) <= a and b;
    outputs(2291) <= not b;
    outputs(2292) <= not (a xor b);
    outputs(2293) <= b;
    outputs(2294) <= not b;
    outputs(2295) <= not a;
    outputs(2296) <= not b;
    outputs(2297) <= not (a or b);
    outputs(2298) <= b and not a;
    outputs(2299) <= a;
    outputs(2300) <= a;
    outputs(2301) <= not b;
    outputs(2302) <= not (a xor b);
    outputs(2303) <= b and not a;
    outputs(2304) <= not (a or b);
    outputs(2305) <= not b;
    outputs(2306) <= not (a or b);
    outputs(2307) <= a and b;
    outputs(2308) <= not (a xor b);
    outputs(2309) <= b and not a;
    outputs(2310) <= a;
    outputs(2311) <= b;
    outputs(2312) <= b;
    outputs(2313) <= b and not a;
    outputs(2314) <= not b;
    outputs(2315) <= not b;
    outputs(2316) <= not (a and b);
    outputs(2317) <= not a;
    outputs(2318) <= not (a xor b);
    outputs(2319) <= not (a xor b);
    outputs(2320) <= a and not b;
    outputs(2321) <= b;
    outputs(2322) <= b;
    outputs(2323) <= not (a or b);
    outputs(2324) <= a or b;
    outputs(2325) <= not a;
    outputs(2326) <= b and not a;
    outputs(2327) <= a;
    outputs(2328) <= a and b;
    outputs(2329) <= not (a or b);
    outputs(2330) <= a;
    outputs(2331) <= a and not b;
    outputs(2332) <= a;
    outputs(2333) <= not b;
    outputs(2334) <= a xor b;
    outputs(2335) <= a and b;
    outputs(2336) <= not (a or b);
    outputs(2337) <= not (a and b);
    outputs(2338) <= not (a or b);
    outputs(2339) <= a and not b;
    outputs(2340) <= not (a or b);
    outputs(2341) <= not b;
    outputs(2342) <= not (a or b);
    outputs(2343) <= a and b;
    outputs(2344) <= not a;
    outputs(2345) <= a and b;
    outputs(2346) <= not a;
    outputs(2347) <= not a;
    outputs(2348) <= not b;
    outputs(2349) <= a xor b;
    outputs(2350) <= b and not a;
    outputs(2351) <= not (a or b);
    outputs(2352) <= b and not a;
    outputs(2353) <= b and not a;
    outputs(2354) <= b and not a;
    outputs(2355) <= a;
    outputs(2356) <= a or b;
    outputs(2357) <= b and not a;
    outputs(2358) <= not (a xor b);
    outputs(2359) <= not b;
    outputs(2360) <= not b;
    outputs(2361) <= not b;
    outputs(2362) <= not b;
    outputs(2363) <= b;
    outputs(2364) <= not (a or b);
    outputs(2365) <= a xor b;
    outputs(2366) <= b and not a;
    outputs(2367) <= not b;
    outputs(2368) <= not (a and b);
    outputs(2369) <= b and not a;
    outputs(2370) <= a xor b;
    outputs(2371) <= not (a or b);
    outputs(2372) <= not a;
    outputs(2373) <= a;
    outputs(2374) <= a;
    outputs(2375) <= b and not a;
    outputs(2376) <= not (a or b);
    outputs(2377) <= b;
    outputs(2378) <= a xor b;
    outputs(2379) <= not b;
    outputs(2380) <= not b;
    outputs(2381) <= not (a and b);
    outputs(2382) <= a and not b;
    outputs(2383) <= a and b;
    outputs(2384) <= b and not a;
    outputs(2385) <= not (a xor b);
    outputs(2386) <= not (a or b);
    outputs(2387) <= not (a xor b);
    outputs(2388) <= not b;
    outputs(2389) <= a and not b;
    outputs(2390) <= not (a or b);
    outputs(2391) <= a and not b;
    outputs(2392) <= not b;
    outputs(2393) <= a xor b;
    outputs(2394) <= not b;
    outputs(2395) <= a and not b;
    outputs(2396) <= not (a and b);
    outputs(2397) <= a;
    outputs(2398) <= a and b;
    outputs(2399) <= not a;
    outputs(2400) <= a;
    outputs(2401) <= b and not a;
    outputs(2402) <= not a;
    outputs(2403) <= a and b;
    outputs(2404) <= a xor b;
    outputs(2405) <= b;
    outputs(2406) <= not a;
    outputs(2407) <= not b;
    outputs(2408) <= a and b;
    outputs(2409) <= not b or a;
    outputs(2410) <= b and not a;
    outputs(2411) <= not a;
    outputs(2412) <= a;
    outputs(2413) <= not (a or b);
    outputs(2414) <= a and not b;
    outputs(2415) <= a;
    outputs(2416) <= not (a or b);
    outputs(2417) <= not (a or b);
    outputs(2418) <= a and not b;
    outputs(2419) <= not (a xor b);
    outputs(2420) <= a and not b;
    outputs(2421) <= not (a or b);
    outputs(2422) <= not (a and b);
    outputs(2423) <= not b;
    outputs(2424) <= not a or b;
    outputs(2425) <= not b;
    outputs(2426) <= not (a or b);
    outputs(2427) <= b;
    outputs(2428) <= not (a or b);
    outputs(2429) <= not b;
    outputs(2430) <= a and not b;
    outputs(2431) <= a and b;
    outputs(2432) <= a xor b;
    outputs(2433) <= b and not a;
    outputs(2434) <= not (a or b);
    outputs(2435) <= a and b;
    outputs(2436) <= a;
    outputs(2437) <= b and not a;
    outputs(2438) <= b;
    outputs(2439) <= a;
    outputs(2440) <= a and b;
    outputs(2441) <= not (a xor b);
    outputs(2442) <= a and not b;
    outputs(2443) <= a and b;
    outputs(2444) <= a and not b;
    outputs(2445) <= not b;
    outputs(2446) <= a;
    outputs(2447) <= a and not b;
    outputs(2448) <= a;
    outputs(2449) <= a and not b;
    outputs(2450) <= not b;
    outputs(2451) <= not (a or b);
    outputs(2452) <= not b;
    outputs(2453) <= a and b;
    outputs(2454) <= b;
    outputs(2455) <= a and b;
    outputs(2456) <= not b;
    outputs(2457) <= not a;
    outputs(2458) <= b and not a;
    outputs(2459) <= b;
    outputs(2460) <= b and not a;
    outputs(2461) <= not (a or b);
    outputs(2462) <= not a;
    outputs(2463) <= not b;
    outputs(2464) <= not a;
    outputs(2465) <= a and not b;
    outputs(2466) <= a and b;
    outputs(2467) <= not b;
    outputs(2468) <= b;
    outputs(2469) <= not b;
    outputs(2470) <= a and b;
    outputs(2471) <= not a;
    outputs(2472) <= not (a xor b);
    outputs(2473) <= b and not a;
    outputs(2474) <= b and not a;
    outputs(2475) <= b;
    outputs(2476) <= b;
    outputs(2477) <= not (a or b);
    outputs(2478) <= not (a or b);
    outputs(2479) <= a and b;
    outputs(2480) <= a and b;
    outputs(2481) <= not b or a;
    outputs(2482) <= not (a or b);
    outputs(2483) <= not (a or b);
    outputs(2484) <= not b;
    outputs(2485) <= not b;
    outputs(2486) <= a and b;
    outputs(2487) <= not a;
    outputs(2488) <= not a;
    outputs(2489) <= b and not a;
    outputs(2490) <= a xor b;
    outputs(2491) <= a and b;
    outputs(2492) <= a;
    outputs(2493) <= a and b;
    outputs(2494) <= b;
    outputs(2495) <= a xor b;
    outputs(2496) <= a and not b;
    outputs(2497) <= a and not b;
    outputs(2498) <= b and not a;
    outputs(2499) <= not b or a;
    outputs(2500) <= a and not b;
    outputs(2501) <= b;
    outputs(2502) <= a and not b;
    outputs(2503) <= b and not a;
    outputs(2504) <= b;
    outputs(2505) <= not a;
    outputs(2506) <= b and not a;
    outputs(2507) <= b;
    outputs(2508) <= a or b;
    outputs(2509) <= not (a xor b);
    outputs(2510) <= a xor b;
    outputs(2511) <= b;
    outputs(2512) <= not (a or b);
    outputs(2513) <= b;
    outputs(2514) <= a and b;
    outputs(2515) <= b and not a;
    outputs(2516) <= a and not b;
    outputs(2517) <= a;
    outputs(2518) <= not b;
    outputs(2519) <= a and not b;
    outputs(2520) <= a and not b;
    outputs(2521) <= not b;
    outputs(2522) <= a and not b;
    outputs(2523) <= not b;
    outputs(2524) <= a xor b;
    outputs(2525) <= a and not b;
    outputs(2526) <= not b;
    outputs(2527) <= a and not b;
    outputs(2528) <= not b;
    outputs(2529) <= a and b;
    outputs(2530) <= a and b;
    outputs(2531) <= a and b;
    outputs(2532) <= not (a and b);
    outputs(2533) <= a;
    outputs(2534) <= a and not b;
    outputs(2535) <= b;
    outputs(2536) <= a and not b;
    outputs(2537) <= a and b;
    outputs(2538) <= not b;
    outputs(2539) <= not a;
    outputs(2540) <= b and not a;
    outputs(2541) <= not (a xor b);
    outputs(2542) <= a and not b;
    outputs(2543) <= b;
    outputs(2544) <= a and not b;
    outputs(2545) <= a xor b;
    outputs(2546) <= not b or a;
    outputs(2547) <= b and not a;
    outputs(2548) <= not (a and b);
    outputs(2549) <= a and b;
    outputs(2550) <= not (a or b);
    outputs(2551) <= a;
    outputs(2552) <= a xor b;
    outputs(2553) <= not (a or b);
    outputs(2554) <= a and not b;
    outputs(2555) <= not b;
    outputs(2556) <= a and b;
    outputs(2557) <= not a;
    outputs(2558) <= a or b;
    outputs(2559) <= a and not b;
end Behavioral;
