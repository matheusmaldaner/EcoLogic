library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(12799 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(12799 downto 0);

begin

    layer0_outputs(0) <= (inputs(183)) or (inputs(44));
    layer0_outputs(1) <= (inputs(172)) xor (inputs(209));
    layer0_outputs(2) <= (inputs(239)) and not (inputs(129));
    layer0_outputs(3) <= not(inputs(200));
    layer0_outputs(4) <= not((inputs(19)) xor (inputs(26)));
    layer0_outputs(5) <= not(inputs(140));
    layer0_outputs(6) <= inputs(181);
    layer0_outputs(7) <= (inputs(103)) and (inputs(186));
    layer0_outputs(8) <= (inputs(106)) xor (inputs(254));
    layer0_outputs(9) <= inputs(170);
    layer0_outputs(10) <= (inputs(116)) or (inputs(5));
    layer0_outputs(11) <= not((inputs(182)) or (inputs(167)));
    layer0_outputs(12) <= not((inputs(115)) or (inputs(15)));
    layer0_outputs(13) <= (inputs(79)) and not (inputs(134));
    layer0_outputs(14) <= not(inputs(229));
    layer0_outputs(15) <= inputs(23);
    layer0_outputs(16) <= not(inputs(152)) or (inputs(92));
    layer0_outputs(17) <= (inputs(126)) xor (inputs(236));
    layer0_outputs(18) <= inputs(45);
    layer0_outputs(19) <= not((inputs(196)) or (inputs(56)));
    layer0_outputs(20) <= (inputs(65)) xor (inputs(29));
    layer0_outputs(21) <= '1';
    layer0_outputs(22) <= not((inputs(93)) or (inputs(12)));
    layer0_outputs(23) <= (inputs(78)) or (inputs(205));
    layer0_outputs(24) <= not(inputs(130));
    layer0_outputs(25) <= (inputs(24)) and not (inputs(204));
    layer0_outputs(26) <= not((inputs(192)) and (inputs(250)));
    layer0_outputs(27) <= not(inputs(212));
    layer0_outputs(28) <= not((inputs(95)) xor (inputs(213)));
    layer0_outputs(29) <= not((inputs(175)) or (inputs(124)));
    layer0_outputs(30) <= not((inputs(194)) and (inputs(87)));
    layer0_outputs(31) <= inputs(250);
    layer0_outputs(32) <= (inputs(16)) or (inputs(8));
    layer0_outputs(33) <= not((inputs(235)) or (inputs(17)));
    layer0_outputs(34) <= inputs(129);
    layer0_outputs(35) <= (inputs(197)) and not (inputs(50));
    layer0_outputs(36) <= inputs(119);
    layer0_outputs(37) <= (inputs(202)) and (inputs(79));
    layer0_outputs(38) <= (inputs(8)) and not (inputs(162));
    layer0_outputs(39) <= not((inputs(62)) or (inputs(48)));
    layer0_outputs(40) <= not(inputs(226)) or (inputs(1));
    layer0_outputs(41) <= not(inputs(177));
    layer0_outputs(42) <= inputs(183);
    layer0_outputs(43) <= inputs(146);
    layer0_outputs(44) <= not(inputs(1));
    layer0_outputs(45) <= not(inputs(237)) or (inputs(179));
    layer0_outputs(46) <= not((inputs(150)) xor (inputs(111)));
    layer0_outputs(47) <= not((inputs(78)) xor (inputs(92)));
    layer0_outputs(48) <= not(inputs(219)) or (inputs(15));
    layer0_outputs(49) <= inputs(10);
    layer0_outputs(50) <= not((inputs(29)) or (inputs(31)));
    layer0_outputs(51) <= (inputs(239)) or (inputs(161));
    layer0_outputs(52) <= inputs(218);
    layer0_outputs(53) <= not((inputs(46)) xor (inputs(233)));
    layer0_outputs(54) <= not((inputs(178)) or (inputs(186)));
    layer0_outputs(55) <= (inputs(81)) or (inputs(254));
    layer0_outputs(56) <= not((inputs(196)) xor (inputs(74)));
    layer0_outputs(57) <= (inputs(154)) xor (inputs(74));
    layer0_outputs(58) <= (inputs(75)) xor (inputs(177));
    layer0_outputs(59) <= not(inputs(70));
    layer0_outputs(60) <= not(inputs(255)) or (inputs(71));
    layer0_outputs(61) <= not((inputs(169)) xor (inputs(234)));
    layer0_outputs(62) <= inputs(162);
    layer0_outputs(63) <= not(inputs(213)) or (inputs(65));
    layer0_outputs(64) <= not((inputs(145)) or (inputs(162)));
    layer0_outputs(65) <= not(inputs(171));
    layer0_outputs(66) <= not(inputs(224));
    layer0_outputs(67) <= '0';
    layer0_outputs(68) <= (inputs(0)) xor (inputs(203));
    layer0_outputs(69) <= inputs(210);
    layer0_outputs(70) <= (inputs(128)) or (inputs(56));
    layer0_outputs(71) <= (inputs(43)) and not (inputs(237));
    layer0_outputs(72) <= (inputs(24)) and not (inputs(131));
    layer0_outputs(73) <= not((inputs(245)) or (inputs(67)));
    layer0_outputs(74) <= (inputs(248)) or (inputs(126));
    layer0_outputs(75) <= (inputs(20)) or (inputs(47));
    layer0_outputs(76) <= (inputs(183)) and not (inputs(48));
    layer0_outputs(77) <= (inputs(29)) xor (inputs(82));
    layer0_outputs(78) <= not((inputs(123)) or (inputs(1)));
    layer0_outputs(79) <= not(inputs(167)) or (inputs(249));
    layer0_outputs(80) <= (inputs(171)) and not (inputs(78));
    layer0_outputs(81) <= (inputs(52)) and not (inputs(227));
    layer0_outputs(82) <= not(inputs(216));
    layer0_outputs(83) <= inputs(18);
    layer0_outputs(84) <= (inputs(11)) or (inputs(127));
    layer0_outputs(85) <= '0';
    layer0_outputs(86) <= not(inputs(110));
    layer0_outputs(87) <= not(inputs(124));
    layer0_outputs(88) <= (inputs(111)) or (inputs(218));
    layer0_outputs(89) <= not((inputs(213)) or (inputs(249)));
    layer0_outputs(90) <= not(inputs(156)) or (inputs(226));
    layer0_outputs(91) <= not(inputs(118)) or (inputs(124));
    layer0_outputs(92) <= not((inputs(47)) and (inputs(87)));
    layer0_outputs(93) <= not(inputs(35)) or (inputs(127));
    layer0_outputs(94) <= not(inputs(147));
    layer0_outputs(95) <= (inputs(109)) and not (inputs(128));
    layer0_outputs(96) <= not(inputs(208));
    layer0_outputs(97) <= not(inputs(52)) or (inputs(193));
    layer0_outputs(98) <= (inputs(146)) or (inputs(85));
    layer0_outputs(99) <= not((inputs(50)) or (inputs(103)));
    layer0_outputs(100) <= not((inputs(179)) xor (inputs(190)));
    layer0_outputs(101) <= not((inputs(152)) or (inputs(52)));
    layer0_outputs(102) <= not(inputs(164)) or (inputs(78));
    layer0_outputs(103) <= not(inputs(98));
    layer0_outputs(104) <= not((inputs(157)) or (inputs(28)));
    layer0_outputs(105) <= (inputs(72)) xor (inputs(52));
    layer0_outputs(106) <= inputs(65);
    layer0_outputs(107) <= inputs(43);
    layer0_outputs(108) <= (inputs(32)) xor (inputs(101));
    layer0_outputs(109) <= not(inputs(108));
    layer0_outputs(110) <= not((inputs(238)) or (inputs(244)));
    layer0_outputs(111) <= not(inputs(41));
    layer0_outputs(112) <= inputs(178);
    layer0_outputs(113) <= inputs(206);
    layer0_outputs(114) <= (inputs(70)) or (inputs(216));
    layer0_outputs(115) <= not((inputs(112)) and (inputs(235)));
    layer0_outputs(116) <= not(inputs(250));
    layer0_outputs(117) <= not(inputs(169));
    layer0_outputs(118) <= (inputs(168)) and not (inputs(200));
    layer0_outputs(119) <= not(inputs(244));
    layer0_outputs(120) <= (inputs(51)) or (inputs(21));
    layer0_outputs(121) <= not(inputs(5)) or (inputs(113));
    layer0_outputs(122) <= not(inputs(97)) or (inputs(16));
    layer0_outputs(123) <= not((inputs(206)) or (inputs(227)));
    layer0_outputs(124) <= not((inputs(159)) or (inputs(78)));
    layer0_outputs(125) <= not((inputs(143)) or (inputs(165)));
    layer0_outputs(126) <= not(inputs(78)) or (inputs(253));
    layer0_outputs(127) <= (inputs(30)) xor (inputs(43));
    layer0_outputs(128) <= (inputs(178)) and not (inputs(15));
    layer0_outputs(129) <= (inputs(82)) and not (inputs(176));
    layer0_outputs(130) <= inputs(102);
    layer0_outputs(131) <= (inputs(236)) xor (inputs(9));
    layer0_outputs(132) <= not((inputs(166)) or (inputs(253)));
    layer0_outputs(133) <= not((inputs(178)) xor (inputs(130)));
    layer0_outputs(134) <= inputs(164);
    layer0_outputs(135) <= not((inputs(222)) xor (inputs(105)));
    layer0_outputs(136) <= not(inputs(229));
    layer0_outputs(137) <= (inputs(3)) or (inputs(32));
    layer0_outputs(138) <= not(inputs(213));
    layer0_outputs(139) <= inputs(233);
    layer0_outputs(140) <= not((inputs(199)) xor (inputs(79)));
    layer0_outputs(141) <= inputs(129);
    layer0_outputs(142) <= not(inputs(82));
    layer0_outputs(143) <= not(inputs(186));
    layer0_outputs(144) <= not(inputs(254));
    layer0_outputs(145) <= (inputs(207)) xor (inputs(227));
    layer0_outputs(146) <= not((inputs(249)) xor (inputs(220)));
    layer0_outputs(147) <= inputs(247);
    layer0_outputs(148) <= not((inputs(68)) or (inputs(129)));
    layer0_outputs(149) <= not((inputs(195)) or (inputs(232)));
    layer0_outputs(150) <= (inputs(108)) xor (inputs(155));
    layer0_outputs(151) <= not(inputs(197)) or (inputs(30));
    layer0_outputs(152) <= not((inputs(6)) and (inputs(155)));
    layer0_outputs(153) <= inputs(148);
    layer0_outputs(154) <= not(inputs(101));
    layer0_outputs(155) <= (inputs(87)) xor (inputs(133));
    layer0_outputs(156) <= not((inputs(177)) or (inputs(247)));
    layer0_outputs(157) <= (inputs(183)) and (inputs(25));
    layer0_outputs(158) <= (inputs(106)) and not (inputs(128));
    layer0_outputs(159) <= not((inputs(154)) xor (inputs(177)));
    layer0_outputs(160) <= not((inputs(190)) xor (inputs(36)));
    layer0_outputs(161) <= (inputs(119)) or (inputs(122));
    layer0_outputs(162) <= not(inputs(235));
    layer0_outputs(163) <= not((inputs(111)) or (inputs(35)));
    layer0_outputs(164) <= (inputs(69)) xor (inputs(49));
    layer0_outputs(165) <= not((inputs(185)) or (inputs(113)));
    layer0_outputs(166) <= not(inputs(133));
    layer0_outputs(167) <= not((inputs(23)) and (inputs(199)));
    layer0_outputs(168) <= (inputs(180)) and not (inputs(96));
    layer0_outputs(169) <= inputs(121);
    layer0_outputs(170) <= not(inputs(255));
    layer0_outputs(171) <= not(inputs(172));
    layer0_outputs(172) <= (inputs(160)) and not (inputs(16));
    layer0_outputs(173) <= inputs(41);
    layer0_outputs(174) <= not(inputs(34)) or (inputs(66));
    layer0_outputs(175) <= not(inputs(225));
    layer0_outputs(176) <= (inputs(125)) xor (inputs(51));
    layer0_outputs(177) <= inputs(230);
    layer0_outputs(178) <= not((inputs(227)) xor (inputs(220)));
    layer0_outputs(179) <= not(inputs(229));
    layer0_outputs(180) <= not(inputs(149));
    layer0_outputs(181) <= (inputs(126)) and not (inputs(252));
    layer0_outputs(182) <= (inputs(168)) or (inputs(71));
    layer0_outputs(183) <= not((inputs(177)) or (inputs(28)));
    layer0_outputs(184) <= inputs(90);
    layer0_outputs(185) <= not(inputs(106)) or (inputs(236));
    layer0_outputs(186) <= not(inputs(234));
    layer0_outputs(187) <= not((inputs(69)) xor (inputs(19)));
    layer0_outputs(188) <= (inputs(153)) and (inputs(168));
    layer0_outputs(189) <= not(inputs(168)) or (inputs(241));
    layer0_outputs(190) <= (inputs(91)) or (inputs(54));
    layer0_outputs(191) <= (inputs(31)) or (inputs(187));
    layer0_outputs(192) <= inputs(210);
    layer0_outputs(193) <= (inputs(60)) xor (inputs(45));
    layer0_outputs(194) <= not(inputs(168)) or (inputs(67));
    layer0_outputs(195) <= (inputs(146)) and not (inputs(90));
    layer0_outputs(196) <= not((inputs(77)) or (inputs(0)));
    layer0_outputs(197) <= inputs(200);
    layer0_outputs(198) <= (inputs(121)) xor (inputs(255));
    layer0_outputs(199) <= not((inputs(161)) or (inputs(77)));
    layer0_outputs(200) <= not(inputs(194));
    layer0_outputs(201) <= not(inputs(122));
    layer0_outputs(202) <= not((inputs(124)) or (inputs(52)));
    layer0_outputs(203) <= not(inputs(140));
    layer0_outputs(204) <= not(inputs(204));
    layer0_outputs(205) <= not(inputs(179));
    layer0_outputs(206) <= (inputs(217)) or (inputs(212));
    layer0_outputs(207) <= (inputs(29)) and not (inputs(143));
    layer0_outputs(208) <= '1';
    layer0_outputs(209) <= (inputs(226)) xor (inputs(21));
    layer0_outputs(210) <= (inputs(247)) and not (inputs(19));
    layer0_outputs(211) <= (inputs(44)) xor (inputs(184));
    layer0_outputs(212) <= inputs(40);
    layer0_outputs(213) <= not(inputs(209)) or (inputs(139));
    layer0_outputs(214) <= inputs(45);
    layer0_outputs(215) <= (inputs(115)) xor (inputs(223));
    layer0_outputs(216) <= (inputs(238)) and not (inputs(13));
    layer0_outputs(217) <= not(inputs(131)) or (inputs(36));
    layer0_outputs(218) <= (inputs(30)) and not (inputs(176));
    layer0_outputs(219) <= not(inputs(121)) or (inputs(159));
    layer0_outputs(220) <= not(inputs(171)) or (inputs(255));
    layer0_outputs(221) <= (inputs(29)) or (inputs(207));
    layer0_outputs(222) <= not((inputs(161)) or (inputs(16)));
    layer0_outputs(223) <= (inputs(46)) xor (inputs(25));
    layer0_outputs(224) <= inputs(98);
    layer0_outputs(225) <= not(inputs(185));
    layer0_outputs(226) <= not(inputs(117));
    layer0_outputs(227) <= not((inputs(1)) or (inputs(100)));
    layer0_outputs(228) <= not(inputs(154));
    layer0_outputs(229) <= (inputs(139)) xor (inputs(101));
    layer0_outputs(230) <= not((inputs(248)) xor (inputs(175)));
    layer0_outputs(231) <= not(inputs(88));
    layer0_outputs(232) <= inputs(162);
    layer0_outputs(233) <= not(inputs(129));
    layer0_outputs(234) <= (inputs(103)) xor (inputs(135));
    layer0_outputs(235) <= not((inputs(173)) and (inputs(188)));
    layer0_outputs(236) <= not(inputs(99)) or (inputs(81));
    layer0_outputs(237) <= inputs(172);
    layer0_outputs(238) <= (inputs(116)) and not (inputs(4));
    layer0_outputs(239) <= (inputs(247)) and not (inputs(166));
    layer0_outputs(240) <= inputs(100);
    layer0_outputs(241) <= not(inputs(223)) or (inputs(40));
    layer0_outputs(242) <= (inputs(170)) or (inputs(133));
    layer0_outputs(243) <= not((inputs(217)) or (inputs(27)));
    layer0_outputs(244) <= (inputs(20)) and (inputs(18));
    layer0_outputs(245) <= (inputs(246)) or (inputs(208));
    layer0_outputs(246) <= not(inputs(174));
    layer0_outputs(247) <= (inputs(195)) xor (inputs(159));
    layer0_outputs(248) <= (inputs(234)) xor (inputs(228));
    layer0_outputs(249) <= not(inputs(59));
    layer0_outputs(250) <= '0';
    layer0_outputs(251) <= not((inputs(211)) and (inputs(45)));
    layer0_outputs(252) <= (inputs(41)) or (inputs(27));
    layer0_outputs(253) <= not((inputs(141)) or (inputs(224)));
    layer0_outputs(254) <= inputs(245);
    layer0_outputs(255) <= not(inputs(220)) or (inputs(10));
    layer0_outputs(256) <= (inputs(21)) and not (inputs(81));
    layer0_outputs(257) <= inputs(6);
    layer0_outputs(258) <= inputs(106);
    layer0_outputs(259) <= (inputs(124)) xor (inputs(103));
    layer0_outputs(260) <= (inputs(167)) or (inputs(174));
    layer0_outputs(261) <= (inputs(187)) and (inputs(126));
    layer0_outputs(262) <= not(inputs(109));
    layer0_outputs(263) <= inputs(8);
    layer0_outputs(264) <= not((inputs(60)) or (inputs(165)));
    layer0_outputs(265) <= (inputs(37)) and (inputs(217));
    layer0_outputs(266) <= (inputs(35)) or (inputs(207));
    layer0_outputs(267) <= inputs(126);
    layer0_outputs(268) <= inputs(127);
    layer0_outputs(269) <= inputs(127);
    layer0_outputs(270) <= (inputs(249)) xor (inputs(42));
    layer0_outputs(271) <= not(inputs(86));
    layer0_outputs(272) <= not(inputs(131)) or (inputs(225));
    layer0_outputs(273) <= (inputs(20)) and not (inputs(44));
    layer0_outputs(274) <= inputs(8);
    layer0_outputs(275) <= not((inputs(69)) xor (inputs(23)));
    layer0_outputs(276) <= not((inputs(244)) or (inputs(225)));
    layer0_outputs(277) <= not(inputs(255)) or (inputs(37));
    layer0_outputs(278) <= not(inputs(196));
    layer0_outputs(279) <= (inputs(132)) xor (inputs(81));
    layer0_outputs(280) <= not(inputs(77));
    layer0_outputs(281) <= inputs(129);
    layer0_outputs(282) <= not((inputs(134)) xor (inputs(164)));
    layer0_outputs(283) <= not(inputs(203));
    layer0_outputs(284) <= not(inputs(179));
    layer0_outputs(285) <= not((inputs(105)) xor (inputs(154)));
    layer0_outputs(286) <= not((inputs(3)) or (inputs(212)));
    layer0_outputs(287) <= inputs(124);
    layer0_outputs(288) <= inputs(31);
    layer0_outputs(289) <= not((inputs(97)) xor (inputs(12)));
    layer0_outputs(290) <= (inputs(79)) or (inputs(134));
    layer0_outputs(291) <= '1';
    layer0_outputs(292) <= (inputs(15)) or (inputs(2));
    layer0_outputs(293) <= (inputs(110)) or (inputs(26));
    layer0_outputs(294) <= (inputs(229)) or (inputs(82));
    layer0_outputs(295) <= not((inputs(216)) xor (inputs(97)));
    layer0_outputs(296) <= not(inputs(131));
    layer0_outputs(297) <= not(inputs(110));
    layer0_outputs(298) <= not((inputs(120)) or (inputs(159)));
    layer0_outputs(299) <= (inputs(38)) and (inputs(87));
    layer0_outputs(300) <= (inputs(207)) and not (inputs(232));
    layer0_outputs(301) <= not(inputs(237));
    layer0_outputs(302) <= not(inputs(15));
    layer0_outputs(303) <= (inputs(74)) and not (inputs(32));
    layer0_outputs(304) <= (inputs(156)) xor (inputs(219));
    layer0_outputs(305) <= not(inputs(114));
    layer0_outputs(306) <= (inputs(200)) and (inputs(198));
    layer0_outputs(307) <= not(inputs(194));
    layer0_outputs(308) <= not(inputs(131));
    layer0_outputs(309) <= not(inputs(98)) or (inputs(49));
    layer0_outputs(310) <= not((inputs(74)) or (inputs(206)));
    layer0_outputs(311) <= (inputs(149)) xor (inputs(31));
    layer0_outputs(312) <= (inputs(172)) and not (inputs(234));
    layer0_outputs(313) <= not((inputs(75)) xor (inputs(96)));
    layer0_outputs(314) <= (inputs(47)) or (inputs(248));
    layer0_outputs(315) <= inputs(161);
    layer0_outputs(316) <= not((inputs(122)) or (inputs(124)));
    layer0_outputs(317) <= not((inputs(232)) and (inputs(5)));
    layer0_outputs(318) <= (inputs(71)) and not (inputs(139));
    layer0_outputs(319) <= (inputs(83)) xor (inputs(161));
    layer0_outputs(320) <= (inputs(40)) and not (inputs(93));
    layer0_outputs(321) <= not((inputs(227)) xor (inputs(8)));
    layer0_outputs(322) <= not((inputs(168)) or (inputs(246)));
    layer0_outputs(323) <= (inputs(189)) xor (inputs(192));
    layer0_outputs(324) <= not(inputs(188));
    layer0_outputs(325) <= not(inputs(149)) or (inputs(45));
    layer0_outputs(326) <= (inputs(195)) and not (inputs(125));
    layer0_outputs(327) <= inputs(74);
    layer0_outputs(328) <= inputs(9);
    layer0_outputs(329) <= not((inputs(185)) or (inputs(76)));
    layer0_outputs(330) <= not((inputs(141)) or (inputs(114)));
    layer0_outputs(331) <= not((inputs(81)) or (inputs(67)));
    layer0_outputs(332) <= not((inputs(150)) or (inputs(132)));
    layer0_outputs(333) <= (inputs(1)) or (inputs(174));
    layer0_outputs(334) <= not((inputs(131)) xor (inputs(188)));
    layer0_outputs(335) <= not((inputs(203)) or (inputs(128)));
    layer0_outputs(336) <= (inputs(103)) and not (inputs(4));
    layer0_outputs(337) <= not(inputs(42));
    layer0_outputs(338) <= not((inputs(255)) or (inputs(163)));
    layer0_outputs(339) <= not((inputs(188)) xor (inputs(136)));
    layer0_outputs(340) <= (inputs(161)) and (inputs(196));
    layer0_outputs(341) <= not((inputs(136)) or (inputs(103)));
    layer0_outputs(342) <= (inputs(224)) xor (inputs(179));
    layer0_outputs(343) <= not(inputs(184)) or (inputs(76));
    layer0_outputs(344) <= (inputs(157)) or (inputs(38));
    layer0_outputs(345) <= (inputs(140)) and not (inputs(94));
    layer0_outputs(346) <= not(inputs(86));
    layer0_outputs(347) <= (inputs(41)) xor (inputs(55));
    layer0_outputs(348) <= not(inputs(27));
    layer0_outputs(349) <= inputs(129);
    layer0_outputs(350) <= inputs(88);
    layer0_outputs(351) <= (inputs(158)) and not (inputs(0));
    layer0_outputs(352) <= inputs(90);
    layer0_outputs(353) <= not(inputs(99));
    layer0_outputs(354) <= (inputs(212)) xor (inputs(226));
    layer0_outputs(355) <= (inputs(42)) and not (inputs(234));
    layer0_outputs(356) <= inputs(198);
    layer0_outputs(357) <= inputs(151);
    layer0_outputs(358) <= inputs(189);
    layer0_outputs(359) <= (inputs(85)) xor (inputs(96));
    layer0_outputs(360) <= not(inputs(71)) or (inputs(136));
    layer0_outputs(361) <= inputs(183);
    layer0_outputs(362) <= (inputs(103)) or (inputs(10));
    layer0_outputs(363) <= not((inputs(137)) and (inputs(196)));
    layer0_outputs(364) <= (inputs(57)) xor (inputs(108));
    layer0_outputs(365) <= (inputs(85)) xor (inputs(86));
    layer0_outputs(366) <= not((inputs(151)) or (inputs(59)));
    layer0_outputs(367) <= not(inputs(85));
    layer0_outputs(368) <= (inputs(149)) or (inputs(206));
    layer0_outputs(369) <= not(inputs(165));
    layer0_outputs(370) <= not((inputs(249)) xor (inputs(201)));
    layer0_outputs(371) <= inputs(157);
    layer0_outputs(372) <= (inputs(221)) xor (inputs(112));
    layer0_outputs(373) <= (inputs(198)) xor (inputs(245));
    layer0_outputs(374) <= (inputs(101)) xor (inputs(39));
    layer0_outputs(375) <= inputs(24);
    layer0_outputs(376) <= not(inputs(173)) or (inputs(125));
    layer0_outputs(377) <= not((inputs(144)) or (inputs(78)));
    layer0_outputs(378) <= (inputs(11)) xor (inputs(174));
    layer0_outputs(379) <= inputs(71);
    layer0_outputs(380) <= not((inputs(156)) or (inputs(68)));
    layer0_outputs(381) <= not((inputs(187)) xor (inputs(19)));
    layer0_outputs(382) <= not(inputs(141));
    layer0_outputs(383) <= not(inputs(26));
    layer0_outputs(384) <= (inputs(196)) or (inputs(99));
    layer0_outputs(385) <= (inputs(144)) or (inputs(212));
    layer0_outputs(386) <= (inputs(80)) and not (inputs(144));
    layer0_outputs(387) <= not((inputs(33)) xor (inputs(192)));
    layer0_outputs(388) <= not((inputs(84)) or (inputs(160)));
    layer0_outputs(389) <= not(inputs(6));
    layer0_outputs(390) <= not(inputs(206));
    layer0_outputs(391) <= '0';
    layer0_outputs(392) <= inputs(87);
    layer0_outputs(393) <= not((inputs(126)) xor (inputs(92)));
    layer0_outputs(394) <= not(inputs(144));
    layer0_outputs(395) <= (inputs(157)) xor (inputs(16));
    layer0_outputs(396) <= inputs(221);
    layer0_outputs(397) <= (inputs(51)) xor (inputs(92));
    layer0_outputs(398) <= (inputs(246)) or (inputs(8));
    layer0_outputs(399) <= inputs(113);
    layer0_outputs(400) <= inputs(40);
    layer0_outputs(401) <= not((inputs(47)) or (inputs(23)));
    layer0_outputs(402) <= not(inputs(228)) or (inputs(97));
    layer0_outputs(403) <= not((inputs(100)) or (inputs(87)));
    layer0_outputs(404) <= not(inputs(249));
    layer0_outputs(405) <= not(inputs(163));
    layer0_outputs(406) <= (inputs(55)) or (inputs(208));
    layer0_outputs(407) <= inputs(215);
    layer0_outputs(408) <= inputs(56);
    layer0_outputs(409) <= (inputs(101)) and not (inputs(176));
    layer0_outputs(410) <= not((inputs(240)) and (inputs(96)));
    layer0_outputs(411) <= inputs(242);
    layer0_outputs(412) <= inputs(255);
    layer0_outputs(413) <= (inputs(89)) and not (inputs(225));
    layer0_outputs(414) <= (inputs(162)) and not (inputs(189));
    layer0_outputs(415) <= not((inputs(76)) or (inputs(21)));
    layer0_outputs(416) <= (inputs(35)) or (inputs(110));
    layer0_outputs(417) <= not((inputs(153)) and (inputs(46)));
    layer0_outputs(418) <= (inputs(204)) or (inputs(46));
    layer0_outputs(419) <= (inputs(41)) or (inputs(205));
    layer0_outputs(420) <= (inputs(65)) xor (inputs(21));
    layer0_outputs(421) <= (inputs(150)) or (inputs(76));
    layer0_outputs(422) <= not(inputs(40)) or (inputs(205));
    layer0_outputs(423) <= (inputs(173)) and not (inputs(32));
    layer0_outputs(424) <= (inputs(171)) xor (inputs(140));
    layer0_outputs(425) <= not(inputs(135)) or (inputs(251));
    layer0_outputs(426) <= inputs(53);
    layer0_outputs(427) <= not(inputs(80));
    layer0_outputs(428) <= (inputs(20)) xor (inputs(134));
    layer0_outputs(429) <= (inputs(114)) or (inputs(83));
    layer0_outputs(430) <= inputs(165);
    layer0_outputs(431) <= not((inputs(96)) xor (inputs(11)));
    layer0_outputs(432) <= not((inputs(144)) and (inputs(210)));
    layer0_outputs(433) <= (inputs(193)) or (inputs(0));
    layer0_outputs(434) <= not(inputs(171));
    layer0_outputs(435) <= (inputs(218)) and (inputs(38));
    layer0_outputs(436) <= (inputs(172)) and not (inputs(217));
    layer0_outputs(437) <= not(inputs(75)) or (inputs(253));
    layer0_outputs(438) <= (inputs(27)) or (inputs(115));
    layer0_outputs(439) <= (inputs(193)) or (inputs(178));
    layer0_outputs(440) <= (inputs(222)) or (inputs(220));
    layer0_outputs(441) <= not((inputs(186)) or (inputs(12)));
    layer0_outputs(442) <= inputs(142);
    layer0_outputs(443) <= not(inputs(177));
    layer0_outputs(444) <= not((inputs(211)) and (inputs(90)));
    layer0_outputs(445) <= inputs(2);
    layer0_outputs(446) <= not(inputs(36));
    layer0_outputs(447) <= (inputs(171)) xor (inputs(23));
    layer0_outputs(448) <= not(inputs(82));
    layer0_outputs(449) <= (inputs(228)) and not (inputs(17));
    layer0_outputs(450) <= (inputs(58)) xor (inputs(26));
    layer0_outputs(451) <= not((inputs(103)) or (inputs(208)));
    layer0_outputs(452) <= inputs(85);
    layer0_outputs(453) <= (inputs(42)) xor (inputs(86));
    layer0_outputs(454) <= not((inputs(153)) or (inputs(154)));
    layer0_outputs(455) <= (inputs(168)) or (inputs(11));
    layer0_outputs(456) <= not(inputs(91));
    layer0_outputs(457) <= inputs(184);
    layer0_outputs(458) <= not(inputs(138));
    layer0_outputs(459) <= not(inputs(157));
    layer0_outputs(460) <= not((inputs(72)) or (inputs(95)));
    layer0_outputs(461) <= not(inputs(74)) or (inputs(67));
    layer0_outputs(462) <= (inputs(153)) xor (inputs(166));
    layer0_outputs(463) <= not((inputs(114)) or (inputs(89)));
    layer0_outputs(464) <= not(inputs(198)) or (inputs(60));
    layer0_outputs(465) <= inputs(231);
    layer0_outputs(466) <= inputs(241);
    layer0_outputs(467) <= inputs(153);
    layer0_outputs(468) <= not((inputs(45)) xor (inputs(78)));
    layer0_outputs(469) <= (inputs(146)) and not (inputs(61));
    layer0_outputs(470) <= not(inputs(110));
    layer0_outputs(471) <= (inputs(117)) or (inputs(145));
    layer0_outputs(472) <= not((inputs(237)) or (inputs(88)));
    layer0_outputs(473) <= inputs(20);
    layer0_outputs(474) <= not(inputs(44));
    layer0_outputs(475) <= not((inputs(212)) xor (inputs(138)));
    layer0_outputs(476) <= not((inputs(38)) xor (inputs(181)));
    layer0_outputs(477) <= (inputs(63)) or (inputs(39));
    layer0_outputs(478) <= (inputs(170)) or (inputs(188));
    layer0_outputs(479) <= not(inputs(197));
    layer0_outputs(480) <= (inputs(10)) or (inputs(182));
    layer0_outputs(481) <= (inputs(136)) and (inputs(222));
    layer0_outputs(482) <= not((inputs(203)) xor (inputs(172)));
    layer0_outputs(483) <= (inputs(18)) and not (inputs(193));
    layer0_outputs(484) <= (inputs(47)) xor (inputs(203));
    layer0_outputs(485) <= not((inputs(132)) xor (inputs(146)));
    layer0_outputs(486) <= not(inputs(146)) or (inputs(72));
    layer0_outputs(487) <= inputs(40);
    layer0_outputs(488) <= not((inputs(34)) or (inputs(169)));
    layer0_outputs(489) <= not((inputs(154)) xor (inputs(81)));
    layer0_outputs(490) <= not((inputs(187)) xor (inputs(131)));
    layer0_outputs(491) <= not(inputs(232));
    layer0_outputs(492) <= (inputs(213)) and not (inputs(156));
    layer0_outputs(493) <= not((inputs(97)) or (inputs(98)));
    layer0_outputs(494) <= (inputs(26)) and (inputs(149));
    layer0_outputs(495) <= not(inputs(102)) or (inputs(163));
    layer0_outputs(496) <= not((inputs(139)) or (inputs(69)));
    layer0_outputs(497) <= inputs(26);
    layer0_outputs(498) <= not(inputs(163)) or (inputs(109));
    layer0_outputs(499) <= not(inputs(171)) or (inputs(18));
    layer0_outputs(500) <= not((inputs(117)) xor (inputs(70)));
    layer0_outputs(501) <= (inputs(66)) xor (inputs(132));
    layer0_outputs(502) <= not((inputs(164)) or (inputs(82)));
    layer0_outputs(503) <= not(inputs(172)) or (inputs(25));
    layer0_outputs(504) <= (inputs(62)) xor (inputs(140));
    layer0_outputs(505) <= (inputs(226)) or (inputs(175));
    layer0_outputs(506) <= (inputs(61)) or (inputs(216));
    layer0_outputs(507) <= (inputs(46)) or (inputs(25));
    layer0_outputs(508) <= inputs(114);
    layer0_outputs(509) <= inputs(104);
    layer0_outputs(510) <= not((inputs(109)) or (inputs(42)));
    layer0_outputs(511) <= not((inputs(74)) or (inputs(132)));
    layer0_outputs(512) <= not(inputs(55)) or (inputs(226));
    layer0_outputs(513) <= not((inputs(125)) xor (inputs(108)));
    layer0_outputs(514) <= (inputs(141)) xor (inputs(192));
    layer0_outputs(515) <= inputs(174);
    layer0_outputs(516) <= not((inputs(116)) xor (inputs(102)));
    layer0_outputs(517) <= not(inputs(214));
    layer0_outputs(518) <= not((inputs(255)) and (inputs(183)));
    layer0_outputs(519) <= (inputs(56)) and (inputs(189));
    layer0_outputs(520) <= not((inputs(227)) or (inputs(216)));
    layer0_outputs(521) <= not(inputs(40));
    layer0_outputs(522) <= inputs(113);
    layer0_outputs(523) <= not((inputs(27)) and (inputs(19)));
    layer0_outputs(524) <= not(inputs(69));
    layer0_outputs(525) <= not((inputs(130)) or (inputs(204)));
    layer0_outputs(526) <= not(inputs(132));
    layer0_outputs(527) <= not((inputs(245)) xor (inputs(224)));
    layer0_outputs(528) <= inputs(35);
    layer0_outputs(529) <= not(inputs(144)) or (inputs(0));
    layer0_outputs(530) <= not(inputs(156));
    layer0_outputs(531) <= (inputs(157)) xor (inputs(101));
    layer0_outputs(532) <= (inputs(223)) xor (inputs(54));
    layer0_outputs(533) <= (inputs(220)) and not (inputs(29));
    layer0_outputs(534) <= not((inputs(192)) or (inputs(248)));
    layer0_outputs(535) <= not((inputs(168)) xor (inputs(86)));
    layer0_outputs(536) <= (inputs(224)) xor (inputs(205));
    layer0_outputs(537) <= (inputs(248)) and not (inputs(50));
    layer0_outputs(538) <= (inputs(69)) or (inputs(125));
    layer0_outputs(539) <= (inputs(228)) or (inputs(148));
    layer0_outputs(540) <= not(inputs(71)) or (inputs(138));
    layer0_outputs(541) <= not((inputs(95)) xor (inputs(65)));
    layer0_outputs(542) <= not(inputs(155));
    layer0_outputs(543) <= not((inputs(58)) xor (inputs(111)));
    layer0_outputs(544) <= '1';
    layer0_outputs(545) <= (inputs(179)) and not (inputs(14));
    layer0_outputs(546) <= not((inputs(126)) or (inputs(144)));
    layer0_outputs(547) <= inputs(3);
    layer0_outputs(548) <= (inputs(184)) and not (inputs(132));
    layer0_outputs(549) <= not(inputs(150)) or (inputs(96));
    layer0_outputs(550) <= (inputs(103)) and not (inputs(1));
    layer0_outputs(551) <= '1';
    layer0_outputs(552) <= not(inputs(229));
    layer0_outputs(553) <= (inputs(174)) xor (inputs(68));
    layer0_outputs(554) <= not(inputs(185)) or (inputs(118));
    layer0_outputs(555) <= (inputs(194)) or (inputs(88));
    layer0_outputs(556) <= (inputs(35)) xor (inputs(122));
    layer0_outputs(557) <= (inputs(26)) or (inputs(173));
    layer0_outputs(558) <= inputs(198);
    layer0_outputs(559) <= inputs(116);
    layer0_outputs(560) <= not(inputs(151));
    layer0_outputs(561) <= (inputs(42)) and not (inputs(145));
    layer0_outputs(562) <= not((inputs(9)) xor (inputs(222)));
    layer0_outputs(563) <= inputs(213);
    layer0_outputs(564) <= inputs(38);
    layer0_outputs(565) <= inputs(233);
    layer0_outputs(566) <= not(inputs(95)) or (inputs(13));
    layer0_outputs(567) <= not((inputs(92)) or (inputs(96)));
    layer0_outputs(568) <= not((inputs(234)) or (inputs(241)));
    layer0_outputs(569) <= (inputs(244)) and not (inputs(60));
    layer0_outputs(570) <= not((inputs(253)) or (inputs(147)));
    layer0_outputs(571) <= not((inputs(182)) or (inputs(160)));
    layer0_outputs(572) <= not(inputs(42)) or (inputs(112));
    layer0_outputs(573) <= (inputs(140)) and not (inputs(14));
    layer0_outputs(574) <= not((inputs(196)) xor (inputs(237)));
    layer0_outputs(575) <= not((inputs(174)) xor (inputs(176)));
    layer0_outputs(576) <= inputs(95);
    layer0_outputs(577) <= (inputs(77)) and not (inputs(13));
    layer0_outputs(578) <= not((inputs(64)) or (inputs(11)));
    layer0_outputs(579) <= not(inputs(44)) or (inputs(108));
    layer0_outputs(580) <= not(inputs(106));
    layer0_outputs(581) <= not((inputs(116)) xor (inputs(36)));
    layer0_outputs(582) <= not(inputs(120));
    layer0_outputs(583) <= (inputs(224)) xor (inputs(252));
    layer0_outputs(584) <= not((inputs(255)) and (inputs(13)));
    layer0_outputs(585) <= (inputs(50)) or (inputs(88));
    layer0_outputs(586) <= not((inputs(185)) or (inputs(217)));
    layer0_outputs(587) <= not(inputs(41));
    layer0_outputs(588) <= not((inputs(39)) and (inputs(186)));
    layer0_outputs(589) <= (inputs(68)) and not (inputs(119));
    layer0_outputs(590) <= not(inputs(200));
    layer0_outputs(591) <= not(inputs(224));
    layer0_outputs(592) <= inputs(214);
    layer0_outputs(593) <= (inputs(235)) or (inputs(216));
    layer0_outputs(594) <= (inputs(88)) xor (inputs(57));
    layer0_outputs(595) <= (inputs(90)) and not (inputs(144));
    layer0_outputs(596) <= not((inputs(117)) xor (inputs(124)));
    layer0_outputs(597) <= not((inputs(85)) xor (inputs(177)));
    layer0_outputs(598) <= not((inputs(222)) or (inputs(82)));
    layer0_outputs(599) <= not(inputs(88));
    layer0_outputs(600) <= (inputs(105)) or (inputs(239));
    layer0_outputs(601) <= not((inputs(181)) xor (inputs(164)));
    layer0_outputs(602) <= (inputs(250)) and not (inputs(222));
    layer0_outputs(603) <= inputs(228);
    layer0_outputs(604) <= inputs(57);
    layer0_outputs(605) <= (inputs(135)) xor (inputs(183));
    layer0_outputs(606) <= not((inputs(210)) and (inputs(203)));
    layer0_outputs(607) <= inputs(114);
    layer0_outputs(608) <= not(inputs(28)) or (inputs(68));
    layer0_outputs(609) <= (inputs(161)) or (inputs(170));
    layer0_outputs(610) <= (inputs(1)) or (inputs(189));
    layer0_outputs(611) <= not(inputs(215)) or (inputs(97));
    layer0_outputs(612) <= (inputs(165)) xor (inputs(151));
    layer0_outputs(613) <= not(inputs(145));
    layer0_outputs(614) <= not((inputs(85)) and (inputs(217)));
    layer0_outputs(615) <= inputs(225);
    layer0_outputs(616) <= inputs(209);
    layer0_outputs(617) <= not(inputs(139));
    layer0_outputs(618) <= not((inputs(17)) or (inputs(21)));
    layer0_outputs(619) <= not((inputs(145)) xor (inputs(100)));
    layer0_outputs(620) <= not((inputs(74)) or (inputs(138)));
    layer0_outputs(621) <= not(inputs(232));
    layer0_outputs(622) <= not(inputs(66));
    layer0_outputs(623) <= inputs(159);
    layer0_outputs(624) <= (inputs(225)) or (inputs(194));
    layer0_outputs(625) <= (inputs(40)) xor (inputs(92));
    layer0_outputs(626) <= not(inputs(189));
    layer0_outputs(627) <= not(inputs(210));
    layer0_outputs(628) <= not(inputs(249)) or (inputs(112));
    layer0_outputs(629) <= inputs(161);
    layer0_outputs(630) <= (inputs(153)) and not (inputs(193));
    layer0_outputs(631) <= (inputs(73)) xor (inputs(214));
    layer0_outputs(632) <= (inputs(224)) xor (inputs(209));
    layer0_outputs(633) <= not((inputs(1)) xor (inputs(139)));
    layer0_outputs(634) <= (inputs(143)) or (inputs(233));
    layer0_outputs(635) <= not(inputs(166));
    layer0_outputs(636) <= (inputs(71)) and not (inputs(140));
    layer0_outputs(637) <= inputs(91);
    layer0_outputs(638) <= not(inputs(34));
    layer0_outputs(639) <= not(inputs(179));
    layer0_outputs(640) <= (inputs(118)) or (inputs(88));
    layer0_outputs(641) <= inputs(98);
    layer0_outputs(642) <= not(inputs(249));
    layer0_outputs(643) <= not(inputs(160));
    layer0_outputs(644) <= inputs(55);
    layer0_outputs(645) <= (inputs(114)) or (inputs(59));
    layer0_outputs(646) <= inputs(85);
    layer0_outputs(647) <= not((inputs(254)) or (inputs(128)));
    layer0_outputs(648) <= (inputs(219)) xor (inputs(211));
    layer0_outputs(649) <= inputs(144);
    layer0_outputs(650) <= not((inputs(162)) or (inputs(113)));
    layer0_outputs(651) <= not(inputs(141)) or (inputs(215));
    layer0_outputs(652) <= not(inputs(104));
    layer0_outputs(653) <= (inputs(2)) or (inputs(6));
    layer0_outputs(654) <= not(inputs(209)) or (inputs(252));
    layer0_outputs(655) <= not(inputs(20));
    layer0_outputs(656) <= not((inputs(24)) or (inputs(21)));
    layer0_outputs(657) <= (inputs(108)) or (inputs(152));
    layer0_outputs(658) <= not((inputs(19)) or (inputs(113)));
    layer0_outputs(659) <= (inputs(240)) and not (inputs(63));
    layer0_outputs(660) <= not(inputs(25));
    layer0_outputs(661) <= (inputs(216)) or (inputs(143));
    layer0_outputs(662) <= not(inputs(241)) or (inputs(223));
    layer0_outputs(663) <= not(inputs(163));
    layer0_outputs(664) <= not(inputs(52));
    layer0_outputs(665) <= not(inputs(200));
    layer0_outputs(666) <= inputs(245);
    layer0_outputs(667) <= (inputs(15)) xor (inputs(170));
    layer0_outputs(668) <= not((inputs(43)) or (inputs(111)));
    layer0_outputs(669) <= (inputs(180)) xor (inputs(27));
    layer0_outputs(670) <= not(inputs(45)) or (inputs(162));
    layer0_outputs(671) <= not(inputs(104));
    layer0_outputs(672) <= (inputs(159)) xor (inputs(197));
    layer0_outputs(673) <= (inputs(100)) and not (inputs(252));
    layer0_outputs(674) <= (inputs(67)) xor (inputs(157));
    layer0_outputs(675) <= (inputs(213)) and not (inputs(243));
    layer0_outputs(676) <= (inputs(169)) xor (inputs(221));
    layer0_outputs(677) <= not((inputs(192)) or (inputs(159)));
    layer0_outputs(678) <= (inputs(198)) or (inputs(33));
    layer0_outputs(679) <= (inputs(109)) or (inputs(251));
    layer0_outputs(680) <= (inputs(194)) and not (inputs(61));
    layer0_outputs(681) <= (inputs(145)) xor (inputs(229));
    layer0_outputs(682) <= not((inputs(150)) or (inputs(166)));
    layer0_outputs(683) <= not(inputs(93));
    layer0_outputs(684) <= not(inputs(101)) or (inputs(191));
    layer0_outputs(685) <= (inputs(62)) xor (inputs(89));
    layer0_outputs(686) <= (inputs(23)) or (inputs(186));
    layer0_outputs(687) <= not((inputs(16)) and (inputs(92)));
    layer0_outputs(688) <= (inputs(190)) or (inputs(76));
    layer0_outputs(689) <= '0';
    layer0_outputs(690) <= not(inputs(232)) or (inputs(118));
    layer0_outputs(691) <= (inputs(255)) xor (inputs(109));
    layer0_outputs(692) <= inputs(228);
    layer0_outputs(693) <= not((inputs(35)) xor (inputs(4)));
    layer0_outputs(694) <= not(inputs(98)) or (inputs(126));
    layer0_outputs(695) <= inputs(95);
    layer0_outputs(696) <= (inputs(10)) or (inputs(213));
    layer0_outputs(697) <= not((inputs(110)) or (inputs(72)));
    layer0_outputs(698) <= (inputs(205)) and (inputs(130));
    layer0_outputs(699) <= (inputs(8)) xor (inputs(194));
    layer0_outputs(700) <= not((inputs(115)) or (inputs(47)));
    layer0_outputs(701) <= not((inputs(208)) or (inputs(229)));
    layer0_outputs(702) <= (inputs(174)) xor (inputs(64));
    layer0_outputs(703) <= (inputs(141)) or (inputs(150));
    layer0_outputs(704) <= not((inputs(1)) or (inputs(58)));
    layer0_outputs(705) <= (inputs(100)) and not (inputs(173));
    layer0_outputs(706) <= not((inputs(35)) or (inputs(18)));
    layer0_outputs(707) <= not((inputs(249)) or (inputs(253)));
    layer0_outputs(708) <= (inputs(97)) or (inputs(140));
    layer0_outputs(709) <= '0';
    layer0_outputs(710) <= (inputs(209)) or (inputs(254));
    layer0_outputs(711) <= not(inputs(216));
    layer0_outputs(712) <= inputs(229);
    layer0_outputs(713) <= not(inputs(227)) or (inputs(82));
    layer0_outputs(714) <= '1';
    layer0_outputs(715) <= (inputs(104)) and not (inputs(204));
    layer0_outputs(716) <= (inputs(179)) or (inputs(141));
    layer0_outputs(717) <= not((inputs(94)) or (inputs(90)));
    layer0_outputs(718) <= (inputs(171)) xor (inputs(125));
    layer0_outputs(719) <= not(inputs(213));
    layer0_outputs(720) <= inputs(29);
    layer0_outputs(721) <= (inputs(198)) or (inputs(84));
    layer0_outputs(722) <= (inputs(16)) or (inputs(2));
    layer0_outputs(723) <= not((inputs(253)) xor (inputs(145)));
    layer0_outputs(724) <= not((inputs(176)) and (inputs(198)));
    layer0_outputs(725) <= not(inputs(20));
    layer0_outputs(726) <= (inputs(209)) xor (inputs(230));
    layer0_outputs(727) <= not(inputs(68)) or (inputs(175));
    layer0_outputs(728) <= not((inputs(251)) or (inputs(212)));
    layer0_outputs(729) <= inputs(40);
    layer0_outputs(730) <= not(inputs(231));
    layer0_outputs(731) <= not(inputs(38));
    layer0_outputs(732) <= '0';
    layer0_outputs(733) <= (inputs(181)) and not (inputs(67));
    layer0_outputs(734) <= inputs(146);
    layer0_outputs(735) <= not(inputs(23));
    layer0_outputs(736) <= (inputs(232)) and not (inputs(26));
    layer0_outputs(737) <= not((inputs(166)) or (inputs(32)));
    layer0_outputs(738) <= not(inputs(189)) or (inputs(121));
    layer0_outputs(739) <= (inputs(135)) and not (inputs(73));
    layer0_outputs(740) <= not((inputs(228)) and (inputs(30)));
    layer0_outputs(741) <= not(inputs(26));
    layer0_outputs(742) <= (inputs(47)) and not (inputs(12));
    layer0_outputs(743) <= (inputs(173)) xor (inputs(141));
    layer0_outputs(744) <= not(inputs(222)) or (inputs(97));
    layer0_outputs(745) <= (inputs(235)) xor (inputs(159));
    layer0_outputs(746) <= (inputs(156)) xor (inputs(116));
    layer0_outputs(747) <= not((inputs(130)) or (inputs(158)));
    layer0_outputs(748) <= (inputs(117)) and not (inputs(206));
    layer0_outputs(749) <= not(inputs(247)) or (inputs(137));
    layer0_outputs(750) <= inputs(42);
    layer0_outputs(751) <= inputs(199);
    layer0_outputs(752) <= (inputs(71)) or (inputs(225));
    layer0_outputs(753) <= not((inputs(116)) xor (inputs(50)));
    layer0_outputs(754) <= not((inputs(40)) or (inputs(120)));
    layer0_outputs(755) <= not((inputs(151)) xor (inputs(131)));
    layer0_outputs(756) <= not(inputs(155));
    layer0_outputs(757) <= '1';
    layer0_outputs(758) <= inputs(186);
    layer0_outputs(759) <= not(inputs(178));
    layer0_outputs(760) <= (inputs(3)) and not (inputs(194));
    layer0_outputs(761) <= not((inputs(22)) xor (inputs(57)));
    layer0_outputs(762) <= (inputs(237)) or (inputs(166));
    layer0_outputs(763) <= (inputs(249)) or (inputs(157));
    layer0_outputs(764) <= (inputs(53)) and not (inputs(174));
    layer0_outputs(765) <= not((inputs(27)) and (inputs(215)));
    layer0_outputs(766) <= (inputs(250)) or (inputs(213));
    layer0_outputs(767) <= not(inputs(87));
    layer0_outputs(768) <= not(inputs(231));
    layer0_outputs(769) <= inputs(230);
    layer0_outputs(770) <= not(inputs(120));
    layer0_outputs(771) <= inputs(232);
    layer0_outputs(772) <= (inputs(33)) xor (inputs(151));
    layer0_outputs(773) <= inputs(228);
    layer0_outputs(774) <= not(inputs(75));
    layer0_outputs(775) <= not(inputs(100));
    layer0_outputs(776) <= not((inputs(115)) xor (inputs(103)));
    layer0_outputs(777) <= not((inputs(121)) xor (inputs(100)));
    layer0_outputs(778) <= inputs(174);
    layer0_outputs(779) <= (inputs(185)) or (inputs(6));
    layer0_outputs(780) <= not(inputs(70)) or (inputs(174));
    layer0_outputs(781) <= (inputs(213)) xor (inputs(248));
    layer0_outputs(782) <= (inputs(202)) xor (inputs(251));
    layer0_outputs(783) <= not(inputs(150)) or (inputs(219));
    layer0_outputs(784) <= not(inputs(26));
    layer0_outputs(785) <= not(inputs(184));
    layer0_outputs(786) <= not((inputs(45)) or (inputs(76)));
    layer0_outputs(787) <= not((inputs(78)) or (inputs(96)));
    layer0_outputs(788) <= not((inputs(45)) or (inputs(78)));
    layer0_outputs(789) <= not(inputs(38)) or (inputs(137));
    layer0_outputs(790) <= (inputs(125)) xor (inputs(94));
    layer0_outputs(791) <= (inputs(206)) and not (inputs(100));
    layer0_outputs(792) <= inputs(86);
    layer0_outputs(793) <= not(inputs(119)) or (inputs(178));
    layer0_outputs(794) <= (inputs(47)) and not (inputs(124));
    layer0_outputs(795) <= inputs(167);
    layer0_outputs(796) <= inputs(59);
    layer0_outputs(797) <= not((inputs(116)) xor (inputs(147)));
    layer0_outputs(798) <= not(inputs(195)) or (inputs(94));
    layer0_outputs(799) <= not(inputs(188));
    layer0_outputs(800) <= not(inputs(193));
    layer0_outputs(801) <= not(inputs(235));
    layer0_outputs(802) <= inputs(22);
    layer0_outputs(803) <= not(inputs(151)) or (inputs(53));
    layer0_outputs(804) <= (inputs(58)) xor (inputs(17));
    layer0_outputs(805) <= (inputs(196)) or (inputs(192));
    layer0_outputs(806) <= (inputs(38)) xor (inputs(89));
    layer0_outputs(807) <= not((inputs(62)) xor (inputs(212)));
    layer0_outputs(808) <= not(inputs(81)) or (inputs(185));
    layer0_outputs(809) <= (inputs(5)) xor (inputs(61));
    layer0_outputs(810) <= not(inputs(1));
    layer0_outputs(811) <= not((inputs(243)) or (inputs(118)));
    layer0_outputs(812) <= (inputs(90)) and (inputs(37));
    layer0_outputs(813) <= not((inputs(87)) or (inputs(72)));
    layer0_outputs(814) <= inputs(9);
    layer0_outputs(815) <= not(inputs(171));
    layer0_outputs(816) <= not((inputs(220)) and (inputs(213)));
    layer0_outputs(817) <= not((inputs(237)) xor (inputs(150)));
    layer0_outputs(818) <= not((inputs(229)) xor (inputs(50)));
    layer0_outputs(819) <= (inputs(214)) and (inputs(107));
    layer0_outputs(820) <= (inputs(253)) or (inputs(67));
    layer0_outputs(821) <= (inputs(24)) xor (inputs(70));
    layer0_outputs(822) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(823) <= '1';
    layer0_outputs(824) <= (inputs(65)) and not (inputs(91));
    layer0_outputs(825) <= not((inputs(149)) xor (inputs(197)));
    layer0_outputs(826) <= (inputs(27)) and not (inputs(141));
    layer0_outputs(827) <= (inputs(184)) or (inputs(125));
    layer0_outputs(828) <= not((inputs(228)) or (inputs(34)));
    layer0_outputs(829) <= not((inputs(196)) xor (inputs(208)));
    layer0_outputs(830) <= not(inputs(25));
    layer0_outputs(831) <= not(inputs(214));
    layer0_outputs(832) <= not(inputs(152));
    layer0_outputs(833) <= (inputs(84)) and not (inputs(247));
    layer0_outputs(834) <= (inputs(107)) or (inputs(60));
    layer0_outputs(835) <= (inputs(189)) xor (inputs(34));
    layer0_outputs(836) <= not((inputs(238)) xor (inputs(143)));
    layer0_outputs(837) <= (inputs(231)) and not (inputs(38));
    layer0_outputs(838) <= inputs(66);
    layer0_outputs(839) <= not(inputs(114));
    layer0_outputs(840) <= not((inputs(15)) or (inputs(160)));
    layer0_outputs(841) <= not(inputs(89));
    layer0_outputs(842) <= not((inputs(92)) and (inputs(44)));
    layer0_outputs(843) <= (inputs(29)) xor (inputs(129));
    layer0_outputs(844) <= inputs(93);
    layer0_outputs(845) <= not((inputs(41)) or (inputs(6)));
    layer0_outputs(846) <= not((inputs(26)) and (inputs(101)));
    layer0_outputs(847) <= not((inputs(101)) xor (inputs(165)));
    layer0_outputs(848) <= (inputs(156)) xor (inputs(62));
    layer0_outputs(849) <= not(inputs(105));
    layer0_outputs(850) <= (inputs(48)) and (inputs(193));
    layer0_outputs(851) <= (inputs(52)) and not (inputs(207));
    layer0_outputs(852) <= (inputs(22)) or (inputs(255));
    layer0_outputs(853) <= (inputs(65)) or (inputs(12));
    layer0_outputs(854) <= (inputs(217)) or (inputs(187));
    layer0_outputs(855) <= not((inputs(19)) xor (inputs(92)));
    layer0_outputs(856) <= (inputs(56)) xor (inputs(1));
    layer0_outputs(857) <= inputs(120);
    layer0_outputs(858) <= not(inputs(242)) or (inputs(35));
    layer0_outputs(859) <= (inputs(18)) or (inputs(2));
    layer0_outputs(860) <= not(inputs(209));
    layer0_outputs(861) <= (inputs(123)) or (inputs(168));
    layer0_outputs(862) <= not(inputs(114));
    layer0_outputs(863) <= not((inputs(121)) xor (inputs(202)));
    layer0_outputs(864) <= not(inputs(89)) or (inputs(68));
    layer0_outputs(865) <= '1';
    layer0_outputs(866) <= (inputs(169)) or (inputs(83));
    layer0_outputs(867) <= not(inputs(192)) or (inputs(234));
    layer0_outputs(868) <= (inputs(218)) and (inputs(117));
    layer0_outputs(869) <= not(inputs(191)) or (inputs(112));
    layer0_outputs(870) <= (inputs(80)) and not (inputs(47));
    layer0_outputs(871) <= (inputs(103)) xor (inputs(31));
    layer0_outputs(872) <= (inputs(64)) or (inputs(22));
    layer0_outputs(873) <= (inputs(202)) and not (inputs(136));
    layer0_outputs(874) <= not(inputs(211));
    layer0_outputs(875) <= (inputs(157)) xor (inputs(223));
    layer0_outputs(876) <= inputs(88);
    layer0_outputs(877) <= not((inputs(233)) xor (inputs(95)));
    layer0_outputs(878) <= (inputs(142)) and (inputs(143));
    layer0_outputs(879) <= (inputs(152)) or (inputs(121));
    layer0_outputs(880) <= not(inputs(108));
    layer0_outputs(881) <= inputs(45);
    layer0_outputs(882) <= not(inputs(179)) or (inputs(57));
    layer0_outputs(883) <= not((inputs(208)) or (inputs(116)));
    layer0_outputs(884) <= inputs(142);
    layer0_outputs(885) <= (inputs(133)) and not (inputs(65));
    layer0_outputs(886) <= inputs(233);
    layer0_outputs(887) <= not((inputs(138)) and (inputs(83)));
    layer0_outputs(888) <= (inputs(237)) or (inputs(220));
    layer0_outputs(889) <= not(inputs(54)) or (inputs(216));
    layer0_outputs(890) <= inputs(55);
    layer0_outputs(891) <= inputs(104);
    layer0_outputs(892) <= not((inputs(220)) or (inputs(38)));
    layer0_outputs(893) <= not((inputs(206)) xor (inputs(28)));
    layer0_outputs(894) <= not((inputs(80)) and (inputs(205)));
    layer0_outputs(895) <= (inputs(197)) and not (inputs(131));
    layer0_outputs(896) <= not(inputs(253)) or (inputs(175));
    layer0_outputs(897) <= not((inputs(82)) xor (inputs(5)));
    layer0_outputs(898) <= not((inputs(241)) or (inputs(237)));
    layer0_outputs(899) <= (inputs(147)) or (inputs(196));
    layer0_outputs(900) <= inputs(43);
    layer0_outputs(901) <= (inputs(126)) and not (inputs(226));
    layer0_outputs(902) <= not(inputs(131)) or (inputs(126));
    layer0_outputs(903) <= not((inputs(5)) xor (inputs(39)));
    layer0_outputs(904) <= (inputs(7)) and not (inputs(184));
    layer0_outputs(905) <= (inputs(174)) or (inputs(230));
    layer0_outputs(906) <= (inputs(209)) or (inputs(160));
    layer0_outputs(907) <= inputs(59);
    layer0_outputs(908) <= not((inputs(251)) or (inputs(93)));
    layer0_outputs(909) <= inputs(237);
    layer0_outputs(910) <= not(inputs(168));
    layer0_outputs(911) <= not((inputs(248)) or (inputs(61)));
    layer0_outputs(912) <= inputs(129);
    layer0_outputs(913) <= (inputs(199)) and not (inputs(60));
    layer0_outputs(914) <= (inputs(105)) xor (inputs(16));
    layer0_outputs(915) <= not((inputs(190)) or (inputs(177)));
    layer0_outputs(916) <= (inputs(155)) and not (inputs(106));
    layer0_outputs(917) <= not(inputs(76));
    layer0_outputs(918) <= not((inputs(212)) or (inputs(96)));
    layer0_outputs(919) <= not((inputs(143)) or (inputs(195)));
    layer0_outputs(920) <= not(inputs(23));
    layer0_outputs(921) <= not(inputs(105)) or (inputs(78));
    layer0_outputs(922) <= not(inputs(203));
    layer0_outputs(923) <= not(inputs(205)) or (inputs(114));
    layer0_outputs(924) <= not((inputs(144)) xor (inputs(168)));
    layer0_outputs(925) <= (inputs(182)) or (inputs(111));
    layer0_outputs(926) <= not((inputs(251)) xor (inputs(5)));
    layer0_outputs(927) <= (inputs(186)) and not (inputs(33));
    layer0_outputs(928) <= not(inputs(137)) or (inputs(31));
    layer0_outputs(929) <= not(inputs(160));
    layer0_outputs(930) <= not(inputs(126));
    layer0_outputs(931) <= (inputs(33)) or (inputs(117));
    layer0_outputs(932) <= not(inputs(47));
    layer0_outputs(933) <= not((inputs(177)) xor (inputs(238)));
    layer0_outputs(934) <= not((inputs(78)) or (inputs(12)));
    layer0_outputs(935) <= inputs(163);
    layer0_outputs(936) <= (inputs(84)) or (inputs(180));
    layer0_outputs(937) <= not(inputs(181)) or (inputs(18));
    layer0_outputs(938) <= (inputs(222)) or (inputs(136));
    layer0_outputs(939) <= not(inputs(68)) or (inputs(154));
    layer0_outputs(940) <= not((inputs(14)) or (inputs(182)));
    layer0_outputs(941) <= (inputs(41)) and (inputs(133));
    layer0_outputs(942) <= not((inputs(123)) xor (inputs(185)));
    layer0_outputs(943) <= not((inputs(29)) or (inputs(101)));
    layer0_outputs(944) <= (inputs(238)) or (inputs(73));
    layer0_outputs(945) <= inputs(21);
    layer0_outputs(946) <= not(inputs(73));
    layer0_outputs(947) <= (inputs(164)) and not (inputs(115));
    layer0_outputs(948) <= (inputs(221)) or (inputs(229));
    layer0_outputs(949) <= not(inputs(53)) or (inputs(127));
    layer0_outputs(950) <= not(inputs(10));
    layer0_outputs(951) <= (inputs(106)) and not (inputs(15));
    layer0_outputs(952) <= not((inputs(228)) or (inputs(217)));
    layer0_outputs(953) <= inputs(136);
    layer0_outputs(954) <= not((inputs(93)) xor (inputs(65)));
    layer0_outputs(955) <= inputs(25);
    layer0_outputs(956) <= inputs(125);
    layer0_outputs(957) <= not(inputs(200)) or (inputs(108));
    layer0_outputs(958) <= inputs(128);
    layer0_outputs(959) <= not(inputs(246));
    layer0_outputs(960) <= (inputs(177)) xor (inputs(118));
    layer0_outputs(961) <= inputs(244);
    layer0_outputs(962) <= not((inputs(200)) and (inputs(254)));
    layer0_outputs(963) <= (inputs(66)) xor (inputs(27));
    layer0_outputs(964) <= (inputs(182)) or (inputs(97));
    layer0_outputs(965) <= not((inputs(28)) and (inputs(233)));
    layer0_outputs(966) <= not((inputs(4)) xor (inputs(90)));
    layer0_outputs(967) <= (inputs(210)) and (inputs(242));
    layer0_outputs(968) <= not((inputs(82)) and (inputs(160)));
    layer0_outputs(969) <= (inputs(204)) or (inputs(113));
    layer0_outputs(970) <= not(inputs(175));
    layer0_outputs(971) <= not(inputs(163));
    layer0_outputs(972) <= (inputs(243)) or (inputs(29));
    layer0_outputs(973) <= (inputs(76)) and not (inputs(97));
    layer0_outputs(974) <= not((inputs(224)) xor (inputs(248)));
    layer0_outputs(975) <= (inputs(62)) or (inputs(105));
    layer0_outputs(976) <= not(inputs(246));
    layer0_outputs(977) <= (inputs(223)) or (inputs(164));
    layer0_outputs(978) <= (inputs(82)) or (inputs(78));
    layer0_outputs(979) <= (inputs(72)) and not (inputs(186));
    layer0_outputs(980) <= not(inputs(108));
    layer0_outputs(981) <= not((inputs(238)) xor (inputs(204)));
    layer0_outputs(982) <= inputs(139);
    layer0_outputs(983) <= (inputs(135)) xor (inputs(216));
    layer0_outputs(984) <= (inputs(135)) or (inputs(104));
    layer0_outputs(985) <= (inputs(110)) xor (inputs(180));
    layer0_outputs(986) <= (inputs(89)) xor (inputs(27));
    layer0_outputs(987) <= inputs(77);
    layer0_outputs(988) <= not(inputs(166)) or (inputs(143));
    layer0_outputs(989) <= (inputs(138)) or (inputs(4));
    layer0_outputs(990) <= (inputs(48)) or (inputs(20));
    layer0_outputs(991) <= not(inputs(67));
    layer0_outputs(992) <= not(inputs(200)) or (inputs(126));
    layer0_outputs(993) <= not(inputs(149)) or (inputs(82));
    layer0_outputs(994) <= not(inputs(102)) or (inputs(185));
    layer0_outputs(995) <= (inputs(52)) and not (inputs(207));
    layer0_outputs(996) <= (inputs(8)) and (inputs(135));
    layer0_outputs(997) <= inputs(217);
    layer0_outputs(998) <= (inputs(10)) or (inputs(5));
    layer0_outputs(999) <= (inputs(83)) or (inputs(146));
    layer0_outputs(1000) <= not(inputs(243));
    layer0_outputs(1001) <= inputs(3);
    layer0_outputs(1002) <= not(inputs(155)) or (inputs(252));
    layer0_outputs(1003) <= not((inputs(93)) or (inputs(135)));
    layer0_outputs(1004) <= not((inputs(153)) or (inputs(130)));
    layer0_outputs(1005) <= not(inputs(133)) or (inputs(223));
    layer0_outputs(1006) <= not(inputs(77));
    layer0_outputs(1007) <= inputs(245);
    layer0_outputs(1008) <= (inputs(19)) or (inputs(32));
    layer0_outputs(1009) <= not(inputs(73));
    layer0_outputs(1010) <= inputs(194);
    layer0_outputs(1011) <= not(inputs(228));
    layer0_outputs(1012) <= not(inputs(100));
    layer0_outputs(1013) <= not(inputs(100));
    layer0_outputs(1014) <= '0';
    layer0_outputs(1015) <= (inputs(69)) and not (inputs(19));
    layer0_outputs(1016) <= (inputs(246)) and not (inputs(109));
    layer0_outputs(1017) <= (inputs(94)) or (inputs(90));
    layer0_outputs(1018) <= (inputs(22)) and not (inputs(147));
    layer0_outputs(1019) <= not(inputs(37)) or (inputs(190));
    layer0_outputs(1020) <= not(inputs(136));
    layer0_outputs(1021) <= not((inputs(190)) xor (inputs(13)));
    layer0_outputs(1022) <= not(inputs(249)) or (inputs(199));
    layer0_outputs(1023) <= not(inputs(25)) or (inputs(30));
    layer0_outputs(1024) <= (inputs(84)) and not (inputs(149));
    layer0_outputs(1025) <= (inputs(255)) or (inputs(207));
    layer0_outputs(1026) <= (inputs(85)) and not (inputs(164));
    layer0_outputs(1027) <= (inputs(247)) and not (inputs(74));
    layer0_outputs(1028) <= not((inputs(150)) or (inputs(6)));
    layer0_outputs(1029) <= (inputs(150)) xor (inputs(197));
    layer0_outputs(1030) <= (inputs(244)) xor (inputs(218));
    layer0_outputs(1031) <= not(inputs(235));
    layer0_outputs(1032) <= not(inputs(217));
    layer0_outputs(1033) <= (inputs(39)) and not (inputs(127));
    layer0_outputs(1034) <= not((inputs(151)) or (inputs(210)));
    layer0_outputs(1035) <= not((inputs(194)) xor (inputs(115)));
    layer0_outputs(1036) <= not(inputs(231)) or (inputs(5));
    layer0_outputs(1037) <= (inputs(95)) or (inputs(215));
    layer0_outputs(1038) <= not(inputs(130)) or (inputs(169));
    layer0_outputs(1039) <= (inputs(14)) and not (inputs(98));
    layer0_outputs(1040) <= (inputs(173)) or (inputs(182));
    layer0_outputs(1041) <= '1';
    layer0_outputs(1042) <= (inputs(171)) or (inputs(138));
    layer0_outputs(1043) <= not(inputs(98)) or (inputs(58));
    layer0_outputs(1044) <= inputs(21);
    layer0_outputs(1045) <= not(inputs(156));
    layer0_outputs(1046) <= not(inputs(224));
    layer0_outputs(1047) <= (inputs(89)) or (inputs(59));
    layer0_outputs(1048) <= (inputs(66)) or (inputs(179));
    layer0_outputs(1049) <= (inputs(217)) xor (inputs(225));
    layer0_outputs(1050) <= inputs(100);
    layer0_outputs(1051) <= not((inputs(176)) or (inputs(194)));
    layer0_outputs(1052) <= (inputs(7)) and not (inputs(98));
    layer0_outputs(1053) <= (inputs(39)) or (inputs(181));
    layer0_outputs(1054) <= (inputs(12)) or (inputs(13));
    layer0_outputs(1055) <= not(inputs(37)) or (inputs(185));
    layer0_outputs(1056) <= not(inputs(133));
    layer0_outputs(1057) <= not((inputs(95)) or (inputs(185)));
    layer0_outputs(1058) <= (inputs(193)) and (inputs(193));
    layer0_outputs(1059) <= not((inputs(29)) xor (inputs(116)));
    layer0_outputs(1060) <= inputs(22);
    layer0_outputs(1061) <= (inputs(36)) and not (inputs(173));
    layer0_outputs(1062) <= (inputs(205)) xor (inputs(207));
    layer0_outputs(1063) <= not(inputs(110));
    layer0_outputs(1064) <= not(inputs(70));
    layer0_outputs(1065) <= not(inputs(116));
    layer0_outputs(1066) <= inputs(193);
    layer0_outputs(1067) <= inputs(58);
    layer0_outputs(1068) <= (inputs(29)) or (inputs(119));
    layer0_outputs(1069) <= not(inputs(165));
    layer0_outputs(1070) <= (inputs(5)) and not (inputs(197));
    layer0_outputs(1071) <= (inputs(208)) and (inputs(109));
    layer0_outputs(1072) <= not((inputs(67)) or (inputs(179)));
    layer0_outputs(1073) <= not((inputs(233)) and (inputs(73)));
    layer0_outputs(1074) <= (inputs(39)) and (inputs(207));
    layer0_outputs(1075) <= not(inputs(8)) or (inputs(80));
    layer0_outputs(1076) <= not(inputs(52)) or (inputs(221));
    layer0_outputs(1077) <= not((inputs(53)) xor (inputs(133)));
    layer0_outputs(1078) <= not(inputs(225));
    layer0_outputs(1079) <= not((inputs(160)) xor (inputs(111)));
    layer0_outputs(1080) <= not(inputs(154));
    layer0_outputs(1081) <= (inputs(65)) or (inputs(103));
    layer0_outputs(1082) <= (inputs(83)) xor (inputs(165));
    layer0_outputs(1083) <= not((inputs(116)) xor (inputs(184)));
    layer0_outputs(1084) <= not(inputs(109));
    layer0_outputs(1085) <= not(inputs(63));
    layer0_outputs(1086) <= not(inputs(142));
    layer0_outputs(1087) <= (inputs(169)) and (inputs(97));
    layer0_outputs(1088) <= (inputs(168)) and not (inputs(136));
    layer0_outputs(1089) <= not(inputs(203));
    layer0_outputs(1090) <= not(inputs(138));
    layer0_outputs(1091) <= not(inputs(74));
    layer0_outputs(1092) <= not((inputs(106)) or (inputs(46)));
    layer0_outputs(1093) <= (inputs(55)) or (inputs(120));
    layer0_outputs(1094) <= (inputs(88)) and not (inputs(192));
    layer0_outputs(1095) <= inputs(219);
    layer0_outputs(1096) <= (inputs(137)) or (inputs(154));
    layer0_outputs(1097) <= (inputs(165)) and not (inputs(151));
    layer0_outputs(1098) <= not(inputs(53)) or (inputs(222));
    layer0_outputs(1099) <= (inputs(175)) or (inputs(89));
    layer0_outputs(1100) <= (inputs(155)) and not (inputs(68));
    layer0_outputs(1101) <= inputs(74);
    layer0_outputs(1102) <= (inputs(186)) or (inputs(32));
    layer0_outputs(1103) <= inputs(58);
    layer0_outputs(1104) <= (inputs(37)) and not (inputs(205));
    layer0_outputs(1105) <= (inputs(238)) or (inputs(93));
    layer0_outputs(1106) <= not((inputs(157)) or (inputs(88)));
    layer0_outputs(1107) <= not(inputs(45));
    layer0_outputs(1108) <= (inputs(211)) and not (inputs(79));
    layer0_outputs(1109) <= not((inputs(253)) or (inputs(101)));
    layer0_outputs(1110) <= not(inputs(227)) or (inputs(253));
    layer0_outputs(1111) <= (inputs(72)) xor (inputs(134));
    layer0_outputs(1112) <= inputs(69);
    layer0_outputs(1113) <= not(inputs(195)) or (inputs(241));
    layer0_outputs(1114) <= not((inputs(150)) xor (inputs(118)));
    layer0_outputs(1115) <= inputs(213);
    layer0_outputs(1116) <= not(inputs(198));
    layer0_outputs(1117) <= (inputs(138)) xor (inputs(233));
    layer0_outputs(1118) <= (inputs(203)) xor (inputs(195));
    layer0_outputs(1119) <= not(inputs(23));
    layer0_outputs(1120) <= not((inputs(120)) or (inputs(123)));
    layer0_outputs(1121) <= not(inputs(120));
    layer0_outputs(1122) <= (inputs(87)) xor (inputs(28));
    layer0_outputs(1123) <= not((inputs(105)) or (inputs(68)));
    layer0_outputs(1124) <= not((inputs(80)) or (inputs(190)));
    layer0_outputs(1125) <= not(inputs(162));
    layer0_outputs(1126) <= (inputs(243)) xor (inputs(177));
    layer0_outputs(1127) <= (inputs(191)) or (inputs(134));
    layer0_outputs(1128) <= (inputs(230)) and not (inputs(112));
    layer0_outputs(1129) <= not(inputs(27));
    layer0_outputs(1130) <= not((inputs(159)) or (inputs(65)));
    layer0_outputs(1131) <= not(inputs(75));
    layer0_outputs(1132) <= inputs(151);
    layer0_outputs(1133) <= (inputs(46)) xor (inputs(73));
    layer0_outputs(1134) <= not(inputs(53)) or (inputs(190));
    layer0_outputs(1135) <= not((inputs(202)) or (inputs(145)));
    layer0_outputs(1136) <= not(inputs(140)) or (inputs(161));
    layer0_outputs(1137) <= not((inputs(185)) or (inputs(21)));
    layer0_outputs(1138) <= (inputs(228)) or (inputs(192));
    layer0_outputs(1139) <= (inputs(222)) or (inputs(81));
    layer0_outputs(1140) <= inputs(138);
    layer0_outputs(1141) <= inputs(248);
    layer0_outputs(1142) <= not(inputs(220));
    layer0_outputs(1143) <= not((inputs(70)) xor (inputs(17)));
    layer0_outputs(1144) <= not(inputs(104));
    layer0_outputs(1145) <= (inputs(205)) and not (inputs(96));
    layer0_outputs(1146) <= (inputs(72)) xor (inputs(2));
    layer0_outputs(1147) <= not(inputs(142));
    layer0_outputs(1148) <= inputs(136);
    layer0_outputs(1149) <= inputs(89);
    layer0_outputs(1150) <= not(inputs(37));
    layer0_outputs(1151) <= not((inputs(53)) xor (inputs(55)));
    layer0_outputs(1152) <= not(inputs(86));
    layer0_outputs(1153) <= not(inputs(21));
    layer0_outputs(1154) <= inputs(125);
    layer0_outputs(1155) <= not(inputs(195)) or (inputs(97));
    layer0_outputs(1156) <= (inputs(35)) and (inputs(0));
    layer0_outputs(1157) <= not(inputs(179));
    layer0_outputs(1158) <= not((inputs(26)) xor (inputs(80)));
    layer0_outputs(1159) <= not(inputs(131));
    layer0_outputs(1160) <= (inputs(40)) and not (inputs(211));
    layer0_outputs(1161) <= (inputs(30)) and not (inputs(33));
    layer0_outputs(1162) <= (inputs(62)) and not (inputs(31));
    layer0_outputs(1163) <= (inputs(237)) xor (inputs(84));
    layer0_outputs(1164) <= not((inputs(78)) or (inputs(54)));
    layer0_outputs(1165) <= (inputs(88)) and (inputs(71));
    layer0_outputs(1166) <= (inputs(235)) or (inputs(97));
    layer0_outputs(1167) <= inputs(57);
    layer0_outputs(1168) <= not((inputs(213)) and (inputs(12)));
    layer0_outputs(1169) <= inputs(99);
    layer0_outputs(1170) <= not((inputs(163)) or (inputs(251)));
    layer0_outputs(1171) <= (inputs(43)) and not (inputs(144));
    layer0_outputs(1172) <= (inputs(192)) and not (inputs(110));
    layer0_outputs(1173) <= (inputs(2)) or (inputs(74));
    layer0_outputs(1174) <= not(inputs(128));
    layer0_outputs(1175) <= not((inputs(112)) xor (inputs(140)));
    layer0_outputs(1176) <= (inputs(128)) or (inputs(86));
    layer0_outputs(1177) <= (inputs(111)) xor (inputs(168));
    layer0_outputs(1178) <= inputs(16);
    layer0_outputs(1179) <= not(inputs(138)) or (inputs(252));
    layer0_outputs(1180) <= (inputs(246)) and not (inputs(199));
    layer0_outputs(1181) <= inputs(177);
    layer0_outputs(1182) <= inputs(226);
    layer0_outputs(1183) <= (inputs(194)) or (inputs(178));
    layer0_outputs(1184) <= (inputs(41)) and not (inputs(226));
    layer0_outputs(1185) <= (inputs(33)) xor (inputs(105));
    layer0_outputs(1186) <= (inputs(42)) and not (inputs(185));
    layer0_outputs(1187) <= not(inputs(117));
    layer0_outputs(1188) <= (inputs(95)) xor (inputs(89));
    layer0_outputs(1189) <= inputs(76);
    layer0_outputs(1190) <= (inputs(139)) or (inputs(245));
    layer0_outputs(1191) <= inputs(249);
    layer0_outputs(1192) <= not(inputs(105));
    layer0_outputs(1193) <= inputs(160);
    layer0_outputs(1194) <= not((inputs(61)) or (inputs(117)));
    layer0_outputs(1195) <= (inputs(69)) and not (inputs(235));
    layer0_outputs(1196) <= not((inputs(247)) or (inputs(62)));
    layer0_outputs(1197) <= not(inputs(215)) or (inputs(34));
    layer0_outputs(1198) <= inputs(184);
    layer0_outputs(1199) <= (inputs(0)) or (inputs(171));
    layer0_outputs(1200) <= inputs(246);
    layer0_outputs(1201) <= inputs(212);
    layer0_outputs(1202) <= not((inputs(153)) and (inputs(157)));
    layer0_outputs(1203) <= not(inputs(166));
    layer0_outputs(1204) <= not(inputs(50)) or (inputs(102));
    layer0_outputs(1205) <= (inputs(35)) and not (inputs(205));
    layer0_outputs(1206) <= not(inputs(254));
    layer0_outputs(1207) <= not(inputs(229)) or (inputs(141));
    layer0_outputs(1208) <= (inputs(119)) and not (inputs(145));
    layer0_outputs(1209) <= not(inputs(57));
    layer0_outputs(1210) <= (inputs(29)) or (inputs(138));
    layer0_outputs(1211) <= not((inputs(130)) or (inputs(129)));
    layer0_outputs(1212) <= not(inputs(84)) or (inputs(225));
    layer0_outputs(1213) <= not(inputs(167));
    layer0_outputs(1214) <= not((inputs(67)) or (inputs(125)));
    layer0_outputs(1215) <= not(inputs(180)) or (inputs(34));
    layer0_outputs(1216) <= not((inputs(124)) xor (inputs(220)));
    layer0_outputs(1217) <= not(inputs(14));
    layer0_outputs(1218) <= not(inputs(131)) or (inputs(181));
    layer0_outputs(1219) <= inputs(90);
    layer0_outputs(1220) <= (inputs(249)) and not (inputs(13));
    layer0_outputs(1221) <= not((inputs(16)) or (inputs(156)));
    layer0_outputs(1222) <= (inputs(25)) or (inputs(140));
    layer0_outputs(1223) <= '0';
    layer0_outputs(1224) <= not((inputs(105)) or (inputs(58)));
    layer0_outputs(1225) <= (inputs(83)) or (inputs(176));
    layer0_outputs(1226) <= inputs(75);
    layer0_outputs(1227) <= (inputs(40)) and not (inputs(171));
    layer0_outputs(1228) <= not((inputs(99)) and (inputs(25)));
    layer0_outputs(1229) <= not(inputs(84)) or (inputs(53));
    layer0_outputs(1230) <= not(inputs(63));
    layer0_outputs(1231) <= not(inputs(197)) or (inputs(94));
    layer0_outputs(1232) <= not(inputs(103));
    layer0_outputs(1233) <= not((inputs(195)) or (inputs(198)));
    layer0_outputs(1234) <= not(inputs(120));
    layer0_outputs(1235) <= (inputs(181)) or (inputs(83));
    layer0_outputs(1236) <= inputs(215);
    layer0_outputs(1237) <= not(inputs(247)) or (inputs(14));
    layer0_outputs(1238) <= (inputs(86)) xor (inputs(115));
    layer0_outputs(1239) <= not((inputs(3)) xor (inputs(32)));
    layer0_outputs(1240) <= inputs(122);
    layer0_outputs(1241) <= (inputs(150)) or (inputs(151));
    layer0_outputs(1242) <= not(inputs(57)) or (inputs(147));
    layer0_outputs(1243) <= '0';
    layer0_outputs(1244) <= (inputs(107)) and not (inputs(132));
    layer0_outputs(1245) <= not(inputs(191)) or (inputs(239));
    layer0_outputs(1246) <= (inputs(109)) and not (inputs(62));
    layer0_outputs(1247) <= (inputs(64)) and (inputs(87));
    layer0_outputs(1248) <= not(inputs(218));
    layer0_outputs(1249) <= not(inputs(148));
    layer0_outputs(1250) <= (inputs(56)) or (inputs(58));
    layer0_outputs(1251) <= (inputs(231)) and not (inputs(78));
    layer0_outputs(1252) <= (inputs(110)) or (inputs(228));
    layer0_outputs(1253) <= not((inputs(130)) or (inputs(160)));
    layer0_outputs(1254) <= not(inputs(83));
    layer0_outputs(1255) <= not((inputs(42)) and (inputs(23)));
    layer0_outputs(1256) <= not((inputs(140)) xor (inputs(234)));
    layer0_outputs(1257) <= inputs(91);
    layer0_outputs(1258) <= (inputs(195)) xor (inputs(47));
    layer0_outputs(1259) <= not(inputs(246)) or (inputs(18));
    layer0_outputs(1260) <= not(inputs(76));
    layer0_outputs(1261) <= not(inputs(225)) or (inputs(56));
    layer0_outputs(1262) <= (inputs(107)) and not (inputs(150));
    layer0_outputs(1263) <= inputs(35);
    layer0_outputs(1264) <= inputs(129);
    layer0_outputs(1265) <= (inputs(18)) xor (inputs(180));
    layer0_outputs(1266) <= inputs(103);
    layer0_outputs(1267) <= not((inputs(101)) or (inputs(66)));
    layer0_outputs(1268) <= not((inputs(221)) and (inputs(249)));
    layer0_outputs(1269) <= (inputs(61)) xor (inputs(92));
    layer0_outputs(1270) <= '1';
    layer0_outputs(1271) <= not(inputs(82));
    layer0_outputs(1272) <= not((inputs(68)) or (inputs(111)));
    layer0_outputs(1273) <= (inputs(125)) xor (inputs(73));
    layer0_outputs(1274) <= not(inputs(246)) or (inputs(96));
    layer0_outputs(1275) <= (inputs(113)) xor (inputs(218));
    layer0_outputs(1276) <= (inputs(27)) and not (inputs(125));
    layer0_outputs(1277) <= (inputs(8)) and (inputs(83));
    layer0_outputs(1278) <= not((inputs(83)) and (inputs(4)));
    layer0_outputs(1279) <= (inputs(49)) or (inputs(80));
    layer0_outputs(1280) <= (inputs(118)) and not (inputs(188));
    layer0_outputs(1281) <= (inputs(37)) and not (inputs(37));
    layer0_outputs(1282) <= not(inputs(228));
    layer0_outputs(1283) <= inputs(179);
    layer0_outputs(1284) <= (inputs(57)) xor (inputs(123));
    layer0_outputs(1285) <= (inputs(127)) or (inputs(196));
    layer0_outputs(1286) <= (inputs(176)) and not (inputs(39));
    layer0_outputs(1287) <= not((inputs(180)) or (inputs(107)));
    layer0_outputs(1288) <= (inputs(116)) or (inputs(62));
    layer0_outputs(1289) <= (inputs(194)) and not (inputs(113));
    layer0_outputs(1290) <= not((inputs(248)) or (inputs(113)));
    layer0_outputs(1291) <= (inputs(10)) and (inputs(82));
    layer0_outputs(1292) <= not(inputs(96)) or (inputs(181));
    layer0_outputs(1293) <= (inputs(29)) xor (inputs(111));
    layer0_outputs(1294) <= not((inputs(236)) or (inputs(149)));
    layer0_outputs(1295) <= inputs(162);
    layer0_outputs(1296) <= not((inputs(112)) or (inputs(231)));
    layer0_outputs(1297) <= (inputs(11)) xor (inputs(128));
    layer0_outputs(1298) <= not((inputs(56)) xor (inputs(5)));
    layer0_outputs(1299) <= inputs(241);
    layer0_outputs(1300) <= not(inputs(105));
    layer0_outputs(1301) <= not(inputs(76)) or (inputs(239));
    layer0_outputs(1302) <= not((inputs(59)) or (inputs(5)));
    layer0_outputs(1303) <= (inputs(221)) and not (inputs(93));
    layer0_outputs(1304) <= not((inputs(7)) or (inputs(85)));
    layer0_outputs(1305) <= not(inputs(18));
    layer0_outputs(1306) <= not((inputs(153)) xor (inputs(243)));
    layer0_outputs(1307) <= not(inputs(11));
    layer0_outputs(1308) <= (inputs(129)) or (inputs(147));
    layer0_outputs(1309) <= (inputs(153)) and (inputs(56));
    layer0_outputs(1310) <= not((inputs(10)) xor (inputs(243)));
    layer0_outputs(1311) <= not((inputs(149)) xor (inputs(56)));
    layer0_outputs(1312) <= not((inputs(236)) xor (inputs(61)));
    layer0_outputs(1313) <= (inputs(65)) and not (inputs(143));
    layer0_outputs(1314) <= (inputs(220)) and not (inputs(0));
    layer0_outputs(1315) <= (inputs(182)) xor (inputs(17));
    layer0_outputs(1316) <= not(inputs(6)) or (inputs(15));
    layer0_outputs(1317) <= (inputs(84)) and not (inputs(210));
    layer0_outputs(1318) <= (inputs(123)) and (inputs(48));
    layer0_outputs(1319) <= (inputs(96)) or (inputs(212));
    layer0_outputs(1320) <= not((inputs(206)) and (inputs(244)));
    layer0_outputs(1321) <= (inputs(55)) xor (inputs(138));
    layer0_outputs(1322) <= not(inputs(84));
    layer0_outputs(1323) <= (inputs(5)) or (inputs(214));
    layer0_outputs(1324) <= (inputs(190)) and not (inputs(47));
    layer0_outputs(1325) <= not((inputs(24)) xor (inputs(56)));
    layer0_outputs(1326) <= (inputs(43)) or (inputs(158));
    layer0_outputs(1327) <= not((inputs(137)) xor (inputs(58)));
    layer0_outputs(1328) <= (inputs(133)) and not (inputs(32));
    layer0_outputs(1329) <= not((inputs(100)) xor (inputs(188)));
    layer0_outputs(1330) <= not(inputs(47));
    layer0_outputs(1331) <= not((inputs(154)) xor (inputs(90)));
    layer0_outputs(1332) <= not((inputs(7)) or (inputs(164)));
    layer0_outputs(1333) <= (inputs(42)) and not (inputs(247));
    layer0_outputs(1334) <= '1';
    layer0_outputs(1335) <= (inputs(171)) xor (inputs(30));
    layer0_outputs(1336) <= (inputs(37)) xor (inputs(5));
    layer0_outputs(1337) <= not(inputs(131)) or (inputs(248));
    layer0_outputs(1338) <= not(inputs(90)) or (inputs(161));
    layer0_outputs(1339) <= not(inputs(204));
    layer0_outputs(1340) <= (inputs(83)) and not (inputs(160));
    layer0_outputs(1341) <= (inputs(113)) or (inputs(195));
    layer0_outputs(1342) <= inputs(246);
    layer0_outputs(1343) <= not(inputs(221));
    layer0_outputs(1344) <= not((inputs(30)) or (inputs(169)));
    layer0_outputs(1345) <= (inputs(121)) and not (inputs(50));
    layer0_outputs(1346) <= not(inputs(86));
    layer0_outputs(1347) <= (inputs(88)) and not (inputs(244));
    layer0_outputs(1348) <= (inputs(117)) and not (inputs(53));
    layer0_outputs(1349) <= (inputs(161)) or (inputs(226));
    layer0_outputs(1350) <= not((inputs(199)) xor (inputs(202)));
    layer0_outputs(1351) <= not((inputs(138)) or (inputs(101)));
    layer0_outputs(1352) <= not((inputs(98)) or (inputs(115)));
    layer0_outputs(1353) <= not((inputs(99)) or (inputs(84)));
    layer0_outputs(1354) <= not(inputs(146));
    layer0_outputs(1355) <= inputs(27);
    layer0_outputs(1356) <= not(inputs(134));
    layer0_outputs(1357) <= not(inputs(246));
    layer0_outputs(1358) <= not(inputs(228)) or (inputs(77));
    layer0_outputs(1359) <= (inputs(104)) and not (inputs(100));
    layer0_outputs(1360) <= (inputs(251)) xor (inputs(240));
    layer0_outputs(1361) <= (inputs(0)) or (inputs(145));
    layer0_outputs(1362) <= (inputs(20)) or (inputs(79));
    layer0_outputs(1363) <= inputs(93);
    layer0_outputs(1364) <= not((inputs(197)) xor (inputs(77)));
    layer0_outputs(1365) <= inputs(9);
    layer0_outputs(1366) <= not((inputs(166)) xor (inputs(246)));
    layer0_outputs(1367) <= (inputs(106)) and not (inputs(53));
    layer0_outputs(1368) <= not(inputs(115));
    layer0_outputs(1369) <= inputs(8);
    layer0_outputs(1370) <= not((inputs(217)) xor (inputs(186)));
    layer0_outputs(1371) <= not(inputs(24));
    layer0_outputs(1372) <= (inputs(158)) xor (inputs(223));
    layer0_outputs(1373) <= not(inputs(243)) or (inputs(217));
    layer0_outputs(1374) <= not(inputs(171)) or (inputs(167));
    layer0_outputs(1375) <= not((inputs(125)) xor (inputs(159)));
    layer0_outputs(1376) <= not((inputs(49)) xor (inputs(177)));
    layer0_outputs(1377) <= not(inputs(152)) or (inputs(0));
    layer0_outputs(1378) <= (inputs(172)) and not (inputs(133));
    layer0_outputs(1379) <= not((inputs(57)) or (inputs(32)));
    layer0_outputs(1380) <= (inputs(170)) and not (inputs(72));
    layer0_outputs(1381) <= (inputs(77)) or (inputs(32));
    layer0_outputs(1382) <= (inputs(224)) xor (inputs(8));
    layer0_outputs(1383) <= (inputs(148)) or (inputs(126));
    layer0_outputs(1384) <= not((inputs(41)) or (inputs(49)));
    layer0_outputs(1385) <= inputs(210);
    layer0_outputs(1386) <= inputs(79);
    layer0_outputs(1387) <= not((inputs(200)) xor (inputs(124)));
    layer0_outputs(1388) <= not((inputs(150)) or (inputs(50)));
    layer0_outputs(1389) <= not(inputs(251));
    layer0_outputs(1390) <= not(inputs(100));
    layer0_outputs(1391) <= not((inputs(243)) xor (inputs(236)));
    layer0_outputs(1392) <= (inputs(110)) or (inputs(152));
    layer0_outputs(1393) <= inputs(152);
    layer0_outputs(1394) <= inputs(63);
    layer0_outputs(1395) <= (inputs(51)) and not (inputs(249));
    layer0_outputs(1396) <= not(inputs(91));
    layer0_outputs(1397) <= inputs(187);
    layer0_outputs(1398) <= (inputs(120)) and not (inputs(177));
    layer0_outputs(1399) <= (inputs(47)) xor (inputs(129));
    layer0_outputs(1400) <= not(inputs(225));
    layer0_outputs(1401) <= not(inputs(247));
    layer0_outputs(1402) <= (inputs(92)) or (inputs(94));
    layer0_outputs(1403) <= not(inputs(39));
    layer0_outputs(1404) <= (inputs(220)) and (inputs(199));
    layer0_outputs(1405) <= inputs(233);
    layer0_outputs(1406) <= (inputs(111)) or (inputs(132));
    layer0_outputs(1407) <= not((inputs(117)) or (inputs(249)));
    layer0_outputs(1408) <= not((inputs(22)) and (inputs(229)));
    layer0_outputs(1409) <= (inputs(103)) xor (inputs(205));
    layer0_outputs(1410) <= not((inputs(149)) xor (inputs(35)));
    layer0_outputs(1411) <= inputs(249);
    layer0_outputs(1412) <= not((inputs(3)) xor (inputs(60)));
    layer0_outputs(1413) <= (inputs(180)) or (inputs(163));
    layer0_outputs(1414) <= not((inputs(218)) xor (inputs(139)));
    layer0_outputs(1415) <= (inputs(209)) xor (inputs(246));
    layer0_outputs(1416) <= (inputs(40)) and (inputs(140));
    layer0_outputs(1417) <= inputs(232);
    layer0_outputs(1418) <= not((inputs(210)) or (inputs(55)));
    layer0_outputs(1419) <= not((inputs(6)) or (inputs(20)));
    layer0_outputs(1420) <= not((inputs(207)) xor (inputs(131)));
    layer0_outputs(1421) <= inputs(210);
    layer0_outputs(1422) <= not(inputs(186)) or (inputs(52));
    layer0_outputs(1423) <= not(inputs(70));
    layer0_outputs(1424) <= inputs(107);
    layer0_outputs(1425) <= not(inputs(125));
    layer0_outputs(1426) <= not(inputs(247)) or (inputs(95));
    layer0_outputs(1427) <= (inputs(45)) xor (inputs(165));
    layer0_outputs(1428) <= not(inputs(12));
    layer0_outputs(1429) <= not((inputs(116)) xor (inputs(169)));
    layer0_outputs(1430) <= not((inputs(41)) xor (inputs(88)));
    layer0_outputs(1431) <= (inputs(227)) or (inputs(239));
    layer0_outputs(1432) <= '0';
    layer0_outputs(1433) <= (inputs(14)) or (inputs(150));
    layer0_outputs(1434) <= not((inputs(232)) xor (inputs(139)));
    layer0_outputs(1435) <= not(inputs(61));
    layer0_outputs(1436) <= not(inputs(83));
    layer0_outputs(1437) <= not(inputs(217));
    layer0_outputs(1438) <= (inputs(230)) and not (inputs(81));
    layer0_outputs(1439) <= (inputs(118)) or (inputs(155));
    layer0_outputs(1440) <= not(inputs(194)) or (inputs(223));
    layer0_outputs(1441) <= (inputs(225)) xor (inputs(186));
    layer0_outputs(1442) <= (inputs(77)) xor (inputs(186));
    layer0_outputs(1443) <= not((inputs(158)) xor (inputs(137)));
    layer0_outputs(1444) <= (inputs(88)) xor (inputs(128));
    layer0_outputs(1445) <= (inputs(173)) xor (inputs(99));
    layer0_outputs(1446) <= (inputs(177)) and not (inputs(244));
    layer0_outputs(1447) <= not(inputs(72));
    layer0_outputs(1448) <= not(inputs(28));
    layer0_outputs(1449) <= not((inputs(249)) or (inputs(146)));
    layer0_outputs(1450) <= (inputs(221)) or (inputs(177));
    layer0_outputs(1451) <= (inputs(247)) or (inputs(195));
    layer0_outputs(1452) <= (inputs(129)) xor (inputs(170));
    layer0_outputs(1453) <= not(inputs(115));
    layer0_outputs(1454) <= not((inputs(180)) or (inputs(221)));
    layer0_outputs(1455) <= '0';
    layer0_outputs(1456) <= not(inputs(33));
    layer0_outputs(1457) <= not(inputs(232));
    layer0_outputs(1458) <= not(inputs(69)) or (inputs(221));
    layer0_outputs(1459) <= inputs(128);
    layer0_outputs(1460) <= (inputs(238)) and not (inputs(93));
    layer0_outputs(1461) <= not(inputs(80));
    layer0_outputs(1462) <= (inputs(5)) or (inputs(135));
    layer0_outputs(1463) <= not(inputs(137));
    layer0_outputs(1464) <= (inputs(93)) and not (inputs(2));
    layer0_outputs(1465) <= not(inputs(85)) or (inputs(62));
    layer0_outputs(1466) <= (inputs(179)) xor (inputs(147));
    layer0_outputs(1467) <= (inputs(81)) or (inputs(10));
    layer0_outputs(1468) <= (inputs(171)) xor (inputs(151));
    layer0_outputs(1469) <= not(inputs(50));
    layer0_outputs(1470) <= not(inputs(151)) or (inputs(206));
    layer0_outputs(1471) <= not((inputs(10)) or (inputs(229)));
    layer0_outputs(1472) <= not((inputs(152)) xor (inputs(217)));
    layer0_outputs(1473) <= not((inputs(55)) or (inputs(46)));
    layer0_outputs(1474) <= '0';
    layer0_outputs(1475) <= not(inputs(32));
    layer0_outputs(1476) <= (inputs(33)) xor (inputs(122));
    layer0_outputs(1477) <= not(inputs(130));
    layer0_outputs(1478) <= inputs(161);
    layer0_outputs(1479) <= inputs(44);
    layer0_outputs(1480) <= not(inputs(117));
    layer0_outputs(1481) <= not((inputs(130)) or (inputs(176)));
    layer0_outputs(1482) <= (inputs(163)) or (inputs(205));
    layer0_outputs(1483) <= not(inputs(182));
    layer0_outputs(1484) <= inputs(129);
    layer0_outputs(1485) <= not((inputs(157)) or (inputs(231)));
    layer0_outputs(1486) <= not(inputs(24)) or (inputs(29));
    layer0_outputs(1487) <= not(inputs(245));
    layer0_outputs(1488) <= inputs(169);
    layer0_outputs(1489) <= not((inputs(226)) or (inputs(224)));
    layer0_outputs(1490) <= inputs(90);
    layer0_outputs(1491) <= not((inputs(55)) xor (inputs(90)));
    layer0_outputs(1492) <= not((inputs(148)) xor (inputs(36)));
    layer0_outputs(1493) <= inputs(117);
    layer0_outputs(1494) <= (inputs(4)) xor (inputs(188));
    layer0_outputs(1495) <= (inputs(120)) and not (inputs(186));
    layer0_outputs(1496) <= not(inputs(117)) or (inputs(244));
    layer0_outputs(1497) <= (inputs(30)) or (inputs(98));
    layer0_outputs(1498) <= (inputs(111)) or (inputs(165));
    layer0_outputs(1499) <= (inputs(237)) and not (inputs(17));
    layer0_outputs(1500) <= not(inputs(213));
    layer0_outputs(1501) <= (inputs(101)) or (inputs(32));
    layer0_outputs(1502) <= inputs(130);
    layer0_outputs(1503) <= (inputs(246)) or (inputs(227));
    layer0_outputs(1504) <= inputs(170);
    layer0_outputs(1505) <= not(inputs(74));
    layer0_outputs(1506) <= not(inputs(12));
    layer0_outputs(1507) <= not((inputs(86)) xor (inputs(60)));
    layer0_outputs(1508) <= not(inputs(100));
    layer0_outputs(1509) <= inputs(207);
    layer0_outputs(1510) <= not(inputs(63));
    layer0_outputs(1511) <= not((inputs(200)) or (inputs(230)));
    layer0_outputs(1512) <= inputs(120);
    layer0_outputs(1513) <= not((inputs(124)) xor (inputs(2)));
    layer0_outputs(1514) <= (inputs(207)) or (inputs(78));
    layer0_outputs(1515) <= not(inputs(203));
    layer0_outputs(1516) <= not(inputs(12));
    layer0_outputs(1517) <= not((inputs(43)) xor (inputs(45)));
    layer0_outputs(1518) <= (inputs(233)) and not (inputs(182));
    layer0_outputs(1519) <= not((inputs(117)) or (inputs(45)));
    layer0_outputs(1520) <= (inputs(69)) xor (inputs(39));
    layer0_outputs(1521) <= not((inputs(174)) or (inputs(250)));
    layer0_outputs(1522) <= (inputs(150)) and not (inputs(238));
    layer0_outputs(1523) <= (inputs(184)) xor (inputs(203));
    layer0_outputs(1524) <= (inputs(4)) xor (inputs(48));
    layer0_outputs(1525) <= (inputs(171)) and not (inputs(191));
    layer0_outputs(1526) <= (inputs(201)) or (inputs(180));
    layer0_outputs(1527) <= (inputs(138)) or (inputs(66));
    layer0_outputs(1528) <= not(inputs(25)) or (inputs(146));
    layer0_outputs(1529) <= not(inputs(177)) or (inputs(185));
    layer0_outputs(1530) <= (inputs(182)) xor (inputs(200));
    layer0_outputs(1531) <= (inputs(94)) or (inputs(120));
    layer0_outputs(1532) <= inputs(106);
    layer0_outputs(1533) <= (inputs(3)) and not (inputs(220));
    layer0_outputs(1534) <= not((inputs(69)) xor (inputs(73)));
    layer0_outputs(1535) <= (inputs(66)) xor (inputs(148));
    layer0_outputs(1536) <= not((inputs(23)) xor (inputs(28)));
    layer0_outputs(1537) <= not(inputs(25)) or (inputs(174));
    layer0_outputs(1538) <= (inputs(109)) and (inputs(175));
    layer0_outputs(1539) <= not((inputs(48)) xor (inputs(12)));
    layer0_outputs(1540) <= not(inputs(51)) or (inputs(217));
    layer0_outputs(1541) <= not(inputs(175)) or (inputs(229));
    layer0_outputs(1542) <= not(inputs(163));
    layer0_outputs(1543) <= not((inputs(49)) xor (inputs(152)));
    layer0_outputs(1544) <= (inputs(167)) and not (inputs(190));
    layer0_outputs(1545) <= not(inputs(176));
    layer0_outputs(1546) <= not((inputs(169)) and (inputs(181)));
    layer0_outputs(1547) <= inputs(205);
    layer0_outputs(1548) <= inputs(198);
    layer0_outputs(1549) <= not(inputs(250)) or (inputs(93));
    layer0_outputs(1550) <= not((inputs(180)) xor (inputs(118)));
    layer0_outputs(1551) <= not(inputs(93)) or (inputs(207));
    layer0_outputs(1552) <= (inputs(19)) or (inputs(39));
    layer0_outputs(1553) <= inputs(103);
    layer0_outputs(1554) <= (inputs(204)) and not (inputs(112));
    layer0_outputs(1555) <= not(inputs(167)) or (inputs(69));
    layer0_outputs(1556) <= inputs(51);
    layer0_outputs(1557) <= (inputs(102)) xor (inputs(6));
    layer0_outputs(1558) <= not(inputs(75));
    layer0_outputs(1559) <= not(inputs(85)) or (inputs(175));
    layer0_outputs(1560) <= inputs(68);
    layer0_outputs(1561) <= (inputs(150)) and not (inputs(236));
    layer0_outputs(1562) <= (inputs(80)) xor (inputs(225));
    layer0_outputs(1563) <= inputs(233);
    layer0_outputs(1564) <= not((inputs(22)) xor (inputs(249)));
    layer0_outputs(1565) <= not(inputs(8));
    layer0_outputs(1566) <= not(inputs(24)) or (inputs(156));
    layer0_outputs(1567) <= not(inputs(207));
    layer0_outputs(1568) <= not((inputs(185)) or (inputs(9)));
    layer0_outputs(1569) <= not((inputs(172)) or (inputs(115)));
    layer0_outputs(1570) <= not(inputs(69)) or (inputs(209));
    layer0_outputs(1571) <= (inputs(238)) xor (inputs(26));
    layer0_outputs(1572) <= inputs(253);
    layer0_outputs(1573) <= inputs(57);
    layer0_outputs(1574) <= not((inputs(142)) or (inputs(141)));
    layer0_outputs(1575) <= not(inputs(211));
    layer0_outputs(1576) <= not(inputs(241));
    layer0_outputs(1577) <= (inputs(156)) xor (inputs(236));
    layer0_outputs(1578) <= not(inputs(132)) or (inputs(50));
    layer0_outputs(1579) <= (inputs(51)) or (inputs(18));
    layer0_outputs(1580) <= not((inputs(183)) xor (inputs(27)));
    layer0_outputs(1581) <= inputs(9);
    layer0_outputs(1582) <= not((inputs(37)) xor (inputs(4)));
    layer0_outputs(1583) <= not(inputs(124));
    layer0_outputs(1584) <= (inputs(200)) xor (inputs(153));
    layer0_outputs(1585) <= (inputs(186)) and not (inputs(5));
    layer0_outputs(1586) <= not(inputs(173));
    layer0_outputs(1587) <= not(inputs(16));
    layer0_outputs(1588) <= not(inputs(90));
    layer0_outputs(1589) <= (inputs(182)) and not (inputs(139));
    layer0_outputs(1590) <= not(inputs(12));
    layer0_outputs(1591) <= not(inputs(92)) or (inputs(157));
    layer0_outputs(1592) <= not(inputs(128)) or (inputs(253));
    layer0_outputs(1593) <= not((inputs(9)) xor (inputs(34)));
    layer0_outputs(1594) <= (inputs(183)) and not (inputs(94));
    layer0_outputs(1595) <= not(inputs(104));
    layer0_outputs(1596) <= not((inputs(91)) and (inputs(119)));
    layer0_outputs(1597) <= not((inputs(31)) xor (inputs(196)));
    layer0_outputs(1598) <= not(inputs(209));
    layer0_outputs(1599) <= not(inputs(65));
    layer0_outputs(1600) <= (inputs(94)) xor (inputs(187));
    layer0_outputs(1601) <= not(inputs(166));
    layer0_outputs(1602) <= inputs(252);
    layer0_outputs(1603) <= (inputs(216)) and not (inputs(2));
    layer0_outputs(1604) <= inputs(172);
    layer0_outputs(1605) <= inputs(252);
    layer0_outputs(1606) <= not(inputs(39)) or (inputs(144));
    layer0_outputs(1607) <= (inputs(197)) xor (inputs(230));
    layer0_outputs(1608) <= not((inputs(130)) xor (inputs(80)));
    layer0_outputs(1609) <= (inputs(4)) and not (inputs(160));
    layer0_outputs(1610) <= inputs(146);
    layer0_outputs(1611) <= not((inputs(109)) xor (inputs(34)));
    layer0_outputs(1612) <= inputs(83);
    layer0_outputs(1613) <= inputs(130);
    layer0_outputs(1614) <= inputs(227);
    layer0_outputs(1615) <= not(inputs(73));
    layer0_outputs(1616) <= not(inputs(107)) or (inputs(14));
    layer0_outputs(1617) <= (inputs(90)) and not (inputs(209));
    layer0_outputs(1618) <= (inputs(140)) and not (inputs(198));
    layer0_outputs(1619) <= (inputs(255)) xor (inputs(249));
    layer0_outputs(1620) <= not((inputs(103)) xor (inputs(134)));
    layer0_outputs(1621) <= not((inputs(17)) or (inputs(129)));
    layer0_outputs(1622) <= not((inputs(67)) xor (inputs(114)));
    layer0_outputs(1623) <= not((inputs(193)) xor (inputs(240)));
    layer0_outputs(1624) <= (inputs(226)) or (inputs(60));
    layer0_outputs(1625) <= (inputs(253)) xor (inputs(130));
    layer0_outputs(1626) <= not((inputs(17)) xor (inputs(46)));
    layer0_outputs(1627) <= (inputs(25)) xor (inputs(75));
    layer0_outputs(1628) <= inputs(78);
    layer0_outputs(1629) <= inputs(226);
    layer0_outputs(1630) <= inputs(90);
    layer0_outputs(1631) <= inputs(155);
    layer0_outputs(1632) <= not((inputs(138)) or (inputs(21)));
    layer0_outputs(1633) <= (inputs(58)) and not (inputs(238));
    layer0_outputs(1634) <= not(inputs(160));
    layer0_outputs(1635) <= not(inputs(70)) or (inputs(242));
    layer0_outputs(1636) <= not((inputs(28)) and (inputs(56)));
    layer0_outputs(1637) <= not((inputs(15)) or (inputs(104)));
    layer0_outputs(1638) <= (inputs(74)) or (inputs(95));
    layer0_outputs(1639) <= not(inputs(240));
    layer0_outputs(1640) <= inputs(91);
    layer0_outputs(1641) <= (inputs(163)) xor (inputs(151));
    layer0_outputs(1642) <= not(inputs(123));
    layer0_outputs(1643) <= not(inputs(117));
    layer0_outputs(1644) <= inputs(118);
    layer0_outputs(1645) <= inputs(220);
    layer0_outputs(1646) <= (inputs(79)) or (inputs(190));
    layer0_outputs(1647) <= (inputs(43)) and not (inputs(32));
    layer0_outputs(1648) <= inputs(148);
    layer0_outputs(1649) <= not(inputs(20)) or (inputs(190));
    layer0_outputs(1650) <= not(inputs(11)) or (inputs(111));
    layer0_outputs(1651) <= (inputs(89)) and not (inputs(252));
    layer0_outputs(1652) <= inputs(57);
    layer0_outputs(1653) <= (inputs(150)) or (inputs(48));
    layer0_outputs(1654) <= inputs(56);
    layer0_outputs(1655) <= not((inputs(188)) or (inputs(10)));
    layer0_outputs(1656) <= (inputs(199)) xor (inputs(123));
    layer0_outputs(1657) <= not(inputs(221)) or (inputs(2));
    layer0_outputs(1658) <= (inputs(74)) and (inputs(57));
    layer0_outputs(1659) <= (inputs(155)) xor (inputs(112));
    layer0_outputs(1660) <= not((inputs(206)) or (inputs(77)));
    layer0_outputs(1661) <= (inputs(106)) xor (inputs(156));
    layer0_outputs(1662) <= not(inputs(136));
    layer0_outputs(1663) <= not((inputs(130)) xor (inputs(65)));
    layer0_outputs(1664) <= not(inputs(248));
    layer0_outputs(1665) <= (inputs(54)) or (inputs(26));
    layer0_outputs(1666) <= not((inputs(214)) or (inputs(237)));
    layer0_outputs(1667) <= (inputs(156)) or (inputs(65));
    layer0_outputs(1668) <= (inputs(231)) xor (inputs(232));
    layer0_outputs(1669) <= (inputs(31)) or (inputs(69));
    layer0_outputs(1670) <= not(inputs(40));
    layer0_outputs(1671) <= not(inputs(151)) or (inputs(113));
    layer0_outputs(1672) <= (inputs(116)) xor (inputs(69));
    layer0_outputs(1673) <= (inputs(83)) or (inputs(203));
    layer0_outputs(1674) <= not((inputs(174)) and (inputs(142)));
    layer0_outputs(1675) <= (inputs(242)) xor (inputs(191));
    layer0_outputs(1676) <= not(inputs(12));
    layer0_outputs(1677) <= not(inputs(66));
    layer0_outputs(1678) <= (inputs(244)) or (inputs(177));
    layer0_outputs(1679) <= not((inputs(151)) or (inputs(70)));
    layer0_outputs(1680) <= inputs(217);
    layer0_outputs(1681) <= inputs(104);
    layer0_outputs(1682) <= (inputs(111)) or (inputs(132));
    layer0_outputs(1683) <= (inputs(179)) and not (inputs(47));
    layer0_outputs(1684) <= not(inputs(74)) or (inputs(127));
    layer0_outputs(1685) <= not((inputs(78)) and (inputs(243)));
    layer0_outputs(1686) <= (inputs(157)) or (inputs(32));
    layer0_outputs(1687) <= (inputs(168)) and not (inputs(251));
    layer0_outputs(1688) <= not((inputs(99)) or (inputs(63)));
    layer0_outputs(1689) <= (inputs(103)) or (inputs(119));
    layer0_outputs(1690) <= not((inputs(73)) xor (inputs(118)));
    layer0_outputs(1691) <= not((inputs(36)) xor (inputs(109)));
    layer0_outputs(1692) <= inputs(142);
    layer0_outputs(1693) <= inputs(128);
    layer0_outputs(1694) <= not((inputs(174)) xor (inputs(6)));
    layer0_outputs(1695) <= (inputs(83)) or (inputs(98));
    layer0_outputs(1696) <= (inputs(227)) and (inputs(23));
    layer0_outputs(1697) <= inputs(106);
    layer0_outputs(1698) <= (inputs(246)) and not (inputs(250));
    layer0_outputs(1699) <= not((inputs(114)) and (inputs(114)));
    layer0_outputs(1700) <= not(inputs(66));
    layer0_outputs(1701) <= not((inputs(114)) or (inputs(192)));
    layer0_outputs(1702) <= (inputs(41)) and not (inputs(142));
    layer0_outputs(1703) <= '1';
    layer0_outputs(1704) <= '0';
    layer0_outputs(1705) <= not((inputs(163)) or (inputs(7)));
    layer0_outputs(1706) <= not(inputs(155)) or (inputs(126));
    layer0_outputs(1707) <= inputs(250);
    layer0_outputs(1708) <= (inputs(82)) and (inputs(162));
    layer0_outputs(1709) <= not(inputs(254)) or (inputs(28));
    layer0_outputs(1710) <= (inputs(91)) and not (inputs(73));
    layer0_outputs(1711) <= inputs(247);
    layer0_outputs(1712) <= not(inputs(139));
    layer0_outputs(1713) <= (inputs(137)) or (inputs(34));
    layer0_outputs(1714) <= inputs(129);
    layer0_outputs(1715) <= (inputs(111)) or (inputs(157));
    layer0_outputs(1716) <= (inputs(52)) or (inputs(120));
    layer0_outputs(1717) <= (inputs(197)) and not (inputs(13));
    layer0_outputs(1718) <= '1';
    layer0_outputs(1719) <= (inputs(175)) and (inputs(19));
    layer0_outputs(1720) <= (inputs(226)) xor (inputs(32));
    layer0_outputs(1721) <= inputs(183);
    layer0_outputs(1722) <= (inputs(146)) and not (inputs(135));
    layer0_outputs(1723) <= (inputs(33)) xor (inputs(67));
    layer0_outputs(1724) <= inputs(168);
    layer0_outputs(1725) <= not(inputs(204));
    layer0_outputs(1726) <= not(inputs(88)) or (inputs(32));
    layer0_outputs(1727) <= not(inputs(24));
    layer0_outputs(1728) <= not(inputs(85)) or (inputs(191));
    layer0_outputs(1729) <= not((inputs(141)) xor (inputs(91)));
    layer0_outputs(1730) <= inputs(102);
    layer0_outputs(1731) <= not(inputs(29));
    layer0_outputs(1732) <= not((inputs(69)) or (inputs(170)));
    layer0_outputs(1733) <= (inputs(111)) and not (inputs(255));
    layer0_outputs(1734) <= (inputs(199)) or (inputs(131));
    layer0_outputs(1735) <= inputs(130);
    layer0_outputs(1736) <= (inputs(116)) and not (inputs(19));
    layer0_outputs(1737) <= not(inputs(15));
    layer0_outputs(1738) <= inputs(239);
    layer0_outputs(1739) <= not((inputs(207)) xor (inputs(22)));
    layer0_outputs(1740) <= not((inputs(246)) xor (inputs(222)));
    layer0_outputs(1741) <= (inputs(112)) xor (inputs(196));
    layer0_outputs(1742) <= not((inputs(106)) xor (inputs(168)));
    layer0_outputs(1743) <= not((inputs(115)) xor (inputs(202)));
    layer0_outputs(1744) <= not((inputs(217)) xor (inputs(32)));
    layer0_outputs(1745) <= (inputs(57)) xor (inputs(7));
    layer0_outputs(1746) <= inputs(47);
    layer0_outputs(1747) <= not((inputs(172)) and (inputs(159)));
    layer0_outputs(1748) <= (inputs(10)) xor (inputs(158));
    layer0_outputs(1749) <= not((inputs(117)) or (inputs(197)));
    layer0_outputs(1750) <= (inputs(219)) or (inputs(171));
    layer0_outputs(1751) <= not(inputs(13));
    layer0_outputs(1752) <= not((inputs(105)) or (inputs(28)));
    layer0_outputs(1753) <= not((inputs(134)) and (inputs(231)));
    layer0_outputs(1754) <= (inputs(75)) xor (inputs(109));
    layer0_outputs(1755) <= not(inputs(211));
    layer0_outputs(1756) <= (inputs(65)) and not (inputs(63));
    layer0_outputs(1757) <= (inputs(187)) or (inputs(193));
    layer0_outputs(1758) <= not(inputs(44));
    layer0_outputs(1759) <= not(inputs(43)) or (inputs(221));
    layer0_outputs(1760) <= not(inputs(234));
    layer0_outputs(1761) <= not((inputs(253)) or (inputs(130)));
    layer0_outputs(1762) <= not(inputs(72));
    layer0_outputs(1763) <= not((inputs(51)) or (inputs(151)));
    layer0_outputs(1764) <= inputs(144);
    layer0_outputs(1765) <= not(inputs(135)) or (inputs(32));
    layer0_outputs(1766) <= not((inputs(108)) xor (inputs(39)));
    layer0_outputs(1767) <= (inputs(247)) or (inputs(100));
    layer0_outputs(1768) <= '0';
    layer0_outputs(1769) <= inputs(133);
    layer0_outputs(1770) <= (inputs(87)) and not (inputs(126));
    layer0_outputs(1771) <= not((inputs(127)) or (inputs(49)));
    layer0_outputs(1772) <= inputs(98);
    layer0_outputs(1773) <= (inputs(210)) and not (inputs(83));
    layer0_outputs(1774) <= not(inputs(39)) or (inputs(195));
    layer0_outputs(1775) <= inputs(145);
    layer0_outputs(1776) <= not((inputs(237)) xor (inputs(172)));
    layer0_outputs(1777) <= not((inputs(201)) or (inputs(195)));
    layer0_outputs(1778) <= not((inputs(114)) or (inputs(70)));
    layer0_outputs(1779) <= not(inputs(83));
    layer0_outputs(1780) <= not(inputs(23)) or (inputs(159));
    layer0_outputs(1781) <= not(inputs(51)) or (inputs(101));
    layer0_outputs(1782) <= inputs(190);
    layer0_outputs(1783) <= not((inputs(71)) or (inputs(89)));
    layer0_outputs(1784) <= (inputs(30)) or (inputs(77));
    layer0_outputs(1785) <= not((inputs(9)) and (inputs(69)));
    layer0_outputs(1786) <= (inputs(78)) or (inputs(45));
    layer0_outputs(1787) <= (inputs(30)) or (inputs(238));
    layer0_outputs(1788) <= not(inputs(55));
    layer0_outputs(1789) <= inputs(78);
    layer0_outputs(1790) <= not(inputs(34)) or (inputs(243));
    layer0_outputs(1791) <= not(inputs(230)) or (inputs(79));
    layer0_outputs(1792) <= inputs(201);
    layer0_outputs(1793) <= inputs(78);
    layer0_outputs(1794) <= inputs(189);
    layer0_outputs(1795) <= (inputs(139)) and not (inputs(40));
    layer0_outputs(1796) <= (inputs(238)) xor (inputs(151));
    layer0_outputs(1797) <= not(inputs(108));
    layer0_outputs(1798) <= not((inputs(172)) xor (inputs(180)));
    layer0_outputs(1799) <= (inputs(137)) and not (inputs(113));
    layer0_outputs(1800) <= (inputs(254)) or (inputs(132));
    layer0_outputs(1801) <= not(inputs(117));
    layer0_outputs(1802) <= not((inputs(0)) or (inputs(91)));
    layer0_outputs(1803) <= not((inputs(254)) or (inputs(68)));
    layer0_outputs(1804) <= not((inputs(37)) or (inputs(227)));
    layer0_outputs(1805) <= not((inputs(229)) or (inputs(243)));
    layer0_outputs(1806) <= not(inputs(186)) or (inputs(31));
    layer0_outputs(1807) <= (inputs(177)) xor (inputs(233));
    layer0_outputs(1808) <= inputs(29);
    layer0_outputs(1809) <= not((inputs(242)) or (inputs(173)));
    layer0_outputs(1810) <= not(inputs(107));
    layer0_outputs(1811) <= inputs(253);
    layer0_outputs(1812) <= not((inputs(162)) or (inputs(122)));
    layer0_outputs(1813) <= (inputs(53)) and not (inputs(238));
    layer0_outputs(1814) <= (inputs(113)) and not (inputs(50));
    layer0_outputs(1815) <= (inputs(99)) and not (inputs(108));
    layer0_outputs(1816) <= not((inputs(234)) or (inputs(184)));
    layer0_outputs(1817) <= not(inputs(68));
    layer0_outputs(1818) <= not((inputs(126)) or (inputs(198)));
    layer0_outputs(1819) <= not((inputs(109)) or (inputs(114)));
    layer0_outputs(1820) <= not((inputs(28)) xor (inputs(129)));
    layer0_outputs(1821) <= (inputs(152)) xor (inputs(139));
    layer0_outputs(1822) <= not((inputs(106)) xor (inputs(95)));
    layer0_outputs(1823) <= (inputs(211)) and not (inputs(46));
    layer0_outputs(1824) <= (inputs(101)) and not (inputs(142));
    layer0_outputs(1825) <= (inputs(191)) xor (inputs(43));
    layer0_outputs(1826) <= inputs(235);
    layer0_outputs(1827) <= not((inputs(114)) or (inputs(198)));
    layer0_outputs(1828) <= not((inputs(124)) xor (inputs(165)));
    layer0_outputs(1829) <= (inputs(62)) and (inputs(62));
    layer0_outputs(1830) <= (inputs(176)) or (inputs(156));
    layer0_outputs(1831) <= '1';
    layer0_outputs(1832) <= (inputs(15)) and not (inputs(26));
    layer0_outputs(1833) <= not(inputs(231)) or (inputs(46));
    layer0_outputs(1834) <= not(inputs(76));
    layer0_outputs(1835) <= not((inputs(41)) xor (inputs(74)));
    layer0_outputs(1836) <= (inputs(219)) xor (inputs(171));
    layer0_outputs(1837) <= (inputs(214)) and (inputs(201));
    layer0_outputs(1838) <= inputs(234);
    layer0_outputs(1839) <= inputs(213);
    layer0_outputs(1840) <= not(inputs(169));
    layer0_outputs(1841) <= inputs(115);
    layer0_outputs(1842) <= (inputs(190)) and (inputs(174));
    layer0_outputs(1843) <= (inputs(253)) and not (inputs(65));
    layer0_outputs(1844) <= inputs(248);
    layer0_outputs(1845) <= inputs(231);
    layer0_outputs(1846) <= inputs(57);
    layer0_outputs(1847) <= (inputs(83)) and not (inputs(87));
    layer0_outputs(1848) <= (inputs(155)) and (inputs(118));
    layer0_outputs(1849) <= not((inputs(143)) xor (inputs(123)));
    layer0_outputs(1850) <= (inputs(24)) and not (inputs(202));
    layer0_outputs(1851) <= not((inputs(130)) xor (inputs(101)));
    layer0_outputs(1852) <= (inputs(79)) and not (inputs(100));
    layer0_outputs(1853) <= (inputs(199)) or (inputs(223));
    layer0_outputs(1854) <= inputs(238);
    layer0_outputs(1855) <= not((inputs(134)) xor (inputs(56)));
    layer0_outputs(1856) <= inputs(211);
    layer0_outputs(1857) <= (inputs(90)) or (inputs(174));
    layer0_outputs(1858) <= (inputs(53)) or (inputs(78));
    layer0_outputs(1859) <= not(inputs(108));
    layer0_outputs(1860) <= not((inputs(80)) or (inputs(99)));
    layer0_outputs(1861) <= not(inputs(51)) or (inputs(242));
    layer0_outputs(1862) <= not(inputs(201)) or (inputs(13));
    layer0_outputs(1863) <= not(inputs(189));
    layer0_outputs(1864) <= not((inputs(81)) xor (inputs(151)));
    layer0_outputs(1865) <= not(inputs(45)) or (inputs(177));
    layer0_outputs(1866) <= not(inputs(194)) or (inputs(159));
    layer0_outputs(1867) <= (inputs(247)) or (inputs(251));
    layer0_outputs(1868) <= (inputs(116)) and not (inputs(159));
    layer0_outputs(1869) <= not(inputs(38)) or (inputs(63));
    layer0_outputs(1870) <= (inputs(179)) and not (inputs(31));
    layer0_outputs(1871) <= (inputs(144)) or (inputs(55));
    layer0_outputs(1872) <= inputs(130);
    layer0_outputs(1873) <= inputs(210);
    layer0_outputs(1874) <= not(inputs(132));
    layer0_outputs(1875) <= not((inputs(99)) xor (inputs(5)));
    layer0_outputs(1876) <= (inputs(247)) and not (inputs(81));
    layer0_outputs(1877) <= not((inputs(5)) or (inputs(215)));
    layer0_outputs(1878) <= (inputs(189)) or (inputs(216));
    layer0_outputs(1879) <= not(inputs(209));
    layer0_outputs(1880) <= not(inputs(14)) or (inputs(210));
    layer0_outputs(1881) <= (inputs(162)) xor (inputs(200));
    layer0_outputs(1882) <= not((inputs(152)) xor (inputs(170)));
    layer0_outputs(1883) <= not((inputs(27)) xor (inputs(186)));
    layer0_outputs(1884) <= (inputs(183)) and not (inputs(158));
    layer0_outputs(1885) <= not(inputs(148)) or (inputs(221));
    layer0_outputs(1886) <= inputs(50);
    layer0_outputs(1887) <= not((inputs(5)) xor (inputs(8)));
    layer0_outputs(1888) <= (inputs(155)) and not (inputs(204));
    layer0_outputs(1889) <= not(inputs(161));
    layer0_outputs(1890) <= not(inputs(176));
    layer0_outputs(1891) <= (inputs(1)) or (inputs(2));
    layer0_outputs(1892) <= not((inputs(149)) or (inputs(243)));
    layer0_outputs(1893) <= (inputs(78)) and not (inputs(54));
    layer0_outputs(1894) <= (inputs(54)) and not (inputs(41));
    layer0_outputs(1895) <= inputs(59);
    layer0_outputs(1896) <= not(inputs(180)) or (inputs(109));
    layer0_outputs(1897) <= (inputs(60)) and not (inputs(182));
    layer0_outputs(1898) <= not((inputs(142)) or (inputs(49)));
    layer0_outputs(1899) <= (inputs(203)) and not (inputs(97));
    layer0_outputs(1900) <= not(inputs(205));
    layer0_outputs(1901) <= not((inputs(70)) xor (inputs(68)));
    layer0_outputs(1902) <= (inputs(75)) xor (inputs(21));
    layer0_outputs(1903) <= (inputs(52)) or (inputs(151));
    layer0_outputs(1904) <= not((inputs(68)) xor (inputs(8)));
    layer0_outputs(1905) <= inputs(76);
    layer0_outputs(1906) <= (inputs(176)) and not (inputs(126));
    layer0_outputs(1907) <= not((inputs(230)) or (inputs(247)));
    layer0_outputs(1908) <= (inputs(251)) and not (inputs(127));
    layer0_outputs(1909) <= not(inputs(103));
    layer0_outputs(1910) <= inputs(104);
    layer0_outputs(1911) <= (inputs(53)) and not (inputs(28));
    layer0_outputs(1912) <= inputs(171);
    layer0_outputs(1913) <= not((inputs(236)) or (inputs(222)));
    layer0_outputs(1914) <= (inputs(219)) xor (inputs(78));
    layer0_outputs(1915) <= not(inputs(94));
    layer0_outputs(1916) <= not((inputs(169)) or (inputs(208)));
    layer0_outputs(1917) <= not((inputs(3)) or (inputs(107)));
    layer0_outputs(1918) <= (inputs(124)) xor (inputs(218));
    layer0_outputs(1919) <= not((inputs(161)) and (inputs(208)));
    layer0_outputs(1920) <= (inputs(122)) and not (inputs(197));
    layer0_outputs(1921) <= (inputs(120)) and not (inputs(179));
    layer0_outputs(1922) <= inputs(163);
    layer0_outputs(1923) <= not((inputs(102)) xor (inputs(56)));
    layer0_outputs(1924) <= (inputs(194)) and not (inputs(45));
    layer0_outputs(1925) <= inputs(21);
    layer0_outputs(1926) <= not((inputs(133)) xor (inputs(181)));
    layer0_outputs(1927) <= not((inputs(132)) or (inputs(232)));
    layer0_outputs(1928) <= (inputs(192)) and (inputs(55));
    layer0_outputs(1929) <= (inputs(127)) or (inputs(171));
    layer0_outputs(1930) <= inputs(86);
    layer0_outputs(1931) <= not(inputs(157)) or (inputs(95));
    layer0_outputs(1932) <= (inputs(168)) or (inputs(201));
    layer0_outputs(1933) <= inputs(200);
    layer0_outputs(1934) <= (inputs(197)) xor (inputs(243));
    layer0_outputs(1935) <= not((inputs(167)) or (inputs(55)));
    layer0_outputs(1936) <= not((inputs(126)) or (inputs(130)));
    layer0_outputs(1937) <= (inputs(153)) xor (inputs(134));
    layer0_outputs(1938) <= not(inputs(151));
    layer0_outputs(1939) <= inputs(208);
    layer0_outputs(1940) <= not(inputs(13)) or (inputs(237));
    layer0_outputs(1941) <= not(inputs(95));
    layer0_outputs(1942) <= not((inputs(97)) or (inputs(62)));
    layer0_outputs(1943) <= not(inputs(137)) or (inputs(127));
    layer0_outputs(1944) <= not(inputs(75)) or (inputs(32));
    layer0_outputs(1945) <= (inputs(132)) xor (inputs(226));
    layer0_outputs(1946) <= not(inputs(86));
    layer0_outputs(1947) <= (inputs(222)) or (inputs(240));
    layer0_outputs(1948) <= not(inputs(13));
    layer0_outputs(1949) <= not((inputs(63)) or (inputs(34)));
    layer0_outputs(1950) <= not(inputs(32)) or (inputs(161));
    layer0_outputs(1951) <= inputs(165);
    layer0_outputs(1952) <= not((inputs(190)) or (inputs(145)));
    layer0_outputs(1953) <= not((inputs(91)) or (inputs(177)));
    layer0_outputs(1954) <= (inputs(199)) xor (inputs(13));
    layer0_outputs(1955) <= inputs(165);
    layer0_outputs(1956) <= not(inputs(217)) or (inputs(0));
    layer0_outputs(1957) <= not(inputs(122)) or (inputs(52));
    layer0_outputs(1958) <= inputs(108);
    layer0_outputs(1959) <= not((inputs(89)) xor (inputs(136)));
    layer0_outputs(1960) <= not(inputs(86));
    layer0_outputs(1961) <= inputs(218);
    layer0_outputs(1962) <= (inputs(99)) or (inputs(231));
    layer0_outputs(1963) <= not(inputs(91));
    layer0_outputs(1964) <= not(inputs(40)) or (inputs(169));
    layer0_outputs(1965) <= not(inputs(12));
    layer0_outputs(1966) <= (inputs(225)) and not (inputs(81));
    layer0_outputs(1967) <= not((inputs(219)) xor (inputs(252)));
    layer0_outputs(1968) <= inputs(249);
    layer0_outputs(1969) <= not(inputs(210)) or (inputs(171));
    layer0_outputs(1970) <= inputs(85);
    layer0_outputs(1971) <= not((inputs(148)) xor (inputs(212)));
    layer0_outputs(1972) <= not(inputs(148));
    layer0_outputs(1973) <= '0';
    layer0_outputs(1974) <= (inputs(44)) or (inputs(168));
    layer0_outputs(1975) <= inputs(110);
    layer0_outputs(1976) <= inputs(245);
    layer0_outputs(1977) <= (inputs(131)) xor (inputs(149));
    layer0_outputs(1978) <= not((inputs(118)) or (inputs(215)));
    layer0_outputs(1979) <= not((inputs(248)) xor (inputs(51)));
    layer0_outputs(1980) <= inputs(0);
    layer0_outputs(1981) <= inputs(179);
    layer0_outputs(1982) <= (inputs(60)) and not (inputs(255));
    layer0_outputs(1983) <= not(inputs(75));
    layer0_outputs(1984) <= not(inputs(28)) or (inputs(86));
    layer0_outputs(1985) <= not((inputs(94)) xor (inputs(46)));
    layer0_outputs(1986) <= not((inputs(138)) xor (inputs(157)));
    layer0_outputs(1987) <= (inputs(199)) and not (inputs(139));
    layer0_outputs(1988) <= not((inputs(153)) or (inputs(203)));
    layer0_outputs(1989) <= inputs(149);
    layer0_outputs(1990) <= (inputs(191)) or (inputs(117));
    layer0_outputs(1991) <= not((inputs(114)) xor (inputs(148)));
    layer0_outputs(1992) <= not(inputs(117)) or (inputs(240));
    layer0_outputs(1993) <= (inputs(212)) and not (inputs(185));
    layer0_outputs(1994) <= not((inputs(81)) and (inputs(130)));
    layer0_outputs(1995) <= (inputs(250)) or (inputs(56));
    layer0_outputs(1996) <= not(inputs(8));
    layer0_outputs(1997) <= inputs(130);
    layer0_outputs(1998) <= not(inputs(179));
    layer0_outputs(1999) <= (inputs(62)) and (inputs(111));
    layer0_outputs(2000) <= not(inputs(96));
    layer0_outputs(2001) <= (inputs(82)) xor (inputs(87));
    layer0_outputs(2002) <= not((inputs(23)) xor (inputs(172)));
    layer0_outputs(2003) <= not(inputs(197));
    layer0_outputs(2004) <= not(inputs(215)) or (inputs(23));
    layer0_outputs(2005) <= (inputs(234)) or (inputs(180));
    layer0_outputs(2006) <= not(inputs(197)) or (inputs(108));
    layer0_outputs(2007) <= not((inputs(150)) xor (inputs(68)));
    layer0_outputs(2008) <= (inputs(132)) xor (inputs(163));
    layer0_outputs(2009) <= not((inputs(103)) xor (inputs(210)));
    layer0_outputs(2010) <= not(inputs(76));
    layer0_outputs(2011) <= (inputs(60)) and not (inputs(49));
    layer0_outputs(2012) <= (inputs(46)) xor (inputs(176));
    layer0_outputs(2013) <= not(inputs(100));
    layer0_outputs(2014) <= not((inputs(1)) and (inputs(174)));
    layer0_outputs(2015) <= not(inputs(11)) or (inputs(61));
    layer0_outputs(2016) <= (inputs(117)) xor (inputs(187));
    layer0_outputs(2017) <= inputs(116);
    layer0_outputs(2018) <= not(inputs(56));
    layer0_outputs(2019) <= (inputs(141)) and (inputs(58));
    layer0_outputs(2020) <= inputs(58);
    layer0_outputs(2021) <= not(inputs(127));
    layer0_outputs(2022) <= not((inputs(109)) xor (inputs(154)));
    layer0_outputs(2023) <= not((inputs(190)) xor (inputs(96)));
    layer0_outputs(2024) <= inputs(248);
    layer0_outputs(2025) <= (inputs(157)) or (inputs(159));
    layer0_outputs(2026) <= not(inputs(106)) or (inputs(128));
    layer0_outputs(2027) <= (inputs(92)) and not (inputs(145));
    layer0_outputs(2028) <= inputs(113);
    layer0_outputs(2029) <= '1';
    layer0_outputs(2030) <= not(inputs(50));
    layer0_outputs(2031) <= (inputs(195)) or (inputs(167));
    layer0_outputs(2032) <= inputs(130);
    layer0_outputs(2033) <= not(inputs(145));
    layer0_outputs(2034) <= inputs(25);
    layer0_outputs(2035) <= inputs(6);
    layer0_outputs(2036) <= (inputs(230)) and not (inputs(85));
    layer0_outputs(2037) <= not(inputs(112));
    layer0_outputs(2038) <= (inputs(184)) and not (inputs(19));
    layer0_outputs(2039) <= not((inputs(226)) or (inputs(40)));
    layer0_outputs(2040) <= (inputs(121)) xor (inputs(182));
    layer0_outputs(2041) <= (inputs(214)) and not (inputs(96));
    layer0_outputs(2042) <= inputs(146);
    layer0_outputs(2043) <= (inputs(135)) xor (inputs(17));
    layer0_outputs(2044) <= (inputs(34)) xor (inputs(244));
    layer0_outputs(2045) <= not((inputs(187)) xor (inputs(111)));
    layer0_outputs(2046) <= (inputs(156)) xor (inputs(186));
    layer0_outputs(2047) <= (inputs(117)) and not (inputs(252));
    layer0_outputs(2048) <= not(inputs(228)) or (inputs(134));
    layer0_outputs(2049) <= (inputs(139)) and not (inputs(182));
    layer0_outputs(2050) <= not(inputs(70));
    layer0_outputs(2051) <= not((inputs(244)) or (inputs(16)));
    layer0_outputs(2052) <= not(inputs(7)) or (inputs(201));
    layer0_outputs(2053) <= '0';
    layer0_outputs(2054) <= (inputs(222)) and (inputs(216));
    layer0_outputs(2055) <= not((inputs(101)) xor (inputs(113)));
    layer0_outputs(2056) <= (inputs(217)) xor (inputs(162));
    layer0_outputs(2057) <= inputs(1);
    layer0_outputs(2058) <= (inputs(88)) xor (inputs(10));
    layer0_outputs(2059) <= (inputs(220)) xor (inputs(150));
    layer0_outputs(2060) <= (inputs(216)) xor (inputs(41));
    layer0_outputs(2061) <= '1';
    layer0_outputs(2062) <= inputs(45);
    layer0_outputs(2063) <= not(inputs(39));
    layer0_outputs(2064) <= (inputs(124)) or (inputs(147));
    layer0_outputs(2065) <= inputs(66);
    layer0_outputs(2066) <= inputs(46);
    layer0_outputs(2067) <= not((inputs(235)) xor (inputs(76)));
    layer0_outputs(2068) <= not(inputs(25)) or (inputs(112));
    layer0_outputs(2069) <= not((inputs(39)) xor (inputs(232)));
    layer0_outputs(2070) <= (inputs(19)) or (inputs(34));
    layer0_outputs(2071) <= not((inputs(96)) xor (inputs(63)));
    layer0_outputs(2072) <= (inputs(63)) or (inputs(193));
    layer0_outputs(2073) <= inputs(162);
    layer0_outputs(2074) <= (inputs(43)) xor (inputs(239));
    layer0_outputs(2075) <= inputs(187);
    layer0_outputs(2076) <= (inputs(67)) and not (inputs(33));
    layer0_outputs(2077) <= (inputs(70)) and not (inputs(22));
    layer0_outputs(2078) <= not(inputs(14));
    layer0_outputs(2079) <= inputs(116);
    layer0_outputs(2080) <= not((inputs(176)) xor (inputs(244)));
    layer0_outputs(2081) <= not(inputs(59)) or (inputs(176));
    layer0_outputs(2082) <= (inputs(205)) xor (inputs(213));
    layer0_outputs(2083) <= (inputs(117)) and not (inputs(36));
    layer0_outputs(2084) <= (inputs(113)) or (inputs(114));
    layer0_outputs(2085) <= (inputs(18)) and (inputs(247));
    layer0_outputs(2086) <= not(inputs(236));
    layer0_outputs(2087) <= not(inputs(186)) or (inputs(251));
    layer0_outputs(2088) <= not((inputs(226)) or (inputs(211)));
    layer0_outputs(2089) <= (inputs(67)) or (inputs(19));
    layer0_outputs(2090) <= not(inputs(208)) or (inputs(58));
    layer0_outputs(2091) <= not(inputs(118));
    layer0_outputs(2092) <= not((inputs(77)) or (inputs(180)));
    layer0_outputs(2093) <= inputs(245);
    layer0_outputs(2094) <= not(inputs(86));
    layer0_outputs(2095) <= (inputs(4)) xor (inputs(120));
    layer0_outputs(2096) <= not((inputs(39)) and (inputs(42)));
    layer0_outputs(2097) <= (inputs(53)) or (inputs(79));
    layer0_outputs(2098) <= not(inputs(41));
    layer0_outputs(2099) <= (inputs(118)) xor (inputs(26));
    layer0_outputs(2100) <= not(inputs(97));
    layer0_outputs(2101) <= not((inputs(248)) xor (inputs(63)));
    layer0_outputs(2102) <= inputs(220);
    layer0_outputs(2103) <= inputs(197);
    layer0_outputs(2104) <= (inputs(52)) and (inputs(233));
    layer0_outputs(2105) <= (inputs(42)) or (inputs(63));
    layer0_outputs(2106) <= (inputs(134)) xor (inputs(204));
    layer0_outputs(2107) <= not(inputs(147)) or (inputs(62));
    layer0_outputs(2108) <= not((inputs(83)) xor (inputs(188)));
    layer0_outputs(2109) <= (inputs(26)) and not (inputs(134));
    layer0_outputs(2110) <= (inputs(137)) and not (inputs(244));
    layer0_outputs(2111) <= (inputs(142)) and not (inputs(176));
    layer0_outputs(2112) <= not(inputs(135));
    layer0_outputs(2113) <= (inputs(129)) or (inputs(189));
    layer0_outputs(2114) <= inputs(163);
    layer0_outputs(2115) <= not((inputs(4)) xor (inputs(119)));
    layer0_outputs(2116) <= not(inputs(85));
    layer0_outputs(2117) <= not(inputs(165)) or (inputs(86));
    layer0_outputs(2118) <= (inputs(171)) and not (inputs(1));
    layer0_outputs(2119) <= not((inputs(161)) or (inputs(72)));
    layer0_outputs(2120) <= '0';
    layer0_outputs(2121) <= not(inputs(43)) or (inputs(178));
    layer0_outputs(2122) <= inputs(231);
    layer0_outputs(2123) <= (inputs(207)) and not (inputs(1));
    layer0_outputs(2124) <= (inputs(16)) xor (inputs(120));
    layer0_outputs(2125) <= not(inputs(177)) or (inputs(186));
    layer0_outputs(2126) <= not(inputs(215)) or (inputs(82));
    layer0_outputs(2127) <= not(inputs(24));
    layer0_outputs(2128) <= not(inputs(138)) or (inputs(32));
    layer0_outputs(2129) <= not(inputs(115)) or (inputs(174));
    layer0_outputs(2130) <= not(inputs(6));
    layer0_outputs(2131) <= (inputs(141)) xor (inputs(191));
    layer0_outputs(2132) <= (inputs(140)) xor (inputs(29));
    layer0_outputs(2133) <= inputs(22);
    layer0_outputs(2134) <= not(inputs(217));
    layer0_outputs(2135) <= not((inputs(228)) and (inputs(169)));
    layer0_outputs(2136) <= not(inputs(35));
    layer0_outputs(2137) <= not(inputs(246)) or (inputs(49));
    layer0_outputs(2138) <= not((inputs(229)) or (inputs(84)));
    layer0_outputs(2139) <= not(inputs(88));
    layer0_outputs(2140) <= (inputs(30)) xor (inputs(131));
    layer0_outputs(2141) <= not(inputs(150)) or (inputs(88));
    layer0_outputs(2142) <= not((inputs(122)) and (inputs(90)));
    layer0_outputs(2143) <= not(inputs(162));
    layer0_outputs(2144) <= not(inputs(107));
    layer0_outputs(2145) <= inputs(238);
    layer0_outputs(2146) <= not((inputs(111)) xor (inputs(33)));
    layer0_outputs(2147) <= (inputs(224)) and (inputs(95));
    layer0_outputs(2148) <= inputs(231);
    layer0_outputs(2149) <= (inputs(39)) and (inputs(33));
    layer0_outputs(2150) <= not(inputs(146)) or (inputs(97));
    layer0_outputs(2151) <= not(inputs(43)) or (inputs(254));
    layer0_outputs(2152) <= not((inputs(212)) xor (inputs(180)));
    layer0_outputs(2153) <= (inputs(33)) or (inputs(38));
    layer0_outputs(2154) <= inputs(201);
    layer0_outputs(2155) <= (inputs(149)) or (inputs(243));
    layer0_outputs(2156) <= not(inputs(110));
    layer0_outputs(2157) <= (inputs(89)) xor (inputs(80));
    layer0_outputs(2158) <= (inputs(53)) and not (inputs(192));
    layer0_outputs(2159) <= not(inputs(196)) or (inputs(49));
    layer0_outputs(2160) <= (inputs(219)) and not (inputs(55));
    layer0_outputs(2161) <= inputs(167);
    layer0_outputs(2162) <= not(inputs(244));
    layer0_outputs(2163) <= not((inputs(192)) xor (inputs(133)));
    layer0_outputs(2164) <= not((inputs(107)) or (inputs(61)));
    layer0_outputs(2165) <= not(inputs(105));
    layer0_outputs(2166) <= '0';
    layer0_outputs(2167) <= (inputs(134)) or (inputs(247));
    layer0_outputs(2168) <= not(inputs(154));
    layer0_outputs(2169) <= not((inputs(37)) or (inputs(194)));
    layer0_outputs(2170) <= not((inputs(145)) or (inputs(51)));
    layer0_outputs(2171) <= inputs(120);
    layer0_outputs(2172) <= inputs(185);
    layer0_outputs(2173) <= (inputs(116)) xor (inputs(87));
    layer0_outputs(2174) <= (inputs(98)) or (inputs(219));
    layer0_outputs(2175) <= not(inputs(229));
    layer0_outputs(2176) <= not(inputs(104));
    layer0_outputs(2177) <= not((inputs(88)) and (inputs(103)));
    layer0_outputs(2178) <= not((inputs(156)) or (inputs(190)));
    layer0_outputs(2179) <= inputs(39);
    layer0_outputs(2180) <= (inputs(126)) or (inputs(26));
    layer0_outputs(2181) <= (inputs(74)) and not (inputs(87));
    layer0_outputs(2182) <= not(inputs(55));
    layer0_outputs(2183) <= not(inputs(8)) or (inputs(148));
    layer0_outputs(2184) <= inputs(192);
    layer0_outputs(2185) <= (inputs(186)) and not (inputs(170));
    layer0_outputs(2186) <= not(inputs(113));
    layer0_outputs(2187) <= not((inputs(202)) xor (inputs(123)));
    layer0_outputs(2188) <= (inputs(2)) or (inputs(190));
    layer0_outputs(2189) <= not((inputs(145)) or (inputs(112)));
    layer0_outputs(2190) <= (inputs(237)) xor (inputs(188));
    layer0_outputs(2191) <= (inputs(211)) or (inputs(33));
    layer0_outputs(2192) <= (inputs(52)) and not (inputs(141));
    layer0_outputs(2193) <= not((inputs(85)) or (inputs(116)));
    layer0_outputs(2194) <= inputs(161);
    layer0_outputs(2195) <= not(inputs(100)) or (inputs(220));
    layer0_outputs(2196) <= inputs(188);
    layer0_outputs(2197) <= inputs(240);
    layer0_outputs(2198) <= not((inputs(4)) or (inputs(140)));
    layer0_outputs(2199) <= (inputs(177)) xor (inputs(243));
    layer0_outputs(2200) <= (inputs(100)) xor (inputs(86));
    layer0_outputs(2201) <= (inputs(107)) or (inputs(171));
    layer0_outputs(2202) <= not((inputs(175)) or (inputs(116)));
    layer0_outputs(2203) <= (inputs(55)) or (inputs(44));
    layer0_outputs(2204) <= not(inputs(58)) or (inputs(81));
    layer0_outputs(2205) <= (inputs(49)) or (inputs(254));
    layer0_outputs(2206) <= inputs(91);
    layer0_outputs(2207) <= (inputs(208)) xor (inputs(12));
    layer0_outputs(2208) <= inputs(100);
    layer0_outputs(2209) <= (inputs(134)) and not (inputs(19));
    layer0_outputs(2210) <= not(inputs(7)) or (inputs(255));
    layer0_outputs(2211) <= inputs(69);
    layer0_outputs(2212) <= (inputs(61)) and (inputs(77));
    layer0_outputs(2213) <= (inputs(24)) and not (inputs(158));
    layer0_outputs(2214) <= not(inputs(28));
    layer0_outputs(2215) <= (inputs(66)) or (inputs(13));
    layer0_outputs(2216) <= (inputs(252)) or (inputs(71));
    layer0_outputs(2217) <= (inputs(167)) or (inputs(73));
    layer0_outputs(2218) <= (inputs(254)) or (inputs(56));
    layer0_outputs(2219) <= inputs(174);
    layer0_outputs(2220) <= (inputs(151)) and not (inputs(0));
    layer0_outputs(2221) <= (inputs(104)) and not (inputs(4));
    layer0_outputs(2222) <= (inputs(6)) and (inputs(242));
    layer0_outputs(2223) <= not((inputs(240)) or (inputs(21)));
    layer0_outputs(2224) <= not((inputs(110)) or (inputs(220)));
    layer0_outputs(2225) <= not((inputs(48)) or (inputs(209)));
    layer0_outputs(2226) <= (inputs(172)) xor (inputs(69));
    layer0_outputs(2227) <= (inputs(145)) and (inputs(66));
    layer0_outputs(2228) <= (inputs(127)) or (inputs(248));
    layer0_outputs(2229) <= not(inputs(220));
    layer0_outputs(2230) <= not(inputs(120)) or (inputs(239));
    layer0_outputs(2231) <= (inputs(201)) or (inputs(206));
    layer0_outputs(2232) <= (inputs(164)) or (inputs(254));
    layer0_outputs(2233) <= not(inputs(235));
    layer0_outputs(2234) <= not(inputs(188));
    layer0_outputs(2235) <= inputs(110);
    layer0_outputs(2236) <= not(inputs(246));
    layer0_outputs(2237) <= (inputs(170)) xor (inputs(110));
    layer0_outputs(2238) <= not((inputs(196)) xor (inputs(209)));
    layer0_outputs(2239) <= (inputs(42)) xor (inputs(69));
    layer0_outputs(2240) <= (inputs(179)) and not (inputs(14));
    layer0_outputs(2241) <= (inputs(112)) or (inputs(12));
    layer0_outputs(2242) <= inputs(102);
    layer0_outputs(2243) <= inputs(3);
    layer0_outputs(2244) <= (inputs(12)) and not (inputs(224));
    layer0_outputs(2245) <= inputs(180);
    layer0_outputs(2246) <= not((inputs(148)) or (inputs(85)));
    layer0_outputs(2247) <= not((inputs(160)) or (inputs(177)));
    layer0_outputs(2248) <= not(inputs(231));
    layer0_outputs(2249) <= not((inputs(61)) or (inputs(115)));
    layer0_outputs(2250) <= (inputs(56)) and not (inputs(157));
    layer0_outputs(2251) <= not(inputs(118)) or (inputs(65));
    layer0_outputs(2252) <= not((inputs(37)) xor (inputs(54)));
    layer0_outputs(2253) <= not(inputs(152));
    layer0_outputs(2254) <= not((inputs(108)) or (inputs(254)));
    layer0_outputs(2255) <= not((inputs(61)) or (inputs(150)));
    layer0_outputs(2256) <= (inputs(232)) xor (inputs(208));
    layer0_outputs(2257) <= inputs(54);
    layer0_outputs(2258) <= inputs(143);
    layer0_outputs(2259) <= not(inputs(164)) or (inputs(17));
    layer0_outputs(2260) <= inputs(245);
    layer0_outputs(2261) <= (inputs(54)) xor (inputs(9));
    layer0_outputs(2262) <= inputs(254);
    layer0_outputs(2263) <= '1';
    layer0_outputs(2264) <= not(inputs(247));
    layer0_outputs(2265) <= (inputs(82)) xor (inputs(85));
    layer0_outputs(2266) <= not(inputs(215)) or (inputs(65));
    layer0_outputs(2267) <= (inputs(132)) xor (inputs(119));
    layer0_outputs(2268) <= (inputs(123)) and not (inputs(29));
    layer0_outputs(2269) <= (inputs(100)) and not (inputs(64));
    layer0_outputs(2270) <= (inputs(100)) and not (inputs(208));
    layer0_outputs(2271) <= not(inputs(245));
    layer0_outputs(2272) <= not(inputs(193));
    layer0_outputs(2273) <= not(inputs(35));
    layer0_outputs(2274) <= not(inputs(70)) or (inputs(254));
    layer0_outputs(2275) <= not(inputs(126));
    layer0_outputs(2276) <= not((inputs(146)) xor (inputs(183)));
    layer0_outputs(2277) <= not((inputs(35)) and (inputs(78)));
    layer0_outputs(2278) <= inputs(104);
    layer0_outputs(2279) <= not((inputs(188)) xor (inputs(186)));
    layer0_outputs(2280) <= not(inputs(76)) or (inputs(216));
    layer0_outputs(2281) <= not((inputs(204)) xor (inputs(250)));
    layer0_outputs(2282) <= inputs(181);
    layer0_outputs(2283) <= (inputs(146)) and (inputs(114));
    layer0_outputs(2284) <= inputs(76);
    layer0_outputs(2285) <= not((inputs(21)) xor (inputs(143)));
    layer0_outputs(2286) <= not(inputs(8)) or (inputs(247));
    layer0_outputs(2287) <= inputs(92);
    layer0_outputs(2288) <= not((inputs(1)) or (inputs(237)));
    layer0_outputs(2289) <= not((inputs(155)) or (inputs(178)));
    layer0_outputs(2290) <= (inputs(215)) xor (inputs(168));
    layer0_outputs(2291) <= (inputs(12)) xor (inputs(241));
    layer0_outputs(2292) <= not(inputs(149));
    layer0_outputs(2293) <= (inputs(129)) xor (inputs(218));
    layer0_outputs(2294) <= inputs(25);
    layer0_outputs(2295) <= (inputs(194)) and not (inputs(162));
    layer0_outputs(2296) <= not(inputs(169)) or (inputs(3));
    layer0_outputs(2297) <= inputs(153);
    layer0_outputs(2298) <= (inputs(173)) or (inputs(176));
    layer0_outputs(2299) <= (inputs(27)) and (inputs(116));
    layer0_outputs(2300) <= inputs(178);
    layer0_outputs(2301) <= (inputs(28)) and not (inputs(197));
    layer0_outputs(2302) <= inputs(146);
    layer0_outputs(2303) <= not(inputs(141));
    layer0_outputs(2304) <= not((inputs(157)) or (inputs(127)));
    layer0_outputs(2305) <= inputs(22);
    layer0_outputs(2306) <= not(inputs(129));
    layer0_outputs(2307) <= (inputs(234)) and (inputs(156));
    layer0_outputs(2308) <= (inputs(47)) or (inputs(172));
    layer0_outputs(2309) <= not(inputs(6));
    layer0_outputs(2310) <= not((inputs(87)) and (inputs(58)));
    layer0_outputs(2311) <= (inputs(155)) or (inputs(46));
    layer0_outputs(2312) <= not(inputs(67));
    layer0_outputs(2313) <= (inputs(238)) or (inputs(194));
    layer0_outputs(2314) <= (inputs(223)) xor (inputs(54));
    layer0_outputs(2315) <= (inputs(24)) and not (inputs(227));
    layer0_outputs(2316) <= not(inputs(174));
    layer0_outputs(2317) <= not((inputs(201)) xor (inputs(156)));
    layer0_outputs(2318) <= not((inputs(173)) or (inputs(19)));
    layer0_outputs(2319) <= (inputs(21)) xor (inputs(190));
    layer0_outputs(2320) <= not((inputs(4)) xor (inputs(101)));
    layer0_outputs(2321) <= not(inputs(193)) or (inputs(18));
    layer0_outputs(2322) <= inputs(14);
    layer0_outputs(2323) <= not((inputs(175)) or (inputs(183)));
    layer0_outputs(2324) <= not((inputs(70)) xor (inputs(83)));
    layer0_outputs(2325) <= (inputs(159)) or (inputs(206));
    layer0_outputs(2326) <= not((inputs(91)) or (inputs(2)));
    layer0_outputs(2327) <= not(inputs(70)) or (inputs(1));
    layer0_outputs(2328) <= (inputs(24)) or (inputs(110));
    layer0_outputs(2329) <= not(inputs(129));
    layer0_outputs(2330) <= '0';
    layer0_outputs(2331) <= inputs(87);
    layer0_outputs(2332) <= (inputs(47)) and not (inputs(176));
    layer0_outputs(2333) <= inputs(22);
    layer0_outputs(2334) <= not(inputs(178)) or (inputs(252));
    layer0_outputs(2335) <= inputs(203);
    layer0_outputs(2336) <= (inputs(236)) xor (inputs(82));
    layer0_outputs(2337) <= not(inputs(52));
    layer0_outputs(2338) <= (inputs(26)) and not (inputs(104));
    layer0_outputs(2339) <= inputs(197);
    layer0_outputs(2340) <= not((inputs(173)) and (inputs(31)));
    layer0_outputs(2341) <= (inputs(9)) and not (inputs(253));
    layer0_outputs(2342) <= not(inputs(237));
    layer0_outputs(2343) <= not(inputs(113));
    layer0_outputs(2344) <= not(inputs(233)) or (inputs(77));
    layer0_outputs(2345) <= not((inputs(203)) or (inputs(231)));
    layer0_outputs(2346) <= not((inputs(102)) and (inputs(90)));
    layer0_outputs(2347) <= inputs(5);
    layer0_outputs(2348) <= not((inputs(157)) xor (inputs(201)));
    layer0_outputs(2349) <= (inputs(28)) xor (inputs(199));
    layer0_outputs(2350) <= (inputs(104)) and (inputs(162));
    layer0_outputs(2351) <= not(inputs(197));
    layer0_outputs(2352) <= inputs(83);
    layer0_outputs(2353) <= not((inputs(136)) or (inputs(36)));
    layer0_outputs(2354) <= (inputs(173)) xor (inputs(212));
    layer0_outputs(2355) <= (inputs(145)) xor (inputs(137));
    layer0_outputs(2356) <= not(inputs(94));
    layer0_outputs(2357) <= not((inputs(135)) or (inputs(82)));
    layer0_outputs(2358) <= (inputs(153)) and not (inputs(144));
    layer0_outputs(2359) <= not(inputs(106)) or (inputs(34));
    layer0_outputs(2360) <= inputs(120);
    layer0_outputs(2361) <= (inputs(241)) xor (inputs(141));
    layer0_outputs(2362) <= not(inputs(63)) or (inputs(123));
    layer0_outputs(2363) <= not(inputs(189));
    layer0_outputs(2364) <= inputs(33);
    layer0_outputs(2365) <= (inputs(26)) and not (inputs(214));
    layer0_outputs(2366) <= inputs(89);
    layer0_outputs(2367) <= not(inputs(54));
    layer0_outputs(2368) <= not(inputs(198));
    layer0_outputs(2369) <= not(inputs(136));
    layer0_outputs(2370) <= (inputs(219)) or (inputs(215));
    layer0_outputs(2371) <= not((inputs(69)) or (inputs(42)));
    layer0_outputs(2372) <= (inputs(166)) and not (inputs(188));
    layer0_outputs(2373) <= not((inputs(176)) or (inputs(249)));
    layer0_outputs(2374) <= (inputs(166)) or (inputs(143));
    layer0_outputs(2375) <= inputs(213);
    layer0_outputs(2376) <= (inputs(197)) and not (inputs(167));
    layer0_outputs(2377) <= inputs(229);
    layer0_outputs(2378) <= not(inputs(56));
    layer0_outputs(2379) <= not(inputs(88));
    layer0_outputs(2380) <= not(inputs(33));
    layer0_outputs(2381) <= not(inputs(169));
    layer0_outputs(2382) <= not(inputs(227)) or (inputs(201));
    layer0_outputs(2383) <= not((inputs(246)) and (inputs(180)));
    layer0_outputs(2384) <= not((inputs(159)) xor (inputs(147)));
    layer0_outputs(2385) <= not(inputs(39));
    layer0_outputs(2386) <= not((inputs(194)) xor (inputs(103)));
    layer0_outputs(2387) <= not((inputs(190)) xor (inputs(154)));
    layer0_outputs(2388) <= (inputs(173)) or (inputs(65));
    layer0_outputs(2389) <= inputs(121);
    layer0_outputs(2390) <= (inputs(120)) xor (inputs(61));
    layer0_outputs(2391) <= not((inputs(189)) or (inputs(220)));
    layer0_outputs(2392) <= not((inputs(146)) xor (inputs(184)));
    layer0_outputs(2393) <= not(inputs(74));
    layer0_outputs(2394) <= inputs(16);
    layer0_outputs(2395) <= inputs(69);
    layer0_outputs(2396) <= (inputs(206)) xor (inputs(187));
    layer0_outputs(2397) <= (inputs(126)) and not (inputs(240));
    layer0_outputs(2398) <= not(inputs(158));
    layer0_outputs(2399) <= not(inputs(25)) or (inputs(146));
    layer0_outputs(2400) <= inputs(228);
    layer0_outputs(2401) <= inputs(184);
    layer0_outputs(2402) <= (inputs(6)) or (inputs(95));
    layer0_outputs(2403) <= (inputs(48)) or (inputs(167));
    layer0_outputs(2404) <= inputs(233);
    layer0_outputs(2405) <= not(inputs(97));
    layer0_outputs(2406) <= (inputs(107)) and not (inputs(82));
    layer0_outputs(2407) <= not((inputs(94)) xor (inputs(204)));
    layer0_outputs(2408) <= not(inputs(104));
    layer0_outputs(2409) <= not(inputs(98));
    layer0_outputs(2410) <= (inputs(126)) xor (inputs(167));
    layer0_outputs(2411) <= inputs(27);
    layer0_outputs(2412) <= '0';
    layer0_outputs(2413) <= not(inputs(40));
    layer0_outputs(2414) <= not((inputs(209)) and (inputs(86)));
    layer0_outputs(2415) <= inputs(26);
    layer0_outputs(2416) <= not(inputs(165));
    layer0_outputs(2417) <= not(inputs(66)) or (inputs(106));
    layer0_outputs(2418) <= not(inputs(145));
    layer0_outputs(2419) <= not((inputs(30)) xor (inputs(17)));
    layer0_outputs(2420) <= not((inputs(164)) or (inputs(143)));
    layer0_outputs(2421) <= inputs(153);
    layer0_outputs(2422) <= not(inputs(88));
    layer0_outputs(2423) <= inputs(204);
    layer0_outputs(2424) <= not(inputs(37)) or (inputs(241));
    layer0_outputs(2425) <= not(inputs(164));
    layer0_outputs(2426) <= not((inputs(62)) or (inputs(123)));
    layer0_outputs(2427) <= not((inputs(104)) xor (inputs(162)));
    layer0_outputs(2428) <= not(inputs(137)) or (inputs(203));
    layer0_outputs(2429) <= not(inputs(72));
    layer0_outputs(2430) <= (inputs(3)) and not (inputs(66));
    layer0_outputs(2431) <= (inputs(213)) and not (inputs(187));
    layer0_outputs(2432) <= not(inputs(101)) or (inputs(16));
    layer0_outputs(2433) <= not((inputs(159)) xor (inputs(72)));
    layer0_outputs(2434) <= not(inputs(17)) or (inputs(29));
    layer0_outputs(2435) <= inputs(113);
    layer0_outputs(2436) <= (inputs(153)) or (inputs(152));
    layer0_outputs(2437) <= not(inputs(104));
    layer0_outputs(2438) <= not((inputs(148)) or (inputs(231)));
    layer0_outputs(2439) <= not((inputs(37)) xor (inputs(244)));
    layer0_outputs(2440) <= (inputs(25)) xor (inputs(193));
    layer0_outputs(2441) <= not(inputs(73));
    layer0_outputs(2442) <= not((inputs(166)) xor (inputs(115)));
    layer0_outputs(2443) <= inputs(25);
    layer0_outputs(2444) <= not(inputs(194));
    layer0_outputs(2445) <= (inputs(172)) and (inputs(75));
    layer0_outputs(2446) <= not((inputs(107)) xor (inputs(172)));
    layer0_outputs(2447) <= not((inputs(121)) or (inputs(163)));
    layer0_outputs(2448) <= (inputs(133)) and not (inputs(227));
    layer0_outputs(2449) <= not(inputs(69));
    layer0_outputs(2450) <= (inputs(202)) or (inputs(161));
    layer0_outputs(2451) <= inputs(34);
    layer0_outputs(2452) <= (inputs(9)) xor (inputs(189));
    layer0_outputs(2453) <= not(inputs(137)) or (inputs(212));
    layer0_outputs(2454) <= not((inputs(239)) xor (inputs(43)));
    layer0_outputs(2455) <= not((inputs(105)) and (inputs(7)));
    layer0_outputs(2456) <= (inputs(159)) xor (inputs(24));
    layer0_outputs(2457) <= inputs(100);
    layer0_outputs(2458) <= not((inputs(176)) or (inputs(204)));
    layer0_outputs(2459) <= (inputs(189)) xor (inputs(186));
    layer0_outputs(2460) <= (inputs(23)) and not (inputs(158));
    layer0_outputs(2461) <= inputs(142);
    layer0_outputs(2462) <= (inputs(112)) xor (inputs(25));
    layer0_outputs(2463) <= (inputs(199)) xor (inputs(186));
    layer0_outputs(2464) <= not((inputs(155)) and (inputs(56)));
    layer0_outputs(2465) <= (inputs(129)) or (inputs(6));
    layer0_outputs(2466) <= not(inputs(188));
    layer0_outputs(2467) <= '1';
    layer0_outputs(2468) <= (inputs(218)) and not (inputs(175));
    layer0_outputs(2469) <= inputs(113);
    layer0_outputs(2470) <= (inputs(255)) or (inputs(21));
    layer0_outputs(2471) <= not((inputs(212)) xor (inputs(219)));
    layer0_outputs(2472) <= not((inputs(227)) or (inputs(248)));
    layer0_outputs(2473) <= not(inputs(13));
    layer0_outputs(2474) <= (inputs(236)) or (inputs(148));
    layer0_outputs(2475) <= (inputs(162)) or (inputs(239));
    layer0_outputs(2476) <= not((inputs(1)) or (inputs(32)));
    layer0_outputs(2477) <= not((inputs(211)) or (inputs(71)));
    layer0_outputs(2478) <= (inputs(89)) and not (inputs(206));
    layer0_outputs(2479) <= inputs(45);
    layer0_outputs(2480) <= not(inputs(200));
    layer0_outputs(2481) <= inputs(55);
    layer0_outputs(2482) <= not(inputs(166)) or (inputs(85));
    layer0_outputs(2483) <= '0';
    layer0_outputs(2484) <= not(inputs(154)) or (inputs(28));
    layer0_outputs(2485) <= not((inputs(14)) or (inputs(252)));
    layer0_outputs(2486) <= (inputs(71)) xor (inputs(100));
    layer0_outputs(2487) <= inputs(56);
    layer0_outputs(2488) <= not(inputs(24));
    layer0_outputs(2489) <= not((inputs(130)) xor (inputs(117)));
    layer0_outputs(2490) <= (inputs(233)) and (inputs(198));
    layer0_outputs(2491) <= (inputs(80)) or (inputs(132));
    layer0_outputs(2492) <= not(inputs(202)) or (inputs(97));
    layer0_outputs(2493) <= (inputs(251)) or (inputs(5));
    layer0_outputs(2494) <= inputs(117);
    layer0_outputs(2495) <= not((inputs(234)) xor (inputs(169)));
    layer0_outputs(2496) <= not((inputs(214)) xor (inputs(244)));
    layer0_outputs(2497) <= not(inputs(173)) or (inputs(29));
    layer0_outputs(2498) <= not((inputs(209)) or (inputs(158)));
    layer0_outputs(2499) <= inputs(114);
    layer0_outputs(2500) <= not(inputs(12)) or (inputs(47));
    layer0_outputs(2501) <= (inputs(22)) and not (inputs(178));
    layer0_outputs(2502) <= not(inputs(42));
    layer0_outputs(2503) <= not(inputs(126));
    layer0_outputs(2504) <= not((inputs(63)) xor (inputs(86)));
    layer0_outputs(2505) <= (inputs(20)) and not (inputs(231));
    layer0_outputs(2506) <= (inputs(34)) or (inputs(188));
    layer0_outputs(2507) <= '0';
    layer0_outputs(2508) <= (inputs(242)) xor (inputs(80));
    layer0_outputs(2509) <= (inputs(27)) xor (inputs(49));
    layer0_outputs(2510) <= (inputs(47)) xor (inputs(126));
    layer0_outputs(2511) <= (inputs(124)) and (inputs(99));
    layer0_outputs(2512) <= inputs(186);
    layer0_outputs(2513) <= (inputs(40)) and (inputs(229));
    layer0_outputs(2514) <= (inputs(44)) xor (inputs(176));
    layer0_outputs(2515) <= '1';
    layer0_outputs(2516) <= inputs(232);
    layer0_outputs(2517) <= (inputs(44)) xor (inputs(71));
    layer0_outputs(2518) <= inputs(245);
    layer0_outputs(2519) <= (inputs(15)) and not (inputs(170));
    layer0_outputs(2520) <= inputs(194);
    layer0_outputs(2521) <= not((inputs(132)) or (inputs(78)));
    layer0_outputs(2522) <= inputs(56);
    layer0_outputs(2523) <= not((inputs(251)) or (inputs(97)));
    layer0_outputs(2524) <= inputs(125);
    layer0_outputs(2525) <= (inputs(23)) or (inputs(189));
    layer0_outputs(2526) <= (inputs(78)) and not (inputs(44));
    layer0_outputs(2527) <= inputs(62);
    layer0_outputs(2528) <= (inputs(106)) and not (inputs(227));
    layer0_outputs(2529) <= (inputs(142)) or (inputs(182));
    layer0_outputs(2530) <= (inputs(218)) xor (inputs(122));
    layer0_outputs(2531) <= (inputs(48)) and not (inputs(238));
    layer0_outputs(2532) <= not((inputs(30)) or (inputs(148)));
    layer0_outputs(2533) <= (inputs(117)) and not (inputs(124));
    layer0_outputs(2534) <= (inputs(0)) and not (inputs(32));
    layer0_outputs(2535) <= (inputs(116)) xor (inputs(111));
    layer0_outputs(2536) <= (inputs(188)) or (inputs(159));
    layer0_outputs(2537) <= (inputs(80)) or (inputs(211));
    layer0_outputs(2538) <= not(inputs(27));
    layer0_outputs(2539) <= inputs(69);
    layer0_outputs(2540) <= not(inputs(20)) or (inputs(199));
    layer0_outputs(2541) <= inputs(154);
    layer0_outputs(2542) <= (inputs(96)) or (inputs(92));
    layer0_outputs(2543) <= (inputs(119)) or (inputs(133));
    layer0_outputs(2544) <= (inputs(62)) xor (inputs(202));
    layer0_outputs(2545) <= not((inputs(55)) or (inputs(245)));
    layer0_outputs(2546) <= inputs(97);
    layer0_outputs(2547) <= (inputs(38)) or (inputs(122));
    layer0_outputs(2548) <= (inputs(10)) xor (inputs(247));
    layer0_outputs(2549) <= inputs(169);
    layer0_outputs(2550) <= (inputs(186)) and not (inputs(154));
    layer0_outputs(2551) <= not(inputs(217)) or (inputs(118));
    layer0_outputs(2552) <= not((inputs(49)) or (inputs(232)));
    layer0_outputs(2553) <= (inputs(192)) xor (inputs(179));
    layer0_outputs(2554) <= not((inputs(185)) or (inputs(77)));
    layer0_outputs(2555) <= inputs(43);
    layer0_outputs(2556) <= not((inputs(231)) or (inputs(79)));
    layer0_outputs(2557) <= not((inputs(87)) or (inputs(136)));
    layer0_outputs(2558) <= (inputs(151)) or (inputs(16));
    layer0_outputs(2559) <= not(inputs(180)) or (inputs(99));
    layer0_outputs(2560) <= inputs(44);
    layer0_outputs(2561) <= not(inputs(20));
    layer0_outputs(2562) <= not(inputs(0));
    layer0_outputs(2563) <= not(inputs(147)) or (inputs(19));
    layer0_outputs(2564) <= not((inputs(194)) or (inputs(51)));
    layer0_outputs(2565) <= not((inputs(115)) or (inputs(171)));
    layer0_outputs(2566) <= not((inputs(40)) and (inputs(120)));
    layer0_outputs(2567) <= inputs(90);
    layer0_outputs(2568) <= (inputs(33)) or (inputs(19));
    layer0_outputs(2569) <= (inputs(200)) xor (inputs(196));
    layer0_outputs(2570) <= (inputs(42)) xor (inputs(71));
    layer0_outputs(2571) <= (inputs(95)) or (inputs(9));
    layer0_outputs(2572) <= not(inputs(152));
    layer0_outputs(2573) <= (inputs(57)) and not (inputs(194));
    layer0_outputs(2574) <= not((inputs(161)) xor (inputs(210)));
    layer0_outputs(2575) <= not(inputs(104));
    layer0_outputs(2576) <= not(inputs(176));
    layer0_outputs(2577) <= inputs(23);
    layer0_outputs(2578) <= inputs(140);
    layer0_outputs(2579) <= inputs(56);
    layer0_outputs(2580) <= inputs(22);
    layer0_outputs(2581) <= inputs(66);
    layer0_outputs(2582) <= inputs(156);
    layer0_outputs(2583) <= not(inputs(107)) or (inputs(221));
    layer0_outputs(2584) <= inputs(227);
    layer0_outputs(2585) <= '1';
    layer0_outputs(2586) <= (inputs(24)) xor (inputs(182));
    layer0_outputs(2587) <= (inputs(152)) and not (inputs(241));
    layer0_outputs(2588) <= not((inputs(131)) or (inputs(109)));
    layer0_outputs(2589) <= not(inputs(232)) or (inputs(70));
    layer0_outputs(2590) <= (inputs(75)) and not (inputs(142));
    layer0_outputs(2591) <= (inputs(87)) xor (inputs(85));
    layer0_outputs(2592) <= not((inputs(147)) or (inputs(69)));
    layer0_outputs(2593) <= inputs(106);
    layer0_outputs(2594) <= not((inputs(46)) xor (inputs(109)));
    layer0_outputs(2595) <= not(inputs(88));
    layer0_outputs(2596) <= not(inputs(59));
    layer0_outputs(2597) <= not(inputs(117));
    layer0_outputs(2598) <= (inputs(136)) and (inputs(132));
    layer0_outputs(2599) <= not(inputs(210)) or (inputs(143));
    layer0_outputs(2600) <= not((inputs(81)) or (inputs(169)));
    layer0_outputs(2601) <= (inputs(231)) and not (inputs(239));
    layer0_outputs(2602) <= not(inputs(216));
    layer0_outputs(2603) <= not((inputs(139)) or (inputs(114)));
    layer0_outputs(2604) <= not(inputs(194)) or (inputs(242));
    layer0_outputs(2605) <= not(inputs(136));
    layer0_outputs(2606) <= (inputs(175)) xor (inputs(219));
    layer0_outputs(2607) <= (inputs(18)) xor (inputs(25));
    layer0_outputs(2608) <= not((inputs(164)) xor (inputs(120)));
    layer0_outputs(2609) <= not((inputs(140)) xor (inputs(123)));
    layer0_outputs(2610) <= (inputs(1)) xor (inputs(118));
    layer0_outputs(2611) <= not(inputs(249)) or (inputs(168));
    layer0_outputs(2612) <= (inputs(113)) and not (inputs(206));
    layer0_outputs(2613) <= not((inputs(123)) xor (inputs(53)));
    layer0_outputs(2614) <= not(inputs(49)) or (inputs(29));
    layer0_outputs(2615) <= not(inputs(59));
    layer0_outputs(2616) <= inputs(21);
    layer0_outputs(2617) <= inputs(12);
    layer0_outputs(2618) <= (inputs(190)) xor (inputs(239));
    layer0_outputs(2619) <= (inputs(217)) and not (inputs(46));
    layer0_outputs(2620) <= not(inputs(61)) or (inputs(172));
    layer0_outputs(2621) <= (inputs(88)) and not (inputs(220));
    layer0_outputs(2622) <= not(inputs(234));
    layer0_outputs(2623) <= (inputs(89)) and not (inputs(77));
    layer0_outputs(2624) <= not((inputs(252)) xor (inputs(32)));
    layer0_outputs(2625) <= inputs(179);
    layer0_outputs(2626) <= not((inputs(190)) or (inputs(183)));
    layer0_outputs(2627) <= not(inputs(149)) or (inputs(207));
    layer0_outputs(2628) <= not(inputs(182)) or (inputs(109));
    layer0_outputs(2629) <= inputs(111);
    layer0_outputs(2630) <= not((inputs(7)) or (inputs(155)));
    layer0_outputs(2631) <= inputs(17);
    layer0_outputs(2632) <= not((inputs(80)) and (inputs(240)));
    layer0_outputs(2633) <= (inputs(60)) and not (inputs(114));
    layer0_outputs(2634) <= not((inputs(60)) or (inputs(2)));
    layer0_outputs(2635) <= not(inputs(165)) or (inputs(169));
    layer0_outputs(2636) <= not(inputs(84));
    layer0_outputs(2637) <= (inputs(109)) xor (inputs(31));
    layer0_outputs(2638) <= (inputs(156)) xor (inputs(113));
    layer0_outputs(2639) <= (inputs(213)) and not (inputs(38));
    layer0_outputs(2640) <= not(inputs(123));
    layer0_outputs(2641) <= not(inputs(78));
    layer0_outputs(2642) <= (inputs(13)) xor (inputs(81));
    layer0_outputs(2643) <= not((inputs(136)) or (inputs(78)));
    layer0_outputs(2644) <= (inputs(225)) and not (inputs(152));
    layer0_outputs(2645) <= (inputs(107)) and (inputs(67));
    layer0_outputs(2646) <= inputs(15);
    layer0_outputs(2647) <= (inputs(59)) or (inputs(143));
    layer0_outputs(2648) <= not(inputs(55));
    layer0_outputs(2649) <= not((inputs(93)) and (inputs(93)));
    layer0_outputs(2650) <= not((inputs(223)) or (inputs(238)));
    layer0_outputs(2651) <= not((inputs(203)) xor (inputs(64)));
    layer0_outputs(2652) <= not(inputs(43)) or (inputs(114));
    layer0_outputs(2653) <= not((inputs(205)) or (inputs(13)));
    layer0_outputs(2654) <= (inputs(192)) or (inputs(16));
    layer0_outputs(2655) <= not((inputs(148)) xor (inputs(86)));
    layer0_outputs(2656) <= not(inputs(107)) or (inputs(245));
    layer0_outputs(2657) <= not((inputs(2)) or (inputs(93)));
    layer0_outputs(2658) <= (inputs(23)) and not (inputs(182));
    layer0_outputs(2659) <= not((inputs(37)) xor (inputs(16)));
    layer0_outputs(2660) <= (inputs(48)) xor (inputs(255));
    layer0_outputs(2661) <= not(inputs(8)) or (inputs(175));
    layer0_outputs(2662) <= (inputs(229)) and not (inputs(17));
    layer0_outputs(2663) <= not(inputs(8)) or (inputs(190));
    layer0_outputs(2664) <= not(inputs(209));
    layer0_outputs(2665) <= (inputs(150)) or (inputs(17));
    layer0_outputs(2666) <= (inputs(58)) or (inputs(14));
    layer0_outputs(2667) <= '1';
    layer0_outputs(2668) <= not(inputs(73));
    layer0_outputs(2669) <= not((inputs(207)) or (inputs(201)));
    layer0_outputs(2670) <= not(inputs(238)) or (inputs(129));
    layer0_outputs(2671) <= not(inputs(26));
    layer0_outputs(2672) <= (inputs(7)) or (inputs(120));
    layer0_outputs(2673) <= (inputs(195)) xor (inputs(237));
    layer0_outputs(2674) <= not(inputs(103)) or (inputs(159));
    layer0_outputs(2675) <= not((inputs(146)) xor (inputs(85)));
    layer0_outputs(2676) <= inputs(209);
    layer0_outputs(2677) <= not((inputs(128)) or (inputs(157)));
    layer0_outputs(2678) <= (inputs(180)) or (inputs(150));
    layer0_outputs(2679) <= inputs(59);
    layer0_outputs(2680) <= (inputs(31)) xor (inputs(60));
    layer0_outputs(2681) <= (inputs(157)) or (inputs(82));
    layer0_outputs(2682) <= not(inputs(220)) or (inputs(191));
    layer0_outputs(2683) <= (inputs(144)) and (inputs(112));
    layer0_outputs(2684) <= inputs(69);
    layer0_outputs(2685) <= not(inputs(22));
    layer0_outputs(2686) <= (inputs(249)) xor (inputs(46));
    layer0_outputs(2687) <= (inputs(61)) xor (inputs(169));
    layer0_outputs(2688) <= (inputs(116)) and not (inputs(191));
    layer0_outputs(2689) <= inputs(198);
    layer0_outputs(2690) <= (inputs(178)) xor (inputs(103));
    layer0_outputs(2691) <= not((inputs(191)) or (inputs(131)));
    layer0_outputs(2692) <= inputs(201);
    layer0_outputs(2693) <= not((inputs(240)) or (inputs(14)));
    layer0_outputs(2694) <= inputs(124);
    layer0_outputs(2695) <= not(inputs(86)) or (inputs(207));
    layer0_outputs(2696) <= not((inputs(136)) or (inputs(151)));
    layer0_outputs(2697) <= not(inputs(155)) or (inputs(16));
    layer0_outputs(2698) <= not(inputs(193));
    layer0_outputs(2699) <= (inputs(166)) and not (inputs(51));
    layer0_outputs(2700) <= not(inputs(195));
    layer0_outputs(2701) <= not(inputs(203)) or (inputs(124));
    layer0_outputs(2702) <= not((inputs(102)) xor (inputs(74)));
    layer0_outputs(2703) <= not(inputs(25)) or (inputs(186));
    layer0_outputs(2704) <= (inputs(208)) or (inputs(172));
    layer0_outputs(2705) <= not(inputs(28));
    layer0_outputs(2706) <= inputs(203);
    layer0_outputs(2707) <= (inputs(64)) and not (inputs(241));
    layer0_outputs(2708) <= not(inputs(142));
    layer0_outputs(2709) <= not((inputs(149)) xor (inputs(171)));
    layer0_outputs(2710) <= inputs(92);
    layer0_outputs(2711) <= (inputs(2)) or (inputs(21));
    layer0_outputs(2712) <= not((inputs(144)) or (inputs(38)));
    layer0_outputs(2713) <= not(inputs(0)) or (inputs(64));
    layer0_outputs(2714) <= not((inputs(242)) or (inputs(22)));
    layer0_outputs(2715) <= inputs(174);
    layer0_outputs(2716) <= (inputs(171)) and (inputs(154));
    layer0_outputs(2717) <= inputs(129);
    layer0_outputs(2718) <= (inputs(77)) and not (inputs(175));
    layer0_outputs(2719) <= not(inputs(36)) or (inputs(219));
    layer0_outputs(2720) <= inputs(231);
    layer0_outputs(2721) <= not(inputs(237));
    layer0_outputs(2722) <= not(inputs(25));
    layer0_outputs(2723) <= not(inputs(255)) or (inputs(42));
    layer0_outputs(2724) <= not(inputs(37)) or (inputs(239));
    layer0_outputs(2725) <= (inputs(23)) and not (inputs(194));
    layer0_outputs(2726) <= (inputs(161)) or (inputs(190));
    layer0_outputs(2727) <= (inputs(9)) and (inputs(87));
    layer0_outputs(2728) <= inputs(10);
    layer0_outputs(2729) <= (inputs(181)) xor (inputs(169));
    layer0_outputs(2730) <= not((inputs(180)) or (inputs(34)));
    layer0_outputs(2731) <= not((inputs(103)) or (inputs(60)));
    layer0_outputs(2732) <= (inputs(139)) xor (inputs(13));
    layer0_outputs(2733) <= not(inputs(210)) or (inputs(232));
    layer0_outputs(2734) <= (inputs(153)) and (inputs(146));
    layer0_outputs(2735) <= not((inputs(59)) or (inputs(3)));
    layer0_outputs(2736) <= not(inputs(153));
    layer0_outputs(2737) <= (inputs(71)) or (inputs(193));
    layer0_outputs(2738) <= not((inputs(200)) xor (inputs(240)));
    layer0_outputs(2739) <= (inputs(158)) and not (inputs(47));
    layer0_outputs(2740) <= not((inputs(35)) or (inputs(237)));
    layer0_outputs(2741) <= not(inputs(199));
    layer0_outputs(2742) <= not(inputs(235));
    layer0_outputs(2743) <= not((inputs(184)) xor (inputs(232)));
    layer0_outputs(2744) <= not(inputs(94)) or (inputs(63));
    layer0_outputs(2745) <= not((inputs(68)) or (inputs(164)));
    layer0_outputs(2746) <= (inputs(28)) or (inputs(16));
    layer0_outputs(2747) <= inputs(170);
    layer0_outputs(2748) <= not(inputs(117)) or (inputs(120));
    layer0_outputs(2749) <= not((inputs(86)) xor (inputs(145)));
    layer0_outputs(2750) <= not((inputs(84)) or (inputs(225)));
    layer0_outputs(2751) <= not(inputs(39));
    layer0_outputs(2752) <= inputs(252);
    layer0_outputs(2753) <= not(inputs(181));
    layer0_outputs(2754) <= not((inputs(168)) xor (inputs(149)));
    layer0_outputs(2755) <= (inputs(194)) and not (inputs(241));
    layer0_outputs(2756) <= (inputs(227)) xor (inputs(193));
    layer0_outputs(2757) <= (inputs(60)) and not (inputs(245));
    layer0_outputs(2758) <= not((inputs(179)) and (inputs(152)));
    layer0_outputs(2759) <= inputs(25);
    layer0_outputs(2760) <= not((inputs(14)) or (inputs(118)));
    layer0_outputs(2761) <= (inputs(210)) or (inputs(105));
    layer0_outputs(2762) <= not((inputs(193)) or (inputs(213)));
    layer0_outputs(2763) <= (inputs(80)) or (inputs(128));
    layer0_outputs(2764) <= not((inputs(44)) xor (inputs(49)));
    layer0_outputs(2765) <= not(inputs(73));
    layer0_outputs(2766) <= (inputs(65)) or (inputs(52));
    layer0_outputs(2767) <= not(inputs(184)) or (inputs(176));
    layer0_outputs(2768) <= not(inputs(125));
    layer0_outputs(2769) <= not(inputs(105)) or (inputs(86));
    layer0_outputs(2770) <= not(inputs(250));
    layer0_outputs(2771) <= not(inputs(192)) or (inputs(156));
    layer0_outputs(2772) <= not(inputs(251));
    layer0_outputs(2773) <= not(inputs(48)) or (inputs(2));
    layer0_outputs(2774) <= inputs(14);
    layer0_outputs(2775) <= (inputs(78)) and (inputs(126));
    layer0_outputs(2776) <= not(inputs(159)) or (inputs(171));
    layer0_outputs(2777) <= not(inputs(12));
    layer0_outputs(2778) <= not(inputs(163));
    layer0_outputs(2779) <= (inputs(109)) and not (inputs(252));
    layer0_outputs(2780) <= not(inputs(166));
    layer0_outputs(2781) <= inputs(35);
    layer0_outputs(2782) <= inputs(236);
    layer0_outputs(2783) <= (inputs(237)) xor (inputs(239));
    layer0_outputs(2784) <= not(inputs(91)) or (inputs(222));
    layer0_outputs(2785) <= inputs(70);
    layer0_outputs(2786) <= inputs(38);
    layer0_outputs(2787) <= not(inputs(244));
    layer0_outputs(2788) <= not(inputs(194)) or (inputs(252));
    layer0_outputs(2789) <= not(inputs(206));
    layer0_outputs(2790) <= not((inputs(246)) xor (inputs(178)));
    layer0_outputs(2791) <= not((inputs(228)) or (inputs(32)));
    layer0_outputs(2792) <= (inputs(91)) and not (inputs(160));
    layer0_outputs(2793) <= (inputs(255)) or (inputs(211));
    layer0_outputs(2794) <= inputs(177);
    layer0_outputs(2795) <= not(inputs(53)) or (inputs(174));
    layer0_outputs(2796) <= (inputs(5)) or (inputs(190));
    layer0_outputs(2797) <= (inputs(149)) and not (inputs(173));
    layer0_outputs(2798) <= inputs(218);
    layer0_outputs(2799) <= (inputs(188)) xor (inputs(20));
    layer0_outputs(2800) <= not(inputs(143));
    layer0_outputs(2801) <= (inputs(113)) xor (inputs(24));
    layer0_outputs(2802) <= (inputs(9)) xor (inputs(74));
    layer0_outputs(2803) <= (inputs(23)) xor (inputs(78));
    layer0_outputs(2804) <= inputs(201);
    layer0_outputs(2805) <= not((inputs(74)) xor (inputs(17)));
    layer0_outputs(2806) <= (inputs(90)) and not (inputs(210));
    layer0_outputs(2807) <= not((inputs(156)) xor (inputs(254)));
    layer0_outputs(2808) <= not(inputs(218)) or (inputs(0));
    layer0_outputs(2809) <= not((inputs(102)) xor (inputs(55)));
    layer0_outputs(2810) <= inputs(40);
    layer0_outputs(2811) <= inputs(248);
    layer0_outputs(2812) <= (inputs(239)) or (inputs(131));
    layer0_outputs(2813) <= inputs(220);
    layer0_outputs(2814) <= inputs(236);
    layer0_outputs(2815) <= (inputs(5)) and not (inputs(174));
    layer0_outputs(2816) <= not(inputs(47));
    layer0_outputs(2817) <= inputs(236);
    layer0_outputs(2818) <= not(inputs(24)) or (inputs(250));
    layer0_outputs(2819) <= not(inputs(119)) or (inputs(176));
    layer0_outputs(2820) <= not((inputs(162)) xor (inputs(208)));
    layer0_outputs(2821) <= inputs(93);
    layer0_outputs(2822) <= not(inputs(56));
    layer0_outputs(2823) <= not((inputs(253)) or (inputs(162)));
    layer0_outputs(2824) <= not((inputs(71)) xor (inputs(2)));
    layer0_outputs(2825) <= not(inputs(36));
    layer0_outputs(2826) <= not(inputs(108));
    layer0_outputs(2827) <= not((inputs(28)) xor (inputs(41)));
    layer0_outputs(2828) <= (inputs(246)) xor (inputs(225));
    layer0_outputs(2829) <= not(inputs(211)) or (inputs(110));
    layer0_outputs(2830) <= not(inputs(8));
    layer0_outputs(2831) <= inputs(135);
    layer0_outputs(2832) <= (inputs(214)) or (inputs(205));
    layer0_outputs(2833) <= not((inputs(177)) xor (inputs(131)));
    layer0_outputs(2834) <= not(inputs(9)) or (inputs(93));
    layer0_outputs(2835) <= inputs(231);
    layer0_outputs(2836) <= not(inputs(218));
    layer0_outputs(2837) <= (inputs(73)) xor (inputs(25));
    layer0_outputs(2838) <= (inputs(89)) and not (inputs(19));
    layer0_outputs(2839) <= inputs(123);
    layer0_outputs(2840) <= (inputs(3)) and not (inputs(30));
    layer0_outputs(2841) <= not(inputs(104));
    layer0_outputs(2842) <= (inputs(246)) xor (inputs(215));
    layer0_outputs(2843) <= (inputs(133)) and not (inputs(191));
    layer0_outputs(2844) <= not(inputs(213));
    layer0_outputs(2845) <= (inputs(22)) xor (inputs(222));
    layer0_outputs(2846) <= inputs(247);
    layer0_outputs(2847) <= (inputs(151)) and not (inputs(236));
    layer0_outputs(2848) <= (inputs(41)) and not (inputs(222));
    layer0_outputs(2849) <= (inputs(170)) and (inputs(251));
    layer0_outputs(2850) <= not(inputs(150));
    layer0_outputs(2851) <= (inputs(226)) and not (inputs(200));
    layer0_outputs(2852) <= not(inputs(23));
    layer0_outputs(2853) <= not((inputs(162)) or (inputs(175)));
    layer0_outputs(2854) <= not(inputs(32)) or (inputs(200));
    layer0_outputs(2855) <= not((inputs(253)) or (inputs(85)));
    layer0_outputs(2856) <= (inputs(132)) or (inputs(19));
    layer0_outputs(2857) <= not((inputs(222)) xor (inputs(77)));
    layer0_outputs(2858) <= (inputs(39)) xor (inputs(70));
    layer0_outputs(2859) <= (inputs(140)) or (inputs(222));
    layer0_outputs(2860) <= not(inputs(116)) or (inputs(44));
    layer0_outputs(2861) <= inputs(161);
    layer0_outputs(2862) <= not((inputs(214)) or (inputs(194)));
    layer0_outputs(2863) <= not((inputs(242)) and (inputs(219)));
    layer0_outputs(2864) <= (inputs(56)) xor (inputs(88));
    layer0_outputs(2865) <= (inputs(45)) and not (inputs(147));
    layer0_outputs(2866) <= '0';
    layer0_outputs(2867) <= (inputs(143)) or (inputs(162));
    layer0_outputs(2868) <= not(inputs(86));
    layer0_outputs(2869) <= inputs(218);
    layer0_outputs(2870) <= not(inputs(15));
    layer0_outputs(2871) <= (inputs(186)) xor (inputs(127));
    layer0_outputs(2872) <= (inputs(34)) or (inputs(25));
    layer0_outputs(2873) <= (inputs(88)) or (inputs(15));
    layer0_outputs(2874) <= not((inputs(0)) or (inputs(172)));
    layer0_outputs(2875) <= not((inputs(195)) xor (inputs(172)));
    layer0_outputs(2876) <= (inputs(70)) and not (inputs(139));
    layer0_outputs(2877) <= (inputs(187)) or (inputs(194));
    layer0_outputs(2878) <= not(inputs(42)) or (inputs(132));
    layer0_outputs(2879) <= not((inputs(150)) xor (inputs(53)));
    layer0_outputs(2880) <= inputs(182);
    layer0_outputs(2881) <= (inputs(181)) or (inputs(172));
    layer0_outputs(2882) <= not((inputs(249)) or (inputs(154)));
    layer0_outputs(2883) <= (inputs(158)) and not (inputs(46));
    layer0_outputs(2884) <= (inputs(160)) or (inputs(169));
    layer0_outputs(2885) <= (inputs(148)) and not (inputs(253));
    layer0_outputs(2886) <= not((inputs(107)) or (inputs(14)));
    layer0_outputs(2887) <= inputs(244);
    layer0_outputs(2888) <= not((inputs(232)) or (inputs(208)));
    layer0_outputs(2889) <= '0';
    layer0_outputs(2890) <= inputs(165);
    layer0_outputs(2891) <= (inputs(86)) xor (inputs(37));
    layer0_outputs(2892) <= not((inputs(73)) xor (inputs(247)));
    layer0_outputs(2893) <= (inputs(185)) or (inputs(160));
    layer0_outputs(2894) <= (inputs(139)) xor (inputs(172));
    layer0_outputs(2895) <= not((inputs(250)) and (inputs(16)));
    layer0_outputs(2896) <= (inputs(245)) and not (inputs(119));
    layer0_outputs(2897) <= (inputs(139)) or (inputs(123));
    layer0_outputs(2898) <= not(inputs(218));
    layer0_outputs(2899) <= not((inputs(219)) xor (inputs(224)));
    layer0_outputs(2900) <= not((inputs(39)) or (inputs(246)));
    layer0_outputs(2901) <= (inputs(115)) and not (inputs(19));
    layer0_outputs(2902) <= not(inputs(151)) or (inputs(63));
    layer0_outputs(2903) <= (inputs(63)) or (inputs(82));
    layer0_outputs(2904) <= not((inputs(246)) or (inputs(130)));
    layer0_outputs(2905) <= not((inputs(224)) or (inputs(253)));
    layer0_outputs(2906) <= inputs(166);
    layer0_outputs(2907) <= not((inputs(80)) xor (inputs(21)));
    layer0_outputs(2908) <= inputs(173);
    layer0_outputs(2909) <= not(inputs(235));
    layer0_outputs(2910) <= not((inputs(224)) or (inputs(5)));
    layer0_outputs(2911) <= not(inputs(179));
    layer0_outputs(2912) <= not(inputs(161)) or (inputs(255));
    layer0_outputs(2913) <= (inputs(194)) xor (inputs(94));
    layer0_outputs(2914) <= (inputs(224)) or (inputs(216));
    layer0_outputs(2915) <= (inputs(223)) or (inputs(205));
    layer0_outputs(2916) <= (inputs(89)) and not (inputs(216));
    layer0_outputs(2917) <= (inputs(239)) and (inputs(245));
    layer0_outputs(2918) <= (inputs(16)) and not (inputs(49));
    layer0_outputs(2919) <= not((inputs(6)) xor (inputs(156)));
    layer0_outputs(2920) <= not(inputs(24)) or (inputs(165));
    layer0_outputs(2921) <= (inputs(206)) or (inputs(242));
    layer0_outputs(2922) <= not(inputs(165));
    layer0_outputs(2923) <= (inputs(53)) or (inputs(212));
    layer0_outputs(2924) <= (inputs(9)) or (inputs(161));
    layer0_outputs(2925) <= (inputs(255)) and (inputs(254));
    layer0_outputs(2926) <= inputs(25);
    layer0_outputs(2927) <= inputs(152);
    layer0_outputs(2928) <= not(inputs(219));
    layer0_outputs(2929) <= not((inputs(25)) xor (inputs(234)));
    layer0_outputs(2930) <= (inputs(89)) and not (inputs(144));
    layer0_outputs(2931) <= inputs(152);
    layer0_outputs(2932) <= inputs(178);
    layer0_outputs(2933) <= not(inputs(216));
    layer0_outputs(2934) <= not((inputs(105)) or (inputs(167)));
    layer0_outputs(2935) <= (inputs(150)) xor (inputs(185));
    layer0_outputs(2936) <= '0';
    layer0_outputs(2937) <= inputs(115);
    layer0_outputs(2938) <= (inputs(46)) and not (inputs(253));
    layer0_outputs(2939) <= not((inputs(49)) or (inputs(150)));
    layer0_outputs(2940) <= not((inputs(73)) xor (inputs(45)));
    layer0_outputs(2941) <= inputs(155);
    layer0_outputs(2942) <= not((inputs(198)) or (inputs(94)));
    layer0_outputs(2943) <= not((inputs(3)) xor (inputs(223)));
    layer0_outputs(2944) <= not((inputs(30)) or (inputs(29)));
    layer0_outputs(2945) <= (inputs(247)) or (inputs(231));
    layer0_outputs(2946) <= inputs(218);
    layer0_outputs(2947) <= not(inputs(252)) or (inputs(214));
    layer0_outputs(2948) <= not((inputs(193)) xor (inputs(86)));
    layer0_outputs(2949) <= not((inputs(246)) xor (inputs(25)));
    layer0_outputs(2950) <= (inputs(51)) or (inputs(36));
    layer0_outputs(2951) <= inputs(72);
    layer0_outputs(2952) <= not((inputs(184)) and (inputs(253)));
    layer0_outputs(2953) <= (inputs(48)) or (inputs(176));
    layer0_outputs(2954) <= inputs(70);
    layer0_outputs(2955) <= inputs(247);
    layer0_outputs(2956) <= not((inputs(235)) xor (inputs(233)));
    layer0_outputs(2957) <= (inputs(157)) or (inputs(4));
    layer0_outputs(2958) <= not(inputs(120)) or (inputs(38));
    layer0_outputs(2959) <= (inputs(146)) or (inputs(112));
    layer0_outputs(2960) <= not((inputs(10)) xor (inputs(43)));
    layer0_outputs(2961) <= (inputs(184)) xor (inputs(88));
    layer0_outputs(2962) <= inputs(81);
    layer0_outputs(2963) <= not(inputs(171));
    layer0_outputs(2964) <= not((inputs(135)) xor (inputs(159)));
    layer0_outputs(2965) <= not(inputs(247));
    layer0_outputs(2966) <= not(inputs(29));
    layer0_outputs(2967) <= not(inputs(27));
    layer0_outputs(2968) <= inputs(92);
    layer0_outputs(2969) <= (inputs(212)) xor (inputs(250));
    layer0_outputs(2970) <= (inputs(7)) or (inputs(81));
    layer0_outputs(2971) <= not((inputs(202)) xor (inputs(89)));
    layer0_outputs(2972) <= (inputs(191)) and not (inputs(143));
    layer0_outputs(2973) <= inputs(243);
    layer0_outputs(2974) <= not((inputs(223)) xor (inputs(98)));
    layer0_outputs(2975) <= not(inputs(115)) or (inputs(205));
    layer0_outputs(2976) <= not((inputs(184)) xor (inputs(69)));
    layer0_outputs(2977) <= (inputs(64)) or (inputs(58));
    layer0_outputs(2978) <= (inputs(132)) and not (inputs(75));
    layer0_outputs(2979) <= inputs(226);
    layer0_outputs(2980) <= not((inputs(18)) xor (inputs(191)));
    layer0_outputs(2981) <= not((inputs(37)) or (inputs(32)));
    layer0_outputs(2982) <= (inputs(26)) xor (inputs(92));
    layer0_outputs(2983) <= not((inputs(115)) xor (inputs(117)));
    layer0_outputs(2984) <= not((inputs(135)) or (inputs(18)));
    layer0_outputs(2985) <= not((inputs(211)) or (inputs(232)));
    layer0_outputs(2986) <= inputs(196);
    layer0_outputs(2987) <= (inputs(151)) and not (inputs(162));
    layer0_outputs(2988) <= (inputs(43)) and not (inputs(255));
    layer0_outputs(2989) <= '1';
    layer0_outputs(2990) <= not(inputs(116));
    layer0_outputs(2991) <= (inputs(229)) or (inputs(233));
    layer0_outputs(2992) <= not((inputs(119)) xor (inputs(94)));
    layer0_outputs(2993) <= not((inputs(112)) xor (inputs(132)));
    layer0_outputs(2994) <= (inputs(8)) and not (inputs(126));
    layer0_outputs(2995) <= not(inputs(39)) or (inputs(87));
    layer0_outputs(2996) <= (inputs(34)) or (inputs(226));
    layer0_outputs(2997) <= not((inputs(61)) xor (inputs(16)));
    layer0_outputs(2998) <= not((inputs(237)) or (inputs(165)));
    layer0_outputs(2999) <= not((inputs(211)) or (inputs(53)));
    layer0_outputs(3000) <= (inputs(121)) and not (inputs(145));
    layer0_outputs(3001) <= not(inputs(189)) or (inputs(60));
    layer0_outputs(3002) <= not((inputs(96)) or (inputs(25)));
    layer0_outputs(3003) <= (inputs(110)) and (inputs(170));
    layer0_outputs(3004) <= (inputs(57)) or (inputs(61));
    layer0_outputs(3005) <= (inputs(78)) and (inputs(113));
    layer0_outputs(3006) <= not((inputs(94)) or (inputs(188)));
    layer0_outputs(3007) <= (inputs(161)) and not (inputs(240));
    layer0_outputs(3008) <= (inputs(102)) and not (inputs(225));
    layer0_outputs(3009) <= inputs(93);
    layer0_outputs(3010) <= inputs(109);
    layer0_outputs(3011) <= (inputs(220)) or (inputs(253));
    layer0_outputs(3012) <= not(inputs(22));
    layer0_outputs(3013) <= not((inputs(2)) xor (inputs(70)));
    layer0_outputs(3014) <= not(inputs(158));
    layer0_outputs(3015) <= not(inputs(174));
    layer0_outputs(3016) <= (inputs(160)) and not (inputs(0));
    layer0_outputs(3017) <= (inputs(202)) or (inputs(130));
    layer0_outputs(3018) <= (inputs(27)) xor (inputs(227));
    layer0_outputs(3019) <= inputs(168);
    layer0_outputs(3020) <= not(inputs(182));
    layer0_outputs(3021) <= inputs(194);
    layer0_outputs(3022) <= not(inputs(245));
    layer0_outputs(3023) <= (inputs(145)) xor (inputs(91));
    layer0_outputs(3024) <= (inputs(26)) and (inputs(9));
    layer0_outputs(3025) <= not((inputs(200)) or (inputs(169)));
    layer0_outputs(3026) <= not(inputs(80)) or (inputs(155));
    layer0_outputs(3027) <= not(inputs(154)) or (inputs(213));
    layer0_outputs(3028) <= (inputs(151)) or (inputs(236));
    layer0_outputs(3029) <= (inputs(81)) or (inputs(71));
    layer0_outputs(3030) <= not(inputs(58));
    layer0_outputs(3031) <= (inputs(203)) and not (inputs(69));
    layer0_outputs(3032) <= (inputs(101)) or (inputs(157));
    layer0_outputs(3033) <= not(inputs(201)) or (inputs(80));
    layer0_outputs(3034) <= (inputs(48)) or (inputs(20));
    layer0_outputs(3035) <= not((inputs(199)) or (inputs(67)));
    layer0_outputs(3036) <= (inputs(6)) and (inputs(7));
    layer0_outputs(3037) <= not((inputs(102)) xor (inputs(144)));
    layer0_outputs(3038) <= not((inputs(251)) xor (inputs(166)));
    layer0_outputs(3039) <= not((inputs(216)) xor (inputs(184)));
    layer0_outputs(3040) <= (inputs(244)) xor (inputs(16));
    layer0_outputs(3041) <= (inputs(190)) and not (inputs(214));
    layer0_outputs(3042) <= not((inputs(4)) or (inputs(216)));
    layer0_outputs(3043) <= inputs(239);
    layer0_outputs(3044) <= (inputs(153)) and not (inputs(21));
    layer0_outputs(3045) <= inputs(63);
    layer0_outputs(3046) <= not((inputs(235)) xor (inputs(220)));
    layer0_outputs(3047) <= inputs(54);
    layer0_outputs(3048) <= not(inputs(187));
    layer0_outputs(3049) <= (inputs(232)) and not (inputs(57));
    layer0_outputs(3050) <= not((inputs(250)) or (inputs(234)));
    layer0_outputs(3051) <= inputs(202);
    layer0_outputs(3052) <= (inputs(225)) xor (inputs(213));
    layer0_outputs(3053) <= not((inputs(172)) xor (inputs(61)));
    layer0_outputs(3054) <= not((inputs(245)) or (inputs(107)));
    layer0_outputs(3055) <= (inputs(202)) and not (inputs(154));
    layer0_outputs(3056) <= (inputs(122)) or (inputs(252));
    layer0_outputs(3057) <= inputs(238);
    layer0_outputs(3058) <= (inputs(33)) xor (inputs(0));
    layer0_outputs(3059) <= not(inputs(86)) or (inputs(1));
    layer0_outputs(3060) <= (inputs(195)) and (inputs(70));
    layer0_outputs(3061) <= (inputs(102)) and not (inputs(14));
    layer0_outputs(3062) <= not(inputs(218));
    layer0_outputs(3063) <= not((inputs(51)) xor (inputs(209)));
    layer0_outputs(3064) <= not(inputs(93)) or (inputs(198));
    layer0_outputs(3065) <= inputs(197);
    layer0_outputs(3066) <= inputs(160);
    layer0_outputs(3067) <= not(inputs(214)) or (inputs(56));
    layer0_outputs(3068) <= (inputs(187)) xor (inputs(195));
    layer0_outputs(3069) <= not((inputs(116)) or (inputs(253)));
    layer0_outputs(3070) <= inputs(39);
    layer0_outputs(3071) <= not((inputs(105)) or (inputs(137)));
    layer0_outputs(3072) <= inputs(129);
    layer0_outputs(3073) <= (inputs(51)) and not (inputs(0));
    layer0_outputs(3074) <= inputs(150);
    layer0_outputs(3075) <= not(inputs(105)) or (inputs(237));
    layer0_outputs(3076) <= not((inputs(213)) or (inputs(21)));
    layer0_outputs(3077) <= not((inputs(22)) and (inputs(87)));
    layer0_outputs(3078) <= not(inputs(97));
    layer0_outputs(3079) <= not((inputs(244)) xor (inputs(201)));
    layer0_outputs(3080) <= not((inputs(123)) or (inputs(138)));
    layer0_outputs(3081) <= not((inputs(140)) xor (inputs(203)));
    layer0_outputs(3082) <= (inputs(245)) and not (inputs(66));
    layer0_outputs(3083) <= not(inputs(74)) or (inputs(88));
    layer0_outputs(3084) <= (inputs(70)) xor (inputs(51));
    layer0_outputs(3085) <= (inputs(51)) xor (inputs(176));
    layer0_outputs(3086) <= inputs(28);
    layer0_outputs(3087) <= (inputs(101)) and not (inputs(16));
    layer0_outputs(3088) <= inputs(119);
    layer0_outputs(3089) <= (inputs(245)) and (inputs(217));
    layer0_outputs(3090) <= (inputs(105)) or (inputs(158));
    layer0_outputs(3091) <= (inputs(112)) and (inputs(149));
    layer0_outputs(3092) <= (inputs(199)) or (inputs(13));
    layer0_outputs(3093) <= inputs(67);
    layer0_outputs(3094) <= not(inputs(86));
    layer0_outputs(3095) <= not(inputs(169));
    layer0_outputs(3096) <= (inputs(222)) xor (inputs(24));
    layer0_outputs(3097) <= not(inputs(210));
    layer0_outputs(3098) <= not((inputs(209)) or (inputs(251)));
    layer0_outputs(3099) <= not((inputs(163)) xor (inputs(202)));
    layer0_outputs(3100) <= (inputs(212)) xor (inputs(118));
    layer0_outputs(3101) <= not(inputs(140)) or (inputs(15));
    layer0_outputs(3102) <= not(inputs(107)) or (inputs(245));
    layer0_outputs(3103) <= not(inputs(74));
    layer0_outputs(3104) <= not(inputs(129)) or (inputs(57));
    layer0_outputs(3105) <= not(inputs(185));
    layer0_outputs(3106) <= not(inputs(1));
    layer0_outputs(3107) <= not(inputs(149)) or (inputs(138));
    layer0_outputs(3108) <= not(inputs(88)) or (inputs(171));
    layer0_outputs(3109) <= not(inputs(64)) or (inputs(28));
    layer0_outputs(3110) <= (inputs(20)) xor (inputs(206));
    layer0_outputs(3111) <= (inputs(118)) and not (inputs(113));
    layer0_outputs(3112) <= not(inputs(149));
    layer0_outputs(3113) <= inputs(249);
    layer0_outputs(3114) <= not((inputs(251)) or (inputs(13)));
    layer0_outputs(3115) <= not(inputs(127));
    layer0_outputs(3116) <= (inputs(106)) xor (inputs(96));
    layer0_outputs(3117) <= (inputs(105)) xor (inputs(141));
    layer0_outputs(3118) <= not((inputs(233)) or (inputs(220)));
    layer0_outputs(3119) <= inputs(137);
    layer0_outputs(3120) <= (inputs(16)) xor (inputs(123));
    layer0_outputs(3121) <= (inputs(119)) and not (inputs(254));
    layer0_outputs(3122) <= not(inputs(37)) or (inputs(234));
    layer0_outputs(3123) <= not(inputs(145));
    layer0_outputs(3124) <= (inputs(154)) xor (inputs(18));
    layer0_outputs(3125) <= (inputs(8)) or (inputs(247));
    layer0_outputs(3126) <= not((inputs(217)) xor (inputs(23)));
    layer0_outputs(3127) <= not(inputs(27));
    layer0_outputs(3128) <= not(inputs(218)) or (inputs(127));
    layer0_outputs(3129) <= not(inputs(219)) or (inputs(80));
    layer0_outputs(3130) <= not(inputs(77));
    layer0_outputs(3131) <= (inputs(55)) or (inputs(31));
    layer0_outputs(3132) <= inputs(180);
    layer0_outputs(3133) <= inputs(135);
    layer0_outputs(3134) <= not(inputs(88));
    layer0_outputs(3135) <= (inputs(79)) or (inputs(68));
    layer0_outputs(3136) <= not((inputs(116)) xor (inputs(43)));
    layer0_outputs(3137) <= not((inputs(180)) xor (inputs(241)));
    layer0_outputs(3138) <= (inputs(8)) and not (inputs(45));
    layer0_outputs(3139) <= (inputs(222)) or (inputs(188));
    layer0_outputs(3140) <= not(inputs(221));
    layer0_outputs(3141) <= not(inputs(102));
    layer0_outputs(3142) <= (inputs(26)) xor (inputs(215));
    layer0_outputs(3143) <= inputs(197);
    layer0_outputs(3144) <= (inputs(21)) and (inputs(24));
    layer0_outputs(3145) <= not(inputs(24));
    layer0_outputs(3146) <= (inputs(26)) xor (inputs(189));
    layer0_outputs(3147) <= inputs(44);
    layer0_outputs(3148) <= not(inputs(183));
    layer0_outputs(3149) <= (inputs(18)) or (inputs(192));
    layer0_outputs(3150) <= not(inputs(247)) or (inputs(73));
    layer0_outputs(3151) <= inputs(242);
    layer0_outputs(3152) <= not((inputs(193)) xor (inputs(217)));
    layer0_outputs(3153) <= not(inputs(21));
    layer0_outputs(3154) <= not(inputs(137));
    layer0_outputs(3155) <= not((inputs(171)) xor (inputs(206)));
    layer0_outputs(3156) <= inputs(251);
    layer0_outputs(3157) <= not(inputs(36));
    layer0_outputs(3158) <= not((inputs(9)) or (inputs(66)));
    layer0_outputs(3159) <= (inputs(54)) and not (inputs(206));
    layer0_outputs(3160) <= not((inputs(15)) or (inputs(106)));
    layer0_outputs(3161) <= not(inputs(89)) or (inputs(128));
    layer0_outputs(3162) <= not(inputs(108));
    layer0_outputs(3163) <= (inputs(238)) or (inputs(239));
    layer0_outputs(3164) <= not((inputs(12)) xor (inputs(29)));
    layer0_outputs(3165) <= inputs(96);
    layer0_outputs(3166) <= not(inputs(52)) or (inputs(93));
    layer0_outputs(3167) <= not(inputs(56)) or (inputs(237));
    layer0_outputs(3168) <= (inputs(7)) xor (inputs(83));
    layer0_outputs(3169) <= not(inputs(162));
    layer0_outputs(3170) <= not((inputs(243)) xor (inputs(64)));
    layer0_outputs(3171) <= (inputs(166)) or (inputs(3));
    layer0_outputs(3172) <= inputs(200);
    layer0_outputs(3173) <= not((inputs(184)) xor (inputs(11)));
    layer0_outputs(3174) <= (inputs(218)) or (inputs(67));
    layer0_outputs(3175) <= not(inputs(230));
    layer0_outputs(3176) <= inputs(57);
    layer0_outputs(3177) <= inputs(39);
    layer0_outputs(3178) <= not(inputs(229));
    layer0_outputs(3179) <= not((inputs(182)) xor (inputs(218)));
    layer0_outputs(3180) <= (inputs(231)) xor (inputs(176));
    layer0_outputs(3181) <= not((inputs(47)) or (inputs(156)));
    layer0_outputs(3182) <= not((inputs(121)) xor (inputs(162)));
    layer0_outputs(3183) <= (inputs(166)) xor (inputs(104));
    layer0_outputs(3184) <= not(inputs(187)) or (inputs(120));
    layer0_outputs(3185) <= not(inputs(115));
    layer0_outputs(3186) <= not((inputs(154)) xor (inputs(225)));
    layer0_outputs(3187) <= inputs(230);
    layer0_outputs(3188) <= (inputs(206)) xor (inputs(141));
    layer0_outputs(3189) <= (inputs(191)) or (inputs(137));
    layer0_outputs(3190) <= (inputs(132)) and not (inputs(16));
    layer0_outputs(3191) <= not(inputs(26)) or (inputs(250));
    layer0_outputs(3192) <= not(inputs(212));
    layer0_outputs(3193) <= (inputs(244)) and not (inputs(80));
    layer0_outputs(3194) <= inputs(128);
    layer0_outputs(3195) <= (inputs(11)) xor (inputs(60));
    layer0_outputs(3196) <= inputs(132);
    layer0_outputs(3197) <= (inputs(220)) xor (inputs(244));
    layer0_outputs(3198) <= not(inputs(74));
    layer0_outputs(3199) <= (inputs(187)) and not (inputs(56));
    layer0_outputs(3200) <= not(inputs(235));
    layer0_outputs(3201) <= not((inputs(45)) or (inputs(202)));
    layer0_outputs(3202) <= not(inputs(178)) or (inputs(17));
    layer0_outputs(3203) <= (inputs(24)) and not (inputs(103));
    layer0_outputs(3204) <= not(inputs(115)) or (inputs(206));
    layer0_outputs(3205) <= (inputs(102)) xor (inputs(72));
    layer0_outputs(3206) <= (inputs(17)) or (inputs(142));
    layer0_outputs(3207) <= not((inputs(96)) xor (inputs(246)));
    layer0_outputs(3208) <= inputs(58);
    layer0_outputs(3209) <= (inputs(126)) or (inputs(135));
    layer0_outputs(3210) <= (inputs(121)) or (inputs(236));
    layer0_outputs(3211) <= (inputs(178)) or (inputs(147));
    layer0_outputs(3212) <= not(inputs(133)) or (inputs(242));
    layer0_outputs(3213) <= (inputs(106)) or (inputs(61));
    layer0_outputs(3214) <= (inputs(146)) or (inputs(187));
    layer0_outputs(3215) <= not(inputs(118));
    layer0_outputs(3216) <= not(inputs(209));
    layer0_outputs(3217) <= (inputs(50)) xor (inputs(183));
    layer0_outputs(3218) <= (inputs(253)) or (inputs(199));
    layer0_outputs(3219) <= (inputs(142)) and not (inputs(14));
    layer0_outputs(3220) <= not(inputs(142));
    layer0_outputs(3221) <= not(inputs(234)) or (inputs(31));
    layer0_outputs(3222) <= not(inputs(179)) or (inputs(47));
    layer0_outputs(3223) <= not((inputs(72)) or (inputs(218)));
    layer0_outputs(3224) <= (inputs(157)) or (inputs(191));
    layer0_outputs(3225) <= (inputs(212)) and not (inputs(149));
    layer0_outputs(3226) <= (inputs(240)) or (inputs(111));
    layer0_outputs(3227) <= (inputs(234)) and not (inputs(47));
    layer0_outputs(3228) <= (inputs(199)) and not (inputs(218));
    layer0_outputs(3229) <= (inputs(93)) or (inputs(192));
    layer0_outputs(3230) <= not((inputs(58)) or (inputs(118)));
    layer0_outputs(3231) <= '0';
    layer0_outputs(3232) <= not(inputs(252));
    layer0_outputs(3233) <= inputs(3);
    layer0_outputs(3234) <= not((inputs(185)) xor (inputs(7)));
    layer0_outputs(3235) <= not(inputs(102));
    layer0_outputs(3236) <= not(inputs(36));
    layer0_outputs(3237) <= not((inputs(194)) or (inputs(111)));
    layer0_outputs(3238) <= (inputs(110)) or (inputs(79));
    layer0_outputs(3239) <= not((inputs(140)) xor (inputs(228)));
    layer0_outputs(3240) <= not(inputs(48));
    layer0_outputs(3241) <= (inputs(199)) and not (inputs(140));
    layer0_outputs(3242) <= (inputs(251)) and not (inputs(98));
    layer0_outputs(3243) <= not(inputs(181));
    layer0_outputs(3244) <= (inputs(204)) xor (inputs(138));
    layer0_outputs(3245) <= (inputs(162)) xor (inputs(212));
    layer0_outputs(3246) <= (inputs(202)) xor (inputs(15));
    layer0_outputs(3247) <= (inputs(154)) and not (inputs(229));
    layer0_outputs(3248) <= not(inputs(243)) or (inputs(158));
    layer0_outputs(3249) <= (inputs(74)) or (inputs(108));
    layer0_outputs(3250) <= (inputs(90)) xor (inputs(108));
    layer0_outputs(3251) <= not((inputs(16)) xor (inputs(65)));
    layer0_outputs(3252) <= not((inputs(130)) or (inputs(197)));
    layer0_outputs(3253) <= not(inputs(163));
    layer0_outputs(3254) <= inputs(6);
    layer0_outputs(3255) <= (inputs(194)) and not (inputs(15));
    layer0_outputs(3256) <= not(inputs(185)) or (inputs(106));
    layer0_outputs(3257) <= not((inputs(53)) xor (inputs(232)));
    layer0_outputs(3258) <= not(inputs(132)) or (inputs(49));
    layer0_outputs(3259) <= (inputs(132)) or (inputs(181));
    layer0_outputs(3260) <= not((inputs(193)) or (inputs(26)));
    layer0_outputs(3261) <= not((inputs(103)) xor (inputs(57)));
    layer0_outputs(3262) <= (inputs(233)) xor (inputs(67));
    layer0_outputs(3263) <= not((inputs(255)) or (inputs(26)));
    layer0_outputs(3264) <= not(inputs(7)) or (inputs(124));
    layer0_outputs(3265) <= inputs(177);
    layer0_outputs(3266) <= (inputs(196)) and (inputs(221));
    layer0_outputs(3267) <= (inputs(108)) and (inputs(156));
    layer0_outputs(3268) <= not(inputs(164));
    layer0_outputs(3269) <= not(inputs(59));
    layer0_outputs(3270) <= not(inputs(224)) or (inputs(241));
    layer0_outputs(3271) <= not(inputs(84)) or (inputs(110));
    layer0_outputs(3272) <= not((inputs(224)) xor (inputs(91)));
    layer0_outputs(3273) <= not(inputs(157));
    layer0_outputs(3274) <= not((inputs(173)) xor (inputs(171)));
    layer0_outputs(3275) <= not(inputs(22)) or (inputs(98));
    layer0_outputs(3276) <= not(inputs(252));
    layer0_outputs(3277) <= not(inputs(140));
    layer0_outputs(3278) <= inputs(114);
    layer0_outputs(3279) <= not(inputs(162));
    layer0_outputs(3280) <= not(inputs(114)) or (inputs(49));
    layer0_outputs(3281) <= inputs(20);
    layer0_outputs(3282) <= (inputs(160)) and not (inputs(9));
    layer0_outputs(3283) <= not(inputs(233)) or (inputs(5));
    layer0_outputs(3284) <= not(inputs(161)) or (inputs(218));
    layer0_outputs(3285) <= '1';
    layer0_outputs(3286) <= not(inputs(43)) or (inputs(97));
    layer0_outputs(3287) <= (inputs(183)) and not (inputs(124));
    layer0_outputs(3288) <= not(inputs(2)) or (inputs(238));
    layer0_outputs(3289) <= not((inputs(10)) xor (inputs(18)));
    layer0_outputs(3290) <= (inputs(140)) xor (inputs(27));
    layer0_outputs(3291) <= not(inputs(105)) or (inputs(210));
    layer0_outputs(3292) <= (inputs(35)) xor (inputs(205));
    layer0_outputs(3293) <= (inputs(59)) or (inputs(104));
    layer0_outputs(3294) <= (inputs(170)) and (inputs(212));
    layer0_outputs(3295) <= not((inputs(27)) or (inputs(248)));
    layer0_outputs(3296) <= (inputs(137)) and not (inputs(181));
    layer0_outputs(3297) <= not(inputs(162));
    layer0_outputs(3298) <= not(inputs(8)) or (inputs(242));
    layer0_outputs(3299) <= (inputs(238)) or (inputs(110));
    layer0_outputs(3300) <= not(inputs(97)) or (inputs(142));
    layer0_outputs(3301) <= (inputs(52)) and not (inputs(128));
    layer0_outputs(3302) <= not((inputs(145)) and (inputs(242)));
    layer0_outputs(3303) <= not(inputs(196)) or (inputs(5));
    layer0_outputs(3304) <= (inputs(101)) xor (inputs(25));
    layer0_outputs(3305) <= not(inputs(221)) or (inputs(19));
    layer0_outputs(3306) <= not(inputs(8)) or (inputs(243));
    layer0_outputs(3307) <= not((inputs(246)) xor (inputs(213)));
    layer0_outputs(3308) <= not((inputs(233)) and (inputs(221)));
    layer0_outputs(3309) <= not((inputs(49)) xor (inputs(71)));
    layer0_outputs(3310) <= not(inputs(229)) or (inputs(114));
    layer0_outputs(3311) <= inputs(59);
    layer0_outputs(3312) <= not(inputs(230));
    layer0_outputs(3313) <= not((inputs(25)) xor (inputs(72)));
    layer0_outputs(3314) <= (inputs(204)) or (inputs(141));
    layer0_outputs(3315) <= not((inputs(250)) or (inputs(230)));
    layer0_outputs(3316) <= not(inputs(57));
    layer0_outputs(3317) <= not((inputs(196)) xor (inputs(244)));
    layer0_outputs(3318) <= (inputs(202)) and not (inputs(159));
    layer0_outputs(3319) <= (inputs(4)) and not (inputs(95));
    layer0_outputs(3320) <= not((inputs(238)) or (inputs(118)));
    layer0_outputs(3321) <= not(inputs(182));
    layer0_outputs(3322) <= not((inputs(227)) xor (inputs(205)));
    layer0_outputs(3323) <= (inputs(90)) and not (inputs(173));
    layer0_outputs(3324) <= (inputs(134)) or (inputs(249));
    layer0_outputs(3325) <= inputs(114);
    layer0_outputs(3326) <= not((inputs(150)) xor (inputs(236)));
    layer0_outputs(3327) <= not((inputs(157)) xor (inputs(106)));
    layer0_outputs(3328) <= not((inputs(232)) or (inputs(243)));
    layer0_outputs(3329) <= (inputs(157)) and not (inputs(65));
    layer0_outputs(3330) <= inputs(224);
    layer0_outputs(3331) <= not((inputs(174)) or (inputs(23)));
    layer0_outputs(3332) <= not((inputs(137)) or (inputs(58)));
    layer0_outputs(3333) <= not(inputs(103));
    layer0_outputs(3334) <= inputs(61);
    layer0_outputs(3335) <= not((inputs(99)) or (inputs(218)));
    layer0_outputs(3336) <= inputs(66);
    layer0_outputs(3337) <= inputs(32);
    layer0_outputs(3338) <= not((inputs(247)) or (inputs(138)));
    layer0_outputs(3339) <= not(inputs(38)) or (inputs(14));
    layer0_outputs(3340) <= not(inputs(139)) or (inputs(254));
    layer0_outputs(3341) <= (inputs(242)) and (inputs(72));
    layer0_outputs(3342) <= not((inputs(113)) or (inputs(15)));
    layer0_outputs(3343) <= (inputs(74)) and not (inputs(71));
    layer0_outputs(3344) <= (inputs(219)) and not (inputs(237));
    layer0_outputs(3345) <= not(inputs(136)) or (inputs(79));
    layer0_outputs(3346) <= not((inputs(253)) and (inputs(86)));
    layer0_outputs(3347) <= not(inputs(205));
    layer0_outputs(3348) <= (inputs(25)) and (inputs(34));
    layer0_outputs(3349) <= (inputs(5)) xor (inputs(202));
    layer0_outputs(3350) <= (inputs(90)) or (inputs(120));
    layer0_outputs(3351) <= not(inputs(230)) or (inputs(41));
    layer0_outputs(3352) <= (inputs(73)) and not (inputs(202));
    layer0_outputs(3353) <= (inputs(26)) xor (inputs(235));
    layer0_outputs(3354) <= not((inputs(179)) xor (inputs(20)));
    layer0_outputs(3355) <= (inputs(63)) and not (inputs(255));
    layer0_outputs(3356) <= not(inputs(165));
    layer0_outputs(3357) <= not(inputs(246));
    layer0_outputs(3358) <= not(inputs(113));
    layer0_outputs(3359) <= not(inputs(114));
    layer0_outputs(3360) <= (inputs(51)) and not (inputs(174));
    layer0_outputs(3361) <= (inputs(221)) or (inputs(146));
    layer0_outputs(3362) <= not((inputs(214)) and (inputs(124)));
    layer0_outputs(3363) <= inputs(247);
    layer0_outputs(3364) <= (inputs(93)) or (inputs(114));
    layer0_outputs(3365) <= not((inputs(138)) and (inputs(173)));
    layer0_outputs(3366) <= not((inputs(167)) xor (inputs(6)));
    layer0_outputs(3367) <= not((inputs(220)) or (inputs(178)));
    layer0_outputs(3368) <= (inputs(96)) and (inputs(5));
    layer0_outputs(3369) <= not((inputs(18)) or (inputs(52)));
    layer0_outputs(3370) <= inputs(41);
    layer0_outputs(3371) <= (inputs(58)) and not (inputs(102));
    layer0_outputs(3372) <= (inputs(60)) xor (inputs(151));
    layer0_outputs(3373) <= (inputs(74)) or (inputs(34));
    layer0_outputs(3374) <= not((inputs(76)) xor (inputs(75)));
    layer0_outputs(3375) <= (inputs(137)) and not (inputs(164));
    layer0_outputs(3376) <= not(inputs(114));
    layer0_outputs(3377) <= not(inputs(43));
    layer0_outputs(3378) <= (inputs(218)) xor (inputs(121));
    layer0_outputs(3379) <= not((inputs(52)) or (inputs(46)));
    layer0_outputs(3380) <= (inputs(187)) and (inputs(238));
    layer0_outputs(3381) <= '1';
    layer0_outputs(3382) <= inputs(1);
    layer0_outputs(3383) <= (inputs(246)) and not (inputs(141));
    layer0_outputs(3384) <= (inputs(192)) xor (inputs(247));
    layer0_outputs(3385) <= not(inputs(183)) or (inputs(249));
    layer0_outputs(3386) <= (inputs(242)) xor (inputs(153));
    layer0_outputs(3387) <= not((inputs(157)) or (inputs(208)));
    layer0_outputs(3388) <= not((inputs(122)) or (inputs(191)));
    layer0_outputs(3389) <= inputs(230);
    layer0_outputs(3390) <= inputs(234);
    layer0_outputs(3391) <= (inputs(89)) xor (inputs(187));
    layer0_outputs(3392) <= not((inputs(189)) or (inputs(155)));
    layer0_outputs(3393) <= not(inputs(251)) or (inputs(61));
    layer0_outputs(3394) <= (inputs(22)) and not (inputs(163));
    layer0_outputs(3395) <= not(inputs(99));
    layer0_outputs(3396) <= not((inputs(78)) xor (inputs(7)));
    layer0_outputs(3397) <= not(inputs(204));
    layer0_outputs(3398) <= not(inputs(182)) or (inputs(136));
    layer0_outputs(3399) <= (inputs(191)) or (inputs(111));
    layer0_outputs(3400) <= not(inputs(67));
    layer0_outputs(3401) <= (inputs(16)) or (inputs(76));
    layer0_outputs(3402) <= (inputs(125)) xor (inputs(44));
    layer0_outputs(3403) <= not(inputs(201));
    layer0_outputs(3404) <= (inputs(193)) xor (inputs(241));
    layer0_outputs(3405) <= not(inputs(107));
    layer0_outputs(3406) <= not((inputs(123)) or (inputs(11)));
    layer0_outputs(3407) <= (inputs(207)) xor (inputs(206));
    layer0_outputs(3408) <= not(inputs(86)) or (inputs(141));
    layer0_outputs(3409) <= not(inputs(116)) or (inputs(57));
    layer0_outputs(3410) <= not((inputs(132)) and (inputs(83)));
    layer0_outputs(3411) <= (inputs(255)) or (inputs(198));
    layer0_outputs(3412) <= (inputs(129)) xor (inputs(163));
    layer0_outputs(3413) <= not((inputs(149)) and (inputs(199)));
    layer0_outputs(3414) <= (inputs(166)) and not (inputs(128));
    layer0_outputs(3415) <= not((inputs(132)) and (inputs(75)));
    layer0_outputs(3416) <= inputs(251);
    layer0_outputs(3417) <= not(inputs(54));
    layer0_outputs(3418) <= not(inputs(179)) or (inputs(240));
    layer0_outputs(3419) <= not(inputs(180));
    layer0_outputs(3420) <= inputs(135);
    layer0_outputs(3421) <= inputs(23);
    layer0_outputs(3422) <= not((inputs(161)) xor (inputs(177)));
    layer0_outputs(3423) <= (inputs(204)) xor (inputs(214));
    layer0_outputs(3424) <= inputs(252);
    layer0_outputs(3425) <= not(inputs(233));
    layer0_outputs(3426) <= (inputs(195)) and not (inputs(63));
    layer0_outputs(3427) <= (inputs(116)) or (inputs(52));
    layer0_outputs(3428) <= not((inputs(62)) or (inputs(254)));
    layer0_outputs(3429) <= (inputs(6)) and (inputs(200));
    layer0_outputs(3430) <= not(inputs(85));
    layer0_outputs(3431) <= not((inputs(153)) and (inputs(152)));
    layer0_outputs(3432) <= inputs(98);
    layer0_outputs(3433) <= not((inputs(172)) xor (inputs(109)));
    layer0_outputs(3434) <= not((inputs(164)) or (inputs(42)));
    layer0_outputs(3435) <= inputs(216);
    layer0_outputs(3436) <= not(inputs(227));
    layer0_outputs(3437) <= not(inputs(21)) or (inputs(144));
    layer0_outputs(3438) <= (inputs(96)) or (inputs(133));
    layer0_outputs(3439) <= inputs(74);
    layer0_outputs(3440) <= not(inputs(129));
    layer0_outputs(3441) <= (inputs(122)) or (inputs(239));
    layer0_outputs(3442) <= not((inputs(71)) or (inputs(35)));
    layer0_outputs(3443) <= not(inputs(179));
    layer0_outputs(3444) <= (inputs(121)) and not (inputs(172));
    layer0_outputs(3445) <= not((inputs(155)) or (inputs(186)));
    layer0_outputs(3446) <= (inputs(232)) xor (inputs(195));
    layer0_outputs(3447) <= (inputs(29)) and not (inputs(178));
    layer0_outputs(3448) <= not(inputs(133));
    layer0_outputs(3449) <= (inputs(188)) and not (inputs(108));
    layer0_outputs(3450) <= inputs(148);
    layer0_outputs(3451) <= inputs(131);
    layer0_outputs(3452) <= inputs(27);
    layer0_outputs(3453) <= not((inputs(108)) and (inputs(34)));
    layer0_outputs(3454) <= inputs(59);
    layer0_outputs(3455) <= (inputs(131)) and not (inputs(94));
    layer0_outputs(3456) <= (inputs(156)) or (inputs(98));
    layer0_outputs(3457) <= not((inputs(109)) and (inputs(146)));
    layer0_outputs(3458) <= (inputs(203)) or (inputs(103));
    layer0_outputs(3459) <= '1';
    layer0_outputs(3460) <= not(inputs(67));
    layer0_outputs(3461) <= not((inputs(84)) xor (inputs(54)));
    layer0_outputs(3462) <= not((inputs(166)) xor (inputs(143)));
    layer0_outputs(3463) <= not(inputs(193));
    layer0_outputs(3464) <= inputs(218);
    layer0_outputs(3465) <= (inputs(96)) and not (inputs(92));
    layer0_outputs(3466) <= inputs(168);
    layer0_outputs(3467) <= (inputs(145)) xor (inputs(223));
    layer0_outputs(3468) <= not(inputs(228)) or (inputs(187));
    layer0_outputs(3469) <= not(inputs(9));
    layer0_outputs(3470) <= inputs(78);
    layer0_outputs(3471) <= inputs(162);
    layer0_outputs(3472) <= not(inputs(39)) or (inputs(241));
    layer0_outputs(3473) <= inputs(225);
    layer0_outputs(3474) <= (inputs(234)) and not (inputs(58));
    layer0_outputs(3475) <= not(inputs(114));
    layer0_outputs(3476) <= (inputs(240)) or (inputs(19));
    layer0_outputs(3477) <= not((inputs(46)) xor (inputs(218)));
    layer0_outputs(3478) <= not((inputs(170)) or (inputs(176)));
    layer0_outputs(3479) <= (inputs(39)) xor (inputs(178));
    layer0_outputs(3480) <= not(inputs(146));
    layer0_outputs(3481) <= not((inputs(84)) and (inputs(106)));
    layer0_outputs(3482) <= not(inputs(141));
    layer0_outputs(3483) <= not(inputs(103));
    layer0_outputs(3484) <= not(inputs(121));
    layer0_outputs(3485) <= (inputs(50)) and not (inputs(149));
    layer0_outputs(3486) <= (inputs(228)) or (inputs(48));
    layer0_outputs(3487) <= (inputs(49)) or (inputs(5));
    layer0_outputs(3488) <= not((inputs(205)) xor (inputs(116)));
    layer0_outputs(3489) <= (inputs(93)) or (inputs(164));
    layer0_outputs(3490) <= not((inputs(231)) xor (inputs(249)));
    layer0_outputs(3491) <= inputs(224);
    layer0_outputs(3492) <= inputs(17);
    layer0_outputs(3493) <= (inputs(44)) xor (inputs(74));
    layer0_outputs(3494) <= not((inputs(85)) xor (inputs(1)));
    layer0_outputs(3495) <= not(inputs(215)) or (inputs(255));
    layer0_outputs(3496) <= not((inputs(206)) xor (inputs(132)));
    layer0_outputs(3497) <= not(inputs(7));
    layer0_outputs(3498) <= not(inputs(160));
    layer0_outputs(3499) <= not(inputs(107)) or (inputs(49));
    layer0_outputs(3500) <= not((inputs(98)) and (inputs(159)));
    layer0_outputs(3501) <= (inputs(15)) and not (inputs(191));
    layer0_outputs(3502) <= (inputs(243)) and not (inputs(28));
    layer0_outputs(3503) <= (inputs(193)) xor (inputs(80));
    layer0_outputs(3504) <= (inputs(98)) and not (inputs(72));
    layer0_outputs(3505) <= not((inputs(0)) xor (inputs(171)));
    layer0_outputs(3506) <= not(inputs(118));
    layer0_outputs(3507) <= not(inputs(98)) or (inputs(184));
    layer0_outputs(3508) <= not(inputs(158)) or (inputs(63));
    layer0_outputs(3509) <= inputs(222);
    layer0_outputs(3510) <= not((inputs(123)) or (inputs(121)));
    layer0_outputs(3511) <= not(inputs(100)) or (inputs(1));
    layer0_outputs(3512) <= (inputs(207)) xor (inputs(134));
    layer0_outputs(3513) <= not(inputs(203)) or (inputs(161));
    layer0_outputs(3514) <= not((inputs(77)) xor (inputs(100)));
    layer0_outputs(3515) <= inputs(102);
    layer0_outputs(3516) <= (inputs(161)) xor (inputs(68));
    layer0_outputs(3517) <= not((inputs(56)) xor (inputs(120)));
    layer0_outputs(3518) <= (inputs(209)) or (inputs(141));
    layer0_outputs(3519) <= not(inputs(72)) or (inputs(59));
    layer0_outputs(3520) <= not((inputs(80)) or (inputs(68)));
    layer0_outputs(3521) <= (inputs(102)) or (inputs(246));
    layer0_outputs(3522) <= not((inputs(133)) xor (inputs(216)));
    layer0_outputs(3523) <= not(inputs(72)) or (inputs(109));
    layer0_outputs(3524) <= inputs(238);
    layer0_outputs(3525) <= not(inputs(152));
    layer0_outputs(3526) <= (inputs(216)) xor (inputs(193));
    layer0_outputs(3527) <= not((inputs(203)) xor (inputs(78)));
    layer0_outputs(3528) <= not((inputs(19)) xor (inputs(65)));
    layer0_outputs(3529) <= not(inputs(42)) or (inputs(235));
    layer0_outputs(3530) <= inputs(85);
    layer0_outputs(3531) <= inputs(128);
    layer0_outputs(3532) <= not(inputs(83));
    layer0_outputs(3533) <= not((inputs(195)) or (inputs(65)));
    layer0_outputs(3534) <= inputs(90);
    layer0_outputs(3535) <= (inputs(210)) and not (inputs(148));
    layer0_outputs(3536) <= (inputs(81)) xor (inputs(75));
    layer0_outputs(3537) <= inputs(92);
    layer0_outputs(3538) <= inputs(230);
    layer0_outputs(3539) <= not((inputs(51)) and (inputs(103)));
    layer0_outputs(3540) <= not((inputs(52)) xor (inputs(86)));
    layer0_outputs(3541) <= inputs(28);
    layer0_outputs(3542) <= (inputs(45)) xor (inputs(60));
    layer0_outputs(3543) <= (inputs(152)) xor (inputs(149));
    layer0_outputs(3544) <= not((inputs(42)) and (inputs(39)));
    layer0_outputs(3545) <= inputs(108);
    layer0_outputs(3546) <= (inputs(235)) and not (inputs(170));
    layer0_outputs(3547) <= not((inputs(8)) xor (inputs(182)));
    layer0_outputs(3548) <= not(inputs(174));
    layer0_outputs(3549) <= (inputs(195)) xor (inputs(72));
    layer0_outputs(3550) <= not(inputs(195)) or (inputs(143));
    layer0_outputs(3551) <= not(inputs(67)) or (inputs(140));
    layer0_outputs(3552) <= not(inputs(198));
    layer0_outputs(3553) <= (inputs(83)) and not (inputs(179));
    layer0_outputs(3554) <= not(inputs(57));
    layer0_outputs(3555) <= (inputs(140)) and (inputs(105));
    layer0_outputs(3556) <= (inputs(116)) and not (inputs(196));
    layer0_outputs(3557) <= not((inputs(121)) and (inputs(99)));
    layer0_outputs(3558) <= (inputs(240)) and not (inputs(220));
    layer0_outputs(3559) <= (inputs(78)) xor (inputs(52));
    layer0_outputs(3560) <= not(inputs(121));
    layer0_outputs(3561) <= (inputs(78)) xor (inputs(186));
    layer0_outputs(3562) <= inputs(206);
    layer0_outputs(3563) <= (inputs(222)) or (inputs(174));
    layer0_outputs(3564) <= (inputs(236)) and not (inputs(240));
    layer0_outputs(3565) <= inputs(194);
    layer0_outputs(3566) <= (inputs(83)) or (inputs(95));
    layer0_outputs(3567) <= not(inputs(14));
    layer0_outputs(3568) <= not(inputs(211));
    layer0_outputs(3569) <= not((inputs(4)) or (inputs(223)));
    layer0_outputs(3570) <= (inputs(151)) and (inputs(31));
    layer0_outputs(3571) <= (inputs(123)) and not (inputs(223));
    layer0_outputs(3572) <= not(inputs(248)) or (inputs(15));
    layer0_outputs(3573) <= not(inputs(54)) or (inputs(163));
    layer0_outputs(3574) <= not((inputs(68)) or (inputs(207)));
    layer0_outputs(3575) <= not((inputs(132)) xor (inputs(143)));
    layer0_outputs(3576) <= not(inputs(185));
    layer0_outputs(3577) <= not(inputs(167));
    layer0_outputs(3578) <= not(inputs(86)) or (inputs(41));
    layer0_outputs(3579) <= inputs(133);
    layer0_outputs(3580) <= not((inputs(255)) or (inputs(110)));
    layer0_outputs(3581) <= not(inputs(34));
    layer0_outputs(3582) <= inputs(247);
    layer0_outputs(3583) <= not((inputs(95)) or (inputs(208)));
    layer0_outputs(3584) <= inputs(226);
    layer0_outputs(3585) <= (inputs(58)) or (inputs(119));
    layer0_outputs(3586) <= inputs(60);
    layer0_outputs(3587) <= not(inputs(29)) or (inputs(248));
    layer0_outputs(3588) <= (inputs(109)) or (inputs(36));
    layer0_outputs(3589) <= inputs(56);
    layer0_outputs(3590) <= (inputs(188)) or (inputs(67));
    layer0_outputs(3591) <= (inputs(47)) or (inputs(181));
    layer0_outputs(3592) <= inputs(105);
    layer0_outputs(3593) <= inputs(186);
    layer0_outputs(3594) <= not((inputs(33)) or (inputs(30)));
    layer0_outputs(3595) <= (inputs(196)) or (inputs(48));
    layer0_outputs(3596) <= not(inputs(7));
    layer0_outputs(3597) <= not((inputs(239)) or (inputs(213)));
    layer0_outputs(3598) <= (inputs(22)) and (inputs(32));
    layer0_outputs(3599) <= inputs(73);
    layer0_outputs(3600) <= not(inputs(144));
    layer0_outputs(3601) <= not((inputs(71)) xor (inputs(98)));
    layer0_outputs(3602) <= not((inputs(77)) xor (inputs(205)));
    layer0_outputs(3603) <= not(inputs(4));
    layer0_outputs(3604) <= (inputs(42)) and not (inputs(181));
    layer0_outputs(3605) <= inputs(28);
    layer0_outputs(3606) <= inputs(205);
    layer0_outputs(3607) <= (inputs(130)) or (inputs(121));
    layer0_outputs(3608) <= '1';
    layer0_outputs(3609) <= not(inputs(93));
    layer0_outputs(3610) <= (inputs(137)) and not (inputs(81));
    layer0_outputs(3611) <= inputs(206);
    layer0_outputs(3612) <= not(inputs(90)) or (inputs(176));
    layer0_outputs(3613) <= (inputs(203)) xor (inputs(79));
    layer0_outputs(3614) <= not(inputs(101));
    layer0_outputs(3615) <= not((inputs(137)) xor (inputs(121)));
    layer0_outputs(3616) <= not((inputs(244)) or (inputs(73)));
    layer0_outputs(3617) <= not(inputs(57));
    layer0_outputs(3618) <= inputs(219);
    layer0_outputs(3619) <= not((inputs(70)) or (inputs(62)));
    layer0_outputs(3620) <= (inputs(105)) and not (inputs(199));
    layer0_outputs(3621) <= '1';
    layer0_outputs(3622) <= not(inputs(98)) or (inputs(170));
    layer0_outputs(3623) <= (inputs(211)) or (inputs(83));
    layer0_outputs(3624) <= not(inputs(248));
    layer0_outputs(3625) <= not((inputs(165)) xor (inputs(147)));
    layer0_outputs(3626) <= (inputs(230)) and not (inputs(0));
    layer0_outputs(3627) <= (inputs(234)) and not (inputs(18));
    layer0_outputs(3628) <= (inputs(213)) or (inputs(23));
    layer0_outputs(3629) <= not((inputs(24)) and (inputs(25)));
    layer0_outputs(3630) <= not(inputs(71)) or (inputs(18));
    layer0_outputs(3631) <= inputs(183);
    layer0_outputs(3632) <= not((inputs(1)) xor (inputs(239)));
    layer0_outputs(3633) <= inputs(167);
    layer0_outputs(3634) <= not((inputs(123)) xor (inputs(160)));
    layer0_outputs(3635) <= (inputs(79)) or (inputs(23));
    layer0_outputs(3636) <= (inputs(4)) and not (inputs(31));
    layer0_outputs(3637) <= not((inputs(236)) or (inputs(94)));
    layer0_outputs(3638) <= not(inputs(193));
    layer0_outputs(3639) <= (inputs(103)) and not (inputs(234));
    layer0_outputs(3640) <= (inputs(193)) or (inputs(85));
    layer0_outputs(3641) <= (inputs(123)) and not (inputs(186));
    layer0_outputs(3642) <= not((inputs(227)) and (inputs(227)));
    layer0_outputs(3643) <= not((inputs(100)) xor (inputs(156)));
    layer0_outputs(3644) <= not((inputs(88)) xor (inputs(86)));
    layer0_outputs(3645) <= not(inputs(169));
    layer0_outputs(3646) <= not((inputs(168)) or (inputs(78)));
    layer0_outputs(3647) <= (inputs(193)) and not (inputs(245));
    layer0_outputs(3648) <= not(inputs(130)) or (inputs(88));
    layer0_outputs(3649) <= not(inputs(105)) or (inputs(3));
    layer0_outputs(3650) <= not(inputs(5));
    layer0_outputs(3651) <= (inputs(214)) and not (inputs(240));
    layer0_outputs(3652) <= inputs(104);
    layer0_outputs(3653) <= (inputs(226)) xor (inputs(22));
    layer0_outputs(3654) <= inputs(40);
    layer0_outputs(3655) <= not((inputs(251)) xor (inputs(89)));
    layer0_outputs(3656) <= not(inputs(10));
    layer0_outputs(3657) <= (inputs(105)) and not (inputs(195));
    layer0_outputs(3658) <= not((inputs(106)) or (inputs(253)));
    layer0_outputs(3659) <= not(inputs(5)) or (inputs(249));
    layer0_outputs(3660) <= inputs(76);
    layer0_outputs(3661) <= (inputs(156)) xor (inputs(37));
    layer0_outputs(3662) <= not((inputs(141)) and (inputs(161)));
    layer0_outputs(3663) <= (inputs(237)) xor (inputs(148));
    layer0_outputs(3664) <= not(inputs(231)) or (inputs(15));
    layer0_outputs(3665) <= not(inputs(38));
    layer0_outputs(3666) <= not(inputs(92));
    layer0_outputs(3667) <= not(inputs(176)) or (inputs(9));
    layer0_outputs(3668) <= (inputs(113)) and (inputs(177));
    layer0_outputs(3669) <= not(inputs(25));
    layer0_outputs(3670) <= not(inputs(105));
    layer0_outputs(3671) <= not(inputs(124)) or (inputs(30));
    layer0_outputs(3672) <= (inputs(205)) and not (inputs(123));
    layer0_outputs(3673) <= (inputs(214)) xor (inputs(246));
    layer0_outputs(3674) <= (inputs(206)) xor (inputs(64));
    layer0_outputs(3675) <= inputs(71);
    layer0_outputs(3676) <= (inputs(107)) and not (inputs(174));
    layer0_outputs(3677) <= (inputs(116)) xor (inputs(43));
    layer0_outputs(3678) <= not(inputs(213));
    layer0_outputs(3679) <= not(inputs(135)) or (inputs(18));
    layer0_outputs(3680) <= not((inputs(80)) xor (inputs(235)));
    layer0_outputs(3681) <= not(inputs(79)) or (inputs(239));
    layer0_outputs(3682) <= (inputs(160)) and (inputs(114));
    layer0_outputs(3683) <= (inputs(150)) xor (inputs(211));
    layer0_outputs(3684) <= not(inputs(177));
    layer0_outputs(3685) <= inputs(72);
    layer0_outputs(3686) <= not((inputs(141)) xor (inputs(120)));
    layer0_outputs(3687) <= (inputs(227)) and not (inputs(103));
    layer0_outputs(3688) <= not(inputs(212)) or (inputs(74));
    layer0_outputs(3689) <= not(inputs(204));
    layer0_outputs(3690) <= (inputs(20)) and not (inputs(31));
    layer0_outputs(3691) <= (inputs(18)) and not (inputs(248));
    layer0_outputs(3692) <= (inputs(226)) and not (inputs(94));
    layer0_outputs(3693) <= not((inputs(42)) or (inputs(56)));
    layer0_outputs(3694) <= not(inputs(227));
    layer0_outputs(3695) <= not(inputs(244)) or (inputs(122));
    layer0_outputs(3696) <= inputs(120);
    layer0_outputs(3697) <= (inputs(168)) or (inputs(116));
    layer0_outputs(3698) <= inputs(105);
    layer0_outputs(3699) <= (inputs(155)) or (inputs(63));
    layer0_outputs(3700) <= not((inputs(87)) and (inputs(58)));
    layer0_outputs(3701) <= not(inputs(99));
    layer0_outputs(3702) <= not(inputs(246));
    layer0_outputs(3703) <= not((inputs(225)) or (inputs(40)));
    layer0_outputs(3704) <= inputs(236);
    layer0_outputs(3705) <= (inputs(182)) xor (inputs(84));
    layer0_outputs(3706) <= not((inputs(131)) and (inputs(209)));
    layer0_outputs(3707) <= not(inputs(182)) or (inputs(33));
    layer0_outputs(3708) <= (inputs(184)) and not (inputs(5));
    layer0_outputs(3709) <= (inputs(148)) xor (inputs(219));
    layer0_outputs(3710) <= (inputs(123)) or (inputs(73));
    layer0_outputs(3711) <= inputs(107);
    layer0_outputs(3712) <= not(inputs(178));
    layer0_outputs(3713) <= not(inputs(163));
    layer0_outputs(3714) <= not((inputs(240)) or (inputs(241)));
    layer0_outputs(3715) <= not(inputs(9));
    layer0_outputs(3716) <= (inputs(28)) xor (inputs(195));
    layer0_outputs(3717) <= not(inputs(195));
    layer0_outputs(3718) <= not(inputs(131));
    layer0_outputs(3719) <= inputs(229);
    layer0_outputs(3720) <= not(inputs(9)) or (inputs(49));
    layer0_outputs(3721) <= not(inputs(123));
    layer0_outputs(3722) <= not((inputs(126)) or (inputs(192)));
    layer0_outputs(3723) <= (inputs(2)) or (inputs(41));
    layer0_outputs(3724) <= not(inputs(147));
    layer0_outputs(3725) <= not((inputs(62)) xor (inputs(75)));
    layer0_outputs(3726) <= not(inputs(152));
    layer0_outputs(3727) <= not(inputs(86));
    layer0_outputs(3728) <= not(inputs(229));
    layer0_outputs(3729) <= inputs(226);
    layer0_outputs(3730) <= (inputs(184)) xor (inputs(134));
    layer0_outputs(3731) <= (inputs(37)) and not (inputs(96));
    layer0_outputs(3732) <= (inputs(243)) and not (inputs(31));
    layer0_outputs(3733) <= (inputs(154)) or (inputs(129));
    layer0_outputs(3734) <= not(inputs(127));
    layer0_outputs(3735) <= (inputs(250)) xor (inputs(91));
    layer0_outputs(3736) <= (inputs(122)) and not (inputs(65));
    layer0_outputs(3737) <= (inputs(50)) or (inputs(108));
    layer0_outputs(3738) <= inputs(89);
    layer0_outputs(3739) <= not(inputs(99));
    layer0_outputs(3740) <= not(inputs(126));
    layer0_outputs(3741) <= (inputs(63)) and not (inputs(239));
    layer0_outputs(3742) <= (inputs(198)) and (inputs(168));
    layer0_outputs(3743) <= (inputs(3)) or (inputs(127));
    layer0_outputs(3744) <= not(inputs(102)) or (inputs(126));
    layer0_outputs(3745) <= (inputs(0)) or (inputs(236));
    layer0_outputs(3746) <= not(inputs(77));
    layer0_outputs(3747) <= not((inputs(59)) or (inputs(198)));
    layer0_outputs(3748) <= not(inputs(97));
    layer0_outputs(3749) <= not(inputs(85));
    layer0_outputs(3750) <= inputs(230);
    layer0_outputs(3751) <= not((inputs(175)) xor (inputs(233)));
    layer0_outputs(3752) <= (inputs(70)) xor (inputs(39));
    layer0_outputs(3753) <= (inputs(191)) and not (inputs(174));
    layer0_outputs(3754) <= not((inputs(167)) or (inputs(102)));
    layer0_outputs(3755) <= inputs(86);
    layer0_outputs(3756) <= not(inputs(69));
    layer0_outputs(3757) <= not(inputs(27));
    layer0_outputs(3758) <= (inputs(17)) and not (inputs(52));
    layer0_outputs(3759) <= not(inputs(184));
    layer0_outputs(3760) <= not(inputs(242));
    layer0_outputs(3761) <= (inputs(126)) or (inputs(1));
    layer0_outputs(3762) <= not((inputs(143)) or (inputs(176)));
    layer0_outputs(3763) <= inputs(34);
    layer0_outputs(3764) <= inputs(50);
    layer0_outputs(3765) <= not((inputs(128)) and (inputs(81)));
    layer0_outputs(3766) <= (inputs(122)) or (inputs(88));
    layer0_outputs(3767) <= not(inputs(76));
    layer0_outputs(3768) <= (inputs(24)) and (inputs(11));
    layer0_outputs(3769) <= not(inputs(65));
    layer0_outputs(3770) <= not(inputs(82));
    layer0_outputs(3771) <= inputs(87);
    layer0_outputs(3772) <= not(inputs(184));
    layer0_outputs(3773) <= not(inputs(110)) or (inputs(7));
    layer0_outputs(3774) <= not((inputs(189)) xor (inputs(227)));
    layer0_outputs(3775) <= (inputs(249)) or (inputs(117));
    layer0_outputs(3776) <= (inputs(217)) or (inputs(196));
    layer0_outputs(3777) <= (inputs(220)) or (inputs(225));
    layer0_outputs(3778) <= (inputs(55)) and not (inputs(74));
    layer0_outputs(3779) <= inputs(15);
    layer0_outputs(3780) <= (inputs(44)) and not (inputs(206));
    layer0_outputs(3781) <= not(inputs(157)) or (inputs(255));
    layer0_outputs(3782) <= not((inputs(41)) or (inputs(16)));
    layer0_outputs(3783) <= (inputs(247)) and (inputs(229));
    layer0_outputs(3784) <= not(inputs(78));
    layer0_outputs(3785) <= not(inputs(248));
    layer0_outputs(3786) <= (inputs(15)) or (inputs(217));
    layer0_outputs(3787) <= not(inputs(103));
    layer0_outputs(3788) <= not(inputs(56)) or (inputs(1));
    layer0_outputs(3789) <= (inputs(188)) or (inputs(204));
    layer0_outputs(3790) <= not(inputs(119));
    layer0_outputs(3791) <= (inputs(204)) and (inputs(150));
    layer0_outputs(3792) <= not(inputs(133));
    layer0_outputs(3793) <= (inputs(120)) and not (inputs(100));
    layer0_outputs(3794) <= not((inputs(17)) and (inputs(98)));
    layer0_outputs(3795) <= (inputs(41)) and not (inputs(207));
    layer0_outputs(3796) <= not((inputs(124)) or (inputs(223)));
    layer0_outputs(3797) <= not((inputs(182)) or (inputs(151)));
    layer0_outputs(3798) <= (inputs(125)) xor (inputs(110));
    layer0_outputs(3799) <= not((inputs(164)) or (inputs(181)));
    layer0_outputs(3800) <= '0';
    layer0_outputs(3801) <= not((inputs(176)) or (inputs(54)));
    layer0_outputs(3802) <= not((inputs(117)) or (inputs(246)));
    layer0_outputs(3803) <= (inputs(107)) xor (inputs(141));
    layer0_outputs(3804) <= inputs(85);
    layer0_outputs(3805) <= not((inputs(37)) xor (inputs(158)));
    layer0_outputs(3806) <= (inputs(22)) and not (inputs(253));
    layer0_outputs(3807) <= (inputs(0)) xor (inputs(116));
    layer0_outputs(3808) <= inputs(248);
    layer0_outputs(3809) <= not((inputs(10)) or (inputs(187)));
    layer0_outputs(3810) <= inputs(183);
    layer0_outputs(3811) <= not(inputs(1));
    layer0_outputs(3812) <= not(inputs(7)) or (inputs(194));
    layer0_outputs(3813) <= not((inputs(195)) xor (inputs(250)));
    layer0_outputs(3814) <= (inputs(43)) and not (inputs(129));
    layer0_outputs(3815) <= not(inputs(145));
    layer0_outputs(3816) <= (inputs(148)) and (inputs(92));
    layer0_outputs(3817) <= (inputs(73)) or (inputs(224));
    layer0_outputs(3818) <= (inputs(47)) or (inputs(168));
    layer0_outputs(3819) <= (inputs(201)) or (inputs(174));
    layer0_outputs(3820) <= inputs(132);
    layer0_outputs(3821) <= not((inputs(12)) or (inputs(109)));
    layer0_outputs(3822) <= not(inputs(2)) or (inputs(2));
    layer0_outputs(3823) <= not((inputs(116)) xor (inputs(80)));
    layer0_outputs(3824) <= not((inputs(152)) xor (inputs(235)));
    layer0_outputs(3825) <= not((inputs(76)) and (inputs(107)));
    layer0_outputs(3826) <= not(inputs(105)) or (inputs(207));
    layer0_outputs(3827) <= (inputs(205)) and not (inputs(102));
    layer0_outputs(3828) <= inputs(111);
    layer0_outputs(3829) <= (inputs(153)) xor (inputs(148));
    layer0_outputs(3830) <= (inputs(37)) or (inputs(177));
    layer0_outputs(3831) <= not((inputs(53)) or (inputs(162)));
    layer0_outputs(3832) <= (inputs(88)) and not (inputs(253));
    layer0_outputs(3833) <= not(inputs(126));
    layer0_outputs(3834) <= (inputs(70)) xor (inputs(49));
    layer0_outputs(3835) <= not((inputs(202)) or (inputs(77)));
    layer0_outputs(3836) <= not(inputs(247));
    layer0_outputs(3837) <= (inputs(14)) and (inputs(74));
    layer0_outputs(3838) <= not(inputs(235)) or (inputs(171));
    layer0_outputs(3839) <= inputs(113);
    layer0_outputs(3840) <= not(inputs(12));
    layer0_outputs(3841) <= inputs(84);
    layer0_outputs(3842) <= (inputs(153)) xor (inputs(177));
    layer0_outputs(3843) <= not((inputs(5)) or (inputs(18)));
    layer0_outputs(3844) <= not(inputs(67));
    layer0_outputs(3845) <= inputs(22);
    layer0_outputs(3846) <= not((inputs(52)) or (inputs(216)));
    layer0_outputs(3847) <= (inputs(146)) or (inputs(183));
    layer0_outputs(3848) <= inputs(57);
    layer0_outputs(3849) <= (inputs(8)) and not (inputs(236));
    layer0_outputs(3850) <= (inputs(62)) xor (inputs(100));
    layer0_outputs(3851) <= not(inputs(42)) or (inputs(40));
    layer0_outputs(3852) <= inputs(181);
    layer0_outputs(3853) <= not(inputs(217)) or (inputs(31));
    layer0_outputs(3854) <= (inputs(151)) and not (inputs(156));
    layer0_outputs(3855) <= not((inputs(66)) or (inputs(162)));
    layer0_outputs(3856) <= inputs(79);
    layer0_outputs(3857) <= (inputs(140)) xor (inputs(155));
    layer0_outputs(3858) <= inputs(75);
    layer0_outputs(3859) <= not((inputs(252)) or (inputs(28)));
    layer0_outputs(3860) <= '0';
    layer0_outputs(3861) <= not(inputs(85)) or (inputs(177));
    layer0_outputs(3862) <= (inputs(2)) or (inputs(22));
    layer0_outputs(3863) <= inputs(128);
    layer0_outputs(3864) <= (inputs(33)) and (inputs(0));
    layer0_outputs(3865) <= not(inputs(68)) or (inputs(232));
    layer0_outputs(3866) <= not((inputs(82)) xor (inputs(174)));
    layer0_outputs(3867) <= inputs(214);
    layer0_outputs(3868) <= (inputs(98)) or (inputs(56));
    layer0_outputs(3869) <= (inputs(218)) and not (inputs(71));
    layer0_outputs(3870) <= (inputs(141)) and (inputs(143));
    layer0_outputs(3871) <= inputs(66);
    layer0_outputs(3872) <= not((inputs(231)) or (inputs(241)));
    layer0_outputs(3873) <= not((inputs(208)) or (inputs(234)));
    layer0_outputs(3874) <= (inputs(214)) and not (inputs(12));
    layer0_outputs(3875) <= not((inputs(32)) or (inputs(133)));
    layer0_outputs(3876) <= (inputs(200)) and not (inputs(26));
    layer0_outputs(3877) <= not((inputs(45)) xor (inputs(208)));
    layer0_outputs(3878) <= (inputs(233)) and not (inputs(1));
    layer0_outputs(3879) <= inputs(142);
    layer0_outputs(3880) <= (inputs(80)) and not (inputs(18));
    layer0_outputs(3881) <= not(inputs(44));
    layer0_outputs(3882) <= (inputs(96)) xor (inputs(92));
    layer0_outputs(3883) <= inputs(147);
    layer0_outputs(3884) <= not((inputs(48)) xor (inputs(185)));
    layer0_outputs(3885) <= '0';
    layer0_outputs(3886) <= (inputs(93)) or (inputs(242));
    layer0_outputs(3887) <= inputs(229);
    layer0_outputs(3888) <= not(inputs(172));
    layer0_outputs(3889) <= not(inputs(221));
    layer0_outputs(3890) <= not((inputs(201)) and (inputs(32)));
    layer0_outputs(3891) <= not((inputs(29)) and (inputs(46)));
    layer0_outputs(3892) <= not(inputs(247)) or (inputs(226));
    layer0_outputs(3893) <= inputs(247);
    layer0_outputs(3894) <= not(inputs(145)) or (inputs(217));
    layer0_outputs(3895) <= (inputs(170)) or (inputs(208));
    layer0_outputs(3896) <= (inputs(142)) and (inputs(128));
    layer0_outputs(3897) <= (inputs(40)) xor (inputs(78));
    layer0_outputs(3898) <= not((inputs(238)) or (inputs(161)));
    layer0_outputs(3899) <= (inputs(101)) and not (inputs(188));
    layer0_outputs(3900) <= not(inputs(68)) or (inputs(151));
    layer0_outputs(3901) <= not(inputs(137));
    layer0_outputs(3902) <= (inputs(58)) and not (inputs(177));
    layer0_outputs(3903) <= (inputs(124)) and not (inputs(225));
    layer0_outputs(3904) <= (inputs(69)) xor (inputs(41));
    layer0_outputs(3905) <= not(inputs(239)) or (inputs(178));
    layer0_outputs(3906) <= not(inputs(141)) or (inputs(253));
    layer0_outputs(3907) <= inputs(28);
    layer0_outputs(3908) <= inputs(121);
    layer0_outputs(3909) <= (inputs(107)) or (inputs(187));
    layer0_outputs(3910) <= not(inputs(22)) or (inputs(46));
    layer0_outputs(3911) <= not(inputs(131));
    layer0_outputs(3912) <= not(inputs(217)) or (inputs(58));
    layer0_outputs(3913) <= not((inputs(178)) or (inputs(150)));
    layer0_outputs(3914) <= (inputs(7)) and not (inputs(64));
    layer0_outputs(3915) <= not((inputs(63)) or (inputs(42)));
    layer0_outputs(3916) <= inputs(88);
    layer0_outputs(3917) <= (inputs(57)) and not (inputs(197));
    layer0_outputs(3918) <= inputs(171);
    layer0_outputs(3919) <= not((inputs(224)) xor (inputs(4)));
    layer0_outputs(3920) <= (inputs(28)) and not (inputs(192));
    layer0_outputs(3921) <= not(inputs(24)) or (inputs(98));
    layer0_outputs(3922) <= not(inputs(55));
    layer0_outputs(3923) <= not(inputs(170));
    layer0_outputs(3924) <= (inputs(125)) or (inputs(7));
    layer0_outputs(3925) <= not(inputs(132)) or (inputs(240));
    layer0_outputs(3926) <= (inputs(56)) and not (inputs(111));
    layer0_outputs(3927) <= not((inputs(205)) or (inputs(23)));
    layer0_outputs(3928) <= inputs(188);
    layer0_outputs(3929) <= not(inputs(10)) or (inputs(4));
    layer0_outputs(3930) <= not((inputs(158)) xor (inputs(3)));
    layer0_outputs(3931) <= not(inputs(229));
    layer0_outputs(3932) <= (inputs(4)) or (inputs(210));
    layer0_outputs(3933) <= (inputs(31)) or (inputs(29));
    layer0_outputs(3934) <= (inputs(86)) xor (inputs(49));
    layer0_outputs(3935) <= inputs(46);
    layer0_outputs(3936) <= inputs(109);
    layer0_outputs(3937) <= not((inputs(189)) or (inputs(185)));
    layer0_outputs(3938) <= not((inputs(214)) xor (inputs(147)));
    layer0_outputs(3939) <= (inputs(134)) and not (inputs(111));
    layer0_outputs(3940) <= not(inputs(122)) or (inputs(96));
    layer0_outputs(3941) <= not(inputs(55)) or (inputs(12));
    layer0_outputs(3942) <= inputs(170);
    layer0_outputs(3943) <= not(inputs(92));
    layer0_outputs(3944) <= not(inputs(162));
    layer0_outputs(3945) <= inputs(133);
    layer0_outputs(3946) <= (inputs(204)) or (inputs(107));
    layer0_outputs(3947) <= not((inputs(238)) xor (inputs(171)));
    layer0_outputs(3948) <= not(inputs(167)) or (inputs(49));
    layer0_outputs(3949) <= (inputs(207)) or (inputs(214));
    layer0_outputs(3950) <= (inputs(105)) and not (inputs(43));
    layer0_outputs(3951) <= not((inputs(204)) xor (inputs(23)));
    layer0_outputs(3952) <= inputs(251);
    layer0_outputs(3953) <= inputs(233);
    layer0_outputs(3954) <= (inputs(100)) and not (inputs(53));
    layer0_outputs(3955) <= inputs(165);
    layer0_outputs(3956) <= inputs(96);
    layer0_outputs(3957) <= not((inputs(69)) xor (inputs(218)));
    layer0_outputs(3958) <= inputs(144);
    layer0_outputs(3959) <= inputs(21);
    layer0_outputs(3960) <= (inputs(182)) and not (inputs(66));
    layer0_outputs(3961) <= (inputs(253)) and not (inputs(55));
    layer0_outputs(3962) <= not(inputs(28)) or (inputs(71));
    layer0_outputs(3963) <= (inputs(58)) or (inputs(48));
    layer0_outputs(3964) <= not(inputs(170));
    layer0_outputs(3965) <= not(inputs(24));
    layer0_outputs(3966) <= (inputs(48)) or (inputs(121));
    layer0_outputs(3967) <= (inputs(23)) xor (inputs(71));
    layer0_outputs(3968) <= not((inputs(192)) or (inputs(22)));
    layer0_outputs(3969) <= (inputs(115)) or (inputs(208));
    layer0_outputs(3970) <= not(inputs(124));
    layer0_outputs(3971) <= (inputs(53)) and (inputs(205));
    layer0_outputs(3972) <= inputs(137);
    layer0_outputs(3973) <= (inputs(57)) or (inputs(32));
    layer0_outputs(3974) <= (inputs(222)) xor (inputs(123));
    layer0_outputs(3975) <= not(inputs(185));
    layer0_outputs(3976) <= not(inputs(121));
    layer0_outputs(3977) <= (inputs(182)) or (inputs(205));
    layer0_outputs(3978) <= '0';
    layer0_outputs(3979) <= (inputs(237)) and not (inputs(179));
    layer0_outputs(3980) <= not(inputs(167)) or (inputs(176));
    layer0_outputs(3981) <= not((inputs(193)) or (inputs(64)));
    layer0_outputs(3982) <= (inputs(214)) and (inputs(41));
    layer0_outputs(3983) <= inputs(146);
    layer0_outputs(3984) <= (inputs(183)) and not (inputs(49));
    layer0_outputs(3985) <= (inputs(146)) xor (inputs(239));
    layer0_outputs(3986) <= (inputs(128)) xor (inputs(181));
    layer0_outputs(3987) <= not(inputs(81));
    layer0_outputs(3988) <= inputs(22);
    layer0_outputs(3989) <= (inputs(87)) xor (inputs(83));
    layer0_outputs(3990) <= not((inputs(117)) or (inputs(142)));
    layer0_outputs(3991) <= inputs(122);
    layer0_outputs(3992) <= (inputs(156)) or (inputs(130));
    layer0_outputs(3993) <= not(inputs(219));
    layer0_outputs(3994) <= not(inputs(176));
    layer0_outputs(3995) <= inputs(140);
    layer0_outputs(3996) <= (inputs(214)) and not (inputs(53));
    layer0_outputs(3997) <= not((inputs(203)) and (inputs(6)));
    layer0_outputs(3998) <= not((inputs(44)) xor (inputs(224)));
    layer0_outputs(3999) <= not(inputs(187));
    layer0_outputs(4000) <= inputs(26);
    layer0_outputs(4001) <= (inputs(133)) and not (inputs(235));
    layer0_outputs(4002) <= (inputs(188)) and not (inputs(78));
    layer0_outputs(4003) <= (inputs(140)) and (inputs(70));
    layer0_outputs(4004) <= '0';
    layer0_outputs(4005) <= not(inputs(99));
    layer0_outputs(4006) <= not((inputs(28)) xor (inputs(46)));
    layer0_outputs(4007) <= inputs(60);
    layer0_outputs(4008) <= (inputs(4)) or (inputs(169));
    layer0_outputs(4009) <= not(inputs(228));
    layer0_outputs(4010) <= not((inputs(231)) or (inputs(11)));
    layer0_outputs(4011) <= not((inputs(167)) xor (inputs(120)));
    layer0_outputs(4012) <= inputs(224);
    layer0_outputs(4013) <= not(inputs(43)) or (inputs(69));
    layer0_outputs(4014) <= not(inputs(166)) or (inputs(220));
    layer0_outputs(4015) <= inputs(200);
    layer0_outputs(4016) <= not((inputs(197)) or (inputs(63)));
    layer0_outputs(4017) <= not(inputs(41)) or (inputs(141));
    layer0_outputs(4018) <= not(inputs(155));
    layer0_outputs(4019) <= not((inputs(5)) xor (inputs(79)));
    layer0_outputs(4020) <= (inputs(112)) xor (inputs(21));
    layer0_outputs(4021) <= not(inputs(134));
    layer0_outputs(4022) <= (inputs(16)) or (inputs(5));
    layer0_outputs(4023) <= not((inputs(39)) or (inputs(158)));
    layer0_outputs(4024) <= (inputs(53)) xor (inputs(244));
    layer0_outputs(4025) <= not(inputs(165)) or (inputs(159));
    layer0_outputs(4026) <= not((inputs(58)) xor (inputs(124)));
    layer0_outputs(4027) <= inputs(102);
    layer0_outputs(4028) <= (inputs(236)) or (inputs(171));
    layer0_outputs(4029) <= not(inputs(252)) or (inputs(31));
    layer0_outputs(4030) <= not(inputs(228));
    layer0_outputs(4031) <= not(inputs(83));
    layer0_outputs(4032) <= not((inputs(96)) or (inputs(205)));
    layer0_outputs(4033) <= (inputs(187)) and not (inputs(9));
    layer0_outputs(4034) <= not((inputs(46)) or (inputs(192)));
    layer0_outputs(4035) <= not(inputs(220));
    layer0_outputs(4036) <= inputs(163);
    layer0_outputs(4037) <= (inputs(137)) or (inputs(156));
    layer0_outputs(4038) <= not(inputs(212));
    layer0_outputs(4039) <= (inputs(141)) xor (inputs(149));
    layer0_outputs(4040) <= (inputs(173)) or (inputs(13));
    layer0_outputs(4041) <= (inputs(141)) and not (inputs(122));
    layer0_outputs(4042) <= (inputs(235)) and (inputs(118));
    layer0_outputs(4043) <= not((inputs(235)) and (inputs(233)));
    layer0_outputs(4044) <= not(inputs(162));
    layer0_outputs(4045) <= inputs(244);
    layer0_outputs(4046) <= not(inputs(103));
    layer0_outputs(4047) <= (inputs(177)) or (inputs(68));
    layer0_outputs(4048) <= (inputs(137)) and not (inputs(175));
    layer0_outputs(4049) <= (inputs(120)) or (inputs(194));
    layer0_outputs(4050) <= not(inputs(27)) or (inputs(75));
    layer0_outputs(4051) <= (inputs(126)) and not (inputs(103));
    layer0_outputs(4052) <= inputs(163);
    layer0_outputs(4053) <= inputs(144);
    layer0_outputs(4054) <= (inputs(56)) or (inputs(24));
    layer0_outputs(4055) <= (inputs(105)) or (inputs(248));
    layer0_outputs(4056) <= inputs(10);
    layer0_outputs(4057) <= (inputs(8)) and not (inputs(128));
    layer0_outputs(4058) <= inputs(90);
    layer0_outputs(4059) <= inputs(181);
    layer0_outputs(4060) <= not(inputs(63));
    layer0_outputs(4061) <= not(inputs(201)) or (inputs(123));
    layer0_outputs(4062) <= not((inputs(174)) xor (inputs(254)));
    layer0_outputs(4063) <= (inputs(61)) xor (inputs(180));
    layer0_outputs(4064) <= inputs(116);
    layer0_outputs(4065) <= not(inputs(232));
    layer0_outputs(4066) <= not((inputs(27)) xor (inputs(0)));
    layer0_outputs(4067) <= not(inputs(39)) or (inputs(241));
    layer0_outputs(4068) <= not((inputs(128)) xor (inputs(163)));
    layer0_outputs(4069) <= not(inputs(57));
    layer0_outputs(4070) <= not(inputs(212)) or (inputs(240));
    layer0_outputs(4071) <= inputs(153);
    layer0_outputs(4072) <= (inputs(32)) or (inputs(162));
    layer0_outputs(4073) <= (inputs(226)) xor (inputs(206));
    layer0_outputs(4074) <= not(inputs(93)) or (inputs(128));
    layer0_outputs(4075) <= not((inputs(147)) or (inputs(40)));
    layer0_outputs(4076) <= '1';
    layer0_outputs(4077) <= not(inputs(180)) or (inputs(249));
    layer0_outputs(4078) <= (inputs(72)) or (inputs(215));
    layer0_outputs(4079) <= not(inputs(66));
    layer0_outputs(4080) <= not(inputs(169));
    layer0_outputs(4081) <= not(inputs(117));
    layer0_outputs(4082) <= not((inputs(110)) xor (inputs(205)));
    layer0_outputs(4083) <= not((inputs(221)) or (inputs(235)));
    layer0_outputs(4084) <= not(inputs(101));
    layer0_outputs(4085) <= not((inputs(134)) or (inputs(177)));
    layer0_outputs(4086) <= inputs(192);
    layer0_outputs(4087) <= inputs(71);
    layer0_outputs(4088) <= not(inputs(46));
    layer0_outputs(4089) <= (inputs(21)) xor (inputs(53));
    layer0_outputs(4090) <= inputs(36);
    layer0_outputs(4091) <= not((inputs(156)) or (inputs(246)));
    layer0_outputs(4092) <= (inputs(209)) and not (inputs(159));
    layer0_outputs(4093) <= (inputs(107)) and not (inputs(66));
    layer0_outputs(4094) <= not(inputs(245));
    layer0_outputs(4095) <= not((inputs(137)) and (inputs(56)));
    layer0_outputs(4096) <= inputs(197);
    layer0_outputs(4097) <= not(inputs(101));
    layer0_outputs(4098) <= (inputs(48)) and not (inputs(239));
    layer0_outputs(4099) <= (inputs(99)) and not (inputs(33));
    layer0_outputs(4100) <= not((inputs(178)) and (inputs(166)));
    layer0_outputs(4101) <= inputs(84);
    layer0_outputs(4102) <= (inputs(218)) and not (inputs(83));
    layer0_outputs(4103) <= not(inputs(213)) or (inputs(46));
    layer0_outputs(4104) <= not(inputs(75));
    layer0_outputs(4105) <= (inputs(161)) xor (inputs(164));
    layer0_outputs(4106) <= inputs(148);
    layer0_outputs(4107) <= not(inputs(114));
    layer0_outputs(4108) <= not((inputs(53)) xor (inputs(148)));
    layer0_outputs(4109) <= (inputs(227)) or (inputs(98));
    layer0_outputs(4110) <= not((inputs(158)) xor (inputs(136)));
    layer0_outputs(4111) <= (inputs(242)) xor (inputs(34));
    layer0_outputs(4112) <= inputs(168);
    layer0_outputs(4113) <= (inputs(41)) and not (inputs(79));
    layer0_outputs(4114) <= (inputs(122)) and not (inputs(232));
    layer0_outputs(4115) <= not((inputs(36)) or (inputs(181)));
    layer0_outputs(4116) <= inputs(87);
    layer0_outputs(4117) <= (inputs(198)) xor (inputs(230));
    layer0_outputs(4118) <= inputs(47);
    layer0_outputs(4119) <= inputs(175);
    layer0_outputs(4120) <= (inputs(121)) and not (inputs(66));
    layer0_outputs(4121) <= not((inputs(3)) xor (inputs(45)));
    layer0_outputs(4122) <= (inputs(103)) xor (inputs(153));
    layer0_outputs(4123) <= not(inputs(99)) or (inputs(35));
    layer0_outputs(4124) <= (inputs(56)) xor (inputs(8));
    layer0_outputs(4125) <= not(inputs(43)) or (inputs(252));
    layer0_outputs(4126) <= not(inputs(122));
    layer0_outputs(4127) <= not(inputs(14));
    layer0_outputs(4128) <= not(inputs(153));
    layer0_outputs(4129) <= (inputs(243)) and not (inputs(65));
    layer0_outputs(4130) <= (inputs(156)) xor (inputs(213));
    layer0_outputs(4131) <= inputs(229);
    layer0_outputs(4132) <= '1';
    layer0_outputs(4133) <= not((inputs(42)) xor (inputs(202)));
    layer0_outputs(4134) <= not(inputs(72)) or (inputs(248));
    layer0_outputs(4135) <= (inputs(165)) xor (inputs(144));
    layer0_outputs(4136) <= (inputs(180)) and not (inputs(46));
    layer0_outputs(4137) <= not(inputs(228)) or (inputs(78));
    layer0_outputs(4138) <= not(inputs(36));
    layer0_outputs(4139) <= not(inputs(85)) or (inputs(191));
    layer0_outputs(4140) <= (inputs(101)) xor (inputs(176));
    layer0_outputs(4141) <= not(inputs(27)) or (inputs(119));
    layer0_outputs(4142) <= (inputs(193)) and not (inputs(140));
    layer0_outputs(4143) <= (inputs(253)) and not (inputs(50));
    layer0_outputs(4144) <= not((inputs(142)) xor (inputs(131)));
    layer0_outputs(4145) <= (inputs(122)) xor (inputs(185));
    layer0_outputs(4146) <= not((inputs(118)) xor (inputs(172)));
    layer0_outputs(4147) <= not(inputs(198));
    layer0_outputs(4148) <= inputs(209);
    layer0_outputs(4149) <= not((inputs(169)) xor (inputs(136)));
    layer0_outputs(4150) <= (inputs(167)) and not (inputs(185));
    layer0_outputs(4151) <= not(inputs(100));
    layer0_outputs(4152) <= inputs(247);
    layer0_outputs(4153) <= not((inputs(62)) and (inputs(62)));
    layer0_outputs(4154) <= inputs(39);
    layer0_outputs(4155) <= not(inputs(198));
    layer0_outputs(4156) <= not(inputs(108));
    layer0_outputs(4157) <= not((inputs(249)) xor (inputs(124)));
    layer0_outputs(4158) <= not(inputs(228)) or (inputs(93));
    layer0_outputs(4159) <= not(inputs(97));
    layer0_outputs(4160) <= not(inputs(183));
    layer0_outputs(4161) <= not(inputs(124)) or (inputs(225));
    layer0_outputs(4162) <= not((inputs(160)) or (inputs(128)));
    layer0_outputs(4163) <= not((inputs(64)) or (inputs(212)));
    layer0_outputs(4164) <= inputs(204);
    layer0_outputs(4165) <= (inputs(83)) and not (inputs(165));
    layer0_outputs(4166) <= inputs(153);
    layer0_outputs(4167) <= not((inputs(71)) or (inputs(187)));
    layer0_outputs(4168) <= not((inputs(222)) and (inputs(132)));
    layer0_outputs(4169) <= not((inputs(90)) or (inputs(4)));
    layer0_outputs(4170) <= not(inputs(245));
    layer0_outputs(4171) <= (inputs(73)) and (inputs(58));
    layer0_outputs(4172) <= not((inputs(203)) xor (inputs(227)));
    layer0_outputs(4173) <= not(inputs(154)) or (inputs(164));
    layer0_outputs(4174) <= (inputs(57)) and not (inputs(80));
    layer0_outputs(4175) <= inputs(106);
    layer0_outputs(4176) <= (inputs(138)) xor (inputs(142));
    layer0_outputs(4177) <= inputs(230);
    layer0_outputs(4178) <= inputs(229);
    layer0_outputs(4179) <= not((inputs(75)) xor (inputs(95)));
    layer0_outputs(4180) <= not(inputs(190));
    layer0_outputs(4181) <= inputs(9);
    layer0_outputs(4182) <= inputs(119);
    layer0_outputs(4183) <= (inputs(229)) or (inputs(220));
    layer0_outputs(4184) <= not((inputs(35)) xor (inputs(81)));
    layer0_outputs(4185) <= not((inputs(111)) xor (inputs(201)));
    layer0_outputs(4186) <= inputs(205);
    layer0_outputs(4187) <= not((inputs(148)) xor (inputs(31)));
    layer0_outputs(4188) <= inputs(56);
    layer0_outputs(4189) <= (inputs(247)) and not (inputs(237));
    layer0_outputs(4190) <= not(inputs(136));
    layer0_outputs(4191) <= not(inputs(122));
    layer0_outputs(4192) <= not(inputs(215));
    layer0_outputs(4193) <= not(inputs(119));
    layer0_outputs(4194) <= not(inputs(158));
    layer0_outputs(4195) <= (inputs(228)) or (inputs(189));
    layer0_outputs(4196) <= not(inputs(104)) or (inputs(142));
    layer0_outputs(4197) <= not(inputs(222)) or (inputs(168));
    layer0_outputs(4198) <= not((inputs(196)) or (inputs(48)));
    layer0_outputs(4199) <= inputs(149);
    layer0_outputs(4200) <= inputs(54);
    layer0_outputs(4201) <= inputs(5);
    layer0_outputs(4202) <= (inputs(199)) and not (inputs(168));
    layer0_outputs(4203) <= not((inputs(51)) xor (inputs(64)));
    layer0_outputs(4204) <= inputs(48);
    layer0_outputs(4205) <= not(inputs(233));
    layer0_outputs(4206) <= not(inputs(156));
    layer0_outputs(4207) <= (inputs(15)) xor (inputs(150));
    layer0_outputs(4208) <= not((inputs(96)) and (inputs(41)));
    layer0_outputs(4209) <= (inputs(14)) and not (inputs(32));
    layer0_outputs(4210) <= (inputs(69)) xor (inputs(206));
    layer0_outputs(4211) <= not((inputs(69)) or (inputs(226)));
    layer0_outputs(4212) <= (inputs(140)) xor (inputs(207));
    layer0_outputs(4213) <= (inputs(105)) xor (inputs(190));
    layer0_outputs(4214) <= not((inputs(39)) and (inputs(170)));
    layer0_outputs(4215) <= not((inputs(221)) or (inputs(169)));
    layer0_outputs(4216) <= (inputs(15)) and not (inputs(155));
    layer0_outputs(4217) <= inputs(161);
    layer0_outputs(4218) <= not((inputs(162)) xor (inputs(219)));
    layer0_outputs(4219) <= not(inputs(89)) or (inputs(202));
    layer0_outputs(4220) <= not(inputs(242)) or (inputs(82));
    layer0_outputs(4221) <= inputs(172);
    layer0_outputs(4222) <= not((inputs(84)) xor (inputs(49)));
    layer0_outputs(4223) <= not(inputs(104));
    layer0_outputs(4224) <= (inputs(170)) xor (inputs(113));
    layer0_outputs(4225) <= (inputs(95)) xor (inputs(203));
    layer0_outputs(4226) <= (inputs(80)) or (inputs(155));
    layer0_outputs(4227) <= (inputs(39)) and not (inputs(141));
    layer0_outputs(4228) <= (inputs(137)) or (inputs(83));
    layer0_outputs(4229) <= (inputs(212)) and not (inputs(59));
    layer0_outputs(4230) <= (inputs(131)) and not (inputs(46));
    layer0_outputs(4231) <= not((inputs(237)) or (inputs(113)));
    layer0_outputs(4232) <= (inputs(72)) or (inputs(50));
    layer0_outputs(4233) <= inputs(26);
    layer0_outputs(4234) <= not((inputs(17)) or (inputs(182)));
    layer0_outputs(4235) <= not((inputs(104)) xor (inputs(152)));
    layer0_outputs(4236) <= not(inputs(158)) or (inputs(68));
    layer0_outputs(4237) <= not((inputs(181)) or (inputs(97)));
    layer0_outputs(4238) <= not(inputs(231));
    layer0_outputs(4239) <= not(inputs(234)) or (inputs(30));
    layer0_outputs(4240) <= inputs(142);
    layer0_outputs(4241) <= inputs(41);
    layer0_outputs(4242) <= not(inputs(81));
    layer0_outputs(4243) <= (inputs(217)) and not (inputs(82));
    layer0_outputs(4244) <= not(inputs(27));
    layer0_outputs(4245) <= not(inputs(234));
    layer0_outputs(4246) <= not(inputs(97));
    layer0_outputs(4247) <= not(inputs(215));
    layer0_outputs(4248) <= not((inputs(240)) xor (inputs(123)));
    layer0_outputs(4249) <= not((inputs(161)) xor (inputs(27)));
    layer0_outputs(4250) <= (inputs(39)) and not (inputs(208));
    layer0_outputs(4251) <= inputs(173);
    layer0_outputs(4252) <= not(inputs(78)) or (inputs(176));
    layer0_outputs(4253) <= (inputs(196)) or (inputs(181));
    layer0_outputs(4254) <= inputs(74);
    layer0_outputs(4255) <= (inputs(238)) and (inputs(195));
    layer0_outputs(4256) <= not(inputs(206));
    layer0_outputs(4257) <= not((inputs(140)) xor (inputs(148)));
    layer0_outputs(4258) <= not(inputs(178)) or (inputs(98));
    layer0_outputs(4259) <= (inputs(8)) and not (inputs(244));
    layer0_outputs(4260) <= inputs(174);
    layer0_outputs(4261) <= not(inputs(6)) or (inputs(203));
    layer0_outputs(4262) <= not(inputs(170)) or (inputs(221));
    layer0_outputs(4263) <= not((inputs(83)) or (inputs(222)));
    layer0_outputs(4264) <= not((inputs(70)) xor (inputs(157)));
    layer0_outputs(4265) <= not((inputs(184)) or (inputs(70)));
    layer0_outputs(4266) <= '1';
    layer0_outputs(4267) <= (inputs(108)) and not (inputs(158));
    layer0_outputs(4268) <= not((inputs(220)) xor (inputs(179)));
    layer0_outputs(4269) <= (inputs(187)) or (inputs(132));
    layer0_outputs(4270) <= inputs(187);
    layer0_outputs(4271) <= (inputs(202)) or (inputs(163));
    layer0_outputs(4272) <= not(inputs(167));
    layer0_outputs(4273) <= not((inputs(30)) xor (inputs(152)));
    layer0_outputs(4274) <= not((inputs(215)) and (inputs(151)));
    layer0_outputs(4275) <= not(inputs(132));
    layer0_outputs(4276) <= (inputs(199)) or (inputs(179));
    layer0_outputs(4277) <= (inputs(255)) or (inputs(193));
    layer0_outputs(4278) <= not(inputs(148));
    layer0_outputs(4279) <= not(inputs(117));
    layer0_outputs(4280) <= not((inputs(94)) xor (inputs(204)));
    layer0_outputs(4281) <= not((inputs(1)) or (inputs(235)));
    layer0_outputs(4282) <= not(inputs(203)) or (inputs(144));
    layer0_outputs(4283) <= (inputs(203)) and not (inputs(49));
    layer0_outputs(4284) <= not((inputs(12)) xor (inputs(182)));
    layer0_outputs(4285) <= not(inputs(214));
    layer0_outputs(4286) <= not((inputs(191)) xor (inputs(53)));
    layer0_outputs(4287) <= (inputs(150)) and not (inputs(248));
    layer0_outputs(4288) <= not((inputs(123)) or (inputs(153)));
    layer0_outputs(4289) <= inputs(105);
    layer0_outputs(4290) <= (inputs(37)) and (inputs(250));
    layer0_outputs(4291) <= inputs(233);
    layer0_outputs(4292) <= not(inputs(163));
    layer0_outputs(4293) <= (inputs(118)) xor (inputs(233));
    layer0_outputs(4294) <= not((inputs(172)) or (inputs(144)));
    layer0_outputs(4295) <= (inputs(150)) or (inputs(7));
    layer0_outputs(4296) <= not(inputs(86)) or (inputs(108));
    layer0_outputs(4297) <= not(inputs(245)) or (inputs(51));
    layer0_outputs(4298) <= (inputs(115)) and not (inputs(40));
    layer0_outputs(4299) <= inputs(99);
    layer0_outputs(4300) <= not(inputs(219));
    layer0_outputs(4301) <= inputs(216);
    layer0_outputs(4302) <= not(inputs(21));
    layer0_outputs(4303) <= inputs(156);
    layer0_outputs(4304) <= not((inputs(219)) or (inputs(234)));
    layer0_outputs(4305) <= (inputs(233)) and not (inputs(1));
    layer0_outputs(4306) <= not(inputs(135));
    layer0_outputs(4307) <= not(inputs(174));
    layer0_outputs(4308) <= (inputs(74)) and not (inputs(206));
    layer0_outputs(4309) <= inputs(23);
    layer0_outputs(4310) <= (inputs(74)) and not (inputs(159));
    layer0_outputs(4311) <= (inputs(246)) and (inputs(187));
    layer0_outputs(4312) <= not((inputs(180)) or (inputs(199)));
    layer0_outputs(4313) <= inputs(204);
    layer0_outputs(4314) <= (inputs(117)) and not (inputs(193));
    layer0_outputs(4315) <= (inputs(196)) xor (inputs(225));
    layer0_outputs(4316) <= (inputs(200)) and not (inputs(0));
    layer0_outputs(4317) <= inputs(228);
    layer0_outputs(4318) <= not(inputs(105)) or (inputs(110));
    layer0_outputs(4319) <= inputs(176);
    layer0_outputs(4320) <= (inputs(207)) xor (inputs(61));
    layer0_outputs(4321) <= (inputs(91)) or (inputs(18));
    layer0_outputs(4322) <= not(inputs(251));
    layer0_outputs(4323) <= not((inputs(37)) or (inputs(30)));
    layer0_outputs(4324) <= not(inputs(123)) or (inputs(112));
    layer0_outputs(4325) <= not((inputs(180)) xor (inputs(47)));
    layer0_outputs(4326) <= (inputs(100)) xor (inputs(146));
    layer0_outputs(4327) <= not(inputs(88)) or (inputs(27));
    layer0_outputs(4328) <= not((inputs(59)) xor (inputs(14)));
    layer0_outputs(4329) <= not(inputs(178));
    layer0_outputs(4330) <= (inputs(99)) and not (inputs(162));
    layer0_outputs(4331) <= not(inputs(184));
    layer0_outputs(4332) <= (inputs(82)) or (inputs(152));
    layer0_outputs(4333) <= not(inputs(21)) or (inputs(204));
    layer0_outputs(4334) <= inputs(36);
    layer0_outputs(4335) <= inputs(101);
    layer0_outputs(4336) <= (inputs(111)) or (inputs(179));
    layer0_outputs(4337) <= (inputs(166)) xor (inputs(69));
    layer0_outputs(4338) <= (inputs(186)) xor (inputs(68));
    layer0_outputs(4339) <= not((inputs(139)) or (inputs(75)));
    layer0_outputs(4340) <= not((inputs(222)) or (inputs(63)));
    layer0_outputs(4341) <= not((inputs(65)) xor (inputs(42)));
    layer0_outputs(4342) <= inputs(76);
    layer0_outputs(4343) <= not((inputs(42)) and (inputs(37)));
    layer0_outputs(4344) <= not(inputs(171));
    layer0_outputs(4345) <= not((inputs(37)) or (inputs(93)));
    layer0_outputs(4346) <= not((inputs(192)) or (inputs(37)));
    layer0_outputs(4347) <= not((inputs(141)) or (inputs(130)));
    layer0_outputs(4348) <= (inputs(26)) xor (inputs(143));
    layer0_outputs(4349) <= (inputs(7)) xor (inputs(242));
    layer0_outputs(4350) <= (inputs(122)) or (inputs(93));
    layer0_outputs(4351) <= inputs(91);
    layer0_outputs(4352) <= (inputs(138)) xor (inputs(200));
    layer0_outputs(4353) <= (inputs(197)) or (inputs(193));
    layer0_outputs(4354) <= (inputs(149)) xor (inputs(229));
    layer0_outputs(4355) <= inputs(181);
    layer0_outputs(4356) <= (inputs(76)) xor (inputs(94));
    layer0_outputs(4357) <= inputs(162);
    layer0_outputs(4358) <= not((inputs(166)) xor (inputs(55)));
    layer0_outputs(4359) <= inputs(147);
    layer0_outputs(4360) <= not(inputs(167));
    layer0_outputs(4361) <= not(inputs(57)) or (inputs(244));
    layer0_outputs(4362) <= not(inputs(249));
    layer0_outputs(4363) <= (inputs(203)) and not (inputs(30));
    layer0_outputs(4364) <= not(inputs(189)) or (inputs(98));
    layer0_outputs(4365) <= not(inputs(138)) or (inputs(212));
    layer0_outputs(4366) <= not(inputs(44)) or (inputs(203));
    layer0_outputs(4367) <= not((inputs(140)) xor (inputs(171)));
    layer0_outputs(4368) <= (inputs(243)) xor (inputs(58));
    layer0_outputs(4369) <= (inputs(181)) or (inputs(43));
    layer0_outputs(4370) <= (inputs(223)) or (inputs(136));
    layer0_outputs(4371) <= (inputs(205)) or (inputs(141));
    layer0_outputs(4372) <= inputs(122);
    layer0_outputs(4373) <= (inputs(89)) and not (inputs(110));
    layer0_outputs(4374) <= inputs(178);
    layer0_outputs(4375) <= not(inputs(168)) or (inputs(132));
    layer0_outputs(4376) <= not(inputs(230)) or (inputs(65));
    layer0_outputs(4377) <= not((inputs(66)) or (inputs(82)));
    layer0_outputs(4378) <= not(inputs(191));
    layer0_outputs(4379) <= not(inputs(213)) or (inputs(23));
    layer0_outputs(4380) <= (inputs(202)) xor (inputs(52));
    layer0_outputs(4381) <= (inputs(220)) and not (inputs(241));
    layer0_outputs(4382) <= not(inputs(109));
    layer0_outputs(4383) <= inputs(141);
    layer0_outputs(4384) <= (inputs(26)) or (inputs(94));
    layer0_outputs(4385) <= not((inputs(255)) xor (inputs(155)));
    layer0_outputs(4386) <= not(inputs(176));
    layer0_outputs(4387) <= (inputs(228)) and not (inputs(91));
    layer0_outputs(4388) <= (inputs(17)) or (inputs(51));
    layer0_outputs(4389) <= (inputs(148)) and (inputs(149));
    layer0_outputs(4390) <= (inputs(188)) or (inputs(164));
    layer0_outputs(4391) <= (inputs(95)) and not (inputs(102));
    layer0_outputs(4392) <= (inputs(234)) or (inputs(192));
    layer0_outputs(4393) <= inputs(148);
    layer0_outputs(4394) <= inputs(53);
    layer0_outputs(4395) <= not(inputs(215));
    layer0_outputs(4396) <= inputs(226);
    layer0_outputs(4397) <= (inputs(211)) and not (inputs(207));
    layer0_outputs(4398) <= not((inputs(175)) xor (inputs(74)));
    layer0_outputs(4399) <= (inputs(96)) or (inputs(230));
    layer0_outputs(4400) <= not(inputs(207)) or (inputs(175));
    layer0_outputs(4401) <= (inputs(161)) xor (inputs(130));
    layer0_outputs(4402) <= not((inputs(73)) xor (inputs(126)));
    layer0_outputs(4403) <= not(inputs(81));
    layer0_outputs(4404) <= (inputs(43)) and not (inputs(207));
    layer0_outputs(4405) <= not(inputs(0)) or (inputs(111));
    layer0_outputs(4406) <= not((inputs(200)) or (inputs(139)));
    layer0_outputs(4407) <= '0';
    layer0_outputs(4408) <= not((inputs(12)) xor (inputs(234)));
    layer0_outputs(4409) <= inputs(240);
    layer0_outputs(4410) <= (inputs(223)) xor (inputs(220));
    layer0_outputs(4411) <= (inputs(108)) and not (inputs(105));
    layer0_outputs(4412) <= (inputs(77)) or (inputs(104));
    layer0_outputs(4413) <= not((inputs(223)) xor (inputs(234)));
    layer0_outputs(4414) <= not((inputs(112)) xor (inputs(224)));
    layer0_outputs(4415) <= not(inputs(210)) or (inputs(47));
    layer0_outputs(4416) <= inputs(118);
    layer0_outputs(4417) <= inputs(10);
    layer0_outputs(4418) <= '1';
    layer0_outputs(4419) <= inputs(179);
    layer0_outputs(4420) <= not(inputs(113));
    layer0_outputs(4421) <= not((inputs(245)) xor (inputs(136)));
    layer0_outputs(4422) <= (inputs(12)) xor (inputs(50));
    layer0_outputs(4423) <= inputs(114);
    layer0_outputs(4424) <= not((inputs(111)) xor (inputs(204)));
    layer0_outputs(4425) <= not(inputs(149));
    layer0_outputs(4426) <= not((inputs(134)) xor (inputs(100)));
    layer0_outputs(4427) <= (inputs(28)) and not (inputs(187));
    layer0_outputs(4428) <= not(inputs(146));
    layer0_outputs(4429) <= not(inputs(209)) or (inputs(142));
    layer0_outputs(4430) <= '1';
    layer0_outputs(4431) <= (inputs(38)) and not (inputs(13));
    layer0_outputs(4432) <= '0';
    layer0_outputs(4433) <= (inputs(105)) xor (inputs(178));
    layer0_outputs(4434) <= not((inputs(57)) or (inputs(85)));
    layer0_outputs(4435) <= '0';
    layer0_outputs(4436) <= inputs(108);
    layer0_outputs(4437) <= (inputs(204)) xor (inputs(120));
    layer0_outputs(4438) <= not((inputs(215)) or (inputs(51)));
    layer0_outputs(4439) <= not((inputs(107)) or (inputs(221)));
    layer0_outputs(4440) <= not((inputs(180)) xor (inputs(52)));
    layer0_outputs(4441) <= inputs(48);
    layer0_outputs(4442) <= not(inputs(236));
    layer0_outputs(4443) <= not((inputs(9)) xor (inputs(123)));
    layer0_outputs(4444) <= not(inputs(86));
    layer0_outputs(4445) <= (inputs(207)) xor (inputs(115));
    layer0_outputs(4446) <= inputs(6);
    layer0_outputs(4447) <= inputs(125);
    layer0_outputs(4448) <= not(inputs(63)) or (inputs(161));
    layer0_outputs(4449) <= inputs(238);
    layer0_outputs(4450) <= not(inputs(42));
    layer0_outputs(4451) <= inputs(22);
    layer0_outputs(4452) <= not(inputs(29)) or (inputs(109));
    layer0_outputs(4453) <= (inputs(67)) and not (inputs(218));
    layer0_outputs(4454) <= not((inputs(69)) xor (inputs(87)));
    layer0_outputs(4455) <= (inputs(152)) or (inputs(5));
    layer0_outputs(4456) <= not((inputs(159)) or (inputs(119)));
    layer0_outputs(4457) <= not(inputs(102)) or (inputs(194));
    layer0_outputs(4458) <= not((inputs(9)) or (inputs(207)));
    layer0_outputs(4459) <= not((inputs(169)) xor (inputs(201)));
    layer0_outputs(4460) <= inputs(211);
    layer0_outputs(4461) <= not((inputs(13)) xor (inputs(202)));
    layer0_outputs(4462) <= (inputs(142)) or (inputs(100));
    layer0_outputs(4463) <= not(inputs(6)) or (inputs(140));
    layer0_outputs(4464) <= not(inputs(11));
    layer0_outputs(4465) <= not((inputs(36)) or (inputs(30)));
    layer0_outputs(4466) <= (inputs(212)) and not (inputs(147));
    layer0_outputs(4467) <= '0';
    layer0_outputs(4468) <= (inputs(71)) or (inputs(31));
    layer0_outputs(4469) <= inputs(220);
    layer0_outputs(4470) <= (inputs(104)) or (inputs(119));
    layer0_outputs(4471) <= (inputs(218)) or (inputs(177));
    layer0_outputs(4472) <= (inputs(227)) or (inputs(218));
    layer0_outputs(4473) <= inputs(110);
    layer0_outputs(4474) <= (inputs(15)) or (inputs(151));
    layer0_outputs(4475) <= (inputs(198)) and not (inputs(190));
    layer0_outputs(4476) <= (inputs(90)) and not (inputs(14));
    layer0_outputs(4477) <= (inputs(205)) and not (inputs(111));
    layer0_outputs(4478) <= not((inputs(117)) xor (inputs(177)));
    layer0_outputs(4479) <= inputs(135);
    layer0_outputs(4480) <= (inputs(33)) and not (inputs(82));
    layer0_outputs(4481) <= (inputs(45)) and (inputs(113));
    layer0_outputs(4482) <= inputs(49);
    layer0_outputs(4483) <= (inputs(55)) or (inputs(50));
    layer0_outputs(4484) <= not((inputs(71)) xor (inputs(133)));
    layer0_outputs(4485) <= inputs(180);
    layer0_outputs(4486) <= not((inputs(190)) or (inputs(69)));
    layer0_outputs(4487) <= not((inputs(107)) or (inputs(1)));
    layer0_outputs(4488) <= not(inputs(222));
    layer0_outputs(4489) <= not(inputs(228));
    layer0_outputs(4490) <= inputs(41);
    layer0_outputs(4491) <= not(inputs(28)) or (inputs(90));
    layer0_outputs(4492) <= not(inputs(162));
    layer0_outputs(4493) <= inputs(175);
    layer0_outputs(4494) <= (inputs(230)) or (inputs(48));
    layer0_outputs(4495) <= not((inputs(101)) xor (inputs(129)));
    layer0_outputs(4496) <= not(inputs(42)) or (inputs(50));
    layer0_outputs(4497) <= (inputs(157)) xor (inputs(221));
    layer0_outputs(4498) <= (inputs(218)) xor (inputs(104));
    layer0_outputs(4499) <= not((inputs(68)) xor (inputs(142)));
    layer0_outputs(4500) <= (inputs(53)) or (inputs(136));
    layer0_outputs(4501) <= inputs(158);
    layer0_outputs(4502) <= not(inputs(148));
    layer0_outputs(4503) <= (inputs(31)) and not (inputs(243));
    layer0_outputs(4504) <= (inputs(87)) xor (inputs(100));
    layer0_outputs(4505) <= (inputs(85)) or (inputs(100));
    layer0_outputs(4506) <= (inputs(254)) xor (inputs(15));
    layer0_outputs(4507) <= (inputs(165)) and not (inputs(3));
    layer0_outputs(4508) <= inputs(4);
    layer0_outputs(4509) <= (inputs(21)) or (inputs(46));
    layer0_outputs(4510) <= (inputs(69)) and not (inputs(242));
    layer0_outputs(4511) <= inputs(252);
    layer0_outputs(4512) <= not((inputs(109)) or (inputs(133)));
    layer0_outputs(4513) <= not(inputs(217));
    layer0_outputs(4514) <= not(inputs(163));
    layer0_outputs(4515) <= not(inputs(92)) or (inputs(71));
    layer0_outputs(4516) <= (inputs(139)) or (inputs(54));
    layer0_outputs(4517) <= not(inputs(231)) or (inputs(237));
    layer0_outputs(4518) <= not(inputs(201));
    layer0_outputs(4519) <= (inputs(199)) and (inputs(152));
    layer0_outputs(4520) <= not((inputs(75)) or (inputs(109)));
    layer0_outputs(4521) <= not(inputs(27));
    layer0_outputs(4522) <= not(inputs(179)) or (inputs(34));
    layer0_outputs(4523) <= (inputs(88)) or (inputs(82));
    layer0_outputs(4524) <= not((inputs(127)) or (inputs(111)));
    layer0_outputs(4525) <= not((inputs(248)) xor (inputs(201)));
    layer0_outputs(4526) <= (inputs(37)) xor (inputs(95));
    layer0_outputs(4527) <= not(inputs(42));
    layer0_outputs(4528) <= inputs(198);
    layer0_outputs(4529) <= inputs(111);
    layer0_outputs(4530) <= (inputs(148)) xor (inputs(113));
    layer0_outputs(4531) <= not((inputs(25)) xor (inputs(2)));
    layer0_outputs(4532) <= inputs(90);
    layer0_outputs(4533) <= (inputs(150)) or (inputs(165));
    layer0_outputs(4534) <= not((inputs(123)) xor (inputs(15)));
    layer0_outputs(4535) <= inputs(211);
    layer0_outputs(4536) <= not(inputs(94));
    layer0_outputs(4537) <= (inputs(115)) xor (inputs(117));
    layer0_outputs(4538) <= not((inputs(87)) xor (inputs(67)));
    layer0_outputs(4539) <= (inputs(136)) or (inputs(238));
    layer0_outputs(4540) <= inputs(246);
    layer0_outputs(4541) <= inputs(202);
    layer0_outputs(4542) <= not(inputs(23)) or (inputs(220));
    layer0_outputs(4543) <= (inputs(110)) or (inputs(104));
    layer0_outputs(4544) <= (inputs(150)) xor (inputs(252));
    layer0_outputs(4545) <= inputs(181);
    layer0_outputs(4546) <= not((inputs(132)) xor (inputs(194)));
    layer0_outputs(4547) <= not(inputs(102));
    layer0_outputs(4548) <= inputs(13);
    layer0_outputs(4549) <= inputs(99);
    layer0_outputs(4550) <= (inputs(91)) xor (inputs(126));
    layer0_outputs(4551) <= (inputs(149)) or (inputs(134));
    layer0_outputs(4552) <= not((inputs(35)) or (inputs(20)));
    layer0_outputs(4553) <= not(inputs(101));
    layer0_outputs(4554) <= not(inputs(207)) or (inputs(234));
    layer0_outputs(4555) <= (inputs(112)) or (inputs(147));
    layer0_outputs(4556) <= (inputs(177)) xor (inputs(41));
    layer0_outputs(4557) <= not((inputs(201)) xor (inputs(94)));
    layer0_outputs(4558) <= (inputs(175)) xor (inputs(229));
    layer0_outputs(4559) <= inputs(164);
    layer0_outputs(4560) <= (inputs(238)) or (inputs(211));
    layer0_outputs(4561) <= not(inputs(18));
    layer0_outputs(4562) <= not(inputs(183));
    layer0_outputs(4563) <= not((inputs(166)) and (inputs(131)));
    layer0_outputs(4564) <= not(inputs(250));
    layer0_outputs(4565) <= not((inputs(75)) and (inputs(155)));
    layer0_outputs(4566) <= (inputs(35)) xor (inputs(54));
    layer0_outputs(4567) <= '1';
    layer0_outputs(4568) <= (inputs(150)) and not (inputs(83));
    layer0_outputs(4569) <= not(inputs(14));
    layer0_outputs(4570) <= not((inputs(62)) or (inputs(170)));
    layer0_outputs(4571) <= inputs(93);
    layer0_outputs(4572) <= (inputs(18)) or (inputs(160));
    layer0_outputs(4573) <= not(inputs(169)) or (inputs(208));
    layer0_outputs(4574) <= (inputs(178)) or (inputs(174));
    layer0_outputs(4575) <= (inputs(41)) or (inputs(210));
    layer0_outputs(4576) <= (inputs(241)) and not (inputs(19));
    layer0_outputs(4577) <= '1';
    layer0_outputs(4578) <= inputs(4);
    layer0_outputs(4579) <= (inputs(192)) xor (inputs(167));
    layer0_outputs(4580) <= not((inputs(197)) xor (inputs(149)));
    layer0_outputs(4581) <= not((inputs(188)) or (inputs(252)));
    layer0_outputs(4582) <= (inputs(132)) and not (inputs(0));
    layer0_outputs(4583) <= (inputs(44)) and not (inputs(120));
    layer0_outputs(4584) <= not((inputs(79)) or (inputs(55)));
    layer0_outputs(4585) <= not((inputs(140)) xor (inputs(207)));
    layer0_outputs(4586) <= (inputs(148)) xor (inputs(52));
    layer0_outputs(4587) <= inputs(32);
    layer0_outputs(4588) <= (inputs(204)) and not (inputs(47));
    layer0_outputs(4589) <= not(inputs(122));
    layer0_outputs(4590) <= not(inputs(103)) or (inputs(21));
    layer0_outputs(4591) <= inputs(234);
    layer0_outputs(4592) <= (inputs(115)) xor (inputs(34));
    layer0_outputs(4593) <= not(inputs(153));
    layer0_outputs(4594) <= (inputs(53)) xor (inputs(249));
    layer0_outputs(4595) <= not(inputs(51)) or (inputs(225));
    layer0_outputs(4596) <= (inputs(154)) and not (inputs(210));
    layer0_outputs(4597) <= inputs(108);
    layer0_outputs(4598) <= (inputs(234)) or (inputs(178));
    layer0_outputs(4599) <= (inputs(92)) and not (inputs(67));
    layer0_outputs(4600) <= inputs(245);
    layer0_outputs(4601) <= inputs(171);
    layer0_outputs(4602) <= not((inputs(135)) and (inputs(36)));
    layer0_outputs(4603) <= (inputs(192)) xor (inputs(65));
    layer0_outputs(4604) <= not((inputs(157)) and (inputs(138)));
    layer0_outputs(4605) <= not(inputs(119));
    layer0_outputs(4606) <= not((inputs(198)) xor (inputs(18)));
    layer0_outputs(4607) <= not(inputs(191));
    layer0_outputs(4608) <= not(inputs(142));
    layer0_outputs(4609) <= not((inputs(202)) xor (inputs(47)));
    layer0_outputs(4610) <= (inputs(89)) and not (inputs(189));
    layer0_outputs(4611) <= (inputs(182)) and (inputs(136));
    layer0_outputs(4612) <= inputs(238);
    layer0_outputs(4613) <= (inputs(59)) xor (inputs(120));
    layer0_outputs(4614) <= inputs(66);
    layer0_outputs(4615) <= inputs(129);
    layer0_outputs(4616) <= inputs(251);
    layer0_outputs(4617) <= not(inputs(139));
    layer0_outputs(4618) <= not(inputs(50)) or (inputs(104));
    layer0_outputs(4619) <= not(inputs(151)) or (inputs(159));
    layer0_outputs(4620) <= not(inputs(21));
    layer0_outputs(4621) <= inputs(119);
    layer0_outputs(4622) <= not((inputs(74)) or (inputs(17)));
    layer0_outputs(4623) <= not(inputs(162));
    layer0_outputs(4624) <= inputs(21);
    layer0_outputs(4625) <= not(inputs(214)) or (inputs(22));
    layer0_outputs(4626) <= not(inputs(82));
    layer0_outputs(4627) <= (inputs(170)) xor (inputs(116));
    layer0_outputs(4628) <= (inputs(248)) and not (inputs(137));
    layer0_outputs(4629) <= (inputs(164)) and not (inputs(31));
    layer0_outputs(4630) <= (inputs(197)) or (inputs(90));
    layer0_outputs(4631) <= (inputs(228)) xor (inputs(189));
    layer0_outputs(4632) <= (inputs(150)) or (inputs(47));
    layer0_outputs(4633) <= (inputs(22)) and not (inputs(97));
    layer0_outputs(4634) <= not(inputs(28));
    layer0_outputs(4635) <= inputs(178);
    layer0_outputs(4636) <= (inputs(135)) xor (inputs(51));
    layer0_outputs(4637) <= inputs(235);
    layer0_outputs(4638) <= not(inputs(84));
    layer0_outputs(4639) <= not((inputs(239)) and (inputs(144)));
    layer0_outputs(4640) <= not((inputs(193)) xor (inputs(213)));
    layer0_outputs(4641) <= inputs(49);
    layer0_outputs(4642) <= not(inputs(43));
    layer0_outputs(4643) <= (inputs(137)) and not (inputs(225));
    layer0_outputs(4644) <= not(inputs(49));
    layer0_outputs(4645) <= not(inputs(165));
    layer0_outputs(4646) <= not((inputs(221)) xor (inputs(38)));
    layer0_outputs(4647) <= not(inputs(183));
    layer0_outputs(4648) <= (inputs(111)) and (inputs(225));
    layer0_outputs(4649) <= not((inputs(162)) or (inputs(238)));
    layer0_outputs(4650) <= inputs(156);
    layer0_outputs(4651) <= not((inputs(102)) and (inputs(89)));
    layer0_outputs(4652) <= inputs(86);
    layer0_outputs(4653) <= (inputs(22)) and not (inputs(30));
    layer0_outputs(4654) <= inputs(236);
    layer0_outputs(4655) <= not((inputs(120)) and (inputs(230)));
    layer0_outputs(4656) <= inputs(75);
    layer0_outputs(4657) <= not(inputs(100)) or (inputs(62));
    layer0_outputs(4658) <= inputs(153);
    layer0_outputs(4659) <= not((inputs(158)) xor (inputs(139)));
    layer0_outputs(4660) <= (inputs(143)) and (inputs(125));
    layer0_outputs(4661) <= not((inputs(156)) or (inputs(228)));
    layer0_outputs(4662) <= (inputs(160)) and not (inputs(186));
    layer0_outputs(4663) <= '0';
    layer0_outputs(4664) <= not((inputs(177)) xor (inputs(190)));
    layer0_outputs(4665) <= inputs(165);
    layer0_outputs(4666) <= (inputs(157)) xor (inputs(33));
    layer0_outputs(4667) <= (inputs(16)) and not (inputs(182));
    layer0_outputs(4668) <= not((inputs(42)) or (inputs(106)));
    layer0_outputs(4669) <= not((inputs(223)) or (inputs(234)));
    layer0_outputs(4670) <= not(inputs(119));
    layer0_outputs(4671) <= not(inputs(61));
    layer0_outputs(4672) <= not((inputs(52)) xor (inputs(208)));
    layer0_outputs(4673) <= not((inputs(143)) or (inputs(249)));
    layer0_outputs(4674) <= (inputs(152)) xor (inputs(202));
    layer0_outputs(4675) <= not((inputs(241)) or (inputs(187)));
    layer0_outputs(4676) <= (inputs(44)) and (inputs(30));
    layer0_outputs(4677) <= not((inputs(129)) or (inputs(83)));
    layer0_outputs(4678) <= (inputs(245)) or (inputs(7));
    layer0_outputs(4679) <= (inputs(237)) xor (inputs(226));
    layer0_outputs(4680) <= not((inputs(23)) xor (inputs(111)));
    layer0_outputs(4681) <= not((inputs(156)) and (inputs(187)));
    layer0_outputs(4682) <= not(inputs(237));
    layer0_outputs(4683) <= not((inputs(142)) xor (inputs(45)));
    layer0_outputs(4684) <= (inputs(50)) and not (inputs(17));
    layer0_outputs(4685) <= (inputs(201)) xor (inputs(248));
    layer0_outputs(4686) <= not(inputs(110)) or (inputs(137));
    layer0_outputs(4687) <= (inputs(16)) xor (inputs(201));
    layer0_outputs(4688) <= (inputs(8)) or (inputs(95));
    layer0_outputs(4689) <= not((inputs(99)) xor (inputs(76)));
    layer0_outputs(4690) <= (inputs(220)) and (inputs(102));
    layer0_outputs(4691) <= not(inputs(68)) or (inputs(165));
    layer0_outputs(4692) <= (inputs(12)) or (inputs(37));
    layer0_outputs(4693) <= not(inputs(120)) or (inputs(80));
    layer0_outputs(4694) <= not((inputs(34)) xor (inputs(4)));
    layer0_outputs(4695) <= (inputs(53)) or (inputs(75));
    layer0_outputs(4696) <= not(inputs(209)) or (inputs(112));
    layer0_outputs(4697) <= (inputs(250)) and (inputs(183));
    layer0_outputs(4698) <= (inputs(118)) xor (inputs(145));
    layer0_outputs(4699) <= inputs(67);
    layer0_outputs(4700) <= inputs(21);
    layer0_outputs(4701) <= inputs(142);
    layer0_outputs(4702) <= (inputs(94)) or (inputs(38));
    layer0_outputs(4703) <= not(inputs(158));
    layer0_outputs(4704) <= not(inputs(104));
    layer0_outputs(4705) <= not(inputs(169));
    layer0_outputs(4706) <= not((inputs(221)) xor (inputs(248)));
    layer0_outputs(4707) <= inputs(98);
    layer0_outputs(4708) <= (inputs(7)) xor (inputs(145));
    layer0_outputs(4709) <= (inputs(199)) and not (inputs(94));
    layer0_outputs(4710) <= not((inputs(218)) or (inputs(172)));
    layer0_outputs(4711) <= (inputs(150)) and not (inputs(83));
    layer0_outputs(4712) <= not((inputs(92)) or (inputs(171)));
    layer0_outputs(4713) <= (inputs(253)) and (inputs(66));
    layer0_outputs(4714) <= (inputs(218)) or (inputs(239));
    layer0_outputs(4715) <= (inputs(203)) or (inputs(10));
    layer0_outputs(4716) <= not((inputs(162)) and (inputs(37)));
    layer0_outputs(4717) <= not((inputs(26)) or (inputs(31)));
    layer0_outputs(4718) <= not(inputs(80));
    layer0_outputs(4719) <= not(inputs(244));
    layer0_outputs(4720) <= (inputs(130)) and not (inputs(175));
    layer0_outputs(4721) <= not(inputs(247));
    layer0_outputs(4722) <= not((inputs(204)) xor (inputs(186)));
    layer0_outputs(4723) <= not((inputs(84)) or (inputs(150)));
    layer0_outputs(4724) <= inputs(43);
    layer0_outputs(4725) <= not((inputs(90)) xor (inputs(104)));
    layer0_outputs(4726) <= (inputs(43)) xor (inputs(130));
    layer0_outputs(4727) <= not((inputs(14)) or (inputs(237)));
    layer0_outputs(4728) <= (inputs(221)) or (inputs(51));
    layer0_outputs(4729) <= not((inputs(161)) xor (inputs(245)));
    layer0_outputs(4730) <= not((inputs(47)) or (inputs(36)));
    layer0_outputs(4731) <= inputs(85);
    layer0_outputs(4732) <= not(inputs(183));
    layer0_outputs(4733) <= inputs(50);
    layer0_outputs(4734) <= (inputs(154)) or (inputs(88));
    layer0_outputs(4735) <= (inputs(197)) or (inputs(142));
    layer0_outputs(4736) <= inputs(232);
    layer0_outputs(4737) <= not(inputs(101)) or (inputs(175));
    layer0_outputs(4738) <= inputs(147);
    layer0_outputs(4739) <= not(inputs(181));
    layer0_outputs(4740) <= (inputs(241)) and (inputs(56));
    layer0_outputs(4741) <= inputs(188);
    layer0_outputs(4742) <= inputs(84);
    layer0_outputs(4743) <= not(inputs(148));
    layer0_outputs(4744) <= not((inputs(249)) or (inputs(210)));
    layer0_outputs(4745) <= (inputs(83)) and not (inputs(63));
    layer0_outputs(4746) <= not((inputs(206)) xor (inputs(211)));
    layer0_outputs(4747) <= not(inputs(43));
    layer0_outputs(4748) <= not(inputs(211));
    layer0_outputs(4749) <= (inputs(195)) and not (inputs(1));
    layer0_outputs(4750) <= not(inputs(24));
    layer0_outputs(4751) <= (inputs(38)) and not (inputs(219));
    layer0_outputs(4752) <= not(inputs(57));
    layer0_outputs(4753) <= not(inputs(178)) or (inputs(31));
    layer0_outputs(4754) <= not(inputs(155)) or (inputs(55));
    layer0_outputs(4755) <= not((inputs(110)) xor (inputs(4)));
    layer0_outputs(4756) <= not(inputs(76)) or (inputs(80));
    layer0_outputs(4757) <= not((inputs(191)) or (inputs(230)));
    layer0_outputs(4758) <= not(inputs(244)) or (inputs(69));
    layer0_outputs(4759) <= not(inputs(31)) or (inputs(139));
    layer0_outputs(4760) <= (inputs(255)) xor (inputs(154));
    layer0_outputs(4761) <= not((inputs(20)) or (inputs(29)));
    layer0_outputs(4762) <= (inputs(150)) or (inputs(118));
    layer0_outputs(4763) <= not((inputs(166)) or (inputs(17)));
    layer0_outputs(4764) <= not((inputs(224)) or (inputs(192)));
    layer0_outputs(4765) <= (inputs(110)) and not (inputs(222));
    layer0_outputs(4766) <= not(inputs(86)) or (inputs(109));
    layer0_outputs(4767) <= not((inputs(243)) or (inputs(2)));
    layer0_outputs(4768) <= not(inputs(198));
    layer0_outputs(4769) <= (inputs(178)) and (inputs(241));
    layer0_outputs(4770) <= (inputs(37)) xor (inputs(79));
    layer0_outputs(4771) <= not(inputs(5));
    layer0_outputs(4772) <= (inputs(124)) xor (inputs(65));
    layer0_outputs(4773) <= not((inputs(9)) xor (inputs(0)));
    layer0_outputs(4774) <= not(inputs(94)) or (inputs(81));
    layer0_outputs(4775) <= not(inputs(120));
    layer0_outputs(4776) <= (inputs(167)) xor (inputs(197));
    layer0_outputs(4777) <= (inputs(61)) xor (inputs(35));
    layer0_outputs(4778) <= (inputs(198)) xor (inputs(84));
    layer0_outputs(4779) <= (inputs(126)) xor (inputs(108));
    layer0_outputs(4780) <= (inputs(186)) and (inputs(147));
    layer0_outputs(4781) <= (inputs(147)) xor (inputs(146));
    layer0_outputs(4782) <= not(inputs(16));
    layer0_outputs(4783) <= (inputs(117)) xor (inputs(133));
    layer0_outputs(4784) <= (inputs(74)) or (inputs(244));
    layer0_outputs(4785) <= not((inputs(165)) xor (inputs(233)));
    layer0_outputs(4786) <= (inputs(62)) and not (inputs(108));
    layer0_outputs(4787) <= not((inputs(195)) xor (inputs(226)));
    layer0_outputs(4788) <= (inputs(229)) xor (inputs(122));
    layer0_outputs(4789) <= inputs(195);
    layer0_outputs(4790) <= inputs(141);
    layer0_outputs(4791) <= (inputs(180)) xor (inputs(145));
    layer0_outputs(4792) <= (inputs(64)) or (inputs(44));
    layer0_outputs(4793) <= (inputs(189)) and not (inputs(43));
    layer0_outputs(4794) <= not((inputs(198)) xor (inputs(208)));
    layer0_outputs(4795) <= not((inputs(164)) or (inputs(149)));
    layer0_outputs(4796) <= inputs(130);
    layer0_outputs(4797) <= not((inputs(35)) or (inputs(142)));
    layer0_outputs(4798) <= not((inputs(230)) or (inputs(162)));
    layer0_outputs(4799) <= not((inputs(233)) or (inputs(0)));
    layer0_outputs(4800) <= not((inputs(96)) or (inputs(147)));
    layer0_outputs(4801) <= inputs(134);
    layer0_outputs(4802) <= (inputs(83)) xor (inputs(54));
    layer0_outputs(4803) <= not(inputs(134)) or (inputs(65));
    layer0_outputs(4804) <= not(inputs(185));
    layer0_outputs(4805) <= (inputs(175)) or (inputs(194));
    layer0_outputs(4806) <= not(inputs(117)) or (inputs(79));
    layer0_outputs(4807) <= not(inputs(232)) or (inputs(119));
    layer0_outputs(4808) <= not(inputs(220));
    layer0_outputs(4809) <= (inputs(212)) and not (inputs(158));
    layer0_outputs(4810) <= (inputs(60)) and not (inputs(160));
    layer0_outputs(4811) <= not((inputs(160)) xor (inputs(16)));
    layer0_outputs(4812) <= inputs(200);
    layer0_outputs(4813) <= (inputs(55)) xor (inputs(200));
    layer0_outputs(4814) <= (inputs(160)) xor (inputs(110));
    layer0_outputs(4815) <= not((inputs(30)) and (inputs(227)));
    layer0_outputs(4816) <= not((inputs(75)) or (inputs(161)));
    layer0_outputs(4817) <= not(inputs(170)) or (inputs(236));
    layer0_outputs(4818) <= inputs(169);
    layer0_outputs(4819) <= (inputs(207)) or (inputs(66));
    layer0_outputs(4820) <= '1';
    layer0_outputs(4821) <= (inputs(75)) and not (inputs(179));
    layer0_outputs(4822) <= not((inputs(55)) or (inputs(111)));
    layer0_outputs(4823) <= inputs(98);
    layer0_outputs(4824) <= (inputs(122)) and (inputs(160));
    layer0_outputs(4825) <= '1';
    layer0_outputs(4826) <= not(inputs(220));
    layer0_outputs(4827) <= not((inputs(96)) xor (inputs(34)));
    layer0_outputs(4828) <= (inputs(252)) xor (inputs(145));
    layer0_outputs(4829) <= not(inputs(85)) or (inputs(0));
    layer0_outputs(4830) <= inputs(220);
    layer0_outputs(4831) <= (inputs(49)) xor (inputs(193));
    layer0_outputs(4832) <= inputs(145);
    layer0_outputs(4833) <= (inputs(227)) and not (inputs(2));
    layer0_outputs(4834) <= not(inputs(242)) or (inputs(244));
    layer0_outputs(4835) <= inputs(40);
    layer0_outputs(4836) <= not(inputs(134)) or (inputs(124));
    layer0_outputs(4837) <= inputs(91);
    layer0_outputs(4838) <= (inputs(44)) and not (inputs(107));
    layer0_outputs(4839) <= (inputs(210)) and not (inputs(94));
    layer0_outputs(4840) <= (inputs(183)) xor (inputs(230));
    layer0_outputs(4841) <= '0';
    layer0_outputs(4842) <= inputs(110);
    layer0_outputs(4843) <= (inputs(231)) xor (inputs(130));
    layer0_outputs(4844) <= (inputs(191)) or (inputs(9));
    layer0_outputs(4845) <= (inputs(253)) or (inputs(48));
    layer0_outputs(4846) <= not((inputs(105)) or (inputs(208)));
    layer0_outputs(4847) <= not((inputs(205)) xor (inputs(155)));
    layer0_outputs(4848) <= (inputs(76)) or (inputs(18));
    layer0_outputs(4849) <= not((inputs(8)) or (inputs(21)));
    layer0_outputs(4850) <= inputs(98);
    layer0_outputs(4851) <= not((inputs(137)) xor (inputs(29)));
    layer0_outputs(4852) <= (inputs(89)) or (inputs(103));
    layer0_outputs(4853) <= not((inputs(145)) xor (inputs(200)));
    layer0_outputs(4854) <= not(inputs(59));
    layer0_outputs(4855) <= inputs(39);
    layer0_outputs(4856) <= '0';
    layer0_outputs(4857) <= not((inputs(38)) and (inputs(228)));
    layer0_outputs(4858) <= not(inputs(74));
    layer0_outputs(4859) <= (inputs(8)) xor (inputs(79));
    layer0_outputs(4860) <= inputs(51);
    layer0_outputs(4861) <= inputs(90);
    layer0_outputs(4862) <= (inputs(12)) and (inputs(225));
    layer0_outputs(4863) <= (inputs(60)) and not (inputs(254));
    layer0_outputs(4864) <= (inputs(43)) or (inputs(107));
    layer0_outputs(4865) <= (inputs(55)) or (inputs(139));
    layer0_outputs(4866) <= not((inputs(211)) or (inputs(52)));
    layer0_outputs(4867) <= (inputs(152)) xor (inputs(214));
    layer0_outputs(4868) <= not(inputs(94)) or (inputs(36));
    layer0_outputs(4869) <= (inputs(189)) and not (inputs(157));
    layer0_outputs(4870) <= (inputs(97)) xor (inputs(149));
    layer0_outputs(4871) <= not((inputs(21)) xor (inputs(175)));
    layer0_outputs(4872) <= (inputs(47)) or (inputs(82));
    layer0_outputs(4873) <= not(inputs(180)) or (inputs(115));
    layer0_outputs(4874) <= not(inputs(163)) or (inputs(33));
    layer0_outputs(4875) <= (inputs(67)) xor (inputs(4));
    layer0_outputs(4876) <= (inputs(42)) xor (inputs(74));
    layer0_outputs(4877) <= (inputs(143)) or (inputs(34));
    layer0_outputs(4878) <= (inputs(227)) xor (inputs(168));
    layer0_outputs(4879) <= (inputs(231)) and not (inputs(141));
    layer0_outputs(4880) <= not(inputs(133));
    layer0_outputs(4881) <= not(inputs(166));
    layer0_outputs(4882) <= not(inputs(84));
    layer0_outputs(4883) <= (inputs(31)) or (inputs(218));
    layer0_outputs(4884) <= (inputs(224)) or (inputs(180));
    layer0_outputs(4885) <= not(inputs(72));
    layer0_outputs(4886) <= not(inputs(57)) or (inputs(66));
    layer0_outputs(4887) <= not((inputs(27)) or (inputs(207)));
    layer0_outputs(4888) <= inputs(122);
    layer0_outputs(4889) <= (inputs(16)) xor (inputs(81));
    layer0_outputs(4890) <= not(inputs(169));
    layer0_outputs(4891) <= (inputs(236)) and not (inputs(96));
    layer0_outputs(4892) <= (inputs(38)) xor (inputs(191));
    layer0_outputs(4893) <= (inputs(53)) xor (inputs(61));
    layer0_outputs(4894) <= not((inputs(95)) xor (inputs(18)));
    layer0_outputs(4895) <= (inputs(102)) xor (inputs(66));
    layer0_outputs(4896) <= not((inputs(208)) xor (inputs(66)));
    layer0_outputs(4897) <= not(inputs(219));
    layer0_outputs(4898) <= (inputs(215)) xor (inputs(232));
    layer0_outputs(4899) <= not(inputs(147));
    layer0_outputs(4900) <= not((inputs(89)) and (inputs(202)));
    layer0_outputs(4901) <= not((inputs(245)) or (inputs(104)));
    layer0_outputs(4902) <= (inputs(196)) xor (inputs(210));
    layer0_outputs(4903) <= not((inputs(34)) xor (inputs(26)));
    layer0_outputs(4904) <= not((inputs(25)) xor (inputs(114)));
    layer0_outputs(4905) <= not(inputs(233));
    layer0_outputs(4906) <= not(inputs(186));
    layer0_outputs(4907) <= inputs(21);
    layer0_outputs(4908) <= (inputs(88)) and not (inputs(234));
    layer0_outputs(4909) <= not(inputs(230)) or (inputs(139));
    layer0_outputs(4910) <= (inputs(107)) or (inputs(63));
    layer0_outputs(4911) <= (inputs(144)) xor (inputs(126));
    layer0_outputs(4912) <= (inputs(58)) xor (inputs(37));
    layer0_outputs(4913) <= (inputs(77)) or (inputs(248));
    layer0_outputs(4914) <= not((inputs(108)) xor (inputs(106)));
    layer0_outputs(4915) <= (inputs(142)) and not (inputs(225));
    layer0_outputs(4916) <= not((inputs(107)) or (inputs(100)));
    layer0_outputs(4917) <= '0';
    layer0_outputs(4918) <= not(inputs(210));
    layer0_outputs(4919) <= inputs(120);
    layer0_outputs(4920) <= not(inputs(198)) or (inputs(13));
    layer0_outputs(4921) <= inputs(76);
    layer0_outputs(4922) <= (inputs(1)) and not (inputs(58));
    layer0_outputs(4923) <= (inputs(251)) xor (inputs(127));
    layer0_outputs(4924) <= '0';
    layer0_outputs(4925) <= inputs(68);
    layer0_outputs(4926) <= not(inputs(234));
    layer0_outputs(4927) <= (inputs(130)) or (inputs(5));
    layer0_outputs(4928) <= inputs(41);
    layer0_outputs(4929) <= not(inputs(217));
    layer0_outputs(4930) <= not(inputs(228));
    layer0_outputs(4931) <= not((inputs(208)) xor (inputs(151)));
    layer0_outputs(4932) <= inputs(99);
    layer0_outputs(4933) <= not((inputs(2)) or (inputs(127)));
    layer0_outputs(4934) <= inputs(57);
    layer0_outputs(4935) <= '1';
    layer0_outputs(4936) <= not(inputs(227)) or (inputs(61));
    layer0_outputs(4937) <= not(inputs(184)) or (inputs(86));
    layer0_outputs(4938) <= (inputs(146)) xor (inputs(171));
    layer0_outputs(4939) <= (inputs(182)) xor (inputs(74));
    layer0_outputs(4940) <= (inputs(251)) and (inputs(244));
    layer0_outputs(4941) <= not(inputs(151)) or (inputs(93));
    layer0_outputs(4942) <= inputs(94);
    layer0_outputs(4943) <= (inputs(77)) and not (inputs(118));
    layer0_outputs(4944) <= (inputs(184)) and not (inputs(26));
    layer0_outputs(4945) <= not((inputs(191)) and (inputs(102)));
    layer0_outputs(4946) <= inputs(197);
    layer0_outputs(4947) <= (inputs(245)) or (inputs(85));
    layer0_outputs(4948) <= inputs(62);
    layer0_outputs(4949) <= not(inputs(41));
    layer0_outputs(4950) <= not(inputs(54)) or (inputs(1));
    layer0_outputs(4951) <= not(inputs(68)) or (inputs(238));
    layer0_outputs(4952) <= (inputs(154)) or (inputs(141));
    layer0_outputs(4953) <= not(inputs(132)) or (inputs(173));
    layer0_outputs(4954) <= (inputs(92)) and not (inputs(2));
    layer0_outputs(4955) <= not((inputs(29)) xor (inputs(237)));
    layer0_outputs(4956) <= not((inputs(50)) or (inputs(158)));
    layer0_outputs(4957) <= inputs(161);
    layer0_outputs(4958) <= (inputs(121)) and not (inputs(18));
    layer0_outputs(4959) <= not((inputs(185)) xor (inputs(250)));
    layer0_outputs(4960) <= not((inputs(244)) or (inputs(24)));
    layer0_outputs(4961) <= inputs(72);
    layer0_outputs(4962) <= not((inputs(11)) or (inputs(204)));
    layer0_outputs(4963) <= inputs(150);
    layer0_outputs(4964) <= inputs(125);
    layer0_outputs(4965) <= not((inputs(57)) xor (inputs(100)));
    layer0_outputs(4966) <= not(inputs(147));
    layer0_outputs(4967) <= (inputs(103)) and not (inputs(253));
    layer0_outputs(4968) <= (inputs(94)) or (inputs(211));
    layer0_outputs(4969) <= not(inputs(141));
    layer0_outputs(4970) <= (inputs(35)) xor (inputs(21));
    layer0_outputs(4971) <= (inputs(81)) or (inputs(228));
    layer0_outputs(4972) <= not((inputs(64)) or (inputs(48)));
    layer0_outputs(4973) <= not((inputs(125)) or (inputs(1)));
    layer0_outputs(4974) <= not(inputs(255)) or (inputs(249));
    layer0_outputs(4975) <= (inputs(219)) and not (inputs(116));
    layer0_outputs(4976) <= not((inputs(5)) or (inputs(188)));
    layer0_outputs(4977) <= (inputs(25)) xor (inputs(209));
    layer0_outputs(4978) <= not(inputs(26)) or (inputs(162));
    layer0_outputs(4979) <= not((inputs(151)) xor (inputs(186)));
    layer0_outputs(4980) <= not(inputs(12)) or (inputs(170));
    layer0_outputs(4981) <= (inputs(61)) and not (inputs(113));
    layer0_outputs(4982) <= not((inputs(44)) xor (inputs(90)));
    layer0_outputs(4983) <= (inputs(14)) xor (inputs(44));
    layer0_outputs(4984) <= not((inputs(199)) or (inputs(184)));
    layer0_outputs(4985) <= (inputs(232)) or (inputs(131));
    layer0_outputs(4986) <= not(inputs(44));
    layer0_outputs(4987) <= (inputs(67)) or (inputs(78));
    layer0_outputs(4988) <= not((inputs(1)) or (inputs(50)));
    layer0_outputs(4989) <= inputs(180);
    layer0_outputs(4990) <= inputs(198);
    layer0_outputs(4991) <= (inputs(46)) or (inputs(78));
    layer0_outputs(4992) <= not((inputs(146)) xor (inputs(46)));
    layer0_outputs(4993) <= (inputs(223)) or (inputs(2));
    layer0_outputs(4994) <= not((inputs(61)) or (inputs(76)));
    layer0_outputs(4995) <= inputs(211);
    layer0_outputs(4996) <= not(inputs(38)) or (inputs(239));
    layer0_outputs(4997) <= not((inputs(173)) xor (inputs(235)));
    layer0_outputs(4998) <= not((inputs(231)) or (inputs(33)));
    layer0_outputs(4999) <= not((inputs(71)) xor (inputs(60)));
    layer0_outputs(5000) <= (inputs(232)) and not (inputs(55));
    layer0_outputs(5001) <= (inputs(10)) and not (inputs(184));
    layer0_outputs(5002) <= (inputs(70)) xor (inputs(231));
    layer0_outputs(5003) <= inputs(226);
    layer0_outputs(5004) <= not(inputs(107));
    layer0_outputs(5005) <= inputs(97);
    layer0_outputs(5006) <= not((inputs(8)) or (inputs(38)));
    layer0_outputs(5007) <= not((inputs(154)) or (inputs(175)));
    layer0_outputs(5008) <= (inputs(151)) xor (inputs(231));
    layer0_outputs(5009) <= not((inputs(252)) or (inputs(161)));
    layer0_outputs(5010) <= not((inputs(160)) xor (inputs(180)));
    layer0_outputs(5011) <= (inputs(149)) and not (inputs(185));
    layer0_outputs(5012) <= (inputs(177)) xor (inputs(107));
    layer0_outputs(5013) <= not(inputs(106));
    layer0_outputs(5014) <= not(inputs(82));
    layer0_outputs(5015) <= not((inputs(10)) or (inputs(84)));
    layer0_outputs(5016) <= inputs(38);
    layer0_outputs(5017) <= (inputs(167)) and not (inputs(235));
    layer0_outputs(5018) <= '0';
    layer0_outputs(5019) <= not(inputs(190));
    layer0_outputs(5020) <= not((inputs(216)) or (inputs(127)));
    layer0_outputs(5021) <= (inputs(39)) or (inputs(251));
    layer0_outputs(5022) <= not(inputs(237)) or (inputs(143));
    layer0_outputs(5023) <= not(inputs(40)) or (inputs(187));
    layer0_outputs(5024) <= not((inputs(194)) or (inputs(24)));
    layer0_outputs(5025) <= not(inputs(133));
    layer0_outputs(5026) <= not(inputs(50)) or (inputs(82));
    layer0_outputs(5027) <= inputs(141);
    layer0_outputs(5028) <= (inputs(28)) xor (inputs(107));
    layer0_outputs(5029) <= not(inputs(214)) or (inputs(93));
    layer0_outputs(5030) <= not(inputs(170)) or (inputs(221));
    layer0_outputs(5031) <= inputs(69);
    layer0_outputs(5032) <= (inputs(131)) and not (inputs(47));
    layer0_outputs(5033) <= (inputs(89)) and not (inputs(48));
    layer0_outputs(5034) <= (inputs(69)) xor (inputs(190));
    layer0_outputs(5035) <= not(inputs(183)) or (inputs(156));
    layer0_outputs(5036) <= not((inputs(63)) or (inputs(64)));
    layer0_outputs(5037) <= (inputs(29)) or (inputs(121));
    layer0_outputs(5038) <= not((inputs(45)) xor (inputs(73)));
    layer0_outputs(5039) <= not(inputs(128)) or (inputs(32));
    layer0_outputs(5040) <= inputs(143);
    layer0_outputs(5041) <= (inputs(244)) or (inputs(4));
    layer0_outputs(5042) <= (inputs(147)) or (inputs(174));
    layer0_outputs(5043) <= inputs(76);
    layer0_outputs(5044) <= not(inputs(102)) or (inputs(55));
    layer0_outputs(5045) <= (inputs(218)) or (inputs(228));
    layer0_outputs(5046) <= (inputs(57)) and (inputs(9));
    layer0_outputs(5047) <= inputs(209);
    layer0_outputs(5048) <= (inputs(150)) or (inputs(236));
    layer0_outputs(5049) <= not((inputs(191)) or (inputs(233)));
    layer0_outputs(5050) <= not((inputs(22)) or (inputs(142)));
    layer0_outputs(5051) <= not((inputs(243)) or (inputs(137)));
    layer0_outputs(5052) <= (inputs(85)) and not (inputs(220));
    layer0_outputs(5053) <= not(inputs(107)) or (inputs(177));
    layer0_outputs(5054) <= (inputs(142)) and (inputs(232));
    layer0_outputs(5055) <= (inputs(82)) and not (inputs(189));
    layer0_outputs(5056) <= (inputs(143)) or (inputs(21));
    layer0_outputs(5057) <= not(inputs(105)) or (inputs(178));
    layer0_outputs(5058) <= not((inputs(95)) xor (inputs(32)));
    layer0_outputs(5059) <= not(inputs(206)) or (inputs(114));
    layer0_outputs(5060) <= (inputs(193)) xor (inputs(151));
    layer0_outputs(5061) <= (inputs(36)) and not (inputs(36));
    layer0_outputs(5062) <= not((inputs(236)) or (inputs(186)));
    layer0_outputs(5063) <= inputs(146);
    layer0_outputs(5064) <= not((inputs(56)) or (inputs(147)));
    layer0_outputs(5065) <= (inputs(171)) and not (inputs(139));
    layer0_outputs(5066) <= (inputs(151)) and not (inputs(46));
    layer0_outputs(5067) <= (inputs(247)) and not (inputs(71));
    layer0_outputs(5068) <= (inputs(69)) and not (inputs(254));
    layer0_outputs(5069) <= not(inputs(232));
    layer0_outputs(5070) <= not((inputs(194)) xor (inputs(117)));
    layer0_outputs(5071) <= not(inputs(146)) or (inputs(192));
    layer0_outputs(5072) <= not((inputs(19)) or (inputs(186)));
    layer0_outputs(5073) <= (inputs(238)) xor (inputs(142));
    layer0_outputs(5074) <= (inputs(249)) xor (inputs(99));
    layer0_outputs(5075) <= not(inputs(179)) or (inputs(185));
    layer0_outputs(5076) <= inputs(228);
    layer0_outputs(5077) <= inputs(134);
    layer0_outputs(5078) <= not(inputs(115));
    layer0_outputs(5079) <= not(inputs(18)) or (inputs(173));
    layer0_outputs(5080) <= (inputs(120)) and not (inputs(110));
    layer0_outputs(5081) <= not(inputs(70));
    layer0_outputs(5082) <= (inputs(101)) or (inputs(163));
    layer0_outputs(5083) <= not(inputs(152));
    layer0_outputs(5084) <= (inputs(151)) and not (inputs(54));
    layer0_outputs(5085) <= not(inputs(82));
    layer0_outputs(5086) <= not((inputs(53)) xor (inputs(86)));
    layer0_outputs(5087) <= '1';
    layer0_outputs(5088) <= not(inputs(45));
    layer0_outputs(5089) <= '0';
    layer0_outputs(5090) <= not(inputs(237));
    layer0_outputs(5091) <= not((inputs(30)) or (inputs(98)));
    layer0_outputs(5092) <= inputs(196);
    layer0_outputs(5093) <= inputs(248);
    layer0_outputs(5094) <= not((inputs(7)) and (inputs(70)));
    layer0_outputs(5095) <= not((inputs(71)) and (inputs(121)));
    layer0_outputs(5096) <= inputs(227);
    layer0_outputs(5097) <= not((inputs(17)) or (inputs(171)));
    layer0_outputs(5098) <= not((inputs(42)) xor (inputs(73)));
    layer0_outputs(5099) <= not((inputs(87)) xor (inputs(107)));
    layer0_outputs(5100) <= not(inputs(168));
    layer0_outputs(5101) <= not((inputs(3)) xor (inputs(86)));
    layer0_outputs(5102) <= (inputs(59)) or (inputs(125));
    layer0_outputs(5103) <= not(inputs(40));
    layer0_outputs(5104) <= (inputs(51)) or (inputs(63));
    layer0_outputs(5105) <= not((inputs(92)) or (inputs(115)));
    layer0_outputs(5106) <= (inputs(178)) xor (inputs(180));
    layer0_outputs(5107) <= (inputs(35)) and (inputs(147));
    layer0_outputs(5108) <= not(inputs(168)) or (inputs(161));
    layer0_outputs(5109) <= not((inputs(167)) or (inputs(202)));
    layer0_outputs(5110) <= not(inputs(61)) or (inputs(222));
    layer0_outputs(5111) <= (inputs(105)) xor (inputs(67));
    layer0_outputs(5112) <= (inputs(245)) or (inputs(144));
    layer0_outputs(5113) <= not(inputs(28)) or (inputs(239));
    layer0_outputs(5114) <= (inputs(158)) xor (inputs(99));
    layer0_outputs(5115) <= not((inputs(193)) or (inputs(133)));
    layer0_outputs(5116) <= not(inputs(106));
    layer0_outputs(5117) <= not(inputs(165));
    layer0_outputs(5118) <= not(inputs(219)) or (inputs(14));
    layer0_outputs(5119) <= inputs(34);
    layer0_outputs(5120) <= not((inputs(65)) and (inputs(0)));
    layer0_outputs(5121) <= not(inputs(54)) or (inputs(190));
    layer0_outputs(5122) <= not(inputs(216));
    layer0_outputs(5123) <= not(inputs(136));
    layer0_outputs(5124) <= (inputs(113)) xor (inputs(51));
    layer0_outputs(5125) <= not(inputs(175));
    layer0_outputs(5126) <= (inputs(196)) xor (inputs(126));
    layer0_outputs(5127) <= inputs(153);
    layer0_outputs(5128) <= inputs(151);
    layer0_outputs(5129) <= not((inputs(177)) or (inputs(174)));
    layer0_outputs(5130) <= not(inputs(228)) or (inputs(59));
    layer0_outputs(5131) <= inputs(124);
    layer0_outputs(5132) <= (inputs(205)) xor (inputs(253));
    layer0_outputs(5133) <= inputs(13);
    layer0_outputs(5134) <= (inputs(24)) or (inputs(78));
    layer0_outputs(5135) <= (inputs(195)) xor (inputs(32));
    layer0_outputs(5136) <= not((inputs(216)) or (inputs(33)));
    layer0_outputs(5137) <= inputs(108);
    layer0_outputs(5138) <= (inputs(98)) and not (inputs(249));
    layer0_outputs(5139) <= not(inputs(169)) or (inputs(213));
    layer0_outputs(5140) <= not((inputs(15)) or (inputs(202)));
    layer0_outputs(5141) <= not(inputs(167));
    layer0_outputs(5142) <= (inputs(38)) xor (inputs(129));
    layer0_outputs(5143) <= (inputs(139)) or (inputs(112));
    layer0_outputs(5144) <= inputs(109);
    layer0_outputs(5145) <= not((inputs(230)) xor (inputs(35)));
    layer0_outputs(5146) <= inputs(190);
    layer0_outputs(5147) <= (inputs(217)) and (inputs(91));
    layer0_outputs(5148) <= not(inputs(98));
    layer0_outputs(5149) <= not(inputs(77));
    layer0_outputs(5150) <= not(inputs(182)) or (inputs(159));
    layer0_outputs(5151) <= not((inputs(62)) xor (inputs(180)));
    layer0_outputs(5152) <= inputs(54);
    layer0_outputs(5153) <= not((inputs(47)) or (inputs(209)));
    layer0_outputs(5154) <= (inputs(37)) and not (inputs(239));
    layer0_outputs(5155) <= not(inputs(76)) or (inputs(126));
    layer0_outputs(5156) <= not((inputs(160)) xor (inputs(253)));
    layer0_outputs(5157) <= (inputs(121)) xor (inputs(206));
    layer0_outputs(5158) <= (inputs(121)) and not (inputs(208));
    layer0_outputs(5159) <= (inputs(79)) or (inputs(227));
    layer0_outputs(5160) <= not((inputs(104)) or (inputs(188)));
    layer0_outputs(5161) <= not(inputs(34)) or (inputs(20));
    layer0_outputs(5162) <= (inputs(231)) and not (inputs(106));
    layer0_outputs(5163) <= not((inputs(146)) or (inputs(252)));
    layer0_outputs(5164) <= (inputs(184)) or (inputs(245));
    layer0_outputs(5165) <= not(inputs(71)) or (inputs(112));
    layer0_outputs(5166) <= not((inputs(95)) xor (inputs(119)));
    layer0_outputs(5167) <= (inputs(183)) and not (inputs(63));
    layer0_outputs(5168) <= not((inputs(224)) or (inputs(87)));
    layer0_outputs(5169) <= inputs(181);
    layer0_outputs(5170) <= not(inputs(224));
    layer0_outputs(5171) <= inputs(101);
    layer0_outputs(5172) <= inputs(252);
    layer0_outputs(5173) <= inputs(166);
    layer0_outputs(5174) <= (inputs(92)) or (inputs(7));
    layer0_outputs(5175) <= '0';
    layer0_outputs(5176) <= (inputs(50)) xor (inputs(113));
    layer0_outputs(5177) <= not((inputs(50)) or (inputs(163)));
    layer0_outputs(5178) <= not((inputs(193)) or (inputs(213)));
    layer0_outputs(5179) <= inputs(173);
    layer0_outputs(5180) <= inputs(250);
    layer0_outputs(5181) <= not(inputs(75));
    layer0_outputs(5182) <= (inputs(247)) or (inputs(79));
    layer0_outputs(5183) <= inputs(49);
    layer0_outputs(5184) <= not(inputs(98));
    layer0_outputs(5185) <= not((inputs(108)) or (inputs(32)));
    layer0_outputs(5186) <= inputs(144);
    layer0_outputs(5187) <= (inputs(153)) and not (inputs(211));
    layer0_outputs(5188) <= not(inputs(26)) or (inputs(254));
    layer0_outputs(5189) <= not(inputs(151));
    layer0_outputs(5190) <= not((inputs(233)) or (inputs(233)));
    layer0_outputs(5191) <= not(inputs(247)) or (inputs(124));
    layer0_outputs(5192) <= (inputs(55)) xor (inputs(24));
    layer0_outputs(5193) <= not(inputs(153));
    layer0_outputs(5194) <= (inputs(29)) xor (inputs(144));
    layer0_outputs(5195) <= (inputs(71)) xor (inputs(100));
    layer0_outputs(5196) <= not(inputs(120));
    layer0_outputs(5197) <= not((inputs(169)) or (inputs(248)));
    layer0_outputs(5198) <= (inputs(60)) xor (inputs(226));
    layer0_outputs(5199) <= not(inputs(121)) or (inputs(143));
    layer0_outputs(5200) <= (inputs(175)) or (inputs(159));
    layer0_outputs(5201) <= (inputs(250)) and not (inputs(1));
    layer0_outputs(5202) <= not(inputs(121));
    layer0_outputs(5203) <= (inputs(127)) or (inputs(204));
    layer0_outputs(5204) <= not(inputs(45)) or (inputs(1));
    layer0_outputs(5205) <= inputs(122);
    layer0_outputs(5206) <= not(inputs(225));
    layer0_outputs(5207) <= not(inputs(42));
    layer0_outputs(5208) <= not((inputs(124)) xor (inputs(240)));
    layer0_outputs(5209) <= (inputs(157)) xor (inputs(210));
    layer0_outputs(5210) <= not(inputs(216)) or (inputs(123));
    layer0_outputs(5211) <= not((inputs(14)) or (inputs(250)));
    layer0_outputs(5212) <= not(inputs(137)) or (inputs(22));
    layer0_outputs(5213) <= inputs(218);
    layer0_outputs(5214) <= (inputs(94)) and not (inputs(97));
    layer0_outputs(5215) <= not(inputs(164)) or (inputs(34));
    layer0_outputs(5216) <= inputs(234);
    layer0_outputs(5217) <= inputs(92);
    layer0_outputs(5218) <= (inputs(77)) or (inputs(127));
    layer0_outputs(5219) <= (inputs(38)) or (inputs(224));
    layer0_outputs(5220) <= inputs(50);
    layer0_outputs(5221) <= not(inputs(91)) or (inputs(208));
    layer0_outputs(5222) <= (inputs(6)) and not (inputs(86));
    layer0_outputs(5223) <= (inputs(113)) or (inputs(177));
    layer0_outputs(5224) <= not(inputs(52)) or (inputs(215));
    layer0_outputs(5225) <= inputs(151);
    layer0_outputs(5226) <= (inputs(217)) and not (inputs(30));
    layer0_outputs(5227) <= not(inputs(39)) or (inputs(104));
    layer0_outputs(5228) <= not((inputs(113)) xor (inputs(218)));
    layer0_outputs(5229) <= not((inputs(246)) or (inputs(226)));
    layer0_outputs(5230) <= not(inputs(99)) or (inputs(3));
    layer0_outputs(5231) <= not((inputs(55)) xor (inputs(29)));
    layer0_outputs(5232) <= not(inputs(31));
    layer0_outputs(5233) <= inputs(165);
    layer0_outputs(5234) <= (inputs(216)) and not (inputs(116));
    layer0_outputs(5235) <= inputs(178);
    layer0_outputs(5236) <= not((inputs(229)) xor (inputs(42)));
    layer0_outputs(5237) <= not(inputs(138));
    layer0_outputs(5238) <= not((inputs(80)) xor (inputs(155)));
    layer0_outputs(5239) <= inputs(167);
    layer0_outputs(5240) <= (inputs(20)) and not (inputs(178));
    layer0_outputs(5241) <= not(inputs(163));
    layer0_outputs(5242) <= (inputs(51)) xor (inputs(241));
    layer0_outputs(5243) <= (inputs(197)) and not (inputs(21));
    layer0_outputs(5244) <= not(inputs(138)) or (inputs(63));
    layer0_outputs(5245) <= (inputs(55)) xor (inputs(66));
    layer0_outputs(5246) <= (inputs(122)) or (inputs(58));
    layer0_outputs(5247) <= not(inputs(211));
    layer0_outputs(5248) <= not((inputs(241)) xor (inputs(195)));
    layer0_outputs(5249) <= not((inputs(188)) xor (inputs(80)));
    layer0_outputs(5250) <= not(inputs(36)) or (inputs(127));
    layer0_outputs(5251) <= not(inputs(162)) or (inputs(125));
    layer0_outputs(5252) <= not(inputs(155)) or (inputs(196));
    layer0_outputs(5253) <= not((inputs(19)) or (inputs(162)));
    layer0_outputs(5254) <= not((inputs(1)) or (inputs(122)));
    layer0_outputs(5255) <= (inputs(6)) or (inputs(2));
    layer0_outputs(5256) <= not(inputs(23));
    layer0_outputs(5257) <= (inputs(4)) xor (inputs(194));
    layer0_outputs(5258) <= not(inputs(59));
    layer0_outputs(5259) <= inputs(28);
    layer0_outputs(5260) <= (inputs(76)) and not (inputs(236));
    layer0_outputs(5261) <= not((inputs(63)) or (inputs(64)));
    layer0_outputs(5262) <= not(inputs(203));
    layer0_outputs(5263) <= not(inputs(179));
    layer0_outputs(5264) <= (inputs(87)) xor (inputs(61));
    layer0_outputs(5265) <= not(inputs(21));
    layer0_outputs(5266) <= (inputs(149)) xor (inputs(0));
    layer0_outputs(5267) <= not(inputs(152));
    layer0_outputs(5268) <= not(inputs(89));
    layer0_outputs(5269) <= not((inputs(197)) or (inputs(1)));
    layer0_outputs(5270) <= not(inputs(164)) or (inputs(255));
    layer0_outputs(5271) <= (inputs(92)) and not (inputs(14));
    layer0_outputs(5272) <= not(inputs(89));
    layer0_outputs(5273) <= not(inputs(193));
    layer0_outputs(5274) <= not(inputs(80)) or (inputs(93));
    layer0_outputs(5275) <= not((inputs(128)) xor (inputs(163)));
    layer0_outputs(5276) <= inputs(136);
    layer0_outputs(5277) <= (inputs(36)) or (inputs(57));
    layer0_outputs(5278) <= not(inputs(35)) or (inputs(145));
    layer0_outputs(5279) <= inputs(89);
    layer0_outputs(5280) <= (inputs(169)) or (inputs(250));
    layer0_outputs(5281) <= not(inputs(228));
    layer0_outputs(5282) <= not((inputs(166)) or (inputs(132)));
    layer0_outputs(5283) <= (inputs(30)) xor (inputs(207));
    layer0_outputs(5284) <= not(inputs(151));
    layer0_outputs(5285) <= inputs(170);
    layer0_outputs(5286) <= inputs(91);
    layer0_outputs(5287) <= not((inputs(13)) or (inputs(54)));
    layer0_outputs(5288) <= (inputs(111)) or (inputs(83));
    layer0_outputs(5289) <= (inputs(72)) and not (inputs(147));
    layer0_outputs(5290) <= not(inputs(200));
    layer0_outputs(5291) <= (inputs(95)) xor (inputs(27));
    layer0_outputs(5292) <= not(inputs(137));
    layer0_outputs(5293) <= inputs(147);
    layer0_outputs(5294) <= not((inputs(132)) or (inputs(16)));
    layer0_outputs(5295) <= not(inputs(72)) or (inputs(32));
    layer0_outputs(5296) <= inputs(68);
    layer0_outputs(5297) <= inputs(28);
    layer0_outputs(5298) <= not(inputs(111));
    layer0_outputs(5299) <= not((inputs(62)) xor (inputs(59)));
    layer0_outputs(5300) <= '1';
    layer0_outputs(5301) <= inputs(244);
    layer0_outputs(5302) <= (inputs(201)) and (inputs(119));
    layer0_outputs(5303) <= (inputs(59)) xor (inputs(89));
    layer0_outputs(5304) <= '1';
    layer0_outputs(5305) <= not((inputs(139)) or (inputs(22)));
    layer0_outputs(5306) <= inputs(19);
    layer0_outputs(5307) <= (inputs(217)) and not (inputs(95));
    layer0_outputs(5308) <= not((inputs(32)) or (inputs(59)));
    layer0_outputs(5309) <= not((inputs(65)) and (inputs(88)));
    layer0_outputs(5310) <= (inputs(78)) or (inputs(101));
    layer0_outputs(5311) <= not(inputs(153));
    layer0_outputs(5312) <= inputs(229);
    layer0_outputs(5313) <= not(inputs(5));
    layer0_outputs(5314) <= not((inputs(155)) xor (inputs(77)));
    layer0_outputs(5315) <= not((inputs(215)) and (inputs(30)));
    layer0_outputs(5316) <= inputs(176);
    layer0_outputs(5317) <= not(inputs(204));
    layer0_outputs(5318) <= (inputs(135)) and not (inputs(116));
    layer0_outputs(5319) <= inputs(142);
    layer0_outputs(5320) <= not((inputs(42)) xor (inputs(179)));
    layer0_outputs(5321) <= not(inputs(48)) or (inputs(78));
    layer0_outputs(5322) <= (inputs(149)) or (inputs(251));
    layer0_outputs(5323) <= inputs(179);
    layer0_outputs(5324) <= not((inputs(114)) or (inputs(21)));
    layer0_outputs(5325) <= (inputs(21)) xor (inputs(142));
    layer0_outputs(5326) <= (inputs(76)) and not (inputs(50));
    layer0_outputs(5327) <= '0';
    layer0_outputs(5328) <= (inputs(135)) and not (inputs(246));
    layer0_outputs(5329) <= (inputs(83)) xor (inputs(39));
    layer0_outputs(5330) <= inputs(100);
    layer0_outputs(5331) <= not(inputs(100));
    layer0_outputs(5332) <= (inputs(55)) or (inputs(65));
    layer0_outputs(5333) <= not(inputs(211));
    layer0_outputs(5334) <= not((inputs(210)) xor (inputs(236)));
    layer0_outputs(5335) <= not((inputs(17)) or (inputs(150)));
    layer0_outputs(5336) <= not(inputs(84));
    layer0_outputs(5337) <= inputs(237);
    layer0_outputs(5338) <= (inputs(76)) and not (inputs(79));
    layer0_outputs(5339) <= not((inputs(49)) or (inputs(77)));
    layer0_outputs(5340) <= not(inputs(29)) or (inputs(227));
    layer0_outputs(5341) <= not(inputs(88)) or (inputs(110));
    layer0_outputs(5342) <= '0';
    layer0_outputs(5343) <= not(inputs(89));
    layer0_outputs(5344) <= (inputs(115)) xor (inputs(177));
    layer0_outputs(5345) <= not((inputs(83)) xor (inputs(87)));
    layer0_outputs(5346) <= not(inputs(104));
    layer0_outputs(5347) <= (inputs(149)) xor (inputs(212));
    layer0_outputs(5348) <= not((inputs(225)) and (inputs(21)));
    layer0_outputs(5349) <= (inputs(66)) and not (inputs(117));
    layer0_outputs(5350) <= not(inputs(43));
    layer0_outputs(5351) <= (inputs(197)) or (inputs(189));
    layer0_outputs(5352) <= not(inputs(97));
    layer0_outputs(5353) <= (inputs(231)) and not (inputs(66));
    layer0_outputs(5354) <= not((inputs(166)) or (inputs(238)));
    layer0_outputs(5355) <= not(inputs(203));
    layer0_outputs(5356) <= (inputs(43)) xor (inputs(75));
    layer0_outputs(5357) <= (inputs(156)) and (inputs(126));
    layer0_outputs(5358) <= not((inputs(155)) xor (inputs(13)));
    layer0_outputs(5359) <= inputs(230);
    layer0_outputs(5360) <= not(inputs(193));
    layer0_outputs(5361) <= not((inputs(220)) or (inputs(120)));
    layer0_outputs(5362) <= inputs(45);
    layer0_outputs(5363) <= inputs(215);
    layer0_outputs(5364) <= not(inputs(251));
    layer0_outputs(5365) <= (inputs(17)) or (inputs(238));
    layer0_outputs(5366) <= not(inputs(2));
    layer0_outputs(5367) <= not((inputs(226)) xor (inputs(53)));
    layer0_outputs(5368) <= not(inputs(157)) or (inputs(112));
    layer0_outputs(5369) <= (inputs(90)) xor (inputs(6));
    layer0_outputs(5370) <= (inputs(213)) and not (inputs(129));
    layer0_outputs(5371) <= (inputs(57)) xor (inputs(30));
    layer0_outputs(5372) <= inputs(58);
    layer0_outputs(5373) <= inputs(6);
    layer0_outputs(5374) <= not((inputs(0)) or (inputs(211)));
    layer0_outputs(5375) <= (inputs(138)) xor (inputs(74));
    layer0_outputs(5376) <= '0';
    layer0_outputs(5377) <= not((inputs(215)) or (inputs(47)));
    layer0_outputs(5378) <= (inputs(188)) and (inputs(122));
    layer0_outputs(5379) <= not((inputs(193)) and (inputs(185)));
    layer0_outputs(5380) <= not(inputs(71));
    layer0_outputs(5381) <= (inputs(181)) and not (inputs(5));
    layer0_outputs(5382) <= not(inputs(52)) or (inputs(145));
    layer0_outputs(5383) <= (inputs(236)) and not (inputs(209));
    layer0_outputs(5384) <= not(inputs(106));
    layer0_outputs(5385) <= (inputs(228)) or (inputs(213));
    layer0_outputs(5386) <= inputs(123);
    layer0_outputs(5387) <= (inputs(89)) and not (inputs(142));
    layer0_outputs(5388) <= not((inputs(203)) xor (inputs(6)));
    layer0_outputs(5389) <= (inputs(183)) xor (inputs(16));
    layer0_outputs(5390) <= not((inputs(153)) and (inputs(90)));
    layer0_outputs(5391) <= not(inputs(56)) or (inputs(205));
    layer0_outputs(5392) <= not((inputs(140)) xor (inputs(46)));
    layer0_outputs(5393) <= (inputs(198)) xor (inputs(11));
    layer0_outputs(5394) <= not((inputs(222)) xor (inputs(89)));
    layer0_outputs(5395) <= not((inputs(191)) or (inputs(7)));
    layer0_outputs(5396) <= (inputs(103)) and not (inputs(165));
    layer0_outputs(5397) <= not((inputs(2)) or (inputs(212)));
    layer0_outputs(5398) <= not(inputs(197)) or (inputs(92));
    layer0_outputs(5399) <= (inputs(101)) and not (inputs(118));
    layer0_outputs(5400) <= not((inputs(244)) xor (inputs(166)));
    layer0_outputs(5401) <= not(inputs(70)) or (inputs(169));
    layer0_outputs(5402) <= not(inputs(116)) or (inputs(240));
    layer0_outputs(5403) <= not((inputs(156)) xor (inputs(246)));
    layer0_outputs(5404) <= not(inputs(10));
    layer0_outputs(5405) <= (inputs(252)) and not (inputs(192));
    layer0_outputs(5406) <= inputs(105);
    layer0_outputs(5407) <= not(inputs(135)) or (inputs(49));
    layer0_outputs(5408) <= (inputs(42)) xor (inputs(49));
    layer0_outputs(5409) <= inputs(118);
    layer0_outputs(5410) <= (inputs(227)) and not (inputs(202));
    layer0_outputs(5411) <= (inputs(226)) xor (inputs(68));
    layer0_outputs(5412) <= not(inputs(172));
    layer0_outputs(5413) <= inputs(62);
    layer0_outputs(5414) <= '1';
    layer0_outputs(5415) <= '0';
    layer0_outputs(5416) <= (inputs(225)) or (inputs(33));
    layer0_outputs(5417) <= (inputs(131)) xor (inputs(25));
    layer0_outputs(5418) <= (inputs(113)) xor (inputs(235));
    layer0_outputs(5419) <= not(inputs(9));
    layer0_outputs(5420) <= inputs(21);
    layer0_outputs(5421) <= not((inputs(122)) or (inputs(1)));
    layer0_outputs(5422) <= not((inputs(92)) xor (inputs(240)));
    layer0_outputs(5423) <= not(inputs(22)) or (inputs(199));
    layer0_outputs(5424) <= not(inputs(213));
    layer0_outputs(5425) <= inputs(21);
    layer0_outputs(5426) <= not(inputs(163));
    layer0_outputs(5427) <= inputs(53);
    layer0_outputs(5428) <= not(inputs(22));
    layer0_outputs(5429) <= not(inputs(164)) or (inputs(190));
    layer0_outputs(5430) <= not(inputs(43)) or (inputs(178));
    layer0_outputs(5431) <= '1';
    layer0_outputs(5432) <= not(inputs(227));
    layer0_outputs(5433) <= inputs(119);
    layer0_outputs(5434) <= not((inputs(3)) or (inputs(139)));
    layer0_outputs(5435) <= not(inputs(105)) or (inputs(24));
    layer0_outputs(5436) <= (inputs(163)) xor (inputs(181));
    layer0_outputs(5437) <= inputs(15);
    layer0_outputs(5438) <= (inputs(171)) and not (inputs(13));
    layer0_outputs(5439) <= not((inputs(180)) and (inputs(76)));
    layer0_outputs(5440) <= (inputs(143)) and not (inputs(242));
    layer0_outputs(5441) <= not(inputs(234)) or (inputs(2));
    layer0_outputs(5442) <= not((inputs(143)) or (inputs(157)));
    layer0_outputs(5443) <= inputs(44);
    layer0_outputs(5444) <= (inputs(168)) xor (inputs(241));
    layer0_outputs(5445) <= (inputs(43)) xor (inputs(236));
    layer0_outputs(5446) <= not(inputs(146));
    layer0_outputs(5447) <= (inputs(248)) and not (inputs(82));
    layer0_outputs(5448) <= (inputs(22)) or (inputs(106));
    layer0_outputs(5449) <= (inputs(239)) or (inputs(93));
    layer0_outputs(5450) <= not((inputs(235)) xor (inputs(167)));
    layer0_outputs(5451) <= (inputs(132)) or (inputs(200));
    layer0_outputs(5452) <= not(inputs(246)) or (inputs(30));
    layer0_outputs(5453) <= not(inputs(254));
    layer0_outputs(5454) <= (inputs(128)) or (inputs(59));
    layer0_outputs(5455) <= not(inputs(197));
    layer0_outputs(5456) <= not((inputs(202)) xor (inputs(171)));
    layer0_outputs(5457) <= (inputs(82)) or (inputs(205));
    layer0_outputs(5458) <= (inputs(58)) xor (inputs(23));
    layer0_outputs(5459) <= (inputs(255)) and not (inputs(142));
    layer0_outputs(5460) <= (inputs(185)) and not (inputs(79));
    layer0_outputs(5461) <= inputs(198);
    layer0_outputs(5462) <= inputs(66);
    layer0_outputs(5463) <= not((inputs(233)) xor (inputs(168)));
    layer0_outputs(5464) <= (inputs(93)) or (inputs(38));
    layer0_outputs(5465) <= (inputs(165)) xor (inputs(237));
    layer0_outputs(5466) <= not(inputs(248));
    layer0_outputs(5467) <= not(inputs(101)) or (inputs(160));
    layer0_outputs(5468) <= not((inputs(185)) xor (inputs(182)));
    layer0_outputs(5469) <= (inputs(153)) and not (inputs(174));
    layer0_outputs(5470) <= not(inputs(47));
    layer0_outputs(5471) <= (inputs(46)) or (inputs(94));
    layer0_outputs(5472) <= inputs(231);
    layer0_outputs(5473) <= not((inputs(183)) or (inputs(183)));
    layer0_outputs(5474) <= (inputs(111)) xor (inputs(125));
    layer0_outputs(5475) <= inputs(232);
    layer0_outputs(5476) <= not(inputs(100)) or (inputs(166));
    layer0_outputs(5477) <= (inputs(151)) xor (inputs(72));
    layer0_outputs(5478) <= not(inputs(47)) or (inputs(181));
    layer0_outputs(5479) <= not(inputs(106));
    layer0_outputs(5480) <= not(inputs(61));
    layer0_outputs(5481) <= not(inputs(119)) or (inputs(153));
    layer0_outputs(5482) <= (inputs(39)) and (inputs(105));
    layer0_outputs(5483) <= inputs(182);
    layer0_outputs(5484) <= (inputs(59)) and not (inputs(32));
    layer0_outputs(5485) <= not(inputs(228));
    layer0_outputs(5486) <= (inputs(241)) xor (inputs(2));
    layer0_outputs(5487) <= not((inputs(35)) and (inputs(124)));
    layer0_outputs(5488) <= inputs(145);
    layer0_outputs(5489) <= inputs(145);
    layer0_outputs(5490) <= inputs(175);
    layer0_outputs(5491) <= not((inputs(12)) or (inputs(145)));
    layer0_outputs(5492) <= inputs(62);
    layer0_outputs(5493) <= inputs(230);
    layer0_outputs(5494) <= not((inputs(79)) or (inputs(43)));
    layer0_outputs(5495) <= (inputs(179)) and not (inputs(74));
    layer0_outputs(5496) <= (inputs(250)) or (inputs(101));
    layer0_outputs(5497) <= not((inputs(114)) or (inputs(14)));
    layer0_outputs(5498) <= inputs(178);
    layer0_outputs(5499) <= not((inputs(10)) and (inputs(199)));
    layer0_outputs(5500) <= not(inputs(102));
    layer0_outputs(5501) <= (inputs(255)) xor (inputs(90));
    layer0_outputs(5502) <= (inputs(193)) and not (inputs(81));
    layer0_outputs(5503) <= inputs(107);
    layer0_outputs(5504) <= not((inputs(84)) xor (inputs(20)));
    layer0_outputs(5505) <= (inputs(96)) xor (inputs(132));
    layer0_outputs(5506) <= inputs(195);
    layer0_outputs(5507) <= not(inputs(75)) or (inputs(85));
    layer0_outputs(5508) <= (inputs(245)) xor (inputs(173));
    layer0_outputs(5509) <= (inputs(151)) xor (inputs(30));
    layer0_outputs(5510) <= not(inputs(101)) or (inputs(196));
    layer0_outputs(5511) <= (inputs(139)) xor (inputs(254));
    layer0_outputs(5512) <= inputs(60);
    layer0_outputs(5513) <= inputs(53);
    layer0_outputs(5514) <= (inputs(192)) or (inputs(118));
    layer0_outputs(5515) <= not((inputs(117)) xor (inputs(160)));
    layer0_outputs(5516) <= not(inputs(31));
    layer0_outputs(5517) <= (inputs(227)) or (inputs(176));
    layer0_outputs(5518) <= (inputs(112)) or (inputs(143));
    layer0_outputs(5519) <= not((inputs(21)) xor (inputs(67)));
    layer0_outputs(5520) <= not(inputs(207));
    layer0_outputs(5521) <= inputs(55);
    layer0_outputs(5522) <= (inputs(0)) and not (inputs(125));
    layer0_outputs(5523) <= (inputs(154)) and not (inputs(225));
    layer0_outputs(5524) <= (inputs(88)) and not (inputs(33));
    layer0_outputs(5525) <= not(inputs(37));
    layer0_outputs(5526) <= inputs(103);
    layer0_outputs(5527) <= not(inputs(196));
    layer0_outputs(5528) <= inputs(217);
    layer0_outputs(5529) <= not(inputs(89));
    layer0_outputs(5530) <= inputs(68);
    layer0_outputs(5531) <= (inputs(50)) or (inputs(82));
    layer0_outputs(5532) <= inputs(50);
    layer0_outputs(5533) <= not(inputs(162)) or (inputs(15));
    layer0_outputs(5534) <= (inputs(201)) or (inputs(78));
    layer0_outputs(5535) <= (inputs(187)) and not (inputs(216));
    layer0_outputs(5536) <= inputs(198);
    layer0_outputs(5537) <= (inputs(209)) or (inputs(226));
    layer0_outputs(5538) <= inputs(135);
    layer0_outputs(5539) <= (inputs(112)) xor (inputs(69));
    layer0_outputs(5540) <= not(inputs(235));
    layer0_outputs(5541) <= not(inputs(69)) or (inputs(93));
    layer0_outputs(5542) <= not((inputs(30)) xor (inputs(92)));
    layer0_outputs(5543) <= not((inputs(208)) or (inputs(144)));
    layer0_outputs(5544) <= not((inputs(203)) xor (inputs(253)));
    layer0_outputs(5545) <= (inputs(76)) and not (inputs(104));
    layer0_outputs(5546) <= (inputs(219)) and not (inputs(31));
    layer0_outputs(5547) <= '0';
    layer0_outputs(5548) <= inputs(108);
    layer0_outputs(5549) <= inputs(245);
    layer0_outputs(5550) <= not((inputs(238)) and (inputs(175)));
    layer0_outputs(5551) <= inputs(238);
    layer0_outputs(5552) <= not((inputs(56)) or (inputs(191)));
    layer0_outputs(5553) <= not((inputs(195)) or (inputs(248)));
    layer0_outputs(5554) <= not(inputs(188));
    layer0_outputs(5555) <= not(inputs(167)) or (inputs(134));
    layer0_outputs(5556) <= inputs(72);
    layer0_outputs(5557) <= inputs(72);
    layer0_outputs(5558) <= not((inputs(230)) or (inputs(52)));
    layer0_outputs(5559) <= not((inputs(61)) or (inputs(37)));
    layer0_outputs(5560) <= not(inputs(188));
    layer0_outputs(5561) <= (inputs(38)) or (inputs(253));
    layer0_outputs(5562) <= not(inputs(10));
    layer0_outputs(5563) <= (inputs(68)) and not (inputs(131));
    layer0_outputs(5564) <= '1';
    layer0_outputs(5565) <= not(inputs(240));
    layer0_outputs(5566) <= (inputs(238)) xor (inputs(238));
    layer0_outputs(5567) <= (inputs(169)) xor (inputs(13));
    layer0_outputs(5568) <= not((inputs(90)) or (inputs(136)));
    layer0_outputs(5569) <= not((inputs(220)) or (inputs(103)));
    layer0_outputs(5570) <= inputs(111);
    layer0_outputs(5571) <= not((inputs(236)) or (inputs(246)));
    layer0_outputs(5572) <= not(inputs(122)) or (inputs(177));
    layer0_outputs(5573) <= not(inputs(86));
    layer0_outputs(5574) <= (inputs(72)) xor (inputs(41));
    layer0_outputs(5575) <= inputs(79);
    layer0_outputs(5576) <= (inputs(192)) and not (inputs(17));
    layer0_outputs(5577) <= not(inputs(88));
    layer0_outputs(5578) <= not((inputs(223)) xor (inputs(62)));
    layer0_outputs(5579) <= (inputs(21)) or (inputs(68));
    layer0_outputs(5580) <= not(inputs(228));
    layer0_outputs(5581) <= (inputs(160)) xor (inputs(242));
    layer0_outputs(5582) <= (inputs(198)) or (inputs(112));
    layer0_outputs(5583) <= inputs(161);
    layer0_outputs(5584) <= not((inputs(79)) or (inputs(74)));
    layer0_outputs(5585) <= (inputs(54)) xor (inputs(231));
    layer0_outputs(5586) <= inputs(136);
    layer0_outputs(5587) <= not(inputs(50));
    layer0_outputs(5588) <= not(inputs(70)) or (inputs(33));
    layer0_outputs(5589) <= not((inputs(26)) or (inputs(239)));
    layer0_outputs(5590) <= (inputs(55)) and (inputs(38));
    layer0_outputs(5591) <= (inputs(84)) and not (inputs(127));
    layer0_outputs(5592) <= (inputs(131)) or (inputs(67));
    layer0_outputs(5593) <= '1';
    layer0_outputs(5594) <= inputs(121);
    layer0_outputs(5595) <= not((inputs(108)) or (inputs(45)));
    layer0_outputs(5596) <= not(inputs(129));
    layer0_outputs(5597) <= (inputs(211)) and not (inputs(64));
    layer0_outputs(5598) <= (inputs(254)) or (inputs(141));
    layer0_outputs(5599) <= not(inputs(232)) or (inputs(89));
    layer0_outputs(5600) <= not(inputs(90)) or (inputs(181));
    layer0_outputs(5601) <= not(inputs(192)) or (inputs(74));
    layer0_outputs(5602) <= (inputs(116)) or (inputs(246));
    layer0_outputs(5603) <= not(inputs(99)) or (inputs(252));
    layer0_outputs(5604) <= inputs(87);
    layer0_outputs(5605) <= not(inputs(119));
    layer0_outputs(5606) <= inputs(141);
    layer0_outputs(5607) <= not(inputs(49)) or (inputs(34));
    layer0_outputs(5608) <= not((inputs(101)) or (inputs(193)));
    layer0_outputs(5609) <= (inputs(80)) xor (inputs(16));
    layer0_outputs(5610) <= not((inputs(168)) or (inputs(164)));
    layer0_outputs(5611) <= not(inputs(57));
    layer0_outputs(5612) <= not(inputs(179)) or (inputs(15));
    layer0_outputs(5613) <= not((inputs(169)) or (inputs(127)));
    layer0_outputs(5614) <= inputs(26);
    layer0_outputs(5615) <= inputs(235);
    layer0_outputs(5616) <= not((inputs(168)) or (inputs(206)));
    layer0_outputs(5617) <= (inputs(235)) or (inputs(23));
    layer0_outputs(5618) <= not((inputs(223)) xor (inputs(224)));
    layer0_outputs(5619) <= not((inputs(190)) xor (inputs(130)));
    layer0_outputs(5620) <= not((inputs(13)) xor (inputs(60)));
    layer0_outputs(5621) <= (inputs(178)) or (inputs(130));
    layer0_outputs(5622) <= not(inputs(181));
    layer0_outputs(5623) <= inputs(102);
    layer0_outputs(5624) <= not(inputs(235));
    layer0_outputs(5625) <= inputs(88);
    layer0_outputs(5626) <= not((inputs(245)) and (inputs(152)));
    layer0_outputs(5627) <= inputs(111);
    layer0_outputs(5628) <= (inputs(48)) and not (inputs(138));
    layer0_outputs(5629) <= inputs(117);
    layer0_outputs(5630) <= (inputs(234)) and (inputs(217));
    layer0_outputs(5631) <= (inputs(195)) and not (inputs(29));
    layer0_outputs(5632) <= (inputs(73)) and (inputs(165));
    layer0_outputs(5633) <= inputs(62);
    layer0_outputs(5634) <= (inputs(56)) and (inputs(182));
    layer0_outputs(5635) <= inputs(108);
    layer0_outputs(5636) <= (inputs(234)) xor (inputs(185));
    layer0_outputs(5637) <= not(inputs(101));
    layer0_outputs(5638) <= not(inputs(152));
    layer0_outputs(5639) <= (inputs(61)) and (inputs(136));
    layer0_outputs(5640) <= not(inputs(234)) or (inputs(113));
    layer0_outputs(5641) <= not(inputs(227)) or (inputs(33));
    layer0_outputs(5642) <= (inputs(164)) and not (inputs(81));
    layer0_outputs(5643) <= (inputs(202)) and not (inputs(60));
    layer0_outputs(5644) <= (inputs(140)) and not (inputs(45));
    layer0_outputs(5645) <= (inputs(107)) xor (inputs(147));
    layer0_outputs(5646) <= inputs(131);
    layer0_outputs(5647) <= inputs(159);
    layer0_outputs(5648) <= inputs(129);
    layer0_outputs(5649) <= not(inputs(41));
    layer0_outputs(5650) <= not(inputs(243));
    layer0_outputs(5651) <= not(inputs(234));
    layer0_outputs(5652) <= (inputs(233)) or (inputs(181));
    layer0_outputs(5653) <= inputs(12);
    layer0_outputs(5654) <= inputs(24);
    layer0_outputs(5655) <= (inputs(134)) xor (inputs(195));
    layer0_outputs(5656) <= not(inputs(28));
    layer0_outputs(5657) <= not(inputs(85));
    layer0_outputs(5658) <= (inputs(111)) and (inputs(59));
    layer0_outputs(5659) <= not((inputs(229)) xor (inputs(177)));
    layer0_outputs(5660) <= (inputs(193)) xor (inputs(94));
    layer0_outputs(5661) <= (inputs(30)) xor (inputs(190));
    layer0_outputs(5662) <= not((inputs(192)) xor (inputs(168)));
    layer0_outputs(5663) <= (inputs(73)) and not (inputs(65));
    layer0_outputs(5664) <= not(inputs(130)) or (inputs(235));
    layer0_outputs(5665) <= (inputs(169)) and not (inputs(30));
    layer0_outputs(5666) <= not(inputs(108));
    layer0_outputs(5667) <= (inputs(129)) or (inputs(10));
    layer0_outputs(5668) <= not((inputs(225)) or (inputs(4)));
    layer0_outputs(5669) <= not(inputs(105));
    layer0_outputs(5670) <= (inputs(3)) or (inputs(168));
    layer0_outputs(5671) <= inputs(71);
    layer0_outputs(5672) <= not(inputs(234));
    layer0_outputs(5673) <= not((inputs(13)) or (inputs(156)));
    layer0_outputs(5674) <= not(inputs(220)) or (inputs(33));
    layer0_outputs(5675) <= (inputs(24)) and not (inputs(12));
    layer0_outputs(5676) <= (inputs(72)) and not (inputs(223));
    layer0_outputs(5677) <= (inputs(25)) xor (inputs(104));
    layer0_outputs(5678) <= not((inputs(83)) xor (inputs(96)));
    layer0_outputs(5679) <= (inputs(83)) xor (inputs(204));
    layer0_outputs(5680) <= (inputs(31)) and not (inputs(94));
    layer0_outputs(5681) <= inputs(221);
    layer0_outputs(5682) <= (inputs(107)) or (inputs(54));
    layer0_outputs(5683) <= (inputs(229)) and not (inputs(61));
    layer0_outputs(5684) <= not(inputs(188)) or (inputs(16));
    layer0_outputs(5685) <= (inputs(32)) xor (inputs(4));
    layer0_outputs(5686) <= (inputs(171)) xor (inputs(113));
    layer0_outputs(5687) <= (inputs(102)) xor (inputs(149));
    layer0_outputs(5688) <= (inputs(69)) xor (inputs(2));
    layer0_outputs(5689) <= (inputs(93)) or (inputs(253));
    layer0_outputs(5690) <= inputs(99);
    layer0_outputs(5691) <= (inputs(187)) or (inputs(35));
    layer0_outputs(5692) <= (inputs(176)) xor (inputs(186));
    layer0_outputs(5693) <= inputs(114);
    layer0_outputs(5694) <= not(inputs(9));
    layer0_outputs(5695) <= not(inputs(98));
    layer0_outputs(5696) <= inputs(30);
    layer0_outputs(5697) <= not((inputs(157)) or (inputs(115)));
    layer0_outputs(5698) <= inputs(102);
    layer0_outputs(5699) <= not(inputs(118)) or (inputs(96));
    layer0_outputs(5700) <= (inputs(112)) or (inputs(47));
    layer0_outputs(5701) <= not(inputs(216));
    layer0_outputs(5702) <= (inputs(102)) and not (inputs(126));
    layer0_outputs(5703) <= (inputs(58)) and not (inputs(204));
    layer0_outputs(5704) <= not(inputs(15));
    layer0_outputs(5705) <= (inputs(43)) or (inputs(22));
    layer0_outputs(5706) <= inputs(184);
    layer0_outputs(5707) <= not(inputs(164)) or (inputs(97));
    layer0_outputs(5708) <= (inputs(136)) or (inputs(2));
    layer0_outputs(5709) <= not(inputs(26));
    layer0_outputs(5710) <= not(inputs(155));
    layer0_outputs(5711) <= not((inputs(223)) or (inputs(61)));
    layer0_outputs(5712) <= (inputs(238)) or (inputs(132));
    layer0_outputs(5713) <= (inputs(8)) xor (inputs(223));
    layer0_outputs(5714) <= not(inputs(148)) or (inputs(19));
    layer0_outputs(5715) <= not((inputs(42)) or (inputs(217)));
    layer0_outputs(5716) <= (inputs(235)) xor (inputs(188));
    layer0_outputs(5717) <= (inputs(76)) and not (inputs(33));
    layer0_outputs(5718) <= not(inputs(40)) or (inputs(226));
    layer0_outputs(5719) <= (inputs(24)) and not (inputs(66));
    layer0_outputs(5720) <= not(inputs(9));
    layer0_outputs(5721) <= not((inputs(238)) xor (inputs(181)));
    layer0_outputs(5722) <= not((inputs(199)) xor (inputs(215)));
    layer0_outputs(5723) <= (inputs(7)) and not (inputs(126));
    layer0_outputs(5724) <= not((inputs(219)) or (inputs(225)));
    layer0_outputs(5725) <= inputs(198);
    layer0_outputs(5726) <= not(inputs(117));
    layer0_outputs(5727) <= (inputs(207)) xor (inputs(87));
    layer0_outputs(5728) <= not((inputs(65)) xor (inputs(67)));
    layer0_outputs(5729) <= not((inputs(247)) or (inputs(252)));
    layer0_outputs(5730) <= inputs(103);
    layer0_outputs(5731) <= not(inputs(99)) or (inputs(122));
    layer0_outputs(5732) <= not(inputs(214));
    layer0_outputs(5733) <= not((inputs(214)) xor (inputs(249)));
    layer0_outputs(5734) <= not(inputs(62)) or (inputs(98));
    layer0_outputs(5735) <= not(inputs(9)) or (inputs(160));
    layer0_outputs(5736) <= (inputs(54)) or (inputs(94));
    layer0_outputs(5737) <= (inputs(160)) and not (inputs(240));
    layer0_outputs(5738) <= not(inputs(26));
    layer0_outputs(5739) <= (inputs(106)) and (inputs(90));
    layer0_outputs(5740) <= (inputs(116)) or (inputs(226));
    layer0_outputs(5741) <= not((inputs(125)) or (inputs(97)));
    layer0_outputs(5742) <= not(inputs(158));
    layer0_outputs(5743) <= (inputs(155)) xor (inputs(169));
    layer0_outputs(5744) <= not(inputs(212)) or (inputs(73));
    layer0_outputs(5745) <= (inputs(190)) or (inputs(67));
    layer0_outputs(5746) <= (inputs(207)) or (inputs(34));
    layer0_outputs(5747) <= inputs(183);
    layer0_outputs(5748) <= not(inputs(235)) or (inputs(112));
    layer0_outputs(5749) <= (inputs(121)) and (inputs(83));
    layer0_outputs(5750) <= (inputs(35)) or (inputs(31));
    layer0_outputs(5751) <= (inputs(252)) xor (inputs(204));
    layer0_outputs(5752) <= not((inputs(31)) xor (inputs(20)));
    layer0_outputs(5753) <= not((inputs(159)) or (inputs(203)));
    layer0_outputs(5754) <= not((inputs(121)) xor (inputs(14)));
    layer0_outputs(5755) <= (inputs(152)) or (inputs(162));
    layer0_outputs(5756) <= (inputs(140)) or (inputs(201));
    layer0_outputs(5757) <= inputs(82);
    layer0_outputs(5758) <= not((inputs(240)) and (inputs(41)));
    layer0_outputs(5759) <= inputs(165);
    layer0_outputs(5760) <= (inputs(133)) xor (inputs(29));
    layer0_outputs(5761) <= inputs(148);
    layer0_outputs(5762) <= inputs(213);
    layer0_outputs(5763) <= (inputs(109)) xor (inputs(227));
    layer0_outputs(5764) <= (inputs(190)) or (inputs(120));
    layer0_outputs(5765) <= (inputs(217)) and not (inputs(56));
    layer0_outputs(5766) <= (inputs(190)) xor (inputs(193));
    layer0_outputs(5767) <= '0';
    layer0_outputs(5768) <= (inputs(247)) and not (inputs(42));
    layer0_outputs(5769) <= (inputs(191)) or (inputs(243));
    layer0_outputs(5770) <= not((inputs(168)) and (inputs(235)));
    layer0_outputs(5771) <= not(inputs(145));
    layer0_outputs(5772) <= not(inputs(59));
    layer0_outputs(5773) <= (inputs(243)) or (inputs(230));
    layer0_outputs(5774) <= not((inputs(10)) xor (inputs(76)));
    layer0_outputs(5775) <= not(inputs(77)) or (inputs(178));
    layer0_outputs(5776) <= not((inputs(16)) xor (inputs(92)));
    layer0_outputs(5777) <= not((inputs(36)) or (inputs(51)));
    layer0_outputs(5778) <= not((inputs(125)) or (inputs(95)));
    layer0_outputs(5779) <= not(inputs(130)) or (inputs(73));
    layer0_outputs(5780) <= not((inputs(136)) xor (inputs(118)));
    layer0_outputs(5781) <= (inputs(209)) and not (inputs(111));
    layer0_outputs(5782) <= not((inputs(111)) xor (inputs(160)));
    layer0_outputs(5783) <= not((inputs(230)) and (inputs(215)));
    layer0_outputs(5784) <= not((inputs(66)) or (inputs(225)));
    layer0_outputs(5785) <= not((inputs(84)) or (inputs(226)));
    layer0_outputs(5786) <= not(inputs(199)) or (inputs(33));
    layer0_outputs(5787) <= not((inputs(241)) and (inputs(170)));
    layer0_outputs(5788) <= not(inputs(45)) or (inputs(7));
    layer0_outputs(5789) <= inputs(219);
    layer0_outputs(5790) <= (inputs(213)) and not (inputs(97));
    layer0_outputs(5791) <= (inputs(208)) or (inputs(251));
    layer0_outputs(5792) <= not(inputs(106));
    layer0_outputs(5793) <= not((inputs(248)) or (inputs(97)));
    layer0_outputs(5794) <= not((inputs(69)) or (inputs(113)));
    layer0_outputs(5795) <= not(inputs(188));
    layer0_outputs(5796) <= (inputs(34)) and not (inputs(97));
    layer0_outputs(5797) <= not((inputs(139)) xor (inputs(248)));
    layer0_outputs(5798) <= not((inputs(219)) or (inputs(210)));
    layer0_outputs(5799) <= not((inputs(78)) xor (inputs(172)));
    layer0_outputs(5800) <= (inputs(88)) and (inputs(132));
    layer0_outputs(5801) <= not(inputs(11));
    layer0_outputs(5802) <= (inputs(3)) and not (inputs(112));
    layer0_outputs(5803) <= (inputs(250)) and not (inputs(62));
    layer0_outputs(5804) <= not((inputs(115)) xor (inputs(53)));
    layer0_outputs(5805) <= inputs(226);
    layer0_outputs(5806) <= (inputs(254)) or (inputs(76));
    layer0_outputs(5807) <= (inputs(64)) xor (inputs(69));
    layer0_outputs(5808) <= inputs(160);
    layer0_outputs(5809) <= not(inputs(53)) or (inputs(181));
    layer0_outputs(5810) <= not((inputs(113)) or (inputs(25)));
    layer0_outputs(5811) <= not(inputs(214));
    layer0_outputs(5812) <= (inputs(155)) and not (inputs(74));
    layer0_outputs(5813) <= inputs(151);
    layer0_outputs(5814) <= (inputs(228)) and not (inputs(143));
    layer0_outputs(5815) <= (inputs(148)) or (inputs(34));
    layer0_outputs(5816) <= not((inputs(159)) and (inputs(241)));
    layer0_outputs(5817) <= (inputs(170)) or (inputs(236));
    layer0_outputs(5818) <= not((inputs(46)) xor (inputs(215)));
    layer0_outputs(5819) <= not((inputs(114)) or (inputs(62)));
    layer0_outputs(5820) <= not(inputs(83));
    layer0_outputs(5821) <= not(inputs(202)) or (inputs(70));
    layer0_outputs(5822) <= inputs(77);
    layer0_outputs(5823) <= not(inputs(105));
    layer0_outputs(5824) <= not(inputs(172));
    layer0_outputs(5825) <= (inputs(103)) and not (inputs(235));
    layer0_outputs(5826) <= not(inputs(246));
    layer0_outputs(5827) <= inputs(74);
    layer0_outputs(5828) <= not(inputs(187)) or (inputs(18));
    layer0_outputs(5829) <= (inputs(160)) xor (inputs(65));
    layer0_outputs(5830) <= not((inputs(134)) xor (inputs(152)));
    layer0_outputs(5831) <= not((inputs(176)) xor (inputs(49)));
    layer0_outputs(5832) <= not((inputs(231)) or (inputs(242)));
    layer0_outputs(5833) <= not(inputs(91)) or (inputs(204));
    layer0_outputs(5834) <= not(inputs(126));
    layer0_outputs(5835) <= (inputs(211)) and not (inputs(240));
    layer0_outputs(5836) <= not(inputs(195));
    layer0_outputs(5837) <= inputs(255);
    layer0_outputs(5838) <= not(inputs(215));
    layer0_outputs(5839) <= (inputs(102)) or (inputs(19));
    layer0_outputs(5840) <= (inputs(43)) or (inputs(223));
    layer0_outputs(5841) <= not((inputs(25)) and (inputs(162)));
    layer0_outputs(5842) <= (inputs(85)) and not (inputs(174));
    layer0_outputs(5843) <= (inputs(160)) and not (inputs(215));
    layer0_outputs(5844) <= (inputs(158)) xor (inputs(89));
    layer0_outputs(5845) <= not(inputs(204)) or (inputs(66));
    layer0_outputs(5846) <= not(inputs(43)) or (inputs(61));
    layer0_outputs(5847) <= not((inputs(175)) or (inputs(147)));
    layer0_outputs(5848) <= (inputs(109)) or (inputs(252));
    layer0_outputs(5849) <= inputs(118);
    layer0_outputs(5850) <= not((inputs(192)) xor (inputs(172)));
    layer0_outputs(5851) <= not(inputs(136)) or (inputs(144));
    layer0_outputs(5852) <= not((inputs(137)) or (inputs(222)));
    layer0_outputs(5853) <= (inputs(172)) and not (inputs(115));
    layer0_outputs(5854) <= not((inputs(52)) xor (inputs(11)));
    layer0_outputs(5855) <= not((inputs(28)) or (inputs(32)));
    layer0_outputs(5856) <= not(inputs(165));
    layer0_outputs(5857) <= not(inputs(102)) or (inputs(206));
    layer0_outputs(5858) <= not(inputs(9));
    layer0_outputs(5859) <= (inputs(140)) or (inputs(37));
    layer0_outputs(5860) <= (inputs(166)) or (inputs(197));
    layer0_outputs(5861) <= (inputs(30)) and not (inputs(229));
    layer0_outputs(5862) <= (inputs(208)) or (inputs(94));
    layer0_outputs(5863) <= not((inputs(88)) and (inputs(60)));
    layer0_outputs(5864) <= inputs(246);
    layer0_outputs(5865) <= inputs(52);
    layer0_outputs(5866) <= not(inputs(124)) or (inputs(118));
    layer0_outputs(5867) <= (inputs(235)) and not (inputs(110));
    layer0_outputs(5868) <= not((inputs(121)) xor (inputs(206)));
    layer0_outputs(5869) <= (inputs(120)) and not (inputs(177));
    layer0_outputs(5870) <= not((inputs(6)) and (inputs(56)));
    layer0_outputs(5871) <= not((inputs(12)) and (inputs(75)));
    layer0_outputs(5872) <= not(inputs(192)) or (inputs(64));
    layer0_outputs(5873) <= inputs(69);
    layer0_outputs(5874) <= (inputs(233)) and not (inputs(110));
    layer0_outputs(5875) <= (inputs(80)) xor (inputs(195));
    layer0_outputs(5876) <= (inputs(137)) xor (inputs(151));
    layer0_outputs(5877) <= not((inputs(236)) xor (inputs(249)));
    layer0_outputs(5878) <= not(inputs(57)) or (inputs(10));
    layer0_outputs(5879) <= inputs(126);
    layer0_outputs(5880) <= not(inputs(211));
    layer0_outputs(5881) <= (inputs(18)) and not (inputs(156));
    layer0_outputs(5882) <= not(inputs(4));
    layer0_outputs(5883) <= (inputs(193)) and not (inputs(153));
    layer0_outputs(5884) <= not(inputs(91)) or (inputs(226));
    layer0_outputs(5885) <= not(inputs(87));
    layer0_outputs(5886) <= (inputs(149)) and not (inputs(60));
    layer0_outputs(5887) <= not((inputs(59)) or (inputs(49)));
    layer0_outputs(5888) <= inputs(22);
    layer0_outputs(5889) <= not((inputs(50)) or (inputs(252)));
    layer0_outputs(5890) <= not(inputs(58));
    layer0_outputs(5891) <= (inputs(184)) or (inputs(126));
    layer0_outputs(5892) <= not((inputs(68)) xor (inputs(59)));
    layer0_outputs(5893) <= not((inputs(152)) or (inputs(189)));
    layer0_outputs(5894) <= inputs(59);
    layer0_outputs(5895) <= (inputs(92)) and not (inputs(179));
    layer0_outputs(5896) <= (inputs(40)) xor (inputs(127));
    layer0_outputs(5897) <= (inputs(17)) or (inputs(223));
    layer0_outputs(5898) <= not(inputs(229));
    layer0_outputs(5899) <= inputs(224);
    layer0_outputs(5900) <= (inputs(118)) and not (inputs(200));
    layer0_outputs(5901) <= not((inputs(197)) or (inputs(219)));
    layer0_outputs(5902) <= not((inputs(123)) xor (inputs(154)));
    layer0_outputs(5903) <= '1';
    layer0_outputs(5904) <= not(inputs(76));
    layer0_outputs(5905) <= not((inputs(95)) xor (inputs(220)));
    layer0_outputs(5906) <= (inputs(180)) or (inputs(61));
    layer0_outputs(5907) <= not(inputs(61));
    layer0_outputs(5908) <= (inputs(118)) xor (inputs(27));
    layer0_outputs(5909) <= (inputs(79)) xor (inputs(247));
    layer0_outputs(5910) <= (inputs(255)) or (inputs(110));
    layer0_outputs(5911) <= (inputs(152)) xor (inputs(106));
    layer0_outputs(5912) <= not((inputs(77)) xor (inputs(47)));
    layer0_outputs(5913) <= not(inputs(149));
    layer0_outputs(5914) <= not(inputs(122)) or (inputs(7));
    layer0_outputs(5915) <= not(inputs(64));
    layer0_outputs(5916) <= not(inputs(172));
    layer0_outputs(5917) <= (inputs(164)) xor (inputs(153));
    layer0_outputs(5918) <= (inputs(221)) or (inputs(138));
    layer0_outputs(5919) <= (inputs(68)) xor (inputs(31));
    layer0_outputs(5920) <= not(inputs(147));
    layer0_outputs(5921) <= not((inputs(17)) or (inputs(207)));
    layer0_outputs(5922) <= not(inputs(13)) or (inputs(105));
    layer0_outputs(5923) <= not((inputs(58)) xor (inputs(26)));
    layer0_outputs(5924) <= not(inputs(146));
    layer0_outputs(5925) <= not(inputs(44)) or (inputs(190));
    layer0_outputs(5926) <= (inputs(245)) or (inputs(230));
    layer0_outputs(5927) <= (inputs(117)) xor (inputs(184));
    layer0_outputs(5928) <= not((inputs(111)) xor (inputs(67)));
    layer0_outputs(5929) <= (inputs(237)) or (inputs(141));
    layer0_outputs(5930) <= (inputs(98)) xor (inputs(69));
    layer0_outputs(5931) <= (inputs(31)) xor (inputs(176));
    layer0_outputs(5932) <= not((inputs(110)) or (inputs(77)));
    layer0_outputs(5933) <= (inputs(130)) or (inputs(68));
    layer0_outputs(5934) <= not(inputs(97));
    layer0_outputs(5935) <= (inputs(108)) xor (inputs(191));
    layer0_outputs(5936) <= not((inputs(56)) xor (inputs(173)));
    layer0_outputs(5937) <= not((inputs(252)) or (inputs(225)));
    layer0_outputs(5938) <= (inputs(70)) xor (inputs(3));
    layer0_outputs(5939) <= (inputs(161)) and not (inputs(138));
    layer0_outputs(5940) <= inputs(131);
    layer0_outputs(5941) <= (inputs(40)) xor (inputs(247));
    layer0_outputs(5942) <= (inputs(38)) xor (inputs(63));
    layer0_outputs(5943) <= (inputs(245)) and not (inputs(207));
    layer0_outputs(5944) <= not((inputs(220)) or (inputs(255)));
    layer0_outputs(5945) <= (inputs(245)) xor (inputs(34));
    layer0_outputs(5946) <= (inputs(255)) and (inputs(129));
    layer0_outputs(5947) <= not((inputs(108)) xor (inputs(17)));
    layer0_outputs(5948) <= not((inputs(205)) or (inputs(172)));
    layer0_outputs(5949) <= not((inputs(69)) xor (inputs(89)));
    layer0_outputs(5950) <= inputs(150);
    layer0_outputs(5951) <= not((inputs(238)) or (inputs(254)));
    layer0_outputs(5952) <= not(inputs(75));
    layer0_outputs(5953) <= (inputs(126)) xor (inputs(107));
    layer0_outputs(5954) <= not(inputs(198));
    layer0_outputs(5955) <= (inputs(122)) and not (inputs(213));
    layer0_outputs(5956) <= not(inputs(198));
    layer0_outputs(5957) <= (inputs(8)) xor (inputs(61));
    layer0_outputs(5958) <= not(inputs(101)) or (inputs(2));
    layer0_outputs(5959) <= (inputs(169)) and (inputs(156));
    layer0_outputs(5960) <= not((inputs(69)) or (inputs(130)));
    layer0_outputs(5961) <= not((inputs(34)) or (inputs(101)));
    layer0_outputs(5962) <= not(inputs(120)) or (inputs(76));
    layer0_outputs(5963) <= (inputs(178)) and (inputs(146));
    layer0_outputs(5964) <= not(inputs(224));
    layer0_outputs(5965) <= not((inputs(57)) or (inputs(62)));
    layer0_outputs(5966) <= (inputs(74)) and not (inputs(164));
    layer0_outputs(5967) <= (inputs(126)) xor (inputs(222));
    layer0_outputs(5968) <= inputs(76);
    layer0_outputs(5969) <= (inputs(244)) and (inputs(48));
    layer0_outputs(5970) <= (inputs(136)) and (inputs(186));
    layer0_outputs(5971) <= (inputs(254)) and not (inputs(138));
    layer0_outputs(5972) <= (inputs(241)) xor (inputs(218));
    layer0_outputs(5973) <= (inputs(117)) or (inputs(143));
    layer0_outputs(5974) <= not(inputs(122)) or (inputs(227));
    layer0_outputs(5975) <= not((inputs(46)) xor (inputs(225)));
    layer0_outputs(5976) <= not(inputs(91)) or (inputs(219));
    layer0_outputs(5977) <= not((inputs(248)) xor (inputs(215)));
    layer0_outputs(5978) <= not(inputs(138)) or (inputs(243));
    layer0_outputs(5979) <= not((inputs(187)) xor (inputs(186)));
    layer0_outputs(5980) <= (inputs(158)) or (inputs(39));
    layer0_outputs(5981) <= not(inputs(20));
    layer0_outputs(5982) <= not((inputs(229)) and (inputs(11)));
    layer0_outputs(5983) <= inputs(168);
    layer0_outputs(5984) <= inputs(180);
    layer0_outputs(5985) <= (inputs(235)) xor (inputs(211));
    layer0_outputs(5986) <= not(inputs(101));
    layer0_outputs(5987) <= not(inputs(118)) or (inputs(224));
    layer0_outputs(5988) <= inputs(59);
    layer0_outputs(5989) <= not(inputs(114));
    layer0_outputs(5990) <= inputs(126);
    layer0_outputs(5991) <= inputs(247);
    layer0_outputs(5992) <= inputs(167);
    layer0_outputs(5993) <= not((inputs(65)) xor (inputs(87)));
    layer0_outputs(5994) <= not((inputs(242)) or (inputs(69)));
    layer0_outputs(5995) <= '1';
    layer0_outputs(5996) <= (inputs(246)) xor (inputs(199));
    layer0_outputs(5997) <= (inputs(126)) or (inputs(29));
    layer0_outputs(5998) <= (inputs(97)) and (inputs(17));
    layer0_outputs(5999) <= not(inputs(135));
    layer0_outputs(6000) <= (inputs(223)) or (inputs(137));
    layer0_outputs(6001) <= not(inputs(96)) or (inputs(97));
    layer0_outputs(6002) <= not((inputs(163)) or (inputs(214)));
    layer0_outputs(6003) <= (inputs(60)) and not (inputs(79));
    layer0_outputs(6004) <= inputs(193);
    layer0_outputs(6005) <= inputs(177);
    layer0_outputs(6006) <= not(inputs(165));
    layer0_outputs(6007) <= not((inputs(220)) or (inputs(167)));
    layer0_outputs(6008) <= not(inputs(115));
    layer0_outputs(6009) <= not(inputs(86));
    layer0_outputs(6010) <= (inputs(249)) or (inputs(165));
    layer0_outputs(6011) <= (inputs(14)) or (inputs(241));
    layer0_outputs(6012) <= (inputs(159)) and not (inputs(56));
    layer0_outputs(6013) <= not((inputs(6)) and (inputs(63)));
    layer0_outputs(6014) <= (inputs(74)) and not (inputs(239));
    layer0_outputs(6015) <= (inputs(186)) or (inputs(208));
    layer0_outputs(6016) <= (inputs(216)) xor (inputs(194));
    layer0_outputs(6017) <= inputs(194);
    layer0_outputs(6018) <= not((inputs(4)) or (inputs(31)));
    layer0_outputs(6019) <= not((inputs(36)) or (inputs(153)));
    layer0_outputs(6020) <= (inputs(220)) xor (inputs(65));
    layer0_outputs(6021) <= not((inputs(241)) xor (inputs(38)));
    layer0_outputs(6022) <= inputs(142);
    layer0_outputs(6023) <= not(inputs(184)) or (inputs(82));
    layer0_outputs(6024) <= not(inputs(122)) or (inputs(207));
    layer0_outputs(6025) <= not((inputs(34)) or (inputs(166)));
    layer0_outputs(6026) <= inputs(158);
    layer0_outputs(6027) <= inputs(93);
    layer0_outputs(6028) <= not(inputs(76));
    layer0_outputs(6029) <= not(inputs(180)) or (inputs(58));
    layer0_outputs(6030) <= not(inputs(9));
    layer0_outputs(6031) <= (inputs(212)) xor (inputs(217));
    layer0_outputs(6032) <= (inputs(220)) xor (inputs(234));
    layer0_outputs(6033) <= not((inputs(203)) or (inputs(158)));
    layer0_outputs(6034) <= not((inputs(60)) or (inputs(75)));
    layer0_outputs(6035) <= (inputs(99)) and not (inputs(174));
    layer0_outputs(6036) <= (inputs(93)) and not (inputs(237));
    layer0_outputs(6037) <= not(inputs(57));
    layer0_outputs(6038) <= inputs(44);
    layer0_outputs(6039) <= (inputs(176)) or (inputs(14));
    layer0_outputs(6040) <= not(inputs(249)) or (inputs(131));
    layer0_outputs(6041) <= not((inputs(139)) xor (inputs(186)));
    layer0_outputs(6042) <= not((inputs(8)) xor (inputs(57)));
    layer0_outputs(6043) <= not(inputs(238));
    layer0_outputs(6044) <= '1';
    layer0_outputs(6045) <= not((inputs(50)) and (inputs(237)));
    layer0_outputs(6046) <= inputs(201);
    layer0_outputs(6047) <= not((inputs(166)) and (inputs(171)));
    layer0_outputs(6048) <= not((inputs(94)) and (inputs(28)));
    layer0_outputs(6049) <= not(inputs(165));
    layer0_outputs(6050) <= (inputs(6)) or (inputs(79));
    layer0_outputs(6051) <= (inputs(32)) and (inputs(237));
    layer0_outputs(6052) <= not(inputs(230)) or (inputs(15));
    layer0_outputs(6053) <= not(inputs(115)) or (inputs(207));
    layer0_outputs(6054) <= '1';
    layer0_outputs(6055) <= (inputs(238)) and not (inputs(171));
    layer0_outputs(6056) <= (inputs(20)) or (inputs(0));
    layer0_outputs(6057) <= (inputs(128)) or (inputs(99));
    layer0_outputs(6058) <= not((inputs(135)) or (inputs(81)));
    layer0_outputs(6059) <= not(inputs(31)) or (inputs(168));
    layer0_outputs(6060) <= not(inputs(120));
    layer0_outputs(6061) <= inputs(93);
    layer0_outputs(6062) <= (inputs(129)) or (inputs(125));
    layer0_outputs(6063) <= (inputs(206)) or (inputs(75));
    layer0_outputs(6064) <= (inputs(241)) or (inputs(22));
    layer0_outputs(6065) <= inputs(146);
    layer0_outputs(6066) <= not(inputs(77)) or (inputs(134));
    layer0_outputs(6067) <= inputs(176);
    layer0_outputs(6068) <= not((inputs(216)) xor (inputs(180)));
    layer0_outputs(6069) <= not((inputs(110)) or (inputs(166)));
    layer0_outputs(6070) <= not(inputs(73));
    layer0_outputs(6071) <= not(inputs(121)) or (inputs(194));
    layer0_outputs(6072) <= not((inputs(2)) xor (inputs(127)));
    layer0_outputs(6073) <= not((inputs(131)) xor (inputs(164)));
    layer0_outputs(6074) <= not(inputs(184)) or (inputs(123));
    layer0_outputs(6075) <= not((inputs(184)) or (inputs(21)));
    layer0_outputs(6076) <= (inputs(172)) xor (inputs(235));
    layer0_outputs(6077) <= not(inputs(8));
    layer0_outputs(6078) <= (inputs(174)) xor (inputs(228));
    layer0_outputs(6079) <= (inputs(183)) xor (inputs(177));
    layer0_outputs(6080) <= not((inputs(241)) or (inputs(184)));
    layer0_outputs(6081) <= not(inputs(242));
    layer0_outputs(6082) <= (inputs(225)) and not (inputs(238));
    layer0_outputs(6083) <= not(inputs(248));
    layer0_outputs(6084) <= not((inputs(139)) or (inputs(94)));
    layer0_outputs(6085) <= not((inputs(29)) xor (inputs(13)));
    layer0_outputs(6086) <= not(inputs(108));
    layer0_outputs(6087) <= (inputs(19)) or (inputs(203));
    layer0_outputs(6088) <= not(inputs(41)) or (inputs(158));
    layer0_outputs(6089) <= '0';
    layer0_outputs(6090) <= inputs(22);
    layer0_outputs(6091) <= (inputs(71)) or (inputs(160));
    layer0_outputs(6092) <= inputs(107);
    layer0_outputs(6093) <= not(inputs(86));
    layer0_outputs(6094) <= inputs(12);
    layer0_outputs(6095) <= (inputs(94)) and not (inputs(254));
    layer0_outputs(6096) <= not(inputs(242)) or (inputs(130));
    layer0_outputs(6097) <= (inputs(105)) and not (inputs(189));
    layer0_outputs(6098) <= not((inputs(237)) or (inputs(244)));
    layer0_outputs(6099) <= (inputs(34)) xor (inputs(6));
    layer0_outputs(6100) <= not((inputs(116)) xor (inputs(70)));
    layer0_outputs(6101) <= inputs(103);
    layer0_outputs(6102) <= not((inputs(232)) xor (inputs(144)));
    layer0_outputs(6103) <= (inputs(60)) xor (inputs(58));
    layer0_outputs(6104) <= not(inputs(18));
    layer0_outputs(6105) <= not((inputs(69)) or (inputs(238)));
    layer0_outputs(6106) <= (inputs(140)) xor (inputs(41));
    layer0_outputs(6107) <= inputs(40);
    layer0_outputs(6108) <= (inputs(56)) and not (inputs(72));
    layer0_outputs(6109) <= inputs(166);
    layer0_outputs(6110) <= not(inputs(74));
    layer0_outputs(6111) <= (inputs(154)) or (inputs(247));
    layer0_outputs(6112) <= (inputs(183)) xor (inputs(119));
    layer0_outputs(6113) <= not((inputs(124)) xor (inputs(74)));
    layer0_outputs(6114) <= (inputs(14)) or (inputs(243));
    layer0_outputs(6115) <= (inputs(24)) and not (inputs(162));
    layer0_outputs(6116) <= not(inputs(59)) or (inputs(32));
    layer0_outputs(6117) <= (inputs(105)) and (inputs(146));
    layer0_outputs(6118) <= not(inputs(70));
    layer0_outputs(6119) <= (inputs(133)) and not (inputs(186));
    layer0_outputs(6120) <= not(inputs(7)) or (inputs(28));
    layer0_outputs(6121) <= (inputs(70)) or (inputs(4));
    layer0_outputs(6122) <= not((inputs(119)) xor (inputs(38)));
    layer0_outputs(6123) <= not((inputs(173)) or (inputs(145)));
    layer0_outputs(6124) <= (inputs(181)) and (inputs(181));
    layer0_outputs(6125) <= not((inputs(250)) or (inputs(5)));
    layer0_outputs(6126) <= (inputs(139)) or (inputs(75));
    layer0_outputs(6127) <= inputs(232);
    layer0_outputs(6128) <= not(inputs(194));
    layer0_outputs(6129) <= inputs(9);
    layer0_outputs(6130) <= not(inputs(217));
    layer0_outputs(6131) <= (inputs(251)) xor (inputs(36));
    layer0_outputs(6132) <= (inputs(165)) or (inputs(198));
    layer0_outputs(6133) <= not((inputs(63)) or (inputs(247)));
    layer0_outputs(6134) <= inputs(172);
    layer0_outputs(6135) <= not(inputs(250));
    layer0_outputs(6136) <= (inputs(231)) or (inputs(215));
    layer0_outputs(6137) <= (inputs(35)) and not (inputs(4));
    layer0_outputs(6138) <= not(inputs(23));
    layer0_outputs(6139) <= not(inputs(106)) or (inputs(177));
    layer0_outputs(6140) <= not(inputs(103));
    layer0_outputs(6141) <= not(inputs(232)) or (inputs(18));
    layer0_outputs(6142) <= not((inputs(18)) xor (inputs(52)));
    layer0_outputs(6143) <= not(inputs(76));
    layer0_outputs(6144) <= not((inputs(169)) xor (inputs(219)));
    layer0_outputs(6145) <= not(inputs(138)) or (inputs(219));
    layer0_outputs(6146) <= not((inputs(64)) or (inputs(136)));
    layer0_outputs(6147) <= not((inputs(87)) or (inputs(159)));
    layer0_outputs(6148) <= inputs(44);
    layer0_outputs(6149) <= not(inputs(120)) or (inputs(224));
    layer0_outputs(6150) <= not(inputs(127));
    layer0_outputs(6151) <= (inputs(180)) xor (inputs(201));
    layer0_outputs(6152) <= inputs(152);
    layer0_outputs(6153) <= not((inputs(51)) or (inputs(206)));
    layer0_outputs(6154) <= not(inputs(218));
    layer0_outputs(6155) <= not((inputs(79)) or (inputs(106)));
    layer0_outputs(6156) <= not(inputs(220)) or (inputs(143));
    layer0_outputs(6157) <= not(inputs(132)) or (inputs(136));
    layer0_outputs(6158) <= (inputs(92)) xor (inputs(36));
    layer0_outputs(6159) <= not((inputs(123)) xor (inputs(137)));
    layer0_outputs(6160) <= inputs(247);
    layer0_outputs(6161) <= (inputs(207)) xor (inputs(31));
    layer0_outputs(6162) <= (inputs(115)) and (inputs(135));
    layer0_outputs(6163) <= (inputs(199)) and not (inputs(118));
    layer0_outputs(6164) <= inputs(101);
    layer0_outputs(6165) <= (inputs(77)) or (inputs(211));
    layer0_outputs(6166) <= (inputs(208)) xor (inputs(249));
    layer0_outputs(6167) <= '0';
    layer0_outputs(6168) <= (inputs(19)) xor (inputs(109));
    layer0_outputs(6169) <= inputs(40);
    layer0_outputs(6170) <= not((inputs(245)) xor (inputs(20)));
    layer0_outputs(6171) <= inputs(230);
    layer0_outputs(6172) <= (inputs(100)) xor (inputs(108));
    layer0_outputs(6173) <= (inputs(167)) xor (inputs(58));
    layer0_outputs(6174) <= not(inputs(118));
    layer0_outputs(6175) <= inputs(132);
    layer0_outputs(6176) <= not(inputs(211)) or (inputs(112));
    layer0_outputs(6177) <= not((inputs(57)) or (inputs(167)));
    layer0_outputs(6178) <= (inputs(152)) xor (inputs(93));
    layer0_outputs(6179) <= not(inputs(82)) or (inputs(49));
    layer0_outputs(6180) <= (inputs(41)) and (inputs(247));
    layer0_outputs(6181) <= (inputs(62)) or (inputs(47));
    layer0_outputs(6182) <= (inputs(125)) xor (inputs(124));
    layer0_outputs(6183) <= inputs(58);
    layer0_outputs(6184) <= not((inputs(233)) xor (inputs(209)));
    layer0_outputs(6185) <= not((inputs(244)) xor (inputs(33)));
    layer0_outputs(6186) <= (inputs(38)) and not (inputs(177));
    layer0_outputs(6187) <= not((inputs(175)) xor (inputs(207)));
    layer0_outputs(6188) <= (inputs(241)) xor (inputs(137));
    layer0_outputs(6189) <= (inputs(79)) and not (inputs(138));
    layer0_outputs(6190) <= not((inputs(1)) and (inputs(203)));
    layer0_outputs(6191) <= (inputs(56)) and not (inputs(49));
    layer0_outputs(6192) <= (inputs(129)) xor (inputs(179));
    layer0_outputs(6193) <= not((inputs(103)) and (inputs(119)));
    layer0_outputs(6194) <= (inputs(75)) or (inputs(33));
    layer0_outputs(6195) <= not(inputs(163)) or (inputs(124));
    layer0_outputs(6196) <= inputs(39);
    layer0_outputs(6197) <= (inputs(176)) xor (inputs(180));
    layer0_outputs(6198) <= inputs(189);
    layer0_outputs(6199) <= not(inputs(66)) or (inputs(231));
    layer0_outputs(6200) <= '1';
    layer0_outputs(6201) <= not((inputs(126)) xor (inputs(104)));
    layer0_outputs(6202) <= '0';
    layer0_outputs(6203) <= (inputs(244)) and not (inputs(1));
    layer0_outputs(6204) <= (inputs(64)) and not (inputs(174));
    layer0_outputs(6205) <= (inputs(211)) or (inputs(35));
    layer0_outputs(6206) <= inputs(128);
    layer0_outputs(6207) <= inputs(237);
    layer0_outputs(6208) <= not(inputs(128));
    layer0_outputs(6209) <= (inputs(81)) xor (inputs(25));
    layer0_outputs(6210) <= not(inputs(146));
    layer0_outputs(6211) <= (inputs(91)) and not (inputs(4));
    layer0_outputs(6212) <= inputs(60);
    layer0_outputs(6213) <= not(inputs(151));
    layer0_outputs(6214) <= not((inputs(220)) xor (inputs(188)));
    layer0_outputs(6215) <= inputs(228);
    layer0_outputs(6216) <= not((inputs(108)) or (inputs(210)));
    layer0_outputs(6217) <= inputs(222);
    layer0_outputs(6218) <= not(inputs(203));
    layer0_outputs(6219) <= (inputs(40)) or (inputs(128));
    layer0_outputs(6220) <= (inputs(157)) or (inputs(112));
    layer0_outputs(6221) <= (inputs(50)) or (inputs(60));
    layer0_outputs(6222) <= not(inputs(50));
    layer0_outputs(6223) <= not((inputs(225)) and (inputs(175)));
    layer0_outputs(6224) <= (inputs(115)) xor (inputs(87));
    layer0_outputs(6225) <= inputs(107);
    layer0_outputs(6226) <= (inputs(251)) and not (inputs(63));
    layer0_outputs(6227) <= not(inputs(248)) or (inputs(130));
    layer0_outputs(6228) <= not((inputs(89)) xor (inputs(72)));
    layer0_outputs(6229) <= (inputs(211)) and (inputs(216));
    layer0_outputs(6230) <= not(inputs(38));
    layer0_outputs(6231) <= (inputs(30)) xor (inputs(140));
    layer0_outputs(6232) <= not((inputs(128)) xor (inputs(211)));
    layer0_outputs(6233) <= (inputs(182)) or (inputs(0));
    layer0_outputs(6234) <= not(inputs(32));
    layer0_outputs(6235) <= not(inputs(80));
    layer0_outputs(6236) <= (inputs(125)) xor (inputs(77));
    layer0_outputs(6237) <= not(inputs(145)) or (inputs(127));
    layer0_outputs(6238) <= inputs(156);
    layer0_outputs(6239) <= inputs(172);
    layer0_outputs(6240) <= (inputs(153)) or (inputs(68));
    layer0_outputs(6241) <= (inputs(6)) or (inputs(80));
    layer0_outputs(6242) <= not((inputs(253)) xor (inputs(230)));
    layer0_outputs(6243) <= inputs(23);
    layer0_outputs(6244) <= not(inputs(9));
    layer0_outputs(6245) <= inputs(55);
    layer0_outputs(6246) <= (inputs(235)) and not (inputs(95));
    layer0_outputs(6247) <= not(inputs(115)) or (inputs(47));
    layer0_outputs(6248) <= not(inputs(248));
    layer0_outputs(6249) <= (inputs(240)) or (inputs(18));
    layer0_outputs(6250) <= not(inputs(116)) or (inputs(110));
    layer0_outputs(6251) <= not(inputs(201));
    layer0_outputs(6252) <= (inputs(58)) or (inputs(109));
    layer0_outputs(6253) <= not((inputs(169)) xor (inputs(6)));
    layer0_outputs(6254) <= (inputs(62)) xor (inputs(0));
    layer0_outputs(6255) <= not(inputs(158));
    layer0_outputs(6256) <= not((inputs(200)) or (inputs(128)));
    layer0_outputs(6257) <= (inputs(97)) or (inputs(94));
    layer0_outputs(6258) <= not((inputs(212)) or (inputs(159)));
    layer0_outputs(6259) <= not(inputs(231)) or (inputs(73));
    layer0_outputs(6260) <= (inputs(130)) xor (inputs(209));
    layer0_outputs(6261) <= not(inputs(244)) or (inputs(181));
    layer0_outputs(6262) <= inputs(215);
    layer0_outputs(6263) <= not(inputs(253)) or (inputs(94));
    layer0_outputs(6264) <= not((inputs(11)) xor (inputs(24)));
    layer0_outputs(6265) <= (inputs(221)) xor (inputs(157));
    layer0_outputs(6266) <= '0';
    layer0_outputs(6267) <= not((inputs(109)) or (inputs(17)));
    layer0_outputs(6268) <= not(inputs(164));
    layer0_outputs(6269) <= (inputs(185)) xor (inputs(180));
    layer0_outputs(6270) <= (inputs(245)) or (inputs(177));
    layer0_outputs(6271) <= not((inputs(97)) or (inputs(220)));
    layer0_outputs(6272) <= not((inputs(44)) xor (inputs(0)));
    layer0_outputs(6273) <= inputs(246);
    layer0_outputs(6274) <= not(inputs(21));
    layer0_outputs(6275) <= inputs(229);
    layer0_outputs(6276) <= (inputs(211)) and (inputs(147));
    layer0_outputs(6277) <= (inputs(132)) xor (inputs(117));
    layer0_outputs(6278) <= not((inputs(184)) or (inputs(198)));
    layer0_outputs(6279) <= not((inputs(97)) or (inputs(217)));
    layer0_outputs(6280) <= not(inputs(84));
    layer0_outputs(6281) <= not((inputs(95)) xor (inputs(20)));
    layer0_outputs(6282) <= not((inputs(251)) and (inputs(206)));
    layer0_outputs(6283) <= (inputs(31)) and not (inputs(174));
    layer0_outputs(6284) <= not((inputs(238)) or (inputs(248)));
    layer0_outputs(6285) <= (inputs(144)) or (inputs(183));
    layer0_outputs(6286) <= not((inputs(133)) xor (inputs(198)));
    layer0_outputs(6287) <= (inputs(19)) and not (inputs(237));
    layer0_outputs(6288) <= inputs(164);
    layer0_outputs(6289) <= not((inputs(8)) xor (inputs(244)));
    layer0_outputs(6290) <= not((inputs(227)) or (inputs(60)));
    layer0_outputs(6291) <= (inputs(116)) xor (inputs(144));
    layer0_outputs(6292) <= (inputs(73)) xor (inputs(196));
    layer0_outputs(6293) <= inputs(87);
    layer0_outputs(6294) <= inputs(77);
    layer0_outputs(6295) <= (inputs(203)) or (inputs(222));
    layer0_outputs(6296) <= not(inputs(149)) or (inputs(202));
    layer0_outputs(6297) <= (inputs(226)) and not (inputs(81));
    layer0_outputs(6298) <= not((inputs(88)) xor (inputs(120)));
    layer0_outputs(6299) <= not(inputs(210));
    layer0_outputs(6300) <= (inputs(109)) and not (inputs(213));
    layer0_outputs(6301) <= (inputs(155)) xor (inputs(2));
    layer0_outputs(6302) <= not((inputs(223)) or (inputs(69)));
    layer0_outputs(6303) <= not(inputs(18));
    layer0_outputs(6304) <= not((inputs(157)) xor (inputs(120)));
    layer0_outputs(6305) <= inputs(123);
    layer0_outputs(6306) <= (inputs(211)) or (inputs(171));
    layer0_outputs(6307) <= not(inputs(167)) or (inputs(55));
    layer0_outputs(6308) <= not(inputs(114));
    layer0_outputs(6309) <= (inputs(119)) and not (inputs(94));
    layer0_outputs(6310) <= inputs(26);
    layer0_outputs(6311) <= not(inputs(231));
    layer0_outputs(6312) <= not((inputs(162)) xor (inputs(101)));
    layer0_outputs(6313) <= inputs(22);
    layer0_outputs(6314) <= not((inputs(191)) or (inputs(123)));
    layer0_outputs(6315) <= not(inputs(3));
    layer0_outputs(6316) <= not((inputs(137)) or (inputs(140)));
    layer0_outputs(6317) <= (inputs(101)) xor (inputs(20));
    layer0_outputs(6318) <= not(inputs(22));
    layer0_outputs(6319) <= not((inputs(51)) xor (inputs(40)));
    layer0_outputs(6320) <= (inputs(173)) or (inputs(126));
    layer0_outputs(6321) <= (inputs(178)) or (inputs(69));
    layer0_outputs(6322) <= inputs(46);
    layer0_outputs(6323) <= inputs(4);
    layer0_outputs(6324) <= (inputs(239)) or (inputs(103));
    layer0_outputs(6325) <= (inputs(44)) and not (inputs(173));
    layer0_outputs(6326) <= (inputs(145)) xor (inputs(165));
    layer0_outputs(6327) <= inputs(182);
    layer0_outputs(6328) <= '1';
    layer0_outputs(6329) <= (inputs(88)) and (inputs(89));
    layer0_outputs(6330) <= (inputs(55)) and not (inputs(247));
    layer0_outputs(6331) <= inputs(137);
    layer0_outputs(6332) <= (inputs(181)) or (inputs(227));
    layer0_outputs(6333) <= not((inputs(155)) or (inputs(240)));
    layer0_outputs(6334) <= '1';
    layer0_outputs(6335) <= not(inputs(202)) or (inputs(192));
    layer0_outputs(6336) <= (inputs(23)) xor (inputs(121));
    layer0_outputs(6337) <= (inputs(66)) and not (inputs(60));
    layer0_outputs(6338) <= (inputs(165)) and not (inputs(224));
    layer0_outputs(6339) <= not(inputs(194));
    layer0_outputs(6340) <= not((inputs(225)) xor (inputs(247)));
    layer0_outputs(6341) <= not(inputs(76)) or (inputs(219));
    layer0_outputs(6342) <= (inputs(12)) or (inputs(173));
    layer0_outputs(6343) <= not((inputs(211)) xor (inputs(135)));
    layer0_outputs(6344) <= not((inputs(81)) xor (inputs(84)));
    layer0_outputs(6345) <= inputs(212);
    layer0_outputs(6346) <= '0';
    layer0_outputs(6347) <= (inputs(1)) or (inputs(32));
    layer0_outputs(6348) <= not(inputs(62)) or (inputs(3));
    layer0_outputs(6349) <= not(inputs(93));
    layer0_outputs(6350) <= (inputs(190)) or (inputs(203));
    layer0_outputs(6351) <= (inputs(49)) xor (inputs(68));
    layer0_outputs(6352) <= inputs(94);
    layer0_outputs(6353) <= not(inputs(85));
    layer0_outputs(6354) <= not((inputs(75)) xor (inputs(128)));
    layer0_outputs(6355) <= (inputs(228)) and not (inputs(159));
    layer0_outputs(6356) <= (inputs(235)) or (inputs(233));
    layer0_outputs(6357) <= not(inputs(177));
    layer0_outputs(6358) <= not(inputs(71)) or (inputs(74));
    layer0_outputs(6359) <= not((inputs(26)) xor (inputs(77)));
    layer0_outputs(6360) <= not((inputs(123)) and (inputs(60)));
    layer0_outputs(6361) <= (inputs(117)) and not (inputs(255));
    layer0_outputs(6362) <= inputs(106);
    layer0_outputs(6363) <= (inputs(24)) xor (inputs(88));
    layer0_outputs(6364) <= not(inputs(209));
    layer0_outputs(6365) <= not(inputs(135));
    layer0_outputs(6366) <= not((inputs(61)) xor (inputs(103)));
    layer0_outputs(6367) <= not((inputs(50)) or (inputs(50)));
    layer0_outputs(6368) <= (inputs(69)) and not (inputs(78));
    layer0_outputs(6369) <= not((inputs(201)) or (inputs(157)));
    layer0_outputs(6370) <= (inputs(187)) and not (inputs(29));
    layer0_outputs(6371) <= not(inputs(32)) or (inputs(236));
    layer0_outputs(6372) <= inputs(99);
    layer0_outputs(6373) <= not(inputs(219)) or (inputs(61));
    layer0_outputs(6374) <= not(inputs(246));
    layer0_outputs(6375) <= not((inputs(2)) or (inputs(15)));
    layer0_outputs(6376) <= (inputs(146)) xor (inputs(165));
    layer0_outputs(6377) <= not((inputs(84)) xor (inputs(135)));
    layer0_outputs(6378) <= (inputs(98)) and not (inputs(235));
    layer0_outputs(6379) <= not((inputs(169)) or (inputs(135)));
    layer0_outputs(6380) <= inputs(99);
    layer0_outputs(6381) <= (inputs(77)) xor (inputs(52));
    layer0_outputs(6382) <= not(inputs(244)) or (inputs(145));
    layer0_outputs(6383) <= inputs(4);
    layer0_outputs(6384) <= not((inputs(158)) and (inputs(210)));
    layer0_outputs(6385) <= not(inputs(250));
    layer0_outputs(6386) <= not((inputs(181)) and (inputs(197)));
    layer0_outputs(6387) <= not(inputs(198));
    layer0_outputs(6388) <= not((inputs(179)) xor (inputs(177)));
    layer0_outputs(6389) <= not(inputs(136));
    layer0_outputs(6390) <= not((inputs(138)) xor (inputs(211)));
    layer0_outputs(6391) <= (inputs(246)) and not (inputs(107));
    layer0_outputs(6392) <= not((inputs(214)) or (inputs(192)));
    layer0_outputs(6393) <= (inputs(196)) or (inputs(228));
    layer0_outputs(6394) <= not(inputs(215));
    layer0_outputs(6395) <= inputs(175);
    layer0_outputs(6396) <= (inputs(18)) and not (inputs(234));
    layer0_outputs(6397) <= inputs(71);
    layer0_outputs(6398) <= inputs(38);
    layer0_outputs(6399) <= (inputs(45)) and (inputs(65));
    layer0_outputs(6400) <= not((inputs(8)) or (inputs(205)));
    layer0_outputs(6401) <= (inputs(229)) and not (inputs(33));
    layer0_outputs(6402) <= not(inputs(209));
    layer0_outputs(6403) <= (inputs(71)) xor (inputs(74));
    layer0_outputs(6404) <= not((inputs(116)) xor (inputs(133)));
    layer0_outputs(6405) <= (inputs(120)) and (inputs(102));
    layer0_outputs(6406) <= '1';
    layer0_outputs(6407) <= inputs(93);
    layer0_outputs(6408) <= not(inputs(32)) or (inputs(221));
    layer0_outputs(6409) <= not((inputs(217)) xor (inputs(253)));
    layer0_outputs(6410) <= not(inputs(167));
    layer0_outputs(6411) <= not(inputs(7)) or (inputs(17));
    layer0_outputs(6412) <= not((inputs(28)) xor (inputs(216)));
    layer0_outputs(6413) <= not((inputs(148)) xor (inputs(151)));
    layer0_outputs(6414) <= (inputs(204)) xor (inputs(195));
    layer0_outputs(6415) <= not(inputs(55));
    layer0_outputs(6416) <= inputs(240);
    layer0_outputs(6417) <= not(inputs(103)) or (inputs(10));
    layer0_outputs(6418) <= (inputs(189)) and (inputs(235));
    layer0_outputs(6419) <= inputs(49);
    layer0_outputs(6420) <= inputs(54);
    layer0_outputs(6421) <= inputs(124);
    layer0_outputs(6422) <= not(inputs(228));
    layer0_outputs(6423) <= (inputs(228)) and not (inputs(173));
    layer0_outputs(6424) <= (inputs(118)) xor (inputs(174));
    layer0_outputs(6425) <= (inputs(180)) or (inputs(250));
    layer0_outputs(6426) <= not(inputs(25));
    layer0_outputs(6427) <= (inputs(145)) or (inputs(196));
    layer0_outputs(6428) <= (inputs(51)) xor (inputs(54));
    layer0_outputs(6429) <= not(inputs(18));
    layer0_outputs(6430) <= inputs(20);
    layer0_outputs(6431) <= not((inputs(207)) and (inputs(232)));
    layer0_outputs(6432) <= not((inputs(20)) xor (inputs(65)));
    layer0_outputs(6433) <= not(inputs(100)) or (inputs(3));
    layer0_outputs(6434) <= not(inputs(195));
    layer0_outputs(6435) <= not((inputs(113)) or (inputs(98)));
    layer0_outputs(6436) <= not(inputs(168)) or (inputs(19));
    layer0_outputs(6437) <= not((inputs(236)) or (inputs(245)));
    layer0_outputs(6438) <= inputs(216);
    layer0_outputs(6439) <= inputs(127);
    layer0_outputs(6440) <= inputs(123);
    layer0_outputs(6441) <= (inputs(91)) or (inputs(130));
    layer0_outputs(6442) <= inputs(60);
    layer0_outputs(6443) <= not(inputs(245));
    layer0_outputs(6444) <= not(inputs(100)) or (inputs(32));
    layer0_outputs(6445) <= (inputs(3)) and not (inputs(76));
    layer0_outputs(6446) <= not(inputs(39)) or (inputs(132));
    layer0_outputs(6447) <= inputs(21);
    layer0_outputs(6448) <= not(inputs(60));
    layer0_outputs(6449) <= (inputs(101)) and not (inputs(128));
    layer0_outputs(6450) <= not(inputs(95));
    layer0_outputs(6451) <= not((inputs(138)) or (inputs(238)));
    layer0_outputs(6452) <= (inputs(38)) and not (inputs(29));
    layer0_outputs(6453) <= not(inputs(231));
    layer0_outputs(6454) <= not(inputs(209));
    layer0_outputs(6455) <= not((inputs(161)) xor (inputs(165)));
    layer0_outputs(6456) <= not(inputs(253));
    layer0_outputs(6457) <= (inputs(193)) or (inputs(87));
    layer0_outputs(6458) <= not(inputs(7)) or (inputs(28));
    layer0_outputs(6459) <= inputs(231);
    layer0_outputs(6460) <= (inputs(239)) xor (inputs(157));
    layer0_outputs(6461) <= not((inputs(217)) xor (inputs(134)));
    layer0_outputs(6462) <= (inputs(223)) or (inputs(242));
    layer0_outputs(6463) <= not((inputs(147)) xor (inputs(159)));
    layer0_outputs(6464) <= not((inputs(211)) and (inputs(230)));
    layer0_outputs(6465) <= (inputs(152)) or (inputs(59));
    layer0_outputs(6466) <= inputs(153);
    layer0_outputs(6467) <= not((inputs(104)) xor (inputs(59)));
    layer0_outputs(6468) <= not(inputs(220));
    layer0_outputs(6469) <= not((inputs(56)) or (inputs(95)));
    layer0_outputs(6470) <= '0';
    layer0_outputs(6471) <= (inputs(201)) and not (inputs(135));
    layer0_outputs(6472) <= not(inputs(22));
    layer0_outputs(6473) <= (inputs(142)) xor (inputs(246));
    layer0_outputs(6474) <= not((inputs(79)) or (inputs(76)));
    layer0_outputs(6475) <= inputs(1);
    layer0_outputs(6476) <= (inputs(114)) and not (inputs(191));
    layer0_outputs(6477) <= (inputs(5)) xor (inputs(219));
    layer0_outputs(6478) <= not((inputs(105)) xor (inputs(237)));
    layer0_outputs(6479) <= inputs(25);
    layer0_outputs(6480) <= (inputs(226)) xor (inputs(48));
    layer0_outputs(6481) <= not(inputs(67)) or (inputs(48));
    layer0_outputs(6482) <= not((inputs(119)) or (inputs(206)));
    layer0_outputs(6483) <= not((inputs(192)) or (inputs(95)));
    layer0_outputs(6484) <= not(inputs(184)) or (inputs(128));
    layer0_outputs(6485) <= not(inputs(163));
    layer0_outputs(6486) <= not((inputs(168)) xor (inputs(124)));
    layer0_outputs(6487) <= (inputs(235)) xor (inputs(193));
    layer0_outputs(6488) <= (inputs(54)) or (inputs(44));
    layer0_outputs(6489) <= not((inputs(77)) or (inputs(150)));
    layer0_outputs(6490) <= inputs(59);
    layer0_outputs(6491) <= (inputs(134)) xor (inputs(212));
    layer0_outputs(6492) <= (inputs(59)) or (inputs(185));
    layer0_outputs(6493) <= not((inputs(228)) and (inputs(140)));
    layer0_outputs(6494) <= (inputs(71)) or (inputs(64));
    layer0_outputs(6495) <= not((inputs(238)) or (inputs(163)));
    layer0_outputs(6496) <= inputs(89);
    layer0_outputs(6497) <= '1';
    layer0_outputs(6498) <= not((inputs(176)) xor (inputs(236)));
    layer0_outputs(6499) <= inputs(132);
    layer0_outputs(6500) <= not((inputs(114)) or (inputs(247)));
    layer0_outputs(6501) <= not((inputs(164)) xor (inputs(157)));
    layer0_outputs(6502) <= not(inputs(118)) or (inputs(14));
    layer0_outputs(6503) <= (inputs(216)) or (inputs(199));
    layer0_outputs(6504) <= '1';
    layer0_outputs(6505) <= (inputs(29)) xor (inputs(47));
    layer0_outputs(6506) <= (inputs(101)) or (inputs(100));
    layer0_outputs(6507) <= (inputs(60)) and not (inputs(239));
    layer0_outputs(6508) <= (inputs(77)) or (inputs(178));
    layer0_outputs(6509) <= not((inputs(111)) or (inputs(111)));
    layer0_outputs(6510) <= (inputs(152)) xor (inputs(189));
    layer0_outputs(6511) <= inputs(228);
    layer0_outputs(6512) <= (inputs(208)) and not (inputs(247));
    layer0_outputs(6513) <= (inputs(108)) xor (inputs(139));
    layer0_outputs(6514) <= not(inputs(75));
    layer0_outputs(6515) <= inputs(128);
    layer0_outputs(6516) <= (inputs(84)) xor (inputs(130));
    layer0_outputs(6517) <= inputs(57);
    layer0_outputs(6518) <= '0';
    layer0_outputs(6519) <= inputs(4);
    layer0_outputs(6520) <= (inputs(220)) and not (inputs(15));
    layer0_outputs(6521) <= (inputs(80)) or (inputs(119));
    layer0_outputs(6522) <= not(inputs(70));
    layer0_outputs(6523) <= not((inputs(221)) or (inputs(179)));
    layer0_outputs(6524) <= (inputs(18)) xor (inputs(146));
    layer0_outputs(6525) <= inputs(133);
    layer0_outputs(6526) <= not(inputs(216));
    layer0_outputs(6527) <= not((inputs(68)) or (inputs(170)));
    layer0_outputs(6528) <= not(inputs(122));
    layer0_outputs(6529) <= not(inputs(79));
    layer0_outputs(6530) <= inputs(244);
    layer0_outputs(6531) <= not(inputs(66)) or (inputs(70));
    layer0_outputs(6532) <= (inputs(236)) xor (inputs(102));
    layer0_outputs(6533) <= inputs(215);
    layer0_outputs(6534) <= inputs(23);
    layer0_outputs(6535) <= '1';
    layer0_outputs(6536) <= (inputs(213)) xor (inputs(184));
    layer0_outputs(6537) <= not(inputs(38));
    layer0_outputs(6538) <= not(inputs(92));
    layer0_outputs(6539) <= not(inputs(224)) or (inputs(125));
    layer0_outputs(6540) <= (inputs(112)) or (inputs(30));
    layer0_outputs(6541) <= (inputs(169)) or (inputs(171));
    layer0_outputs(6542) <= not((inputs(107)) xor (inputs(3)));
    layer0_outputs(6543) <= (inputs(33)) or (inputs(59));
    layer0_outputs(6544) <= not(inputs(103)) or (inputs(190));
    layer0_outputs(6545) <= not(inputs(68));
    layer0_outputs(6546) <= (inputs(10)) or (inputs(116));
    layer0_outputs(6547) <= (inputs(27)) or (inputs(51));
    layer0_outputs(6548) <= not((inputs(205)) and (inputs(48)));
    layer0_outputs(6549) <= (inputs(223)) xor (inputs(219));
    layer0_outputs(6550) <= inputs(3);
    layer0_outputs(6551) <= inputs(5);
    layer0_outputs(6552) <= (inputs(220)) xor (inputs(14));
    layer0_outputs(6553) <= not((inputs(3)) or (inputs(121)));
    layer0_outputs(6554) <= not(inputs(72)) or (inputs(55));
    layer0_outputs(6555) <= not(inputs(89)) or (inputs(221));
    layer0_outputs(6556) <= not(inputs(109));
    layer0_outputs(6557) <= not((inputs(146)) or (inputs(167)));
    layer0_outputs(6558) <= (inputs(187)) xor (inputs(121));
    layer0_outputs(6559) <= not((inputs(161)) and (inputs(250)));
    layer0_outputs(6560) <= not((inputs(246)) xor (inputs(214)));
    layer0_outputs(6561) <= (inputs(23)) xor (inputs(38));
    layer0_outputs(6562) <= inputs(214);
    layer0_outputs(6563) <= not((inputs(109)) or (inputs(128)));
    layer0_outputs(6564) <= not(inputs(169));
    layer0_outputs(6565) <= (inputs(185)) and not (inputs(90));
    layer0_outputs(6566) <= not(inputs(236));
    layer0_outputs(6567) <= not(inputs(201)) or (inputs(72));
    layer0_outputs(6568) <= inputs(59);
    layer0_outputs(6569) <= not((inputs(211)) xor (inputs(107)));
    layer0_outputs(6570) <= (inputs(131)) and not (inputs(94));
    layer0_outputs(6571) <= not((inputs(28)) or (inputs(242)));
    layer0_outputs(6572) <= (inputs(100)) and not (inputs(144));
    layer0_outputs(6573) <= not(inputs(124)) or (inputs(198));
    layer0_outputs(6574) <= not((inputs(148)) xor (inputs(118)));
    layer0_outputs(6575) <= not(inputs(253));
    layer0_outputs(6576) <= (inputs(150)) and not (inputs(175));
    layer0_outputs(6577) <= (inputs(109)) or (inputs(20));
    layer0_outputs(6578) <= not((inputs(254)) xor (inputs(154)));
    layer0_outputs(6579) <= not(inputs(8));
    layer0_outputs(6580) <= not((inputs(13)) xor (inputs(22)));
    layer0_outputs(6581) <= not((inputs(14)) and (inputs(202)));
    layer0_outputs(6582) <= inputs(144);
    layer0_outputs(6583) <= (inputs(183)) and not (inputs(97));
    layer0_outputs(6584) <= (inputs(178)) and not (inputs(242));
    layer0_outputs(6585) <= inputs(161);
    layer0_outputs(6586) <= inputs(255);
    layer0_outputs(6587) <= (inputs(170)) or (inputs(153));
    layer0_outputs(6588) <= not(inputs(220));
    layer0_outputs(6589) <= (inputs(55)) and not (inputs(134));
    layer0_outputs(6590) <= (inputs(68)) or (inputs(148));
    layer0_outputs(6591) <= inputs(176);
    layer0_outputs(6592) <= (inputs(249)) or (inputs(64));
    layer0_outputs(6593) <= inputs(245);
    layer0_outputs(6594) <= inputs(66);
    layer0_outputs(6595) <= (inputs(60)) or (inputs(241));
    layer0_outputs(6596) <= (inputs(62)) and not (inputs(118));
    layer0_outputs(6597) <= not(inputs(250)) or (inputs(3));
    layer0_outputs(6598) <= not((inputs(130)) or (inputs(132)));
    layer0_outputs(6599) <= (inputs(187)) xor (inputs(132));
    layer0_outputs(6600) <= (inputs(232)) or (inputs(103));
    layer0_outputs(6601) <= not(inputs(196));
    layer0_outputs(6602) <= (inputs(246)) or (inputs(62));
    layer0_outputs(6603) <= (inputs(63)) xor (inputs(19));
    layer0_outputs(6604) <= not(inputs(165)) or (inputs(50));
    layer0_outputs(6605) <= not((inputs(239)) xor (inputs(210)));
    layer0_outputs(6606) <= '0';
    layer0_outputs(6607) <= (inputs(154)) xor (inputs(106));
    layer0_outputs(6608) <= not(inputs(93));
    layer0_outputs(6609) <= not(inputs(151)) or (inputs(112));
    layer0_outputs(6610) <= inputs(233);
    layer0_outputs(6611) <= (inputs(172)) or (inputs(144));
    layer0_outputs(6612) <= inputs(101);
    layer0_outputs(6613) <= inputs(185);
    layer0_outputs(6614) <= not(inputs(190));
    layer0_outputs(6615) <= not((inputs(210)) and (inputs(216)));
    layer0_outputs(6616) <= (inputs(228)) and not (inputs(245));
    layer0_outputs(6617) <= (inputs(90)) xor (inputs(219));
    layer0_outputs(6618) <= not((inputs(227)) or (inputs(155)));
    layer0_outputs(6619) <= not(inputs(199));
    layer0_outputs(6620) <= (inputs(14)) and not (inputs(45));
    layer0_outputs(6621) <= inputs(61);
    layer0_outputs(6622) <= not(inputs(107)) or (inputs(95));
    layer0_outputs(6623) <= not((inputs(235)) xor (inputs(186)));
    layer0_outputs(6624) <= not((inputs(229)) or (inputs(213)));
    layer0_outputs(6625) <= not((inputs(37)) xor (inputs(5)));
    layer0_outputs(6626) <= (inputs(173)) xor (inputs(139));
    layer0_outputs(6627) <= not(inputs(29)) or (inputs(253));
    layer0_outputs(6628) <= not(inputs(205));
    layer0_outputs(6629) <= inputs(249);
    layer0_outputs(6630) <= (inputs(16)) or (inputs(208));
    layer0_outputs(6631) <= not((inputs(67)) or (inputs(166)));
    layer0_outputs(6632) <= not((inputs(181)) xor (inputs(184)));
    layer0_outputs(6633) <= not((inputs(251)) or (inputs(40)));
    layer0_outputs(6634) <= (inputs(206)) xor (inputs(86));
    layer0_outputs(6635) <= not(inputs(135));
    layer0_outputs(6636) <= not(inputs(117));
    layer0_outputs(6637) <= (inputs(105)) and not (inputs(31));
    layer0_outputs(6638) <= not(inputs(25)) or (inputs(147));
    layer0_outputs(6639) <= not(inputs(13));
    layer0_outputs(6640) <= (inputs(76)) and not (inputs(1));
    layer0_outputs(6641) <= not((inputs(74)) xor (inputs(72)));
    layer0_outputs(6642) <= not((inputs(95)) xor (inputs(177)));
    layer0_outputs(6643) <= inputs(36);
    layer0_outputs(6644) <= not(inputs(103));
    layer0_outputs(6645) <= not(inputs(104)) or (inputs(3));
    layer0_outputs(6646) <= (inputs(121)) and not (inputs(114));
    layer0_outputs(6647) <= not((inputs(117)) xor (inputs(171)));
    layer0_outputs(6648) <= not(inputs(124)) or (inputs(118));
    layer0_outputs(6649) <= not(inputs(119));
    layer0_outputs(6650) <= inputs(193);
    layer0_outputs(6651) <= not((inputs(216)) and (inputs(181)));
    layer0_outputs(6652) <= not(inputs(135)) or (inputs(193));
    layer0_outputs(6653) <= not(inputs(214));
    layer0_outputs(6654) <= (inputs(74)) and not (inputs(110));
    layer0_outputs(6655) <= (inputs(137)) and not (inputs(49));
    layer0_outputs(6656) <= not((inputs(219)) xor (inputs(87)));
    layer0_outputs(6657) <= not((inputs(63)) xor (inputs(246)));
    layer0_outputs(6658) <= (inputs(42)) and (inputs(244));
    layer0_outputs(6659) <= (inputs(9)) or (inputs(3));
    layer0_outputs(6660) <= inputs(73);
    layer0_outputs(6661) <= (inputs(157)) or (inputs(85));
    layer0_outputs(6662) <= (inputs(39)) or (inputs(130));
    layer0_outputs(6663) <= (inputs(191)) and (inputs(11));
    layer0_outputs(6664) <= not(inputs(38));
    layer0_outputs(6665) <= not((inputs(178)) xor (inputs(90)));
    layer0_outputs(6666) <= not(inputs(193)) or (inputs(249));
    layer0_outputs(6667) <= not((inputs(120)) xor (inputs(127)));
    layer0_outputs(6668) <= not((inputs(233)) or (inputs(63)));
    layer0_outputs(6669) <= not((inputs(182)) xor (inputs(137)));
    layer0_outputs(6670) <= inputs(124);
    layer0_outputs(6671) <= inputs(234);
    layer0_outputs(6672) <= inputs(13);
    layer0_outputs(6673) <= not(inputs(173)) or (inputs(76));
    layer0_outputs(6674) <= not(inputs(235)) or (inputs(12));
    layer0_outputs(6675) <= not((inputs(137)) xor (inputs(233)));
    layer0_outputs(6676) <= (inputs(137)) and not (inputs(117));
    layer0_outputs(6677) <= not((inputs(22)) or (inputs(134)));
    layer0_outputs(6678) <= not((inputs(176)) or (inputs(9)));
    layer0_outputs(6679) <= not(inputs(53)) or (inputs(157));
    layer0_outputs(6680) <= not(inputs(14)) or (inputs(190));
    layer0_outputs(6681) <= not(inputs(23));
    layer0_outputs(6682) <= not((inputs(234)) xor (inputs(171)));
    layer0_outputs(6683) <= not(inputs(207)) or (inputs(186));
    layer0_outputs(6684) <= inputs(119);
    layer0_outputs(6685) <= (inputs(60)) or (inputs(238));
    layer0_outputs(6686) <= not((inputs(112)) xor (inputs(99)));
    layer0_outputs(6687) <= not((inputs(1)) and (inputs(1)));
    layer0_outputs(6688) <= (inputs(153)) and not (inputs(25));
    layer0_outputs(6689) <= (inputs(181)) and not (inputs(171));
    layer0_outputs(6690) <= inputs(59);
    layer0_outputs(6691) <= not((inputs(162)) xor (inputs(64)));
    layer0_outputs(6692) <= not((inputs(25)) or (inputs(95)));
    layer0_outputs(6693) <= inputs(219);
    layer0_outputs(6694) <= not(inputs(230));
    layer0_outputs(6695) <= '1';
    layer0_outputs(6696) <= not((inputs(26)) and (inputs(166)));
    layer0_outputs(6697) <= (inputs(219)) or (inputs(62));
    layer0_outputs(6698) <= not(inputs(32)) or (inputs(17));
    layer0_outputs(6699) <= not((inputs(2)) or (inputs(17)));
    layer0_outputs(6700) <= (inputs(224)) or (inputs(16));
    layer0_outputs(6701) <= not((inputs(56)) and (inputs(144)));
    layer0_outputs(6702) <= inputs(28);
    layer0_outputs(6703) <= not((inputs(221)) xor (inputs(10)));
    layer0_outputs(6704) <= (inputs(125)) or (inputs(99));
    layer0_outputs(6705) <= not(inputs(214));
    layer0_outputs(6706) <= not(inputs(115));
    layer0_outputs(6707) <= not(inputs(101)) or (inputs(1));
    layer0_outputs(6708) <= (inputs(170)) and (inputs(65));
    layer0_outputs(6709) <= not(inputs(125)) or (inputs(152));
    layer0_outputs(6710) <= (inputs(134)) or (inputs(153));
    layer0_outputs(6711) <= not(inputs(72));
    layer0_outputs(6712) <= (inputs(185)) and not (inputs(111));
    layer0_outputs(6713) <= not((inputs(50)) xor (inputs(218)));
    layer0_outputs(6714) <= '1';
    layer0_outputs(6715) <= (inputs(41)) and not (inputs(101));
    layer0_outputs(6716) <= not(inputs(150)) or (inputs(158));
    layer0_outputs(6717) <= inputs(46);
    layer0_outputs(6718) <= not(inputs(98));
    layer0_outputs(6719) <= not((inputs(100)) xor (inputs(143)));
    layer0_outputs(6720) <= inputs(161);
    layer0_outputs(6721) <= (inputs(194)) and not (inputs(14));
    layer0_outputs(6722) <= not(inputs(92));
    layer0_outputs(6723) <= (inputs(90)) xor (inputs(89));
    layer0_outputs(6724) <= not(inputs(220)) or (inputs(62));
    layer0_outputs(6725) <= not(inputs(74));
    layer0_outputs(6726) <= (inputs(225)) or (inputs(192));
    layer0_outputs(6727) <= not(inputs(63));
    layer0_outputs(6728) <= (inputs(26)) xor (inputs(223));
    layer0_outputs(6729) <= not(inputs(229));
    layer0_outputs(6730) <= (inputs(100)) and not (inputs(217));
    layer0_outputs(6731) <= not(inputs(167));
    layer0_outputs(6732) <= (inputs(41)) or (inputs(123));
    layer0_outputs(6733) <= (inputs(62)) xor (inputs(27));
    layer0_outputs(6734) <= not(inputs(118));
    layer0_outputs(6735) <= (inputs(27)) and not (inputs(168));
    layer0_outputs(6736) <= (inputs(4)) xor (inputs(68));
    layer0_outputs(6737) <= not(inputs(237));
    layer0_outputs(6738) <= not((inputs(45)) or (inputs(30)));
    layer0_outputs(6739) <= (inputs(181)) or (inputs(184));
    layer0_outputs(6740) <= inputs(151);
    layer0_outputs(6741) <= (inputs(119)) and (inputs(69));
    layer0_outputs(6742) <= (inputs(125)) or (inputs(6));
    layer0_outputs(6743) <= not((inputs(131)) or (inputs(112)));
    layer0_outputs(6744) <= (inputs(22)) and not (inputs(55));
    layer0_outputs(6745) <= inputs(215);
    layer0_outputs(6746) <= not((inputs(139)) or (inputs(157)));
    layer0_outputs(6747) <= inputs(72);
    layer0_outputs(6748) <= not((inputs(36)) xor (inputs(25)));
    layer0_outputs(6749) <= (inputs(135)) and not (inputs(236));
    layer0_outputs(6750) <= (inputs(119)) and not (inputs(81));
    layer0_outputs(6751) <= not(inputs(107));
    layer0_outputs(6752) <= not((inputs(59)) or (inputs(138)));
    layer0_outputs(6753) <= not(inputs(235));
    layer0_outputs(6754) <= (inputs(125)) xor (inputs(243));
    layer0_outputs(6755) <= (inputs(188)) and not (inputs(120));
    layer0_outputs(6756) <= not(inputs(132));
    layer0_outputs(6757) <= inputs(15);
    layer0_outputs(6758) <= not((inputs(44)) or (inputs(221)));
    layer0_outputs(6759) <= inputs(81);
    layer0_outputs(6760) <= (inputs(69)) xor (inputs(22));
    layer0_outputs(6761) <= not(inputs(116));
    layer0_outputs(6762) <= inputs(95);
    layer0_outputs(6763) <= not((inputs(62)) xor (inputs(186)));
    layer0_outputs(6764) <= (inputs(120)) or (inputs(114));
    layer0_outputs(6765) <= (inputs(135)) xor (inputs(172));
    layer0_outputs(6766) <= (inputs(203)) xor (inputs(105));
    layer0_outputs(6767) <= not(inputs(114));
    layer0_outputs(6768) <= not(inputs(29)) or (inputs(101));
    layer0_outputs(6769) <= (inputs(158)) and not (inputs(51));
    layer0_outputs(6770) <= not((inputs(220)) xor (inputs(241)));
    layer0_outputs(6771) <= (inputs(2)) xor (inputs(32));
    layer0_outputs(6772) <= inputs(19);
    layer0_outputs(6773) <= not((inputs(32)) or (inputs(20)));
    layer0_outputs(6774) <= '1';
    layer0_outputs(6775) <= (inputs(54)) and not (inputs(156));
    layer0_outputs(6776) <= (inputs(76)) or (inputs(128));
    layer0_outputs(6777) <= not((inputs(143)) xor (inputs(123)));
    layer0_outputs(6778) <= not((inputs(195)) or (inputs(106)));
    layer0_outputs(6779) <= not(inputs(227)) or (inputs(49));
    layer0_outputs(6780) <= not((inputs(168)) or (inputs(146)));
    layer0_outputs(6781) <= not(inputs(27)) or (inputs(113));
    layer0_outputs(6782) <= not((inputs(1)) or (inputs(130)));
    layer0_outputs(6783) <= not((inputs(207)) or (inputs(225)));
    layer0_outputs(6784) <= (inputs(89)) or (inputs(223));
    layer0_outputs(6785) <= not((inputs(161)) or (inputs(163)));
    layer0_outputs(6786) <= (inputs(1)) or (inputs(125));
    layer0_outputs(6787) <= not(inputs(54));
    layer0_outputs(6788) <= inputs(125);
    layer0_outputs(6789) <= (inputs(162)) and not (inputs(97));
    layer0_outputs(6790) <= inputs(83);
    layer0_outputs(6791) <= not((inputs(73)) xor (inputs(166)));
    layer0_outputs(6792) <= not((inputs(81)) or (inputs(144)));
    layer0_outputs(6793) <= (inputs(38)) and not (inputs(75));
    layer0_outputs(6794) <= (inputs(47)) xor (inputs(243));
    layer0_outputs(6795) <= not(inputs(166)) or (inputs(143));
    layer0_outputs(6796) <= not((inputs(189)) and (inputs(132)));
    layer0_outputs(6797) <= not(inputs(85));
    layer0_outputs(6798) <= (inputs(100)) and not (inputs(16));
    layer0_outputs(6799) <= inputs(41);
    layer0_outputs(6800) <= (inputs(156)) and not (inputs(30));
    layer0_outputs(6801) <= (inputs(30)) or (inputs(50));
    layer0_outputs(6802) <= not(inputs(166));
    layer0_outputs(6803) <= not(inputs(203));
    layer0_outputs(6804) <= (inputs(5)) or (inputs(58));
    layer0_outputs(6805) <= inputs(166);
    layer0_outputs(6806) <= inputs(33);
    layer0_outputs(6807) <= (inputs(55)) xor (inputs(9));
    layer0_outputs(6808) <= (inputs(254)) and not (inputs(0));
    layer0_outputs(6809) <= (inputs(249)) and not (inputs(78));
    layer0_outputs(6810) <= not((inputs(56)) xor (inputs(43)));
    layer0_outputs(6811) <= not(inputs(23)) or (inputs(162));
    layer0_outputs(6812) <= (inputs(164)) and not (inputs(35));
    layer0_outputs(6813) <= (inputs(190)) xor (inputs(70));
    layer0_outputs(6814) <= (inputs(69)) xor (inputs(81));
    layer0_outputs(6815) <= not((inputs(143)) xor (inputs(131)));
    layer0_outputs(6816) <= not(inputs(234));
    layer0_outputs(6817) <= inputs(165);
    layer0_outputs(6818) <= not(inputs(209)) or (inputs(240));
    layer0_outputs(6819) <= not(inputs(119));
    layer0_outputs(6820) <= inputs(195);
    layer0_outputs(6821) <= not(inputs(140)) or (inputs(251));
    layer0_outputs(6822) <= inputs(24);
    layer0_outputs(6823) <= not((inputs(30)) xor (inputs(194)));
    layer0_outputs(6824) <= not(inputs(205)) or (inputs(22));
    layer0_outputs(6825) <= inputs(93);
    layer0_outputs(6826) <= not(inputs(167)) or (inputs(217));
    layer0_outputs(6827) <= not(inputs(187)) or (inputs(143));
    layer0_outputs(6828) <= (inputs(241)) and (inputs(239));
    layer0_outputs(6829) <= not((inputs(203)) xor (inputs(106)));
    layer0_outputs(6830) <= not(inputs(223));
    layer0_outputs(6831) <= not((inputs(120)) or (inputs(135)));
    layer0_outputs(6832) <= not(inputs(159)) or (inputs(15));
    layer0_outputs(6833) <= (inputs(106)) and (inputs(21));
    layer0_outputs(6834) <= not((inputs(171)) or (inputs(41)));
    layer0_outputs(6835) <= (inputs(148)) xor (inputs(163));
    layer0_outputs(6836) <= (inputs(34)) or (inputs(194));
    layer0_outputs(6837) <= not((inputs(229)) or (inputs(175)));
    layer0_outputs(6838) <= (inputs(201)) and (inputs(225));
    layer0_outputs(6839) <= not((inputs(249)) or (inputs(164)));
    layer0_outputs(6840) <= not((inputs(245)) or (inputs(145)));
    layer0_outputs(6841) <= (inputs(118)) or (inputs(244));
    layer0_outputs(6842) <= inputs(216);
    layer0_outputs(6843) <= not(inputs(88)) or (inputs(145));
    layer0_outputs(6844) <= not(inputs(244)) or (inputs(65));
    layer0_outputs(6845) <= (inputs(177)) xor (inputs(141));
    layer0_outputs(6846) <= (inputs(52)) and not (inputs(142));
    layer0_outputs(6847) <= not(inputs(182));
    layer0_outputs(6848) <= inputs(91);
    layer0_outputs(6849) <= not(inputs(114));
    layer0_outputs(6850) <= inputs(108);
    layer0_outputs(6851) <= not((inputs(75)) xor (inputs(45)));
    layer0_outputs(6852) <= not(inputs(13));
    layer0_outputs(6853) <= not(inputs(62));
    layer0_outputs(6854) <= inputs(90);
    layer0_outputs(6855) <= (inputs(113)) or (inputs(139));
    layer0_outputs(6856) <= not(inputs(160)) or (inputs(86));
    layer0_outputs(6857) <= (inputs(79)) or (inputs(121));
    layer0_outputs(6858) <= not((inputs(198)) or (inputs(96)));
    layer0_outputs(6859) <= (inputs(50)) or (inputs(239));
    layer0_outputs(6860) <= (inputs(150)) and (inputs(194));
    layer0_outputs(6861) <= not(inputs(162));
    layer0_outputs(6862) <= inputs(73);
    layer0_outputs(6863) <= (inputs(163)) xor (inputs(64));
    layer0_outputs(6864) <= not(inputs(52));
    layer0_outputs(6865) <= not((inputs(52)) xor (inputs(117)));
    layer0_outputs(6866) <= not((inputs(120)) xor (inputs(108)));
    layer0_outputs(6867) <= (inputs(188)) or (inputs(160));
    layer0_outputs(6868) <= (inputs(101)) and not (inputs(198));
    layer0_outputs(6869) <= (inputs(148)) and (inputs(14));
    layer0_outputs(6870) <= not((inputs(124)) or (inputs(157)));
    layer0_outputs(6871) <= (inputs(173)) xor (inputs(19));
    layer0_outputs(6872) <= not((inputs(188)) or (inputs(0)));
    layer0_outputs(6873) <= inputs(7);
    layer0_outputs(6874) <= (inputs(37)) or (inputs(19));
    layer0_outputs(6875) <= (inputs(245)) xor (inputs(33));
    layer0_outputs(6876) <= (inputs(33)) xor (inputs(218));
    layer0_outputs(6877) <= (inputs(167)) or (inputs(243));
    layer0_outputs(6878) <= not((inputs(7)) and (inputs(83)));
    layer0_outputs(6879) <= inputs(43);
    layer0_outputs(6880) <= not(inputs(59));
    layer0_outputs(6881) <= not(inputs(163));
    layer0_outputs(6882) <= not(inputs(255));
    layer0_outputs(6883) <= not(inputs(243)) or (inputs(66));
    layer0_outputs(6884) <= '1';
    layer0_outputs(6885) <= '0';
    layer0_outputs(6886) <= not(inputs(121)) or (inputs(160));
    layer0_outputs(6887) <= inputs(123);
    layer0_outputs(6888) <= inputs(41);
    layer0_outputs(6889) <= not(inputs(216)) or (inputs(94));
    layer0_outputs(6890) <= (inputs(49)) xor (inputs(24));
    layer0_outputs(6891) <= inputs(174);
    layer0_outputs(6892) <= not(inputs(165)) or (inputs(115));
    layer0_outputs(6893) <= (inputs(11)) and (inputs(38));
    layer0_outputs(6894) <= not((inputs(168)) or (inputs(167)));
    layer0_outputs(6895) <= not((inputs(29)) xor (inputs(117)));
    layer0_outputs(6896) <= (inputs(18)) xor (inputs(158));
    layer0_outputs(6897) <= not((inputs(37)) and (inputs(230)));
    layer0_outputs(6898) <= (inputs(46)) xor (inputs(111));
    layer0_outputs(6899) <= not((inputs(93)) or (inputs(17)));
    layer0_outputs(6900) <= not(inputs(39));
    layer0_outputs(6901) <= (inputs(49)) xor (inputs(22));
    layer0_outputs(6902) <= (inputs(146)) and (inputs(209));
    layer0_outputs(6903) <= (inputs(156)) and not (inputs(206));
    layer0_outputs(6904) <= (inputs(12)) xor (inputs(72));
    layer0_outputs(6905) <= not((inputs(56)) or (inputs(95)));
    layer0_outputs(6906) <= (inputs(240)) xor (inputs(14));
    layer0_outputs(6907) <= not(inputs(10));
    layer0_outputs(6908) <= (inputs(76)) and (inputs(122));
    layer0_outputs(6909) <= inputs(115);
    layer0_outputs(6910) <= inputs(217);
    layer0_outputs(6911) <= not(inputs(165)) or (inputs(57));
    layer0_outputs(6912) <= (inputs(4)) and not (inputs(161));
    layer0_outputs(6913) <= (inputs(189)) or (inputs(18));
    layer0_outputs(6914) <= not(inputs(201));
    layer0_outputs(6915) <= (inputs(105)) or (inputs(112));
    layer0_outputs(6916) <= (inputs(136)) or (inputs(191));
    layer0_outputs(6917) <= inputs(211);
    layer0_outputs(6918) <= (inputs(181)) or (inputs(94));
    layer0_outputs(6919) <= not((inputs(217)) or (inputs(188)));
    layer0_outputs(6920) <= (inputs(209)) or (inputs(176));
    layer0_outputs(6921) <= not((inputs(36)) and (inputs(149)));
    layer0_outputs(6922) <= (inputs(195)) and not (inputs(95));
    layer0_outputs(6923) <= not((inputs(254)) xor (inputs(10)));
    layer0_outputs(6924) <= not((inputs(0)) or (inputs(46)));
    layer0_outputs(6925) <= not((inputs(210)) or (inputs(175)));
    layer0_outputs(6926) <= not(inputs(231));
    layer0_outputs(6927) <= not(inputs(42)) or (inputs(72));
    layer0_outputs(6928) <= (inputs(228)) and not (inputs(82));
    layer0_outputs(6929) <= (inputs(140)) and not (inputs(73));
    layer0_outputs(6930) <= not(inputs(138));
    layer0_outputs(6931) <= inputs(210);
    layer0_outputs(6932) <= (inputs(140)) and not (inputs(45));
    layer0_outputs(6933) <= (inputs(177)) or (inputs(143));
    layer0_outputs(6934) <= not((inputs(38)) or (inputs(161)));
    layer0_outputs(6935) <= not(inputs(130));
    layer0_outputs(6936) <= (inputs(79)) or (inputs(132));
    layer0_outputs(6937) <= (inputs(237)) and not (inputs(15));
    layer0_outputs(6938) <= not((inputs(61)) or (inputs(211)));
    layer0_outputs(6939) <= inputs(246);
    layer0_outputs(6940) <= (inputs(100)) and not (inputs(24));
    layer0_outputs(6941) <= (inputs(88)) xor (inputs(225));
    layer0_outputs(6942) <= (inputs(54)) xor (inputs(64));
    layer0_outputs(6943) <= (inputs(231)) xor (inputs(160));
    layer0_outputs(6944) <= not(inputs(21));
    layer0_outputs(6945) <= (inputs(4)) or (inputs(147));
    layer0_outputs(6946) <= not(inputs(164));
    layer0_outputs(6947) <= inputs(252);
    layer0_outputs(6948) <= not(inputs(116)) or (inputs(236));
    layer0_outputs(6949) <= (inputs(108)) and not (inputs(194));
    layer0_outputs(6950) <= not(inputs(59)) or (inputs(224));
    layer0_outputs(6951) <= not(inputs(47));
    layer0_outputs(6952) <= inputs(99);
    layer0_outputs(6953) <= (inputs(156)) xor (inputs(66));
    layer0_outputs(6954) <= not((inputs(153)) or (inputs(118)));
    layer0_outputs(6955) <= (inputs(33)) and not (inputs(224));
    layer0_outputs(6956) <= not(inputs(61));
    layer0_outputs(6957) <= (inputs(58)) and (inputs(40));
    layer0_outputs(6958) <= not(inputs(138)) or (inputs(108));
    layer0_outputs(6959) <= not(inputs(98)) or (inputs(192));
    layer0_outputs(6960) <= (inputs(99)) or (inputs(24));
    layer0_outputs(6961) <= (inputs(233)) and not (inputs(103));
    layer0_outputs(6962) <= not((inputs(228)) or (inputs(235)));
    layer0_outputs(6963) <= not(inputs(218));
    layer0_outputs(6964) <= inputs(155);
    layer0_outputs(6965) <= (inputs(70)) and not (inputs(111));
    layer0_outputs(6966) <= (inputs(253)) and (inputs(197));
    layer0_outputs(6967) <= inputs(60);
    layer0_outputs(6968) <= (inputs(220)) or (inputs(250));
    layer0_outputs(6969) <= inputs(39);
    layer0_outputs(6970) <= inputs(202);
    layer0_outputs(6971) <= (inputs(203)) xor (inputs(193));
    layer0_outputs(6972) <= inputs(177);
    layer0_outputs(6973) <= not((inputs(57)) or (inputs(177)));
    layer0_outputs(6974) <= (inputs(138)) or (inputs(237));
    layer0_outputs(6975) <= not((inputs(106)) xor (inputs(154)));
    layer0_outputs(6976) <= inputs(88);
    layer0_outputs(6977) <= not(inputs(54)) or (inputs(13));
    layer0_outputs(6978) <= not((inputs(33)) xor (inputs(235)));
    layer0_outputs(6979) <= not(inputs(236));
    layer0_outputs(6980) <= not(inputs(167));
    layer0_outputs(6981) <= not((inputs(19)) or (inputs(182)));
    layer0_outputs(6982) <= not(inputs(151)) or (inputs(158));
    layer0_outputs(6983) <= (inputs(6)) xor (inputs(176));
    layer0_outputs(6984) <= not(inputs(245)) or (inputs(122));
    layer0_outputs(6985) <= not(inputs(116)) or (inputs(249));
    layer0_outputs(6986) <= (inputs(61)) or (inputs(41));
    layer0_outputs(6987) <= inputs(25);
    layer0_outputs(6988) <= not(inputs(145)) or (inputs(188));
    layer0_outputs(6989) <= not((inputs(9)) xor (inputs(3)));
    layer0_outputs(6990) <= (inputs(114)) xor (inputs(138));
    layer0_outputs(6991) <= not((inputs(180)) xor (inputs(109)));
    layer0_outputs(6992) <= inputs(116);
    layer0_outputs(6993) <= (inputs(38)) or (inputs(1));
    layer0_outputs(6994) <= not((inputs(244)) or (inputs(94)));
    layer0_outputs(6995) <= not(inputs(167)) or (inputs(230));
    layer0_outputs(6996) <= (inputs(124)) or (inputs(163));
    layer0_outputs(6997) <= '1';
    layer0_outputs(6998) <= (inputs(255)) or (inputs(68));
    layer0_outputs(6999) <= not(inputs(117)) or (inputs(140));
    layer0_outputs(7000) <= (inputs(94)) or (inputs(151));
    layer0_outputs(7001) <= not((inputs(113)) or (inputs(76)));
    layer0_outputs(7002) <= (inputs(103)) xor (inputs(35));
    layer0_outputs(7003) <= not((inputs(102)) xor (inputs(35)));
    layer0_outputs(7004) <= not((inputs(34)) xor (inputs(216)));
    layer0_outputs(7005) <= (inputs(22)) and (inputs(202));
    layer0_outputs(7006) <= not((inputs(53)) xor (inputs(78)));
    layer0_outputs(7007) <= (inputs(37)) and not (inputs(190));
    layer0_outputs(7008) <= not((inputs(64)) xor (inputs(54)));
    layer0_outputs(7009) <= (inputs(61)) or (inputs(109));
    layer0_outputs(7010) <= not(inputs(76));
    layer0_outputs(7011) <= (inputs(180)) or (inputs(236));
    layer0_outputs(7012) <= not(inputs(175)) or (inputs(15));
    layer0_outputs(7013) <= not((inputs(20)) or (inputs(160)));
    layer0_outputs(7014) <= (inputs(74)) xor (inputs(98));
    layer0_outputs(7015) <= inputs(26);
    layer0_outputs(7016) <= (inputs(239)) and not (inputs(0));
    layer0_outputs(7017) <= (inputs(92)) and not (inputs(72));
    layer0_outputs(7018) <= not(inputs(38)) or (inputs(173));
    layer0_outputs(7019) <= not(inputs(111));
    layer0_outputs(7020) <= not(inputs(121)) or (inputs(220));
    layer0_outputs(7021) <= not(inputs(163)) or (inputs(77));
    layer0_outputs(7022) <= not(inputs(59));
    layer0_outputs(7023) <= (inputs(134)) xor (inputs(130));
    layer0_outputs(7024) <= not((inputs(77)) xor (inputs(135)));
    layer0_outputs(7025) <= (inputs(87)) and not (inputs(15));
    layer0_outputs(7026) <= not((inputs(39)) and (inputs(225)));
    layer0_outputs(7027) <= inputs(155);
    layer0_outputs(7028) <= not((inputs(55)) or (inputs(112)));
    layer0_outputs(7029) <= not((inputs(38)) xor (inputs(56)));
    layer0_outputs(7030) <= (inputs(118)) or (inputs(137));
    layer0_outputs(7031) <= (inputs(12)) xor (inputs(135));
    layer0_outputs(7032) <= (inputs(150)) and not (inputs(35));
    layer0_outputs(7033) <= (inputs(91)) or (inputs(80));
    layer0_outputs(7034) <= not((inputs(213)) or (inputs(135)));
    layer0_outputs(7035) <= not((inputs(99)) and (inputs(115)));
    layer0_outputs(7036) <= inputs(214);
    layer0_outputs(7037) <= not((inputs(223)) or (inputs(212)));
    layer0_outputs(7038) <= (inputs(43)) xor (inputs(198));
    layer0_outputs(7039) <= (inputs(23)) xor (inputs(85));
    layer0_outputs(7040) <= (inputs(61)) and not (inputs(64));
    layer0_outputs(7041) <= not(inputs(98));
    layer0_outputs(7042) <= inputs(125);
    layer0_outputs(7043) <= inputs(39);
    layer0_outputs(7044) <= inputs(170);
    layer0_outputs(7045) <= (inputs(149)) and not (inputs(75));
    layer0_outputs(7046) <= not(inputs(121));
    layer0_outputs(7047) <= not(inputs(95));
    layer0_outputs(7048) <= not((inputs(154)) xor (inputs(123)));
    layer0_outputs(7049) <= '1';
    layer0_outputs(7050) <= not(inputs(71));
    layer0_outputs(7051) <= not((inputs(84)) or (inputs(211)));
    layer0_outputs(7052) <= not(inputs(192)) or (inputs(223));
    layer0_outputs(7053) <= (inputs(61)) and (inputs(194));
    layer0_outputs(7054) <= not(inputs(91));
    layer0_outputs(7055) <= not((inputs(212)) and (inputs(11)));
    layer0_outputs(7056) <= (inputs(154)) and not (inputs(97));
    layer0_outputs(7057) <= inputs(137);
    layer0_outputs(7058) <= not((inputs(156)) or (inputs(27)));
    layer0_outputs(7059) <= not(inputs(97));
    layer0_outputs(7060) <= (inputs(6)) and not (inputs(99));
    layer0_outputs(7061) <= inputs(88);
    layer0_outputs(7062) <= not(inputs(83));
    layer0_outputs(7063) <= (inputs(122)) and not (inputs(182));
    layer0_outputs(7064) <= not(inputs(227));
    layer0_outputs(7065) <= inputs(72);
    layer0_outputs(7066) <= not(inputs(107));
    layer0_outputs(7067) <= (inputs(36)) and not (inputs(96));
    layer0_outputs(7068) <= (inputs(127)) or (inputs(215));
    layer0_outputs(7069) <= not((inputs(98)) xor (inputs(72)));
    layer0_outputs(7070) <= (inputs(160)) or (inputs(64));
    layer0_outputs(7071) <= not(inputs(148));
    layer0_outputs(7072) <= not(inputs(68));
    layer0_outputs(7073) <= not((inputs(45)) or (inputs(204)));
    layer0_outputs(7074) <= not(inputs(143)) or (inputs(9));
    layer0_outputs(7075) <= not((inputs(93)) and (inputs(64)));
    layer0_outputs(7076) <= '0';
    layer0_outputs(7077) <= not(inputs(167)) or (inputs(15));
    layer0_outputs(7078) <= not((inputs(254)) xor (inputs(242)));
    layer0_outputs(7079) <= not(inputs(201));
    layer0_outputs(7080) <= not(inputs(94));
    layer0_outputs(7081) <= not(inputs(148)) or (inputs(100));
    layer0_outputs(7082) <= not(inputs(70));
    layer0_outputs(7083) <= inputs(146);
    layer0_outputs(7084) <= (inputs(208)) or (inputs(247));
    layer0_outputs(7085) <= (inputs(65)) or (inputs(230));
    layer0_outputs(7086) <= inputs(175);
    layer0_outputs(7087) <= inputs(150);
    layer0_outputs(7088) <= not(inputs(126)) or (inputs(35));
    layer0_outputs(7089) <= (inputs(92)) or (inputs(45));
    layer0_outputs(7090) <= (inputs(6)) and not (inputs(130));
    layer0_outputs(7091) <= not(inputs(7));
    layer0_outputs(7092) <= not(inputs(74));
    layer0_outputs(7093) <= not(inputs(180));
    layer0_outputs(7094) <= not((inputs(38)) or (inputs(98)));
    layer0_outputs(7095) <= inputs(23);
    layer0_outputs(7096) <= inputs(163);
    layer0_outputs(7097) <= (inputs(82)) and (inputs(72));
    layer0_outputs(7098) <= inputs(57);
    layer0_outputs(7099) <= not((inputs(8)) or (inputs(159)));
    layer0_outputs(7100) <= not(inputs(79));
    layer0_outputs(7101) <= (inputs(46)) or (inputs(39));
    layer0_outputs(7102) <= not((inputs(34)) or (inputs(12)));
    layer0_outputs(7103) <= not((inputs(207)) xor (inputs(123)));
    layer0_outputs(7104) <= '1';
    layer0_outputs(7105) <= not(inputs(168)) or (inputs(249));
    layer0_outputs(7106) <= (inputs(235)) or (inputs(253));
    layer0_outputs(7107) <= (inputs(26)) and not (inputs(144));
    layer0_outputs(7108) <= (inputs(107)) and not (inputs(9));
    layer0_outputs(7109) <= not(inputs(3));
    layer0_outputs(7110) <= not((inputs(249)) and (inputs(173)));
    layer0_outputs(7111) <= (inputs(79)) or (inputs(62));
    layer0_outputs(7112) <= not(inputs(10)) or (inputs(242));
    layer0_outputs(7113) <= not((inputs(90)) and (inputs(100)));
    layer0_outputs(7114) <= not((inputs(17)) and (inputs(96)));
    layer0_outputs(7115) <= inputs(124);
    layer0_outputs(7116) <= (inputs(173)) and not (inputs(32));
    layer0_outputs(7117) <= not((inputs(79)) or (inputs(178)));
    layer0_outputs(7118) <= not(inputs(201));
    layer0_outputs(7119) <= not(inputs(167));
    layer0_outputs(7120) <= not(inputs(2)) or (inputs(239));
    layer0_outputs(7121) <= not((inputs(19)) or (inputs(56)));
    layer0_outputs(7122) <= inputs(135);
    layer0_outputs(7123) <= not((inputs(95)) and (inputs(61)));
    layer0_outputs(7124) <= (inputs(171)) and not (inputs(66));
    layer0_outputs(7125) <= (inputs(52)) xor (inputs(209));
    layer0_outputs(7126) <= not((inputs(26)) and (inputs(190)));
    layer0_outputs(7127) <= (inputs(101)) and not (inputs(3));
    layer0_outputs(7128) <= not((inputs(203)) or (inputs(97)));
    layer0_outputs(7129) <= (inputs(202)) xor (inputs(217));
    layer0_outputs(7130) <= (inputs(211)) xor (inputs(58));
    layer0_outputs(7131) <= not(inputs(249)) or (inputs(59));
    layer0_outputs(7132) <= (inputs(123)) and (inputs(83));
    layer0_outputs(7133) <= (inputs(92)) and not (inputs(65));
    layer0_outputs(7134) <= (inputs(160)) and not (inputs(9));
    layer0_outputs(7135) <= (inputs(8)) and not (inputs(241));
    layer0_outputs(7136) <= (inputs(99)) and not (inputs(174));
    layer0_outputs(7137) <= (inputs(236)) or (inputs(168));
    layer0_outputs(7138) <= (inputs(3)) or (inputs(45));
    layer0_outputs(7139) <= not((inputs(63)) and (inputs(15)));
    layer0_outputs(7140) <= inputs(196);
    layer0_outputs(7141) <= (inputs(85)) and not (inputs(234));
    layer0_outputs(7142) <= inputs(228);
    layer0_outputs(7143) <= not((inputs(8)) xor (inputs(10)));
    layer0_outputs(7144) <= not((inputs(85)) or (inputs(66)));
    layer0_outputs(7145) <= '1';
    layer0_outputs(7146) <= not(inputs(178));
    layer0_outputs(7147) <= (inputs(215)) and (inputs(203));
    layer0_outputs(7148) <= (inputs(154)) and not (inputs(20));
    layer0_outputs(7149) <= (inputs(168)) and not (inputs(36));
    layer0_outputs(7150) <= not(inputs(13));
    layer0_outputs(7151) <= inputs(120);
    layer0_outputs(7152) <= inputs(100);
    layer0_outputs(7153) <= not((inputs(203)) or (inputs(134)));
    layer0_outputs(7154) <= not((inputs(202)) or (inputs(233)));
    layer0_outputs(7155) <= not((inputs(195)) or (inputs(128)));
    layer0_outputs(7156) <= inputs(172);
    layer0_outputs(7157) <= (inputs(226)) and (inputs(157));
    layer0_outputs(7158) <= not(inputs(129));
    layer0_outputs(7159) <= (inputs(84)) and not (inputs(18));
    layer0_outputs(7160) <= not(inputs(178)) or (inputs(15));
    layer0_outputs(7161) <= not(inputs(214));
    layer0_outputs(7162) <= (inputs(167)) or (inputs(89));
    layer0_outputs(7163) <= (inputs(172)) or (inputs(69));
    layer0_outputs(7164) <= not(inputs(215)) or (inputs(111));
    layer0_outputs(7165) <= inputs(81);
    layer0_outputs(7166) <= not(inputs(75)) or (inputs(9));
    layer0_outputs(7167) <= not(inputs(101));
    layer0_outputs(7168) <= not(inputs(214));
    layer0_outputs(7169) <= (inputs(177)) and not (inputs(39));
    layer0_outputs(7170) <= (inputs(234)) or (inputs(230));
    layer0_outputs(7171) <= not((inputs(110)) and (inputs(12)));
    layer0_outputs(7172) <= (inputs(229)) and not (inputs(38));
    layer0_outputs(7173) <= inputs(83);
    layer0_outputs(7174) <= (inputs(29)) and (inputs(26));
    layer0_outputs(7175) <= not((inputs(100)) or (inputs(192)));
    layer0_outputs(7176) <= (inputs(26)) and not (inputs(2));
    layer0_outputs(7177) <= not(inputs(231));
    layer0_outputs(7178) <= (inputs(54)) xor (inputs(150));
    layer0_outputs(7179) <= (inputs(80)) or (inputs(231));
    layer0_outputs(7180) <= '1';
    layer0_outputs(7181) <= not(inputs(77)) or (inputs(99));
    layer0_outputs(7182) <= not(inputs(116));
    layer0_outputs(7183) <= (inputs(111)) and not (inputs(255));
    layer0_outputs(7184) <= not(inputs(183)) or (inputs(118));
    layer0_outputs(7185) <= (inputs(11)) and (inputs(48));
    layer0_outputs(7186) <= not((inputs(241)) xor (inputs(213)));
    layer0_outputs(7187) <= (inputs(179)) and not (inputs(175));
    layer0_outputs(7188) <= not(inputs(112));
    layer0_outputs(7189) <= inputs(101);
    layer0_outputs(7190) <= inputs(88);
    layer0_outputs(7191) <= inputs(49);
    layer0_outputs(7192) <= not((inputs(172)) or (inputs(234)));
    layer0_outputs(7193) <= (inputs(210)) xor (inputs(85));
    layer0_outputs(7194) <= (inputs(5)) or (inputs(90));
    layer0_outputs(7195) <= not(inputs(82));
    layer0_outputs(7196) <= inputs(201);
    layer0_outputs(7197) <= (inputs(210)) and not (inputs(15));
    layer0_outputs(7198) <= not(inputs(52)) or (inputs(158));
    layer0_outputs(7199) <= not((inputs(15)) and (inputs(20)));
    layer0_outputs(7200) <= not(inputs(153)) or (inputs(78));
    layer0_outputs(7201) <= not(inputs(85)) or (inputs(126));
    layer0_outputs(7202) <= (inputs(71)) xor (inputs(36));
    layer0_outputs(7203) <= (inputs(133)) and not (inputs(239));
    layer0_outputs(7204) <= (inputs(142)) and not (inputs(33));
    layer0_outputs(7205) <= not(inputs(56));
    layer0_outputs(7206) <= inputs(37);
    layer0_outputs(7207) <= not(inputs(148));
    layer0_outputs(7208) <= (inputs(39)) xor (inputs(211));
    layer0_outputs(7209) <= (inputs(174)) xor (inputs(156));
    layer0_outputs(7210) <= inputs(168);
    layer0_outputs(7211) <= (inputs(154)) and (inputs(185));
    layer0_outputs(7212) <= not(inputs(143)) or (inputs(136));
    layer0_outputs(7213) <= not((inputs(36)) and (inputs(149)));
    layer0_outputs(7214) <= (inputs(84)) and not (inputs(49));
    layer0_outputs(7215) <= not(inputs(51));
    layer0_outputs(7216) <= not((inputs(73)) xor (inputs(8)));
    layer0_outputs(7217) <= not(inputs(180)) or (inputs(20));
    layer0_outputs(7218) <= inputs(92);
    layer0_outputs(7219) <= not(inputs(72));
    layer0_outputs(7220) <= (inputs(173)) and not (inputs(64));
    layer0_outputs(7221) <= (inputs(176)) and not (inputs(139));
    layer0_outputs(7222) <= not(inputs(54)) or (inputs(236));
    layer0_outputs(7223) <= not(inputs(164));
    layer0_outputs(7224) <= (inputs(122)) xor (inputs(169));
    layer0_outputs(7225) <= not((inputs(212)) and (inputs(147)));
    layer0_outputs(7226) <= (inputs(206)) or (inputs(177));
    layer0_outputs(7227) <= not((inputs(144)) xor (inputs(236)));
    layer0_outputs(7228) <= (inputs(166)) xor (inputs(36));
    layer0_outputs(7229) <= inputs(218);
    layer0_outputs(7230) <= not((inputs(222)) or (inputs(137)));
    layer0_outputs(7231) <= (inputs(148)) xor (inputs(159));
    layer0_outputs(7232) <= not((inputs(249)) and (inputs(225)));
    layer0_outputs(7233) <= inputs(120);
    layer0_outputs(7234) <= inputs(178);
    layer0_outputs(7235) <= not(inputs(211));
    layer0_outputs(7236) <= not(inputs(104));
    layer0_outputs(7237) <= not((inputs(173)) or (inputs(233)));
    layer0_outputs(7238) <= not(inputs(19));
    layer0_outputs(7239) <= not(inputs(137));
    layer0_outputs(7240) <= not(inputs(8)) or (inputs(4));
    layer0_outputs(7241) <= not((inputs(89)) xor (inputs(118)));
    layer0_outputs(7242) <= (inputs(192)) xor (inputs(88));
    layer0_outputs(7243) <= inputs(30);
    layer0_outputs(7244) <= inputs(146);
    layer0_outputs(7245) <= not(inputs(222));
    layer0_outputs(7246) <= (inputs(84)) or (inputs(146));
    layer0_outputs(7247) <= not((inputs(29)) or (inputs(19)));
    layer0_outputs(7248) <= not((inputs(233)) xor (inputs(189)));
    layer0_outputs(7249) <= (inputs(25)) or (inputs(93));
    layer0_outputs(7250) <= (inputs(248)) and not (inputs(92));
    layer0_outputs(7251) <= not(inputs(138)) or (inputs(244));
    layer0_outputs(7252) <= not(inputs(183));
    layer0_outputs(7253) <= not((inputs(83)) or (inputs(204)));
    layer0_outputs(7254) <= not(inputs(218)) or (inputs(7));
    layer0_outputs(7255) <= not(inputs(133)) or (inputs(142));
    layer0_outputs(7256) <= not(inputs(215));
    layer0_outputs(7257) <= inputs(130);
    layer0_outputs(7258) <= inputs(27);
    layer0_outputs(7259) <= inputs(57);
    layer0_outputs(7260) <= (inputs(147)) and not (inputs(63));
    layer0_outputs(7261) <= inputs(61);
    layer0_outputs(7262) <= (inputs(27)) xor (inputs(61));
    layer0_outputs(7263) <= (inputs(133)) xor (inputs(119));
    layer0_outputs(7264) <= (inputs(171)) or (inputs(165));
    layer0_outputs(7265) <= not(inputs(248));
    layer0_outputs(7266) <= not(inputs(13));
    layer0_outputs(7267) <= not(inputs(171));
    layer0_outputs(7268) <= (inputs(91)) or (inputs(92));
    layer0_outputs(7269) <= (inputs(68)) xor (inputs(177));
    layer0_outputs(7270) <= not(inputs(23)) or (inputs(113));
    layer0_outputs(7271) <= not(inputs(154)) or (inputs(136));
    layer0_outputs(7272) <= inputs(152);
    layer0_outputs(7273) <= (inputs(61)) xor (inputs(93));
    layer0_outputs(7274) <= inputs(122);
    layer0_outputs(7275) <= not(inputs(34));
    layer0_outputs(7276) <= not((inputs(81)) or (inputs(185)));
    layer0_outputs(7277) <= not(inputs(182)) or (inputs(227));
    layer0_outputs(7278) <= not(inputs(104)) or (inputs(80));
    layer0_outputs(7279) <= not((inputs(75)) or (inputs(154)));
    layer0_outputs(7280) <= not(inputs(20)) or (inputs(182));
    layer0_outputs(7281) <= not((inputs(127)) xor (inputs(251)));
    layer0_outputs(7282) <= inputs(118);
    layer0_outputs(7283) <= inputs(99);
    layer0_outputs(7284) <= (inputs(33)) xor (inputs(3));
    layer0_outputs(7285) <= inputs(109);
    layer0_outputs(7286) <= (inputs(106)) and not (inputs(32));
    layer0_outputs(7287) <= not((inputs(170)) xor (inputs(89)));
    layer0_outputs(7288) <= not((inputs(38)) xor (inputs(48)));
    layer0_outputs(7289) <= inputs(185);
    layer0_outputs(7290) <= (inputs(201)) or (inputs(222));
    layer0_outputs(7291) <= (inputs(16)) xor (inputs(240));
    layer0_outputs(7292) <= (inputs(172)) xor (inputs(253));
    layer0_outputs(7293) <= not(inputs(136)) or (inputs(130));
    layer0_outputs(7294) <= (inputs(13)) and not (inputs(184));
    layer0_outputs(7295) <= not((inputs(234)) or (inputs(151)));
    layer0_outputs(7296) <= (inputs(71)) or (inputs(176));
    layer0_outputs(7297) <= inputs(22);
    layer0_outputs(7298) <= not(inputs(50));
    layer0_outputs(7299) <= not((inputs(112)) or (inputs(163)));
    layer0_outputs(7300) <= not(inputs(40));
    layer0_outputs(7301) <= not((inputs(166)) or (inputs(15)));
    layer0_outputs(7302) <= inputs(121);
    layer0_outputs(7303) <= not((inputs(198)) and (inputs(197)));
    layer0_outputs(7304) <= (inputs(88)) xor (inputs(81));
    layer0_outputs(7305) <= not((inputs(76)) and (inputs(123)));
    layer0_outputs(7306) <= not(inputs(14)) or (inputs(252));
    layer0_outputs(7307) <= (inputs(8)) xor (inputs(233));
    layer0_outputs(7308) <= not(inputs(220)) or (inputs(115));
    layer0_outputs(7309) <= not((inputs(52)) or (inputs(84)));
    layer0_outputs(7310) <= (inputs(186)) and (inputs(71));
    layer0_outputs(7311) <= inputs(37);
    layer0_outputs(7312) <= not((inputs(45)) xor (inputs(88)));
    layer0_outputs(7313) <= (inputs(144)) xor (inputs(12));
    layer0_outputs(7314) <= (inputs(216)) and not (inputs(178));
    layer0_outputs(7315) <= not((inputs(194)) or (inputs(254)));
    layer0_outputs(7316) <= not(inputs(53)) or (inputs(114));
    layer0_outputs(7317) <= (inputs(164)) or (inputs(253));
    layer0_outputs(7318) <= inputs(55);
    layer0_outputs(7319) <= (inputs(83)) xor (inputs(1));
    layer0_outputs(7320) <= not((inputs(88)) or (inputs(99)));
    layer0_outputs(7321) <= (inputs(215)) and not (inputs(5));
    layer0_outputs(7322) <= not(inputs(153));
    layer0_outputs(7323) <= not(inputs(23)) or (inputs(15));
    layer0_outputs(7324) <= inputs(182);
    layer0_outputs(7325) <= not((inputs(194)) or (inputs(37)));
    layer0_outputs(7326) <= not((inputs(232)) or (inputs(94)));
    layer0_outputs(7327) <= not((inputs(236)) or (inputs(140)));
    layer0_outputs(7328) <= (inputs(10)) and not (inputs(140));
    layer0_outputs(7329) <= inputs(40);
    layer0_outputs(7330) <= (inputs(236)) xor (inputs(218));
    layer0_outputs(7331) <= not((inputs(223)) or (inputs(134)));
    layer0_outputs(7332) <= (inputs(170)) xor (inputs(86));
    layer0_outputs(7333) <= not(inputs(153));
    layer0_outputs(7334) <= not(inputs(19));
    layer0_outputs(7335) <= not((inputs(86)) xor (inputs(82)));
    layer0_outputs(7336) <= inputs(185);
    layer0_outputs(7337) <= inputs(95);
    layer0_outputs(7338) <= not((inputs(169)) xor (inputs(26)));
    layer0_outputs(7339) <= inputs(35);
    layer0_outputs(7340) <= (inputs(98)) and not (inputs(40));
    layer0_outputs(7341) <= inputs(77);
    layer0_outputs(7342) <= not(inputs(21));
    layer0_outputs(7343) <= (inputs(205)) or (inputs(170));
    layer0_outputs(7344) <= inputs(14);
    layer0_outputs(7345) <= not((inputs(42)) xor (inputs(245)));
    layer0_outputs(7346) <= not((inputs(72)) xor (inputs(107)));
    layer0_outputs(7347) <= not(inputs(143));
    layer0_outputs(7348) <= not(inputs(195));
    layer0_outputs(7349) <= (inputs(121)) or (inputs(2));
    layer0_outputs(7350) <= not(inputs(59));
    layer0_outputs(7351) <= not(inputs(247));
    layer0_outputs(7352) <= not(inputs(248));
    layer0_outputs(7353) <= (inputs(0)) and (inputs(79));
    layer0_outputs(7354) <= (inputs(82)) or (inputs(159));
    layer0_outputs(7355) <= not(inputs(185)) or (inputs(2));
    layer0_outputs(7356) <= inputs(150);
    layer0_outputs(7357) <= not(inputs(243)) or (inputs(3));
    layer0_outputs(7358) <= not(inputs(69));
    layer0_outputs(7359) <= not(inputs(135));
    layer0_outputs(7360) <= not(inputs(197)) or (inputs(42));
    layer0_outputs(7361) <= not(inputs(213));
    layer0_outputs(7362) <= not((inputs(243)) xor (inputs(178)));
    layer0_outputs(7363) <= (inputs(231)) xor (inputs(215));
    layer0_outputs(7364) <= inputs(40);
    layer0_outputs(7365) <= (inputs(72)) xor (inputs(12));
    layer0_outputs(7366) <= (inputs(192)) and not (inputs(51));
    layer0_outputs(7367) <= (inputs(88)) and not (inputs(236));
    layer0_outputs(7368) <= not(inputs(133)) or (inputs(64));
    layer0_outputs(7369) <= not(inputs(102));
    layer0_outputs(7370) <= not(inputs(35)) or (inputs(134));
    layer0_outputs(7371) <= inputs(206);
    layer0_outputs(7372) <= (inputs(225)) and (inputs(109));
    layer0_outputs(7373) <= not(inputs(215));
    layer0_outputs(7374) <= (inputs(18)) or (inputs(45));
    layer0_outputs(7375) <= not(inputs(122));
    layer0_outputs(7376) <= (inputs(125)) xor (inputs(165));
    layer0_outputs(7377) <= (inputs(174)) xor (inputs(133));
    layer0_outputs(7378) <= not(inputs(104)) or (inputs(181));
    layer0_outputs(7379) <= (inputs(195)) and (inputs(61));
    layer0_outputs(7380) <= (inputs(31)) or (inputs(114));
    layer0_outputs(7381) <= (inputs(122)) xor (inputs(11));
    layer0_outputs(7382) <= (inputs(249)) and (inputs(5));
    layer0_outputs(7383) <= not(inputs(248)) or (inputs(90));
    layer0_outputs(7384) <= (inputs(200)) xor (inputs(86));
    layer0_outputs(7385) <= inputs(200);
    layer0_outputs(7386) <= (inputs(64)) xor (inputs(167));
    layer0_outputs(7387) <= inputs(64);
    layer0_outputs(7388) <= not(inputs(3)) or (inputs(51));
    layer0_outputs(7389) <= not(inputs(212)) or (inputs(51));
    layer0_outputs(7390) <= not((inputs(217)) or (inputs(204)));
    layer0_outputs(7391) <= (inputs(27)) or (inputs(40));
    layer0_outputs(7392) <= (inputs(53)) and (inputs(206));
    layer0_outputs(7393) <= (inputs(42)) and not (inputs(18));
    layer0_outputs(7394) <= (inputs(166)) and not (inputs(16));
    layer0_outputs(7395) <= (inputs(94)) and (inputs(134));
    layer0_outputs(7396) <= not((inputs(43)) or (inputs(50)));
    layer0_outputs(7397) <= not(inputs(32));
    layer0_outputs(7398) <= (inputs(26)) and not (inputs(207));
    layer0_outputs(7399) <= (inputs(112)) or (inputs(98));
    layer0_outputs(7400) <= (inputs(249)) and (inputs(51));
    layer0_outputs(7401) <= not((inputs(123)) xor (inputs(79)));
    layer0_outputs(7402) <= (inputs(243)) xor (inputs(19));
    layer0_outputs(7403) <= inputs(240);
    layer0_outputs(7404) <= not((inputs(65)) or (inputs(106)));
    layer0_outputs(7405) <= inputs(231);
    layer0_outputs(7406) <= inputs(82);
    layer0_outputs(7407) <= not((inputs(163)) xor (inputs(255)));
    layer0_outputs(7408) <= not((inputs(87)) xor (inputs(115)));
    layer0_outputs(7409) <= not(inputs(36));
    layer0_outputs(7410) <= '1';
    layer0_outputs(7411) <= not((inputs(155)) xor (inputs(170)));
    layer0_outputs(7412) <= inputs(235);
    layer0_outputs(7413) <= not(inputs(234));
    layer0_outputs(7414) <= not((inputs(105)) xor (inputs(185)));
    layer0_outputs(7415) <= not(inputs(94));
    layer0_outputs(7416) <= not(inputs(31)) or (inputs(236));
    layer0_outputs(7417) <= (inputs(197)) or (inputs(142));
    layer0_outputs(7418) <= not(inputs(229)) or (inputs(107));
    layer0_outputs(7419) <= (inputs(42)) or (inputs(255));
    layer0_outputs(7420) <= not(inputs(243));
    layer0_outputs(7421) <= not(inputs(85));
    layer0_outputs(7422) <= not((inputs(95)) or (inputs(25)));
    layer0_outputs(7423) <= not(inputs(181)) or (inputs(208));
    layer0_outputs(7424) <= inputs(218);
    layer0_outputs(7425) <= not(inputs(146)) or (inputs(173));
    layer0_outputs(7426) <= not(inputs(73));
    layer0_outputs(7427) <= not(inputs(38)) or (inputs(113));
    layer0_outputs(7428) <= not(inputs(1));
    layer0_outputs(7429) <= inputs(14);
    layer0_outputs(7430) <= (inputs(163)) or (inputs(81));
    layer0_outputs(7431) <= not(inputs(94));
    layer0_outputs(7432) <= (inputs(224)) and not (inputs(99));
    layer0_outputs(7433) <= not(inputs(232));
    layer0_outputs(7434) <= not(inputs(39));
    layer0_outputs(7435) <= not((inputs(164)) xor (inputs(16)));
    layer0_outputs(7436) <= not((inputs(224)) and (inputs(8)));
    layer0_outputs(7437) <= inputs(186);
    layer0_outputs(7438) <= (inputs(85)) xor (inputs(145));
    layer0_outputs(7439) <= inputs(51);
    layer0_outputs(7440) <= inputs(29);
    layer0_outputs(7441) <= not((inputs(248)) or (inputs(185)));
    layer0_outputs(7442) <= (inputs(70)) and not (inputs(146));
    layer0_outputs(7443) <= (inputs(19)) or (inputs(52));
    layer0_outputs(7444) <= (inputs(38)) and not (inputs(127));
    layer0_outputs(7445) <= (inputs(211)) or (inputs(5));
    layer0_outputs(7446) <= not(inputs(83)) or (inputs(134));
    layer0_outputs(7447) <= (inputs(191)) or (inputs(113));
    layer0_outputs(7448) <= inputs(106);
    layer0_outputs(7449) <= inputs(12);
    layer0_outputs(7450) <= (inputs(213)) xor (inputs(182));
    layer0_outputs(7451) <= not(inputs(81));
    layer0_outputs(7452) <= inputs(98);
    layer0_outputs(7453) <= not(inputs(42));
    layer0_outputs(7454) <= not((inputs(107)) or (inputs(2)));
    layer0_outputs(7455) <= inputs(70);
    layer0_outputs(7456) <= (inputs(102)) xor (inputs(56));
    layer0_outputs(7457) <= not((inputs(66)) or (inputs(239)));
    layer0_outputs(7458) <= not(inputs(2));
    layer0_outputs(7459) <= not(inputs(24));
    layer0_outputs(7460) <= not((inputs(174)) xor (inputs(222)));
    layer0_outputs(7461) <= not((inputs(210)) or (inputs(193)));
    layer0_outputs(7462) <= inputs(156);
    layer0_outputs(7463) <= not(inputs(143)) or (inputs(48));
    layer0_outputs(7464) <= not((inputs(229)) xor (inputs(124)));
    layer0_outputs(7465) <= inputs(78);
    layer0_outputs(7466) <= inputs(228);
    layer0_outputs(7467) <= not(inputs(47)) or (inputs(113));
    layer0_outputs(7468) <= (inputs(142)) and not (inputs(153));
    layer0_outputs(7469) <= not(inputs(90)) or (inputs(30));
    layer0_outputs(7470) <= (inputs(192)) and not (inputs(205));
    layer0_outputs(7471) <= (inputs(183)) and (inputs(246));
    layer0_outputs(7472) <= '0';
    layer0_outputs(7473) <= not(inputs(188));
    layer0_outputs(7474) <= not((inputs(141)) xor (inputs(187)));
    layer0_outputs(7475) <= not(inputs(123)) or (inputs(77));
    layer0_outputs(7476) <= inputs(67);
    layer0_outputs(7477) <= inputs(222);
    layer0_outputs(7478) <= not(inputs(111));
    layer0_outputs(7479) <= (inputs(211)) and not (inputs(0));
    layer0_outputs(7480) <= not(inputs(122));
    layer0_outputs(7481) <= not(inputs(151));
    layer0_outputs(7482) <= (inputs(84)) xor (inputs(145));
    layer0_outputs(7483) <= not((inputs(161)) or (inputs(245)));
    layer0_outputs(7484) <= not((inputs(131)) xor (inputs(165)));
    layer0_outputs(7485) <= not(inputs(71));
    layer0_outputs(7486) <= not(inputs(133));
    layer0_outputs(7487) <= (inputs(235)) xor (inputs(220));
    layer0_outputs(7488) <= not((inputs(17)) or (inputs(238)));
    layer0_outputs(7489) <= not((inputs(27)) and (inputs(84)));
    layer0_outputs(7490) <= not(inputs(209));
    layer0_outputs(7491) <= not(inputs(28));
    layer0_outputs(7492) <= not((inputs(64)) or (inputs(131)));
    layer0_outputs(7493) <= not(inputs(123)) or (inputs(215));
    layer0_outputs(7494) <= not(inputs(230)) or (inputs(94));
    layer0_outputs(7495) <= (inputs(2)) or (inputs(225));
    layer0_outputs(7496) <= inputs(238);
    layer0_outputs(7497) <= not(inputs(131)) or (inputs(7));
    layer0_outputs(7498) <= (inputs(194)) and not (inputs(97));
    layer0_outputs(7499) <= (inputs(20)) and (inputs(43));
    layer0_outputs(7500) <= '1';
    layer0_outputs(7501) <= inputs(19);
    layer0_outputs(7502) <= not(inputs(20));
    layer0_outputs(7503) <= inputs(214);
    layer0_outputs(7504) <= (inputs(214)) or (inputs(241));
    layer0_outputs(7505) <= not(inputs(113)) or (inputs(224));
    layer0_outputs(7506) <= (inputs(244)) or (inputs(147));
    layer0_outputs(7507) <= (inputs(51)) or (inputs(202));
    layer0_outputs(7508) <= (inputs(102)) and not (inputs(5));
    layer0_outputs(7509) <= not((inputs(218)) and (inputs(169)));
    layer0_outputs(7510) <= not(inputs(165));
    layer0_outputs(7511) <= (inputs(24)) and not (inputs(168));
    layer0_outputs(7512) <= (inputs(20)) xor (inputs(229));
    layer0_outputs(7513) <= inputs(216);
    layer0_outputs(7514) <= not((inputs(26)) xor (inputs(144)));
    layer0_outputs(7515) <= (inputs(241)) xor (inputs(45));
    layer0_outputs(7516) <= inputs(235);
    layer0_outputs(7517) <= not((inputs(205)) xor (inputs(62)));
    layer0_outputs(7518) <= not(inputs(11));
    layer0_outputs(7519) <= not(inputs(97));
    layer0_outputs(7520) <= (inputs(214)) or (inputs(163));
    layer0_outputs(7521) <= (inputs(206)) or (inputs(149));
    layer0_outputs(7522) <= not((inputs(130)) or (inputs(184)));
    layer0_outputs(7523) <= not(inputs(199));
    layer0_outputs(7524) <= not(inputs(230));
    layer0_outputs(7525) <= not(inputs(188));
    layer0_outputs(7526) <= not((inputs(91)) or (inputs(106)));
    layer0_outputs(7527) <= not(inputs(229));
    layer0_outputs(7528) <= not(inputs(116));
    layer0_outputs(7529) <= not((inputs(237)) or (inputs(196)));
    layer0_outputs(7530) <= (inputs(46)) xor (inputs(55));
    layer0_outputs(7531) <= (inputs(163)) or (inputs(125));
    layer0_outputs(7532) <= inputs(91);
    layer0_outputs(7533) <= not(inputs(172)) or (inputs(242));
    layer0_outputs(7534) <= not((inputs(37)) xor (inputs(71)));
    layer0_outputs(7535) <= '1';
    layer0_outputs(7536) <= (inputs(193)) and not (inputs(20));
    layer0_outputs(7537) <= not((inputs(56)) xor (inputs(49)));
    layer0_outputs(7538) <= (inputs(50)) xor (inputs(18));
    layer0_outputs(7539) <= (inputs(166)) or (inputs(32));
    layer0_outputs(7540) <= not(inputs(9));
    layer0_outputs(7541) <= inputs(229);
    layer0_outputs(7542) <= (inputs(118)) and not (inputs(78));
    layer0_outputs(7543) <= (inputs(24)) xor (inputs(230));
    layer0_outputs(7544) <= not((inputs(218)) or (inputs(235)));
    layer0_outputs(7545) <= not((inputs(96)) or (inputs(98)));
    layer0_outputs(7546) <= not(inputs(217)) or (inputs(141));
    layer0_outputs(7547) <= not(inputs(67));
    layer0_outputs(7548) <= not((inputs(168)) xor (inputs(135)));
    layer0_outputs(7549) <= inputs(136);
    layer0_outputs(7550) <= inputs(201);
    layer0_outputs(7551) <= not(inputs(227));
    layer0_outputs(7552) <= (inputs(54)) and not (inputs(96));
    layer0_outputs(7553) <= (inputs(255)) xor (inputs(137));
    layer0_outputs(7554) <= inputs(87);
    layer0_outputs(7555) <= (inputs(11)) xor (inputs(255));
    layer0_outputs(7556) <= (inputs(3)) or (inputs(159));
    layer0_outputs(7557) <= (inputs(102)) and not (inputs(62));
    layer0_outputs(7558) <= not(inputs(208));
    layer0_outputs(7559) <= (inputs(189)) and not (inputs(168));
    layer0_outputs(7560) <= not((inputs(18)) or (inputs(221)));
    layer0_outputs(7561) <= (inputs(164)) and not (inputs(33));
    layer0_outputs(7562) <= not(inputs(126));
    layer0_outputs(7563) <= not((inputs(64)) xor (inputs(86)));
    layer0_outputs(7564) <= (inputs(90)) and not (inputs(0));
    layer0_outputs(7565) <= inputs(5);
    layer0_outputs(7566) <= (inputs(83)) xor (inputs(158));
    layer0_outputs(7567) <= not(inputs(131));
    layer0_outputs(7568) <= '1';
    layer0_outputs(7569) <= not((inputs(214)) or (inputs(175)));
    layer0_outputs(7570) <= (inputs(97)) or (inputs(99));
    layer0_outputs(7571) <= (inputs(72)) and not (inputs(192));
    layer0_outputs(7572) <= inputs(50);
    layer0_outputs(7573) <= not((inputs(228)) or (inputs(130)));
    layer0_outputs(7574) <= (inputs(194)) or (inputs(23));
    layer0_outputs(7575) <= (inputs(255)) or (inputs(45));
    layer0_outputs(7576) <= not(inputs(112));
    layer0_outputs(7577) <= not(inputs(65)) or (inputs(109));
    layer0_outputs(7578) <= (inputs(248)) xor (inputs(2));
    layer0_outputs(7579) <= (inputs(222)) xor (inputs(244));
    layer0_outputs(7580) <= not(inputs(235));
    layer0_outputs(7581) <= not(inputs(17));
    layer0_outputs(7582) <= (inputs(205)) xor (inputs(206));
    layer0_outputs(7583) <= (inputs(203)) and not (inputs(235));
    layer0_outputs(7584) <= inputs(212);
    layer0_outputs(7585) <= not(inputs(112));
    layer0_outputs(7586) <= not((inputs(36)) or (inputs(107)));
    layer0_outputs(7587) <= not((inputs(92)) or (inputs(59)));
    layer0_outputs(7588) <= not((inputs(202)) or (inputs(18)));
    layer0_outputs(7589) <= (inputs(157)) xor (inputs(193));
    layer0_outputs(7590) <= (inputs(37)) and (inputs(206));
    layer0_outputs(7591) <= not((inputs(28)) xor (inputs(184)));
    layer0_outputs(7592) <= not(inputs(71));
    layer0_outputs(7593) <= not(inputs(84));
    layer0_outputs(7594) <= not((inputs(242)) or (inputs(227)));
    layer0_outputs(7595) <= not(inputs(208));
    layer0_outputs(7596) <= not(inputs(228));
    layer0_outputs(7597) <= (inputs(173)) xor (inputs(220));
    layer0_outputs(7598) <= (inputs(131)) and not (inputs(65));
    layer0_outputs(7599) <= not(inputs(90));
    layer0_outputs(7600) <= inputs(197);
    layer0_outputs(7601) <= not((inputs(105)) xor (inputs(87)));
    layer0_outputs(7602) <= (inputs(159)) or (inputs(197));
    layer0_outputs(7603) <= (inputs(0)) and not (inputs(251));
    layer0_outputs(7604) <= not((inputs(81)) or (inputs(134)));
    layer0_outputs(7605) <= inputs(251);
    layer0_outputs(7606) <= (inputs(195)) or (inputs(28));
    layer0_outputs(7607) <= (inputs(5)) or (inputs(240));
    layer0_outputs(7608) <= (inputs(168)) or (inputs(68));
    layer0_outputs(7609) <= not(inputs(152));
    layer0_outputs(7610) <= not(inputs(166));
    layer0_outputs(7611) <= '1';
    layer0_outputs(7612) <= (inputs(134)) and not (inputs(65));
    layer0_outputs(7613) <= not((inputs(166)) xor (inputs(148)));
    layer0_outputs(7614) <= not((inputs(241)) or (inputs(162)));
    layer0_outputs(7615) <= inputs(238);
    layer0_outputs(7616) <= (inputs(97)) or (inputs(175));
    layer0_outputs(7617) <= not(inputs(212)) or (inputs(128));
    layer0_outputs(7618) <= not(inputs(202));
    layer0_outputs(7619) <= not((inputs(90)) and (inputs(198)));
    layer0_outputs(7620) <= (inputs(86)) xor (inputs(198));
    layer0_outputs(7621) <= (inputs(91)) xor (inputs(127));
    layer0_outputs(7622) <= inputs(89);
    layer0_outputs(7623) <= not((inputs(189)) or (inputs(124)));
    layer0_outputs(7624) <= not((inputs(24)) and (inputs(104)));
    layer0_outputs(7625) <= not((inputs(132)) or (inputs(97)));
    layer0_outputs(7626) <= (inputs(81)) and not (inputs(125));
    layer0_outputs(7627) <= (inputs(26)) or (inputs(121));
    layer0_outputs(7628) <= (inputs(228)) and (inputs(171));
    layer0_outputs(7629) <= not(inputs(221));
    layer0_outputs(7630) <= not((inputs(204)) xor (inputs(59)));
    layer0_outputs(7631) <= (inputs(147)) xor (inputs(240));
    layer0_outputs(7632) <= (inputs(130)) or (inputs(132));
    layer0_outputs(7633) <= not(inputs(115));
    layer0_outputs(7634) <= inputs(65);
    layer0_outputs(7635) <= (inputs(204)) and not (inputs(146));
    layer0_outputs(7636) <= '1';
    layer0_outputs(7637) <= (inputs(222)) and not (inputs(131));
    layer0_outputs(7638) <= not((inputs(70)) xor (inputs(235)));
    layer0_outputs(7639) <= (inputs(174)) and not (inputs(220));
    layer0_outputs(7640) <= not((inputs(50)) and (inputs(42)));
    layer0_outputs(7641) <= not(inputs(40)) or (inputs(170));
    layer0_outputs(7642) <= not(inputs(189));
    layer0_outputs(7643) <= not(inputs(97));
    layer0_outputs(7644) <= (inputs(61)) or (inputs(14));
    layer0_outputs(7645) <= not(inputs(214)) or (inputs(58));
    layer0_outputs(7646) <= inputs(167);
    layer0_outputs(7647) <= not(inputs(31));
    layer0_outputs(7648) <= (inputs(167)) and not (inputs(100));
    layer0_outputs(7649) <= inputs(180);
    layer0_outputs(7650) <= (inputs(186)) xor (inputs(233));
    layer0_outputs(7651) <= not(inputs(164));
    layer0_outputs(7652) <= '0';
    layer0_outputs(7653) <= (inputs(86)) or (inputs(104));
    layer0_outputs(7654) <= not((inputs(141)) or (inputs(2)));
    layer0_outputs(7655) <= not(inputs(97));
    layer0_outputs(7656) <= inputs(116);
    layer0_outputs(7657) <= not((inputs(47)) xor (inputs(29)));
    layer0_outputs(7658) <= not(inputs(156)) or (inputs(29));
    layer0_outputs(7659) <= (inputs(104)) and not (inputs(86));
    layer0_outputs(7660) <= inputs(128);
    layer0_outputs(7661) <= (inputs(96)) xor (inputs(115));
    layer0_outputs(7662) <= not(inputs(188));
    layer0_outputs(7663) <= (inputs(244)) xor (inputs(98));
    layer0_outputs(7664) <= not(inputs(164)) or (inputs(111));
    layer0_outputs(7665) <= (inputs(164)) xor (inputs(130));
    layer0_outputs(7666) <= (inputs(6)) xor (inputs(11));
    layer0_outputs(7667) <= '0';
    layer0_outputs(7668) <= not(inputs(254)) or (inputs(167));
    layer0_outputs(7669) <= not((inputs(175)) xor (inputs(208)));
    layer0_outputs(7670) <= (inputs(246)) or (inputs(78));
    layer0_outputs(7671) <= (inputs(105)) xor (inputs(74));
    layer0_outputs(7672) <= not(inputs(211));
    layer0_outputs(7673) <= (inputs(194)) or (inputs(191));
    layer0_outputs(7674) <= inputs(248);
    layer0_outputs(7675) <= not((inputs(6)) or (inputs(62)));
    layer0_outputs(7676) <= not(inputs(164)) or (inputs(33));
    layer0_outputs(7677) <= inputs(25);
    layer0_outputs(7678) <= not((inputs(52)) xor (inputs(53)));
    layer0_outputs(7679) <= inputs(61);
    layer0_outputs(7680) <= not((inputs(137)) and (inputs(51)));
    layer0_outputs(7681) <= inputs(86);
    layer0_outputs(7682) <= not(inputs(152));
    layer0_outputs(7683) <= inputs(50);
    layer0_outputs(7684) <= not(inputs(176)) or (inputs(79));
    layer0_outputs(7685) <= (inputs(247)) or (inputs(242));
    layer0_outputs(7686) <= not(inputs(142));
    layer0_outputs(7687) <= (inputs(237)) or (inputs(236));
    layer0_outputs(7688) <= not((inputs(84)) or (inputs(87)));
    layer0_outputs(7689) <= not(inputs(173)) or (inputs(242));
    layer0_outputs(7690) <= not(inputs(119)) or (inputs(210));
    layer0_outputs(7691) <= not(inputs(163));
    layer0_outputs(7692) <= not((inputs(10)) and (inputs(232)));
    layer0_outputs(7693) <= (inputs(207)) xor (inputs(213));
    layer0_outputs(7694) <= (inputs(198)) and not (inputs(108));
    layer0_outputs(7695) <= not(inputs(5)) or (inputs(225));
    layer0_outputs(7696) <= not((inputs(211)) xor (inputs(66)));
    layer0_outputs(7697) <= (inputs(122)) xor (inputs(134));
    layer0_outputs(7698) <= (inputs(118)) or (inputs(251));
    layer0_outputs(7699) <= inputs(112);
    layer0_outputs(7700) <= not(inputs(21));
    layer0_outputs(7701) <= (inputs(10)) xor (inputs(92));
    layer0_outputs(7702) <= not(inputs(195)) or (inputs(2));
    layer0_outputs(7703) <= not((inputs(79)) or (inputs(189)));
    layer0_outputs(7704) <= not(inputs(189));
    layer0_outputs(7705) <= not((inputs(238)) xor (inputs(230)));
    layer0_outputs(7706) <= not((inputs(178)) or (inputs(79)));
    layer0_outputs(7707) <= not(inputs(200)) or (inputs(116));
    layer0_outputs(7708) <= (inputs(110)) or (inputs(145));
    layer0_outputs(7709) <= (inputs(37)) or (inputs(107));
    layer0_outputs(7710) <= (inputs(208)) xor (inputs(174));
    layer0_outputs(7711) <= inputs(150);
    layer0_outputs(7712) <= not(inputs(196));
    layer0_outputs(7713) <= inputs(139);
    layer0_outputs(7714) <= (inputs(87)) and not (inputs(208));
    layer0_outputs(7715) <= (inputs(40)) xor (inputs(26));
    layer0_outputs(7716) <= not((inputs(118)) or (inputs(142)));
    layer0_outputs(7717) <= (inputs(145)) or (inputs(124));
    layer0_outputs(7718) <= (inputs(210)) and (inputs(74));
    layer0_outputs(7719) <= inputs(150);
    layer0_outputs(7720) <= not(inputs(24)) or (inputs(88));
    layer0_outputs(7721) <= not((inputs(85)) xor (inputs(249)));
    layer0_outputs(7722) <= not(inputs(162)) or (inputs(14));
    layer0_outputs(7723) <= (inputs(98)) and (inputs(113));
    layer0_outputs(7724) <= not((inputs(179)) xor (inputs(200)));
    layer0_outputs(7725) <= not(inputs(105));
    layer0_outputs(7726) <= inputs(114);
    layer0_outputs(7727) <= not((inputs(202)) xor (inputs(139)));
    layer0_outputs(7728) <= not((inputs(71)) xor (inputs(197)));
    layer0_outputs(7729) <= (inputs(211)) and not (inputs(97));
    layer0_outputs(7730) <= not(inputs(27));
    layer0_outputs(7731) <= inputs(210);
    layer0_outputs(7732) <= not((inputs(124)) xor (inputs(191)));
    layer0_outputs(7733) <= (inputs(185)) and not (inputs(113));
    layer0_outputs(7734) <= (inputs(1)) or (inputs(123));
    layer0_outputs(7735) <= not(inputs(76));
    layer0_outputs(7736) <= not(inputs(131));
    layer0_outputs(7737) <= (inputs(200)) and not (inputs(94));
    layer0_outputs(7738) <= not((inputs(232)) and (inputs(235)));
    layer0_outputs(7739) <= (inputs(172)) and not (inputs(117));
    layer0_outputs(7740) <= not(inputs(179)) or (inputs(15));
    layer0_outputs(7741) <= not((inputs(121)) xor (inputs(251)));
    layer0_outputs(7742) <= not(inputs(25));
    layer0_outputs(7743) <= (inputs(118)) and not (inputs(209));
    layer0_outputs(7744) <= not((inputs(137)) or (inputs(133)));
    layer0_outputs(7745) <= inputs(86);
    layer0_outputs(7746) <= not(inputs(179));
    layer0_outputs(7747) <= not((inputs(204)) or (inputs(30)));
    layer0_outputs(7748) <= not((inputs(40)) and (inputs(91)));
    layer0_outputs(7749) <= (inputs(185)) xor (inputs(120));
    layer0_outputs(7750) <= inputs(209);
    layer0_outputs(7751) <= not((inputs(133)) xor (inputs(221)));
    layer0_outputs(7752) <= (inputs(77)) or (inputs(112));
    layer0_outputs(7753) <= (inputs(25)) or (inputs(191));
    layer0_outputs(7754) <= not(inputs(21));
    layer0_outputs(7755) <= (inputs(82)) or (inputs(58));
    layer0_outputs(7756) <= inputs(91);
    layer0_outputs(7757) <= (inputs(37)) or (inputs(142));
    layer0_outputs(7758) <= not(inputs(62)) or (inputs(205));
    layer0_outputs(7759) <= not((inputs(188)) xor (inputs(210)));
    layer0_outputs(7760) <= (inputs(191)) and (inputs(146));
    layer0_outputs(7761) <= not(inputs(129));
    layer0_outputs(7762) <= not((inputs(135)) xor (inputs(179)));
    layer0_outputs(7763) <= (inputs(56)) and not (inputs(55));
    layer0_outputs(7764) <= inputs(98);
    layer0_outputs(7765) <= inputs(7);
    layer0_outputs(7766) <= not((inputs(188)) xor (inputs(108)));
    layer0_outputs(7767) <= not((inputs(58)) xor (inputs(185)));
    layer0_outputs(7768) <= not(inputs(201)) or (inputs(82));
    layer0_outputs(7769) <= inputs(88);
    layer0_outputs(7770) <= (inputs(119)) or (inputs(31));
    layer0_outputs(7771) <= not((inputs(66)) and (inputs(116)));
    layer0_outputs(7772) <= (inputs(119)) and not (inputs(14));
    layer0_outputs(7773) <= not((inputs(91)) and (inputs(133)));
    layer0_outputs(7774) <= (inputs(91)) and not (inputs(181));
    layer0_outputs(7775) <= (inputs(7)) and (inputs(7));
    layer0_outputs(7776) <= (inputs(221)) and not (inputs(16));
    layer0_outputs(7777) <= (inputs(51)) or (inputs(140));
    layer0_outputs(7778) <= not(inputs(98)) or (inputs(80));
    layer0_outputs(7779) <= inputs(144);
    layer0_outputs(7780) <= not((inputs(198)) xor (inputs(165)));
    layer0_outputs(7781) <= not(inputs(231));
    layer0_outputs(7782) <= (inputs(193)) or (inputs(167));
    layer0_outputs(7783) <= not((inputs(237)) or (inputs(229)));
    layer0_outputs(7784) <= (inputs(109)) or (inputs(251));
    layer0_outputs(7785) <= not((inputs(105)) or (inputs(105)));
    layer0_outputs(7786) <= not((inputs(254)) or (inputs(199)));
    layer0_outputs(7787) <= (inputs(161)) xor (inputs(96));
    layer0_outputs(7788) <= (inputs(124)) or (inputs(34));
    layer0_outputs(7789) <= (inputs(45)) and not (inputs(9));
    layer0_outputs(7790) <= (inputs(205)) xor (inputs(225));
    layer0_outputs(7791) <= not((inputs(72)) or (inputs(159)));
    layer0_outputs(7792) <= not((inputs(204)) or (inputs(159)));
    layer0_outputs(7793) <= not((inputs(135)) xor (inputs(18)));
    layer0_outputs(7794) <= not((inputs(180)) xor (inputs(31)));
    layer0_outputs(7795) <= (inputs(141)) xor (inputs(254));
    layer0_outputs(7796) <= inputs(61);
    layer0_outputs(7797) <= (inputs(171)) xor (inputs(140));
    layer0_outputs(7798) <= inputs(80);
    layer0_outputs(7799) <= (inputs(109)) xor (inputs(61));
    layer0_outputs(7800) <= not(inputs(170));
    layer0_outputs(7801) <= (inputs(121)) and not (inputs(252));
    layer0_outputs(7802) <= not(inputs(51));
    layer0_outputs(7803) <= inputs(199);
    layer0_outputs(7804) <= inputs(60);
    layer0_outputs(7805) <= (inputs(243)) and not (inputs(158));
    layer0_outputs(7806) <= not(inputs(164));
    layer0_outputs(7807) <= not(inputs(40));
    layer0_outputs(7808) <= (inputs(147)) and not (inputs(51));
    layer0_outputs(7809) <= (inputs(130)) and (inputs(114));
    layer0_outputs(7810) <= '0';
    layer0_outputs(7811) <= not(inputs(104));
    layer0_outputs(7812) <= not(inputs(71)) or (inputs(81));
    layer0_outputs(7813) <= (inputs(221)) xor (inputs(139));
    layer0_outputs(7814) <= (inputs(19)) or (inputs(212));
    layer0_outputs(7815) <= not((inputs(246)) and (inputs(172)));
    layer0_outputs(7816) <= not((inputs(33)) xor (inputs(96)));
    layer0_outputs(7817) <= not((inputs(162)) or (inputs(151)));
    layer0_outputs(7818) <= (inputs(73)) or (inputs(64));
    layer0_outputs(7819) <= (inputs(203)) or (inputs(224));
    layer0_outputs(7820) <= (inputs(166)) xor (inputs(129));
    layer0_outputs(7821) <= (inputs(177)) and not (inputs(253));
    layer0_outputs(7822) <= inputs(209);
    layer0_outputs(7823) <= (inputs(58)) xor (inputs(170));
    layer0_outputs(7824) <= not((inputs(117)) or (inputs(197)));
    layer0_outputs(7825) <= not(inputs(231));
    layer0_outputs(7826) <= inputs(149);
    layer0_outputs(7827) <= (inputs(218)) and not (inputs(115));
    layer0_outputs(7828) <= (inputs(32)) or (inputs(81));
    layer0_outputs(7829) <= (inputs(27)) xor (inputs(59));
    layer0_outputs(7830) <= inputs(247);
    layer0_outputs(7831) <= not(inputs(103));
    layer0_outputs(7832) <= (inputs(118)) xor (inputs(3));
    layer0_outputs(7833) <= not(inputs(3));
    layer0_outputs(7834) <= inputs(191);
    layer0_outputs(7835) <= not((inputs(203)) xor (inputs(172)));
    layer0_outputs(7836) <= (inputs(1)) and (inputs(1));
    layer0_outputs(7837) <= '1';
    layer0_outputs(7838) <= not((inputs(88)) or (inputs(141)));
    layer0_outputs(7839) <= (inputs(242)) or (inputs(9));
    layer0_outputs(7840) <= not((inputs(21)) or (inputs(183)));
    layer0_outputs(7841) <= not(inputs(202)) or (inputs(144));
    layer0_outputs(7842) <= (inputs(78)) xor (inputs(126));
    layer0_outputs(7843) <= not((inputs(79)) or (inputs(125)));
    layer0_outputs(7844) <= inputs(200);
    layer0_outputs(7845) <= (inputs(4)) xor (inputs(81));
    layer0_outputs(7846) <= not((inputs(141)) or (inputs(76)));
    layer0_outputs(7847) <= not(inputs(232)) or (inputs(61));
    layer0_outputs(7848) <= not((inputs(158)) xor (inputs(154)));
    layer0_outputs(7849) <= (inputs(227)) xor (inputs(145));
    layer0_outputs(7850) <= not(inputs(233)) or (inputs(81));
    layer0_outputs(7851) <= (inputs(198)) and not (inputs(15));
    layer0_outputs(7852) <= (inputs(54)) or (inputs(95));
    layer0_outputs(7853) <= not(inputs(13)) or (inputs(242));
    layer0_outputs(7854) <= not((inputs(80)) xor (inputs(252)));
    layer0_outputs(7855) <= inputs(108);
    layer0_outputs(7856) <= not((inputs(152)) or (inputs(28)));
    layer0_outputs(7857) <= inputs(147);
    layer0_outputs(7858) <= not(inputs(121));
    layer0_outputs(7859) <= (inputs(20)) or (inputs(193));
    layer0_outputs(7860) <= (inputs(229)) and not (inputs(137));
    layer0_outputs(7861) <= (inputs(3)) and not (inputs(236));
    layer0_outputs(7862) <= (inputs(86)) and not (inputs(126));
    layer0_outputs(7863) <= not(inputs(9));
    layer0_outputs(7864) <= (inputs(66)) or (inputs(181));
    layer0_outputs(7865) <= not(inputs(146));
    layer0_outputs(7866) <= (inputs(236)) and not (inputs(229));
    layer0_outputs(7867) <= not(inputs(62));
    layer0_outputs(7868) <= inputs(235);
    layer0_outputs(7869) <= (inputs(196)) or (inputs(65));
    layer0_outputs(7870) <= not(inputs(212));
    layer0_outputs(7871) <= not(inputs(74)) or (inputs(130));
    layer0_outputs(7872) <= not((inputs(60)) or (inputs(177)));
    layer0_outputs(7873) <= not(inputs(103));
    layer0_outputs(7874) <= not(inputs(185)) or (inputs(97));
    layer0_outputs(7875) <= not((inputs(250)) or (inputs(31)));
    layer0_outputs(7876) <= (inputs(159)) or (inputs(29));
    layer0_outputs(7877) <= (inputs(153)) or (inputs(165));
    layer0_outputs(7878) <= inputs(244);
    layer0_outputs(7879) <= (inputs(75)) and not (inputs(125));
    layer0_outputs(7880) <= not((inputs(83)) xor (inputs(52)));
    layer0_outputs(7881) <= not((inputs(114)) xor (inputs(100)));
    layer0_outputs(7882) <= not(inputs(196)) or (inputs(70));
    layer0_outputs(7883) <= inputs(84);
    layer0_outputs(7884) <= not(inputs(25)) or (inputs(176));
    layer0_outputs(7885) <= '0';
    layer0_outputs(7886) <= not(inputs(114));
    layer0_outputs(7887) <= not((inputs(238)) or (inputs(70)));
    layer0_outputs(7888) <= not((inputs(177)) or (inputs(3)));
    layer0_outputs(7889) <= not(inputs(249)) or (inputs(254));
    layer0_outputs(7890) <= inputs(87);
    layer0_outputs(7891) <= not(inputs(69));
    layer0_outputs(7892) <= not((inputs(228)) and (inputs(168)));
    layer0_outputs(7893) <= not(inputs(87));
    layer0_outputs(7894) <= (inputs(45)) or (inputs(139));
    layer0_outputs(7895) <= inputs(156);
    layer0_outputs(7896) <= not(inputs(193));
    layer0_outputs(7897) <= not(inputs(188));
    layer0_outputs(7898) <= inputs(126);
    layer0_outputs(7899) <= not((inputs(148)) xor (inputs(139)));
    layer0_outputs(7900) <= not((inputs(134)) or (inputs(44)));
    layer0_outputs(7901) <= not(inputs(186)) or (inputs(220));
    layer0_outputs(7902) <= inputs(131);
    layer0_outputs(7903) <= not(inputs(93));
    layer0_outputs(7904) <= inputs(165);
    layer0_outputs(7905) <= not((inputs(4)) xor (inputs(49)));
    layer0_outputs(7906) <= not((inputs(80)) and (inputs(146)));
    layer0_outputs(7907) <= not((inputs(138)) xor (inputs(51)));
    layer0_outputs(7908) <= (inputs(3)) xor (inputs(175));
    layer0_outputs(7909) <= (inputs(255)) or (inputs(190));
    layer0_outputs(7910) <= inputs(231);
    layer0_outputs(7911) <= not((inputs(35)) xor (inputs(229)));
    layer0_outputs(7912) <= not(inputs(70)) or (inputs(227));
    layer0_outputs(7913) <= inputs(39);
    layer0_outputs(7914) <= not(inputs(89)) or (inputs(212));
    layer0_outputs(7915) <= not(inputs(199));
    layer0_outputs(7916) <= not(inputs(251)) or (inputs(181));
    layer0_outputs(7917) <= (inputs(80)) or (inputs(86));
    layer0_outputs(7918) <= not(inputs(20));
    layer0_outputs(7919) <= not(inputs(186));
    layer0_outputs(7920) <= not((inputs(87)) xor (inputs(74)));
    layer0_outputs(7921) <= not(inputs(11));
    layer0_outputs(7922) <= not((inputs(213)) or (inputs(101)));
    layer0_outputs(7923) <= not((inputs(60)) or (inputs(90)));
    layer0_outputs(7924) <= not(inputs(194));
    layer0_outputs(7925) <= not((inputs(67)) xor (inputs(121)));
    layer0_outputs(7926) <= (inputs(162)) or (inputs(79));
    layer0_outputs(7927) <= not((inputs(208)) and (inputs(115)));
    layer0_outputs(7928) <= inputs(10);
    layer0_outputs(7929) <= not(inputs(102)) or (inputs(33));
    layer0_outputs(7930) <= not(inputs(189)) or (inputs(103));
    layer0_outputs(7931) <= not((inputs(22)) and (inputs(60)));
    layer0_outputs(7932) <= (inputs(64)) and not (inputs(7));
    layer0_outputs(7933) <= inputs(234);
    layer0_outputs(7934) <= '1';
    layer0_outputs(7935) <= not((inputs(251)) or (inputs(116)));
    layer0_outputs(7936) <= (inputs(128)) or (inputs(77));
    layer0_outputs(7937) <= not((inputs(158)) or (inputs(100)));
    layer0_outputs(7938) <= (inputs(0)) xor (inputs(213));
    layer0_outputs(7939) <= not((inputs(54)) or (inputs(226)));
    layer0_outputs(7940) <= not(inputs(152)) or (inputs(126));
    layer0_outputs(7941) <= not((inputs(19)) xor (inputs(155)));
    layer0_outputs(7942) <= (inputs(6)) or (inputs(107));
    layer0_outputs(7943) <= not(inputs(72));
    layer0_outputs(7944) <= not((inputs(200)) xor (inputs(8)));
    layer0_outputs(7945) <= (inputs(214)) xor (inputs(216));
    layer0_outputs(7946) <= not((inputs(16)) and (inputs(8)));
    layer0_outputs(7947) <= '1';
    layer0_outputs(7948) <= not(inputs(10)) or (inputs(9));
    layer0_outputs(7949) <= inputs(219);
    layer0_outputs(7950) <= (inputs(235)) or (inputs(197));
    layer0_outputs(7951) <= not(inputs(161)) or (inputs(172));
    layer0_outputs(7952) <= not(inputs(8)) or (inputs(2));
    layer0_outputs(7953) <= not((inputs(152)) or (inputs(207)));
    layer0_outputs(7954) <= inputs(13);
    layer0_outputs(7955) <= (inputs(176)) and not (inputs(221));
    layer0_outputs(7956) <= not((inputs(26)) or (inputs(26)));
    layer0_outputs(7957) <= (inputs(27)) xor (inputs(208));
    layer0_outputs(7958) <= not(inputs(9));
    layer0_outputs(7959) <= (inputs(146)) xor (inputs(132));
    layer0_outputs(7960) <= not(inputs(17));
    layer0_outputs(7961) <= not(inputs(131)) or (inputs(255));
    layer0_outputs(7962) <= (inputs(44)) xor (inputs(204));
    layer0_outputs(7963) <= inputs(70);
    layer0_outputs(7964) <= '0';
    layer0_outputs(7965) <= not(inputs(210)) or (inputs(113));
    layer0_outputs(7966) <= not((inputs(162)) xor (inputs(154)));
    layer0_outputs(7967) <= (inputs(139)) xor (inputs(158));
    layer0_outputs(7968) <= (inputs(146)) xor (inputs(168));
    layer0_outputs(7969) <= not(inputs(240)) or (inputs(242));
    layer0_outputs(7970) <= not((inputs(148)) xor (inputs(133)));
    layer0_outputs(7971) <= (inputs(216)) and not (inputs(141));
    layer0_outputs(7972) <= (inputs(136)) and (inputs(51));
    layer0_outputs(7973) <= inputs(64);
    layer0_outputs(7974) <= not(inputs(211));
    layer0_outputs(7975) <= inputs(39);
    layer0_outputs(7976) <= (inputs(104)) xor (inputs(111));
    layer0_outputs(7977) <= inputs(232);
    layer0_outputs(7978) <= not((inputs(119)) xor (inputs(88)));
    layer0_outputs(7979) <= (inputs(237)) or (inputs(236));
    layer0_outputs(7980) <= (inputs(221)) xor (inputs(100));
    layer0_outputs(7981) <= not((inputs(241)) or (inputs(117)));
    layer0_outputs(7982) <= not((inputs(102)) or (inputs(253)));
    layer0_outputs(7983) <= not(inputs(51));
    layer0_outputs(7984) <= not((inputs(233)) or (inputs(186)));
    layer0_outputs(7985) <= not(inputs(154)) or (inputs(212));
    layer0_outputs(7986) <= (inputs(106)) and not (inputs(190));
    layer0_outputs(7987) <= inputs(178);
    layer0_outputs(7988) <= not(inputs(159)) or (inputs(250));
    layer0_outputs(7989) <= inputs(167);
    layer0_outputs(7990) <= inputs(102);
    layer0_outputs(7991) <= not(inputs(67));
    layer0_outputs(7992) <= not(inputs(98));
    layer0_outputs(7993) <= '1';
    layer0_outputs(7994) <= not((inputs(23)) or (inputs(231)));
    layer0_outputs(7995) <= not(inputs(215));
    layer0_outputs(7996) <= (inputs(191)) or (inputs(253));
    layer0_outputs(7997) <= not(inputs(44));
    layer0_outputs(7998) <= not(inputs(252));
    layer0_outputs(7999) <= not(inputs(25)) or (inputs(119));
    layer0_outputs(8000) <= not(inputs(231)) or (inputs(91));
    layer0_outputs(8001) <= (inputs(176)) or (inputs(186));
    layer0_outputs(8002) <= not(inputs(218));
    layer0_outputs(8003) <= inputs(23);
    layer0_outputs(8004) <= not(inputs(227)) or (inputs(61));
    layer0_outputs(8005) <= inputs(223);
    layer0_outputs(8006) <= inputs(132);
    layer0_outputs(8007) <= not((inputs(209)) or (inputs(14)));
    layer0_outputs(8008) <= not((inputs(36)) xor (inputs(72)));
    layer0_outputs(8009) <= not((inputs(174)) xor (inputs(83)));
    layer0_outputs(8010) <= (inputs(12)) xor (inputs(58));
    layer0_outputs(8011) <= not(inputs(177)) or (inputs(171));
    layer0_outputs(8012) <= (inputs(107)) xor (inputs(11));
    layer0_outputs(8013) <= inputs(202);
    layer0_outputs(8014) <= '1';
    layer0_outputs(8015) <= inputs(229);
    layer0_outputs(8016) <= (inputs(85)) or (inputs(96));
    layer0_outputs(8017) <= (inputs(114)) xor (inputs(230));
    layer0_outputs(8018) <= (inputs(227)) xor (inputs(91));
    layer0_outputs(8019) <= (inputs(248)) xor (inputs(85));
    layer0_outputs(8020) <= (inputs(84)) and not (inputs(33));
    layer0_outputs(8021) <= inputs(22);
    layer0_outputs(8022) <= (inputs(249)) xor (inputs(220));
    layer0_outputs(8023) <= (inputs(212)) xor (inputs(228));
    layer0_outputs(8024) <= inputs(129);
    layer0_outputs(8025) <= not((inputs(80)) or (inputs(69)));
    layer0_outputs(8026) <= (inputs(250)) xor (inputs(95));
    layer0_outputs(8027) <= inputs(149);
    layer0_outputs(8028) <= (inputs(185)) and (inputs(227));
    layer0_outputs(8029) <= not(inputs(219));
    layer0_outputs(8030) <= not((inputs(233)) or (inputs(95)));
    layer0_outputs(8031) <= not(inputs(108));
    layer0_outputs(8032) <= (inputs(135)) xor (inputs(52));
    layer0_outputs(8033) <= (inputs(102)) xor (inputs(131));
    layer0_outputs(8034) <= not((inputs(92)) or (inputs(91)));
    layer0_outputs(8035) <= (inputs(180)) and not (inputs(98));
    layer0_outputs(8036) <= inputs(53);
    layer0_outputs(8037) <= not((inputs(99)) and (inputs(229)));
    layer0_outputs(8038) <= '1';
    layer0_outputs(8039) <= not(inputs(145));
    layer0_outputs(8040) <= not(inputs(180));
    layer0_outputs(8041) <= not(inputs(232));
    layer0_outputs(8042) <= inputs(105);
    layer0_outputs(8043) <= inputs(234);
    layer0_outputs(8044) <= not((inputs(2)) xor (inputs(255)));
    layer0_outputs(8045) <= not(inputs(134)) or (inputs(126));
    layer0_outputs(8046) <= not((inputs(91)) xor (inputs(3)));
    layer0_outputs(8047) <= (inputs(234)) xor (inputs(187));
    layer0_outputs(8048) <= (inputs(192)) or (inputs(146));
    layer0_outputs(8049) <= (inputs(28)) xor (inputs(44));
    layer0_outputs(8050) <= not(inputs(163));
    layer0_outputs(8051) <= not((inputs(67)) or (inputs(47)));
    layer0_outputs(8052) <= not((inputs(203)) xor (inputs(8)));
    layer0_outputs(8053) <= not((inputs(202)) xor (inputs(236)));
    layer0_outputs(8054) <= (inputs(6)) xor (inputs(54));
    layer0_outputs(8055) <= (inputs(166)) and not (inputs(49));
    layer0_outputs(8056) <= (inputs(222)) or (inputs(246));
    layer0_outputs(8057) <= not(inputs(191)) or (inputs(156));
    layer0_outputs(8058) <= inputs(99);
    layer0_outputs(8059) <= (inputs(209)) or (inputs(171));
    layer0_outputs(8060) <= not((inputs(46)) xor (inputs(75)));
    layer0_outputs(8061) <= (inputs(167)) and not (inputs(76));
    layer0_outputs(8062) <= (inputs(26)) and not (inputs(13));
    layer0_outputs(8063) <= not(inputs(18));
    layer0_outputs(8064) <= inputs(210);
    layer0_outputs(8065) <= (inputs(1)) or (inputs(189));
    layer0_outputs(8066) <= not(inputs(196));
    layer0_outputs(8067) <= (inputs(198)) xor (inputs(233));
    layer0_outputs(8068) <= '0';
    layer0_outputs(8069) <= (inputs(106)) and not (inputs(189));
    layer0_outputs(8070) <= (inputs(197)) and not (inputs(219));
    layer0_outputs(8071) <= (inputs(18)) xor (inputs(46));
    layer0_outputs(8072) <= inputs(122);
    layer0_outputs(8073) <= not((inputs(110)) or (inputs(84)));
    layer0_outputs(8074) <= (inputs(146)) and not (inputs(236));
    layer0_outputs(8075) <= (inputs(17)) and (inputs(174));
    layer0_outputs(8076) <= not(inputs(43));
    layer0_outputs(8077) <= not((inputs(32)) or (inputs(151)));
    layer0_outputs(8078) <= not((inputs(235)) xor (inputs(188)));
    layer0_outputs(8079) <= (inputs(17)) xor (inputs(184));
    layer0_outputs(8080) <= not((inputs(96)) xor (inputs(165)));
    layer0_outputs(8081) <= not(inputs(162)) or (inputs(77));
    layer0_outputs(8082) <= (inputs(254)) or (inputs(165));
    layer0_outputs(8083) <= (inputs(19)) xor (inputs(122));
    layer0_outputs(8084) <= inputs(145);
    layer0_outputs(8085) <= not(inputs(131));
    layer0_outputs(8086) <= not(inputs(67));
    layer0_outputs(8087) <= not((inputs(120)) xor (inputs(195)));
    layer0_outputs(8088) <= inputs(79);
    layer0_outputs(8089) <= not((inputs(76)) xor (inputs(10)));
    layer0_outputs(8090) <= not((inputs(46)) or (inputs(102)));
    layer0_outputs(8091) <= (inputs(133)) and (inputs(33));
    layer0_outputs(8092) <= not(inputs(203));
    layer0_outputs(8093) <= not((inputs(133)) and (inputs(227)));
    layer0_outputs(8094) <= not(inputs(249));
    layer0_outputs(8095) <= not(inputs(198)) or (inputs(111));
    layer0_outputs(8096) <= not(inputs(141)) or (inputs(253));
    layer0_outputs(8097) <= (inputs(87)) and not (inputs(254));
    layer0_outputs(8098) <= not((inputs(95)) xor (inputs(40)));
    layer0_outputs(8099) <= (inputs(195)) xor (inputs(120));
    layer0_outputs(8100) <= inputs(116);
    layer0_outputs(8101) <= not(inputs(118)) or (inputs(49));
    layer0_outputs(8102) <= (inputs(206)) xor (inputs(146));
    layer0_outputs(8103) <= inputs(61);
    layer0_outputs(8104) <= not(inputs(75));
    layer0_outputs(8105) <= (inputs(250)) or (inputs(147));
    layer0_outputs(8106) <= not((inputs(193)) and (inputs(135)));
    layer0_outputs(8107) <= not(inputs(190));
    layer0_outputs(8108) <= not((inputs(12)) and (inputs(121)));
    layer0_outputs(8109) <= inputs(105);
    layer0_outputs(8110) <= not(inputs(211));
    layer0_outputs(8111) <= (inputs(158)) xor (inputs(237));
    layer0_outputs(8112) <= not(inputs(17));
    layer0_outputs(8113) <= inputs(97);
    layer0_outputs(8114) <= inputs(225);
    layer0_outputs(8115) <= not((inputs(179)) xor (inputs(72)));
    layer0_outputs(8116) <= (inputs(170)) and not (inputs(160));
    layer0_outputs(8117) <= (inputs(118)) xor (inputs(183));
    layer0_outputs(8118) <= not(inputs(164));
    layer0_outputs(8119) <= (inputs(169)) xor (inputs(180));
    layer0_outputs(8120) <= inputs(187);
    layer0_outputs(8121) <= not(inputs(73));
    layer0_outputs(8122) <= not(inputs(38)) or (inputs(85));
    layer0_outputs(8123) <= not(inputs(181));
    layer0_outputs(8124) <= (inputs(20)) and (inputs(40));
    layer0_outputs(8125) <= not(inputs(112));
    layer0_outputs(8126) <= not((inputs(17)) or (inputs(36)));
    layer0_outputs(8127) <= (inputs(195)) and (inputs(76));
    layer0_outputs(8128) <= not(inputs(174));
    layer0_outputs(8129) <= not((inputs(238)) xor (inputs(34)));
    layer0_outputs(8130) <= (inputs(173)) or (inputs(43));
    layer0_outputs(8131) <= inputs(87);
    layer0_outputs(8132) <= inputs(107);
    layer0_outputs(8133) <= not(inputs(91));
    layer0_outputs(8134) <= (inputs(148)) and not (inputs(28));
    layer0_outputs(8135) <= (inputs(35)) xor (inputs(114));
    layer0_outputs(8136) <= not(inputs(137));
    layer0_outputs(8137) <= (inputs(90)) or (inputs(182));
    layer0_outputs(8138) <= (inputs(152)) and not (inputs(239));
    layer0_outputs(8139) <= inputs(89);
    layer0_outputs(8140) <= inputs(139);
    layer0_outputs(8141) <= not(inputs(177));
    layer0_outputs(8142) <= inputs(107);
    layer0_outputs(8143) <= inputs(209);
    layer0_outputs(8144) <= inputs(194);
    layer0_outputs(8145) <= (inputs(69)) and not (inputs(191));
    layer0_outputs(8146) <= not(inputs(244)) or (inputs(1));
    layer0_outputs(8147) <= not((inputs(106)) xor (inputs(141)));
    layer0_outputs(8148) <= not(inputs(109)) or (inputs(237));
    layer0_outputs(8149) <= (inputs(182)) and not (inputs(235));
    layer0_outputs(8150) <= not((inputs(95)) xor (inputs(104)));
    layer0_outputs(8151) <= '1';
    layer0_outputs(8152) <= (inputs(84)) and not (inputs(144));
    layer0_outputs(8153) <= (inputs(228)) and not (inputs(64));
    layer0_outputs(8154) <= inputs(163);
    layer0_outputs(8155) <= (inputs(182)) and (inputs(247));
    layer0_outputs(8156) <= (inputs(46)) or (inputs(84));
    layer0_outputs(8157) <= not((inputs(147)) or (inputs(225)));
    layer0_outputs(8158) <= inputs(34);
    layer0_outputs(8159) <= (inputs(152)) and not (inputs(204));
    layer0_outputs(8160) <= (inputs(6)) xor (inputs(158));
    layer0_outputs(8161) <= not(inputs(110)) or (inputs(0));
    layer0_outputs(8162) <= (inputs(254)) or (inputs(121));
    layer0_outputs(8163) <= not(inputs(227));
    layer0_outputs(8164) <= not((inputs(163)) or (inputs(201)));
    layer0_outputs(8165) <= not(inputs(124)) or (inputs(20));
    layer0_outputs(8166) <= not(inputs(126));
    layer0_outputs(8167) <= (inputs(191)) xor (inputs(95));
    layer0_outputs(8168) <= (inputs(53)) or (inputs(173));
    layer0_outputs(8169) <= not((inputs(166)) or (inputs(248)));
    layer0_outputs(8170) <= not((inputs(147)) and (inputs(147)));
    layer0_outputs(8171) <= not((inputs(48)) xor (inputs(25)));
    layer0_outputs(8172) <= (inputs(109)) or (inputs(36));
    layer0_outputs(8173) <= inputs(164);
    layer0_outputs(8174) <= inputs(102);
    layer0_outputs(8175) <= not(inputs(89));
    layer0_outputs(8176) <= not(inputs(41)) or (inputs(207));
    layer0_outputs(8177) <= (inputs(76)) xor (inputs(72));
    layer0_outputs(8178) <= inputs(230);
    layer0_outputs(8179) <= (inputs(7)) xor (inputs(52));
    layer0_outputs(8180) <= not((inputs(0)) xor (inputs(125)));
    layer0_outputs(8181) <= not(inputs(231));
    layer0_outputs(8182) <= not((inputs(44)) and (inputs(105)));
    layer0_outputs(8183) <= (inputs(230)) and not (inputs(255));
    layer0_outputs(8184) <= (inputs(112)) and not (inputs(192));
    layer0_outputs(8185) <= not(inputs(23));
    layer0_outputs(8186) <= (inputs(123)) or (inputs(167));
    layer0_outputs(8187) <= (inputs(9)) or (inputs(236));
    layer0_outputs(8188) <= not(inputs(60)) or (inputs(97));
    layer0_outputs(8189) <= not(inputs(93));
    layer0_outputs(8190) <= (inputs(214)) or (inputs(233));
    layer0_outputs(8191) <= not((inputs(233)) xor (inputs(245)));
    layer0_outputs(8192) <= not((inputs(93)) or (inputs(21)));
    layer0_outputs(8193) <= (inputs(118)) xor (inputs(72));
    layer0_outputs(8194) <= (inputs(243)) or (inputs(149));
    layer0_outputs(8195) <= not(inputs(121));
    layer0_outputs(8196) <= inputs(219);
    layer0_outputs(8197) <= (inputs(13)) xor (inputs(30));
    layer0_outputs(8198) <= '0';
    layer0_outputs(8199) <= not(inputs(198));
    layer0_outputs(8200) <= (inputs(89)) xor (inputs(38));
    layer0_outputs(8201) <= inputs(210);
    layer0_outputs(8202) <= inputs(171);
    layer0_outputs(8203) <= '1';
    layer0_outputs(8204) <= (inputs(177)) and not (inputs(107));
    layer0_outputs(8205) <= inputs(100);
    layer0_outputs(8206) <= not(inputs(230));
    layer0_outputs(8207) <= not(inputs(94));
    layer0_outputs(8208) <= '0';
    layer0_outputs(8209) <= not((inputs(162)) or (inputs(185)));
    layer0_outputs(8210) <= not(inputs(216)) or (inputs(20));
    layer0_outputs(8211) <= not((inputs(106)) or (inputs(137)));
    layer0_outputs(8212) <= (inputs(109)) xor (inputs(95));
    layer0_outputs(8213) <= inputs(76);
    layer0_outputs(8214) <= not(inputs(209));
    layer0_outputs(8215) <= '1';
    layer0_outputs(8216) <= not((inputs(190)) or (inputs(215)));
    layer0_outputs(8217) <= (inputs(93)) xor (inputs(76));
    layer0_outputs(8218) <= (inputs(178)) and not (inputs(170));
    layer0_outputs(8219) <= (inputs(115)) xor (inputs(85));
    layer0_outputs(8220) <= inputs(121);
    layer0_outputs(8221) <= not((inputs(100)) xor (inputs(10)));
    layer0_outputs(8222) <= not((inputs(164)) or (inputs(65)));
    layer0_outputs(8223) <= not(inputs(133)) or (inputs(18));
    layer0_outputs(8224) <= not(inputs(155)) or (inputs(224));
    layer0_outputs(8225) <= (inputs(27)) and not (inputs(239));
    layer0_outputs(8226) <= (inputs(91)) and not (inputs(232));
    layer0_outputs(8227) <= (inputs(85)) or (inputs(48));
    layer0_outputs(8228) <= (inputs(108)) or (inputs(121));
    layer0_outputs(8229) <= (inputs(35)) or (inputs(213));
    layer0_outputs(8230) <= (inputs(158)) or (inputs(68));
    layer0_outputs(8231) <= (inputs(226)) or (inputs(190));
    layer0_outputs(8232) <= (inputs(97)) or (inputs(52));
    layer0_outputs(8233) <= (inputs(82)) or (inputs(212));
    layer0_outputs(8234) <= not((inputs(48)) or (inputs(65)));
    layer0_outputs(8235) <= (inputs(151)) and not (inputs(31));
    layer0_outputs(8236) <= not((inputs(200)) or (inputs(225)));
    layer0_outputs(8237) <= not(inputs(145)) or (inputs(191));
    layer0_outputs(8238) <= not((inputs(212)) or (inputs(214)));
    layer0_outputs(8239) <= not((inputs(3)) or (inputs(30)));
    layer0_outputs(8240) <= (inputs(83)) and not (inputs(127));
    layer0_outputs(8241) <= not(inputs(27)) or (inputs(245));
    layer0_outputs(8242) <= not(inputs(104));
    layer0_outputs(8243) <= (inputs(46)) xor (inputs(242));
    layer0_outputs(8244) <= not(inputs(16));
    layer0_outputs(8245) <= not(inputs(205));
    layer0_outputs(8246) <= (inputs(232)) and not (inputs(155));
    layer0_outputs(8247) <= not(inputs(230));
    layer0_outputs(8248) <= not((inputs(79)) or (inputs(26)));
    layer0_outputs(8249) <= (inputs(88)) and not (inputs(219));
    layer0_outputs(8250) <= not((inputs(180)) or (inputs(232)));
    layer0_outputs(8251) <= (inputs(143)) or (inputs(46));
    layer0_outputs(8252) <= (inputs(210)) or (inputs(223));
    layer0_outputs(8253) <= not(inputs(92)) or (inputs(252));
    layer0_outputs(8254) <= not(inputs(61)) or (inputs(240));
    layer0_outputs(8255) <= (inputs(154)) and not (inputs(223));
    layer0_outputs(8256) <= not((inputs(77)) xor (inputs(60)));
    layer0_outputs(8257) <= (inputs(89)) xor (inputs(23));
    layer0_outputs(8258) <= not(inputs(10));
    layer0_outputs(8259) <= not((inputs(64)) or (inputs(32)));
    layer0_outputs(8260) <= not(inputs(200)) or (inputs(196));
    layer0_outputs(8261) <= (inputs(218)) and not (inputs(30));
    layer0_outputs(8262) <= (inputs(115)) or (inputs(236));
    layer0_outputs(8263) <= not(inputs(156)) or (inputs(213));
    layer0_outputs(8264) <= not(inputs(90));
    layer0_outputs(8265) <= not(inputs(9));
    layer0_outputs(8266) <= (inputs(140)) xor (inputs(251));
    layer0_outputs(8267) <= not((inputs(48)) and (inputs(48)));
    layer0_outputs(8268) <= (inputs(102)) or (inputs(58));
    layer0_outputs(8269) <= not(inputs(24));
    layer0_outputs(8270) <= not((inputs(21)) or (inputs(110)));
    layer0_outputs(8271) <= inputs(25);
    layer0_outputs(8272) <= inputs(88);
    layer0_outputs(8273) <= not((inputs(160)) xor (inputs(247)));
    layer0_outputs(8274) <= not(inputs(121)) or (inputs(193));
    layer0_outputs(8275) <= not(inputs(162)) or (inputs(110));
    layer0_outputs(8276) <= inputs(101);
    layer0_outputs(8277) <= (inputs(47)) and not (inputs(169));
    layer0_outputs(8278) <= not(inputs(232));
    layer0_outputs(8279) <= (inputs(34)) xor (inputs(85));
    layer0_outputs(8280) <= not((inputs(2)) and (inputs(25)));
    layer0_outputs(8281) <= inputs(101);
    layer0_outputs(8282) <= not(inputs(11)) or (inputs(183));
    layer0_outputs(8283) <= inputs(119);
    layer0_outputs(8284) <= (inputs(34)) or (inputs(89));
    layer0_outputs(8285) <= (inputs(24)) and not (inputs(122));
    layer0_outputs(8286) <= (inputs(161)) or (inputs(102));
    layer0_outputs(8287) <= not((inputs(42)) xor (inputs(249)));
    layer0_outputs(8288) <= (inputs(150)) and not (inputs(79));
    layer0_outputs(8289) <= not(inputs(122));
    layer0_outputs(8290) <= (inputs(59)) xor (inputs(93));
    layer0_outputs(8291) <= '0';
    layer0_outputs(8292) <= not(inputs(243)) or (inputs(125));
    layer0_outputs(8293) <= '0';
    layer0_outputs(8294) <= not((inputs(123)) or (inputs(22)));
    layer0_outputs(8295) <= not(inputs(235));
    layer0_outputs(8296) <= not((inputs(161)) xor (inputs(193)));
    layer0_outputs(8297) <= (inputs(135)) and not (inputs(41));
    layer0_outputs(8298) <= (inputs(73)) xor (inputs(76));
    layer0_outputs(8299) <= (inputs(164)) and not (inputs(123));
    layer0_outputs(8300) <= not((inputs(160)) or (inputs(58)));
    layer0_outputs(8301) <= (inputs(36)) or (inputs(21));
    layer0_outputs(8302) <= not(inputs(114));
    layer0_outputs(8303) <= inputs(167);
    layer0_outputs(8304) <= not((inputs(24)) and (inputs(104)));
    layer0_outputs(8305) <= not(inputs(18));
    layer0_outputs(8306) <= not(inputs(180));
    layer0_outputs(8307) <= (inputs(231)) and not (inputs(112));
    layer0_outputs(8308) <= (inputs(168)) and not (inputs(173));
    layer0_outputs(8309) <= not((inputs(226)) and (inputs(28)));
    layer0_outputs(8310) <= not(inputs(158));
    layer0_outputs(8311) <= (inputs(184)) xor (inputs(3));
    layer0_outputs(8312) <= (inputs(229)) and not (inputs(143));
    layer0_outputs(8313) <= (inputs(153)) and not (inputs(26));
    layer0_outputs(8314) <= (inputs(114)) xor (inputs(56));
    layer0_outputs(8315) <= (inputs(74)) xor (inputs(137));
    layer0_outputs(8316) <= not(inputs(159)) or (inputs(240));
    layer0_outputs(8317) <= not(inputs(159));
    layer0_outputs(8318) <= '1';
    layer0_outputs(8319) <= not(inputs(131));
    layer0_outputs(8320) <= not((inputs(180)) or (inputs(234)));
    layer0_outputs(8321) <= inputs(87);
    layer0_outputs(8322) <= (inputs(232)) xor (inputs(186));
    layer0_outputs(8323) <= (inputs(238)) or (inputs(65));
    layer0_outputs(8324) <= not((inputs(150)) xor (inputs(243)));
    layer0_outputs(8325) <= not(inputs(109));
    layer0_outputs(8326) <= (inputs(29)) and (inputs(20));
    layer0_outputs(8327) <= not((inputs(0)) xor (inputs(220)));
    layer0_outputs(8328) <= not((inputs(86)) or (inputs(188)));
    layer0_outputs(8329) <= inputs(218);
    layer0_outputs(8330) <= not(inputs(229));
    layer0_outputs(8331) <= not(inputs(14));
    layer0_outputs(8332) <= inputs(145);
    layer0_outputs(8333) <= (inputs(86)) xor (inputs(158));
    layer0_outputs(8334) <= (inputs(140)) or (inputs(125));
    layer0_outputs(8335) <= (inputs(36)) or (inputs(247));
    layer0_outputs(8336) <= (inputs(68)) xor (inputs(64));
    layer0_outputs(8337) <= inputs(60);
    layer0_outputs(8338) <= inputs(82);
    layer0_outputs(8339) <= (inputs(38)) or (inputs(20));
    layer0_outputs(8340) <= not(inputs(174)) or (inputs(181));
    layer0_outputs(8341) <= (inputs(119)) or (inputs(225));
    layer0_outputs(8342) <= (inputs(56)) or (inputs(177));
    layer0_outputs(8343) <= not((inputs(103)) and (inputs(67)));
    layer0_outputs(8344) <= (inputs(171)) xor (inputs(250));
    layer0_outputs(8345) <= not((inputs(79)) or (inputs(55)));
    layer0_outputs(8346) <= inputs(82);
    layer0_outputs(8347) <= not(inputs(147)) or (inputs(189));
    layer0_outputs(8348) <= (inputs(92)) or (inputs(89));
    layer0_outputs(8349) <= inputs(37);
    layer0_outputs(8350) <= (inputs(46)) and not (inputs(223));
    layer0_outputs(8351) <= (inputs(253)) or (inputs(93));
    layer0_outputs(8352) <= not(inputs(186));
    layer0_outputs(8353) <= (inputs(81)) and not (inputs(154));
    layer0_outputs(8354) <= not(inputs(196)) or (inputs(185));
    layer0_outputs(8355) <= not((inputs(69)) or (inputs(36)));
    layer0_outputs(8356) <= not((inputs(5)) xor (inputs(177)));
    layer0_outputs(8357) <= not((inputs(118)) xor (inputs(179)));
    layer0_outputs(8358) <= (inputs(116)) or (inputs(17));
    layer0_outputs(8359) <= (inputs(107)) and not (inputs(173));
    layer0_outputs(8360) <= not(inputs(71));
    layer0_outputs(8361) <= not(inputs(197));
    layer0_outputs(8362) <= not(inputs(179));
    layer0_outputs(8363) <= (inputs(20)) xor (inputs(30));
    layer0_outputs(8364) <= (inputs(45)) xor (inputs(26));
    layer0_outputs(8365) <= (inputs(216)) and not (inputs(45));
    layer0_outputs(8366) <= '0';
    layer0_outputs(8367) <= not((inputs(59)) or (inputs(3)));
    layer0_outputs(8368) <= inputs(168);
    layer0_outputs(8369) <= not(inputs(134));
    layer0_outputs(8370) <= not(inputs(178)) or (inputs(18));
    layer0_outputs(8371) <= inputs(76);
    layer0_outputs(8372) <= not((inputs(6)) or (inputs(94)));
    layer0_outputs(8373) <= not(inputs(36));
    layer0_outputs(8374) <= (inputs(185)) or (inputs(199));
    layer0_outputs(8375) <= not((inputs(178)) xor (inputs(155)));
    layer0_outputs(8376) <= (inputs(182)) xor (inputs(61));
    layer0_outputs(8377) <= (inputs(216)) or (inputs(35));
    layer0_outputs(8378) <= (inputs(23)) xor (inputs(53));
    layer0_outputs(8379) <= not(inputs(53)) or (inputs(63));
    layer0_outputs(8380) <= not(inputs(33)) or (inputs(110));
    layer0_outputs(8381) <= (inputs(226)) or (inputs(202));
    layer0_outputs(8382) <= not(inputs(42));
    layer0_outputs(8383) <= not((inputs(121)) or (inputs(79)));
    layer0_outputs(8384) <= not(inputs(195)) or (inputs(29));
    layer0_outputs(8385) <= (inputs(35)) and (inputs(204));
    layer0_outputs(8386) <= inputs(160);
    layer0_outputs(8387) <= not(inputs(42)) or (inputs(34));
    layer0_outputs(8388) <= (inputs(136)) or (inputs(248));
    layer0_outputs(8389) <= not((inputs(225)) xor (inputs(181)));
    layer0_outputs(8390) <= inputs(217);
    layer0_outputs(8391) <= (inputs(5)) or (inputs(38));
    layer0_outputs(8392) <= not(inputs(210)) or (inputs(174));
    layer0_outputs(8393) <= inputs(247);
    layer0_outputs(8394) <= not(inputs(234)) or (inputs(65));
    layer0_outputs(8395) <= not((inputs(11)) xor (inputs(160)));
    layer0_outputs(8396) <= (inputs(63)) or (inputs(71));
    layer0_outputs(8397) <= not((inputs(204)) or (inputs(64)));
    layer0_outputs(8398) <= (inputs(83)) or (inputs(182));
    layer0_outputs(8399) <= inputs(75);
    layer0_outputs(8400) <= (inputs(109)) or (inputs(125));
    layer0_outputs(8401) <= inputs(108);
    layer0_outputs(8402) <= (inputs(156)) or (inputs(21));
    layer0_outputs(8403) <= inputs(129);
    layer0_outputs(8404) <= (inputs(103)) xor (inputs(46));
    layer0_outputs(8405) <= not((inputs(4)) xor (inputs(160)));
    layer0_outputs(8406) <= inputs(127);
    layer0_outputs(8407) <= not((inputs(123)) or (inputs(115)));
    layer0_outputs(8408) <= not((inputs(172)) xor (inputs(244)));
    layer0_outputs(8409) <= not((inputs(195)) xor (inputs(250)));
    layer0_outputs(8410) <= not(inputs(42)) or (inputs(114));
    layer0_outputs(8411) <= not((inputs(233)) xor (inputs(161)));
    layer0_outputs(8412) <= (inputs(203)) and not (inputs(253));
    layer0_outputs(8413) <= not((inputs(246)) or (inputs(49)));
    layer0_outputs(8414) <= (inputs(163)) or (inputs(223));
    layer0_outputs(8415) <= (inputs(222)) or (inputs(63));
    layer0_outputs(8416) <= not((inputs(41)) or (inputs(110)));
    layer0_outputs(8417) <= not(inputs(167));
    layer0_outputs(8418) <= (inputs(8)) xor (inputs(111));
    layer0_outputs(8419) <= not((inputs(208)) xor (inputs(184)));
    layer0_outputs(8420) <= inputs(192);
    layer0_outputs(8421) <= not((inputs(183)) xor (inputs(193)));
    layer0_outputs(8422) <= not(inputs(97));
    layer0_outputs(8423) <= not((inputs(120)) xor (inputs(164)));
    layer0_outputs(8424) <= not(inputs(147));
    layer0_outputs(8425) <= (inputs(142)) xor (inputs(103));
    layer0_outputs(8426) <= not(inputs(163));
    layer0_outputs(8427) <= (inputs(186)) or (inputs(52));
    layer0_outputs(8428) <= not((inputs(2)) xor (inputs(237)));
    layer0_outputs(8429) <= inputs(70);
    layer0_outputs(8430) <= not(inputs(114));
    layer0_outputs(8431) <= not(inputs(206));
    layer0_outputs(8432) <= not((inputs(21)) or (inputs(94)));
    layer0_outputs(8433) <= (inputs(70)) or (inputs(149));
    layer0_outputs(8434) <= inputs(19);
    layer0_outputs(8435) <= inputs(83);
    layer0_outputs(8436) <= not((inputs(206)) or (inputs(76)));
    layer0_outputs(8437) <= (inputs(22)) and not (inputs(165));
    layer0_outputs(8438) <= (inputs(229)) and (inputs(105));
    layer0_outputs(8439) <= not(inputs(62));
    layer0_outputs(8440) <= not(inputs(115));
    layer0_outputs(8441) <= not((inputs(250)) or (inputs(161)));
    layer0_outputs(8442) <= not((inputs(250)) xor (inputs(42)));
    layer0_outputs(8443) <= (inputs(228)) xor (inputs(109));
    layer0_outputs(8444) <= '1';
    layer0_outputs(8445) <= (inputs(13)) and not (inputs(208));
    layer0_outputs(8446) <= not(inputs(213)) or (inputs(65));
    layer0_outputs(8447) <= inputs(99);
    layer0_outputs(8448) <= not((inputs(146)) xor (inputs(206)));
    layer0_outputs(8449) <= not((inputs(208)) xor (inputs(100)));
    layer0_outputs(8450) <= not((inputs(95)) xor (inputs(203)));
    layer0_outputs(8451) <= not(inputs(24));
    layer0_outputs(8452) <= not(inputs(234)) or (inputs(76));
    layer0_outputs(8453) <= not(inputs(117)) or (inputs(75));
    layer0_outputs(8454) <= not((inputs(121)) and (inputs(71)));
    layer0_outputs(8455) <= (inputs(238)) or (inputs(66));
    layer0_outputs(8456) <= (inputs(144)) and not (inputs(216));
    layer0_outputs(8457) <= (inputs(102)) and not (inputs(155));
    layer0_outputs(8458) <= (inputs(154)) xor (inputs(201));
    layer0_outputs(8459) <= (inputs(86)) xor (inputs(188));
    layer0_outputs(8460) <= not((inputs(212)) xor (inputs(65)));
    layer0_outputs(8461) <= (inputs(60)) and (inputs(41));
    layer0_outputs(8462) <= not((inputs(196)) or (inputs(16)));
    layer0_outputs(8463) <= not(inputs(133));
    layer0_outputs(8464) <= inputs(135);
    layer0_outputs(8465) <= inputs(130);
    layer0_outputs(8466) <= not(inputs(212)) or (inputs(63));
    layer0_outputs(8467) <= not((inputs(203)) or (inputs(164)));
    layer0_outputs(8468) <= not(inputs(52)) or (inputs(215));
    layer0_outputs(8469) <= (inputs(105)) xor (inputs(75));
    layer0_outputs(8470) <= inputs(144);
    layer0_outputs(8471) <= not((inputs(232)) xor (inputs(109)));
    layer0_outputs(8472) <= not((inputs(88)) or (inputs(213)));
    layer0_outputs(8473) <= inputs(81);
    layer0_outputs(8474) <= (inputs(172)) xor (inputs(170));
    layer0_outputs(8475) <= inputs(71);
    layer0_outputs(8476) <= not(inputs(244)) or (inputs(3));
    layer0_outputs(8477) <= not((inputs(148)) or (inputs(220)));
    layer0_outputs(8478) <= not((inputs(245)) xor (inputs(156)));
    layer0_outputs(8479) <= inputs(195);
    layer0_outputs(8480) <= inputs(236);
    layer0_outputs(8481) <= (inputs(162)) xor (inputs(196));
    layer0_outputs(8482) <= not((inputs(109)) xor (inputs(91)));
    layer0_outputs(8483) <= (inputs(118)) and not (inputs(127));
    layer0_outputs(8484) <= inputs(193);
    layer0_outputs(8485) <= inputs(157);
    layer0_outputs(8486) <= not(inputs(38)) or (inputs(139));
    layer0_outputs(8487) <= not(inputs(133));
    layer0_outputs(8488) <= (inputs(212)) and (inputs(164));
    layer0_outputs(8489) <= (inputs(25)) xor (inputs(68));
    layer0_outputs(8490) <= (inputs(147)) xor (inputs(68));
    layer0_outputs(8491) <= '1';
    layer0_outputs(8492) <= not((inputs(108)) xor (inputs(82)));
    layer0_outputs(8493) <= not(inputs(184)) or (inputs(29));
    layer0_outputs(8494) <= inputs(104);
    layer0_outputs(8495) <= (inputs(135)) and not (inputs(159));
    layer0_outputs(8496) <= not((inputs(49)) xor (inputs(25)));
    layer0_outputs(8497) <= not(inputs(82));
    layer0_outputs(8498) <= not(inputs(211));
    layer0_outputs(8499) <= (inputs(64)) or (inputs(172));
    layer0_outputs(8500) <= not(inputs(174)) or (inputs(170));
    layer0_outputs(8501) <= not((inputs(68)) or (inputs(76)));
    layer0_outputs(8502) <= not(inputs(8));
    layer0_outputs(8503) <= (inputs(45)) and not (inputs(136));
    layer0_outputs(8504) <= '0';
    layer0_outputs(8505) <= not(inputs(7)) or (inputs(128));
    layer0_outputs(8506) <= (inputs(100)) xor (inputs(119));
    layer0_outputs(8507) <= inputs(130);
    layer0_outputs(8508) <= not((inputs(176)) or (inputs(242)));
    layer0_outputs(8509) <= not(inputs(42));
    layer0_outputs(8510) <= not(inputs(120)) or (inputs(39));
    layer0_outputs(8511) <= not(inputs(113));
    layer0_outputs(8512) <= (inputs(45)) or (inputs(59));
    layer0_outputs(8513) <= inputs(212);
    layer0_outputs(8514) <= inputs(11);
    layer0_outputs(8515) <= (inputs(176)) or (inputs(73));
    layer0_outputs(8516) <= not(inputs(45));
    layer0_outputs(8517) <= not(inputs(75));
    layer0_outputs(8518) <= not(inputs(145));
    layer0_outputs(8519) <= not(inputs(178)) or (inputs(37));
    layer0_outputs(8520) <= (inputs(90)) xor (inputs(237));
    layer0_outputs(8521) <= not((inputs(201)) or (inputs(80)));
    layer0_outputs(8522) <= not(inputs(63));
    layer0_outputs(8523) <= inputs(189);
    layer0_outputs(8524) <= not(inputs(229));
    layer0_outputs(8525) <= (inputs(112)) or (inputs(205));
    layer0_outputs(8526) <= (inputs(171)) and not (inputs(110));
    layer0_outputs(8527) <= not((inputs(48)) xor (inputs(250)));
    layer0_outputs(8528) <= not(inputs(172)) or (inputs(42));
    layer0_outputs(8529) <= not(inputs(76));
    layer0_outputs(8530) <= not(inputs(44));
    layer0_outputs(8531) <= not(inputs(149)) or (inputs(181));
    layer0_outputs(8532) <= not((inputs(54)) xor (inputs(42)));
    layer0_outputs(8533) <= not(inputs(155));
    layer0_outputs(8534) <= not((inputs(154)) and (inputs(11)));
    layer0_outputs(8535) <= not((inputs(65)) xor (inputs(24)));
    layer0_outputs(8536) <= (inputs(161)) xor (inputs(115));
    layer0_outputs(8537) <= not(inputs(63)) or (inputs(241));
    layer0_outputs(8538) <= (inputs(114)) xor (inputs(133));
    layer0_outputs(8539) <= not(inputs(22)) or (inputs(243));
    layer0_outputs(8540) <= not(inputs(29));
    layer0_outputs(8541) <= (inputs(49)) and not (inputs(239));
    layer0_outputs(8542) <= (inputs(103)) and not (inputs(91));
    layer0_outputs(8543) <= inputs(162);
    layer0_outputs(8544) <= not((inputs(52)) xor (inputs(73)));
    layer0_outputs(8545) <= not((inputs(255)) or (inputs(14)));
    layer0_outputs(8546) <= inputs(10);
    layer0_outputs(8547) <= (inputs(202)) or (inputs(185));
    layer0_outputs(8548) <= (inputs(5)) and not (inputs(97));
    layer0_outputs(8549) <= inputs(46);
    layer0_outputs(8550) <= not(inputs(227));
    layer0_outputs(8551) <= (inputs(161)) or (inputs(36));
    layer0_outputs(8552) <= (inputs(32)) or (inputs(124));
    layer0_outputs(8553) <= not(inputs(67)) or (inputs(149));
    layer0_outputs(8554) <= inputs(124);
    layer0_outputs(8555) <= not(inputs(37)) or (inputs(118));
    layer0_outputs(8556) <= not(inputs(233)) or (inputs(15));
    layer0_outputs(8557) <= (inputs(183)) xor (inputs(210));
    layer0_outputs(8558) <= not(inputs(223));
    layer0_outputs(8559) <= (inputs(194)) and not (inputs(110));
    layer0_outputs(8560) <= inputs(188);
    layer0_outputs(8561) <= (inputs(64)) xor (inputs(222));
    layer0_outputs(8562) <= not(inputs(57)) or (inputs(172));
    layer0_outputs(8563) <= (inputs(16)) xor (inputs(63));
    layer0_outputs(8564) <= not(inputs(231)) or (inputs(253));
    layer0_outputs(8565) <= not((inputs(127)) or (inputs(223)));
    layer0_outputs(8566) <= inputs(153);
    layer0_outputs(8567) <= not((inputs(18)) and (inputs(175)));
    layer0_outputs(8568) <= not(inputs(46));
    layer0_outputs(8569) <= (inputs(176)) xor (inputs(233));
    layer0_outputs(8570) <= (inputs(54)) or (inputs(40));
    layer0_outputs(8571) <= not(inputs(23)) or (inputs(246));
    layer0_outputs(8572) <= inputs(7);
    layer0_outputs(8573) <= (inputs(6)) and not (inputs(126));
    layer0_outputs(8574) <= (inputs(172)) xor (inputs(228));
    layer0_outputs(8575) <= not(inputs(210));
    layer0_outputs(8576) <= not((inputs(110)) or (inputs(71)));
    layer0_outputs(8577) <= not(inputs(116)) or (inputs(140));
    layer0_outputs(8578) <= not((inputs(165)) or (inputs(87)));
    layer0_outputs(8579) <= inputs(117);
    layer0_outputs(8580) <= not(inputs(114)) or (inputs(141));
    layer0_outputs(8581) <= not(inputs(139));
    layer0_outputs(8582) <= not(inputs(254));
    layer0_outputs(8583) <= not(inputs(232)) or (inputs(96));
    layer0_outputs(8584) <= not(inputs(240)) or (inputs(31));
    layer0_outputs(8585) <= (inputs(75)) and (inputs(105));
    layer0_outputs(8586) <= inputs(81);
    layer0_outputs(8587) <= not((inputs(34)) xor (inputs(26)));
    layer0_outputs(8588) <= not(inputs(28)) or (inputs(81));
    layer0_outputs(8589) <= (inputs(98)) xor (inputs(22));
    layer0_outputs(8590) <= not((inputs(254)) or (inputs(73)));
    layer0_outputs(8591) <= (inputs(220)) xor (inputs(121));
    layer0_outputs(8592) <= not(inputs(10));
    layer0_outputs(8593) <= not((inputs(177)) or (inputs(48)));
    layer0_outputs(8594) <= not(inputs(85));
    layer0_outputs(8595) <= not(inputs(93));
    layer0_outputs(8596) <= inputs(187);
    layer0_outputs(8597) <= (inputs(247)) xor (inputs(238));
    layer0_outputs(8598) <= not(inputs(174));
    layer0_outputs(8599) <= not(inputs(134)) or (inputs(126));
    layer0_outputs(8600) <= (inputs(229)) and not (inputs(165));
    layer0_outputs(8601) <= not(inputs(51)) or (inputs(204));
    layer0_outputs(8602) <= (inputs(68)) or (inputs(202));
    layer0_outputs(8603) <= not((inputs(143)) or (inputs(204)));
    layer0_outputs(8604) <= (inputs(160)) or (inputs(33));
    layer0_outputs(8605) <= not((inputs(226)) or (inputs(210)));
    layer0_outputs(8606) <= (inputs(230)) and not (inputs(239));
    layer0_outputs(8607) <= not((inputs(8)) xor (inputs(64)));
    layer0_outputs(8608) <= (inputs(95)) or (inputs(243));
    layer0_outputs(8609) <= not((inputs(9)) and (inputs(31)));
    layer0_outputs(8610) <= inputs(201);
    layer0_outputs(8611) <= not(inputs(26));
    layer0_outputs(8612) <= (inputs(40)) or (inputs(47));
    layer0_outputs(8613) <= (inputs(241)) xor (inputs(195));
    layer0_outputs(8614) <= (inputs(120)) xor (inputs(69));
    layer0_outputs(8615) <= not(inputs(88)) or (inputs(190));
    layer0_outputs(8616) <= inputs(49);
    layer0_outputs(8617) <= not(inputs(229));
    layer0_outputs(8618) <= (inputs(131)) xor (inputs(86));
    layer0_outputs(8619) <= not((inputs(227)) xor (inputs(161)));
    layer0_outputs(8620) <= not(inputs(117));
    layer0_outputs(8621) <= inputs(4);
    layer0_outputs(8622) <= (inputs(173)) xor (inputs(188));
    layer0_outputs(8623) <= (inputs(110)) or (inputs(38));
    layer0_outputs(8624) <= not(inputs(101)) or (inputs(58));
    layer0_outputs(8625) <= not((inputs(48)) or (inputs(50)));
    layer0_outputs(8626) <= inputs(61);
    layer0_outputs(8627) <= (inputs(4)) or (inputs(132));
    layer0_outputs(8628) <= not((inputs(48)) or (inputs(250)));
    layer0_outputs(8629) <= inputs(138);
    layer0_outputs(8630) <= not((inputs(228)) xor (inputs(81)));
    layer0_outputs(8631) <= (inputs(104)) and not (inputs(63));
    layer0_outputs(8632) <= not((inputs(138)) or (inputs(63)));
    layer0_outputs(8633) <= not(inputs(100));
    layer0_outputs(8634) <= not(inputs(38));
    layer0_outputs(8635) <= not(inputs(155));
    layer0_outputs(8636) <= not(inputs(231));
    layer0_outputs(8637) <= not((inputs(152)) and (inputs(220)));
    layer0_outputs(8638) <= (inputs(102)) xor (inputs(53));
    layer0_outputs(8639) <= inputs(110);
    layer0_outputs(8640) <= (inputs(127)) or (inputs(196));
    layer0_outputs(8641) <= not((inputs(122)) or (inputs(82)));
    layer0_outputs(8642) <= inputs(127);
    layer0_outputs(8643) <= not(inputs(11));
    layer0_outputs(8644) <= not(inputs(187));
    layer0_outputs(8645) <= (inputs(221)) and not (inputs(79));
    layer0_outputs(8646) <= not((inputs(2)) or (inputs(197)));
    layer0_outputs(8647) <= (inputs(190)) and not (inputs(144));
    layer0_outputs(8648) <= not(inputs(160));
    layer0_outputs(8649) <= not(inputs(108)) or (inputs(143));
    layer0_outputs(8650) <= (inputs(11)) xor (inputs(39));
    layer0_outputs(8651) <= not((inputs(69)) xor (inputs(134)));
    layer0_outputs(8652) <= (inputs(30)) or (inputs(133));
    layer0_outputs(8653) <= not((inputs(220)) and (inputs(189)));
    layer0_outputs(8654) <= not(inputs(195));
    layer0_outputs(8655) <= not(inputs(10));
    layer0_outputs(8656) <= (inputs(213)) and not (inputs(63));
    layer0_outputs(8657) <= (inputs(173)) or (inputs(202));
    layer0_outputs(8658) <= not((inputs(18)) or (inputs(126)));
    layer0_outputs(8659) <= not((inputs(158)) or (inputs(83)));
    layer0_outputs(8660) <= not((inputs(145)) or (inputs(214)));
    layer0_outputs(8661) <= inputs(73);
    layer0_outputs(8662) <= not(inputs(203));
    layer0_outputs(8663) <= not((inputs(149)) xor (inputs(63)));
    layer0_outputs(8664) <= (inputs(197)) or (inputs(145));
    layer0_outputs(8665) <= not(inputs(229)) or (inputs(224));
    layer0_outputs(8666) <= not((inputs(84)) or (inputs(83)));
    layer0_outputs(8667) <= not(inputs(18)) or (inputs(83));
    layer0_outputs(8668) <= not((inputs(2)) xor (inputs(149)));
    layer0_outputs(8669) <= inputs(132);
    layer0_outputs(8670) <= not((inputs(103)) xor (inputs(195)));
    layer0_outputs(8671) <= not((inputs(160)) xor (inputs(129)));
    layer0_outputs(8672) <= (inputs(154)) and (inputs(204));
    layer0_outputs(8673) <= inputs(127);
    layer0_outputs(8674) <= not((inputs(154)) or (inputs(123)));
    layer0_outputs(8675) <= (inputs(147)) or (inputs(204));
    layer0_outputs(8676) <= (inputs(253)) xor (inputs(250));
    layer0_outputs(8677) <= inputs(26);
    layer0_outputs(8678) <= (inputs(132)) xor (inputs(123));
    layer0_outputs(8679) <= (inputs(106)) or (inputs(138));
    layer0_outputs(8680) <= inputs(38);
    layer0_outputs(8681) <= not((inputs(117)) xor (inputs(142)));
    layer0_outputs(8682) <= (inputs(231)) and (inputs(77));
    layer0_outputs(8683) <= (inputs(252)) and not (inputs(159));
    layer0_outputs(8684) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(8685) <= not(inputs(78));
    layer0_outputs(8686) <= not(inputs(58)) or (inputs(193));
    layer0_outputs(8687) <= not((inputs(75)) and (inputs(41)));
    layer0_outputs(8688) <= not(inputs(234));
    layer0_outputs(8689) <= not((inputs(128)) or (inputs(193)));
    layer0_outputs(8690) <= not(inputs(22));
    layer0_outputs(8691) <= not((inputs(167)) xor (inputs(26)));
    layer0_outputs(8692) <= not(inputs(246)) or (inputs(34));
    layer0_outputs(8693) <= (inputs(49)) or (inputs(166));
    layer0_outputs(8694) <= (inputs(204)) or (inputs(216));
    layer0_outputs(8695) <= (inputs(103)) xor (inputs(17));
    layer0_outputs(8696) <= not((inputs(145)) and (inputs(184)));
    layer0_outputs(8697) <= not((inputs(208)) or (inputs(197)));
    layer0_outputs(8698) <= (inputs(130)) xor (inputs(206));
    layer0_outputs(8699) <= '0';
    layer0_outputs(8700) <= (inputs(253)) xor (inputs(137));
    layer0_outputs(8701) <= not((inputs(2)) or (inputs(160)));
    layer0_outputs(8702) <= '0';
    layer0_outputs(8703) <= not(inputs(21));
    layer0_outputs(8704) <= inputs(106);
    layer0_outputs(8705) <= not(inputs(67)) or (inputs(162));
    layer0_outputs(8706) <= not(inputs(111));
    layer0_outputs(8707) <= not((inputs(172)) or (inputs(208)));
    layer0_outputs(8708) <= not((inputs(29)) and (inputs(37)));
    layer0_outputs(8709) <= not((inputs(12)) or (inputs(198)));
    layer0_outputs(8710) <= not(inputs(105)) or (inputs(200));
    layer0_outputs(8711) <= not(inputs(54));
    layer0_outputs(8712) <= inputs(221);
    layer0_outputs(8713) <= (inputs(225)) or (inputs(6));
    layer0_outputs(8714) <= '0';
    layer0_outputs(8715) <= not(inputs(243)) or (inputs(13));
    layer0_outputs(8716) <= '0';
    layer0_outputs(8717) <= (inputs(104)) and not (inputs(239));
    layer0_outputs(8718) <= not((inputs(181)) xor (inputs(253)));
    layer0_outputs(8719) <= inputs(247);
    layer0_outputs(8720) <= (inputs(35)) or (inputs(179));
    layer0_outputs(8721) <= not((inputs(228)) or (inputs(253)));
    layer0_outputs(8722) <= (inputs(218)) and not (inputs(62));
    layer0_outputs(8723) <= not(inputs(139)) or (inputs(171));
    layer0_outputs(8724) <= inputs(60);
    layer0_outputs(8725) <= inputs(23);
    layer0_outputs(8726) <= inputs(83);
    layer0_outputs(8727) <= not(inputs(108));
    layer0_outputs(8728) <= not(inputs(84));
    layer0_outputs(8729) <= not(inputs(238));
    layer0_outputs(8730) <= not((inputs(104)) xor (inputs(169)));
    layer0_outputs(8731) <= (inputs(250)) or (inputs(166));
    layer0_outputs(8732) <= not(inputs(132)) or (inputs(50));
    layer0_outputs(8733) <= (inputs(220)) and not (inputs(119));
    layer0_outputs(8734) <= (inputs(3)) xor (inputs(9));
    layer0_outputs(8735) <= not(inputs(139));
    layer0_outputs(8736) <= not(inputs(106));
    layer0_outputs(8737) <= not(inputs(172)) or (inputs(106));
    layer0_outputs(8738) <= (inputs(134)) xor (inputs(196));
    layer0_outputs(8739) <= not((inputs(28)) and (inputs(120)));
    layer0_outputs(8740) <= not((inputs(47)) xor (inputs(68)));
    layer0_outputs(8741) <= '0';
    layer0_outputs(8742) <= (inputs(122)) and not (inputs(187));
    layer0_outputs(8743) <= not(inputs(201));
    layer0_outputs(8744) <= not(inputs(134)) or (inputs(158));
    layer0_outputs(8745) <= (inputs(44)) or (inputs(7));
    layer0_outputs(8746) <= not((inputs(155)) or (inputs(159)));
    layer0_outputs(8747) <= (inputs(241)) or (inputs(255));
    layer0_outputs(8748) <= inputs(6);
    layer0_outputs(8749) <= (inputs(185)) and (inputs(186));
    layer0_outputs(8750) <= not(inputs(107)) or (inputs(114));
    layer0_outputs(8751) <= (inputs(205)) xor (inputs(132));
    layer0_outputs(8752) <= (inputs(179)) xor (inputs(162));
    layer0_outputs(8753) <= not((inputs(149)) xor (inputs(119)));
    layer0_outputs(8754) <= (inputs(118)) xor (inputs(245));
    layer0_outputs(8755) <= (inputs(188)) xor (inputs(104));
    layer0_outputs(8756) <= (inputs(238)) and not (inputs(108));
    layer0_outputs(8757) <= not(inputs(57)) or (inputs(134));
    layer0_outputs(8758) <= not((inputs(20)) or (inputs(218)));
    layer0_outputs(8759) <= not(inputs(40)) or (inputs(33));
    layer0_outputs(8760) <= (inputs(140)) xor (inputs(9));
    layer0_outputs(8761) <= '0';
    layer0_outputs(8762) <= (inputs(158)) and not (inputs(125));
    layer0_outputs(8763) <= (inputs(69)) xor (inputs(83));
    layer0_outputs(8764) <= (inputs(239)) or (inputs(75));
    layer0_outputs(8765) <= not(inputs(59));
    layer0_outputs(8766) <= not((inputs(169)) or (inputs(146)));
    layer0_outputs(8767) <= (inputs(88)) xor (inputs(93));
    layer0_outputs(8768) <= (inputs(245)) xor (inputs(125));
    layer0_outputs(8769) <= not(inputs(79)) or (inputs(219));
    layer0_outputs(8770) <= inputs(2);
    layer0_outputs(8771) <= not((inputs(133)) xor (inputs(118)));
    layer0_outputs(8772) <= not(inputs(209));
    layer0_outputs(8773) <= not((inputs(95)) xor (inputs(73)));
    layer0_outputs(8774) <= (inputs(230)) and (inputs(91));
    layer0_outputs(8775) <= not((inputs(36)) xor (inputs(251)));
    layer0_outputs(8776) <= inputs(221);
    layer0_outputs(8777) <= '0';
    layer0_outputs(8778) <= inputs(103);
    layer0_outputs(8779) <= not(inputs(182)) or (inputs(143));
    layer0_outputs(8780) <= not(inputs(240));
    layer0_outputs(8781) <= not(inputs(232)) or (inputs(125));
    layer0_outputs(8782) <= not((inputs(250)) or (inputs(230)));
    layer0_outputs(8783) <= inputs(121);
    layer0_outputs(8784) <= (inputs(250)) xor (inputs(217));
    layer0_outputs(8785) <= inputs(227);
    layer0_outputs(8786) <= not(inputs(73));
    layer0_outputs(8787) <= not((inputs(178)) or (inputs(175)));
    layer0_outputs(8788) <= inputs(229);
    layer0_outputs(8789) <= (inputs(65)) xor (inputs(226));
    layer0_outputs(8790) <= (inputs(115)) xor (inputs(193));
    layer0_outputs(8791) <= not((inputs(89)) xor (inputs(41)));
    layer0_outputs(8792) <= (inputs(107)) xor (inputs(227));
    layer0_outputs(8793) <= not((inputs(7)) or (inputs(21)));
    layer0_outputs(8794) <= not(inputs(147));
    layer0_outputs(8795) <= (inputs(29)) xor (inputs(224));
    layer0_outputs(8796) <= (inputs(197)) and not (inputs(98));
    layer0_outputs(8797) <= not(inputs(45));
    layer0_outputs(8798) <= not(inputs(38));
    layer0_outputs(8799) <= (inputs(213)) or (inputs(219));
    layer0_outputs(8800) <= (inputs(151)) and not (inputs(232));
    layer0_outputs(8801) <= inputs(34);
    layer0_outputs(8802) <= not(inputs(198)) or (inputs(30));
    layer0_outputs(8803) <= (inputs(202)) and not (inputs(123));
    layer0_outputs(8804) <= (inputs(228)) and not (inputs(138));
    layer0_outputs(8805) <= not((inputs(133)) xor (inputs(83)));
    layer0_outputs(8806) <= (inputs(173)) or (inputs(177));
    layer0_outputs(8807) <= inputs(114);
    layer0_outputs(8808) <= (inputs(65)) or (inputs(135));
    layer0_outputs(8809) <= not(inputs(30));
    layer0_outputs(8810) <= not((inputs(131)) or (inputs(245)));
    layer0_outputs(8811) <= not((inputs(21)) or (inputs(126)));
    layer0_outputs(8812) <= not((inputs(115)) xor (inputs(17)));
    layer0_outputs(8813) <= not(inputs(164)) or (inputs(207));
    layer0_outputs(8814) <= (inputs(181)) and not (inputs(21));
    layer0_outputs(8815) <= inputs(49);
    layer0_outputs(8816) <= not(inputs(22));
    layer0_outputs(8817) <= (inputs(75)) xor (inputs(186));
    layer0_outputs(8818) <= not(inputs(231));
    layer0_outputs(8819) <= (inputs(3)) xor (inputs(153));
    layer0_outputs(8820) <= not(inputs(99)) or (inputs(206));
    layer0_outputs(8821) <= not(inputs(120));
    layer0_outputs(8822) <= (inputs(126)) and not (inputs(220));
    layer0_outputs(8823) <= not(inputs(210));
    layer0_outputs(8824) <= not((inputs(139)) or (inputs(203)));
    layer0_outputs(8825) <= inputs(148);
    layer0_outputs(8826) <= not(inputs(234)) or (inputs(112));
    layer0_outputs(8827) <= not(inputs(3));
    layer0_outputs(8828) <= (inputs(4)) and not (inputs(149));
    layer0_outputs(8829) <= not((inputs(70)) or (inputs(39)));
    layer0_outputs(8830) <= not((inputs(101)) or (inputs(90)));
    layer0_outputs(8831) <= (inputs(239)) xor (inputs(117));
    layer0_outputs(8832) <= not(inputs(186));
    layer0_outputs(8833) <= not(inputs(156)) or (inputs(28));
    layer0_outputs(8834) <= (inputs(51)) and not (inputs(161));
    layer0_outputs(8835) <= not(inputs(222)) or (inputs(96));
    layer0_outputs(8836) <= (inputs(185)) and (inputs(41));
    layer0_outputs(8837) <= (inputs(246)) and not (inputs(88));
    layer0_outputs(8838) <= not((inputs(28)) xor (inputs(153)));
    layer0_outputs(8839) <= (inputs(61)) and not (inputs(130));
    layer0_outputs(8840) <= (inputs(106)) and (inputs(122));
    layer0_outputs(8841) <= not(inputs(172)) or (inputs(251));
    layer0_outputs(8842) <= not(inputs(105)) or (inputs(132));
    layer0_outputs(8843) <= (inputs(217)) and not (inputs(50));
    layer0_outputs(8844) <= not(inputs(166));
    layer0_outputs(8845) <= inputs(156);
    layer0_outputs(8846) <= not(inputs(253));
    layer0_outputs(8847) <= inputs(76);
    layer0_outputs(8848) <= inputs(50);
    layer0_outputs(8849) <= (inputs(5)) or (inputs(186));
    layer0_outputs(8850) <= not(inputs(225));
    layer0_outputs(8851) <= (inputs(150)) or (inputs(158));
    layer0_outputs(8852) <= not((inputs(42)) xor (inputs(170)));
    layer0_outputs(8853) <= (inputs(192)) or (inputs(58));
    layer0_outputs(8854) <= not(inputs(3));
    layer0_outputs(8855) <= (inputs(210)) xor (inputs(203));
    layer0_outputs(8856) <= not((inputs(142)) or (inputs(204)));
    layer0_outputs(8857) <= (inputs(127)) and not (inputs(4));
    layer0_outputs(8858) <= not(inputs(179));
    layer0_outputs(8859) <= not(inputs(150));
    layer0_outputs(8860) <= (inputs(20)) xor (inputs(72));
    layer0_outputs(8861) <= not((inputs(23)) or (inputs(156)));
    layer0_outputs(8862) <= not(inputs(155));
    layer0_outputs(8863) <= not((inputs(132)) or (inputs(97)));
    layer0_outputs(8864) <= (inputs(225)) or (inputs(254));
    layer0_outputs(8865) <= (inputs(46)) xor (inputs(23));
    layer0_outputs(8866) <= (inputs(52)) or (inputs(7));
    layer0_outputs(8867) <= not(inputs(224)) or (inputs(252));
    layer0_outputs(8868) <= '0';
    layer0_outputs(8869) <= (inputs(242)) and not (inputs(120));
    layer0_outputs(8870) <= inputs(19);
    layer0_outputs(8871) <= (inputs(157)) xor (inputs(88));
    layer0_outputs(8872) <= (inputs(104)) and not (inputs(215));
    layer0_outputs(8873) <= not((inputs(245)) or (inputs(144)));
    layer0_outputs(8874) <= not(inputs(246)) or (inputs(142));
    layer0_outputs(8875) <= inputs(202);
    layer0_outputs(8876) <= not(inputs(183)) or (inputs(14));
    layer0_outputs(8877) <= (inputs(97)) or (inputs(238));
    layer0_outputs(8878) <= not((inputs(188)) or (inputs(64)));
    layer0_outputs(8879) <= (inputs(156)) xor (inputs(182));
    layer0_outputs(8880) <= not((inputs(181)) xor (inputs(33)));
    layer0_outputs(8881) <= (inputs(19)) and not (inputs(141));
    layer0_outputs(8882) <= not(inputs(102));
    layer0_outputs(8883) <= not((inputs(242)) xor (inputs(210)));
    layer0_outputs(8884) <= not(inputs(99));
    layer0_outputs(8885) <= (inputs(133)) and not (inputs(138));
    layer0_outputs(8886) <= (inputs(72)) and not (inputs(238));
    layer0_outputs(8887) <= not(inputs(233)) or (inputs(57));
    layer0_outputs(8888) <= inputs(189);
    layer0_outputs(8889) <= (inputs(37)) or (inputs(64));
    layer0_outputs(8890) <= inputs(165);
    layer0_outputs(8891) <= not(inputs(231));
    layer0_outputs(8892) <= not(inputs(212));
    layer0_outputs(8893) <= (inputs(236)) or (inputs(183));
    layer0_outputs(8894) <= not((inputs(66)) xor (inputs(212)));
    layer0_outputs(8895) <= not(inputs(113));
    layer0_outputs(8896) <= (inputs(113)) or (inputs(182));
    layer0_outputs(8897) <= inputs(25);
    layer0_outputs(8898) <= not((inputs(44)) or (inputs(129)));
    layer0_outputs(8899) <= (inputs(73)) xor (inputs(243));
    layer0_outputs(8900) <= (inputs(21)) and not (inputs(61));
    layer0_outputs(8901) <= not(inputs(85)) or (inputs(163));
    layer0_outputs(8902) <= not(inputs(5)) or (inputs(145));
    layer0_outputs(8903) <= not(inputs(131));
    layer0_outputs(8904) <= inputs(192);
    layer0_outputs(8905) <= not((inputs(96)) or (inputs(161)));
    layer0_outputs(8906) <= not(inputs(233)) or (inputs(224));
    layer0_outputs(8907) <= (inputs(135)) xor (inputs(103));
    layer0_outputs(8908) <= not((inputs(41)) or (inputs(2)));
    layer0_outputs(8909) <= not((inputs(186)) xor (inputs(219)));
    layer0_outputs(8910) <= inputs(199);
    layer0_outputs(8911) <= (inputs(50)) and not (inputs(139));
    layer0_outputs(8912) <= (inputs(72)) or (inputs(55));
    layer0_outputs(8913) <= inputs(154);
    layer0_outputs(8914) <= (inputs(81)) or (inputs(208));
    layer0_outputs(8915) <= not(inputs(194));
    layer0_outputs(8916) <= (inputs(4)) xor (inputs(136));
    layer0_outputs(8917) <= not(inputs(20)) or (inputs(199));
    layer0_outputs(8918) <= (inputs(62)) and not (inputs(175));
    layer0_outputs(8919) <= (inputs(247)) xor (inputs(144));
    layer0_outputs(8920) <= not((inputs(186)) xor (inputs(234)));
    layer0_outputs(8921) <= (inputs(249)) or (inputs(161));
    layer0_outputs(8922) <= (inputs(193)) xor (inputs(207));
    layer0_outputs(8923) <= (inputs(237)) or (inputs(238));
    layer0_outputs(8924) <= (inputs(166)) and not (inputs(159));
    layer0_outputs(8925) <= not((inputs(207)) or (inputs(49)));
    layer0_outputs(8926) <= (inputs(11)) and (inputs(77));
    layer0_outputs(8927) <= not((inputs(189)) or (inputs(242)));
    layer0_outputs(8928) <= (inputs(78)) xor (inputs(171));
    layer0_outputs(8929) <= not((inputs(202)) or (inputs(219)));
    layer0_outputs(8930) <= not(inputs(144));
    layer0_outputs(8931) <= not((inputs(217)) and (inputs(216)));
    layer0_outputs(8932) <= (inputs(137)) and not (inputs(250));
    layer0_outputs(8933) <= not(inputs(248));
    layer0_outputs(8934) <= not(inputs(38)) or (inputs(207));
    layer0_outputs(8935) <= (inputs(226)) or (inputs(132));
    layer0_outputs(8936) <= not((inputs(136)) xor (inputs(128)));
    layer0_outputs(8937) <= not(inputs(77));
    layer0_outputs(8938) <= (inputs(155)) and not (inputs(66));
    layer0_outputs(8939) <= (inputs(15)) and not (inputs(252));
    layer0_outputs(8940) <= not(inputs(142));
    layer0_outputs(8941) <= not(inputs(6)) or (inputs(84));
    layer0_outputs(8942) <= not(inputs(56));
    layer0_outputs(8943) <= (inputs(65)) or (inputs(121));
    layer0_outputs(8944) <= not((inputs(248)) or (inputs(192)));
    layer0_outputs(8945) <= (inputs(174)) or (inputs(246));
    layer0_outputs(8946) <= (inputs(134)) xor (inputs(22));
    layer0_outputs(8947) <= not(inputs(248)) or (inputs(27));
    layer0_outputs(8948) <= not(inputs(218)) or (inputs(127));
    layer0_outputs(8949) <= not(inputs(23));
    layer0_outputs(8950) <= (inputs(190)) and (inputs(110));
    layer0_outputs(8951) <= (inputs(199)) and not (inputs(29));
    layer0_outputs(8952) <= not((inputs(89)) or (inputs(18)));
    layer0_outputs(8953) <= inputs(47);
    layer0_outputs(8954) <= inputs(66);
    layer0_outputs(8955) <= not((inputs(40)) xor (inputs(8)));
    layer0_outputs(8956) <= not(inputs(35));
    layer0_outputs(8957) <= (inputs(192)) or (inputs(250));
    layer0_outputs(8958) <= (inputs(34)) and not (inputs(129));
    layer0_outputs(8959) <= not((inputs(91)) or (inputs(73)));
    layer0_outputs(8960) <= not(inputs(119));
    layer0_outputs(8961) <= '1';
    layer0_outputs(8962) <= not(inputs(229));
    layer0_outputs(8963) <= inputs(96);
    layer0_outputs(8964) <= (inputs(152)) or (inputs(190));
    layer0_outputs(8965) <= not(inputs(134));
    layer0_outputs(8966) <= inputs(110);
    layer0_outputs(8967) <= not((inputs(190)) or (inputs(203)));
    layer0_outputs(8968) <= not(inputs(91)) or (inputs(242));
    layer0_outputs(8969) <= not(inputs(168));
    layer0_outputs(8970) <= not(inputs(115)) or (inputs(176));
    layer0_outputs(8971) <= '0';
    layer0_outputs(8972) <= (inputs(23)) xor (inputs(34));
    layer0_outputs(8973) <= (inputs(84)) and not (inputs(181));
    layer0_outputs(8974) <= not((inputs(191)) and (inputs(70)));
    layer0_outputs(8975) <= (inputs(196)) and not (inputs(252));
    layer0_outputs(8976) <= not(inputs(39));
    layer0_outputs(8977) <= not(inputs(121)) or (inputs(161));
    layer0_outputs(8978) <= inputs(103);
    layer0_outputs(8979) <= not((inputs(25)) and (inputs(99)));
    layer0_outputs(8980) <= not(inputs(187)) or (inputs(48));
    layer0_outputs(8981) <= not(inputs(245));
    layer0_outputs(8982) <= inputs(113);
    layer0_outputs(8983) <= (inputs(123)) and not (inputs(161));
    layer0_outputs(8984) <= not(inputs(182));
    layer0_outputs(8985) <= not(inputs(152));
    layer0_outputs(8986) <= (inputs(59)) xor (inputs(48));
    layer0_outputs(8987) <= (inputs(129)) or (inputs(7));
    layer0_outputs(8988) <= not((inputs(192)) or (inputs(222)));
    layer0_outputs(8989) <= not(inputs(148));
    layer0_outputs(8990) <= '0';
    layer0_outputs(8991) <= inputs(198);
    layer0_outputs(8992) <= inputs(61);
    layer0_outputs(8993) <= (inputs(19)) and not (inputs(95));
    layer0_outputs(8994) <= not(inputs(251));
    layer0_outputs(8995) <= not((inputs(16)) or (inputs(55)));
    layer0_outputs(8996) <= not((inputs(170)) or (inputs(166)));
    layer0_outputs(8997) <= not(inputs(151)) or (inputs(142));
    layer0_outputs(8998) <= not((inputs(5)) xor (inputs(50)));
    layer0_outputs(8999) <= not(inputs(58));
    layer0_outputs(9000) <= (inputs(103)) or (inputs(223));
    layer0_outputs(9001) <= not((inputs(111)) xor (inputs(83)));
    layer0_outputs(9002) <= not(inputs(20)) or (inputs(163));
    layer0_outputs(9003) <= (inputs(47)) or (inputs(226));
    layer0_outputs(9004) <= not(inputs(196)) or (inputs(113));
    layer0_outputs(9005) <= inputs(14);
    layer0_outputs(9006) <= (inputs(248)) and not (inputs(62));
    layer0_outputs(9007) <= not((inputs(128)) or (inputs(126)));
    layer0_outputs(9008) <= not((inputs(101)) or (inputs(221)));
    layer0_outputs(9009) <= (inputs(60)) and not (inputs(205));
    layer0_outputs(9010) <= inputs(213);
    layer0_outputs(9011) <= not(inputs(22));
    layer0_outputs(9012) <= not(inputs(16));
    layer0_outputs(9013) <= (inputs(132)) xor (inputs(145));
    layer0_outputs(9014) <= not(inputs(131));
    layer0_outputs(9015) <= not((inputs(184)) or (inputs(73)));
    layer0_outputs(9016) <= (inputs(114)) and not (inputs(179));
    layer0_outputs(9017) <= not((inputs(168)) or (inputs(99)));
    layer0_outputs(9018) <= inputs(72);
    layer0_outputs(9019) <= not((inputs(105)) xor (inputs(83)));
    layer0_outputs(9020) <= not(inputs(231)) or (inputs(255));
    layer0_outputs(9021) <= not((inputs(73)) or (inputs(75)));
    layer0_outputs(9022) <= not(inputs(75));
    layer0_outputs(9023) <= not(inputs(144)) or (inputs(15));
    layer0_outputs(9024) <= not(inputs(205)) or (inputs(97));
    layer0_outputs(9025) <= not((inputs(127)) xor (inputs(133)));
    layer0_outputs(9026) <= not(inputs(23));
    layer0_outputs(9027) <= (inputs(179)) xor (inputs(245));
    layer0_outputs(9028) <= (inputs(112)) or (inputs(195));
    layer0_outputs(9029) <= not(inputs(122));
    layer0_outputs(9030) <= not(inputs(74));
    layer0_outputs(9031) <= inputs(94);
    layer0_outputs(9032) <= (inputs(74)) or (inputs(75));
    layer0_outputs(9033) <= not((inputs(210)) or (inputs(214)));
    layer0_outputs(9034) <= not(inputs(138));
    layer0_outputs(9035) <= inputs(120);
    layer0_outputs(9036) <= inputs(161);
    layer0_outputs(9037) <= (inputs(25)) and (inputs(122));
    layer0_outputs(9038) <= (inputs(64)) or (inputs(67));
    layer0_outputs(9039) <= inputs(82);
    layer0_outputs(9040) <= not((inputs(214)) and (inputs(215)));
    layer0_outputs(9041) <= (inputs(210)) and not (inputs(239));
    layer0_outputs(9042) <= not(inputs(205)) or (inputs(82));
    layer0_outputs(9043) <= not((inputs(138)) or (inputs(35)));
    layer0_outputs(9044) <= not(inputs(168)) or (inputs(205));
    layer0_outputs(9045) <= '1';
    layer0_outputs(9046) <= '0';
    layer0_outputs(9047) <= not((inputs(36)) or (inputs(197)));
    layer0_outputs(9048) <= inputs(37);
    layer0_outputs(9049) <= (inputs(143)) or (inputs(154));
    layer0_outputs(9050) <= not((inputs(144)) or (inputs(72)));
    layer0_outputs(9051) <= not((inputs(92)) xor (inputs(17)));
    layer0_outputs(9052) <= inputs(200);
    layer0_outputs(9053) <= inputs(41);
    layer0_outputs(9054) <= inputs(199);
    layer0_outputs(9055) <= '1';
    layer0_outputs(9056) <= (inputs(217)) xor (inputs(181));
    layer0_outputs(9057) <= not(inputs(28)) or (inputs(238));
    layer0_outputs(9058) <= (inputs(160)) or (inputs(140));
    layer0_outputs(9059) <= not((inputs(226)) xor (inputs(79)));
    layer0_outputs(9060) <= not(inputs(110));
    layer0_outputs(9061) <= (inputs(232)) and not (inputs(114));
    layer0_outputs(9062) <= inputs(187);
    layer0_outputs(9063) <= (inputs(22)) xor (inputs(75));
    layer0_outputs(9064) <= inputs(194);
    layer0_outputs(9065) <= not((inputs(149)) xor (inputs(119)));
    layer0_outputs(9066) <= not((inputs(122)) or (inputs(27)));
    layer0_outputs(9067) <= not(inputs(43));
    layer0_outputs(9068) <= not((inputs(44)) or (inputs(254)));
    layer0_outputs(9069) <= not((inputs(238)) xor (inputs(226)));
    layer0_outputs(9070) <= not(inputs(149)) or (inputs(230));
    layer0_outputs(9071) <= not((inputs(138)) or (inputs(34)));
    layer0_outputs(9072) <= (inputs(22)) xor (inputs(126));
    layer0_outputs(9073) <= not(inputs(113)) or (inputs(139));
    layer0_outputs(9074) <= inputs(70);
    layer0_outputs(9075) <= (inputs(5)) xor (inputs(19));
    layer0_outputs(9076) <= '0';
    layer0_outputs(9077) <= not(inputs(20)) or (inputs(83));
    layer0_outputs(9078) <= inputs(115);
    layer0_outputs(9079) <= not((inputs(65)) xor (inputs(121)));
    layer0_outputs(9080) <= (inputs(249)) and not (inputs(254));
    layer0_outputs(9081) <= not((inputs(235)) or (inputs(141)));
    layer0_outputs(9082) <= not((inputs(54)) or (inputs(20)));
    layer0_outputs(9083) <= not((inputs(229)) and (inputs(101)));
    layer0_outputs(9084) <= inputs(140);
    layer0_outputs(9085) <= (inputs(159)) or (inputs(19));
    layer0_outputs(9086) <= (inputs(180)) xor (inputs(252));
    layer0_outputs(9087) <= not((inputs(45)) or (inputs(201)));
    layer0_outputs(9088) <= not(inputs(26)) or (inputs(178));
    layer0_outputs(9089) <= (inputs(227)) and not (inputs(3));
    layer0_outputs(9090) <= not((inputs(139)) or (inputs(58)));
    layer0_outputs(9091) <= not((inputs(22)) or (inputs(103)));
    layer0_outputs(9092) <= (inputs(52)) xor (inputs(202));
    layer0_outputs(9093) <= not((inputs(33)) xor (inputs(249)));
    layer0_outputs(9094) <= not((inputs(146)) or (inputs(184)));
    layer0_outputs(9095) <= not(inputs(6)) or (inputs(80));
    layer0_outputs(9096) <= not((inputs(87)) or (inputs(204)));
    layer0_outputs(9097) <= not(inputs(230));
    layer0_outputs(9098) <= (inputs(203)) and not (inputs(96));
    layer0_outputs(9099) <= (inputs(95)) or (inputs(243));
    layer0_outputs(9100) <= not((inputs(192)) or (inputs(100)));
    layer0_outputs(9101) <= not((inputs(173)) or (inputs(204)));
    layer0_outputs(9102) <= (inputs(21)) and not (inputs(254));
    layer0_outputs(9103) <= (inputs(17)) xor (inputs(85));
    layer0_outputs(9104) <= (inputs(122)) and not (inputs(81));
    layer0_outputs(9105) <= inputs(58);
    layer0_outputs(9106) <= (inputs(89)) xor (inputs(171));
    layer0_outputs(9107) <= not(inputs(248));
    layer0_outputs(9108) <= not((inputs(14)) xor (inputs(44)));
    layer0_outputs(9109) <= (inputs(209)) and not (inputs(127));
    layer0_outputs(9110) <= not((inputs(130)) xor (inputs(214)));
    layer0_outputs(9111) <= not(inputs(133));
    layer0_outputs(9112) <= not(inputs(119)) or (inputs(129));
    layer0_outputs(9113) <= inputs(8);
    layer0_outputs(9114) <= not(inputs(248));
    layer0_outputs(9115) <= '1';
    layer0_outputs(9116) <= not((inputs(112)) or (inputs(212)));
    layer0_outputs(9117) <= (inputs(99)) or (inputs(125));
    layer0_outputs(9118) <= not(inputs(245));
    layer0_outputs(9119) <= not((inputs(96)) xor (inputs(71)));
    layer0_outputs(9120) <= not((inputs(53)) and (inputs(65)));
    layer0_outputs(9121) <= not((inputs(234)) or (inputs(231)));
    layer0_outputs(9122) <= inputs(217);
    layer0_outputs(9123) <= not((inputs(11)) or (inputs(219)));
    layer0_outputs(9124) <= not(inputs(217));
    layer0_outputs(9125) <= (inputs(168)) xor (inputs(60));
    layer0_outputs(9126) <= not((inputs(172)) and (inputs(184)));
    layer0_outputs(9127) <= not((inputs(132)) or (inputs(169)));
    layer0_outputs(9128) <= not(inputs(167)) or (inputs(213));
    layer0_outputs(9129) <= (inputs(245)) xor (inputs(221));
    layer0_outputs(9130) <= not((inputs(72)) xor (inputs(73)));
    layer0_outputs(9131) <= not((inputs(152)) xor (inputs(41)));
    layer0_outputs(9132) <= (inputs(202)) or (inputs(115));
    layer0_outputs(9133) <= not((inputs(254)) or (inputs(141)));
    layer0_outputs(9134) <= not(inputs(155)) or (inputs(109));
    layer0_outputs(9135) <= not((inputs(6)) or (inputs(252)));
    layer0_outputs(9136) <= not(inputs(139));
    layer0_outputs(9137) <= (inputs(175)) or (inputs(180));
    layer0_outputs(9138) <= (inputs(42)) xor (inputs(31));
    layer0_outputs(9139) <= (inputs(213)) and not (inputs(9));
    layer0_outputs(9140) <= not((inputs(149)) xor (inputs(166)));
    layer0_outputs(9141) <= not((inputs(239)) or (inputs(222)));
    layer0_outputs(9142) <= not((inputs(92)) or (inputs(144)));
    layer0_outputs(9143) <= not(inputs(28));
    layer0_outputs(9144) <= not((inputs(215)) or (inputs(15)));
    layer0_outputs(9145) <= not(inputs(21));
    layer0_outputs(9146) <= inputs(151);
    layer0_outputs(9147) <= (inputs(133)) or (inputs(141));
    layer0_outputs(9148) <= (inputs(35)) xor (inputs(173));
    layer0_outputs(9149) <= (inputs(119)) xor (inputs(19));
    layer0_outputs(9150) <= (inputs(123)) and (inputs(200));
    layer0_outputs(9151) <= inputs(15);
    layer0_outputs(9152) <= not(inputs(33));
    layer0_outputs(9153) <= not((inputs(202)) xor (inputs(33)));
    layer0_outputs(9154) <= not(inputs(238));
    layer0_outputs(9155) <= not(inputs(101));
    layer0_outputs(9156) <= (inputs(68)) or (inputs(246));
    layer0_outputs(9157) <= not(inputs(28)) or (inputs(146));
    layer0_outputs(9158) <= not(inputs(143)) or (inputs(6));
    layer0_outputs(9159) <= inputs(9);
    layer0_outputs(9160) <= not(inputs(254)) or (inputs(33));
    layer0_outputs(9161) <= not((inputs(54)) xor (inputs(22)));
    layer0_outputs(9162) <= (inputs(181)) or (inputs(199));
    layer0_outputs(9163) <= (inputs(255)) or (inputs(233));
    layer0_outputs(9164) <= not(inputs(200)) or (inputs(110));
    layer0_outputs(9165) <= not(inputs(216));
    layer0_outputs(9166) <= not(inputs(4));
    layer0_outputs(9167) <= not((inputs(68)) xor (inputs(85)));
    layer0_outputs(9168) <= not(inputs(129)) or (inputs(251));
    layer0_outputs(9169) <= inputs(219);
    layer0_outputs(9170) <= not(inputs(112)) or (inputs(238));
    layer0_outputs(9171) <= (inputs(104)) and (inputs(104));
    layer0_outputs(9172) <= not((inputs(84)) or (inputs(92)));
    layer0_outputs(9173) <= not((inputs(116)) xor (inputs(3)));
    layer0_outputs(9174) <= not(inputs(43));
    layer0_outputs(9175) <= not(inputs(115));
    layer0_outputs(9176) <= (inputs(203)) and (inputs(38));
    layer0_outputs(9177) <= not((inputs(8)) or (inputs(215)));
    layer0_outputs(9178) <= not(inputs(102));
    layer0_outputs(9179) <= not(inputs(166));
    layer0_outputs(9180) <= not((inputs(92)) or (inputs(75)));
    layer0_outputs(9181) <= (inputs(165)) or (inputs(6));
    layer0_outputs(9182) <= not(inputs(68));
    layer0_outputs(9183) <= not(inputs(34));
    layer0_outputs(9184) <= not(inputs(91));
    layer0_outputs(9185) <= (inputs(156)) xor (inputs(123));
    layer0_outputs(9186) <= (inputs(75)) xor (inputs(233));
    layer0_outputs(9187) <= (inputs(88)) or (inputs(226));
    layer0_outputs(9188) <= not(inputs(72));
    layer0_outputs(9189) <= '1';
    layer0_outputs(9190) <= not(inputs(188)) or (inputs(94));
    layer0_outputs(9191) <= not((inputs(238)) or (inputs(198)));
    layer0_outputs(9192) <= not(inputs(204));
    layer0_outputs(9193) <= not(inputs(7));
    layer0_outputs(9194) <= (inputs(20)) xor (inputs(216));
    layer0_outputs(9195) <= not(inputs(205));
    layer0_outputs(9196) <= not(inputs(132)) or (inputs(2));
    layer0_outputs(9197) <= (inputs(95)) and not (inputs(34));
    layer0_outputs(9198) <= not(inputs(216)) or (inputs(1));
    layer0_outputs(9199) <= '0';
    layer0_outputs(9200) <= inputs(211);
    layer0_outputs(9201) <= (inputs(91)) or (inputs(50));
    layer0_outputs(9202) <= (inputs(14)) or (inputs(107));
    layer0_outputs(9203) <= inputs(63);
    layer0_outputs(9204) <= not(inputs(246));
    layer0_outputs(9205) <= not((inputs(206)) xor (inputs(110)));
    layer0_outputs(9206) <= not(inputs(119)) or (inputs(96));
    layer0_outputs(9207) <= inputs(24);
    layer0_outputs(9208) <= inputs(170);
    layer0_outputs(9209) <= not((inputs(69)) and (inputs(157)));
    layer0_outputs(9210) <= inputs(129);
    layer0_outputs(9211) <= (inputs(137)) xor (inputs(57));
    layer0_outputs(9212) <= not(inputs(229)) or (inputs(63));
    layer0_outputs(9213) <= not((inputs(250)) xor (inputs(179)));
    layer0_outputs(9214) <= '1';
    layer0_outputs(9215) <= (inputs(161)) or (inputs(245));
    layer0_outputs(9216) <= not((inputs(2)) and (inputs(153)));
    layer0_outputs(9217) <= (inputs(117)) or (inputs(182));
    layer0_outputs(9218) <= (inputs(215)) and not (inputs(82));
    layer0_outputs(9219) <= inputs(9);
    layer0_outputs(9220) <= (inputs(131)) xor (inputs(53));
    layer0_outputs(9221) <= (inputs(138)) xor (inputs(199));
    layer0_outputs(9222) <= (inputs(119)) and not (inputs(62));
    layer0_outputs(9223) <= not(inputs(227)) or (inputs(224));
    layer0_outputs(9224) <= inputs(21);
    layer0_outputs(9225) <= (inputs(121)) or (inputs(110));
    layer0_outputs(9226) <= not((inputs(43)) or (inputs(155)));
    layer0_outputs(9227) <= inputs(16);
    layer0_outputs(9228) <= (inputs(136)) and not (inputs(130));
    layer0_outputs(9229) <= not(inputs(111)) or (inputs(3));
    layer0_outputs(9230) <= (inputs(153)) xor (inputs(242));
    layer0_outputs(9231) <= (inputs(207)) xor (inputs(26));
    layer0_outputs(9232) <= not((inputs(154)) xor (inputs(119)));
    layer0_outputs(9233) <= not(inputs(88)) or (inputs(34));
    layer0_outputs(9234) <= not(inputs(148));
    layer0_outputs(9235) <= not(inputs(123));
    layer0_outputs(9236) <= not(inputs(83));
    layer0_outputs(9237) <= '0';
    layer0_outputs(9238) <= not(inputs(36));
    layer0_outputs(9239) <= (inputs(205)) xor (inputs(171));
    layer0_outputs(9240) <= not(inputs(164)) or (inputs(99));
    layer0_outputs(9241) <= inputs(144);
    layer0_outputs(9242) <= (inputs(105)) or (inputs(241));
    layer0_outputs(9243) <= (inputs(105)) and not (inputs(177));
    layer0_outputs(9244) <= not((inputs(218)) or (inputs(252)));
    layer0_outputs(9245) <= (inputs(54)) xor (inputs(53));
    layer0_outputs(9246) <= inputs(135);
    layer0_outputs(9247) <= (inputs(228)) xor (inputs(162));
    layer0_outputs(9248) <= (inputs(56)) and not (inputs(22));
    layer0_outputs(9249) <= not(inputs(6));
    layer0_outputs(9250) <= not(inputs(57)) or (inputs(3));
    layer0_outputs(9251) <= not(inputs(184));
    layer0_outputs(9252) <= inputs(62);
    layer0_outputs(9253) <= inputs(180);
    layer0_outputs(9254) <= not(inputs(136));
    layer0_outputs(9255) <= not(inputs(165)) or (inputs(223));
    layer0_outputs(9256) <= (inputs(215)) xor (inputs(176));
    layer0_outputs(9257) <= '1';
    layer0_outputs(9258) <= (inputs(24)) or (inputs(24));
    layer0_outputs(9259) <= (inputs(4)) and not (inputs(80));
    layer0_outputs(9260) <= (inputs(252)) or (inputs(252));
    layer0_outputs(9261) <= (inputs(206)) xor (inputs(33));
    layer0_outputs(9262) <= (inputs(229)) and not (inputs(136));
    layer0_outputs(9263) <= (inputs(200)) and not (inputs(15));
    layer0_outputs(9264) <= (inputs(209)) and not (inputs(128));
    layer0_outputs(9265) <= not(inputs(166)) or (inputs(30));
    layer0_outputs(9266) <= (inputs(131)) or (inputs(80));
    layer0_outputs(9267) <= (inputs(4)) or (inputs(61));
    layer0_outputs(9268) <= not((inputs(171)) or (inputs(188)));
    layer0_outputs(9269) <= (inputs(164)) xor (inputs(211));
    layer0_outputs(9270) <= not(inputs(158));
    layer0_outputs(9271) <= not(inputs(178));
    layer0_outputs(9272) <= not((inputs(193)) or (inputs(25)));
    layer0_outputs(9273) <= not(inputs(113));
    layer0_outputs(9274) <= inputs(129);
    layer0_outputs(9275) <= not((inputs(165)) and (inputs(199)));
    layer0_outputs(9276) <= not(inputs(126));
    layer0_outputs(9277) <= not((inputs(251)) or (inputs(223)));
    layer0_outputs(9278) <= not(inputs(218));
    layer0_outputs(9279) <= (inputs(133)) and not (inputs(48));
    layer0_outputs(9280) <= (inputs(66)) xor (inputs(62));
    layer0_outputs(9281) <= inputs(212);
    layer0_outputs(9282) <= not(inputs(20)) or (inputs(188));
    layer0_outputs(9283) <= not((inputs(192)) or (inputs(43)));
    layer0_outputs(9284) <= inputs(247);
    layer0_outputs(9285) <= inputs(79);
    layer0_outputs(9286) <= not(inputs(67)) or (inputs(205));
    layer0_outputs(9287) <= not(inputs(102)) or (inputs(14));
    layer0_outputs(9288) <= inputs(69);
    layer0_outputs(9289) <= not(inputs(215));
    layer0_outputs(9290) <= not((inputs(26)) xor (inputs(74)));
    layer0_outputs(9291) <= (inputs(71)) and not (inputs(80));
    layer0_outputs(9292) <= inputs(145);
    layer0_outputs(9293) <= not(inputs(64));
    layer0_outputs(9294) <= (inputs(146)) xor (inputs(120));
    layer0_outputs(9295) <= '1';
    layer0_outputs(9296) <= not(inputs(114));
    layer0_outputs(9297) <= not((inputs(40)) or (inputs(142)));
    layer0_outputs(9298) <= not(inputs(149)) or (inputs(76));
    layer0_outputs(9299) <= not(inputs(223));
    layer0_outputs(9300) <= (inputs(205)) xor (inputs(16));
    layer0_outputs(9301) <= inputs(70);
    layer0_outputs(9302) <= (inputs(7)) or (inputs(84));
    layer0_outputs(9303) <= (inputs(24)) and not (inputs(197));
    layer0_outputs(9304) <= inputs(163);
    layer0_outputs(9305) <= '0';
    layer0_outputs(9306) <= (inputs(154)) xor (inputs(153));
    layer0_outputs(9307) <= inputs(102);
    layer0_outputs(9308) <= (inputs(89)) and not (inputs(97));
    layer0_outputs(9309) <= (inputs(212)) or (inputs(32));
    layer0_outputs(9310) <= not(inputs(29));
    layer0_outputs(9311) <= (inputs(219)) xor (inputs(231));
    layer0_outputs(9312) <= inputs(117);
    layer0_outputs(9313) <= (inputs(117)) xor (inputs(181));
    layer0_outputs(9314) <= (inputs(103)) and (inputs(92));
    layer0_outputs(9315) <= not(inputs(211));
    layer0_outputs(9316) <= not((inputs(240)) xor (inputs(5)));
    layer0_outputs(9317) <= not((inputs(164)) xor (inputs(134)));
    layer0_outputs(9318) <= not((inputs(178)) or (inputs(22)));
    layer0_outputs(9319) <= not((inputs(69)) xor (inputs(97)));
    layer0_outputs(9320) <= (inputs(98)) and (inputs(22));
    layer0_outputs(9321) <= inputs(251);
    layer0_outputs(9322) <= inputs(65);
    layer0_outputs(9323) <= (inputs(186)) and (inputs(109));
    layer0_outputs(9324) <= not((inputs(204)) or (inputs(196)));
    layer0_outputs(9325) <= inputs(231);
    layer0_outputs(9326) <= not((inputs(179)) xor (inputs(86)));
    layer0_outputs(9327) <= '1';
    layer0_outputs(9328) <= not(inputs(214));
    layer0_outputs(9329) <= (inputs(255)) or (inputs(188));
    layer0_outputs(9330) <= not((inputs(198)) xor (inputs(183)));
    layer0_outputs(9331) <= not((inputs(247)) xor (inputs(77)));
    layer0_outputs(9332) <= not(inputs(18)) or (inputs(114));
    layer0_outputs(9333) <= inputs(25);
    layer0_outputs(9334) <= (inputs(80)) and not (inputs(39));
    layer0_outputs(9335) <= inputs(94);
    layer0_outputs(9336) <= (inputs(73)) or (inputs(129));
    layer0_outputs(9337) <= (inputs(166)) and (inputs(148));
    layer0_outputs(9338) <= not((inputs(83)) or (inputs(47)));
    layer0_outputs(9339) <= not((inputs(173)) xor (inputs(223)));
    layer0_outputs(9340) <= (inputs(248)) and not (inputs(82));
    layer0_outputs(9341) <= inputs(164);
    layer0_outputs(9342) <= not(inputs(234));
    layer0_outputs(9343) <= not((inputs(203)) or (inputs(86)));
    layer0_outputs(9344) <= not(inputs(154)) or (inputs(193));
    layer0_outputs(9345) <= not(inputs(203));
    layer0_outputs(9346) <= (inputs(127)) and (inputs(13));
    layer0_outputs(9347) <= inputs(101);
    layer0_outputs(9348) <= not((inputs(91)) or (inputs(216)));
    layer0_outputs(9349) <= not(inputs(46));
    layer0_outputs(9350) <= inputs(88);
    layer0_outputs(9351) <= inputs(68);
    layer0_outputs(9352) <= (inputs(198)) xor (inputs(38));
    layer0_outputs(9353) <= (inputs(40)) and (inputs(54));
    layer0_outputs(9354) <= not((inputs(177)) xor (inputs(149)));
    layer0_outputs(9355) <= inputs(166);
    layer0_outputs(9356) <= inputs(246);
    layer0_outputs(9357) <= inputs(87);
    layer0_outputs(9358) <= not(inputs(58));
    layer0_outputs(9359) <= not(inputs(126));
    layer0_outputs(9360) <= not((inputs(242)) or (inputs(182)));
    layer0_outputs(9361) <= inputs(212);
    layer0_outputs(9362) <= not((inputs(103)) or (inputs(111)));
    layer0_outputs(9363) <= not(inputs(11)) or (inputs(191));
    layer0_outputs(9364) <= (inputs(212)) and (inputs(149));
    layer0_outputs(9365) <= (inputs(131)) or (inputs(235));
    layer0_outputs(9366) <= (inputs(57)) and not (inputs(79));
    layer0_outputs(9367) <= not((inputs(17)) or (inputs(159)));
    layer0_outputs(9368) <= not(inputs(131)) or (inputs(214));
    layer0_outputs(9369) <= not((inputs(54)) xor (inputs(89)));
    layer0_outputs(9370) <= not((inputs(115)) xor (inputs(252)));
    layer0_outputs(9371) <= not(inputs(12)) or (inputs(154));
    layer0_outputs(9372) <= not((inputs(7)) or (inputs(229)));
    layer0_outputs(9373) <= inputs(170);
    layer0_outputs(9374) <= inputs(231);
    layer0_outputs(9375) <= (inputs(222)) xor (inputs(209));
    layer0_outputs(9376) <= not(inputs(170)) or (inputs(63));
    layer0_outputs(9377) <= not(inputs(103)) or (inputs(174));
    layer0_outputs(9378) <= not(inputs(51));
    layer0_outputs(9379) <= (inputs(210)) or (inputs(195));
    layer0_outputs(9380) <= not(inputs(148));
    layer0_outputs(9381) <= (inputs(23)) or (inputs(59));
    layer0_outputs(9382) <= (inputs(141)) and not (inputs(66));
    layer0_outputs(9383) <= not(inputs(114));
    layer0_outputs(9384) <= (inputs(157)) xor (inputs(140));
    layer0_outputs(9385) <= not((inputs(139)) xor (inputs(172)));
    layer0_outputs(9386) <= not(inputs(13)) or (inputs(208));
    layer0_outputs(9387) <= (inputs(201)) and (inputs(155));
    layer0_outputs(9388) <= not((inputs(119)) and (inputs(40)));
    layer0_outputs(9389) <= not((inputs(230)) xor (inputs(251)));
    layer0_outputs(9390) <= not((inputs(63)) xor (inputs(133)));
    layer0_outputs(9391) <= not((inputs(61)) and (inputs(107)));
    layer0_outputs(9392) <= (inputs(249)) xor (inputs(187));
    layer0_outputs(9393) <= inputs(172);
    layer0_outputs(9394) <= (inputs(106)) and not (inputs(28));
    layer0_outputs(9395) <= (inputs(43)) and (inputs(8));
    layer0_outputs(9396) <= inputs(65);
    layer0_outputs(9397) <= (inputs(57)) and not (inputs(97));
    layer0_outputs(9398) <= not((inputs(131)) xor (inputs(195)));
    layer0_outputs(9399) <= not(inputs(64));
    layer0_outputs(9400) <= not((inputs(90)) xor (inputs(170)));
    layer0_outputs(9401) <= inputs(76);
    layer0_outputs(9402) <= not(inputs(53));
    layer0_outputs(9403) <= inputs(216);
    layer0_outputs(9404) <= not(inputs(207)) or (inputs(236));
    layer0_outputs(9405) <= not(inputs(25));
    layer0_outputs(9406) <= (inputs(127)) and not (inputs(238));
    layer0_outputs(9407) <= (inputs(48)) xor (inputs(110));
    layer0_outputs(9408) <= (inputs(146)) xor (inputs(117));
    layer0_outputs(9409) <= not(inputs(254));
    layer0_outputs(9410) <= inputs(102);
    layer0_outputs(9411) <= inputs(142);
    layer0_outputs(9412) <= (inputs(155)) or (inputs(18));
    layer0_outputs(9413) <= (inputs(135)) and (inputs(115));
    layer0_outputs(9414) <= not(inputs(39)) or (inputs(77));
    layer0_outputs(9415) <= not((inputs(215)) or (inputs(118)));
    layer0_outputs(9416) <= not(inputs(72));
    layer0_outputs(9417) <= not(inputs(192)) or (inputs(202));
    layer0_outputs(9418) <= (inputs(3)) and not (inputs(160));
    layer0_outputs(9419) <= not((inputs(186)) or (inputs(17)));
    layer0_outputs(9420) <= (inputs(138)) or (inputs(113));
    layer0_outputs(9421) <= not((inputs(53)) xor (inputs(14)));
    layer0_outputs(9422) <= inputs(137);
    layer0_outputs(9423) <= not(inputs(55));
    layer0_outputs(9424) <= not((inputs(41)) or (inputs(189)));
    layer0_outputs(9425) <= (inputs(39)) or (inputs(53));
    layer0_outputs(9426) <= (inputs(157)) or (inputs(173));
    layer0_outputs(9427) <= (inputs(45)) xor (inputs(92));
    layer0_outputs(9428) <= not(inputs(136)) or (inputs(248));
    layer0_outputs(9429) <= not((inputs(55)) or (inputs(79)));
    layer0_outputs(9430) <= not(inputs(8)) or (inputs(41));
    layer0_outputs(9431) <= not(inputs(177));
    layer0_outputs(9432) <= (inputs(157)) or (inputs(195));
    layer0_outputs(9433) <= (inputs(232)) or (inputs(206));
    layer0_outputs(9434) <= inputs(117);
    layer0_outputs(9435) <= not(inputs(221));
    layer0_outputs(9436) <= not(inputs(48)) or (inputs(10));
    layer0_outputs(9437) <= not(inputs(22));
    layer0_outputs(9438) <= not((inputs(135)) or (inputs(3)));
    layer0_outputs(9439) <= (inputs(36)) and not (inputs(79));
    layer0_outputs(9440) <= not(inputs(84));
    layer0_outputs(9441) <= not(inputs(66));
    layer0_outputs(9442) <= inputs(88);
    layer0_outputs(9443) <= (inputs(51)) and not (inputs(191));
    layer0_outputs(9444) <= inputs(228);
    layer0_outputs(9445) <= (inputs(106)) or (inputs(200));
    layer0_outputs(9446) <= inputs(182);
    layer0_outputs(9447) <= inputs(18);
    layer0_outputs(9448) <= inputs(249);
    layer0_outputs(9449) <= not((inputs(168)) and (inputs(143)));
    layer0_outputs(9450) <= not(inputs(143)) or (inputs(135));
    layer0_outputs(9451) <= (inputs(175)) xor (inputs(90));
    layer0_outputs(9452) <= inputs(115);
    layer0_outputs(9453) <= not(inputs(49));
    layer0_outputs(9454) <= not(inputs(184));
    layer0_outputs(9455) <= inputs(94);
    layer0_outputs(9456) <= not(inputs(93));
    layer0_outputs(9457) <= not(inputs(250)) or (inputs(140));
    layer0_outputs(9458) <= not((inputs(143)) or (inputs(126)));
    layer0_outputs(9459) <= not((inputs(97)) xor (inputs(88)));
    layer0_outputs(9460) <= inputs(92);
    layer0_outputs(9461) <= not(inputs(245));
    layer0_outputs(9462) <= (inputs(44)) xor (inputs(208));
    layer0_outputs(9463) <= (inputs(75)) and not (inputs(223));
    layer0_outputs(9464) <= not(inputs(74)) or (inputs(48));
    layer0_outputs(9465) <= inputs(36);
    layer0_outputs(9466) <= inputs(137);
    layer0_outputs(9467) <= not((inputs(27)) or (inputs(172)));
    layer0_outputs(9468) <= inputs(92);
    layer0_outputs(9469) <= not(inputs(101));
    layer0_outputs(9470) <= (inputs(50)) and not (inputs(173));
    layer0_outputs(9471) <= (inputs(67)) xor (inputs(80));
    layer0_outputs(9472) <= (inputs(244)) and not (inputs(15));
    layer0_outputs(9473) <= not(inputs(12)) or (inputs(91));
    layer0_outputs(9474) <= (inputs(205)) or (inputs(241));
    layer0_outputs(9475) <= not(inputs(221));
    layer0_outputs(9476) <= not(inputs(9));
    layer0_outputs(9477) <= not(inputs(166));
    layer0_outputs(9478) <= (inputs(101)) xor (inputs(170));
    layer0_outputs(9479) <= (inputs(17)) xor (inputs(21));
    layer0_outputs(9480) <= (inputs(53)) xor (inputs(62));
    layer0_outputs(9481) <= not((inputs(164)) xor (inputs(181)));
    layer0_outputs(9482) <= not((inputs(135)) or (inputs(250)));
    layer0_outputs(9483) <= not(inputs(85));
    layer0_outputs(9484) <= not((inputs(31)) or (inputs(242)));
    layer0_outputs(9485) <= not((inputs(188)) xor (inputs(162)));
    layer0_outputs(9486) <= not(inputs(152));
    layer0_outputs(9487) <= not(inputs(222));
    layer0_outputs(9488) <= not(inputs(102)) or (inputs(214));
    layer0_outputs(9489) <= not((inputs(34)) xor (inputs(189)));
    layer0_outputs(9490) <= inputs(51);
    layer0_outputs(9491) <= not((inputs(192)) and (inputs(224)));
    layer0_outputs(9492) <= (inputs(195)) and not (inputs(184));
    layer0_outputs(9493) <= not((inputs(229)) xor (inputs(248)));
    layer0_outputs(9494) <= (inputs(196)) or (inputs(104));
    layer0_outputs(9495) <= not(inputs(145));
    layer0_outputs(9496) <= not((inputs(226)) xor (inputs(103)));
    layer0_outputs(9497) <= not((inputs(4)) xor (inputs(35)));
    layer0_outputs(9498) <= not(inputs(23));
    layer0_outputs(9499) <= (inputs(189)) xor (inputs(129));
    layer0_outputs(9500) <= (inputs(231)) or (inputs(253));
    layer0_outputs(9501) <= not(inputs(133)) or (inputs(3));
    layer0_outputs(9502) <= not((inputs(241)) or (inputs(109)));
    layer0_outputs(9503) <= (inputs(39)) xor (inputs(212));
    layer0_outputs(9504) <= not(inputs(98)) or (inputs(147));
    layer0_outputs(9505) <= not(inputs(37)) or (inputs(164));
    layer0_outputs(9506) <= inputs(77);
    layer0_outputs(9507) <= inputs(245);
    layer0_outputs(9508) <= not(inputs(66));
    layer0_outputs(9509) <= not((inputs(134)) and (inputs(206)));
    layer0_outputs(9510) <= not(inputs(238)) or (inputs(110));
    layer0_outputs(9511) <= not((inputs(175)) xor (inputs(164)));
    layer0_outputs(9512) <= not(inputs(52));
    layer0_outputs(9513) <= inputs(248);
    layer0_outputs(9514) <= not(inputs(224)) or (inputs(196));
    layer0_outputs(9515) <= (inputs(21)) and (inputs(148));
    layer0_outputs(9516) <= not(inputs(167));
    layer0_outputs(9517) <= not(inputs(233));
    layer0_outputs(9518) <= (inputs(199)) and not (inputs(94));
    layer0_outputs(9519) <= inputs(222);
    layer0_outputs(9520) <= not((inputs(95)) or (inputs(219)));
    layer0_outputs(9521) <= not(inputs(154)) or (inputs(103));
    layer0_outputs(9522) <= not(inputs(65));
    layer0_outputs(9523) <= (inputs(137)) and not (inputs(178));
    layer0_outputs(9524) <= not(inputs(67)) or (inputs(181));
    layer0_outputs(9525) <= (inputs(104)) or (inputs(117));
    layer0_outputs(9526) <= (inputs(108)) or (inputs(59));
    layer0_outputs(9527) <= (inputs(19)) xor (inputs(189));
    layer0_outputs(9528) <= not((inputs(204)) or (inputs(155)));
    layer0_outputs(9529) <= not((inputs(225)) xor (inputs(91)));
    layer0_outputs(9530) <= inputs(60);
    layer0_outputs(9531) <= not(inputs(22));
    layer0_outputs(9532) <= not(inputs(36)) or (inputs(152));
    layer0_outputs(9533) <= not(inputs(13));
    layer0_outputs(9534) <= not(inputs(95));
    layer0_outputs(9535) <= '0';
    layer0_outputs(9536) <= inputs(165);
    layer0_outputs(9537) <= not((inputs(212)) or (inputs(147)));
    layer0_outputs(9538) <= (inputs(208)) and (inputs(168));
    layer0_outputs(9539) <= not(inputs(166));
    layer0_outputs(9540) <= inputs(119);
    layer0_outputs(9541) <= not(inputs(28));
    layer0_outputs(9542) <= not((inputs(54)) xor (inputs(171)));
    layer0_outputs(9543) <= (inputs(174)) xor (inputs(131));
    layer0_outputs(9544) <= inputs(228);
    layer0_outputs(9545) <= not((inputs(144)) xor (inputs(92)));
    layer0_outputs(9546) <= inputs(246);
    layer0_outputs(9547) <= (inputs(44)) and not (inputs(206));
    layer0_outputs(9548) <= inputs(177);
    layer0_outputs(9549) <= inputs(148);
    layer0_outputs(9550) <= (inputs(41)) or (inputs(105));
    layer0_outputs(9551) <= not(inputs(181));
    layer0_outputs(9552) <= (inputs(216)) and not (inputs(109));
    layer0_outputs(9553) <= not((inputs(176)) xor (inputs(228)));
    layer0_outputs(9554) <= (inputs(56)) and not (inputs(254));
    layer0_outputs(9555) <= not((inputs(1)) or (inputs(205)));
    layer0_outputs(9556) <= not((inputs(157)) or (inputs(128)));
    layer0_outputs(9557) <= '1';
    layer0_outputs(9558) <= (inputs(140)) and not (inputs(112));
    layer0_outputs(9559) <= inputs(166);
    layer0_outputs(9560) <= not((inputs(80)) and (inputs(243)));
    layer0_outputs(9561) <= inputs(10);
    layer0_outputs(9562) <= not((inputs(197)) xor (inputs(164)));
    layer0_outputs(9563) <= (inputs(117)) and not (inputs(159));
    layer0_outputs(9564) <= not(inputs(236)) or (inputs(144));
    layer0_outputs(9565) <= not(inputs(54));
    layer0_outputs(9566) <= not((inputs(122)) and (inputs(85)));
    layer0_outputs(9567) <= not(inputs(244)) or (inputs(253));
    layer0_outputs(9568) <= not(inputs(107));
    layer0_outputs(9569) <= not((inputs(148)) xor (inputs(36)));
    layer0_outputs(9570) <= not(inputs(12));
    layer0_outputs(9571) <= not((inputs(128)) or (inputs(154)));
    layer0_outputs(9572) <= (inputs(27)) or (inputs(239));
    layer0_outputs(9573) <= not((inputs(183)) or (inputs(101)));
    layer0_outputs(9574) <= not((inputs(156)) xor (inputs(51)));
    layer0_outputs(9575) <= (inputs(210)) and not (inputs(87));
    layer0_outputs(9576) <= not(inputs(189)) or (inputs(91));
    layer0_outputs(9577) <= (inputs(42)) and not (inputs(45));
    layer0_outputs(9578) <= not(inputs(226));
    layer0_outputs(9579) <= not(inputs(133));
    layer0_outputs(9580) <= inputs(247);
    layer0_outputs(9581) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(9582) <= (inputs(44)) xor (inputs(141));
    layer0_outputs(9583) <= not(inputs(231));
    layer0_outputs(9584) <= (inputs(11)) or (inputs(75));
    layer0_outputs(9585) <= (inputs(177)) xor (inputs(228));
    layer0_outputs(9586) <= (inputs(8)) and not (inputs(98));
    layer0_outputs(9587) <= not((inputs(1)) or (inputs(195)));
    layer0_outputs(9588) <= inputs(39);
    layer0_outputs(9589) <= not(inputs(23)) or (inputs(35));
    layer0_outputs(9590) <= not(inputs(23));
    layer0_outputs(9591) <= inputs(70);
    layer0_outputs(9592) <= not((inputs(244)) or (inputs(218)));
    layer0_outputs(9593) <= not((inputs(65)) xor (inputs(118)));
    layer0_outputs(9594) <= not((inputs(131)) or (inputs(190)));
    layer0_outputs(9595) <= (inputs(68)) and not (inputs(225));
    layer0_outputs(9596) <= inputs(234);
    layer0_outputs(9597) <= not(inputs(27)) or (inputs(186));
    layer0_outputs(9598) <= not((inputs(66)) or (inputs(120)));
    layer0_outputs(9599) <= not((inputs(237)) or (inputs(13)));
    layer0_outputs(9600) <= (inputs(232)) and not (inputs(63));
    layer0_outputs(9601) <= not((inputs(216)) and (inputs(89)));
    layer0_outputs(9602) <= inputs(17);
    layer0_outputs(9603) <= (inputs(201)) xor (inputs(193));
    layer0_outputs(9604) <= inputs(57);
    layer0_outputs(9605) <= not((inputs(112)) or (inputs(120)));
    layer0_outputs(9606) <= (inputs(102)) xor (inputs(141));
    layer0_outputs(9607) <= not(inputs(24));
    layer0_outputs(9608) <= (inputs(35)) and not (inputs(232));
    layer0_outputs(9609) <= (inputs(175)) xor (inputs(107));
    layer0_outputs(9610) <= (inputs(104)) and not (inputs(97));
    layer0_outputs(9611) <= not(inputs(25));
    layer0_outputs(9612) <= inputs(145);
    layer0_outputs(9613) <= (inputs(247)) xor (inputs(244));
    layer0_outputs(9614) <= (inputs(24)) and (inputs(25));
    layer0_outputs(9615) <= not((inputs(132)) xor (inputs(98)));
    layer0_outputs(9616) <= not((inputs(130)) or (inputs(81)));
    layer0_outputs(9617) <= inputs(130);
    layer0_outputs(9618) <= (inputs(115)) xor (inputs(32));
    layer0_outputs(9619) <= not((inputs(128)) or (inputs(6)));
    layer0_outputs(9620) <= inputs(252);
    layer0_outputs(9621) <= (inputs(55)) and not (inputs(146));
    layer0_outputs(9622) <= not((inputs(170)) and (inputs(158)));
    layer0_outputs(9623) <= not((inputs(213)) and (inputs(230)));
    layer0_outputs(9624) <= not((inputs(157)) and (inputs(94)));
    layer0_outputs(9625) <= not((inputs(41)) xor (inputs(159)));
    layer0_outputs(9626) <= not((inputs(80)) or (inputs(236)));
    layer0_outputs(9627) <= not((inputs(27)) xor (inputs(39)));
    layer0_outputs(9628) <= (inputs(166)) and not (inputs(46));
    layer0_outputs(9629) <= not((inputs(12)) or (inputs(41)));
    layer0_outputs(9630) <= not(inputs(46));
    layer0_outputs(9631) <= inputs(182);
    layer0_outputs(9632) <= (inputs(191)) xor (inputs(99));
    layer0_outputs(9633) <= (inputs(49)) or (inputs(61));
    layer0_outputs(9634) <= not((inputs(213)) or (inputs(17)));
    layer0_outputs(9635) <= not(inputs(237)) or (inputs(142));
    layer0_outputs(9636) <= not(inputs(195)) or (inputs(79));
    layer0_outputs(9637) <= (inputs(229)) xor (inputs(165));
    layer0_outputs(9638) <= not(inputs(134)) or (inputs(159));
    layer0_outputs(9639) <= not((inputs(183)) xor (inputs(136)));
    layer0_outputs(9640) <= (inputs(216)) and not (inputs(77));
    layer0_outputs(9641) <= not((inputs(214)) xor (inputs(37)));
    layer0_outputs(9642) <= not((inputs(171)) xor (inputs(247)));
    layer0_outputs(9643) <= (inputs(253)) or (inputs(169));
    layer0_outputs(9644) <= inputs(85);
    layer0_outputs(9645) <= not((inputs(158)) or (inputs(106)));
    layer0_outputs(9646) <= (inputs(156)) xor (inputs(130));
    layer0_outputs(9647) <= (inputs(77)) or (inputs(239));
    layer0_outputs(9648) <= (inputs(206)) xor (inputs(63));
    layer0_outputs(9649) <= (inputs(140)) and not (inputs(63));
    layer0_outputs(9650) <= (inputs(46)) xor (inputs(58));
    layer0_outputs(9651) <= (inputs(25)) xor (inputs(64));
    layer0_outputs(9652) <= inputs(70);
    layer0_outputs(9653) <= not(inputs(92));
    layer0_outputs(9654) <= (inputs(255)) or (inputs(234));
    layer0_outputs(9655) <= not(inputs(210)) or (inputs(64));
    layer0_outputs(9656) <= (inputs(4)) xor (inputs(26));
    layer0_outputs(9657) <= not((inputs(89)) and (inputs(169)));
    layer0_outputs(9658) <= not(inputs(160));
    layer0_outputs(9659) <= inputs(197);
    layer0_outputs(9660) <= inputs(162);
    layer0_outputs(9661) <= (inputs(112)) or (inputs(246));
    layer0_outputs(9662) <= inputs(181);
    layer0_outputs(9663) <= inputs(226);
    layer0_outputs(9664) <= (inputs(15)) xor (inputs(190));
    layer0_outputs(9665) <= not((inputs(158)) or (inputs(185)));
    layer0_outputs(9666) <= inputs(221);
    layer0_outputs(9667) <= not(inputs(99));
    layer0_outputs(9668) <= inputs(108);
    layer0_outputs(9669) <= not(inputs(169)) or (inputs(197));
    layer0_outputs(9670) <= (inputs(189)) or (inputs(174));
    layer0_outputs(9671) <= not(inputs(118)) or (inputs(228));
    layer0_outputs(9672) <= not((inputs(71)) xor (inputs(133)));
    layer0_outputs(9673) <= inputs(19);
    layer0_outputs(9674) <= not((inputs(123)) xor (inputs(117)));
    layer0_outputs(9675) <= (inputs(180)) and not (inputs(78));
    layer0_outputs(9676) <= (inputs(143)) or (inputs(41));
    layer0_outputs(9677) <= not((inputs(36)) and (inputs(102)));
    layer0_outputs(9678) <= not(inputs(145));
    layer0_outputs(9679) <= not((inputs(46)) xor (inputs(88)));
    layer0_outputs(9680) <= (inputs(157)) or (inputs(69));
    layer0_outputs(9681) <= (inputs(236)) xor (inputs(157));
    layer0_outputs(9682) <= (inputs(181)) or (inputs(92));
    layer0_outputs(9683) <= not(inputs(167));
    layer0_outputs(9684) <= not((inputs(234)) or (inputs(48)));
    layer0_outputs(9685) <= (inputs(186)) and not (inputs(62));
    layer0_outputs(9686) <= not(inputs(120)) or (inputs(56));
    layer0_outputs(9687) <= (inputs(209)) or (inputs(194));
    layer0_outputs(9688) <= inputs(127);
    layer0_outputs(9689) <= (inputs(151)) or (inputs(64));
    layer0_outputs(9690) <= (inputs(109)) or (inputs(42));
    layer0_outputs(9691) <= inputs(128);
    layer0_outputs(9692) <= not(inputs(59)) or (inputs(174));
    layer0_outputs(9693) <= inputs(171);
    layer0_outputs(9694) <= (inputs(199)) or (inputs(169));
    layer0_outputs(9695) <= (inputs(185)) and (inputs(227));
    layer0_outputs(9696) <= inputs(136);
    layer0_outputs(9697) <= not(inputs(20));
    layer0_outputs(9698) <= (inputs(7)) or (inputs(185));
    layer0_outputs(9699) <= (inputs(145)) or (inputs(25));
    layer0_outputs(9700) <= inputs(129);
    layer0_outputs(9701) <= not(inputs(208));
    layer0_outputs(9702) <= not(inputs(141)) or (inputs(23));
    layer0_outputs(9703) <= not(inputs(28)) or (inputs(240));
    layer0_outputs(9704) <= (inputs(33)) xor (inputs(4));
    layer0_outputs(9705) <= (inputs(213)) xor (inputs(224));
    layer0_outputs(9706) <= not((inputs(36)) xor (inputs(84)));
    layer0_outputs(9707) <= not((inputs(78)) or (inputs(3)));
    layer0_outputs(9708) <= not((inputs(155)) and (inputs(189)));
    layer0_outputs(9709) <= not(inputs(106));
    layer0_outputs(9710) <= not((inputs(86)) or (inputs(253)));
    layer0_outputs(9711) <= (inputs(47)) xor (inputs(168));
    layer0_outputs(9712) <= not(inputs(41)) or (inputs(80));
    layer0_outputs(9713) <= not((inputs(106)) xor (inputs(108)));
    layer0_outputs(9714) <= (inputs(12)) xor (inputs(72));
    layer0_outputs(9715) <= (inputs(196)) or (inputs(244));
    layer0_outputs(9716) <= (inputs(244)) and not (inputs(255));
    layer0_outputs(9717) <= not((inputs(103)) xor (inputs(154)));
    layer0_outputs(9718) <= (inputs(197)) and not (inputs(111));
    layer0_outputs(9719) <= (inputs(227)) and not (inputs(159));
    layer0_outputs(9720) <= not(inputs(26));
    layer0_outputs(9721) <= not((inputs(166)) or (inputs(34)));
    layer0_outputs(9722) <= (inputs(64)) xor (inputs(23));
    layer0_outputs(9723) <= (inputs(83)) and not (inputs(187));
    layer0_outputs(9724) <= not(inputs(146));
    layer0_outputs(9725) <= (inputs(54)) or (inputs(17));
    layer0_outputs(9726) <= (inputs(192)) xor (inputs(160));
    layer0_outputs(9727) <= not(inputs(90));
    layer0_outputs(9728) <= not((inputs(211)) or (inputs(208)));
    layer0_outputs(9729) <= not(inputs(78));
    layer0_outputs(9730) <= not(inputs(248));
    layer0_outputs(9731) <= (inputs(147)) or (inputs(149));
    layer0_outputs(9732) <= not(inputs(153));
    layer0_outputs(9733) <= (inputs(187)) and not (inputs(16));
    layer0_outputs(9734) <= not(inputs(100));
    layer0_outputs(9735) <= (inputs(49)) xor (inputs(43));
    layer0_outputs(9736) <= not(inputs(107));
    layer0_outputs(9737) <= (inputs(102)) xor (inputs(201));
    layer0_outputs(9738) <= (inputs(251)) or (inputs(175));
    layer0_outputs(9739) <= (inputs(193)) or (inputs(144));
    layer0_outputs(9740) <= (inputs(162)) xor (inputs(213));
    layer0_outputs(9741) <= not(inputs(1)) or (inputs(178));
    layer0_outputs(9742) <= not((inputs(106)) or (inputs(163)));
    layer0_outputs(9743) <= not(inputs(166));
    layer0_outputs(9744) <= not((inputs(117)) xor (inputs(222)));
    layer0_outputs(9745) <= not(inputs(227));
    layer0_outputs(9746) <= (inputs(76)) and not (inputs(84));
    layer0_outputs(9747) <= not((inputs(184)) or (inputs(79)));
    layer0_outputs(9748) <= not(inputs(5));
    layer0_outputs(9749) <= (inputs(37)) or (inputs(105));
    layer0_outputs(9750) <= (inputs(54)) or (inputs(191));
    layer0_outputs(9751) <= (inputs(11)) or (inputs(43));
    layer0_outputs(9752) <= (inputs(119)) and not (inputs(56));
    layer0_outputs(9753) <= not(inputs(163));
    layer0_outputs(9754) <= (inputs(47)) or (inputs(254));
    layer0_outputs(9755) <= not((inputs(182)) or (inputs(103)));
    layer0_outputs(9756) <= not((inputs(32)) xor (inputs(226)));
    layer0_outputs(9757) <= not((inputs(52)) or (inputs(112)));
    layer0_outputs(9758) <= (inputs(199)) and not (inputs(158));
    layer0_outputs(9759) <= not(inputs(134)) or (inputs(15));
    layer0_outputs(9760) <= (inputs(119)) and not (inputs(141));
    layer0_outputs(9761) <= inputs(38);
    layer0_outputs(9762) <= inputs(134);
    layer0_outputs(9763) <= not(inputs(239));
    layer0_outputs(9764) <= not(inputs(229));
    layer0_outputs(9765) <= (inputs(108)) and not (inputs(254));
    layer0_outputs(9766) <= not((inputs(206)) and (inputs(208)));
    layer0_outputs(9767) <= not(inputs(225));
    layer0_outputs(9768) <= inputs(88);
    layer0_outputs(9769) <= (inputs(54)) xor (inputs(48));
    layer0_outputs(9770) <= not((inputs(8)) xor (inputs(51)));
    layer0_outputs(9771) <= inputs(168);
    layer0_outputs(9772) <= not((inputs(222)) xor (inputs(211)));
    layer0_outputs(9773) <= (inputs(70)) xor (inputs(207));
    layer0_outputs(9774) <= not(inputs(19));
    layer0_outputs(9775) <= (inputs(176)) or (inputs(128));
    layer0_outputs(9776) <= inputs(244);
    layer0_outputs(9777) <= inputs(252);
    layer0_outputs(9778) <= inputs(130);
    layer0_outputs(9779) <= not(inputs(74));
    layer0_outputs(9780) <= not((inputs(84)) or (inputs(51)));
    layer0_outputs(9781) <= not((inputs(163)) and (inputs(48)));
    layer0_outputs(9782) <= not(inputs(33));
    layer0_outputs(9783) <= inputs(8);
    layer0_outputs(9784) <= not(inputs(67)) or (inputs(228));
    layer0_outputs(9785) <= not((inputs(209)) or (inputs(66)));
    layer0_outputs(9786) <= (inputs(65)) xor (inputs(51));
    layer0_outputs(9787) <= not(inputs(140));
    layer0_outputs(9788) <= not(inputs(203));
    layer0_outputs(9789) <= inputs(53);
    layer0_outputs(9790) <= not((inputs(38)) xor (inputs(30)));
    layer0_outputs(9791) <= not((inputs(5)) or (inputs(207)));
    layer0_outputs(9792) <= (inputs(137)) and (inputs(12));
    layer0_outputs(9793) <= (inputs(216)) and not (inputs(27));
    layer0_outputs(9794) <= (inputs(219)) or (inputs(172));
    layer0_outputs(9795) <= (inputs(82)) or (inputs(162));
    layer0_outputs(9796) <= (inputs(180)) xor (inputs(242));
    layer0_outputs(9797) <= inputs(82);
    layer0_outputs(9798) <= inputs(199);
    layer0_outputs(9799) <= not((inputs(219)) xor (inputs(66)));
    layer0_outputs(9800) <= inputs(99);
    layer0_outputs(9801) <= not((inputs(240)) or (inputs(124)));
    layer0_outputs(9802) <= not(inputs(58)) or (inputs(188));
    layer0_outputs(9803) <= '1';
    layer0_outputs(9804) <= not(inputs(60));
    layer0_outputs(9805) <= not(inputs(23)) or (inputs(131));
    layer0_outputs(9806) <= not((inputs(110)) and (inputs(49)));
    layer0_outputs(9807) <= not((inputs(90)) xor (inputs(127)));
    layer0_outputs(9808) <= (inputs(0)) and not (inputs(186));
    layer0_outputs(9809) <= (inputs(201)) or (inputs(181));
    layer0_outputs(9810) <= '0';
    layer0_outputs(9811) <= not((inputs(47)) or (inputs(250)));
    layer0_outputs(9812) <= not((inputs(35)) or (inputs(192)));
    layer0_outputs(9813) <= (inputs(231)) or (inputs(215));
    layer0_outputs(9814) <= inputs(21);
    layer0_outputs(9815) <= (inputs(128)) and not (inputs(245));
    layer0_outputs(9816) <= not(inputs(11));
    layer0_outputs(9817) <= not(inputs(101));
    layer0_outputs(9818) <= not((inputs(143)) or (inputs(125)));
    layer0_outputs(9819) <= not(inputs(249));
    layer0_outputs(9820) <= not((inputs(21)) xor (inputs(55)));
    layer0_outputs(9821) <= (inputs(221)) xor (inputs(135));
    layer0_outputs(9822) <= not(inputs(210));
    layer0_outputs(9823) <= not((inputs(134)) or (inputs(119)));
    layer0_outputs(9824) <= (inputs(170)) xor (inputs(171));
    layer0_outputs(9825) <= not(inputs(123));
    layer0_outputs(9826) <= (inputs(195)) or (inputs(220));
    layer0_outputs(9827) <= not((inputs(18)) or (inputs(150)));
    layer0_outputs(9828) <= (inputs(23)) or (inputs(220));
    layer0_outputs(9829) <= inputs(219);
    layer0_outputs(9830) <= (inputs(245)) and (inputs(25));
    layer0_outputs(9831) <= (inputs(151)) or (inputs(232));
    layer0_outputs(9832) <= not((inputs(250)) and (inputs(55)));
    layer0_outputs(9833) <= not(inputs(138)) or (inputs(101));
    layer0_outputs(9834) <= not(inputs(35));
    layer0_outputs(9835) <= not(inputs(132));
    layer0_outputs(9836) <= (inputs(121)) xor (inputs(71));
    layer0_outputs(9837) <= not((inputs(1)) xor (inputs(222)));
    layer0_outputs(9838) <= not((inputs(60)) or (inputs(165)));
    layer0_outputs(9839) <= (inputs(108)) or (inputs(20));
    layer0_outputs(9840) <= '0';
    layer0_outputs(9841) <= (inputs(149)) xor (inputs(235));
    layer0_outputs(9842) <= (inputs(165)) and not (inputs(113));
    layer0_outputs(9843) <= not((inputs(98)) or (inputs(27)));
    layer0_outputs(9844) <= not((inputs(82)) xor (inputs(48)));
    layer0_outputs(9845) <= not(inputs(248)) or (inputs(206));
    layer0_outputs(9846) <= not((inputs(133)) xor (inputs(161)));
    layer0_outputs(9847) <= not(inputs(44));
    layer0_outputs(9848) <= not((inputs(10)) or (inputs(61)));
    layer0_outputs(9849) <= not(inputs(43)) or (inputs(186));
    layer0_outputs(9850) <= not(inputs(135)) or (inputs(172));
    layer0_outputs(9851) <= not((inputs(219)) xor (inputs(80)));
    layer0_outputs(9852) <= (inputs(17)) or (inputs(255));
    layer0_outputs(9853) <= not((inputs(220)) or (inputs(120)));
    layer0_outputs(9854) <= not(inputs(247)) or (inputs(44));
    layer0_outputs(9855) <= (inputs(36)) and not (inputs(240));
    layer0_outputs(9856) <= not(inputs(223));
    layer0_outputs(9857) <= (inputs(13)) xor (inputs(17));
    layer0_outputs(9858) <= not(inputs(22));
    layer0_outputs(9859) <= (inputs(59)) xor (inputs(35));
    layer0_outputs(9860) <= not((inputs(211)) xor (inputs(111)));
    layer0_outputs(9861) <= inputs(193);
    layer0_outputs(9862) <= not((inputs(211)) or (inputs(238)));
    layer0_outputs(9863) <= (inputs(172)) or (inputs(69));
    layer0_outputs(9864) <= (inputs(109)) or (inputs(136));
    layer0_outputs(9865) <= not((inputs(148)) or (inputs(185)));
    layer0_outputs(9866) <= (inputs(115)) xor (inputs(36));
    layer0_outputs(9867) <= not(inputs(42));
    layer0_outputs(9868) <= (inputs(8)) and not (inputs(249));
    layer0_outputs(9869) <= (inputs(148)) or (inputs(98));
    layer0_outputs(9870) <= (inputs(152)) and not (inputs(58));
    layer0_outputs(9871) <= inputs(7);
    layer0_outputs(9872) <= (inputs(47)) xor (inputs(232));
    layer0_outputs(9873) <= not((inputs(138)) or (inputs(6)));
    layer0_outputs(9874) <= inputs(111);
    layer0_outputs(9875) <= not(inputs(43));
    layer0_outputs(9876) <= inputs(75);
    layer0_outputs(9877) <= not(inputs(0)) or (inputs(28));
    layer0_outputs(9878) <= not((inputs(86)) or (inputs(202)));
    layer0_outputs(9879) <= not((inputs(107)) or (inputs(55)));
    layer0_outputs(9880) <= inputs(161);
    layer0_outputs(9881) <= (inputs(169)) and not (inputs(15));
    layer0_outputs(9882) <= (inputs(207)) or (inputs(80));
    layer0_outputs(9883) <= (inputs(12)) and (inputs(46));
    layer0_outputs(9884) <= not(inputs(201)) or (inputs(123));
    layer0_outputs(9885) <= not((inputs(60)) or (inputs(96)));
    layer0_outputs(9886) <= not((inputs(152)) xor (inputs(194)));
    layer0_outputs(9887) <= not(inputs(198)) or (inputs(37));
    layer0_outputs(9888) <= not(inputs(6)) or (inputs(112));
    layer0_outputs(9889) <= inputs(230);
    layer0_outputs(9890) <= (inputs(194)) or (inputs(183));
    layer0_outputs(9891) <= (inputs(66)) and not (inputs(46));
    layer0_outputs(9892) <= not((inputs(23)) or (inputs(3)));
    layer0_outputs(9893) <= (inputs(118)) xor (inputs(178));
    layer0_outputs(9894) <= not((inputs(11)) and (inputs(13)));
    layer0_outputs(9895) <= not(inputs(56));
    layer0_outputs(9896) <= inputs(87);
    layer0_outputs(9897) <= not((inputs(31)) and (inputs(212)));
    layer0_outputs(9898) <= (inputs(148)) or (inputs(249));
    layer0_outputs(9899) <= not(inputs(235)) or (inputs(0));
    layer0_outputs(9900) <= (inputs(92)) and not (inputs(175));
    layer0_outputs(9901) <= not((inputs(10)) xor (inputs(60)));
    layer0_outputs(9902) <= inputs(89);
    layer0_outputs(9903) <= inputs(152);
    layer0_outputs(9904) <= not((inputs(10)) xor (inputs(39)));
    layer0_outputs(9905) <= not(inputs(41));
    layer0_outputs(9906) <= not((inputs(253)) and (inputs(159)));
    layer0_outputs(9907) <= (inputs(30)) and not (inputs(246));
    layer0_outputs(9908) <= inputs(216);
    layer0_outputs(9909) <= not(inputs(58));
    layer0_outputs(9910) <= inputs(23);
    layer0_outputs(9911) <= (inputs(123)) xor (inputs(125));
    layer0_outputs(9912) <= (inputs(121)) or (inputs(29));
    layer0_outputs(9913) <= not((inputs(17)) or (inputs(72)));
    layer0_outputs(9914) <= not(inputs(148));
    layer0_outputs(9915) <= not(inputs(181));
    layer0_outputs(9916) <= inputs(158);
    layer0_outputs(9917) <= not(inputs(41)) or (inputs(16));
    layer0_outputs(9918) <= (inputs(144)) or (inputs(128));
    layer0_outputs(9919) <= (inputs(190)) xor (inputs(142));
    layer0_outputs(9920) <= not((inputs(104)) xor (inputs(186)));
    layer0_outputs(9921) <= not(inputs(106));
    layer0_outputs(9922) <= not((inputs(74)) xor (inputs(42)));
    layer0_outputs(9923) <= inputs(168);
    layer0_outputs(9924) <= not(inputs(53));
    layer0_outputs(9925) <= inputs(56);
    layer0_outputs(9926) <= (inputs(124)) and (inputs(73));
    layer0_outputs(9927) <= (inputs(220)) and not (inputs(14));
    layer0_outputs(9928) <= not(inputs(147)) or (inputs(195));
    layer0_outputs(9929) <= not(inputs(52));
    layer0_outputs(9930) <= not(inputs(231)) or (inputs(224));
    layer0_outputs(9931) <= (inputs(230)) xor (inputs(123));
    layer0_outputs(9932) <= (inputs(73)) and not (inputs(19));
    layer0_outputs(9933) <= (inputs(188)) and not (inputs(125));
    layer0_outputs(9934) <= inputs(180);
    layer0_outputs(9935) <= not(inputs(19));
    layer0_outputs(9936) <= (inputs(117)) xor (inputs(254));
    layer0_outputs(9937) <= inputs(113);
    layer0_outputs(9938) <= not((inputs(16)) xor (inputs(69)));
    layer0_outputs(9939) <= (inputs(106)) and not (inputs(228));
    layer0_outputs(9940) <= (inputs(83)) xor (inputs(23));
    layer0_outputs(9941) <= not((inputs(196)) and (inputs(164)));
    layer0_outputs(9942) <= (inputs(131)) and not (inputs(249));
    layer0_outputs(9943) <= not(inputs(74));
    layer0_outputs(9944) <= inputs(157);
    layer0_outputs(9945) <= (inputs(71)) and not (inputs(35));
    layer0_outputs(9946) <= not((inputs(173)) and (inputs(162)));
    layer0_outputs(9947) <= not(inputs(91)) or (inputs(112));
    layer0_outputs(9948) <= not((inputs(62)) xor (inputs(78)));
    layer0_outputs(9949) <= inputs(122);
    layer0_outputs(9950) <= not(inputs(182));
    layer0_outputs(9951) <= not(inputs(246)) or (inputs(147));
    layer0_outputs(9952) <= inputs(56);
    layer0_outputs(9953) <= not(inputs(183));
    layer0_outputs(9954) <= not(inputs(149));
    layer0_outputs(9955) <= not((inputs(83)) or (inputs(131)));
    layer0_outputs(9956) <= (inputs(163)) or (inputs(1));
    layer0_outputs(9957) <= not((inputs(36)) or (inputs(136)));
    layer0_outputs(9958) <= not(inputs(106));
    layer0_outputs(9959) <= (inputs(86)) or (inputs(31));
    layer0_outputs(9960) <= (inputs(140)) and (inputs(228));
    layer0_outputs(9961) <= not((inputs(118)) and (inputs(65)));
    layer0_outputs(9962) <= not((inputs(205)) or (inputs(55)));
    layer0_outputs(9963) <= not(inputs(217));
    layer0_outputs(9964) <= (inputs(144)) xor (inputs(82));
    layer0_outputs(9965) <= not(inputs(171));
    layer0_outputs(9966) <= inputs(113);
    layer0_outputs(9967) <= (inputs(53)) and not (inputs(204));
    layer0_outputs(9968) <= not(inputs(166));
    layer0_outputs(9969) <= (inputs(168)) and not (inputs(48));
    layer0_outputs(9970) <= not(inputs(155)) or (inputs(140));
    layer0_outputs(9971) <= not(inputs(68));
    layer0_outputs(9972) <= (inputs(59)) or (inputs(125));
    layer0_outputs(9973) <= (inputs(44)) xor (inputs(99));
    layer0_outputs(9974) <= (inputs(56)) and not (inputs(120));
    layer0_outputs(9975) <= (inputs(77)) and not (inputs(251));
    layer0_outputs(9976) <= (inputs(138)) or (inputs(187));
    layer0_outputs(9977) <= not(inputs(104));
    layer0_outputs(9978) <= not(inputs(110));
    layer0_outputs(9979) <= not(inputs(170)) or (inputs(36));
    layer0_outputs(9980) <= (inputs(138)) and (inputs(75));
    layer0_outputs(9981) <= inputs(175);
    layer0_outputs(9982) <= not((inputs(134)) or (inputs(185)));
    layer0_outputs(9983) <= not((inputs(180)) and (inputs(200)));
    layer0_outputs(9984) <= (inputs(154)) or (inputs(120));
    layer0_outputs(9985) <= inputs(230);
    layer0_outputs(9986) <= not(inputs(23));
    layer0_outputs(9987) <= (inputs(83)) or (inputs(189));
    layer0_outputs(9988) <= (inputs(225)) and not (inputs(78));
    layer0_outputs(9989) <= not((inputs(137)) or (inputs(14)));
    layer0_outputs(9990) <= not((inputs(50)) xor (inputs(150)));
    layer0_outputs(9991) <= (inputs(136)) and not (inputs(111));
    layer0_outputs(9992) <= (inputs(72)) and not (inputs(253));
    layer0_outputs(9993) <= not((inputs(87)) xor (inputs(52)));
    layer0_outputs(9994) <= inputs(30);
    layer0_outputs(9995) <= inputs(84);
    layer0_outputs(9996) <= not((inputs(255)) xor (inputs(240)));
    layer0_outputs(9997) <= (inputs(125)) xor (inputs(239));
    layer0_outputs(9998) <= (inputs(145)) or (inputs(50));
    layer0_outputs(9999) <= (inputs(203)) and not (inputs(16));
    layer0_outputs(10000) <= (inputs(110)) or (inputs(138));
    layer0_outputs(10001) <= not((inputs(92)) xor (inputs(225)));
    layer0_outputs(10002) <= inputs(131);
    layer0_outputs(10003) <= not(inputs(94));
    layer0_outputs(10004) <= (inputs(196)) or (inputs(245));
    layer0_outputs(10005) <= (inputs(127)) xor (inputs(104));
    layer0_outputs(10006) <= not((inputs(246)) or (inputs(213)));
    layer0_outputs(10007) <= not(inputs(150));
    layer0_outputs(10008) <= not((inputs(254)) xor (inputs(46)));
    layer0_outputs(10009) <= (inputs(235)) xor (inputs(105));
    layer0_outputs(10010) <= '0';
    layer0_outputs(10011) <= not(inputs(80));
    layer0_outputs(10012) <= not(inputs(91));
    layer0_outputs(10013) <= inputs(31);
    layer0_outputs(10014) <= inputs(118);
    layer0_outputs(10015) <= not(inputs(35)) or (inputs(200));
    layer0_outputs(10016) <= not(inputs(242)) or (inputs(130));
    layer0_outputs(10017) <= (inputs(143)) or (inputs(198));
    layer0_outputs(10018) <= inputs(146);
    layer0_outputs(10019) <= (inputs(180)) and not (inputs(90));
    layer0_outputs(10020) <= not(inputs(14));
    layer0_outputs(10021) <= (inputs(33)) or (inputs(77));
    layer0_outputs(10022) <= (inputs(150)) and not (inputs(49));
    layer0_outputs(10023) <= (inputs(240)) or (inputs(226));
    layer0_outputs(10024) <= (inputs(184)) or (inputs(113));
    layer0_outputs(10025) <= inputs(225);
    layer0_outputs(10026) <= (inputs(209)) and not (inputs(224));
    layer0_outputs(10027) <= inputs(28);
    layer0_outputs(10028) <= (inputs(46)) xor (inputs(247));
    layer0_outputs(10029) <= inputs(89);
    layer0_outputs(10030) <= not((inputs(195)) or (inputs(132)));
    layer0_outputs(10031) <= (inputs(254)) xor (inputs(244));
    layer0_outputs(10032) <= not((inputs(72)) xor (inputs(32)));
    layer0_outputs(10033) <= (inputs(169)) or (inputs(46));
    layer0_outputs(10034) <= inputs(222);
    layer0_outputs(10035) <= not((inputs(68)) xor (inputs(159)));
    layer0_outputs(10036) <= inputs(179);
    layer0_outputs(10037) <= (inputs(113)) or (inputs(184));
    layer0_outputs(10038) <= inputs(169);
    layer0_outputs(10039) <= not(inputs(176)) or (inputs(150));
    layer0_outputs(10040) <= (inputs(235)) xor (inputs(13));
    layer0_outputs(10041) <= not(inputs(24));
    layer0_outputs(10042) <= (inputs(255)) and (inputs(161));
    layer0_outputs(10043) <= not(inputs(143));
    layer0_outputs(10044) <= (inputs(181)) or (inputs(1));
    layer0_outputs(10045) <= not(inputs(59));
    layer0_outputs(10046) <= inputs(99);
    layer0_outputs(10047) <= not(inputs(231)) or (inputs(50));
    layer0_outputs(10048) <= not(inputs(54));
    layer0_outputs(10049) <= (inputs(255)) xor (inputs(57));
    layer0_outputs(10050) <= (inputs(161)) or (inputs(189));
    layer0_outputs(10051) <= not((inputs(101)) xor (inputs(86)));
    layer0_outputs(10052) <= (inputs(46)) and not (inputs(254));
    layer0_outputs(10053) <= (inputs(93)) or (inputs(237));
    layer0_outputs(10054) <= not((inputs(212)) or (inputs(81)));
    layer0_outputs(10055) <= inputs(20);
    layer0_outputs(10056) <= (inputs(199)) xor (inputs(224));
    layer0_outputs(10057) <= not((inputs(175)) or (inputs(180)));
    layer0_outputs(10058) <= inputs(24);
    layer0_outputs(10059) <= not((inputs(175)) or (inputs(163)));
    layer0_outputs(10060) <= inputs(77);
    layer0_outputs(10061) <= (inputs(209)) or (inputs(158));
    layer0_outputs(10062) <= inputs(100);
    layer0_outputs(10063) <= not(inputs(230));
    layer0_outputs(10064) <= (inputs(190)) and not (inputs(84));
    layer0_outputs(10065) <= not(inputs(168)) or (inputs(87));
    layer0_outputs(10066) <= not((inputs(149)) xor (inputs(192)));
    layer0_outputs(10067) <= (inputs(20)) xor (inputs(27));
    layer0_outputs(10068) <= not(inputs(248));
    layer0_outputs(10069) <= not(inputs(231));
    layer0_outputs(10070) <= not((inputs(52)) or (inputs(154)));
    layer0_outputs(10071) <= (inputs(160)) xor (inputs(117));
    layer0_outputs(10072) <= not(inputs(22));
    layer0_outputs(10073) <= not(inputs(3));
    layer0_outputs(10074) <= (inputs(45)) and (inputs(121));
    layer0_outputs(10075) <= not(inputs(236));
    layer0_outputs(10076) <= not(inputs(103));
    layer0_outputs(10077) <= not((inputs(41)) and (inputs(132)));
    layer0_outputs(10078) <= not(inputs(94)) or (inputs(2));
    layer0_outputs(10079) <= not(inputs(246)) or (inputs(29));
    layer0_outputs(10080) <= (inputs(69)) xor (inputs(184));
    layer0_outputs(10081) <= (inputs(198)) xor (inputs(205));
    layer0_outputs(10082) <= not(inputs(182));
    layer0_outputs(10083) <= not(inputs(232));
    layer0_outputs(10084) <= not(inputs(55)) or (inputs(235));
    layer0_outputs(10085) <= not(inputs(148));
    layer0_outputs(10086) <= not((inputs(187)) xor (inputs(152)));
    layer0_outputs(10087) <= (inputs(127)) or (inputs(6));
    layer0_outputs(10088) <= not(inputs(203));
    layer0_outputs(10089) <= inputs(246);
    layer0_outputs(10090) <= not(inputs(129));
    layer0_outputs(10091) <= (inputs(177)) and not (inputs(35));
    layer0_outputs(10092) <= (inputs(153)) and not (inputs(162));
    layer0_outputs(10093) <= inputs(83);
    layer0_outputs(10094) <= not(inputs(137));
    layer0_outputs(10095) <= not((inputs(219)) and (inputs(217)));
    layer0_outputs(10096) <= inputs(44);
    layer0_outputs(10097) <= not(inputs(34));
    layer0_outputs(10098) <= inputs(212);
    layer0_outputs(10099) <= not((inputs(247)) and (inputs(164)));
    layer0_outputs(10100) <= not((inputs(80)) xor (inputs(134)));
    layer0_outputs(10101) <= not(inputs(158));
    layer0_outputs(10102) <= not((inputs(212)) xor (inputs(243)));
    layer0_outputs(10103) <= not(inputs(23)) or (inputs(222));
    layer0_outputs(10104) <= not(inputs(32));
    layer0_outputs(10105) <= not(inputs(227)) or (inputs(109));
    layer0_outputs(10106) <= inputs(162);
    layer0_outputs(10107) <= not((inputs(149)) or (inputs(67)));
    layer0_outputs(10108) <= not((inputs(43)) xor (inputs(102)));
    layer0_outputs(10109) <= (inputs(235)) and (inputs(110));
    layer0_outputs(10110) <= not(inputs(253));
    layer0_outputs(10111) <= not(inputs(248)) or (inputs(114));
    layer0_outputs(10112) <= not(inputs(141));
    layer0_outputs(10113) <= not(inputs(17));
    layer0_outputs(10114) <= not((inputs(77)) or (inputs(37)));
    layer0_outputs(10115) <= not((inputs(0)) or (inputs(122)));
    layer0_outputs(10116) <= (inputs(213)) and (inputs(217));
    layer0_outputs(10117) <= not((inputs(183)) xor (inputs(31)));
    layer0_outputs(10118) <= not(inputs(90));
    layer0_outputs(10119) <= inputs(67);
    layer0_outputs(10120) <= (inputs(49)) and not (inputs(57));
    layer0_outputs(10121) <= (inputs(42)) xor (inputs(129));
    layer0_outputs(10122) <= inputs(79);
    layer0_outputs(10123) <= (inputs(57)) and (inputs(105));
    layer0_outputs(10124) <= (inputs(144)) xor (inputs(211));
    layer0_outputs(10125) <= (inputs(124)) and (inputs(108));
    layer0_outputs(10126) <= not((inputs(28)) xor (inputs(72)));
    layer0_outputs(10127) <= (inputs(215)) xor (inputs(226));
    layer0_outputs(10128) <= not(inputs(76));
    layer0_outputs(10129) <= not(inputs(27)) or (inputs(145));
    layer0_outputs(10130) <= (inputs(7)) xor (inputs(181));
    layer0_outputs(10131) <= not(inputs(181));
    layer0_outputs(10132) <= not((inputs(79)) or (inputs(42)));
    layer0_outputs(10133) <= not((inputs(109)) xor (inputs(32)));
    layer0_outputs(10134) <= not(inputs(43));
    layer0_outputs(10135) <= inputs(153);
    layer0_outputs(10136) <= (inputs(52)) or (inputs(13));
    layer0_outputs(10137) <= not(inputs(18));
    layer0_outputs(10138) <= not((inputs(67)) or (inputs(158)));
    layer0_outputs(10139) <= not((inputs(114)) or (inputs(157)));
    layer0_outputs(10140) <= not(inputs(58));
    layer0_outputs(10141) <= not((inputs(185)) or (inputs(208)));
    layer0_outputs(10142) <= (inputs(187)) xor (inputs(84));
    layer0_outputs(10143) <= (inputs(86)) or (inputs(82));
    layer0_outputs(10144) <= not(inputs(170)) or (inputs(91));
    layer0_outputs(10145) <= (inputs(187)) and not (inputs(93));
    layer0_outputs(10146) <= not(inputs(131));
    layer0_outputs(10147) <= (inputs(137)) xor (inputs(218));
    layer0_outputs(10148) <= inputs(227);
    layer0_outputs(10149) <= (inputs(41)) or (inputs(6));
    layer0_outputs(10150) <= inputs(125);
    layer0_outputs(10151) <= (inputs(192)) and not (inputs(59));
    layer0_outputs(10152) <= not((inputs(66)) xor (inputs(106)));
    layer0_outputs(10153) <= not(inputs(108));
    layer0_outputs(10154) <= '0';
    layer0_outputs(10155) <= (inputs(143)) or (inputs(252));
    layer0_outputs(10156) <= not((inputs(118)) xor (inputs(172)));
    layer0_outputs(10157) <= inputs(70);
    layer0_outputs(10158) <= (inputs(20)) xor (inputs(222));
    layer0_outputs(10159) <= inputs(35);
    layer0_outputs(10160) <= not(inputs(232)) or (inputs(73));
    layer0_outputs(10161) <= not((inputs(149)) or (inputs(66)));
    layer0_outputs(10162) <= inputs(163);
    layer0_outputs(10163) <= not((inputs(148)) or (inputs(140)));
    layer0_outputs(10164) <= not(inputs(232)) or (inputs(123));
    layer0_outputs(10165) <= not(inputs(128));
    layer0_outputs(10166) <= not((inputs(99)) and (inputs(83)));
    layer0_outputs(10167) <= (inputs(59)) and not (inputs(241));
    layer0_outputs(10168) <= inputs(118);
    layer0_outputs(10169) <= (inputs(123)) or (inputs(16));
    layer0_outputs(10170) <= not((inputs(91)) or (inputs(145)));
    layer0_outputs(10171) <= inputs(241);
    layer0_outputs(10172) <= not((inputs(8)) xor (inputs(225)));
    layer0_outputs(10173) <= not(inputs(179)) or (inputs(16));
    layer0_outputs(10174) <= (inputs(196)) and not (inputs(63));
    layer0_outputs(10175) <= not(inputs(38)) or (inputs(175));
    layer0_outputs(10176) <= inputs(55);
    layer0_outputs(10177) <= not((inputs(240)) xor (inputs(136)));
    layer0_outputs(10178) <= inputs(112);
    layer0_outputs(10179) <= not((inputs(13)) or (inputs(190)));
    layer0_outputs(10180) <= not(inputs(110));
    layer0_outputs(10181) <= not(inputs(120)) or (inputs(2));
    layer0_outputs(10182) <= '0';
    layer0_outputs(10183) <= not((inputs(253)) xor (inputs(207)));
    layer0_outputs(10184) <= not(inputs(89)) or (inputs(19));
    layer0_outputs(10185) <= (inputs(243)) or (inputs(86));
    layer0_outputs(10186) <= '1';
    layer0_outputs(10187) <= not((inputs(134)) and (inputs(216)));
    layer0_outputs(10188) <= not((inputs(126)) xor (inputs(79)));
    layer0_outputs(10189) <= not(inputs(97));
    layer0_outputs(10190) <= not(inputs(43)) or (inputs(173));
    layer0_outputs(10191) <= (inputs(148)) xor (inputs(122));
    layer0_outputs(10192) <= not(inputs(136)) or (inputs(73));
    layer0_outputs(10193) <= '0';
    layer0_outputs(10194) <= inputs(19);
    layer0_outputs(10195) <= (inputs(108)) and (inputs(71));
    layer0_outputs(10196) <= (inputs(175)) or (inputs(133));
    layer0_outputs(10197) <= (inputs(56)) and not (inputs(254));
    layer0_outputs(10198) <= not((inputs(37)) and (inputs(187)));
    layer0_outputs(10199) <= (inputs(176)) xor (inputs(167));
    layer0_outputs(10200) <= not((inputs(194)) or (inputs(180)));
    layer0_outputs(10201) <= not(inputs(187)) or (inputs(80));
    layer0_outputs(10202) <= not(inputs(162)) or (inputs(114));
    layer0_outputs(10203) <= not((inputs(31)) or (inputs(114)));
    layer0_outputs(10204) <= inputs(15);
    layer0_outputs(10205) <= (inputs(42)) xor (inputs(31));
    layer0_outputs(10206) <= '1';
    layer0_outputs(10207) <= inputs(46);
    layer0_outputs(10208) <= not(inputs(77));
    layer0_outputs(10209) <= (inputs(161)) or (inputs(194));
    layer0_outputs(10210) <= (inputs(199)) and not (inputs(243));
    layer0_outputs(10211) <= not((inputs(75)) or (inputs(74)));
    layer0_outputs(10212) <= (inputs(64)) or (inputs(178));
    layer0_outputs(10213) <= not((inputs(36)) xor (inputs(100)));
    layer0_outputs(10214) <= inputs(93);
    layer0_outputs(10215) <= not(inputs(29));
    layer0_outputs(10216) <= (inputs(230)) or (inputs(78));
    layer0_outputs(10217) <= not(inputs(112));
    layer0_outputs(10218) <= not((inputs(71)) xor (inputs(148)));
    layer0_outputs(10219) <= (inputs(67)) or (inputs(113));
    layer0_outputs(10220) <= not((inputs(91)) xor (inputs(93)));
    layer0_outputs(10221) <= not((inputs(41)) or (inputs(175)));
    layer0_outputs(10222) <= not((inputs(61)) or (inputs(47)));
    layer0_outputs(10223) <= not(inputs(122));
    layer0_outputs(10224) <= not((inputs(157)) xor (inputs(103)));
    layer0_outputs(10225) <= (inputs(219)) xor (inputs(141));
    layer0_outputs(10226) <= inputs(140);
    layer0_outputs(10227) <= not(inputs(57));
    layer0_outputs(10228) <= not((inputs(108)) and (inputs(214)));
    layer0_outputs(10229) <= not(inputs(187));
    layer0_outputs(10230) <= (inputs(153)) xor (inputs(43));
    layer0_outputs(10231) <= (inputs(66)) and not (inputs(191));
    layer0_outputs(10232) <= (inputs(96)) or (inputs(149));
    layer0_outputs(10233) <= not((inputs(19)) xor (inputs(87)));
    layer0_outputs(10234) <= (inputs(183)) or (inputs(220));
    layer0_outputs(10235) <= inputs(164);
    layer0_outputs(10236) <= not(inputs(24)) or (inputs(165));
    layer0_outputs(10237) <= not((inputs(20)) or (inputs(77)));
    layer0_outputs(10238) <= not(inputs(74));
    layer0_outputs(10239) <= (inputs(15)) xor (inputs(98));
    layer0_outputs(10240) <= (inputs(7)) or (inputs(237));
    layer0_outputs(10241) <= not(inputs(133)) or (inputs(205));
    layer0_outputs(10242) <= (inputs(177)) or (inputs(179));
    layer0_outputs(10243) <= (inputs(10)) xor (inputs(244));
    layer0_outputs(10244) <= not((inputs(73)) or (inputs(216)));
    layer0_outputs(10245) <= inputs(8);
    layer0_outputs(10246) <= inputs(151);
    layer0_outputs(10247) <= inputs(120);
    layer0_outputs(10248) <= (inputs(199)) and not (inputs(219));
    layer0_outputs(10249) <= not(inputs(42)) or (inputs(223));
    layer0_outputs(10250) <= (inputs(20)) or (inputs(8));
    layer0_outputs(10251) <= not(inputs(244)) or (inputs(112));
    layer0_outputs(10252) <= not((inputs(30)) or (inputs(157)));
    layer0_outputs(10253) <= not(inputs(86)) or (inputs(110));
    layer0_outputs(10254) <= inputs(119);
    layer0_outputs(10255) <= '0';
    layer0_outputs(10256) <= not((inputs(96)) xor (inputs(88)));
    layer0_outputs(10257) <= (inputs(176)) and not (inputs(31));
    layer0_outputs(10258) <= not(inputs(184));
    layer0_outputs(10259) <= not(inputs(75));
    layer0_outputs(10260) <= not((inputs(168)) xor (inputs(138)));
    layer0_outputs(10261) <= not(inputs(10));
    layer0_outputs(10262) <= not(inputs(161)) or (inputs(237));
    layer0_outputs(10263) <= (inputs(207)) and not (inputs(13));
    layer0_outputs(10264) <= not(inputs(191));
    layer0_outputs(10265) <= not(inputs(52));
    layer0_outputs(10266) <= not((inputs(89)) or (inputs(62)));
    layer0_outputs(10267) <= (inputs(189)) xor (inputs(24));
    layer0_outputs(10268) <= (inputs(49)) xor (inputs(53));
    layer0_outputs(10269) <= not(inputs(61));
    layer0_outputs(10270) <= (inputs(160)) or (inputs(201));
    layer0_outputs(10271) <= (inputs(160)) or (inputs(125));
    layer0_outputs(10272) <= not(inputs(203)) or (inputs(3));
    layer0_outputs(10273) <= not(inputs(151));
    layer0_outputs(10274) <= not((inputs(163)) or (inputs(91)));
    layer0_outputs(10275) <= (inputs(173)) and not (inputs(159));
    layer0_outputs(10276) <= inputs(45);
    layer0_outputs(10277) <= inputs(35);
    layer0_outputs(10278) <= not((inputs(82)) or (inputs(123)));
    layer0_outputs(10279) <= not(inputs(130)) or (inputs(220));
    layer0_outputs(10280) <= not((inputs(223)) xor (inputs(172)));
    layer0_outputs(10281) <= (inputs(93)) or (inputs(143));
    layer0_outputs(10282) <= not((inputs(59)) or (inputs(58)));
    layer0_outputs(10283) <= (inputs(243)) and not (inputs(105));
    layer0_outputs(10284) <= (inputs(29)) and not (inputs(124));
    layer0_outputs(10285) <= inputs(66);
    layer0_outputs(10286) <= '0';
    layer0_outputs(10287) <= not(inputs(194)) or (inputs(150));
    layer0_outputs(10288) <= not(inputs(106));
    layer0_outputs(10289) <= (inputs(253)) or (inputs(233));
    layer0_outputs(10290) <= inputs(69);
    layer0_outputs(10291) <= (inputs(230)) and not (inputs(59));
    layer0_outputs(10292) <= not(inputs(20));
    layer0_outputs(10293) <= (inputs(216)) and not (inputs(44));
    layer0_outputs(10294) <= (inputs(17)) or (inputs(75));
    layer0_outputs(10295) <= inputs(144);
    layer0_outputs(10296) <= inputs(18);
    layer0_outputs(10297) <= (inputs(218)) xor (inputs(154));
    layer0_outputs(10298) <= inputs(148);
    layer0_outputs(10299) <= (inputs(54)) xor (inputs(101));
    layer0_outputs(10300) <= not((inputs(141)) xor (inputs(195)));
    layer0_outputs(10301) <= inputs(180);
    layer0_outputs(10302) <= inputs(200);
    layer0_outputs(10303) <= not(inputs(12));
    layer0_outputs(10304) <= not((inputs(141)) xor (inputs(215)));
    layer0_outputs(10305) <= not((inputs(134)) xor (inputs(152)));
    layer0_outputs(10306) <= not((inputs(50)) xor (inputs(213)));
    layer0_outputs(10307) <= (inputs(14)) or (inputs(47));
    layer0_outputs(10308) <= (inputs(74)) xor (inputs(47));
    layer0_outputs(10309) <= (inputs(57)) xor (inputs(55));
    layer0_outputs(10310) <= inputs(1);
    layer0_outputs(10311) <= (inputs(108)) and not (inputs(244));
    layer0_outputs(10312) <= not(inputs(42));
    layer0_outputs(10313) <= (inputs(187)) and not (inputs(71));
    layer0_outputs(10314) <= not(inputs(176)) or (inputs(49));
    layer0_outputs(10315) <= not(inputs(147));
    layer0_outputs(10316) <= inputs(63);
    layer0_outputs(10317) <= not(inputs(202)) or (inputs(247));
    layer0_outputs(10318) <= not((inputs(47)) and (inputs(63)));
    layer0_outputs(10319) <= not(inputs(21));
    layer0_outputs(10320) <= inputs(108);
    layer0_outputs(10321) <= (inputs(101)) and not (inputs(111));
    layer0_outputs(10322) <= inputs(102);
    layer0_outputs(10323) <= (inputs(254)) or (inputs(17));
    layer0_outputs(10324) <= not(inputs(102));
    layer0_outputs(10325) <= not(inputs(20));
    layer0_outputs(10326) <= inputs(252);
    layer0_outputs(10327) <= (inputs(230)) and not (inputs(158));
    layer0_outputs(10328) <= (inputs(79)) or (inputs(61));
    layer0_outputs(10329) <= not((inputs(189)) xor (inputs(209)));
    layer0_outputs(10330) <= not(inputs(238));
    layer0_outputs(10331) <= (inputs(158)) and not (inputs(128));
    layer0_outputs(10332) <= inputs(113);
    layer0_outputs(10333) <= (inputs(189)) or (inputs(172));
    layer0_outputs(10334) <= not((inputs(153)) and (inputs(37)));
    layer0_outputs(10335) <= (inputs(139)) and (inputs(182));
    layer0_outputs(10336) <= (inputs(10)) and not (inputs(208));
    layer0_outputs(10337) <= (inputs(95)) or (inputs(12));
    layer0_outputs(10338) <= not((inputs(206)) or (inputs(209)));
    layer0_outputs(10339) <= '1';
    layer0_outputs(10340) <= inputs(64);
    layer0_outputs(10341) <= not((inputs(86)) or (inputs(89)));
    layer0_outputs(10342) <= not((inputs(226)) xor (inputs(43)));
    layer0_outputs(10343) <= not(inputs(152));
    layer0_outputs(10344) <= (inputs(227)) and not (inputs(127));
    layer0_outputs(10345) <= inputs(145);
    layer0_outputs(10346) <= inputs(45);
    layer0_outputs(10347) <= inputs(105);
    layer0_outputs(10348) <= not((inputs(36)) or (inputs(15)));
    layer0_outputs(10349) <= not((inputs(223)) or (inputs(90)));
    layer0_outputs(10350) <= (inputs(205)) or (inputs(200));
    layer0_outputs(10351) <= (inputs(150)) xor (inputs(161));
    layer0_outputs(10352) <= inputs(113);
    layer0_outputs(10353) <= (inputs(223)) or (inputs(88));
    layer0_outputs(10354) <= (inputs(155)) or (inputs(192));
    layer0_outputs(10355) <= not((inputs(205)) or (inputs(25)));
    layer0_outputs(10356) <= not(inputs(249));
    layer0_outputs(10357) <= inputs(213);
    layer0_outputs(10358) <= not(inputs(229));
    layer0_outputs(10359) <= (inputs(117)) and not (inputs(242));
    layer0_outputs(10360) <= not((inputs(222)) xor (inputs(89)));
    layer0_outputs(10361) <= not((inputs(94)) or (inputs(160)));
    layer0_outputs(10362) <= not(inputs(23)) or (inputs(85));
    layer0_outputs(10363) <= inputs(25);
    layer0_outputs(10364) <= not((inputs(229)) or (inputs(226)));
    layer0_outputs(10365) <= not(inputs(122));
    layer0_outputs(10366) <= not(inputs(102)) or (inputs(47));
    layer0_outputs(10367) <= not(inputs(24)) or (inputs(190));
    layer0_outputs(10368) <= not(inputs(148)) or (inputs(141));
    layer0_outputs(10369) <= (inputs(72)) xor (inputs(126));
    layer0_outputs(10370) <= (inputs(143)) or (inputs(76));
    layer0_outputs(10371) <= not((inputs(38)) or (inputs(16)));
    layer0_outputs(10372) <= not(inputs(108));
    layer0_outputs(10373) <= not((inputs(220)) xor (inputs(171)));
    layer0_outputs(10374) <= '1';
    layer0_outputs(10375) <= (inputs(54)) or (inputs(222));
    layer0_outputs(10376) <= (inputs(184)) and not (inputs(128));
    layer0_outputs(10377) <= not((inputs(116)) or (inputs(103)));
    layer0_outputs(10378) <= not((inputs(28)) and (inputs(226)));
    layer0_outputs(10379) <= not(inputs(20));
    layer0_outputs(10380) <= not(inputs(216));
    layer0_outputs(10381) <= '1';
    layer0_outputs(10382) <= inputs(114);
    layer0_outputs(10383) <= (inputs(69)) and not (inputs(64));
    layer0_outputs(10384) <= (inputs(75)) xor (inputs(174));
    layer0_outputs(10385) <= not(inputs(26));
    layer0_outputs(10386) <= not((inputs(177)) or (inputs(230)));
    layer0_outputs(10387) <= not(inputs(188)) or (inputs(10));
    layer0_outputs(10388) <= not((inputs(23)) xor (inputs(211)));
    layer0_outputs(10389) <= not(inputs(98));
    layer0_outputs(10390) <= not(inputs(26)) or (inputs(206));
    layer0_outputs(10391) <= not((inputs(136)) xor (inputs(74)));
    layer0_outputs(10392) <= (inputs(152)) and (inputs(200));
    layer0_outputs(10393) <= (inputs(222)) xor (inputs(189));
    layer0_outputs(10394) <= not(inputs(248)) or (inputs(123));
    layer0_outputs(10395) <= inputs(93);
    layer0_outputs(10396) <= (inputs(123)) and (inputs(27));
    layer0_outputs(10397) <= inputs(78);
    layer0_outputs(10398) <= (inputs(248)) or (inputs(176));
    layer0_outputs(10399) <= inputs(249);
    layer0_outputs(10400) <= (inputs(4)) and (inputs(135));
    layer0_outputs(10401) <= not((inputs(75)) xor (inputs(240)));
    layer0_outputs(10402) <= not((inputs(63)) xor (inputs(47)));
    layer0_outputs(10403) <= not((inputs(173)) xor (inputs(197)));
    layer0_outputs(10404) <= not((inputs(39)) or (inputs(34)));
    layer0_outputs(10405) <= not((inputs(20)) xor (inputs(155)));
    layer0_outputs(10406) <= (inputs(146)) or (inputs(235));
    layer0_outputs(10407) <= (inputs(160)) or (inputs(33));
    layer0_outputs(10408) <= (inputs(205)) or (inputs(115));
    layer0_outputs(10409) <= not(inputs(211)) or (inputs(56));
    layer0_outputs(10410) <= (inputs(106)) or (inputs(157));
    layer0_outputs(10411) <= (inputs(50)) xor (inputs(188));
    layer0_outputs(10412) <= (inputs(233)) and not (inputs(125));
    layer0_outputs(10413) <= not((inputs(56)) xor (inputs(224)));
    layer0_outputs(10414) <= not(inputs(113));
    layer0_outputs(10415) <= not((inputs(30)) xor (inputs(239)));
    layer0_outputs(10416) <= (inputs(72)) or (inputs(42));
    layer0_outputs(10417) <= (inputs(187)) and not (inputs(73));
    layer0_outputs(10418) <= not(inputs(51));
    layer0_outputs(10419) <= (inputs(102)) or (inputs(242));
    layer0_outputs(10420) <= (inputs(223)) xor (inputs(122));
    layer0_outputs(10421) <= (inputs(59)) or (inputs(129));
    layer0_outputs(10422) <= (inputs(195)) and not (inputs(7));
    layer0_outputs(10423) <= (inputs(116)) or (inputs(128));
    layer0_outputs(10424) <= inputs(23);
    layer0_outputs(10425) <= not((inputs(203)) and (inputs(218)));
    layer0_outputs(10426) <= (inputs(8)) xor (inputs(164));
    layer0_outputs(10427) <= (inputs(225)) and not (inputs(137));
    layer0_outputs(10428) <= not(inputs(182));
    layer0_outputs(10429) <= inputs(116);
    layer0_outputs(10430) <= inputs(204);
    layer0_outputs(10431) <= inputs(163);
    layer0_outputs(10432) <= not(inputs(215));
    layer0_outputs(10433) <= not(inputs(45)) or (inputs(137));
    layer0_outputs(10434) <= not(inputs(41)) or (inputs(158));
    layer0_outputs(10435) <= (inputs(200)) and not (inputs(226));
    layer0_outputs(10436) <= not((inputs(154)) xor (inputs(138)));
    layer0_outputs(10437) <= inputs(170);
    layer0_outputs(10438) <= not((inputs(121)) or (inputs(67)));
    layer0_outputs(10439) <= (inputs(157)) or (inputs(109));
    layer0_outputs(10440) <= not(inputs(63));
    layer0_outputs(10441) <= inputs(230);
    layer0_outputs(10442) <= not((inputs(104)) or (inputs(78)));
    layer0_outputs(10443) <= not((inputs(66)) or (inputs(133)));
    layer0_outputs(10444) <= not((inputs(233)) xor (inputs(215)));
    layer0_outputs(10445) <= not((inputs(141)) xor (inputs(119)));
    layer0_outputs(10446) <= not((inputs(51)) xor (inputs(23)));
    layer0_outputs(10447) <= (inputs(16)) and not (inputs(9));
    layer0_outputs(10448) <= inputs(227);
    layer0_outputs(10449) <= inputs(196);
    layer0_outputs(10450) <= not(inputs(222)) or (inputs(159));
    layer0_outputs(10451) <= (inputs(116)) and not (inputs(207));
    layer0_outputs(10452) <= (inputs(78)) and (inputs(142));
    layer0_outputs(10453) <= not((inputs(135)) or (inputs(194)));
    layer0_outputs(10454) <= inputs(129);
    layer0_outputs(10455) <= '1';
    layer0_outputs(10456) <= not((inputs(0)) or (inputs(30)));
    layer0_outputs(10457) <= not(inputs(150)) or (inputs(192));
    layer0_outputs(10458) <= (inputs(88)) and not (inputs(48));
    layer0_outputs(10459) <= not(inputs(200));
    layer0_outputs(10460) <= (inputs(46)) and not (inputs(148));
    layer0_outputs(10461) <= (inputs(134)) and not (inputs(139));
    layer0_outputs(10462) <= not((inputs(199)) or (inputs(134)));
    layer0_outputs(10463) <= (inputs(8)) xor (inputs(112));
    layer0_outputs(10464) <= not(inputs(45));
    layer0_outputs(10465) <= not((inputs(189)) xor (inputs(233)));
    layer0_outputs(10466) <= inputs(165);
    layer0_outputs(10467) <= not((inputs(52)) and (inputs(41)));
    layer0_outputs(10468) <= not(inputs(23));
    layer0_outputs(10469) <= not((inputs(207)) xor (inputs(127)));
    layer0_outputs(10470) <= not((inputs(118)) xor (inputs(179)));
    layer0_outputs(10471) <= not(inputs(236)) or (inputs(1));
    layer0_outputs(10472) <= (inputs(147)) and not (inputs(15));
    layer0_outputs(10473) <= (inputs(123)) and not (inputs(21));
    layer0_outputs(10474) <= not(inputs(118)) or (inputs(6));
    layer0_outputs(10475) <= (inputs(117)) xor (inputs(186));
    layer0_outputs(10476) <= (inputs(33)) and not (inputs(197));
    layer0_outputs(10477) <= inputs(131);
    layer0_outputs(10478) <= not(inputs(32)) or (inputs(201));
    layer0_outputs(10479) <= (inputs(248)) or (inputs(5));
    layer0_outputs(10480) <= (inputs(104)) xor (inputs(239));
    layer0_outputs(10481) <= not((inputs(152)) or (inputs(1)));
    layer0_outputs(10482) <= (inputs(49)) and (inputs(79));
    layer0_outputs(10483) <= not(inputs(147));
    layer0_outputs(10484) <= inputs(212);
    layer0_outputs(10485) <= inputs(68);
    layer0_outputs(10486) <= (inputs(5)) or (inputs(230));
    layer0_outputs(10487) <= '0';
    layer0_outputs(10488) <= (inputs(161)) xor (inputs(133));
    layer0_outputs(10489) <= not((inputs(174)) or (inputs(178)));
    layer0_outputs(10490) <= (inputs(215)) and (inputs(201));
    layer0_outputs(10491) <= (inputs(213)) and not (inputs(109));
    layer0_outputs(10492) <= inputs(89);
    layer0_outputs(10493) <= not(inputs(59));
    layer0_outputs(10494) <= not((inputs(44)) xor (inputs(57)));
    layer0_outputs(10495) <= not(inputs(198));
    layer0_outputs(10496) <= (inputs(215)) and not (inputs(52));
    layer0_outputs(10497) <= (inputs(75)) xor (inputs(37));
    layer0_outputs(10498) <= not(inputs(103));
    layer0_outputs(10499) <= (inputs(170)) xor (inputs(208));
    layer0_outputs(10500) <= not(inputs(100)) or (inputs(166));
    layer0_outputs(10501) <= not((inputs(147)) or (inputs(132)));
    layer0_outputs(10502) <= not((inputs(10)) xor (inputs(57)));
    layer0_outputs(10503) <= inputs(26);
    layer0_outputs(10504) <= inputs(127);
    layer0_outputs(10505) <= (inputs(153)) or (inputs(81));
    layer0_outputs(10506) <= not(inputs(202)) or (inputs(126));
    layer0_outputs(10507) <= not(inputs(19)) or (inputs(85));
    layer0_outputs(10508) <= not(inputs(63)) or (inputs(110));
    layer0_outputs(10509) <= inputs(164);
    layer0_outputs(10510) <= not((inputs(139)) xor (inputs(111)));
    layer0_outputs(10511) <= (inputs(224)) xor (inputs(105));
    layer0_outputs(10512) <= (inputs(196)) or (inputs(248));
    layer0_outputs(10513) <= (inputs(85)) and not (inputs(50));
    layer0_outputs(10514) <= (inputs(70)) xor (inputs(139));
    layer0_outputs(10515) <= (inputs(246)) and not (inputs(239));
    layer0_outputs(10516) <= not(inputs(229));
    layer0_outputs(10517) <= (inputs(197)) and not (inputs(70));
    layer0_outputs(10518) <= not(inputs(35)) or (inputs(113));
    layer0_outputs(10519) <= (inputs(181)) and (inputs(122));
    layer0_outputs(10520) <= not((inputs(128)) xor (inputs(11)));
    layer0_outputs(10521) <= inputs(70);
    layer0_outputs(10522) <= not((inputs(241)) or (inputs(255)));
    layer0_outputs(10523) <= not(inputs(75));
    layer0_outputs(10524) <= inputs(3);
    layer0_outputs(10525) <= not((inputs(93)) or (inputs(68)));
    layer0_outputs(10526) <= (inputs(220)) or (inputs(191));
    layer0_outputs(10527) <= not((inputs(4)) and (inputs(60)));
    layer0_outputs(10528) <= not((inputs(168)) and (inputs(232)));
    layer0_outputs(10529) <= (inputs(51)) and not (inputs(159));
    layer0_outputs(10530) <= inputs(81);
    layer0_outputs(10531) <= inputs(66);
    layer0_outputs(10532) <= not((inputs(78)) xor (inputs(173)));
    layer0_outputs(10533) <= inputs(30);
    layer0_outputs(10534) <= inputs(92);
    layer0_outputs(10535) <= not(inputs(218)) or (inputs(164));
    layer0_outputs(10536) <= not(inputs(35));
    layer0_outputs(10537) <= not(inputs(102)) or (inputs(126));
    layer0_outputs(10538) <= (inputs(23)) and (inputs(9));
    layer0_outputs(10539) <= not(inputs(65));
    layer0_outputs(10540) <= not((inputs(165)) xor (inputs(45)));
    layer0_outputs(10541) <= inputs(41);
    layer0_outputs(10542) <= not((inputs(162)) xor (inputs(179)));
    layer0_outputs(10543) <= (inputs(96)) or (inputs(191));
    layer0_outputs(10544) <= (inputs(68)) and not (inputs(119));
    layer0_outputs(10545) <= inputs(8);
    layer0_outputs(10546) <= not(inputs(97));
    layer0_outputs(10547) <= inputs(111);
    layer0_outputs(10548) <= inputs(181);
    layer0_outputs(10549) <= not(inputs(91));
    layer0_outputs(10550) <= inputs(84);
    layer0_outputs(10551) <= (inputs(26)) and not (inputs(220));
    layer0_outputs(10552) <= not(inputs(6)) or (inputs(106));
    layer0_outputs(10553) <= not((inputs(208)) xor (inputs(103)));
    layer0_outputs(10554) <= (inputs(45)) and not (inputs(7));
    layer0_outputs(10555) <= not((inputs(66)) xor (inputs(244)));
    layer0_outputs(10556) <= inputs(122);
    layer0_outputs(10557) <= inputs(43);
    layer0_outputs(10558) <= not(inputs(252));
    layer0_outputs(10559) <= (inputs(67)) xor (inputs(8));
    layer0_outputs(10560) <= inputs(190);
    layer0_outputs(10561) <= not((inputs(37)) xor (inputs(7)));
    layer0_outputs(10562) <= not(inputs(146));
    layer0_outputs(10563) <= not(inputs(219));
    layer0_outputs(10564) <= not((inputs(1)) or (inputs(56)));
    layer0_outputs(10565) <= inputs(35);
    layer0_outputs(10566) <= '0';
    layer0_outputs(10567) <= (inputs(22)) and not (inputs(130));
    layer0_outputs(10568) <= inputs(142);
    layer0_outputs(10569) <= not((inputs(213)) xor (inputs(176)));
    layer0_outputs(10570) <= (inputs(138)) or (inputs(174));
    layer0_outputs(10571) <= not(inputs(115));
    layer0_outputs(10572) <= not(inputs(59));
    layer0_outputs(10573) <= (inputs(179)) or (inputs(250));
    layer0_outputs(10574) <= (inputs(65)) xor (inputs(62));
    layer0_outputs(10575) <= (inputs(58)) and not (inputs(101));
    layer0_outputs(10576) <= not((inputs(89)) xor (inputs(207)));
    layer0_outputs(10577) <= not(inputs(27));
    layer0_outputs(10578) <= not((inputs(199)) or (inputs(206)));
    layer0_outputs(10579) <= inputs(76);
    layer0_outputs(10580) <= not((inputs(190)) xor (inputs(4)));
    layer0_outputs(10581) <= not((inputs(200)) xor (inputs(188)));
    layer0_outputs(10582) <= not(inputs(229));
    layer0_outputs(10583) <= not(inputs(70)) or (inputs(48));
    layer0_outputs(10584) <= (inputs(205)) xor (inputs(203));
    layer0_outputs(10585) <= not(inputs(102));
    layer0_outputs(10586) <= inputs(154);
    layer0_outputs(10587) <= inputs(21);
    layer0_outputs(10588) <= not(inputs(93));
    layer0_outputs(10589) <= inputs(87);
    layer0_outputs(10590) <= not((inputs(168)) xor (inputs(144)));
    layer0_outputs(10591) <= not((inputs(71)) xor (inputs(59)));
    layer0_outputs(10592) <= (inputs(49)) or (inputs(110));
    layer0_outputs(10593) <= not((inputs(43)) or (inputs(172)));
    layer0_outputs(10594) <= inputs(81);
    layer0_outputs(10595) <= (inputs(146)) and not (inputs(58));
    layer0_outputs(10596) <= not((inputs(133)) xor (inputs(87)));
    layer0_outputs(10597) <= (inputs(53)) and (inputs(54));
    layer0_outputs(10598) <= (inputs(94)) xor (inputs(107));
    layer0_outputs(10599) <= not(inputs(167)) or (inputs(242));
    layer0_outputs(10600) <= not(inputs(128));
    layer0_outputs(10601) <= not((inputs(19)) or (inputs(77)));
    layer0_outputs(10602) <= not(inputs(80));
    layer0_outputs(10603) <= (inputs(196)) xor (inputs(159));
    layer0_outputs(10604) <= not(inputs(135));
    layer0_outputs(10605) <= not((inputs(119)) xor (inputs(32)));
    layer0_outputs(10606) <= not((inputs(10)) xor (inputs(192)));
    layer0_outputs(10607) <= not(inputs(204));
    layer0_outputs(10608) <= not(inputs(54));
    layer0_outputs(10609) <= inputs(198);
    layer0_outputs(10610) <= (inputs(22)) and not (inputs(183));
    layer0_outputs(10611) <= (inputs(242)) or (inputs(137));
    layer0_outputs(10612) <= (inputs(80)) and not (inputs(12));
    layer0_outputs(10613) <= (inputs(173)) xor (inputs(255));
    layer0_outputs(10614) <= not(inputs(146));
    layer0_outputs(10615) <= not(inputs(214));
    layer0_outputs(10616) <= not(inputs(68)) or (inputs(48));
    layer0_outputs(10617) <= (inputs(155)) and not (inputs(135));
    layer0_outputs(10618) <= (inputs(182)) and (inputs(155));
    layer0_outputs(10619) <= (inputs(60)) xor (inputs(150));
    layer0_outputs(10620) <= (inputs(254)) or (inputs(110));
    layer0_outputs(10621) <= not(inputs(23));
    layer0_outputs(10622) <= (inputs(33)) or (inputs(195));
    layer0_outputs(10623) <= not(inputs(231)) or (inputs(105));
    layer0_outputs(10624) <= not(inputs(147)) or (inputs(190));
    layer0_outputs(10625) <= not(inputs(105));
    layer0_outputs(10626) <= (inputs(113)) or (inputs(53));
    layer0_outputs(10627) <= not((inputs(54)) xor (inputs(184)));
    layer0_outputs(10628) <= (inputs(62)) or (inputs(19));
    layer0_outputs(10629) <= (inputs(135)) and not (inputs(34));
    layer0_outputs(10630) <= (inputs(208)) and not (inputs(143));
    layer0_outputs(10631) <= not((inputs(165)) or (inputs(141)));
    layer0_outputs(10632) <= not(inputs(135));
    layer0_outputs(10633) <= not(inputs(205));
    layer0_outputs(10634) <= (inputs(58)) or (inputs(107));
    layer0_outputs(10635) <= (inputs(125)) or (inputs(232));
    layer0_outputs(10636) <= (inputs(149)) and (inputs(106));
    layer0_outputs(10637) <= inputs(184);
    layer0_outputs(10638) <= not(inputs(141));
    layer0_outputs(10639) <= inputs(208);
    layer0_outputs(10640) <= (inputs(114)) and not (inputs(251));
    layer0_outputs(10641) <= inputs(89);
    layer0_outputs(10642) <= not((inputs(129)) xor (inputs(139)));
    layer0_outputs(10643) <= not(inputs(6)) or (inputs(57));
    layer0_outputs(10644) <= inputs(197);
    layer0_outputs(10645) <= not(inputs(194));
    layer0_outputs(10646) <= not((inputs(64)) xor (inputs(228)));
    layer0_outputs(10647) <= not((inputs(192)) or (inputs(244)));
    layer0_outputs(10648) <= not((inputs(237)) or (inputs(110)));
    layer0_outputs(10649) <= (inputs(244)) xor (inputs(153));
    layer0_outputs(10650) <= (inputs(122)) and (inputs(119));
    layer0_outputs(10651) <= inputs(166);
    layer0_outputs(10652) <= not(inputs(226)) or (inputs(149));
    layer0_outputs(10653) <= inputs(130);
    layer0_outputs(10654) <= not((inputs(80)) xor (inputs(48)));
    layer0_outputs(10655) <= not((inputs(155)) xor (inputs(131)));
    layer0_outputs(10656) <= (inputs(159)) xor (inputs(23));
    layer0_outputs(10657) <= (inputs(111)) and (inputs(49));
    layer0_outputs(10658) <= (inputs(0)) xor (inputs(6));
    layer0_outputs(10659) <= not(inputs(93)) or (inputs(236));
    layer0_outputs(10660) <= not((inputs(195)) or (inputs(175)));
    layer0_outputs(10661) <= '0';
    layer0_outputs(10662) <= (inputs(13)) and not (inputs(39));
    layer0_outputs(10663) <= inputs(199);
    layer0_outputs(10664) <= (inputs(78)) xor (inputs(195));
    layer0_outputs(10665) <= not((inputs(27)) xor (inputs(28)));
    layer0_outputs(10666) <= (inputs(70)) and not (inputs(190));
    layer0_outputs(10667) <= not((inputs(227)) xor (inputs(207)));
    layer0_outputs(10668) <= not((inputs(30)) xor (inputs(109)));
    layer0_outputs(10669) <= inputs(128);
    layer0_outputs(10670) <= not((inputs(103)) and (inputs(167)));
    layer0_outputs(10671) <= (inputs(159)) and not (inputs(11));
    layer0_outputs(10672) <= not(inputs(105));
    layer0_outputs(10673) <= (inputs(129)) xor (inputs(85));
    layer0_outputs(10674) <= not(inputs(123));
    layer0_outputs(10675) <= not(inputs(25));
    layer0_outputs(10676) <= not(inputs(106));
    layer0_outputs(10677) <= not((inputs(0)) or (inputs(54)));
    layer0_outputs(10678) <= (inputs(7)) or (inputs(18));
    layer0_outputs(10679) <= not(inputs(103));
    layer0_outputs(10680) <= not(inputs(24)) or (inputs(181));
    layer0_outputs(10681) <= inputs(195);
    layer0_outputs(10682) <= (inputs(79)) xor (inputs(82));
    layer0_outputs(10683) <= (inputs(175)) xor (inputs(110));
    layer0_outputs(10684) <= not(inputs(209));
    layer0_outputs(10685) <= not(inputs(162));
    layer0_outputs(10686) <= not(inputs(57)) or (inputs(174));
    layer0_outputs(10687) <= inputs(41);
    layer0_outputs(10688) <= not(inputs(138)) or (inputs(179));
    layer0_outputs(10689) <= not(inputs(176));
    layer0_outputs(10690) <= not(inputs(100));
    layer0_outputs(10691) <= (inputs(99)) or (inputs(172));
    layer0_outputs(10692) <= not(inputs(17));
    layer0_outputs(10693) <= not((inputs(91)) xor (inputs(125)));
    layer0_outputs(10694) <= inputs(197);
    layer0_outputs(10695) <= inputs(116);
    layer0_outputs(10696) <= not((inputs(137)) or (inputs(20)));
    layer0_outputs(10697) <= not(inputs(173)) or (inputs(31));
    layer0_outputs(10698) <= not((inputs(112)) or (inputs(25)));
    layer0_outputs(10699) <= inputs(55);
    layer0_outputs(10700) <= not((inputs(64)) and (inputs(140)));
    layer0_outputs(10701) <= not((inputs(237)) or (inputs(14)));
    layer0_outputs(10702) <= not((inputs(175)) xor (inputs(18)));
    layer0_outputs(10703) <= inputs(9);
    layer0_outputs(10704) <= (inputs(188)) xor (inputs(107));
    layer0_outputs(10705) <= not(inputs(7));
    layer0_outputs(10706) <= inputs(226);
    layer0_outputs(10707) <= inputs(233);
    layer0_outputs(10708) <= not(inputs(124)) or (inputs(151));
    layer0_outputs(10709) <= '0';
    layer0_outputs(10710) <= (inputs(189)) or (inputs(159));
    layer0_outputs(10711) <= not(inputs(148)) or (inputs(17));
    layer0_outputs(10712) <= not(inputs(57));
    layer0_outputs(10713) <= not(inputs(233));
    layer0_outputs(10714) <= inputs(127);
    layer0_outputs(10715) <= (inputs(144)) or (inputs(178));
    layer0_outputs(10716) <= (inputs(106)) and not (inputs(127));
    layer0_outputs(10717) <= (inputs(17)) xor (inputs(134));
    layer0_outputs(10718) <= inputs(137);
    layer0_outputs(10719) <= not((inputs(200)) xor (inputs(214)));
    layer0_outputs(10720) <= (inputs(121)) xor (inputs(132));
    layer0_outputs(10721) <= inputs(172);
    layer0_outputs(10722) <= not((inputs(210)) or (inputs(3)));
    layer0_outputs(10723) <= (inputs(208)) and not (inputs(241));
    layer0_outputs(10724) <= inputs(25);
    layer0_outputs(10725) <= not((inputs(204)) xor (inputs(11)));
    layer0_outputs(10726) <= (inputs(49)) and not (inputs(175));
    layer0_outputs(10727) <= not(inputs(51));
    layer0_outputs(10728) <= not((inputs(134)) and (inputs(39)));
    layer0_outputs(10729) <= not(inputs(40));
    layer0_outputs(10730) <= not(inputs(51));
    layer0_outputs(10731) <= not(inputs(153));
    layer0_outputs(10732) <= (inputs(7)) or (inputs(96));
    layer0_outputs(10733) <= not((inputs(134)) and (inputs(144)));
    layer0_outputs(10734) <= (inputs(173)) and not (inputs(134));
    layer0_outputs(10735) <= inputs(230);
    layer0_outputs(10736) <= (inputs(195)) xor (inputs(240));
    layer0_outputs(10737) <= inputs(91);
    layer0_outputs(10738) <= (inputs(13)) and not (inputs(254));
    layer0_outputs(10739) <= inputs(233);
    layer0_outputs(10740) <= (inputs(126)) or (inputs(231));
    layer0_outputs(10741) <= not((inputs(52)) and (inputs(29)));
    layer0_outputs(10742) <= not(inputs(24));
    layer0_outputs(10743) <= not(inputs(8)) or (inputs(131));
    layer0_outputs(10744) <= not(inputs(124));
    layer0_outputs(10745) <= not(inputs(59));
    layer0_outputs(10746) <= not(inputs(107));
    layer0_outputs(10747) <= not(inputs(89)) or (inputs(176));
    layer0_outputs(10748) <= not(inputs(146));
    layer0_outputs(10749) <= (inputs(25)) xor (inputs(72));
    layer0_outputs(10750) <= not(inputs(10));
    layer0_outputs(10751) <= inputs(161);
    layer0_outputs(10752) <= not(inputs(10));
    layer0_outputs(10753) <= not(inputs(8));
    layer0_outputs(10754) <= not(inputs(153));
    layer0_outputs(10755) <= inputs(101);
    layer0_outputs(10756) <= not((inputs(41)) xor (inputs(80)));
    layer0_outputs(10757) <= not((inputs(93)) xor (inputs(175)));
    layer0_outputs(10758) <= (inputs(140)) and not (inputs(88));
    layer0_outputs(10759) <= (inputs(28)) xor (inputs(37));
    layer0_outputs(10760) <= not((inputs(217)) or (inputs(226)));
    layer0_outputs(10761) <= inputs(29);
    layer0_outputs(10762) <= (inputs(115)) xor (inputs(117));
    layer0_outputs(10763) <= (inputs(174)) xor (inputs(241));
    layer0_outputs(10764) <= (inputs(190)) and not (inputs(78));
    layer0_outputs(10765) <= (inputs(197)) and not (inputs(120));
    layer0_outputs(10766) <= (inputs(64)) and not (inputs(151));
    layer0_outputs(10767) <= (inputs(157)) and not (inputs(65));
    layer0_outputs(10768) <= not(inputs(72)) or (inputs(209));
    layer0_outputs(10769) <= not(inputs(27));
    layer0_outputs(10770) <= (inputs(122)) xor (inputs(141));
    layer0_outputs(10771) <= not(inputs(96));
    layer0_outputs(10772) <= not(inputs(44)) or (inputs(97));
    layer0_outputs(10773) <= not(inputs(147));
    layer0_outputs(10774) <= (inputs(232)) and not (inputs(24));
    layer0_outputs(10775) <= (inputs(24)) xor (inputs(1));
    layer0_outputs(10776) <= inputs(219);
    layer0_outputs(10777) <= inputs(198);
    layer0_outputs(10778) <= not(inputs(214));
    layer0_outputs(10779) <= (inputs(138)) or (inputs(176));
    layer0_outputs(10780) <= not(inputs(133));
    layer0_outputs(10781) <= (inputs(175)) or (inputs(187));
    layer0_outputs(10782) <= not(inputs(99)) or (inputs(168));
    layer0_outputs(10783) <= inputs(129);
    layer0_outputs(10784) <= (inputs(133)) xor (inputs(178));
    layer0_outputs(10785) <= (inputs(116)) and not (inputs(251));
    layer0_outputs(10786) <= not(inputs(212));
    layer0_outputs(10787) <= not(inputs(24));
    layer0_outputs(10788) <= (inputs(97)) xor (inputs(85));
    layer0_outputs(10789) <= not(inputs(180)) or (inputs(221));
    layer0_outputs(10790) <= not((inputs(165)) xor (inputs(167)));
    layer0_outputs(10791) <= inputs(144);
    layer0_outputs(10792) <= (inputs(87)) and not (inputs(94));
    layer0_outputs(10793) <= not((inputs(84)) xor (inputs(34)));
    layer0_outputs(10794) <= not(inputs(123)) or (inputs(199));
    layer0_outputs(10795) <= not((inputs(221)) or (inputs(157)));
    layer0_outputs(10796) <= not(inputs(90)) or (inputs(173));
    layer0_outputs(10797) <= (inputs(154)) and not (inputs(97));
    layer0_outputs(10798) <= not(inputs(30));
    layer0_outputs(10799) <= not(inputs(5)) or (inputs(255));
    layer0_outputs(10800) <= '0';
    layer0_outputs(10801) <= not(inputs(145));
    layer0_outputs(10802) <= inputs(82);
    layer0_outputs(10803) <= not((inputs(65)) or (inputs(71)));
    layer0_outputs(10804) <= inputs(85);
    layer0_outputs(10805) <= not((inputs(30)) or (inputs(73)));
    layer0_outputs(10806) <= inputs(230);
    layer0_outputs(10807) <= inputs(140);
    layer0_outputs(10808) <= (inputs(208)) or (inputs(62));
    layer0_outputs(10809) <= not(inputs(99)) or (inputs(80));
    layer0_outputs(10810) <= not(inputs(130));
    layer0_outputs(10811) <= not(inputs(243));
    layer0_outputs(10812) <= (inputs(84)) and not (inputs(38));
    layer0_outputs(10813) <= not(inputs(231));
    layer0_outputs(10814) <= not(inputs(0)) or (inputs(123));
    layer0_outputs(10815) <= not(inputs(185)) or (inputs(3));
    layer0_outputs(10816) <= not((inputs(203)) or (inputs(36)));
    layer0_outputs(10817) <= inputs(22);
    layer0_outputs(10818) <= not(inputs(195)) or (inputs(20));
    layer0_outputs(10819) <= not(inputs(42)) or (inputs(206));
    layer0_outputs(10820) <= (inputs(222)) or (inputs(123));
    layer0_outputs(10821) <= not(inputs(165));
    layer0_outputs(10822) <= inputs(30);
    layer0_outputs(10823) <= inputs(65);
    layer0_outputs(10824) <= not((inputs(115)) or (inputs(252)));
    layer0_outputs(10825) <= (inputs(214)) and not (inputs(4));
    layer0_outputs(10826) <= inputs(96);
    layer0_outputs(10827) <= (inputs(92)) xor (inputs(31));
    layer0_outputs(10828) <= not((inputs(54)) xor (inputs(27)));
    layer0_outputs(10829) <= not(inputs(194)) or (inputs(64));
    layer0_outputs(10830) <= not(inputs(93)) or (inputs(253));
    layer0_outputs(10831) <= inputs(63);
    layer0_outputs(10832) <= not((inputs(73)) or (inputs(113)));
    layer0_outputs(10833) <= '0';
    layer0_outputs(10834) <= not(inputs(82));
    layer0_outputs(10835) <= (inputs(126)) or (inputs(34));
    layer0_outputs(10836) <= inputs(150);
    layer0_outputs(10837) <= not(inputs(230));
    layer0_outputs(10838) <= not((inputs(180)) and (inputs(202)));
    layer0_outputs(10839) <= (inputs(61)) or (inputs(176));
    layer0_outputs(10840) <= inputs(64);
    layer0_outputs(10841) <= inputs(56);
    layer0_outputs(10842) <= (inputs(181)) and not (inputs(172));
    layer0_outputs(10843) <= (inputs(41)) xor (inputs(14));
    layer0_outputs(10844) <= (inputs(214)) or (inputs(0));
    layer0_outputs(10845) <= not(inputs(164));
    layer0_outputs(10846) <= (inputs(73)) and not (inputs(176));
    layer0_outputs(10847) <= not(inputs(86)) or (inputs(193));
    layer0_outputs(10848) <= not(inputs(114));
    layer0_outputs(10849) <= not((inputs(16)) or (inputs(132)));
    layer0_outputs(10850) <= not(inputs(42)) or (inputs(0));
    layer0_outputs(10851) <= inputs(202);
    layer0_outputs(10852) <= (inputs(132)) and (inputs(67));
    layer0_outputs(10853) <= (inputs(216)) and not (inputs(48));
    layer0_outputs(10854) <= not((inputs(198)) or (inputs(209)));
    layer0_outputs(10855) <= not(inputs(45)) or (inputs(169));
    layer0_outputs(10856) <= inputs(104);
    layer0_outputs(10857) <= not((inputs(255)) or (inputs(236)));
    layer0_outputs(10858) <= not((inputs(107)) xor (inputs(210)));
    layer0_outputs(10859) <= inputs(254);
    layer0_outputs(10860) <= not(inputs(172)) or (inputs(85));
    layer0_outputs(10861) <= not(inputs(28));
    layer0_outputs(10862) <= inputs(19);
    layer0_outputs(10863) <= not((inputs(151)) xor (inputs(93)));
    layer0_outputs(10864) <= not((inputs(125)) xor (inputs(176)));
    layer0_outputs(10865) <= not((inputs(255)) xor (inputs(199)));
    layer0_outputs(10866) <= inputs(62);
    layer0_outputs(10867) <= not(inputs(125));
    layer0_outputs(10868) <= not(inputs(180)) or (inputs(62));
    layer0_outputs(10869) <= (inputs(88)) xor (inputs(76));
    layer0_outputs(10870) <= (inputs(194)) or (inputs(89));
    layer0_outputs(10871) <= (inputs(217)) and not (inputs(150));
    layer0_outputs(10872) <= inputs(229);
    layer0_outputs(10873) <= not((inputs(147)) or (inputs(65)));
    layer0_outputs(10874) <= not((inputs(24)) or (inputs(48)));
    layer0_outputs(10875) <= not(inputs(181));
    layer0_outputs(10876) <= (inputs(243)) or (inputs(46));
    layer0_outputs(10877) <= (inputs(226)) xor (inputs(163));
    layer0_outputs(10878) <= not(inputs(208)) or (inputs(185));
    layer0_outputs(10879) <= (inputs(117)) and not (inputs(96));
    layer0_outputs(10880) <= not(inputs(201)) or (inputs(120));
    layer0_outputs(10881) <= not(inputs(203));
    layer0_outputs(10882) <= (inputs(6)) and not (inputs(195));
    layer0_outputs(10883) <= inputs(83);
    layer0_outputs(10884) <= (inputs(191)) and not (inputs(65));
    layer0_outputs(10885) <= not(inputs(86));
    layer0_outputs(10886) <= not(inputs(81));
    layer0_outputs(10887) <= not((inputs(89)) xor (inputs(64)));
    layer0_outputs(10888) <= (inputs(163)) and not (inputs(11));
    layer0_outputs(10889) <= inputs(119);
    layer0_outputs(10890) <= inputs(222);
    layer0_outputs(10891) <= not((inputs(116)) xor (inputs(117)));
    layer0_outputs(10892) <= not((inputs(108)) xor (inputs(106)));
    layer0_outputs(10893) <= (inputs(162)) xor (inputs(90));
    layer0_outputs(10894) <= not((inputs(174)) xor (inputs(107)));
    layer0_outputs(10895) <= (inputs(51)) or (inputs(128));
    layer0_outputs(10896) <= not((inputs(164)) xor (inputs(36)));
    layer0_outputs(10897) <= (inputs(37)) or (inputs(158));
    layer0_outputs(10898) <= (inputs(229)) and (inputs(85));
    layer0_outputs(10899) <= inputs(38);
    layer0_outputs(10900) <= inputs(137);
    layer0_outputs(10901) <= not((inputs(48)) xor (inputs(98)));
    layer0_outputs(10902) <= not(inputs(34)) or (inputs(84));
    layer0_outputs(10903) <= not((inputs(180)) or (inputs(26)));
    layer0_outputs(10904) <= inputs(209);
    layer0_outputs(10905) <= inputs(122);
    layer0_outputs(10906) <= (inputs(55)) or (inputs(251));
    layer0_outputs(10907) <= not((inputs(13)) or (inputs(239)));
    layer0_outputs(10908) <= (inputs(121)) or (inputs(182));
    layer0_outputs(10909) <= not(inputs(112)) or (inputs(67));
    layer0_outputs(10910) <= (inputs(247)) or (inputs(93));
    layer0_outputs(10911) <= not((inputs(214)) xor (inputs(223)));
    layer0_outputs(10912) <= (inputs(80)) or (inputs(105));
    layer0_outputs(10913) <= '0';
    layer0_outputs(10914) <= (inputs(207)) and not (inputs(63));
    layer0_outputs(10915) <= (inputs(25)) xor (inputs(35));
    layer0_outputs(10916) <= not(inputs(218));
    layer0_outputs(10917) <= inputs(183);
    layer0_outputs(10918) <= not(inputs(27)) or (inputs(185));
    layer0_outputs(10919) <= not((inputs(176)) xor (inputs(80)));
    layer0_outputs(10920) <= (inputs(193)) and not (inputs(44));
    layer0_outputs(10921) <= (inputs(9)) and not (inputs(235));
    layer0_outputs(10922) <= not(inputs(41)) or (inputs(222));
    layer0_outputs(10923) <= (inputs(105)) and not (inputs(204));
    layer0_outputs(10924) <= not(inputs(136));
    layer0_outputs(10925) <= (inputs(203)) or (inputs(34));
    layer0_outputs(10926) <= not((inputs(42)) xor (inputs(55)));
    layer0_outputs(10927) <= not(inputs(43));
    layer0_outputs(10928) <= not((inputs(219)) xor (inputs(252)));
    layer0_outputs(10929) <= not(inputs(71)) or (inputs(50));
    layer0_outputs(10930) <= not((inputs(81)) xor (inputs(121)));
    layer0_outputs(10931) <= inputs(149);
    layer0_outputs(10932) <= (inputs(201)) and not (inputs(236));
    layer0_outputs(10933) <= not(inputs(49)) or (inputs(150));
    layer0_outputs(10934) <= (inputs(172)) xor (inputs(109));
    layer0_outputs(10935) <= not((inputs(95)) or (inputs(48)));
    layer0_outputs(10936) <= (inputs(204)) and not (inputs(35));
    layer0_outputs(10937) <= not(inputs(210));
    layer0_outputs(10938) <= not((inputs(71)) xor (inputs(218)));
    layer0_outputs(10939) <= not((inputs(73)) or (inputs(142)));
    layer0_outputs(10940) <= not((inputs(70)) and (inputs(218)));
    layer0_outputs(10941) <= (inputs(197)) and not (inputs(140));
    layer0_outputs(10942) <= inputs(56);
    layer0_outputs(10943) <= not((inputs(127)) and (inputs(127)));
    layer0_outputs(10944) <= not(inputs(176)) or (inputs(48));
    layer0_outputs(10945) <= (inputs(164)) xor (inputs(237));
    layer0_outputs(10946) <= not(inputs(13)) or (inputs(192));
    layer0_outputs(10947) <= (inputs(152)) and not (inputs(50));
    layer0_outputs(10948) <= '0';
    layer0_outputs(10949) <= not(inputs(193));
    layer0_outputs(10950) <= not(inputs(172));
    layer0_outputs(10951) <= '0';
    layer0_outputs(10952) <= (inputs(135)) and not (inputs(86));
    layer0_outputs(10953) <= (inputs(99)) and (inputs(187));
    layer0_outputs(10954) <= inputs(57);
    layer0_outputs(10955) <= (inputs(209)) and not (inputs(115));
    layer0_outputs(10956) <= (inputs(141)) or (inputs(112));
    layer0_outputs(10957) <= not(inputs(39));
    layer0_outputs(10958) <= (inputs(235)) xor (inputs(154));
    layer0_outputs(10959) <= not(inputs(167)) or (inputs(101));
    layer0_outputs(10960) <= not((inputs(214)) or (inputs(163)));
    layer0_outputs(10961) <= (inputs(210)) and not (inputs(76));
    layer0_outputs(10962) <= inputs(99);
    layer0_outputs(10963) <= inputs(11);
    layer0_outputs(10964) <= (inputs(122)) xor (inputs(58));
    layer0_outputs(10965) <= not((inputs(81)) xor (inputs(19)));
    layer0_outputs(10966) <= inputs(174);
    layer0_outputs(10967) <= (inputs(117)) xor (inputs(138));
    layer0_outputs(10968) <= inputs(215);
    layer0_outputs(10969) <= not(inputs(97));
    layer0_outputs(10970) <= not((inputs(19)) xor (inputs(136)));
    layer0_outputs(10971) <= (inputs(111)) and not (inputs(144));
    layer0_outputs(10972) <= not((inputs(224)) xor (inputs(189)));
    layer0_outputs(10973) <= (inputs(50)) xor (inputs(34));
    layer0_outputs(10974) <= inputs(151);
    layer0_outputs(10975) <= not(inputs(5)) or (inputs(1));
    layer0_outputs(10976) <= inputs(127);
    layer0_outputs(10977) <= not(inputs(250));
    layer0_outputs(10978) <= (inputs(202)) or (inputs(128));
    layer0_outputs(10979) <= not((inputs(178)) or (inputs(4)));
    layer0_outputs(10980) <= inputs(92);
    layer0_outputs(10981) <= (inputs(91)) or (inputs(66));
    layer0_outputs(10982) <= (inputs(135)) and (inputs(125));
    layer0_outputs(10983) <= not((inputs(85)) or (inputs(37)));
    layer0_outputs(10984) <= not(inputs(98)) or (inputs(15));
    layer0_outputs(10985) <= (inputs(252)) or (inputs(193));
    layer0_outputs(10986) <= not(inputs(152)) or (inputs(81));
    layer0_outputs(10987) <= not(inputs(31));
    layer0_outputs(10988) <= inputs(140);
    layer0_outputs(10989) <= not((inputs(179)) or (inputs(188)));
    layer0_outputs(10990) <= inputs(232);
    layer0_outputs(10991) <= not(inputs(117)) or (inputs(244));
    layer0_outputs(10992) <= inputs(164);
    layer0_outputs(10993) <= inputs(170);
    layer0_outputs(10994) <= (inputs(244)) or (inputs(191));
    layer0_outputs(10995) <= (inputs(196)) and not (inputs(30));
    layer0_outputs(10996) <= not((inputs(46)) xor (inputs(12)));
    layer0_outputs(10997) <= (inputs(211)) and not (inputs(113));
    layer0_outputs(10998) <= (inputs(63)) and not (inputs(240));
    layer0_outputs(10999) <= not(inputs(232));
    layer0_outputs(11000) <= (inputs(30)) or (inputs(120));
    layer0_outputs(11001) <= (inputs(21)) and not (inputs(37));
    layer0_outputs(11002) <= not((inputs(229)) xor (inputs(95)));
    layer0_outputs(11003) <= inputs(253);
    layer0_outputs(11004) <= not(inputs(110));
    layer0_outputs(11005) <= '0';
    layer0_outputs(11006) <= inputs(137);
    layer0_outputs(11007) <= not(inputs(127));
    layer0_outputs(11008) <= inputs(5);
    layer0_outputs(11009) <= inputs(71);
    layer0_outputs(11010) <= (inputs(40)) xor (inputs(177));
    layer0_outputs(11011) <= (inputs(28)) and not (inputs(132));
    layer0_outputs(11012) <= not(inputs(198)) or (inputs(114));
    layer0_outputs(11013) <= not((inputs(225)) or (inputs(181)));
    layer0_outputs(11014) <= inputs(98);
    layer0_outputs(11015) <= (inputs(31)) xor (inputs(67));
    layer0_outputs(11016) <= not((inputs(229)) and (inputs(131)));
    layer0_outputs(11017) <= (inputs(232)) and not (inputs(5));
    layer0_outputs(11018) <= not((inputs(223)) and (inputs(57)));
    layer0_outputs(11019) <= inputs(189);
    layer0_outputs(11020) <= not(inputs(222)) or (inputs(13));
    layer0_outputs(11021) <= (inputs(73)) and not (inputs(28));
    layer0_outputs(11022) <= '1';
    layer0_outputs(11023) <= (inputs(72)) and not (inputs(67));
    layer0_outputs(11024) <= not((inputs(41)) or (inputs(31)));
    layer0_outputs(11025) <= (inputs(112)) and not (inputs(48));
    layer0_outputs(11026) <= not(inputs(209)) or (inputs(252));
    layer0_outputs(11027) <= not(inputs(130)) or (inputs(15));
    layer0_outputs(11028) <= not((inputs(227)) xor (inputs(181)));
    layer0_outputs(11029) <= (inputs(43)) xor (inputs(90));
    layer0_outputs(11030) <= not(inputs(98));
    layer0_outputs(11031) <= (inputs(146)) xor (inputs(116));
    layer0_outputs(11032) <= not((inputs(184)) and (inputs(64)));
    layer0_outputs(11033) <= not(inputs(14));
    layer0_outputs(11034) <= (inputs(104)) and (inputs(214));
    layer0_outputs(11035) <= not((inputs(21)) xor (inputs(54)));
    layer0_outputs(11036) <= inputs(113);
    layer0_outputs(11037) <= (inputs(104)) or (inputs(206));
    layer0_outputs(11038) <= not((inputs(166)) xor (inputs(234)));
    layer0_outputs(11039) <= not((inputs(85)) xor (inputs(58)));
    layer0_outputs(11040) <= (inputs(107)) or (inputs(60));
    layer0_outputs(11041) <= (inputs(215)) or (inputs(190));
    layer0_outputs(11042) <= (inputs(225)) or (inputs(253));
    layer0_outputs(11043) <= (inputs(58)) xor (inputs(192));
    layer0_outputs(11044) <= (inputs(32)) or (inputs(121));
    layer0_outputs(11045) <= not(inputs(182));
    layer0_outputs(11046) <= not(inputs(83)) or (inputs(60));
    layer0_outputs(11047) <= (inputs(69)) xor (inputs(82));
    layer0_outputs(11048) <= not(inputs(110));
    layer0_outputs(11049) <= (inputs(60)) and (inputs(27));
    layer0_outputs(11050) <= not((inputs(81)) xor (inputs(86)));
    layer0_outputs(11051) <= inputs(218);
    layer0_outputs(11052) <= not((inputs(104)) xor (inputs(124)));
    layer0_outputs(11053) <= (inputs(156)) or (inputs(12));
    layer0_outputs(11054) <= (inputs(41)) and not (inputs(112));
    layer0_outputs(11055) <= not(inputs(13));
    layer0_outputs(11056) <= (inputs(104)) or (inputs(219));
    layer0_outputs(11057) <= not((inputs(190)) or (inputs(81)));
    layer0_outputs(11058) <= not(inputs(213));
    layer0_outputs(11059) <= not((inputs(19)) and (inputs(34)));
    layer0_outputs(11060) <= not(inputs(169));
    layer0_outputs(11061) <= (inputs(210)) xor (inputs(194));
    layer0_outputs(11062) <= inputs(147);
    layer0_outputs(11063) <= not((inputs(186)) xor (inputs(155)));
    layer0_outputs(11064) <= not(inputs(130)) or (inputs(191));
    layer0_outputs(11065) <= inputs(71);
    layer0_outputs(11066) <= not(inputs(236)) or (inputs(127));
    layer0_outputs(11067) <= not((inputs(171)) xor (inputs(185)));
    layer0_outputs(11068) <= not(inputs(33)) or (inputs(232));
    layer0_outputs(11069) <= not(inputs(12));
    layer0_outputs(11070) <= inputs(169);
    layer0_outputs(11071) <= not((inputs(239)) or (inputs(76)));
    layer0_outputs(11072) <= inputs(191);
    layer0_outputs(11073) <= not(inputs(7));
    layer0_outputs(11074) <= (inputs(228)) or (inputs(247));
    layer0_outputs(11075) <= inputs(107);
    layer0_outputs(11076) <= not((inputs(203)) xor (inputs(232)));
    layer0_outputs(11077) <= not(inputs(123));
    layer0_outputs(11078) <= not(inputs(146));
    layer0_outputs(11079) <= inputs(60);
    layer0_outputs(11080) <= (inputs(51)) and not (inputs(210));
    layer0_outputs(11081) <= not((inputs(61)) and (inputs(76)));
    layer0_outputs(11082) <= (inputs(28)) or (inputs(71));
    layer0_outputs(11083) <= not(inputs(57));
    layer0_outputs(11084) <= not((inputs(175)) or (inputs(40)));
    layer0_outputs(11085) <= not(inputs(38));
    layer0_outputs(11086) <= inputs(100);
    layer0_outputs(11087) <= not(inputs(163)) or (inputs(74));
    layer0_outputs(11088) <= not(inputs(210));
    layer0_outputs(11089) <= (inputs(167)) xor (inputs(164));
    layer0_outputs(11090) <= (inputs(114)) or (inputs(117));
    layer0_outputs(11091) <= not(inputs(225)) or (inputs(47));
    layer0_outputs(11092) <= not(inputs(150));
    layer0_outputs(11093) <= (inputs(53)) or (inputs(119));
    layer0_outputs(11094) <= inputs(231);
    layer0_outputs(11095) <= inputs(185);
    layer0_outputs(11096) <= inputs(10);
    layer0_outputs(11097) <= (inputs(98)) or (inputs(161));
    layer0_outputs(11098) <= (inputs(227)) and not (inputs(19));
    layer0_outputs(11099) <= not((inputs(12)) xor (inputs(59)));
    layer0_outputs(11100) <= inputs(152);
    layer0_outputs(11101) <= (inputs(204)) xor (inputs(46));
    layer0_outputs(11102) <= not(inputs(101));
    layer0_outputs(11103) <= not((inputs(16)) xor (inputs(216)));
    layer0_outputs(11104) <= '0';
    layer0_outputs(11105) <= not(inputs(108)) or (inputs(175));
    layer0_outputs(11106) <= (inputs(124)) and not (inputs(223));
    layer0_outputs(11107) <= not(inputs(216));
    layer0_outputs(11108) <= (inputs(100)) xor (inputs(160));
    layer0_outputs(11109) <= not((inputs(210)) or (inputs(214)));
    layer0_outputs(11110) <= not(inputs(54));
    layer0_outputs(11111) <= not((inputs(241)) xor (inputs(32)));
    layer0_outputs(11112) <= (inputs(34)) xor (inputs(237));
    layer0_outputs(11113) <= (inputs(229)) and not (inputs(52));
    layer0_outputs(11114) <= inputs(91);
    layer0_outputs(11115) <= inputs(52);
    layer0_outputs(11116) <= not((inputs(166)) or (inputs(253)));
    layer0_outputs(11117) <= (inputs(233)) and not (inputs(20));
    layer0_outputs(11118) <= (inputs(51)) or (inputs(191));
    layer0_outputs(11119) <= (inputs(46)) xor (inputs(42));
    layer0_outputs(11120) <= not(inputs(12)) or (inputs(153));
    layer0_outputs(11121) <= (inputs(68)) and not (inputs(209));
    layer0_outputs(11122) <= (inputs(21)) or (inputs(45));
    layer0_outputs(11123) <= not(inputs(83)) or (inputs(1));
    layer0_outputs(11124) <= inputs(5);
    layer0_outputs(11125) <= inputs(18);
    layer0_outputs(11126) <= not((inputs(73)) and (inputs(110)));
    layer0_outputs(11127) <= not(inputs(214));
    layer0_outputs(11128) <= (inputs(143)) or (inputs(81));
    layer0_outputs(11129) <= not(inputs(7)) or (inputs(163));
    layer0_outputs(11130) <= not(inputs(6));
    layer0_outputs(11131) <= (inputs(141)) or (inputs(226));
    layer0_outputs(11132) <= (inputs(162)) or (inputs(125));
    layer0_outputs(11133) <= not((inputs(20)) or (inputs(221)));
    layer0_outputs(11134) <= (inputs(84)) and not (inputs(194));
    layer0_outputs(11135) <= not(inputs(195));
    layer0_outputs(11136) <= (inputs(138)) xor (inputs(186));
    layer0_outputs(11137) <= not((inputs(35)) xor (inputs(11)));
    layer0_outputs(11138) <= not(inputs(100));
    layer0_outputs(11139) <= not(inputs(25));
    layer0_outputs(11140) <= not(inputs(62)) or (inputs(251));
    layer0_outputs(11141) <= not(inputs(44)) or (inputs(16));
    layer0_outputs(11142) <= not(inputs(44)) or (inputs(144));
    layer0_outputs(11143) <= inputs(230);
    layer0_outputs(11144) <= (inputs(4)) and not (inputs(241));
    layer0_outputs(11145) <= (inputs(172)) and not (inputs(3));
    layer0_outputs(11146) <= (inputs(225)) and not (inputs(113));
    layer0_outputs(11147) <= '0';
    layer0_outputs(11148) <= not((inputs(192)) or (inputs(243)));
    layer0_outputs(11149) <= not(inputs(245));
    layer0_outputs(11150) <= (inputs(198)) and not (inputs(94));
    layer0_outputs(11151) <= inputs(239);
    layer0_outputs(11152) <= not(inputs(147));
    layer0_outputs(11153) <= (inputs(48)) or (inputs(200));
    layer0_outputs(11154) <= (inputs(176)) or (inputs(161));
    layer0_outputs(11155) <= inputs(235);
    layer0_outputs(11156) <= not(inputs(227)) or (inputs(47));
    layer0_outputs(11157) <= (inputs(238)) and not (inputs(46));
    layer0_outputs(11158) <= (inputs(33)) xor (inputs(20));
    layer0_outputs(11159) <= not(inputs(93));
    layer0_outputs(11160) <= inputs(234);
    layer0_outputs(11161) <= inputs(79);
    layer0_outputs(11162) <= not((inputs(60)) and (inputs(218)));
    layer0_outputs(11163) <= (inputs(7)) xor (inputs(10));
    layer0_outputs(11164) <= (inputs(143)) or (inputs(64));
    layer0_outputs(11165) <= not((inputs(127)) or (inputs(48)));
    layer0_outputs(11166) <= (inputs(90)) or (inputs(223));
    layer0_outputs(11167) <= not((inputs(234)) and (inputs(35)));
    layer0_outputs(11168) <= inputs(143);
    layer0_outputs(11169) <= inputs(90);
    layer0_outputs(11170) <= inputs(249);
    layer0_outputs(11171) <= not(inputs(248)) or (inputs(81));
    layer0_outputs(11172) <= not((inputs(253)) or (inputs(0)));
    layer0_outputs(11173) <= not(inputs(199));
    layer0_outputs(11174) <= not((inputs(223)) or (inputs(168)));
    layer0_outputs(11175) <= inputs(107);
    layer0_outputs(11176) <= not((inputs(100)) or (inputs(180)));
    layer0_outputs(11177) <= (inputs(244)) and not (inputs(173));
    layer0_outputs(11178) <= not((inputs(144)) or (inputs(136)));
    layer0_outputs(11179) <= not(inputs(24));
    layer0_outputs(11180) <= inputs(9);
    layer0_outputs(11181) <= (inputs(115)) xor (inputs(112));
    layer0_outputs(11182) <= (inputs(16)) or (inputs(158));
    layer0_outputs(11183) <= (inputs(191)) or (inputs(6));
    layer0_outputs(11184) <= not((inputs(216)) xor (inputs(0)));
    layer0_outputs(11185) <= (inputs(41)) or (inputs(39));
    layer0_outputs(11186) <= (inputs(133)) or (inputs(129));
    layer0_outputs(11187) <= not(inputs(115));
    layer0_outputs(11188) <= not(inputs(37)) or (inputs(128));
    layer0_outputs(11189) <= (inputs(227)) and not (inputs(240));
    layer0_outputs(11190) <= (inputs(142)) or (inputs(162));
    layer0_outputs(11191) <= (inputs(71)) and not (inputs(78));
    layer0_outputs(11192) <= not((inputs(20)) or (inputs(40)));
    layer0_outputs(11193) <= (inputs(250)) or (inputs(223));
    layer0_outputs(11194) <= (inputs(44)) and not (inputs(237));
    layer0_outputs(11195) <= (inputs(147)) or (inputs(30));
    layer0_outputs(11196) <= not((inputs(73)) xor (inputs(226)));
    layer0_outputs(11197) <= not((inputs(11)) xor (inputs(153)));
    layer0_outputs(11198) <= inputs(214);
    layer0_outputs(11199) <= inputs(41);
    layer0_outputs(11200) <= not((inputs(166)) or (inputs(180)));
    layer0_outputs(11201) <= not(inputs(183)) or (inputs(155));
    layer0_outputs(11202) <= (inputs(248)) xor (inputs(12));
    layer0_outputs(11203) <= inputs(136);
    layer0_outputs(11204) <= inputs(78);
    layer0_outputs(11205) <= inputs(163);
    layer0_outputs(11206) <= (inputs(234)) xor (inputs(162));
    layer0_outputs(11207) <= (inputs(67)) xor (inputs(68));
    layer0_outputs(11208) <= (inputs(249)) or (inputs(129));
    layer0_outputs(11209) <= not((inputs(131)) or (inputs(197)));
    layer0_outputs(11210) <= (inputs(24)) and not (inputs(243));
    layer0_outputs(11211) <= not((inputs(223)) and (inputs(226)));
    layer0_outputs(11212) <= (inputs(108)) and not (inputs(175));
    layer0_outputs(11213) <= inputs(70);
    layer0_outputs(11214) <= inputs(25);
    layer0_outputs(11215) <= not((inputs(131)) or (inputs(246)));
    layer0_outputs(11216) <= not(inputs(179)) or (inputs(109));
    layer0_outputs(11217) <= (inputs(84)) xor (inputs(184));
    layer0_outputs(11218) <= (inputs(97)) or (inputs(72));
    layer0_outputs(11219) <= (inputs(64)) xor (inputs(79));
    layer0_outputs(11220) <= not(inputs(181));
    layer0_outputs(11221) <= (inputs(43)) or (inputs(43));
    layer0_outputs(11222) <= not(inputs(161));
    layer0_outputs(11223) <= not(inputs(28));
    layer0_outputs(11224) <= not(inputs(27));
    layer0_outputs(11225) <= inputs(121);
    layer0_outputs(11226) <= (inputs(90)) xor (inputs(25));
    layer0_outputs(11227) <= not(inputs(130));
    layer0_outputs(11228) <= (inputs(167)) xor (inputs(95));
    layer0_outputs(11229) <= (inputs(45)) and not (inputs(252));
    layer0_outputs(11230) <= (inputs(7)) and not (inputs(167));
    layer0_outputs(11231) <= not(inputs(216)) or (inputs(140));
    layer0_outputs(11232) <= (inputs(76)) and not (inputs(29));
    layer0_outputs(11233) <= not((inputs(140)) and (inputs(140)));
    layer0_outputs(11234) <= not(inputs(40));
    layer0_outputs(11235) <= not((inputs(253)) or (inputs(151)));
    layer0_outputs(11236) <= (inputs(251)) or (inputs(236));
    layer0_outputs(11237) <= inputs(93);
    layer0_outputs(11238) <= (inputs(177)) or (inputs(173));
    layer0_outputs(11239) <= not((inputs(137)) xor (inputs(117)));
    layer0_outputs(11240) <= not((inputs(87)) xor (inputs(99)));
    layer0_outputs(11241) <= (inputs(129)) and not (inputs(20));
    layer0_outputs(11242) <= not((inputs(175)) xor (inputs(50)));
    layer0_outputs(11243) <= not(inputs(52));
    layer0_outputs(11244) <= not(inputs(9));
    layer0_outputs(11245) <= (inputs(90)) and not (inputs(233));
    layer0_outputs(11246) <= not(inputs(21));
    layer0_outputs(11247) <= (inputs(163)) and not (inputs(62));
    layer0_outputs(11248) <= not((inputs(131)) xor (inputs(58)));
    layer0_outputs(11249) <= not(inputs(183)) or (inputs(52));
    layer0_outputs(11250) <= not(inputs(132));
    layer0_outputs(11251) <= (inputs(116)) or (inputs(220));
    layer0_outputs(11252) <= (inputs(183)) and (inputs(141));
    layer0_outputs(11253) <= (inputs(22)) or (inputs(91));
    layer0_outputs(11254) <= (inputs(52)) xor (inputs(16));
    layer0_outputs(11255) <= not((inputs(151)) and (inputs(27)));
    layer0_outputs(11256) <= (inputs(52)) or (inputs(114));
    layer0_outputs(11257) <= not((inputs(104)) or (inputs(122)));
    layer0_outputs(11258) <= not(inputs(129));
    layer0_outputs(11259) <= inputs(197);
    layer0_outputs(11260) <= (inputs(173)) and not (inputs(167));
    layer0_outputs(11261) <= not((inputs(165)) xor (inputs(119)));
    layer0_outputs(11262) <= (inputs(106)) and not (inputs(179));
    layer0_outputs(11263) <= (inputs(228)) and not (inputs(95));
    layer0_outputs(11264) <= not((inputs(232)) and (inputs(134)));
    layer0_outputs(11265) <= not((inputs(226)) or (inputs(7)));
    layer0_outputs(11266) <= not(inputs(82)) or (inputs(191));
    layer0_outputs(11267) <= (inputs(9)) and not (inputs(29));
    layer0_outputs(11268) <= not(inputs(228));
    layer0_outputs(11269) <= not((inputs(73)) xor (inputs(68)));
    layer0_outputs(11270) <= not((inputs(205)) or (inputs(116)));
    layer0_outputs(11271) <= not((inputs(6)) xor (inputs(110)));
    layer0_outputs(11272) <= not(inputs(136));
    layer0_outputs(11273) <= inputs(211);
    layer0_outputs(11274) <= inputs(98);
    layer0_outputs(11275) <= inputs(107);
    layer0_outputs(11276) <= (inputs(72)) or (inputs(201));
    layer0_outputs(11277) <= inputs(236);
    layer0_outputs(11278) <= not(inputs(77)) or (inputs(240));
    layer0_outputs(11279) <= inputs(101);
    layer0_outputs(11280) <= not((inputs(217)) or (inputs(233)));
    layer0_outputs(11281) <= not((inputs(234)) and (inputs(248)));
    layer0_outputs(11282) <= not((inputs(57)) xor (inputs(74)));
    layer0_outputs(11283) <= not((inputs(102)) or (inputs(248)));
    layer0_outputs(11284) <= '0';
    layer0_outputs(11285) <= (inputs(109)) xor (inputs(64));
    layer0_outputs(11286) <= inputs(231);
    layer0_outputs(11287) <= inputs(163);
    layer0_outputs(11288) <= inputs(168);
    layer0_outputs(11289) <= (inputs(112)) and not (inputs(70));
    layer0_outputs(11290) <= inputs(229);
    layer0_outputs(11291) <= not((inputs(42)) and (inputs(205)));
    layer0_outputs(11292) <= (inputs(200)) and not (inputs(158));
    layer0_outputs(11293) <= inputs(231);
    layer0_outputs(11294) <= not(inputs(245));
    layer0_outputs(11295) <= not(inputs(197)) or (inputs(254));
    layer0_outputs(11296) <= (inputs(85)) xor (inputs(4));
    layer0_outputs(11297) <= not(inputs(170));
    layer0_outputs(11298) <= not((inputs(192)) or (inputs(227)));
    layer0_outputs(11299) <= inputs(8);
    layer0_outputs(11300) <= not((inputs(70)) and (inputs(218)));
    layer0_outputs(11301) <= (inputs(196)) or (inputs(47));
    layer0_outputs(11302) <= (inputs(146)) or (inputs(81));
    layer0_outputs(11303) <= not((inputs(246)) or (inputs(249)));
    layer0_outputs(11304) <= not((inputs(133)) xor (inputs(130)));
    layer0_outputs(11305) <= inputs(206);
    layer0_outputs(11306) <= not(inputs(77)) or (inputs(16));
    layer0_outputs(11307) <= not(inputs(183));
    layer0_outputs(11308) <= (inputs(31)) or (inputs(138));
    layer0_outputs(11309) <= not((inputs(47)) or (inputs(25)));
    layer0_outputs(11310) <= not((inputs(97)) xor (inputs(24)));
    layer0_outputs(11311) <= (inputs(78)) xor (inputs(66));
    layer0_outputs(11312) <= (inputs(64)) xor (inputs(199));
    layer0_outputs(11313) <= not(inputs(189));
    layer0_outputs(11314) <= not((inputs(188)) or (inputs(180)));
    layer0_outputs(11315) <= not((inputs(220)) xor (inputs(173)));
    layer0_outputs(11316) <= (inputs(73)) xor (inputs(0));
    layer0_outputs(11317) <= not(inputs(156)) or (inputs(15));
    layer0_outputs(11318) <= not((inputs(11)) xor (inputs(160)));
    layer0_outputs(11319) <= not((inputs(112)) or (inputs(90)));
    layer0_outputs(11320) <= not(inputs(2));
    layer0_outputs(11321) <= not((inputs(85)) xor (inputs(252)));
    layer0_outputs(11322) <= inputs(115);
    layer0_outputs(11323) <= not(inputs(187)) or (inputs(6));
    layer0_outputs(11324) <= not((inputs(116)) or (inputs(11)));
    layer0_outputs(11325) <= (inputs(89)) or (inputs(132));
    layer0_outputs(11326) <= (inputs(194)) or (inputs(167));
    layer0_outputs(11327) <= not((inputs(78)) xor (inputs(222)));
    layer0_outputs(11328) <= inputs(51);
    layer0_outputs(11329) <= not(inputs(148)) or (inputs(64));
    layer0_outputs(11330) <= (inputs(179)) and not (inputs(31));
    layer0_outputs(11331) <= not((inputs(202)) xor (inputs(11)));
    layer0_outputs(11332) <= not((inputs(228)) or (inputs(221)));
    layer0_outputs(11333) <= not((inputs(83)) xor (inputs(115)));
    layer0_outputs(11334) <= (inputs(240)) or (inputs(56));
    layer0_outputs(11335) <= (inputs(5)) and not (inputs(126));
    layer0_outputs(11336) <= (inputs(235)) or (inputs(95));
    layer0_outputs(11337) <= inputs(154);
    layer0_outputs(11338) <= inputs(132);
    layer0_outputs(11339) <= (inputs(73)) or (inputs(204));
    layer0_outputs(11340) <= not((inputs(64)) and (inputs(228)));
    layer0_outputs(11341) <= inputs(64);
    layer0_outputs(11342) <= (inputs(94)) or (inputs(176));
    layer0_outputs(11343) <= not(inputs(221)) or (inputs(224));
    layer0_outputs(11344) <= (inputs(248)) or (inputs(159));
    layer0_outputs(11345) <= (inputs(232)) and (inputs(163));
    layer0_outputs(11346) <= (inputs(184)) or (inputs(224));
    layer0_outputs(11347) <= inputs(125);
    layer0_outputs(11348) <= (inputs(210)) or (inputs(179));
    layer0_outputs(11349) <= (inputs(34)) and not (inputs(128));
    layer0_outputs(11350) <= not(inputs(190)) or (inputs(253));
    layer0_outputs(11351) <= not(inputs(231));
    layer0_outputs(11352) <= '0';
    layer0_outputs(11353) <= not((inputs(207)) or (inputs(98)));
    layer0_outputs(11354) <= not((inputs(164)) xor (inputs(162)));
    layer0_outputs(11355) <= not((inputs(23)) xor (inputs(119)));
    layer0_outputs(11356) <= not(inputs(58)) or (inputs(242));
    layer0_outputs(11357) <= inputs(62);
    layer0_outputs(11358) <= not((inputs(96)) and (inputs(75)));
    layer0_outputs(11359) <= not(inputs(210));
    layer0_outputs(11360) <= inputs(42);
    layer0_outputs(11361) <= (inputs(214)) and not (inputs(39));
    layer0_outputs(11362) <= (inputs(77)) or (inputs(96));
    layer0_outputs(11363) <= (inputs(85)) and not (inputs(250));
    layer0_outputs(11364) <= not((inputs(35)) xor (inputs(140)));
    layer0_outputs(11365) <= not((inputs(137)) or (inputs(109)));
    layer0_outputs(11366) <= not(inputs(33)) or (inputs(152));
    layer0_outputs(11367) <= not(inputs(87));
    layer0_outputs(11368) <= (inputs(43)) xor (inputs(13));
    layer0_outputs(11369) <= (inputs(125)) or (inputs(103));
    layer0_outputs(11370) <= inputs(110);
    layer0_outputs(11371) <= not(inputs(19)) or (inputs(81));
    layer0_outputs(11372) <= (inputs(104)) and not (inputs(62));
    layer0_outputs(11373) <= not(inputs(212)) or (inputs(19));
    layer0_outputs(11374) <= (inputs(7)) and not (inputs(87));
    layer0_outputs(11375) <= not(inputs(230));
    layer0_outputs(11376) <= not((inputs(12)) or (inputs(24)));
    layer0_outputs(11377) <= inputs(156);
    layer0_outputs(11378) <= inputs(53);
    layer0_outputs(11379) <= not(inputs(77)) or (inputs(16));
    layer0_outputs(11380) <= (inputs(147)) or (inputs(148));
    layer0_outputs(11381) <= (inputs(120)) and (inputs(123));
    layer0_outputs(11382) <= not((inputs(173)) or (inputs(155)));
    layer0_outputs(11383) <= not((inputs(18)) or (inputs(154)));
    layer0_outputs(11384) <= not(inputs(164));
    layer0_outputs(11385) <= inputs(9);
    layer0_outputs(11386) <= (inputs(253)) and not (inputs(143));
    layer0_outputs(11387) <= not(inputs(140));
    layer0_outputs(11388) <= (inputs(31)) xor (inputs(114));
    layer0_outputs(11389) <= not(inputs(182)) or (inputs(84));
    layer0_outputs(11390) <= (inputs(73)) and not (inputs(66));
    layer0_outputs(11391) <= not((inputs(243)) or (inputs(193)));
    layer0_outputs(11392) <= (inputs(180)) xor (inputs(106));
    layer0_outputs(11393) <= not((inputs(22)) and (inputs(26)));
    layer0_outputs(11394) <= not((inputs(66)) or (inputs(103)));
    layer0_outputs(11395) <= not((inputs(137)) or (inputs(46)));
    layer0_outputs(11396) <= not((inputs(152)) and (inputs(25)));
    layer0_outputs(11397) <= not(inputs(30));
    layer0_outputs(11398) <= not(inputs(191)) or (inputs(2));
    layer0_outputs(11399) <= not((inputs(83)) or (inputs(29)));
    layer0_outputs(11400) <= not((inputs(30)) xor (inputs(94)));
    layer0_outputs(11401) <= (inputs(45)) or (inputs(127));
    layer0_outputs(11402) <= inputs(226);
    layer0_outputs(11403) <= (inputs(219)) and not (inputs(207));
    layer0_outputs(11404) <= not(inputs(106)) or (inputs(138));
    layer0_outputs(11405) <= (inputs(198)) and (inputs(198));
    layer0_outputs(11406) <= not(inputs(0));
    layer0_outputs(11407) <= not((inputs(176)) xor (inputs(234)));
    layer0_outputs(11408) <= not(inputs(133)) or (inputs(35));
    layer0_outputs(11409) <= (inputs(177)) and not (inputs(68));
    layer0_outputs(11410) <= inputs(99);
    layer0_outputs(11411) <= (inputs(38)) and not (inputs(205));
    layer0_outputs(11412) <= not((inputs(251)) or (inputs(97)));
    layer0_outputs(11413) <= (inputs(74)) or (inputs(235));
    layer0_outputs(11414) <= not((inputs(114)) or (inputs(236)));
    layer0_outputs(11415) <= not((inputs(168)) xor (inputs(210)));
    layer0_outputs(11416) <= (inputs(182)) and not (inputs(221));
    layer0_outputs(11417) <= not(inputs(84)) or (inputs(185));
    layer0_outputs(11418) <= (inputs(209)) and not (inputs(116));
    layer0_outputs(11419) <= not(inputs(55)) or (inputs(111));
    layer0_outputs(11420) <= not(inputs(142));
    layer0_outputs(11421) <= (inputs(128)) or (inputs(138));
    layer0_outputs(11422) <= not((inputs(119)) or (inputs(34)));
    layer0_outputs(11423) <= (inputs(24)) and not (inputs(115));
    layer0_outputs(11424) <= not((inputs(237)) or (inputs(137)));
    layer0_outputs(11425) <= inputs(168);
    layer0_outputs(11426) <= not((inputs(147)) or (inputs(199)));
    layer0_outputs(11427) <= not(inputs(121)) or (inputs(191));
    layer0_outputs(11428) <= not(inputs(8)) or (inputs(80));
    layer0_outputs(11429) <= (inputs(208)) xor (inputs(86));
    layer0_outputs(11430) <= (inputs(199)) and not (inputs(129));
    layer0_outputs(11431) <= not((inputs(159)) or (inputs(13)));
    layer0_outputs(11432) <= not(inputs(32));
    layer0_outputs(11433) <= not(inputs(25));
    layer0_outputs(11434) <= not((inputs(169)) or (inputs(68)));
    layer0_outputs(11435) <= inputs(148);
    layer0_outputs(11436) <= (inputs(90)) or (inputs(62));
    layer0_outputs(11437) <= not((inputs(85)) or (inputs(190)));
    layer0_outputs(11438) <= (inputs(199)) xor (inputs(245));
    layer0_outputs(11439) <= not(inputs(114));
    layer0_outputs(11440) <= (inputs(142)) xor (inputs(221));
    layer0_outputs(11441) <= not(inputs(118)) or (inputs(32));
    layer0_outputs(11442) <= not(inputs(108));
    layer0_outputs(11443) <= inputs(63);
    layer0_outputs(11444) <= not(inputs(210)) or (inputs(80));
    layer0_outputs(11445) <= not(inputs(153));
    layer0_outputs(11446) <= (inputs(182)) or (inputs(166));
    layer0_outputs(11447) <= (inputs(86)) and not (inputs(147));
    layer0_outputs(11448) <= (inputs(189)) xor (inputs(63));
    layer0_outputs(11449) <= not((inputs(211)) or (inputs(247)));
    layer0_outputs(11450) <= inputs(115);
    layer0_outputs(11451) <= not(inputs(139));
    layer0_outputs(11452) <= (inputs(117)) or (inputs(8));
    layer0_outputs(11453) <= (inputs(129)) or (inputs(231));
    layer0_outputs(11454) <= not(inputs(210));
    layer0_outputs(11455) <= (inputs(47)) or (inputs(44));
    layer0_outputs(11456) <= (inputs(128)) or (inputs(108));
    layer0_outputs(11457) <= (inputs(251)) xor (inputs(212));
    layer0_outputs(11458) <= not((inputs(105)) or (inputs(125)));
    layer0_outputs(11459) <= not((inputs(95)) or (inputs(177)));
    layer0_outputs(11460) <= inputs(27);
    layer0_outputs(11461) <= inputs(24);
    layer0_outputs(11462) <= not(inputs(179)) or (inputs(17));
    layer0_outputs(11463) <= not((inputs(116)) xor (inputs(211)));
    layer0_outputs(11464) <= not(inputs(67)) or (inputs(227));
    layer0_outputs(11465) <= inputs(41);
    layer0_outputs(11466) <= not((inputs(210)) or (inputs(205)));
    layer0_outputs(11467) <= not((inputs(68)) or (inputs(134)));
    layer0_outputs(11468) <= (inputs(179)) and (inputs(114));
    layer0_outputs(11469) <= inputs(192);
    layer0_outputs(11470) <= (inputs(191)) or (inputs(24));
    layer0_outputs(11471) <= not((inputs(142)) or (inputs(58)));
    layer0_outputs(11472) <= not((inputs(177)) or (inputs(148)));
    layer0_outputs(11473) <= not(inputs(197)) or (inputs(28));
    layer0_outputs(11474) <= (inputs(47)) or (inputs(19));
    layer0_outputs(11475) <= (inputs(142)) and not (inputs(12));
    layer0_outputs(11476) <= (inputs(17)) or (inputs(55));
    layer0_outputs(11477) <= not(inputs(191));
    layer0_outputs(11478) <= (inputs(113)) or (inputs(16));
    layer0_outputs(11479) <= inputs(120);
    layer0_outputs(11480) <= not(inputs(200));
    layer0_outputs(11481) <= not((inputs(68)) or (inputs(94)));
    layer0_outputs(11482) <= not(inputs(59));
    layer0_outputs(11483) <= (inputs(108)) or (inputs(83));
    layer0_outputs(11484) <= (inputs(251)) xor (inputs(149));
    layer0_outputs(11485) <= (inputs(115)) or (inputs(246));
    layer0_outputs(11486) <= not((inputs(20)) or (inputs(146)));
    layer0_outputs(11487) <= not((inputs(109)) xor (inputs(83)));
    layer0_outputs(11488) <= not((inputs(145)) or (inputs(197)));
    layer0_outputs(11489) <= not((inputs(19)) xor (inputs(93)));
    layer0_outputs(11490) <= not(inputs(247)) or (inputs(239));
    layer0_outputs(11491) <= (inputs(162)) xor (inputs(231));
    layer0_outputs(11492) <= not((inputs(29)) xor (inputs(171)));
    layer0_outputs(11493) <= not(inputs(145));
    layer0_outputs(11494) <= inputs(204);
    layer0_outputs(11495) <= not((inputs(165)) or (inputs(92)));
    layer0_outputs(11496) <= not((inputs(237)) xor (inputs(46)));
    layer0_outputs(11497) <= not((inputs(49)) or (inputs(48)));
    layer0_outputs(11498) <= (inputs(243)) or (inputs(143));
    layer0_outputs(11499) <= not(inputs(43)) or (inputs(92));
    layer0_outputs(11500) <= (inputs(164)) and not (inputs(114));
    layer0_outputs(11501) <= (inputs(122)) and (inputs(129));
    layer0_outputs(11502) <= not(inputs(43));
    layer0_outputs(11503) <= not(inputs(112)) or (inputs(237));
    layer0_outputs(11504) <= (inputs(251)) or (inputs(222));
    layer0_outputs(11505) <= (inputs(49)) xor (inputs(201));
    layer0_outputs(11506) <= (inputs(219)) and not (inputs(117));
    layer0_outputs(11507) <= not((inputs(101)) xor (inputs(133)));
    layer0_outputs(11508) <= not((inputs(183)) xor (inputs(63)));
    layer0_outputs(11509) <= inputs(242);
    layer0_outputs(11510) <= (inputs(42)) or (inputs(58));
    layer0_outputs(11511) <= not((inputs(87)) xor (inputs(145)));
    layer0_outputs(11512) <= not(inputs(109)) or (inputs(227));
    layer0_outputs(11513) <= not((inputs(6)) xor (inputs(130)));
    layer0_outputs(11514) <= (inputs(119)) and not (inputs(20));
    layer0_outputs(11515) <= not(inputs(10));
    layer0_outputs(11516) <= inputs(226);
    layer0_outputs(11517) <= (inputs(35)) xor (inputs(27));
    layer0_outputs(11518) <= (inputs(254)) xor (inputs(165));
    layer0_outputs(11519) <= not((inputs(75)) xor (inputs(26)));
    layer0_outputs(11520) <= not((inputs(236)) or (inputs(220)));
    layer0_outputs(11521) <= inputs(228);
    layer0_outputs(11522) <= not(inputs(202)) or (inputs(79));
    layer0_outputs(11523) <= not(inputs(53)) or (inputs(217));
    layer0_outputs(11524) <= (inputs(228)) and not (inputs(90));
    layer0_outputs(11525) <= not((inputs(124)) or (inputs(99)));
    layer0_outputs(11526) <= (inputs(77)) xor (inputs(65));
    layer0_outputs(11527) <= not(inputs(152));
    layer0_outputs(11528) <= not((inputs(6)) xor (inputs(53)));
    layer0_outputs(11529) <= (inputs(40)) and not (inputs(102));
    layer0_outputs(11530) <= not((inputs(139)) or (inputs(220)));
    layer0_outputs(11531) <= inputs(26);
    layer0_outputs(11532) <= (inputs(100)) xor (inputs(119));
    layer0_outputs(11533) <= not(inputs(40));
    layer0_outputs(11534) <= not(inputs(184));
    layer0_outputs(11535) <= (inputs(249)) and not (inputs(102));
    layer0_outputs(11536) <= (inputs(61)) and not (inputs(135));
    layer0_outputs(11537) <= (inputs(233)) and (inputs(30));
    layer0_outputs(11538) <= not((inputs(28)) or (inputs(84)));
    layer0_outputs(11539) <= not((inputs(52)) or (inputs(77)));
    layer0_outputs(11540) <= not((inputs(12)) and (inputs(99)));
    layer0_outputs(11541) <= (inputs(98)) and not (inputs(56));
    layer0_outputs(11542) <= (inputs(92)) and not (inputs(192));
    layer0_outputs(11543) <= not((inputs(56)) xor (inputs(41)));
    layer0_outputs(11544) <= (inputs(181)) and not (inputs(207));
    layer0_outputs(11545) <= (inputs(100)) and (inputs(9));
    layer0_outputs(11546) <= (inputs(47)) and not (inputs(109));
    layer0_outputs(11547) <= (inputs(22)) and not (inputs(68));
    layer0_outputs(11548) <= inputs(78);
    layer0_outputs(11549) <= not((inputs(173)) xor (inputs(165)));
    layer0_outputs(11550) <= not(inputs(236)) or (inputs(158));
    layer0_outputs(11551) <= inputs(155);
    layer0_outputs(11552) <= not(inputs(152));
    layer0_outputs(11553) <= not(inputs(124));
    layer0_outputs(11554) <= not(inputs(39));
    layer0_outputs(11555) <= not((inputs(209)) xor (inputs(33)));
    layer0_outputs(11556) <= not((inputs(162)) xor (inputs(230)));
    layer0_outputs(11557) <= (inputs(187)) and not (inputs(63));
    layer0_outputs(11558) <= inputs(74);
    layer0_outputs(11559) <= (inputs(178)) xor (inputs(234));
    layer0_outputs(11560) <= (inputs(177)) or (inputs(127));
    layer0_outputs(11561) <= (inputs(10)) and not (inputs(195));
    layer0_outputs(11562) <= (inputs(85)) and not (inputs(17));
    layer0_outputs(11563) <= not((inputs(91)) xor (inputs(160)));
    layer0_outputs(11564) <= inputs(24);
    layer0_outputs(11565) <= not(inputs(136));
    layer0_outputs(11566) <= not((inputs(160)) xor (inputs(219)));
    layer0_outputs(11567) <= (inputs(179)) xor (inputs(250));
    layer0_outputs(11568) <= not((inputs(178)) xor (inputs(246)));
    layer0_outputs(11569) <= (inputs(6)) and not (inputs(218));
    layer0_outputs(11570) <= not(inputs(15));
    layer0_outputs(11571) <= not((inputs(186)) or (inputs(86)));
    layer0_outputs(11572) <= inputs(222);
    layer0_outputs(11573) <= not(inputs(108));
    layer0_outputs(11574) <= inputs(208);
    layer0_outputs(11575) <= not((inputs(2)) xor (inputs(123)));
    layer0_outputs(11576) <= not((inputs(30)) or (inputs(233)));
    layer0_outputs(11577) <= not(inputs(141)) or (inputs(243));
    layer0_outputs(11578) <= not((inputs(4)) xor (inputs(100)));
    layer0_outputs(11579) <= not(inputs(128));
    layer0_outputs(11580) <= (inputs(17)) or (inputs(58));
    layer0_outputs(11581) <= not((inputs(128)) or (inputs(182)));
    layer0_outputs(11582) <= not(inputs(148)) or (inputs(31));
    layer0_outputs(11583) <= (inputs(188)) xor (inputs(77));
    layer0_outputs(11584) <= not((inputs(22)) xor (inputs(242)));
    layer0_outputs(11585) <= inputs(162);
    layer0_outputs(11586) <= inputs(146);
    layer0_outputs(11587) <= not((inputs(214)) and (inputs(166)));
    layer0_outputs(11588) <= (inputs(209)) or (inputs(239));
    layer0_outputs(11589) <= (inputs(171)) xor (inputs(123));
    layer0_outputs(11590) <= not((inputs(170)) or (inputs(243)));
    layer0_outputs(11591) <= (inputs(233)) and (inputs(181));
    layer0_outputs(11592) <= not(inputs(106));
    layer0_outputs(11593) <= (inputs(75)) or (inputs(174));
    layer0_outputs(11594) <= (inputs(151)) and not (inputs(170));
    layer0_outputs(11595) <= (inputs(46)) and not (inputs(252));
    layer0_outputs(11596) <= not((inputs(170)) xor (inputs(5)));
    layer0_outputs(11597) <= not(inputs(23));
    layer0_outputs(11598) <= not((inputs(106)) xor (inputs(73)));
    layer0_outputs(11599) <= (inputs(226)) xor (inputs(99));
    layer0_outputs(11600) <= (inputs(178)) xor (inputs(191));
    layer0_outputs(11601) <= not(inputs(217));
    layer0_outputs(11602) <= (inputs(106)) and not (inputs(166));
    layer0_outputs(11603) <= inputs(190);
    layer0_outputs(11604) <= (inputs(120)) or (inputs(124));
    layer0_outputs(11605) <= (inputs(98)) or (inputs(42));
    layer0_outputs(11606) <= (inputs(222)) xor (inputs(95));
    layer0_outputs(11607) <= inputs(187);
    layer0_outputs(11608) <= inputs(233);
    layer0_outputs(11609) <= not(inputs(249));
    layer0_outputs(11610) <= not((inputs(44)) or (inputs(174)));
    layer0_outputs(11611) <= not(inputs(186)) or (inputs(50));
    layer0_outputs(11612) <= not((inputs(65)) or (inputs(27)));
    layer0_outputs(11613) <= '1';
    layer0_outputs(11614) <= (inputs(210)) or (inputs(26));
    layer0_outputs(11615) <= (inputs(59)) and not (inputs(4));
    layer0_outputs(11616) <= inputs(94);
    layer0_outputs(11617) <= inputs(217);
    layer0_outputs(11618) <= not(inputs(166));
    layer0_outputs(11619) <= not(inputs(158)) or (inputs(243));
    layer0_outputs(11620) <= not((inputs(173)) or (inputs(185)));
    layer0_outputs(11621) <= not((inputs(192)) or (inputs(171)));
    layer0_outputs(11622) <= not(inputs(222));
    layer0_outputs(11623) <= (inputs(231)) and not (inputs(117));
    layer0_outputs(11624) <= (inputs(61)) or (inputs(115));
    layer0_outputs(11625) <= (inputs(202)) and (inputs(133));
    layer0_outputs(11626) <= not((inputs(83)) xor (inputs(19)));
    layer0_outputs(11627) <= (inputs(42)) and not (inputs(183));
    layer0_outputs(11628) <= not((inputs(59)) and (inputs(55)));
    layer0_outputs(11629) <= (inputs(162)) or (inputs(93));
    layer0_outputs(11630) <= inputs(229);
    layer0_outputs(11631) <= not((inputs(190)) xor (inputs(116)));
    layer0_outputs(11632) <= not(inputs(245)) or (inputs(112));
    layer0_outputs(11633) <= not(inputs(231)) or (inputs(238));
    layer0_outputs(11634) <= not(inputs(248));
    layer0_outputs(11635) <= not(inputs(193)) or (inputs(255));
    layer0_outputs(11636) <= not(inputs(24));
    layer0_outputs(11637) <= not((inputs(5)) or (inputs(85)));
    layer0_outputs(11638) <= (inputs(148)) or (inputs(31));
    layer0_outputs(11639) <= not((inputs(200)) or (inputs(167)));
    layer0_outputs(11640) <= (inputs(65)) xor (inputs(102));
    layer0_outputs(11641) <= not(inputs(5)) or (inputs(212));
    layer0_outputs(11642) <= not(inputs(113));
    layer0_outputs(11643) <= not(inputs(171));
    layer0_outputs(11644) <= inputs(42);
    layer0_outputs(11645) <= not((inputs(158)) or (inputs(27)));
    layer0_outputs(11646) <= not((inputs(228)) xor (inputs(82)));
    layer0_outputs(11647) <= (inputs(55)) and not (inputs(176));
    layer0_outputs(11648) <= inputs(165);
    layer0_outputs(11649) <= not(inputs(65));
    layer0_outputs(11650) <= (inputs(232)) xor (inputs(199));
    layer0_outputs(11651) <= not((inputs(85)) xor (inputs(255)));
    layer0_outputs(11652) <= not((inputs(81)) or (inputs(98)));
    layer0_outputs(11653) <= not(inputs(246));
    layer0_outputs(11654) <= (inputs(35)) or (inputs(140));
    layer0_outputs(11655) <= not((inputs(199)) or (inputs(175)));
    layer0_outputs(11656) <= not(inputs(148));
    layer0_outputs(11657) <= not(inputs(131));
    layer0_outputs(11658) <= (inputs(63)) or (inputs(72));
    layer0_outputs(11659) <= not(inputs(184)) or (inputs(244));
    layer0_outputs(11660) <= (inputs(126)) xor (inputs(206));
    layer0_outputs(11661) <= inputs(32);
    layer0_outputs(11662) <= inputs(223);
    layer0_outputs(11663) <= (inputs(196)) and not (inputs(186));
    layer0_outputs(11664) <= (inputs(119)) and not (inputs(227));
    layer0_outputs(11665) <= inputs(170);
    layer0_outputs(11666) <= inputs(24);
    layer0_outputs(11667) <= not(inputs(107));
    layer0_outputs(11668) <= (inputs(48)) xor (inputs(149));
    layer0_outputs(11669) <= (inputs(68)) or (inputs(38));
    layer0_outputs(11670) <= not((inputs(38)) and (inputs(35)));
    layer0_outputs(11671) <= (inputs(206)) or (inputs(30));
    layer0_outputs(11672) <= not((inputs(128)) xor (inputs(161)));
    layer0_outputs(11673) <= (inputs(36)) or (inputs(174));
    layer0_outputs(11674) <= inputs(17);
    layer0_outputs(11675) <= (inputs(129)) or (inputs(84));
    layer0_outputs(11676) <= not(inputs(58));
    layer0_outputs(11677) <= inputs(226);
    layer0_outputs(11678) <= (inputs(129)) or (inputs(91));
    layer0_outputs(11679) <= (inputs(66)) xor (inputs(131));
    layer0_outputs(11680) <= not((inputs(224)) or (inputs(238)));
    layer0_outputs(11681) <= (inputs(27)) xor (inputs(134));
    layer0_outputs(11682) <= not(inputs(243));
    layer0_outputs(11683) <= not((inputs(156)) xor (inputs(7)));
    layer0_outputs(11684) <= not(inputs(45));
    layer0_outputs(11685) <= not(inputs(93));
    layer0_outputs(11686) <= not((inputs(129)) or (inputs(50)));
    layer0_outputs(11687) <= not((inputs(46)) and (inputs(54)));
    layer0_outputs(11688) <= (inputs(51)) xor (inputs(9));
    layer0_outputs(11689) <= inputs(62);
    layer0_outputs(11690) <= not((inputs(15)) and (inputs(251)));
    layer0_outputs(11691) <= (inputs(136)) and not (inputs(12));
    layer0_outputs(11692) <= (inputs(202)) and not (inputs(241));
    layer0_outputs(11693) <= inputs(171);
    layer0_outputs(11694) <= (inputs(28)) and not (inputs(116));
    layer0_outputs(11695) <= not((inputs(224)) or (inputs(124)));
    layer0_outputs(11696) <= (inputs(87)) or (inputs(116));
    layer0_outputs(11697) <= not(inputs(221));
    layer0_outputs(11698) <= not(inputs(137));
    layer0_outputs(11699) <= (inputs(46)) or (inputs(19));
    layer0_outputs(11700) <= not((inputs(4)) or (inputs(249)));
    layer0_outputs(11701) <= inputs(202);
    layer0_outputs(11702) <= (inputs(238)) or (inputs(126));
    layer0_outputs(11703) <= (inputs(239)) xor (inputs(195));
    layer0_outputs(11704) <= not(inputs(175));
    layer0_outputs(11705) <= (inputs(35)) and not (inputs(1));
    layer0_outputs(11706) <= (inputs(30)) xor (inputs(43));
    layer0_outputs(11707) <= inputs(211);
    layer0_outputs(11708) <= inputs(234);
    layer0_outputs(11709) <= (inputs(0)) and not (inputs(75));
    layer0_outputs(11710) <= not((inputs(191)) and (inputs(81)));
    layer0_outputs(11711) <= inputs(70);
    layer0_outputs(11712) <= (inputs(164)) xor (inputs(102));
    layer0_outputs(11713) <= not((inputs(189)) or (inputs(43)));
    layer0_outputs(11714) <= not(inputs(103)) or (inputs(11));
    layer0_outputs(11715) <= not(inputs(156)) or (inputs(244));
    layer0_outputs(11716) <= (inputs(246)) and not (inputs(200));
    layer0_outputs(11717) <= inputs(205);
    layer0_outputs(11718) <= not(inputs(213)) or (inputs(60));
    layer0_outputs(11719) <= not(inputs(94));
    layer0_outputs(11720) <= '0';
    layer0_outputs(11721) <= (inputs(86)) and not (inputs(142));
    layer0_outputs(11722) <= inputs(157);
    layer0_outputs(11723) <= not((inputs(231)) and (inputs(217)));
    layer0_outputs(11724) <= inputs(109);
    layer0_outputs(11725) <= not((inputs(32)) or (inputs(228)));
    layer0_outputs(11726) <= not(inputs(201)) or (inputs(209));
    layer0_outputs(11727) <= (inputs(97)) and not (inputs(123));
    layer0_outputs(11728) <= inputs(199);
    layer0_outputs(11729) <= not(inputs(168)) or (inputs(244));
    layer0_outputs(11730) <= (inputs(124)) and not (inputs(16));
    layer0_outputs(11731) <= inputs(230);
    layer0_outputs(11732) <= not(inputs(97)) or (inputs(80));
    layer0_outputs(11733) <= not((inputs(246)) or (inputs(42)));
    layer0_outputs(11734) <= not(inputs(174));
    layer0_outputs(11735) <= (inputs(0)) xor (inputs(78));
    layer0_outputs(11736) <= (inputs(44)) and not (inputs(208));
    layer0_outputs(11737) <= not(inputs(174));
    layer0_outputs(11738) <= inputs(42);
    layer0_outputs(11739) <= '0';
    layer0_outputs(11740) <= not(inputs(242)) or (inputs(208));
    layer0_outputs(11741) <= not((inputs(186)) or (inputs(78)));
    layer0_outputs(11742) <= not(inputs(102));
    layer0_outputs(11743) <= not((inputs(124)) or (inputs(22)));
    layer0_outputs(11744) <= not((inputs(255)) xor (inputs(209)));
    layer0_outputs(11745) <= (inputs(104)) and not (inputs(50));
    layer0_outputs(11746) <= (inputs(95)) or (inputs(23));
    layer0_outputs(11747) <= not((inputs(26)) or (inputs(3)));
    layer0_outputs(11748) <= not((inputs(57)) or (inputs(253)));
    layer0_outputs(11749) <= inputs(232);
    layer0_outputs(11750) <= inputs(135);
    layer0_outputs(11751) <= not((inputs(166)) or (inputs(167)));
    layer0_outputs(11752) <= not(inputs(232));
    layer0_outputs(11753) <= (inputs(239)) xor (inputs(110));
    layer0_outputs(11754) <= inputs(92);
    layer0_outputs(11755) <= (inputs(245)) and not (inputs(91));
    layer0_outputs(11756) <= (inputs(40)) and not (inputs(252));
    layer0_outputs(11757) <= (inputs(48)) or (inputs(180));
    layer0_outputs(11758) <= not(inputs(98));
    layer0_outputs(11759) <= not((inputs(154)) and (inputs(156)));
    layer0_outputs(11760) <= not(inputs(103));
    layer0_outputs(11761) <= (inputs(213)) or (inputs(142));
    layer0_outputs(11762) <= (inputs(57)) and not (inputs(80));
    layer0_outputs(11763) <= not(inputs(32));
    layer0_outputs(11764) <= (inputs(94)) xor (inputs(49));
    layer0_outputs(11765) <= (inputs(186)) and (inputs(143));
    layer0_outputs(11766) <= not(inputs(58)) or (inputs(209));
    layer0_outputs(11767) <= inputs(40);
    layer0_outputs(11768) <= not((inputs(213)) xor (inputs(200)));
    layer0_outputs(11769) <= (inputs(82)) and not (inputs(62));
    layer0_outputs(11770) <= (inputs(21)) and not (inputs(252));
    layer0_outputs(11771) <= inputs(122);
    layer0_outputs(11772) <= inputs(40);
    layer0_outputs(11773) <= (inputs(219)) xor (inputs(36));
    layer0_outputs(11774) <= not(inputs(109));
    layer0_outputs(11775) <= not((inputs(139)) or (inputs(14)));
    layer0_outputs(11776) <= not(inputs(69));
    layer0_outputs(11777) <= (inputs(205)) xor (inputs(92));
    layer0_outputs(11778) <= not(inputs(104)) or (inputs(49));
    layer0_outputs(11779) <= inputs(102);
    layer0_outputs(11780) <= inputs(47);
    layer0_outputs(11781) <= '0';
    layer0_outputs(11782) <= not(inputs(253));
    layer0_outputs(11783) <= not((inputs(138)) or (inputs(9)));
    layer0_outputs(11784) <= (inputs(205)) or (inputs(18));
    layer0_outputs(11785) <= not((inputs(85)) xor (inputs(122)));
    layer0_outputs(11786) <= (inputs(253)) and not (inputs(206));
    layer0_outputs(11787) <= (inputs(150)) or (inputs(19));
    layer0_outputs(11788) <= not(inputs(54));
    layer0_outputs(11789) <= not((inputs(145)) or (inputs(125)));
    layer0_outputs(11790) <= not(inputs(179));
    layer0_outputs(11791) <= not((inputs(169)) xor (inputs(141)));
    layer0_outputs(11792) <= not((inputs(160)) or (inputs(194)));
    layer0_outputs(11793) <= not(inputs(93)) or (inputs(222));
    layer0_outputs(11794) <= (inputs(210)) and (inputs(168));
    layer0_outputs(11795) <= (inputs(28)) xor (inputs(17));
    layer0_outputs(11796) <= (inputs(25)) or (inputs(57));
    layer0_outputs(11797) <= not((inputs(168)) or (inputs(32)));
    layer0_outputs(11798) <= not((inputs(106)) and (inputs(28)));
    layer0_outputs(11799) <= (inputs(236)) and not (inputs(196));
    layer0_outputs(11800) <= not(inputs(176)) or (inputs(204));
    layer0_outputs(11801) <= not((inputs(159)) xor (inputs(234)));
    layer0_outputs(11802) <= not(inputs(225));
    layer0_outputs(11803) <= not(inputs(198)) or (inputs(190));
    layer0_outputs(11804) <= not((inputs(117)) or (inputs(190)));
    layer0_outputs(11805) <= not(inputs(77)) or (inputs(121));
    layer0_outputs(11806) <= not((inputs(120)) xor (inputs(147)));
    layer0_outputs(11807) <= not(inputs(129));
    layer0_outputs(11808) <= not((inputs(210)) or (inputs(147)));
    layer0_outputs(11809) <= inputs(19);
    layer0_outputs(11810) <= (inputs(203)) or (inputs(119));
    layer0_outputs(11811) <= not(inputs(16)) or (inputs(222));
    layer0_outputs(11812) <= (inputs(19)) and not (inputs(206));
    layer0_outputs(11813) <= '1';
    layer0_outputs(11814) <= not(inputs(165));
    layer0_outputs(11815) <= (inputs(142)) xor (inputs(25));
    layer0_outputs(11816) <= not((inputs(155)) xor (inputs(246)));
    layer0_outputs(11817) <= (inputs(196)) xor (inputs(178));
    layer0_outputs(11818) <= (inputs(247)) and not (inputs(92));
    layer0_outputs(11819) <= not((inputs(167)) xor (inputs(131)));
    layer0_outputs(11820) <= not(inputs(84)) or (inputs(47));
    layer0_outputs(11821) <= not(inputs(252)) or (inputs(65));
    layer0_outputs(11822) <= inputs(9);
    layer0_outputs(11823) <= (inputs(2)) or (inputs(38));
    layer0_outputs(11824) <= inputs(215);
    layer0_outputs(11825) <= not((inputs(185)) xor (inputs(250)));
    layer0_outputs(11826) <= (inputs(125)) and not (inputs(221));
    layer0_outputs(11827) <= not(inputs(145));
    layer0_outputs(11828) <= not((inputs(141)) and (inputs(87)));
    layer0_outputs(11829) <= (inputs(189)) and (inputs(248));
    layer0_outputs(11830) <= (inputs(109)) and not (inputs(163));
    layer0_outputs(11831) <= not((inputs(74)) xor (inputs(58)));
    layer0_outputs(11832) <= not(inputs(82)) or (inputs(159));
    layer0_outputs(11833) <= (inputs(121)) and not (inputs(49));
    layer0_outputs(11834) <= (inputs(24)) xor (inputs(82));
    layer0_outputs(11835) <= inputs(8);
    layer0_outputs(11836) <= not(inputs(96));
    layer0_outputs(11837) <= not(inputs(125));
    layer0_outputs(11838) <= (inputs(210)) or (inputs(150));
    layer0_outputs(11839) <= not((inputs(33)) or (inputs(56)));
    layer0_outputs(11840) <= (inputs(148)) and not (inputs(32));
    layer0_outputs(11841) <= (inputs(254)) xor (inputs(206));
    layer0_outputs(11842) <= (inputs(3)) and not (inputs(63));
    layer0_outputs(11843) <= not(inputs(100));
    layer0_outputs(11844) <= (inputs(129)) or (inputs(182));
    layer0_outputs(11845) <= not(inputs(163));
    layer0_outputs(11846) <= (inputs(122)) and not (inputs(70));
    layer0_outputs(11847) <= not(inputs(150));
    layer0_outputs(11848) <= not(inputs(250)) or (inputs(125));
    layer0_outputs(11849) <= (inputs(189)) and (inputs(85));
    layer0_outputs(11850) <= (inputs(182)) and not (inputs(223));
    layer0_outputs(11851) <= not((inputs(148)) and (inputs(178)));
    layer0_outputs(11852) <= not((inputs(113)) or (inputs(216)));
    layer0_outputs(11853) <= (inputs(133)) and not (inputs(4));
    layer0_outputs(11854) <= not(inputs(56)) or (inputs(254));
    layer0_outputs(11855) <= (inputs(36)) or (inputs(150));
    layer0_outputs(11856) <= not((inputs(82)) xor (inputs(84)));
    layer0_outputs(11857) <= (inputs(147)) and not (inputs(3));
    layer0_outputs(11858) <= (inputs(23)) or (inputs(209));
    layer0_outputs(11859) <= (inputs(90)) and not (inputs(222));
    layer0_outputs(11860) <= not(inputs(93));
    layer0_outputs(11861) <= inputs(247);
    layer0_outputs(11862) <= (inputs(235)) or (inputs(228));
    layer0_outputs(11863) <= (inputs(209)) xor (inputs(195));
    layer0_outputs(11864) <= (inputs(29)) and not (inputs(230));
    layer0_outputs(11865) <= not(inputs(162));
    layer0_outputs(11866) <= (inputs(161)) xor (inputs(188));
    layer0_outputs(11867) <= (inputs(239)) or (inputs(113));
    layer0_outputs(11868) <= (inputs(237)) and (inputs(252));
    layer0_outputs(11869) <= not(inputs(117)) or (inputs(51));
    layer0_outputs(11870) <= (inputs(124)) xor (inputs(142));
    layer0_outputs(11871) <= (inputs(179)) and not (inputs(2));
    layer0_outputs(11872) <= (inputs(6)) and not (inputs(220));
    layer0_outputs(11873) <= (inputs(216)) or (inputs(222));
    layer0_outputs(11874) <= not(inputs(146)) or (inputs(69));
    layer0_outputs(11875) <= (inputs(135)) and not (inputs(14));
    layer0_outputs(11876) <= inputs(248);
    layer0_outputs(11877) <= (inputs(75)) and not (inputs(160));
    layer0_outputs(11878) <= not((inputs(50)) or (inputs(40)));
    layer0_outputs(11879) <= (inputs(37)) and not (inputs(50));
    layer0_outputs(11880) <= inputs(198);
    layer0_outputs(11881) <= (inputs(197)) xor (inputs(3));
    layer0_outputs(11882) <= (inputs(33)) xor (inputs(52));
    layer0_outputs(11883) <= (inputs(204)) and not (inputs(241));
    layer0_outputs(11884) <= (inputs(40)) and not (inputs(139));
    layer0_outputs(11885) <= not(inputs(164));
    layer0_outputs(11886) <= '0';
    layer0_outputs(11887) <= not((inputs(112)) xor (inputs(172)));
    layer0_outputs(11888) <= not(inputs(181));
    layer0_outputs(11889) <= (inputs(16)) or (inputs(176));
    layer0_outputs(11890) <= (inputs(112)) or (inputs(116));
    layer0_outputs(11891) <= inputs(192);
    layer0_outputs(11892) <= not(inputs(243));
    layer0_outputs(11893) <= (inputs(52)) or (inputs(56));
    layer0_outputs(11894) <= (inputs(73)) or (inputs(237));
    layer0_outputs(11895) <= (inputs(98)) or (inputs(155));
    layer0_outputs(11896) <= not((inputs(13)) xor (inputs(186)));
    layer0_outputs(11897) <= (inputs(190)) xor (inputs(98));
    layer0_outputs(11898) <= (inputs(83)) xor (inputs(111));
    layer0_outputs(11899) <= (inputs(255)) xor (inputs(15));
    layer0_outputs(11900) <= inputs(188);
    layer0_outputs(11901) <= not(inputs(7));
    layer0_outputs(11902) <= (inputs(156)) or (inputs(44));
    layer0_outputs(11903) <= not(inputs(9)) or (inputs(114));
    layer0_outputs(11904) <= (inputs(236)) xor (inputs(34));
    layer0_outputs(11905) <= not((inputs(138)) or (inputs(231)));
    layer0_outputs(11906) <= not(inputs(90)) or (inputs(226));
    layer0_outputs(11907) <= not((inputs(175)) or (inputs(95)));
    layer0_outputs(11908) <= (inputs(65)) or (inputs(149));
    layer0_outputs(11909) <= (inputs(148)) or (inputs(52));
    layer0_outputs(11910) <= (inputs(217)) and not (inputs(1));
    layer0_outputs(11911) <= (inputs(87)) or (inputs(205));
    layer0_outputs(11912) <= (inputs(187)) xor (inputs(250));
    layer0_outputs(11913) <= not(inputs(247)) or (inputs(88));
    layer0_outputs(11914) <= not(inputs(89));
    layer0_outputs(11915) <= (inputs(255)) and not (inputs(103));
    layer0_outputs(11916) <= not((inputs(167)) and (inputs(124)));
    layer0_outputs(11917) <= (inputs(71)) xor (inputs(25));
    layer0_outputs(11918) <= not((inputs(161)) or (inputs(178)));
    layer0_outputs(11919) <= not(inputs(88));
    layer0_outputs(11920) <= (inputs(139)) or (inputs(14));
    layer0_outputs(11921) <= not(inputs(51)) or (inputs(62));
    layer0_outputs(11922) <= not((inputs(124)) or (inputs(59)));
    layer0_outputs(11923) <= (inputs(210)) and not (inputs(20));
    layer0_outputs(11924) <= inputs(146);
    layer0_outputs(11925) <= (inputs(10)) xor (inputs(156));
    layer0_outputs(11926) <= not((inputs(165)) or (inputs(14)));
    layer0_outputs(11927) <= (inputs(56)) xor (inputs(57));
    layer0_outputs(11928) <= (inputs(43)) and not (inputs(18));
    layer0_outputs(11929) <= not(inputs(246)) or (inputs(157));
    layer0_outputs(11930) <= (inputs(212)) xor (inputs(183));
    layer0_outputs(11931) <= not((inputs(120)) or (inputs(33)));
    layer0_outputs(11932) <= not((inputs(128)) or (inputs(95)));
    layer0_outputs(11933) <= inputs(71);
    layer0_outputs(11934) <= not(inputs(6));
    layer0_outputs(11935) <= not((inputs(24)) or (inputs(7)));
    layer0_outputs(11936) <= (inputs(110)) xor (inputs(27));
    layer0_outputs(11937) <= (inputs(29)) and (inputs(101));
    layer0_outputs(11938) <= (inputs(74)) and not (inputs(205));
    layer0_outputs(11939) <= not((inputs(187)) or (inputs(130)));
    layer0_outputs(11940) <= (inputs(18)) xor (inputs(80));
    layer0_outputs(11941) <= inputs(67);
    layer0_outputs(11942) <= inputs(230);
    layer0_outputs(11943) <= not(inputs(179));
    layer0_outputs(11944) <= not((inputs(170)) xor (inputs(141)));
    layer0_outputs(11945) <= not((inputs(57)) or (inputs(77)));
    layer0_outputs(11946) <= not((inputs(199)) or (inputs(234)));
    layer0_outputs(11947) <= not(inputs(10));
    layer0_outputs(11948) <= not(inputs(127)) or (inputs(187));
    layer0_outputs(11949) <= not((inputs(24)) or (inputs(23)));
    layer0_outputs(11950) <= (inputs(115)) and not (inputs(62));
    layer0_outputs(11951) <= inputs(168);
    layer0_outputs(11952) <= (inputs(39)) xor (inputs(123));
    layer0_outputs(11953) <= inputs(82);
    layer0_outputs(11954) <= not((inputs(242)) xor (inputs(36)));
    layer0_outputs(11955) <= (inputs(17)) xor (inputs(101));
    layer0_outputs(11956) <= (inputs(180)) xor (inputs(174));
    layer0_outputs(11957) <= (inputs(230)) xor (inputs(4));
    layer0_outputs(11958) <= not(inputs(94));
    layer0_outputs(11959) <= not((inputs(184)) xor (inputs(200)));
    layer0_outputs(11960) <= (inputs(35)) xor (inputs(67));
    layer0_outputs(11961) <= (inputs(234)) xor (inputs(163));
    layer0_outputs(11962) <= (inputs(78)) and not (inputs(0));
    layer0_outputs(11963) <= not((inputs(223)) or (inputs(216)));
    layer0_outputs(11964) <= (inputs(27)) xor (inputs(100));
    layer0_outputs(11965) <= not((inputs(190)) xor (inputs(166)));
    layer0_outputs(11966) <= not((inputs(209)) xor (inputs(4)));
    layer0_outputs(11967) <= not((inputs(46)) or (inputs(26)));
    layer0_outputs(11968) <= inputs(11);
    layer0_outputs(11969) <= inputs(48);
    layer0_outputs(11970) <= (inputs(89)) xor (inputs(164));
    layer0_outputs(11971) <= not((inputs(99)) or (inputs(12)));
    layer0_outputs(11972) <= inputs(152);
    layer0_outputs(11973) <= not(inputs(183)) or (inputs(175));
    layer0_outputs(11974) <= not(inputs(77));
    layer0_outputs(11975) <= (inputs(2)) and (inputs(37));
    layer0_outputs(11976) <= not((inputs(189)) xor (inputs(240)));
    layer0_outputs(11977) <= not(inputs(245)) or (inputs(68));
    layer0_outputs(11978) <= not(inputs(216)) or (inputs(189));
    layer0_outputs(11979) <= inputs(103);
    layer0_outputs(11980) <= not((inputs(30)) or (inputs(81)));
    layer0_outputs(11981) <= not(inputs(154)) or (inputs(62));
    layer0_outputs(11982) <= not(inputs(162));
    layer0_outputs(11983) <= (inputs(85)) and not (inputs(236));
    layer0_outputs(11984) <= not((inputs(133)) xor (inputs(139)));
    layer0_outputs(11985) <= (inputs(168)) xor (inputs(138));
    layer0_outputs(11986) <= not(inputs(184));
    layer0_outputs(11987) <= (inputs(231)) and not (inputs(124));
    layer0_outputs(11988) <= (inputs(128)) xor (inputs(101));
    layer0_outputs(11989) <= not(inputs(213)) or (inputs(4));
    layer0_outputs(11990) <= (inputs(62)) or (inputs(6));
    layer0_outputs(11991) <= not(inputs(5));
    layer0_outputs(11992) <= not((inputs(133)) or (inputs(118)));
    layer0_outputs(11993) <= (inputs(89)) xor (inputs(167));
    layer0_outputs(11994) <= (inputs(166)) and (inputs(136));
    layer0_outputs(11995) <= inputs(221);
    layer0_outputs(11996) <= not(inputs(164)) or (inputs(177));
    layer0_outputs(11997) <= not(inputs(37)) or (inputs(103));
    layer0_outputs(11998) <= not(inputs(65));
    layer0_outputs(11999) <= inputs(5);
    layer0_outputs(12000) <= (inputs(157)) and (inputs(207));
    layer0_outputs(12001) <= not((inputs(214)) or (inputs(193)));
    layer0_outputs(12002) <= inputs(120);
    layer0_outputs(12003) <= (inputs(176)) or (inputs(191));
    layer0_outputs(12004) <= not((inputs(96)) or (inputs(161)));
    layer0_outputs(12005) <= inputs(152);
    layer0_outputs(12006) <= (inputs(101)) xor (inputs(72));
    layer0_outputs(12007) <= (inputs(139)) or (inputs(30));
    layer0_outputs(12008) <= inputs(106);
    layer0_outputs(12009) <= not((inputs(55)) xor (inputs(125)));
    layer0_outputs(12010) <= not(inputs(146));
    layer0_outputs(12011) <= not((inputs(80)) xor (inputs(216)));
    layer0_outputs(12012) <= (inputs(221)) and not (inputs(33));
    layer0_outputs(12013) <= not((inputs(44)) xor (inputs(227)));
    layer0_outputs(12014) <= not(inputs(122));
    layer0_outputs(12015) <= (inputs(27)) and not (inputs(159));
    layer0_outputs(12016) <= (inputs(207)) and not (inputs(254));
    layer0_outputs(12017) <= inputs(104);
    layer0_outputs(12018) <= not((inputs(108)) or (inputs(30)));
    layer0_outputs(12019) <= (inputs(121)) xor (inputs(179));
    layer0_outputs(12020) <= not(inputs(38));
    layer0_outputs(12021) <= not(inputs(87));
    layer0_outputs(12022) <= (inputs(177)) xor (inputs(192));
    layer0_outputs(12023) <= not((inputs(252)) or (inputs(169)));
    layer0_outputs(12024) <= inputs(152);
    layer0_outputs(12025) <= (inputs(240)) or (inputs(244));
    layer0_outputs(12026) <= (inputs(19)) xor (inputs(204));
    layer0_outputs(12027) <= not((inputs(243)) or (inputs(247)));
    layer0_outputs(12028) <= not(inputs(34)) or (inputs(84));
    layer0_outputs(12029) <= not((inputs(110)) or (inputs(223)));
    layer0_outputs(12030) <= (inputs(226)) and not (inputs(187));
    layer0_outputs(12031) <= '0';
    layer0_outputs(12032) <= (inputs(200)) or (inputs(160));
    layer0_outputs(12033) <= (inputs(44)) and (inputs(61));
    layer0_outputs(12034) <= not(inputs(167)) or (inputs(201));
    layer0_outputs(12035) <= not((inputs(207)) xor (inputs(40)));
    layer0_outputs(12036) <= inputs(202);
    layer0_outputs(12037) <= not(inputs(104)) or (inputs(229));
    layer0_outputs(12038) <= not(inputs(193));
    layer0_outputs(12039) <= inputs(233);
    layer0_outputs(12040) <= not(inputs(92)) or (inputs(160));
    layer0_outputs(12041) <= not(inputs(195));
    layer0_outputs(12042) <= (inputs(87)) xor (inputs(224));
    layer0_outputs(12043) <= not(inputs(129));
    layer0_outputs(12044) <= not(inputs(219)) or (inputs(3));
    layer0_outputs(12045) <= inputs(15);
    layer0_outputs(12046) <= not((inputs(247)) or (inputs(42)));
    layer0_outputs(12047) <= not(inputs(74));
    layer0_outputs(12048) <= not(inputs(89));
    layer0_outputs(12049) <= not((inputs(191)) xor (inputs(222)));
    layer0_outputs(12050) <= (inputs(205)) and not (inputs(142));
    layer0_outputs(12051) <= (inputs(75)) xor (inputs(109));
    layer0_outputs(12052) <= (inputs(223)) or (inputs(251));
    layer0_outputs(12053) <= inputs(53);
    layer0_outputs(12054) <= inputs(30);
    layer0_outputs(12055) <= not(inputs(196));
    layer0_outputs(12056) <= not(inputs(24)) or (inputs(146));
    layer0_outputs(12057) <= (inputs(228)) xor (inputs(134));
    layer0_outputs(12058) <= not((inputs(110)) or (inputs(13)));
    layer0_outputs(12059) <= not(inputs(232)) or (inputs(178));
    layer0_outputs(12060) <= not(inputs(226));
    layer0_outputs(12061) <= (inputs(224)) or (inputs(211));
    layer0_outputs(12062) <= not((inputs(211)) and (inputs(70)));
    layer0_outputs(12063) <= not(inputs(13));
    layer0_outputs(12064) <= not((inputs(200)) or (inputs(83)));
    layer0_outputs(12065) <= not(inputs(153));
    layer0_outputs(12066) <= (inputs(117)) xor (inputs(173));
    layer0_outputs(12067) <= (inputs(115)) and not (inputs(239));
    layer0_outputs(12068) <= not(inputs(162));
    layer0_outputs(12069) <= not(inputs(166)) or (inputs(208));
    layer0_outputs(12070) <= (inputs(231)) xor (inputs(224));
    layer0_outputs(12071) <= (inputs(42)) and not (inputs(165));
    layer0_outputs(12072) <= (inputs(144)) and not (inputs(136));
    layer0_outputs(12073) <= inputs(172);
    layer0_outputs(12074) <= inputs(214);
    layer0_outputs(12075) <= inputs(147);
    layer0_outputs(12076) <= (inputs(235)) xor (inputs(184));
    layer0_outputs(12077) <= (inputs(186)) xor (inputs(142));
    layer0_outputs(12078) <= inputs(148);
    layer0_outputs(12079) <= (inputs(32)) and not (inputs(127));
    layer0_outputs(12080) <= not((inputs(146)) xor (inputs(182)));
    layer0_outputs(12081) <= (inputs(86)) or (inputs(181));
    layer0_outputs(12082) <= not(inputs(249));
    layer0_outputs(12083) <= inputs(134);
    layer0_outputs(12084) <= not((inputs(81)) or (inputs(117)));
    layer0_outputs(12085) <= (inputs(109)) or (inputs(183));
    layer0_outputs(12086) <= inputs(71);
    layer0_outputs(12087) <= not((inputs(193)) xor (inputs(8)));
    layer0_outputs(12088) <= not(inputs(22)) or (inputs(160));
    layer0_outputs(12089) <= (inputs(40)) and not (inputs(210));
    layer0_outputs(12090) <= (inputs(59)) and not (inputs(4));
    layer0_outputs(12091) <= (inputs(34)) xor (inputs(7));
    layer0_outputs(12092) <= not(inputs(44));
    layer0_outputs(12093) <= not(inputs(99));
    layer0_outputs(12094) <= inputs(145);
    layer0_outputs(12095) <= not((inputs(178)) and (inputs(83)));
    layer0_outputs(12096) <= (inputs(74)) or (inputs(143));
    layer0_outputs(12097) <= not((inputs(170)) or (inputs(16)));
    layer0_outputs(12098) <= inputs(180);
    layer0_outputs(12099) <= (inputs(241)) or (inputs(107));
    layer0_outputs(12100) <= (inputs(10)) xor (inputs(59));
    layer0_outputs(12101) <= inputs(178);
    layer0_outputs(12102) <= not(inputs(88));
    layer0_outputs(12103) <= (inputs(150)) and not (inputs(5));
    layer0_outputs(12104) <= (inputs(18)) xor (inputs(100));
    layer0_outputs(12105) <= not(inputs(15));
    layer0_outputs(12106) <= (inputs(170)) or (inputs(199));
    layer0_outputs(12107) <= (inputs(25)) and not (inputs(237));
    layer0_outputs(12108) <= (inputs(194)) or (inputs(175));
    layer0_outputs(12109) <= (inputs(178)) xor (inputs(142));
    layer0_outputs(12110) <= (inputs(209)) and not (inputs(10));
    layer0_outputs(12111) <= not((inputs(161)) xor (inputs(182)));
    layer0_outputs(12112) <= not((inputs(11)) xor (inputs(96)));
    layer0_outputs(12113) <= not(inputs(176));
    layer0_outputs(12114) <= not((inputs(59)) or (inputs(3)));
    layer0_outputs(12115) <= not((inputs(115)) or (inputs(56)));
    layer0_outputs(12116) <= inputs(212);
    layer0_outputs(12117) <= not(inputs(253));
    layer0_outputs(12118) <= not(inputs(218)) or (inputs(76));
    layer0_outputs(12119) <= not((inputs(244)) or (inputs(188)));
    layer0_outputs(12120) <= (inputs(165)) or (inputs(206));
    layer0_outputs(12121) <= (inputs(245)) and not (inputs(47));
    layer0_outputs(12122) <= (inputs(215)) and not (inputs(120));
    layer0_outputs(12123) <= (inputs(37)) xor (inputs(70));
    layer0_outputs(12124) <= not((inputs(33)) xor (inputs(118)));
    layer0_outputs(12125) <= not(inputs(224));
    layer0_outputs(12126) <= not((inputs(61)) xor (inputs(156)));
    layer0_outputs(12127) <= (inputs(217)) and not (inputs(76));
    layer0_outputs(12128) <= not((inputs(18)) or (inputs(94)));
    layer0_outputs(12129) <= (inputs(12)) xor (inputs(43));
    layer0_outputs(12130) <= (inputs(240)) or (inputs(57));
    layer0_outputs(12131) <= not(inputs(221));
    layer0_outputs(12132) <= (inputs(232)) or (inputs(113));
    layer0_outputs(12133) <= not(inputs(95));
    layer0_outputs(12134) <= inputs(154);
    layer0_outputs(12135) <= (inputs(80)) and not (inputs(17));
    layer0_outputs(12136) <= inputs(229);
    layer0_outputs(12137) <= not((inputs(211)) or (inputs(232)));
    layer0_outputs(12138) <= (inputs(11)) and (inputs(253));
    layer0_outputs(12139) <= '1';
    layer0_outputs(12140) <= inputs(76);
    layer0_outputs(12141) <= (inputs(190)) xor (inputs(185));
    layer0_outputs(12142) <= not(inputs(142));
    layer0_outputs(12143) <= not((inputs(207)) xor (inputs(145)));
    layer0_outputs(12144) <= not((inputs(223)) or (inputs(172)));
    layer0_outputs(12145) <= not((inputs(64)) or (inputs(151)));
    layer0_outputs(12146) <= not(inputs(233)) or (inputs(238));
    layer0_outputs(12147) <= not((inputs(229)) and (inputs(165)));
    layer0_outputs(12148) <= not(inputs(177));
    layer0_outputs(12149) <= (inputs(7)) xor (inputs(51));
    layer0_outputs(12150) <= (inputs(166)) and not (inputs(245));
    layer0_outputs(12151) <= inputs(128);
    layer0_outputs(12152) <= not((inputs(15)) or (inputs(1)));
    layer0_outputs(12153) <= not(inputs(111));
    layer0_outputs(12154) <= not(inputs(159));
    layer0_outputs(12155) <= (inputs(121)) or (inputs(209));
    layer0_outputs(12156) <= (inputs(91)) xor (inputs(89));
    layer0_outputs(12157) <= (inputs(200)) or (inputs(251));
    layer0_outputs(12158) <= not(inputs(57));
    layer0_outputs(12159) <= inputs(90);
    layer0_outputs(12160) <= (inputs(140)) and not (inputs(243));
    layer0_outputs(12161) <= inputs(142);
    layer0_outputs(12162) <= (inputs(119)) xor (inputs(91));
    layer0_outputs(12163) <= not(inputs(194));
    layer0_outputs(12164) <= (inputs(8)) xor (inputs(198));
    layer0_outputs(12165) <= inputs(147);
    layer0_outputs(12166) <= not(inputs(13));
    layer0_outputs(12167) <= not((inputs(142)) xor (inputs(12)));
    layer0_outputs(12168) <= not(inputs(116));
    layer0_outputs(12169) <= not((inputs(243)) xor (inputs(51)));
    layer0_outputs(12170) <= not(inputs(107));
    layer0_outputs(12171) <= not(inputs(164)) or (inputs(17));
    layer0_outputs(12172) <= inputs(38);
    layer0_outputs(12173) <= inputs(122);
    layer0_outputs(12174) <= (inputs(3)) and not (inputs(81));
    layer0_outputs(12175) <= (inputs(14)) xor (inputs(247));
    layer0_outputs(12176) <= (inputs(40)) and not (inputs(55));
    layer0_outputs(12177) <= (inputs(191)) xor (inputs(25));
    layer0_outputs(12178) <= (inputs(144)) or (inputs(99));
    layer0_outputs(12179) <= not((inputs(78)) or (inputs(95)));
    layer0_outputs(12180) <= (inputs(70)) and not (inputs(157));
    layer0_outputs(12181) <= not((inputs(223)) xor (inputs(176)));
    layer0_outputs(12182) <= not(inputs(24));
    layer0_outputs(12183) <= (inputs(5)) xor (inputs(189));
    layer0_outputs(12184) <= not(inputs(84));
    layer0_outputs(12185) <= (inputs(168)) and not (inputs(35));
    layer0_outputs(12186) <= not((inputs(85)) or (inputs(163)));
    layer0_outputs(12187) <= not((inputs(123)) or (inputs(172)));
    layer0_outputs(12188) <= not((inputs(190)) xor (inputs(51)));
    layer0_outputs(12189) <= inputs(219);
    layer0_outputs(12190) <= (inputs(144)) and not (inputs(26));
    layer0_outputs(12191) <= inputs(195);
    layer0_outputs(12192) <= inputs(82);
    layer0_outputs(12193) <= not((inputs(68)) xor (inputs(131)));
    layer0_outputs(12194) <= (inputs(167)) xor (inputs(160));
    layer0_outputs(12195) <= (inputs(136)) or (inputs(106));
    layer0_outputs(12196) <= not((inputs(113)) and (inputs(14)));
    layer0_outputs(12197) <= (inputs(55)) xor (inputs(216));
    layer0_outputs(12198) <= (inputs(12)) and not (inputs(140));
    layer0_outputs(12199) <= not((inputs(84)) or (inputs(190)));
    layer0_outputs(12200) <= not(inputs(116));
    layer0_outputs(12201) <= not(inputs(104));
    layer0_outputs(12202) <= not((inputs(246)) xor (inputs(41)));
    layer0_outputs(12203) <= inputs(151);
    layer0_outputs(12204) <= not((inputs(40)) or (inputs(208)));
    layer0_outputs(12205) <= not((inputs(13)) xor (inputs(88)));
    layer0_outputs(12206) <= inputs(203);
    layer0_outputs(12207) <= not((inputs(152)) or (inputs(208)));
    layer0_outputs(12208) <= not((inputs(99)) xor (inputs(47)));
    layer0_outputs(12209) <= (inputs(129)) and not (inputs(249));
    layer0_outputs(12210) <= not(inputs(9));
    layer0_outputs(12211) <= not(inputs(160));
    layer0_outputs(12212) <= inputs(93);
    layer0_outputs(12213) <= not(inputs(27)) or (inputs(174));
    layer0_outputs(12214) <= inputs(24);
    layer0_outputs(12215) <= not((inputs(201)) xor (inputs(117)));
    layer0_outputs(12216) <= not((inputs(210)) or (inputs(237)));
    layer0_outputs(12217) <= (inputs(25)) or (inputs(250));
    layer0_outputs(12218) <= not(inputs(42));
    layer0_outputs(12219) <= not((inputs(95)) xor (inputs(91)));
    layer0_outputs(12220) <= not(inputs(146));
    layer0_outputs(12221) <= not((inputs(141)) or (inputs(54)));
    layer0_outputs(12222) <= inputs(166);
    layer0_outputs(12223) <= not((inputs(99)) or (inputs(198)));
    layer0_outputs(12224) <= inputs(139);
    layer0_outputs(12225) <= inputs(219);
    layer0_outputs(12226) <= not((inputs(87)) xor (inputs(91)));
    layer0_outputs(12227) <= not(inputs(18));
    layer0_outputs(12228) <= not(inputs(73));
    layer0_outputs(12229) <= not(inputs(167)) or (inputs(255));
    layer0_outputs(12230) <= (inputs(32)) or (inputs(24));
    layer0_outputs(12231) <= (inputs(244)) and (inputs(205));
    layer0_outputs(12232) <= (inputs(105)) and not (inputs(196));
    layer0_outputs(12233) <= not((inputs(163)) xor (inputs(147)));
    layer0_outputs(12234) <= '1';
    layer0_outputs(12235) <= not((inputs(147)) xor (inputs(234)));
    layer0_outputs(12236) <= not((inputs(198)) xor (inputs(170)));
    layer0_outputs(12237) <= (inputs(238)) or (inputs(222));
    layer0_outputs(12238) <= not(inputs(75)) or (inputs(10));
    layer0_outputs(12239) <= not(inputs(89)) or (inputs(81));
    layer0_outputs(12240) <= (inputs(6)) and not (inputs(52));
    layer0_outputs(12241) <= (inputs(198)) and not (inputs(239));
    layer0_outputs(12242) <= not((inputs(245)) xor (inputs(167)));
    layer0_outputs(12243) <= not((inputs(189)) xor (inputs(106)));
    layer0_outputs(12244) <= inputs(218);
    layer0_outputs(12245) <= not((inputs(165)) or (inputs(31)));
    layer0_outputs(12246) <= '0';
    layer0_outputs(12247) <= inputs(204);
    layer0_outputs(12248) <= inputs(124);
    layer0_outputs(12249) <= (inputs(241)) xor (inputs(182));
    layer0_outputs(12250) <= not(inputs(88)) or (inputs(144));
    layer0_outputs(12251) <= not(inputs(125)) or (inputs(73));
    layer0_outputs(12252) <= not(inputs(40));
    layer0_outputs(12253) <= (inputs(232)) xor (inputs(169));
    layer0_outputs(12254) <= not(inputs(99));
    layer0_outputs(12255) <= not(inputs(11));
    layer0_outputs(12256) <= not((inputs(53)) xor (inputs(73)));
    layer0_outputs(12257) <= (inputs(62)) or (inputs(224));
    layer0_outputs(12258) <= not(inputs(194));
    layer0_outputs(12259) <= inputs(179);
    layer0_outputs(12260) <= (inputs(58)) xor (inputs(149));
    layer0_outputs(12261) <= not(inputs(100));
    layer0_outputs(12262) <= not((inputs(160)) xor (inputs(6)));
    layer0_outputs(12263) <= (inputs(207)) and not (inputs(62));
    layer0_outputs(12264) <= inputs(36);
    layer0_outputs(12265) <= not((inputs(179)) xor (inputs(224)));
    layer0_outputs(12266) <= not(inputs(135)) or (inputs(252));
    layer0_outputs(12267) <= (inputs(156)) and not (inputs(42));
    layer0_outputs(12268) <= inputs(183);
    layer0_outputs(12269) <= not(inputs(110));
    layer0_outputs(12270) <= not((inputs(127)) or (inputs(237)));
    layer0_outputs(12271) <= not(inputs(130));
    layer0_outputs(12272) <= not((inputs(14)) or (inputs(201)));
    layer0_outputs(12273) <= (inputs(129)) or (inputs(61));
    layer0_outputs(12274) <= not(inputs(116));
    layer0_outputs(12275) <= not(inputs(222));
    layer0_outputs(12276) <= inputs(43);
    layer0_outputs(12277) <= not((inputs(230)) or (inputs(192)));
    layer0_outputs(12278) <= not(inputs(22));
    layer0_outputs(12279) <= inputs(125);
    layer0_outputs(12280) <= (inputs(39)) and not (inputs(237));
    layer0_outputs(12281) <= (inputs(147)) or (inputs(94));
    layer0_outputs(12282) <= (inputs(236)) or (inputs(64));
    layer0_outputs(12283) <= (inputs(97)) and not (inputs(56));
    layer0_outputs(12284) <= not((inputs(95)) or (inputs(52)));
    layer0_outputs(12285) <= (inputs(105)) or (inputs(20));
    layer0_outputs(12286) <= not((inputs(221)) xor (inputs(208)));
    layer0_outputs(12287) <= inputs(213);
    layer0_outputs(12288) <= '1';
    layer0_outputs(12289) <= inputs(179);
    layer0_outputs(12290) <= inputs(202);
    layer0_outputs(12291) <= not((inputs(165)) xor (inputs(162)));
    layer0_outputs(12292) <= not(inputs(73));
    layer0_outputs(12293) <= not(inputs(196)) or (inputs(254));
    layer0_outputs(12294) <= (inputs(207)) xor (inputs(116));
    layer0_outputs(12295) <= (inputs(243)) xor (inputs(206));
    layer0_outputs(12296) <= not((inputs(87)) or (inputs(200)));
    layer0_outputs(12297) <= inputs(181);
    layer0_outputs(12298) <= not((inputs(212)) and (inputs(92)));
    layer0_outputs(12299) <= not((inputs(202)) xor (inputs(4)));
    layer0_outputs(12300) <= not((inputs(160)) xor (inputs(132)));
    layer0_outputs(12301) <= not(inputs(209));
    layer0_outputs(12302) <= (inputs(192)) xor (inputs(167));
    layer0_outputs(12303) <= not(inputs(222));
    layer0_outputs(12304) <= inputs(77);
    layer0_outputs(12305) <= not(inputs(128)) or (inputs(72));
    layer0_outputs(12306) <= inputs(104);
    layer0_outputs(12307) <= not((inputs(23)) or (inputs(219)));
    layer0_outputs(12308) <= (inputs(130)) or (inputs(85));
    layer0_outputs(12309) <= (inputs(171)) xor (inputs(217));
    layer0_outputs(12310) <= not(inputs(243)) or (inputs(95));
    layer0_outputs(12311) <= inputs(249);
    layer0_outputs(12312) <= not(inputs(130));
    layer0_outputs(12313) <= not(inputs(103));
    layer0_outputs(12314) <= not((inputs(63)) or (inputs(69)));
    layer0_outputs(12315) <= (inputs(168)) and not (inputs(79));
    layer0_outputs(12316) <= not((inputs(0)) xor (inputs(35)));
    layer0_outputs(12317) <= (inputs(67)) xor (inputs(235));
    layer0_outputs(12318) <= not(inputs(221));
    layer0_outputs(12319) <= (inputs(144)) xor (inputs(58));
    layer0_outputs(12320) <= inputs(167);
    layer0_outputs(12321) <= inputs(85);
    layer0_outputs(12322) <= (inputs(130)) and not (inputs(72));
    layer0_outputs(12323) <= not(inputs(29));
    layer0_outputs(12324) <= inputs(114);
    layer0_outputs(12325) <= (inputs(221)) or (inputs(95));
    layer0_outputs(12326) <= inputs(176);
    layer0_outputs(12327) <= (inputs(133)) xor (inputs(93));
    layer0_outputs(12328) <= not((inputs(74)) xor (inputs(35)));
    layer0_outputs(12329) <= not((inputs(28)) xor (inputs(72)));
    layer0_outputs(12330) <= not((inputs(204)) or (inputs(223)));
    layer0_outputs(12331) <= (inputs(34)) xor (inputs(255));
    layer0_outputs(12332) <= (inputs(77)) and not (inputs(226));
    layer0_outputs(12333) <= not((inputs(0)) or (inputs(207)));
    layer0_outputs(12334) <= not(inputs(197)) or (inputs(182));
    layer0_outputs(12335) <= not(inputs(77));
    layer0_outputs(12336) <= not((inputs(130)) or (inputs(13)));
    layer0_outputs(12337) <= not(inputs(137)) or (inputs(94));
    layer0_outputs(12338) <= not(inputs(6));
    layer0_outputs(12339) <= inputs(56);
    layer0_outputs(12340) <= (inputs(251)) xor (inputs(202));
    layer0_outputs(12341) <= inputs(182);
    layer0_outputs(12342) <= not((inputs(47)) or (inputs(228)));
    layer0_outputs(12343) <= (inputs(135)) and not (inputs(109));
    layer0_outputs(12344) <= (inputs(122)) or (inputs(214));
    layer0_outputs(12345) <= not(inputs(167));
    layer0_outputs(12346) <= not((inputs(149)) xor (inputs(246)));
    layer0_outputs(12347) <= not(inputs(200)) or (inputs(133));
    layer0_outputs(12348) <= (inputs(66)) and not (inputs(222));
    layer0_outputs(12349) <= not((inputs(182)) xor (inputs(217)));
    layer0_outputs(12350) <= inputs(55);
    layer0_outputs(12351) <= (inputs(132)) and not (inputs(244));
    layer0_outputs(12352) <= not(inputs(234));
    layer0_outputs(12353) <= not((inputs(19)) xor (inputs(194)));
    layer0_outputs(12354) <= (inputs(237)) or (inputs(229));
    layer0_outputs(12355) <= (inputs(181)) or (inputs(188));
    layer0_outputs(12356) <= inputs(7);
    layer0_outputs(12357) <= (inputs(180)) or (inputs(202));
    layer0_outputs(12358) <= not(inputs(218));
    layer0_outputs(12359) <= (inputs(211)) and not (inputs(12));
    layer0_outputs(12360) <= (inputs(172)) xor (inputs(151));
    layer0_outputs(12361) <= not(inputs(6));
    layer0_outputs(12362) <= (inputs(223)) and (inputs(33));
    layer0_outputs(12363) <= (inputs(94)) xor (inputs(35));
    layer0_outputs(12364) <= not(inputs(237));
    layer0_outputs(12365) <= not((inputs(54)) xor (inputs(52)));
    layer0_outputs(12366) <= (inputs(238)) or (inputs(79));
    layer0_outputs(12367) <= not((inputs(224)) xor (inputs(136)));
    layer0_outputs(12368) <= not(inputs(32));
    layer0_outputs(12369) <= (inputs(176)) or (inputs(240));
    layer0_outputs(12370) <= (inputs(148)) and not (inputs(81));
    layer0_outputs(12371) <= not(inputs(82)) or (inputs(161));
    layer0_outputs(12372) <= (inputs(226)) and (inputs(14));
    layer0_outputs(12373) <= inputs(110);
    layer0_outputs(12374) <= (inputs(146)) and not (inputs(238));
    layer0_outputs(12375) <= not(inputs(21)) or (inputs(240));
    layer0_outputs(12376) <= inputs(236);
    layer0_outputs(12377) <= (inputs(199)) or (inputs(11));
    layer0_outputs(12378) <= not(inputs(244)) or (inputs(125));
    layer0_outputs(12379) <= (inputs(45)) xor (inputs(190));
    layer0_outputs(12380) <= not((inputs(199)) or (inputs(180)));
    layer0_outputs(12381) <= not(inputs(105)) or (inputs(173));
    layer0_outputs(12382) <= (inputs(23)) and not (inputs(30));
    layer0_outputs(12383) <= (inputs(131)) xor (inputs(67));
    layer0_outputs(12384) <= not(inputs(224));
    layer0_outputs(12385) <= not(inputs(36)) or (inputs(194));
    layer0_outputs(12386) <= inputs(22);
    layer0_outputs(12387) <= not(inputs(217)) or (inputs(16));
    layer0_outputs(12388) <= (inputs(195)) xor (inputs(12));
    layer0_outputs(12389) <= inputs(95);
    layer0_outputs(12390) <= inputs(120);
    layer0_outputs(12391) <= not(inputs(58));
    layer0_outputs(12392) <= inputs(37);
    layer0_outputs(12393) <= (inputs(169)) or (inputs(124));
    layer0_outputs(12394) <= inputs(228);
    layer0_outputs(12395) <= (inputs(105)) and (inputs(28));
    layer0_outputs(12396) <= not(inputs(195));
    layer0_outputs(12397) <= inputs(101);
    layer0_outputs(12398) <= (inputs(99)) xor (inputs(55));
    layer0_outputs(12399) <= inputs(150);
    layer0_outputs(12400) <= not((inputs(199)) and (inputs(152)));
    layer0_outputs(12401) <= (inputs(22)) and not (inputs(42));
    layer0_outputs(12402) <= not(inputs(94)) or (inputs(254));
    layer0_outputs(12403) <= not((inputs(190)) or (inputs(18)));
    layer0_outputs(12404) <= not(inputs(138));
    layer0_outputs(12405) <= not(inputs(71));
    layer0_outputs(12406) <= inputs(73);
    layer0_outputs(12407) <= (inputs(96)) or (inputs(171));
    layer0_outputs(12408) <= inputs(127);
    layer0_outputs(12409) <= not(inputs(87));
    layer0_outputs(12410) <= not(inputs(64)) or (inputs(54));
    layer0_outputs(12411) <= not(inputs(196));
    layer0_outputs(12412) <= not((inputs(145)) or (inputs(19)));
    layer0_outputs(12413) <= not((inputs(197)) or (inputs(65)));
    layer0_outputs(12414) <= not(inputs(250));
    layer0_outputs(12415) <= (inputs(135)) and not (inputs(85));
    layer0_outputs(12416) <= not((inputs(93)) xor (inputs(186)));
    layer0_outputs(12417) <= not((inputs(158)) or (inputs(162)));
    layer0_outputs(12418) <= inputs(116);
    layer0_outputs(12419) <= (inputs(102)) or (inputs(40));
    layer0_outputs(12420) <= not(inputs(174)) or (inputs(255));
    layer0_outputs(12421) <= (inputs(169)) and not (inputs(112));
    layer0_outputs(12422) <= not(inputs(234));
    layer0_outputs(12423) <= not((inputs(76)) or (inputs(142)));
    layer0_outputs(12424) <= inputs(170);
    layer0_outputs(12425) <= inputs(225);
    layer0_outputs(12426) <= (inputs(60)) and not (inputs(136));
    layer0_outputs(12427) <= inputs(164);
    layer0_outputs(12428) <= (inputs(54)) xor (inputs(57));
    layer0_outputs(12429) <= inputs(30);
    layer0_outputs(12430) <= (inputs(139)) xor (inputs(115));
    layer0_outputs(12431) <= inputs(133);
    layer0_outputs(12432) <= inputs(22);
    layer0_outputs(12433) <= not((inputs(104)) or (inputs(111)));
    layer0_outputs(12434) <= not((inputs(90)) xor (inputs(34)));
    layer0_outputs(12435) <= inputs(84);
    layer0_outputs(12436) <= not((inputs(169)) or (inputs(200)));
    layer0_outputs(12437) <= not(inputs(201)) or (inputs(96));
    layer0_outputs(12438) <= inputs(35);
    layer0_outputs(12439) <= (inputs(238)) xor (inputs(101));
    layer0_outputs(12440) <= not((inputs(106)) or (inputs(64)));
    layer0_outputs(12441) <= (inputs(147)) xor (inputs(158));
    layer0_outputs(12442) <= (inputs(60)) or (inputs(66));
    layer0_outputs(12443) <= not(inputs(139));
    layer0_outputs(12444) <= not((inputs(185)) xor (inputs(177)));
    layer0_outputs(12445) <= (inputs(173)) xor (inputs(105));
    layer0_outputs(12446) <= (inputs(68)) or (inputs(21));
    layer0_outputs(12447) <= (inputs(219)) xor (inputs(255));
    layer0_outputs(12448) <= (inputs(140)) and (inputs(165));
    layer0_outputs(12449) <= not(inputs(226)) or (inputs(150));
    layer0_outputs(12450) <= not(inputs(60));
    layer0_outputs(12451) <= not((inputs(66)) xor (inputs(242)));
    layer0_outputs(12452) <= not((inputs(13)) or (inputs(125)));
    layer0_outputs(12453) <= inputs(197);
    layer0_outputs(12454) <= (inputs(164)) and not (inputs(31));
    layer0_outputs(12455) <= not((inputs(35)) and (inputs(36)));
    layer0_outputs(12456) <= (inputs(159)) and not (inputs(172));
    layer0_outputs(12457) <= inputs(9);
    layer0_outputs(12458) <= (inputs(112)) and not (inputs(84));
    layer0_outputs(12459) <= (inputs(97)) xor (inputs(254));
    layer0_outputs(12460) <= not((inputs(24)) xor (inputs(86)));
    layer0_outputs(12461) <= not(inputs(122)) or (inputs(190));
    layer0_outputs(12462) <= '1';
    layer0_outputs(12463) <= inputs(129);
    layer0_outputs(12464) <= (inputs(55)) or (inputs(109));
    layer0_outputs(12465) <= (inputs(253)) and not (inputs(253));
    layer0_outputs(12466) <= not((inputs(163)) xor (inputs(246)));
    layer0_outputs(12467) <= inputs(162);
    layer0_outputs(12468) <= (inputs(24)) and not (inputs(15));
    layer0_outputs(12469) <= not(inputs(109));
    layer0_outputs(12470) <= not((inputs(156)) or (inputs(248)));
    layer0_outputs(12471) <= inputs(170);
    layer0_outputs(12472) <= (inputs(201)) or (inputs(225));
    layer0_outputs(12473) <= not(inputs(148));
    layer0_outputs(12474) <= (inputs(237)) or (inputs(178));
    layer0_outputs(12475) <= '0';
    layer0_outputs(12476) <= not((inputs(136)) xor (inputs(240)));
    layer0_outputs(12477) <= not((inputs(123)) or (inputs(238)));
    layer0_outputs(12478) <= (inputs(70)) or (inputs(108));
    layer0_outputs(12479) <= not(inputs(61));
    layer0_outputs(12480) <= not(inputs(121)) or (inputs(22));
    layer0_outputs(12481) <= (inputs(215)) xor (inputs(161));
    layer0_outputs(12482) <= (inputs(163)) or (inputs(90));
    layer0_outputs(12483) <= (inputs(242)) xor (inputs(145));
    layer0_outputs(12484) <= (inputs(109)) xor (inputs(24));
    layer0_outputs(12485) <= not(inputs(133)) or (inputs(225));
    layer0_outputs(12486) <= not(inputs(232));
    layer0_outputs(12487) <= not((inputs(17)) xor (inputs(3)));
    layer0_outputs(12488) <= inputs(27);
    layer0_outputs(12489) <= (inputs(222)) or (inputs(236));
    layer0_outputs(12490) <= inputs(215);
    layer0_outputs(12491) <= not(inputs(70)) or (inputs(143));
    layer0_outputs(12492) <= (inputs(105)) and not (inputs(1));
    layer0_outputs(12493) <= (inputs(164)) and not (inputs(250));
    layer0_outputs(12494) <= (inputs(163)) or (inputs(77));
    layer0_outputs(12495) <= not((inputs(181)) and (inputs(7)));
    layer0_outputs(12496) <= inputs(66);
    layer0_outputs(12497) <= not(inputs(30));
    layer0_outputs(12498) <= (inputs(172)) and (inputs(53));
    layer0_outputs(12499) <= not(inputs(145)) or (inputs(138));
    layer0_outputs(12500) <= (inputs(44)) or (inputs(29));
    layer0_outputs(12501) <= not(inputs(0));
    layer0_outputs(12502) <= (inputs(237)) and (inputs(94));
    layer0_outputs(12503) <= not(inputs(79));
    layer0_outputs(12504) <= (inputs(221)) xor (inputs(4));
    layer0_outputs(12505) <= not(inputs(81));
    layer0_outputs(12506) <= inputs(61);
    layer0_outputs(12507) <= (inputs(8)) xor (inputs(6));
    layer0_outputs(12508) <= not(inputs(254)) or (inputs(185));
    layer0_outputs(12509) <= not(inputs(91));
    layer0_outputs(12510) <= not(inputs(84));
    layer0_outputs(12511) <= '0';
    layer0_outputs(12512) <= not(inputs(164));
    layer0_outputs(12513) <= (inputs(84)) or (inputs(184));
    layer0_outputs(12514) <= inputs(99);
    layer0_outputs(12515) <= (inputs(103)) and not (inputs(160));
    layer0_outputs(12516) <= not((inputs(46)) or (inputs(234)));
    layer0_outputs(12517) <= not(inputs(46));
    layer0_outputs(12518) <= (inputs(31)) xor (inputs(193));
    layer0_outputs(12519) <= not(inputs(215));
    layer0_outputs(12520) <= inputs(230);
    layer0_outputs(12521) <= not(inputs(63));
    layer0_outputs(12522) <= (inputs(155)) and not (inputs(183));
    layer0_outputs(12523) <= not((inputs(119)) xor (inputs(246)));
    layer0_outputs(12524) <= not(inputs(0)) or (inputs(146));
    layer0_outputs(12525) <= (inputs(202)) and not (inputs(60));
    layer0_outputs(12526) <= not(inputs(244));
    layer0_outputs(12527) <= (inputs(32)) and (inputs(79));
    layer0_outputs(12528) <= inputs(34);
    layer0_outputs(12529) <= not(inputs(205));
    layer0_outputs(12530) <= inputs(246);
    layer0_outputs(12531) <= not(inputs(146));
    layer0_outputs(12532) <= (inputs(100)) and not (inputs(55));
    layer0_outputs(12533) <= (inputs(223)) or (inputs(171));
    layer0_outputs(12534) <= not(inputs(154));
    layer0_outputs(12535) <= not(inputs(90));
    layer0_outputs(12536) <= (inputs(138)) or (inputs(52));
    layer0_outputs(12537) <= inputs(10);
    layer0_outputs(12538) <= not(inputs(105)) or (inputs(16));
    layer0_outputs(12539) <= (inputs(147)) xor (inputs(217));
    layer0_outputs(12540) <= inputs(37);
    layer0_outputs(12541) <= not(inputs(207)) or (inputs(61));
    layer0_outputs(12542) <= not((inputs(78)) xor (inputs(20)));
    layer0_outputs(12543) <= not(inputs(39));
    layer0_outputs(12544) <= inputs(82);
    layer0_outputs(12545) <= not((inputs(182)) xor (inputs(183)));
    layer0_outputs(12546) <= (inputs(85)) or (inputs(205));
    layer0_outputs(12547) <= inputs(115);
    layer0_outputs(12548) <= (inputs(109)) and not (inputs(241));
    layer0_outputs(12549) <= (inputs(38)) and not (inputs(141));
    layer0_outputs(12550) <= (inputs(193)) or (inputs(129));
    layer0_outputs(12551) <= not((inputs(187)) xor (inputs(77)));
    layer0_outputs(12552) <= (inputs(148)) and not (inputs(96));
    layer0_outputs(12553) <= '1';
    layer0_outputs(12554) <= not((inputs(50)) or (inputs(104)));
    layer0_outputs(12555) <= not(inputs(61)) or (inputs(13));
    layer0_outputs(12556) <= not(inputs(213));
    layer0_outputs(12557) <= (inputs(92)) xor (inputs(134));
    layer0_outputs(12558) <= not((inputs(246)) xor (inputs(127)));
    layer0_outputs(12559) <= not((inputs(207)) xor (inputs(218)));
    layer0_outputs(12560) <= not(inputs(27));
    layer0_outputs(12561) <= not((inputs(216)) or (inputs(70)));
    layer0_outputs(12562) <= inputs(119);
    layer0_outputs(12563) <= not(inputs(40));
    layer0_outputs(12564) <= inputs(203);
    layer0_outputs(12565) <= (inputs(216)) or (inputs(195));
    layer0_outputs(12566) <= not((inputs(200)) or (inputs(238)));
    layer0_outputs(12567) <= not((inputs(197)) or (inputs(78)));
    layer0_outputs(12568) <= (inputs(216)) xor (inputs(190));
    layer0_outputs(12569) <= not((inputs(67)) xor (inputs(14)));
    layer0_outputs(12570) <= inputs(91);
    layer0_outputs(12571) <= (inputs(158)) or (inputs(79));
    layer0_outputs(12572) <= not(inputs(180));
    layer0_outputs(12573) <= not(inputs(83)) or (inputs(56));
    layer0_outputs(12574) <= inputs(203);
    layer0_outputs(12575) <= not(inputs(29));
    layer0_outputs(12576) <= not(inputs(7)) or (inputs(190));
    layer0_outputs(12577) <= (inputs(110)) or (inputs(212));
    layer0_outputs(12578) <= (inputs(22)) and not (inputs(155));
    layer0_outputs(12579) <= not((inputs(87)) xor (inputs(139)));
    layer0_outputs(12580) <= not(inputs(249));
    layer0_outputs(12581) <= not(inputs(66)) or (inputs(243));
    layer0_outputs(12582) <= not((inputs(4)) xor (inputs(224)));
    layer0_outputs(12583) <= (inputs(126)) xor (inputs(172));
    layer0_outputs(12584) <= (inputs(44)) or (inputs(14));
    layer0_outputs(12585) <= not((inputs(217)) xor (inputs(153)));
    layer0_outputs(12586) <= not((inputs(172)) or (inputs(11)));
    layer0_outputs(12587) <= not(inputs(7)) or (inputs(209));
    layer0_outputs(12588) <= not(inputs(177));
    layer0_outputs(12589) <= not((inputs(199)) xor (inputs(225)));
    layer0_outputs(12590) <= (inputs(72)) and not (inputs(67));
    layer0_outputs(12591) <= not((inputs(183)) or (inputs(173)));
    layer0_outputs(12592) <= (inputs(126)) or (inputs(178));
    layer0_outputs(12593) <= (inputs(230)) or (inputs(92));
    layer0_outputs(12594) <= inputs(23);
    layer0_outputs(12595) <= inputs(252);
    layer0_outputs(12596) <= not(inputs(229));
    layer0_outputs(12597) <= not((inputs(62)) or (inputs(213)));
    layer0_outputs(12598) <= not(inputs(45)) or (inputs(111));
    layer0_outputs(12599) <= (inputs(189)) xor (inputs(152));
    layer0_outputs(12600) <= (inputs(40)) or (inputs(30));
    layer0_outputs(12601) <= not(inputs(113));
    layer0_outputs(12602) <= inputs(81);
    layer0_outputs(12603) <= (inputs(224)) xor (inputs(14));
    layer0_outputs(12604) <= not(inputs(201)) or (inputs(221));
    layer0_outputs(12605) <= not(inputs(212)) or (inputs(4));
    layer0_outputs(12606) <= not(inputs(94)) or (inputs(208));
    layer0_outputs(12607) <= not(inputs(104)) or (inputs(98));
    layer0_outputs(12608) <= (inputs(124)) or (inputs(117));
    layer0_outputs(12609) <= not(inputs(13)) or (inputs(38));
    layer0_outputs(12610) <= not((inputs(47)) xor (inputs(106)));
    layer0_outputs(12611) <= '1';
    layer0_outputs(12612) <= not(inputs(207));
    layer0_outputs(12613) <= '0';
    layer0_outputs(12614) <= inputs(142);
    layer0_outputs(12615) <= (inputs(94)) xor (inputs(124));
    layer0_outputs(12616) <= (inputs(106)) or (inputs(183));
    layer0_outputs(12617) <= (inputs(250)) or (inputs(188));
    layer0_outputs(12618) <= not((inputs(186)) and (inputs(87)));
    layer0_outputs(12619) <= not((inputs(246)) xor (inputs(62)));
    layer0_outputs(12620) <= (inputs(152)) xor (inputs(229));
    layer0_outputs(12621) <= not((inputs(73)) xor (inputs(227)));
    layer0_outputs(12622) <= not(inputs(4));
    layer0_outputs(12623) <= not((inputs(68)) or (inputs(142)));
    layer0_outputs(12624) <= not(inputs(143));
    layer0_outputs(12625) <= not(inputs(53));
    layer0_outputs(12626) <= not((inputs(147)) xor (inputs(88)));
    layer0_outputs(12627) <= (inputs(4)) or (inputs(58));
    layer0_outputs(12628) <= (inputs(235)) and not (inputs(94));
    layer0_outputs(12629) <= not(inputs(248));
    layer0_outputs(12630) <= (inputs(166)) and not (inputs(51));
    layer0_outputs(12631) <= not(inputs(21));
    layer0_outputs(12632) <= inputs(20);
    layer0_outputs(12633) <= (inputs(57)) and not (inputs(192));
    layer0_outputs(12634) <= not(inputs(52)) or (inputs(244));
    layer0_outputs(12635) <= not((inputs(122)) or (inputs(159)));
    layer0_outputs(12636) <= not(inputs(223)) or (inputs(82));
    layer0_outputs(12637) <= not(inputs(59));
    layer0_outputs(12638) <= (inputs(151)) xor (inputs(130));
    layer0_outputs(12639) <= (inputs(232)) and (inputs(89));
    layer0_outputs(12640) <= inputs(147);
    layer0_outputs(12641) <= (inputs(121)) and not (inputs(227));
    layer0_outputs(12642) <= inputs(148);
    layer0_outputs(12643) <= (inputs(251)) or (inputs(50));
    layer0_outputs(12644) <= not(inputs(200));
    layer0_outputs(12645) <= not(inputs(207));
    layer0_outputs(12646) <= not((inputs(129)) xor (inputs(164)));
    layer0_outputs(12647) <= (inputs(250)) and not (inputs(127));
    layer0_outputs(12648) <= (inputs(217)) xor (inputs(255));
    layer0_outputs(12649) <= (inputs(239)) xor (inputs(11));
    layer0_outputs(12650) <= not((inputs(201)) xor (inputs(18)));
    layer0_outputs(12651) <= inputs(44);
    layer0_outputs(12652) <= not(inputs(199)) or (inputs(79));
    layer0_outputs(12653) <= not(inputs(59)) or (inputs(114));
    layer0_outputs(12654) <= (inputs(183)) or (inputs(143));
    layer0_outputs(12655) <= not(inputs(133));
    layer0_outputs(12656) <= not(inputs(114));
    layer0_outputs(12657) <= (inputs(118)) xor (inputs(182));
    layer0_outputs(12658) <= not((inputs(241)) xor (inputs(138)));
    layer0_outputs(12659) <= not(inputs(219));
    layer0_outputs(12660) <= not(inputs(174)) or (inputs(169));
    layer0_outputs(12661) <= (inputs(110)) and (inputs(33));
    layer0_outputs(12662) <= not((inputs(240)) xor (inputs(225)));
    layer0_outputs(12663) <= '0';
    layer0_outputs(12664) <= not(inputs(92));
    layer0_outputs(12665) <= inputs(10);
    layer0_outputs(12666) <= (inputs(18)) or (inputs(231));
    layer0_outputs(12667) <= inputs(248);
    layer0_outputs(12668) <= not((inputs(208)) or (inputs(183)));
    layer0_outputs(12669) <= (inputs(54)) or (inputs(93));
    layer0_outputs(12670) <= not((inputs(17)) or (inputs(19)));
    layer0_outputs(12671) <= not((inputs(214)) or (inputs(140)));
    layer0_outputs(12672) <= inputs(203);
    layer0_outputs(12673) <= inputs(27);
    layer0_outputs(12674) <= (inputs(247)) and not (inputs(134));
    layer0_outputs(12675) <= not((inputs(245)) or (inputs(209)));
    layer0_outputs(12676) <= not(inputs(84));
    layer0_outputs(12677) <= (inputs(99)) and not (inputs(79));
    layer0_outputs(12678) <= (inputs(79)) or (inputs(128));
    layer0_outputs(12679) <= not((inputs(150)) and (inputs(145)));
    layer0_outputs(12680) <= not(inputs(245)) or (inputs(136));
    layer0_outputs(12681) <= not(inputs(182));
    layer0_outputs(12682) <= inputs(139);
    layer0_outputs(12683) <= not((inputs(68)) or (inputs(49)));
    layer0_outputs(12684) <= not(inputs(254));
    layer0_outputs(12685) <= not(inputs(242)) or (inputs(169));
    layer0_outputs(12686) <= not(inputs(164));
    layer0_outputs(12687) <= (inputs(52)) and not (inputs(190));
    layer0_outputs(12688) <= not((inputs(24)) or (inputs(160)));
    layer0_outputs(12689) <= (inputs(225)) and not (inputs(1));
    layer0_outputs(12690) <= inputs(250);
    layer0_outputs(12691) <= not(inputs(41)) or (inputs(184));
    layer0_outputs(12692) <= not((inputs(14)) or (inputs(34)));
    layer0_outputs(12693) <= not(inputs(127));
    layer0_outputs(12694) <= (inputs(196)) and not (inputs(130));
    layer0_outputs(12695) <= (inputs(151)) and not (inputs(98));
    layer0_outputs(12696) <= not((inputs(227)) or (inputs(148)));
    layer0_outputs(12697) <= not((inputs(20)) or (inputs(81)));
    layer0_outputs(12698) <= (inputs(110)) xor (inputs(74));
    layer0_outputs(12699) <= inputs(80);
    layer0_outputs(12700) <= (inputs(236)) or (inputs(191));
    layer0_outputs(12701) <= (inputs(98)) xor (inputs(29));
    layer0_outputs(12702) <= not(inputs(149)) or (inputs(221));
    layer0_outputs(12703) <= not(inputs(91));
    layer0_outputs(12704) <= (inputs(219)) xor (inputs(96));
    layer0_outputs(12705) <= not(inputs(131));
    layer0_outputs(12706) <= not(inputs(181));
    layer0_outputs(12707) <= not((inputs(187)) xor (inputs(37)));
    layer0_outputs(12708) <= (inputs(82)) xor (inputs(187));
    layer0_outputs(12709) <= (inputs(101)) and (inputs(227));
    layer0_outputs(12710) <= not((inputs(18)) xor (inputs(65)));
    layer0_outputs(12711) <= not(inputs(102));
    layer0_outputs(12712) <= (inputs(183)) and not (inputs(117));
    layer0_outputs(12713) <= (inputs(192)) and not (inputs(15));
    layer0_outputs(12714) <= (inputs(104)) or (inputs(2));
    layer0_outputs(12715) <= (inputs(109)) xor (inputs(80));
    layer0_outputs(12716) <= (inputs(49)) or (inputs(126));
    layer0_outputs(12717) <= not(inputs(183));
    layer0_outputs(12718) <= (inputs(233)) xor (inputs(62));
    layer0_outputs(12719) <= not(inputs(211));
    layer0_outputs(12720) <= not((inputs(254)) xor (inputs(33)));
    layer0_outputs(12721) <= not((inputs(198)) xor (inputs(224)));
    layer0_outputs(12722) <= not(inputs(61));
    layer0_outputs(12723) <= not(inputs(132)) or (inputs(19));
    layer0_outputs(12724) <= not((inputs(146)) or (inputs(194)));
    layer0_outputs(12725) <= (inputs(147)) and not (inputs(33));
    layer0_outputs(12726) <= not(inputs(65)) or (inputs(111));
    layer0_outputs(12727) <= not((inputs(214)) xor (inputs(9)));
    layer0_outputs(12728) <= not(inputs(233)) or (inputs(105));
    layer0_outputs(12729) <= (inputs(201)) xor (inputs(233));
    layer0_outputs(12730) <= inputs(215);
    layer0_outputs(12731) <= not(inputs(252));
    layer0_outputs(12732) <= (inputs(188)) or (inputs(248));
    layer0_outputs(12733) <= not(inputs(100)) or (inputs(111));
    layer0_outputs(12734) <= not((inputs(5)) or (inputs(3)));
    layer0_outputs(12735) <= not((inputs(26)) and (inputs(124)));
    layer0_outputs(12736) <= (inputs(233)) and (inputs(154));
    layer0_outputs(12737) <= not(inputs(217));
    layer0_outputs(12738) <= (inputs(181)) xor (inputs(237));
    layer0_outputs(12739) <= not((inputs(8)) and (inputs(169)));
    layer0_outputs(12740) <= not((inputs(25)) or (inputs(95)));
    layer0_outputs(12741) <= not(inputs(181)) or (inputs(124));
    layer0_outputs(12742) <= not(inputs(38)) or (inputs(115));
    layer0_outputs(12743) <= not(inputs(84)) or (inputs(159));
    layer0_outputs(12744) <= not(inputs(8));
    layer0_outputs(12745) <= not(inputs(163));
    layer0_outputs(12746) <= not((inputs(211)) or (inputs(188)));
    layer0_outputs(12747) <= not((inputs(194)) or (inputs(185)));
    layer0_outputs(12748) <= (inputs(211)) and not (inputs(137));
    layer0_outputs(12749) <= inputs(212);
    layer0_outputs(12750) <= not((inputs(170)) xor (inputs(98)));
    layer0_outputs(12751) <= not(inputs(84));
    layer0_outputs(12752) <= not(inputs(178)) or (inputs(124));
    layer0_outputs(12753) <= not((inputs(116)) or (inputs(253)));
    layer0_outputs(12754) <= (inputs(203)) xor (inputs(232));
    layer0_outputs(12755) <= not(inputs(208)) or (inputs(84));
    layer0_outputs(12756) <= not((inputs(164)) or (inputs(254)));
    layer0_outputs(12757) <= not(inputs(180));
    layer0_outputs(12758) <= (inputs(213)) and (inputs(194));
    layer0_outputs(12759) <= not((inputs(178)) or (inputs(54)));
    layer0_outputs(12760) <= inputs(137);
    layer0_outputs(12761) <= not((inputs(8)) xor (inputs(69)));
    layer0_outputs(12762) <= not((inputs(129)) xor (inputs(158)));
    layer0_outputs(12763) <= inputs(199);
    layer0_outputs(12764) <= not((inputs(214)) xor (inputs(80)));
    layer0_outputs(12765) <= not(inputs(240));
    layer0_outputs(12766) <= '0';
    layer0_outputs(12767) <= inputs(136);
    layer0_outputs(12768) <= not((inputs(170)) xor (inputs(217)));
    layer0_outputs(12769) <= (inputs(106)) and not (inputs(243));
    layer0_outputs(12770) <= (inputs(217)) or (inputs(217));
    layer0_outputs(12771) <= '1';
    layer0_outputs(12772) <= not(inputs(131));
    layer0_outputs(12773) <= (inputs(84)) or (inputs(18));
    layer0_outputs(12774) <= not(inputs(70)) or (inputs(243));
    layer0_outputs(12775) <= (inputs(63)) xor (inputs(102));
    layer0_outputs(12776) <= not((inputs(31)) or (inputs(64)));
    layer0_outputs(12777) <= not(inputs(196)) or (inputs(1));
    layer0_outputs(12778) <= not((inputs(251)) or (inputs(184)));
    layer0_outputs(12779) <= not((inputs(144)) or (inputs(80)));
    layer0_outputs(12780) <= (inputs(141)) and not (inputs(143));
    layer0_outputs(12781) <= (inputs(26)) and not (inputs(104));
    layer0_outputs(12782) <= not(inputs(161));
    layer0_outputs(12783) <= inputs(77);
    layer0_outputs(12784) <= not(inputs(136)) or (inputs(255));
    layer0_outputs(12785) <= inputs(101);
    layer0_outputs(12786) <= not(inputs(174)) or (inputs(29));
    layer0_outputs(12787) <= not((inputs(105)) xor (inputs(9)));
    layer0_outputs(12788) <= (inputs(199)) and (inputs(205));
    layer0_outputs(12789) <= (inputs(75)) and not (inputs(152));
    layer0_outputs(12790) <= not(inputs(243)) or (inputs(254));
    layer0_outputs(12791) <= inputs(152);
    layer0_outputs(12792) <= not((inputs(23)) or (inputs(190)));
    layer0_outputs(12793) <= not(inputs(138));
    layer0_outputs(12794) <= not((inputs(252)) xor (inputs(50)));
    layer0_outputs(12795) <= not(inputs(216));
    layer0_outputs(12796) <= (inputs(159)) or (inputs(157));
    layer0_outputs(12797) <= inputs(124);
    layer0_outputs(12798) <= inputs(194);
    layer0_outputs(12799) <= (inputs(105)) and not (inputs(254));
    outputs(0) <= layer0_outputs(3077);
    outputs(1) <= layer0_outputs(4276);
    outputs(2) <= not((layer0_outputs(2875)) xor (layer0_outputs(8415)));
    outputs(3) <= (layer0_outputs(7184)) and (layer0_outputs(8018));
    outputs(4) <= (layer0_outputs(2071)) xor (layer0_outputs(3468));
    outputs(5) <= layer0_outputs(6286);
    outputs(6) <= not(layer0_outputs(3496));
    outputs(7) <= not(layer0_outputs(7946)) or (layer0_outputs(12729));
    outputs(8) <= (layer0_outputs(4014)) and (layer0_outputs(3095));
    outputs(9) <= layer0_outputs(11610);
    outputs(10) <= layer0_outputs(2767);
    outputs(11) <= not((layer0_outputs(8277)) xor (layer0_outputs(9779)));
    outputs(12) <= not(layer0_outputs(721)) or (layer0_outputs(3589));
    outputs(13) <= not(layer0_outputs(6289));
    outputs(14) <= (layer0_outputs(1038)) xor (layer0_outputs(3037));
    outputs(15) <= not(layer0_outputs(4016));
    outputs(16) <= not(layer0_outputs(10706));
    outputs(17) <= (layer0_outputs(2317)) xor (layer0_outputs(4491));
    outputs(18) <= layer0_outputs(1922);
    outputs(19) <= not((layer0_outputs(7064)) xor (layer0_outputs(10666)));
    outputs(20) <= layer0_outputs(5761);
    outputs(21) <= not(layer0_outputs(10278)) or (layer0_outputs(4447));
    outputs(22) <= (layer0_outputs(9534)) xor (layer0_outputs(10938));
    outputs(23) <= not(layer0_outputs(1373)) or (layer0_outputs(958));
    outputs(24) <= (layer0_outputs(8369)) xor (layer0_outputs(10362));
    outputs(25) <= not((layer0_outputs(3923)) xor (layer0_outputs(4670)));
    outputs(26) <= not(layer0_outputs(7774));
    outputs(27) <= not(layer0_outputs(11064));
    outputs(28) <= not(layer0_outputs(11361)) or (layer0_outputs(10573));
    outputs(29) <= (layer0_outputs(7287)) and (layer0_outputs(3021));
    outputs(30) <= layer0_outputs(11759);
    outputs(31) <= not(layer0_outputs(230)) or (layer0_outputs(2779));
    outputs(32) <= not((layer0_outputs(3483)) xor (layer0_outputs(4502)));
    outputs(33) <= layer0_outputs(5910);
    outputs(34) <= not(layer0_outputs(10974));
    outputs(35) <= not((layer0_outputs(10171)) xor (layer0_outputs(5812)));
    outputs(36) <= layer0_outputs(7346);
    outputs(37) <= (layer0_outputs(11826)) and not (layer0_outputs(5429));
    outputs(38) <= not((layer0_outputs(2014)) xor (layer0_outputs(3589)));
    outputs(39) <= not((layer0_outputs(6985)) xor (layer0_outputs(824)));
    outputs(40) <= not(layer0_outputs(11269));
    outputs(41) <= (layer0_outputs(8455)) xor (layer0_outputs(9084));
    outputs(42) <= (layer0_outputs(3646)) xor (layer0_outputs(480));
    outputs(43) <= not((layer0_outputs(12507)) xor (layer0_outputs(5281)));
    outputs(44) <= not(layer0_outputs(9250));
    outputs(45) <= not((layer0_outputs(10665)) xor (layer0_outputs(6723)));
    outputs(46) <= not((layer0_outputs(9156)) xor (layer0_outputs(7558)));
    outputs(47) <= not(layer0_outputs(7722));
    outputs(48) <= (layer0_outputs(3777)) xor (layer0_outputs(8122));
    outputs(49) <= (layer0_outputs(1015)) and not (layer0_outputs(3293));
    outputs(50) <= (layer0_outputs(9954)) and not (layer0_outputs(9984));
    outputs(51) <= (layer0_outputs(2671)) xor (layer0_outputs(11734));
    outputs(52) <= (layer0_outputs(4088)) xor (layer0_outputs(7093));
    outputs(53) <= not(layer0_outputs(12068)) or (layer0_outputs(58));
    outputs(54) <= layer0_outputs(5686);
    outputs(55) <= layer0_outputs(7229);
    outputs(56) <= layer0_outputs(3100);
    outputs(57) <= not(layer0_outputs(12438));
    outputs(58) <= (layer0_outputs(1390)) xor (layer0_outputs(1801));
    outputs(59) <= (layer0_outputs(12178)) and (layer0_outputs(8020));
    outputs(60) <= (layer0_outputs(10842)) xor (layer0_outputs(8736));
    outputs(61) <= (layer0_outputs(2580)) xor (layer0_outputs(5849));
    outputs(62) <= (layer0_outputs(2019)) or (layer0_outputs(2683));
    outputs(63) <= not(layer0_outputs(12637));
    outputs(64) <= layer0_outputs(6762);
    outputs(65) <= not((layer0_outputs(8050)) and (layer0_outputs(9158)));
    outputs(66) <= not((layer0_outputs(9439)) xor (layer0_outputs(2575)));
    outputs(67) <= not(layer0_outputs(10373));
    outputs(68) <= layer0_outputs(248);
    outputs(69) <= layer0_outputs(11550);
    outputs(70) <= (layer0_outputs(3682)) and (layer0_outputs(6491));
    outputs(71) <= not((layer0_outputs(4229)) or (layer0_outputs(11355)));
    outputs(72) <= (layer0_outputs(6825)) or (layer0_outputs(7400));
    outputs(73) <= not((layer0_outputs(12703)) xor (layer0_outputs(3576)));
    outputs(74) <= not(layer0_outputs(5239));
    outputs(75) <= (layer0_outputs(5316)) and not (layer0_outputs(8430));
    outputs(76) <= not((layer0_outputs(5706)) xor (layer0_outputs(4575)));
    outputs(77) <= not(layer0_outputs(9696));
    outputs(78) <= (layer0_outputs(2425)) xor (layer0_outputs(3551));
    outputs(79) <= not(layer0_outputs(9173));
    outputs(80) <= not(layer0_outputs(10247));
    outputs(81) <= layer0_outputs(652);
    outputs(82) <= layer0_outputs(8089);
    outputs(83) <= layer0_outputs(12715);
    outputs(84) <= not(layer0_outputs(1578)) or (layer0_outputs(6197));
    outputs(85) <= (layer0_outputs(12477)) xor (layer0_outputs(3006));
    outputs(86) <= not(layer0_outputs(12002));
    outputs(87) <= (layer0_outputs(11597)) and not (layer0_outputs(10593));
    outputs(88) <= not((layer0_outputs(1946)) or (layer0_outputs(5149)));
    outputs(89) <= not(layer0_outputs(746));
    outputs(90) <= layer0_outputs(9650);
    outputs(91) <= not(layer0_outputs(7957));
    outputs(92) <= not(layer0_outputs(2161));
    outputs(93) <= not((layer0_outputs(2004)) xor (layer0_outputs(9280)));
    outputs(94) <= (layer0_outputs(5339)) xor (layer0_outputs(2074));
    outputs(95) <= (layer0_outputs(12571)) or (layer0_outputs(1101));
    outputs(96) <= '1';
    outputs(97) <= not(layer0_outputs(11304));
    outputs(98) <= not(layer0_outputs(4901));
    outputs(99) <= layer0_outputs(1564);
    outputs(100) <= not((layer0_outputs(4609)) xor (layer0_outputs(1356)));
    outputs(101) <= (layer0_outputs(8917)) and (layer0_outputs(2885));
    outputs(102) <= not(layer0_outputs(1811));
    outputs(103) <= not(layer0_outputs(73));
    outputs(104) <= (layer0_outputs(9406)) and (layer0_outputs(9071));
    outputs(105) <= not(layer0_outputs(4207));
    outputs(106) <= layer0_outputs(597);
    outputs(107) <= layer0_outputs(3461);
    outputs(108) <= (layer0_outputs(6213)) xor (layer0_outputs(8404));
    outputs(109) <= layer0_outputs(2846);
    outputs(110) <= (layer0_outputs(576)) xor (layer0_outputs(11285));
    outputs(111) <= layer0_outputs(9401);
    outputs(112) <= (layer0_outputs(2060)) xor (layer0_outputs(6628));
    outputs(113) <= not((layer0_outputs(2130)) xor (layer0_outputs(9512)));
    outputs(114) <= layer0_outputs(7417);
    outputs(115) <= not((layer0_outputs(8397)) xor (layer0_outputs(7027)));
    outputs(116) <= not((layer0_outputs(12011)) xor (layer0_outputs(10904)));
    outputs(117) <= not((layer0_outputs(998)) xor (layer0_outputs(3074)));
    outputs(118) <= layer0_outputs(4257);
    outputs(119) <= not(layer0_outputs(10929));
    outputs(120) <= not(layer0_outputs(7881));
    outputs(121) <= (layer0_outputs(7143)) xor (layer0_outputs(11420));
    outputs(122) <= not((layer0_outputs(7751)) xor (layer0_outputs(10069)));
    outputs(123) <= not((layer0_outputs(8136)) xor (layer0_outputs(11045)));
    outputs(124) <= (layer0_outputs(3890)) and not (layer0_outputs(2616));
    outputs(125) <= (layer0_outputs(4717)) xor (layer0_outputs(283));
    outputs(126) <= layer0_outputs(3680);
    outputs(127) <= (layer0_outputs(8386)) or (layer0_outputs(12498));
    outputs(128) <= not((layer0_outputs(7478)) and (layer0_outputs(8243)));
    outputs(129) <= (layer0_outputs(6831)) and (layer0_outputs(10071));
    outputs(130) <= not((layer0_outputs(8973)) or (layer0_outputs(5127)));
    outputs(131) <= not((layer0_outputs(2248)) and (layer0_outputs(7812)));
    outputs(132) <= not((layer0_outputs(6917)) xor (layer0_outputs(7113)));
    outputs(133) <= not((layer0_outputs(562)) and (layer0_outputs(9882)));
    outputs(134) <= not(layer0_outputs(2080)) or (layer0_outputs(3885));
    outputs(135) <= not((layer0_outputs(9589)) xor (layer0_outputs(1324)));
    outputs(136) <= not((layer0_outputs(6546)) xor (layer0_outputs(5039)));
    outputs(137) <= not((layer0_outputs(7770)) xor (layer0_outputs(9498)));
    outputs(138) <= (layer0_outputs(11317)) xor (layer0_outputs(7022));
    outputs(139) <= not(layer0_outputs(4470));
    outputs(140) <= not(layer0_outputs(3312));
    outputs(141) <= not(layer0_outputs(3318));
    outputs(142) <= not((layer0_outputs(6466)) and (layer0_outputs(1636)));
    outputs(143) <= (layer0_outputs(10422)) and not (layer0_outputs(10249));
    outputs(144) <= not(layer0_outputs(11563));
    outputs(145) <= layer0_outputs(9997);
    outputs(146) <= layer0_outputs(1763);
    outputs(147) <= not(layer0_outputs(7443));
    outputs(148) <= not((layer0_outputs(5323)) xor (layer0_outputs(10039)));
    outputs(149) <= not((layer0_outputs(5557)) xor (layer0_outputs(6092)));
    outputs(150) <= not(layer0_outputs(9615));
    outputs(151) <= not(layer0_outputs(11741));
    outputs(152) <= layer0_outputs(6669);
    outputs(153) <= not(layer0_outputs(10973));
    outputs(154) <= not(layer0_outputs(9653)) or (layer0_outputs(8507));
    outputs(155) <= not(layer0_outputs(12675));
    outputs(156) <= layer0_outputs(442);
    outputs(157) <= not(layer0_outputs(9846));
    outputs(158) <= not((layer0_outputs(4506)) or (layer0_outputs(8284)));
    outputs(159) <= not(layer0_outputs(10475));
    outputs(160) <= not(layer0_outputs(9838));
    outputs(161) <= (layer0_outputs(6936)) and (layer0_outputs(10666));
    outputs(162) <= layer0_outputs(5737);
    outputs(163) <= not(layer0_outputs(12769));
    outputs(164) <= not((layer0_outputs(7288)) xor (layer0_outputs(2172)));
    outputs(165) <= (layer0_outputs(2313)) and not (layer0_outputs(7160));
    outputs(166) <= layer0_outputs(4779);
    outputs(167) <= (layer0_outputs(7182)) xor (layer0_outputs(11711));
    outputs(168) <= not(layer0_outputs(313));
    outputs(169) <= layer0_outputs(133);
    outputs(170) <= not(layer0_outputs(4133));
    outputs(171) <= layer0_outputs(10907);
    outputs(172) <= not(layer0_outputs(7123)) or (layer0_outputs(9872));
    outputs(173) <= layer0_outputs(12374);
    outputs(174) <= not((layer0_outputs(5837)) xor (layer0_outputs(2587)));
    outputs(175) <= not(layer0_outputs(113));
    outputs(176) <= not(layer0_outputs(9142));
    outputs(177) <= not((layer0_outputs(12081)) xor (layer0_outputs(10993)));
    outputs(178) <= not(layer0_outputs(5084));
    outputs(179) <= (layer0_outputs(11386)) xor (layer0_outputs(10115));
    outputs(180) <= not((layer0_outputs(12135)) or (layer0_outputs(11949)));
    outputs(181) <= layer0_outputs(9438);
    outputs(182) <= not(layer0_outputs(5867));
    outputs(183) <= layer0_outputs(3385);
    outputs(184) <= (layer0_outputs(9034)) xor (layer0_outputs(600));
    outputs(185) <= not((layer0_outputs(11899)) or (layer0_outputs(4227)));
    outputs(186) <= not(layer0_outputs(1149));
    outputs(187) <= not(layer0_outputs(5424));
    outputs(188) <= not((layer0_outputs(140)) xor (layer0_outputs(5726)));
    outputs(189) <= not(layer0_outputs(1656));
    outputs(190) <= not(layer0_outputs(8686));
    outputs(191) <= not(layer0_outputs(1290));
    outputs(192) <= not((layer0_outputs(11935)) xor (layer0_outputs(12017)));
    outputs(193) <= layer0_outputs(6206);
    outputs(194) <= (layer0_outputs(8439)) and not (layer0_outputs(11933));
    outputs(195) <= not(layer0_outputs(1175)) or (layer0_outputs(11630));
    outputs(196) <= layer0_outputs(3099);
    outputs(197) <= layer0_outputs(11052);
    outputs(198) <= layer0_outputs(3982);
    outputs(199) <= not((layer0_outputs(4998)) or (layer0_outputs(437)));
    outputs(200) <= layer0_outputs(2375);
    outputs(201) <= (layer0_outputs(8779)) and not (layer0_outputs(5055));
    outputs(202) <= (layer0_outputs(7808)) xor (layer0_outputs(3344));
    outputs(203) <= not((layer0_outputs(10850)) or (layer0_outputs(5931)));
    outputs(204) <= (layer0_outputs(7618)) xor (layer0_outputs(10772));
    outputs(205) <= not(layer0_outputs(9087)) or (layer0_outputs(9632));
    outputs(206) <= layer0_outputs(8966);
    outputs(207) <= not(layer0_outputs(10922)) or (layer0_outputs(11571));
    outputs(208) <= not(layer0_outputs(12024));
    outputs(209) <= layer0_outputs(4234);
    outputs(210) <= (layer0_outputs(1385)) or (layer0_outputs(1842));
    outputs(211) <= layer0_outputs(3050);
    outputs(212) <= not(layer0_outputs(9491));
    outputs(213) <= (layer0_outputs(3507)) and not (layer0_outputs(10204));
    outputs(214) <= (layer0_outputs(11857)) xor (layer0_outputs(12740));
    outputs(215) <= layer0_outputs(2548);
    outputs(216) <= not(layer0_outputs(10246));
    outputs(217) <= (layer0_outputs(4732)) and (layer0_outputs(50));
    outputs(218) <= (layer0_outputs(4399)) and not (layer0_outputs(6607));
    outputs(219) <= not((layer0_outputs(12674)) xor (layer0_outputs(1344)));
    outputs(220) <= layer0_outputs(12389);
    outputs(221) <= (layer0_outputs(7172)) or (layer0_outputs(2166));
    outputs(222) <= (layer0_outputs(12312)) xor (layer0_outputs(5515));
    outputs(223) <= layer0_outputs(4765);
    outputs(224) <= not(layer0_outputs(9385));
    outputs(225) <= (layer0_outputs(6797)) xor (layer0_outputs(11296));
    outputs(226) <= layer0_outputs(8386);
    outputs(227) <= not((layer0_outputs(2606)) and (layer0_outputs(10793)));
    outputs(228) <= (layer0_outputs(9193)) xor (layer0_outputs(8611));
    outputs(229) <= not((layer0_outputs(1196)) xor (layer0_outputs(12377)));
    outputs(230) <= (layer0_outputs(7689)) xor (layer0_outputs(4745));
    outputs(231) <= (layer0_outputs(4581)) and (layer0_outputs(9267));
    outputs(232) <= (layer0_outputs(10055)) xor (layer0_outputs(11523));
    outputs(233) <= not(layer0_outputs(6011));
    outputs(234) <= not(layer0_outputs(9142));
    outputs(235) <= (layer0_outputs(5503)) xor (layer0_outputs(5305));
    outputs(236) <= layer0_outputs(10995);
    outputs(237) <= layer0_outputs(1115);
    outputs(238) <= (layer0_outputs(7364)) xor (layer0_outputs(9572));
    outputs(239) <= not(layer0_outputs(4686));
    outputs(240) <= (layer0_outputs(10807)) xor (layer0_outputs(1233));
    outputs(241) <= not(layer0_outputs(1903));
    outputs(242) <= layer0_outputs(7359);
    outputs(243) <= not(layer0_outputs(10685));
    outputs(244) <= layer0_outputs(2228);
    outputs(245) <= not(layer0_outputs(8717)) or (layer0_outputs(11079));
    outputs(246) <= not(layer0_outputs(8892));
    outputs(247) <= (layer0_outputs(12313)) xor (layer0_outputs(9054));
    outputs(248) <= not(layer0_outputs(10507)) or (layer0_outputs(6238));
    outputs(249) <= (layer0_outputs(10607)) xor (layer0_outputs(5888));
    outputs(250) <= not((layer0_outputs(4641)) xor (layer0_outputs(1572)));
    outputs(251) <= (layer0_outputs(9940)) xor (layer0_outputs(2789));
    outputs(252) <= not(layer0_outputs(4658));
    outputs(253) <= not(layer0_outputs(9678));
    outputs(254) <= not(layer0_outputs(7646));
    outputs(255) <= not(layer0_outputs(7705));
    outputs(256) <= (layer0_outputs(11182)) xor (layer0_outputs(11668));
    outputs(257) <= not(layer0_outputs(5553));
    outputs(258) <= layer0_outputs(8428);
    outputs(259) <= not(layer0_outputs(3892));
    outputs(260) <= layer0_outputs(5626);
    outputs(261) <= layer0_outputs(10144);
    outputs(262) <= layer0_outputs(947);
    outputs(263) <= layer0_outputs(1427);
    outputs(264) <= not(layer0_outputs(10160));
    outputs(265) <= not(layer0_outputs(12320));
    outputs(266) <= not((layer0_outputs(7648)) or (layer0_outputs(6870)));
    outputs(267) <= (layer0_outputs(4182)) xor (layer0_outputs(5268));
    outputs(268) <= layer0_outputs(5963);
    outputs(269) <= layer0_outputs(1638);
    outputs(270) <= not((layer0_outputs(4983)) xor (layer0_outputs(380)));
    outputs(271) <= not(layer0_outputs(6463)) or (layer0_outputs(2237));
    outputs(272) <= not((layer0_outputs(11177)) xor (layer0_outputs(2416)));
    outputs(273) <= (layer0_outputs(7650)) or (layer0_outputs(3963));
    outputs(274) <= (layer0_outputs(270)) xor (layer0_outputs(4724));
    outputs(275) <= layer0_outputs(105);
    outputs(276) <= layer0_outputs(5347);
    outputs(277) <= not(layer0_outputs(5586));
    outputs(278) <= layer0_outputs(10704);
    outputs(279) <= layer0_outputs(4730);
    outputs(280) <= not((layer0_outputs(11631)) and (layer0_outputs(9023)));
    outputs(281) <= not(layer0_outputs(6692)) or (layer0_outputs(11151));
    outputs(282) <= not((layer0_outputs(7042)) xor (layer0_outputs(6041)));
    outputs(283) <= not(layer0_outputs(888));
    outputs(284) <= not(layer0_outputs(8589));
    outputs(285) <= layer0_outputs(8018);
    outputs(286) <= layer0_outputs(6352);
    outputs(287) <= not(layer0_outputs(12771)) or (layer0_outputs(4375));
    outputs(288) <= not(layer0_outputs(8375));
    outputs(289) <= layer0_outputs(8469);
    outputs(290) <= not((layer0_outputs(4494)) xor (layer0_outputs(11358)));
    outputs(291) <= (layer0_outputs(4615)) and not (layer0_outputs(12381));
    outputs(292) <= not(layer0_outputs(8345));
    outputs(293) <= not((layer0_outputs(3319)) and (layer0_outputs(233)));
    outputs(294) <= not(layer0_outputs(5912));
    outputs(295) <= not((layer0_outputs(9304)) xor (layer0_outputs(10898)));
    outputs(296) <= (layer0_outputs(12151)) and not (layer0_outputs(7698));
    outputs(297) <= (layer0_outputs(4434)) xor (layer0_outputs(7013));
    outputs(298) <= (layer0_outputs(12598)) and not (layer0_outputs(4919));
    outputs(299) <= layer0_outputs(6978);
    outputs(300) <= not(layer0_outputs(4999)) or (layer0_outputs(9960));
    outputs(301) <= layer0_outputs(6939);
    outputs(302) <= (layer0_outputs(695)) xor (layer0_outputs(8733));
    outputs(303) <= layer0_outputs(1503);
    outputs(304) <= not(layer0_outputs(6466));
    outputs(305) <= not(layer0_outputs(10851)) or (layer0_outputs(3534));
    outputs(306) <= layer0_outputs(6410);
    outputs(307) <= (layer0_outputs(3004)) and not (layer0_outputs(581));
    outputs(308) <= layer0_outputs(9103);
    outputs(309) <= (layer0_outputs(2794)) xor (layer0_outputs(10721));
    outputs(310) <= not((layer0_outputs(3895)) and (layer0_outputs(10500)));
    outputs(311) <= not((layer0_outputs(2615)) and (layer0_outputs(7931)));
    outputs(312) <= not(layer0_outputs(1453));
    outputs(313) <= not((layer0_outputs(1428)) xor (layer0_outputs(8522)));
    outputs(314) <= not(layer0_outputs(6676));
    outputs(315) <= not((layer0_outputs(5375)) and (layer0_outputs(2586)));
    outputs(316) <= (layer0_outputs(5642)) and (layer0_outputs(5945));
    outputs(317) <= not(layer0_outputs(12686));
    outputs(318) <= (layer0_outputs(8072)) xor (layer0_outputs(458));
    outputs(319) <= (layer0_outputs(5100)) xor (layer0_outputs(8149));
    outputs(320) <= not(layer0_outputs(9764));
    outputs(321) <= not((layer0_outputs(9657)) and (layer0_outputs(6977)));
    outputs(322) <= (layer0_outputs(4913)) and not (layer0_outputs(11671));
    outputs(323) <= not(layer0_outputs(8872));
    outputs(324) <= not(layer0_outputs(9050));
    outputs(325) <= not((layer0_outputs(12464)) or (layer0_outputs(8178)));
    outputs(326) <= layer0_outputs(10598);
    outputs(327) <= not(layer0_outputs(4122));
    outputs(328) <= not(layer0_outputs(11000));
    outputs(329) <= (layer0_outputs(2354)) xor (layer0_outputs(6217));
    outputs(330) <= not(layer0_outputs(2189));
    outputs(331) <= not((layer0_outputs(9466)) xor (layer0_outputs(3043)));
    outputs(332) <= not((layer0_outputs(2418)) and (layer0_outputs(1157)));
    outputs(333) <= not(layer0_outputs(9376)) or (layer0_outputs(9031));
    outputs(334) <= not(layer0_outputs(919));
    outputs(335) <= not((layer0_outputs(9977)) xor (layer0_outputs(12469)));
    outputs(336) <= layer0_outputs(832);
    outputs(337) <= (layer0_outputs(9262)) and not (layer0_outputs(10833));
    outputs(338) <= not(layer0_outputs(12293));
    outputs(339) <= layer0_outputs(7230);
    outputs(340) <= (layer0_outputs(522)) xor (layer0_outputs(10680));
    outputs(341) <= not((layer0_outputs(9963)) xor (layer0_outputs(10697)));
    outputs(342) <= not((layer0_outputs(9124)) xor (layer0_outputs(9367)));
    outputs(343) <= layer0_outputs(11069);
    outputs(344) <= not((layer0_outputs(2128)) xor (layer0_outputs(9047)));
    outputs(345) <= (layer0_outputs(83)) xor (layer0_outputs(9154));
    outputs(346) <= layer0_outputs(8853);
    outputs(347) <= not((layer0_outputs(5666)) or (layer0_outputs(11254)));
    outputs(348) <= not(layer0_outputs(10444));
    outputs(349) <= not(layer0_outputs(9754));
    outputs(350) <= not((layer0_outputs(11671)) or (layer0_outputs(10627)));
    outputs(351) <= (layer0_outputs(7310)) or (layer0_outputs(6103));
    outputs(352) <= not(layer0_outputs(11827));
    outputs(353) <= (layer0_outputs(5883)) xor (layer0_outputs(8141));
    outputs(354) <= layer0_outputs(5975);
    outputs(355) <= layer0_outputs(3055);
    outputs(356) <= layer0_outputs(5582);
    outputs(357) <= not(layer0_outputs(460)) or (layer0_outputs(8682));
    outputs(358) <= (layer0_outputs(7322)) and (layer0_outputs(7717));
    outputs(359) <= layer0_outputs(5271);
    outputs(360) <= layer0_outputs(11650);
    outputs(361) <= not(layer0_outputs(1759));
    outputs(362) <= layer0_outputs(3052);
    outputs(363) <= layer0_outputs(6478);
    outputs(364) <= layer0_outputs(1923);
    outputs(365) <= not(layer0_outputs(587));
    outputs(366) <= layer0_outputs(790);
    outputs(367) <= layer0_outputs(7768);
    outputs(368) <= not((layer0_outputs(11990)) and (layer0_outputs(3034)));
    outputs(369) <= not((layer0_outputs(3023)) xor (layer0_outputs(7404)));
    outputs(370) <= not((layer0_outputs(10111)) and (layer0_outputs(9213)));
    outputs(371) <= layer0_outputs(4053);
    outputs(372) <= (layer0_outputs(11096)) xor (layer0_outputs(10133));
    outputs(373) <= not(layer0_outputs(8930));
    outputs(374) <= not((layer0_outputs(9058)) xor (layer0_outputs(5442)));
    outputs(375) <= layer0_outputs(4893);
    outputs(376) <= not(layer0_outputs(12052));
    outputs(377) <= layer0_outputs(2837);
    outputs(378) <= (layer0_outputs(2424)) xor (layer0_outputs(7452));
    outputs(379) <= layer0_outputs(10335);
    outputs(380) <= layer0_outputs(7239);
    outputs(381) <= not(layer0_outputs(5239));
    outputs(382) <= not((layer0_outputs(7675)) xor (layer0_outputs(12797)));
    outputs(383) <= layer0_outputs(4808);
    outputs(384) <= not((layer0_outputs(3268)) xor (layer0_outputs(8762)));
    outputs(385) <= layer0_outputs(7512);
    outputs(386) <= not(layer0_outputs(747));
    outputs(387) <= layer0_outputs(3389);
    outputs(388) <= not((layer0_outputs(7045)) or (layer0_outputs(470)));
    outputs(389) <= not(layer0_outputs(1724)) or (layer0_outputs(8169));
    outputs(390) <= (layer0_outputs(4569)) and (layer0_outputs(5026));
    outputs(391) <= layer0_outputs(8627);
    outputs(392) <= not((layer0_outputs(11788)) xor (layer0_outputs(11540)));
    outputs(393) <= (layer0_outputs(11422)) and not (layer0_outputs(5630));
    outputs(394) <= (layer0_outputs(4644)) xor (layer0_outputs(10326));
    outputs(395) <= layer0_outputs(8129);
    outputs(396) <= (layer0_outputs(4018)) xor (layer0_outputs(8706));
    outputs(397) <= not(layer0_outputs(1591)) or (layer0_outputs(9866));
    outputs(398) <= (layer0_outputs(12082)) xor (layer0_outputs(724));
    outputs(399) <= (layer0_outputs(10829)) xor (layer0_outputs(6724));
    outputs(400) <= (layer0_outputs(796)) xor (layer0_outputs(1974));
    outputs(401) <= not(layer0_outputs(7407));
    outputs(402) <= (layer0_outputs(11051)) xor (layer0_outputs(3452));
    outputs(403) <= not(layer0_outputs(613));
    outputs(404) <= not(layer0_outputs(8176));
    outputs(405) <= layer0_outputs(7936);
    outputs(406) <= not(layer0_outputs(1849));
    outputs(407) <= not(layer0_outputs(6688));
    outputs(408) <= layer0_outputs(5505);
    outputs(409) <= (layer0_outputs(4263)) xor (layer0_outputs(166));
    outputs(410) <= layer0_outputs(11370);
    outputs(411) <= not(layer0_outputs(8237)) or (layer0_outputs(10449));
    outputs(412) <= not(layer0_outputs(12499));
    outputs(413) <= layer0_outputs(1442);
    outputs(414) <= not(layer0_outputs(2470));
    outputs(415) <= (layer0_outputs(10953)) and not (layer0_outputs(8714));
    outputs(416) <= not((layer0_outputs(8332)) xor (layer0_outputs(4743)));
    outputs(417) <= (layer0_outputs(10640)) or (layer0_outputs(268));
    outputs(418) <= not(layer0_outputs(8378));
    outputs(419) <= not(layer0_outputs(756)) or (layer0_outputs(11826));
    outputs(420) <= (layer0_outputs(2869)) xor (layer0_outputs(12797));
    outputs(421) <= (layer0_outputs(2484)) and not (layer0_outputs(10159));
    outputs(422) <= (layer0_outputs(10972)) xor (layer0_outputs(11176));
    outputs(423) <= not((layer0_outputs(12789)) xor (layer0_outputs(8519)));
    outputs(424) <= (layer0_outputs(9755)) xor (layer0_outputs(5524));
    outputs(425) <= not(layer0_outputs(7195));
    outputs(426) <= (layer0_outputs(12247)) xor (layer0_outputs(4270));
    outputs(427) <= not(layer0_outputs(9838));
    outputs(428) <= not((layer0_outputs(8723)) xor (layer0_outputs(4471)));
    outputs(429) <= layer0_outputs(699);
    outputs(430) <= not(layer0_outputs(8443)) or (layer0_outputs(8062));
    outputs(431) <= layer0_outputs(7873);
    outputs(432) <= not(layer0_outputs(1486));
    outputs(433) <= not(layer0_outputs(989));
    outputs(434) <= not(layer0_outputs(4755));
    outputs(435) <= not(layer0_outputs(8319));
    outputs(436) <= (layer0_outputs(8837)) xor (layer0_outputs(7036));
    outputs(437) <= not((layer0_outputs(8786)) xor (layer0_outputs(11184)));
    outputs(438) <= layer0_outputs(6058);
    outputs(439) <= layer0_outputs(414);
    outputs(440) <= not(layer0_outputs(9540));
    outputs(441) <= (layer0_outputs(5475)) xor (layer0_outputs(4535));
    outputs(442) <= (layer0_outputs(2602)) xor (layer0_outputs(1769));
    outputs(443) <= (layer0_outputs(10571)) xor (layer0_outputs(2704));
    outputs(444) <= (layer0_outputs(6744)) xor (layer0_outputs(6800));
    outputs(445) <= not((layer0_outputs(2273)) xor (layer0_outputs(11363)));
    outputs(446) <= (layer0_outputs(11220)) xor (layer0_outputs(7550));
    outputs(447) <= not((layer0_outputs(12398)) and (layer0_outputs(11159)));
    outputs(448) <= not((layer0_outputs(11265)) and (layer0_outputs(11951)));
    outputs(449) <= not(layer0_outputs(9174));
    outputs(450) <= not(layer0_outputs(11918));
    outputs(451) <= not(layer0_outputs(3280));
    outputs(452) <= not(layer0_outputs(437));
    outputs(453) <= not(layer0_outputs(5225));
    outputs(454) <= not(layer0_outputs(6664)) or (layer0_outputs(8019));
    outputs(455) <= (layer0_outputs(2720)) and not (layer0_outputs(9242));
    outputs(456) <= layer0_outputs(1893);
    outputs(457) <= not((layer0_outputs(9556)) and (layer0_outputs(11733)));
    outputs(458) <= layer0_outputs(501);
    outputs(459) <= not(layer0_outputs(11472));
    outputs(460) <= (layer0_outputs(11311)) or (layer0_outputs(4708));
    outputs(461) <= (layer0_outputs(7978)) and not (layer0_outputs(3610));
    outputs(462) <= layer0_outputs(2835);
    outputs(463) <= not(layer0_outputs(8783));
    outputs(464) <= not(layer0_outputs(12010));
    outputs(465) <= layer0_outputs(3651);
    outputs(466) <= layer0_outputs(9893);
    outputs(467) <= (layer0_outputs(10416)) xor (layer0_outputs(296));
    outputs(468) <= not((layer0_outputs(5733)) xor (layer0_outputs(2786)));
    outputs(469) <= not(layer0_outputs(8207));
    outputs(470) <= layer0_outputs(4651);
    outputs(471) <= (layer0_outputs(10660)) xor (layer0_outputs(799));
    outputs(472) <= not((layer0_outputs(7639)) xor (layer0_outputs(9903)));
    outputs(473) <= (layer0_outputs(12569)) xor (layer0_outputs(9915));
    outputs(474) <= not(layer0_outputs(8162));
    outputs(475) <= not(layer0_outputs(3712));
    outputs(476) <= not((layer0_outputs(12102)) xor (layer0_outputs(3387)));
    outputs(477) <= layer0_outputs(4957);
    outputs(478) <= not((layer0_outputs(12366)) and (layer0_outputs(5483)));
    outputs(479) <= not((layer0_outputs(8632)) xor (layer0_outputs(5659)));
    outputs(480) <= (layer0_outputs(8340)) and not (layer0_outputs(12343));
    outputs(481) <= not((layer0_outputs(4020)) xor (layer0_outputs(6437)));
    outputs(482) <= (layer0_outputs(12776)) and (layer0_outputs(4080));
    outputs(483) <= (layer0_outputs(6255)) xor (layer0_outputs(4244));
    outputs(484) <= not((layer0_outputs(6247)) xor (layer0_outputs(3717)));
    outputs(485) <= not((layer0_outputs(5954)) xor (layer0_outputs(187)));
    outputs(486) <= layer0_outputs(5193);
    outputs(487) <= (layer0_outputs(10651)) xor (layer0_outputs(7850));
    outputs(488) <= not((layer0_outputs(3275)) xor (layer0_outputs(6022)));
    outputs(489) <= not((layer0_outputs(3636)) xor (layer0_outputs(9465)));
    outputs(490) <= not(layer0_outputs(6829));
    outputs(491) <= layer0_outputs(2780);
    outputs(492) <= not(layer0_outputs(9947));
    outputs(493) <= not(layer0_outputs(2912));
    outputs(494) <= not((layer0_outputs(5679)) or (layer0_outputs(4642)));
    outputs(495) <= layer0_outputs(4315);
    outputs(496) <= not(layer0_outputs(10066));
    outputs(497) <= not(layer0_outputs(12768));
    outputs(498) <= not(layer0_outputs(1110)) or (layer0_outputs(4540));
    outputs(499) <= not(layer0_outputs(8389));
    outputs(500) <= (layer0_outputs(4411)) and not (layer0_outputs(5060));
    outputs(501) <= not((layer0_outputs(2787)) xor (layer0_outputs(8003)));
    outputs(502) <= (layer0_outputs(5047)) xor (layer0_outputs(4701));
    outputs(503) <= not(layer0_outputs(8962));
    outputs(504) <= not(layer0_outputs(2275));
    outputs(505) <= not(layer0_outputs(7225));
    outputs(506) <= not(layer0_outputs(12599));
    outputs(507) <= (layer0_outputs(6171)) and not (layer0_outputs(6947));
    outputs(508) <= not(layer0_outputs(3823));
    outputs(509) <= not(layer0_outputs(178));
    outputs(510) <= not((layer0_outputs(10226)) xor (layer0_outputs(3327)));
    outputs(511) <= not((layer0_outputs(5024)) xor (layer0_outputs(11187)));
    outputs(512) <= not(layer0_outputs(1492));
    outputs(513) <= not((layer0_outputs(235)) and (layer0_outputs(3781)));
    outputs(514) <= not(layer0_outputs(9551)) or (layer0_outputs(1868));
    outputs(515) <= layer0_outputs(11698);
    outputs(516) <= not(layer0_outputs(774));
    outputs(517) <= not((layer0_outputs(1280)) and (layer0_outputs(5181)));
    outputs(518) <= not((layer0_outputs(3839)) xor (layer0_outputs(526)));
    outputs(519) <= not((layer0_outputs(244)) or (layer0_outputs(9845)));
    outputs(520) <= layer0_outputs(8982);
    outputs(521) <= layer0_outputs(1114);
    outputs(522) <= layer0_outputs(5254);
    outputs(523) <= (layer0_outputs(3253)) xor (layer0_outputs(10695));
    outputs(524) <= not((layer0_outputs(3629)) xor (layer0_outputs(7952)));
    outputs(525) <= layer0_outputs(1213);
    outputs(526) <= not((layer0_outputs(6129)) and (layer0_outputs(4416)));
    outputs(527) <= not(layer0_outputs(5433)) or (layer0_outputs(7578));
    outputs(528) <= not(layer0_outputs(2126)) or (layer0_outputs(4648));
    outputs(529) <= not((layer0_outputs(2722)) xor (layer0_outputs(2788)));
    outputs(530) <= layer0_outputs(1682);
    outputs(531) <= (layer0_outputs(7521)) xor (layer0_outputs(9570));
    outputs(532) <= not((layer0_outputs(4539)) xor (layer0_outputs(10914)));
    outputs(533) <= not(layer0_outputs(9737));
    outputs(534) <= (layer0_outputs(9065)) or (layer0_outputs(3974));
    outputs(535) <= not(layer0_outputs(5111));
    outputs(536) <= (layer0_outputs(1997)) and (layer0_outputs(10841));
    outputs(537) <= not((layer0_outputs(6178)) and (layer0_outputs(12115)));
    outputs(538) <= layer0_outputs(6982);
    outputs(539) <= layer0_outputs(10179);
    outputs(540) <= not((layer0_outputs(1356)) xor (layer0_outputs(2963)));
    outputs(541) <= (layer0_outputs(2298)) xor (layer0_outputs(11652));
    outputs(542) <= layer0_outputs(7468);
    outputs(543) <= layer0_outputs(923);
    outputs(544) <= not((layer0_outputs(7695)) xor (layer0_outputs(9263)));
    outputs(545) <= layer0_outputs(12626);
    outputs(546) <= not((layer0_outputs(5315)) xor (layer0_outputs(10777)));
    outputs(547) <= (layer0_outputs(4413)) xor (layer0_outputs(2906));
    outputs(548) <= not((layer0_outputs(5707)) or (layer0_outputs(3728)));
    outputs(549) <= (layer0_outputs(2750)) xor (layer0_outputs(12290));
    outputs(550) <= (layer0_outputs(5899)) xor (layer0_outputs(7858));
    outputs(551) <= not(layer0_outputs(517));
    outputs(552) <= (layer0_outputs(7557)) xor (layer0_outputs(7610));
    outputs(553) <= not(layer0_outputs(2831)) or (layer0_outputs(1464));
    outputs(554) <= layer0_outputs(8837);
    outputs(555) <= layer0_outputs(4253);
    outputs(556) <= not((layer0_outputs(11450)) xor (layer0_outputs(11888)));
    outputs(557) <= layer0_outputs(12329);
    outputs(558) <= not(layer0_outputs(8253));
    outputs(559) <= not(layer0_outputs(9355));
    outputs(560) <= layer0_outputs(7898);
    outputs(561) <= not((layer0_outputs(6356)) xor (layer0_outputs(863)));
    outputs(562) <= (layer0_outputs(10370)) and (layer0_outputs(2905));
    outputs(563) <= not((layer0_outputs(3955)) xor (layer0_outputs(12724)));
    outputs(564) <= layer0_outputs(10672);
    outputs(565) <= layer0_outputs(4766);
    outputs(566) <= layer0_outputs(3072);
    outputs(567) <= layer0_outputs(5677);
    outputs(568) <= not((layer0_outputs(1430)) and (layer0_outputs(10084)));
    outputs(569) <= not(layer0_outputs(3966));
    outputs(570) <= layer0_outputs(9435);
    outputs(571) <= not(layer0_outputs(933));
    outputs(572) <= not(layer0_outputs(8722)) or (layer0_outputs(3856));
    outputs(573) <= layer0_outputs(4336);
    outputs(574) <= layer0_outputs(10770);
    outputs(575) <= (layer0_outputs(5947)) xor (layer0_outputs(10992));
    outputs(576) <= layer0_outputs(2629);
    outputs(577) <= not(layer0_outputs(4993));
    outputs(578) <= not(layer0_outputs(4075));
    outputs(579) <= (layer0_outputs(8788)) and not (layer0_outputs(7349));
    outputs(580) <= not(layer0_outputs(6832)) or (layer0_outputs(6804));
    outputs(581) <= layer0_outputs(5474);
    outputs(582) <= (layer0_outputs(4342)) or (layer0_outputs(2461));
    outputs(583) <= (layer0_outputs(2797)) and (layer0_outputs(941));
    outputs(584) <= (layer0_outputs(4605)) xor (layer0_outputs(1098));
    outputs(585) <= not(layer0_outputs(8370)) or (layer0_outputs(12591));
    outputs(586) <= not((layer0_outputs(7052)) and (layer0_outputs(2175)));
    outputs(587) <= (layer0_outputs(890)) xor (layer0_outputs(12734));
    outputs(588) <= not(layer0_outputs(3633));
    outputs(589) <= (layer0_outputs(3828)) and (layer0_outputs(5758));
    outputs(590) <= not(layer0_outputs(12312));
    outputs(591) <= not(layer0_outputs(7088));
    outputs(592) <= layer0_outputs(5196);
    outputs(593) <= layer0_outputs(6113);
    outputs(594) <= not(layer0_outputs(602));
    outputs(595) <= not(layer0_outputs(968));
    outputs(596) <= (layer0_outputs(6626)) and not (layer0_outputs(2095));
    outputs(597) <= (layer0_outputs(11194)) xor (layer0_outputs(7578));
    outputs(598) <= (layer0_outputs(1306)) and (layer0_outputs(3719));
    outputs(599) <= not((layer0_outputs(11118)) xor (layer0_outputs(6157)));
    outputs(600) <= not(layer0_outputs(5158));
    outputs(601) <= (layer0_outputs(12056)) and not (layer0_outputs(6703));
    outputs(602) <= not(layer0_outputs(9870));
    outputs(603) <= not(layer0_outputs(10331));
    outputs(604) <= layer0_outputs(7860);
    outputs(605) <= (layer0_outputs(8312)) and not (layer0_outputs(6805));
    outputs(606) <= not((layer0_outputs(4153)) xor (layer0_outputs(5485)));
    outputs(607) <= (layer0_outputs(8479)) or (layer0_outputs(379));
    outputs(608) <= (layer0_outputs(1619)) xor (layer0_outputs(1530));
    outputs(609) <= not(layer0_outputs(6880));
    outputs(610) <= not(layer0_outputs(3818));
    outputs(611) <= layer0_outputs(8033);
    outputs(612) <= not((layer0_outputs(5994)) or (layer0_outputs(3718)));
    outputs(613) <= not(layer0_outputs(9495));
    outputs(614) <= (layer0_outputs(4861)) xor (layer0_outputs(1840));
    outputs(615) <= not(layer0_outputs(9495));
    outputs(616) <= not((layer0_outputs(10714)) xor (layer0_outputs(12298)));
    outputs(617) <= (layer0_outputs(7133)) and not (layer0_outputs(4830));
    outputs(618) <= (layer0_outputs(74)) and (layer0_outputs(7682));
    outputs(619) <= (layer0_outputs(9581)) and not (layer0_outputs(8370));
    outputs(620) <= (layer0_outputs(6869)) xor (layer0_outputs(2205));
    outputs(621) <= layer0_outputs(8969);
    outputs(622) <= not(layer0_outputs(10269));
    outputs(623) <= layer0_outputs(2001);
    outputs(624) <= (layer0_outputs(4834)) and not (layer0_outputs(5378));
    outputs(625) <= layer0_outputs(7856);
    outputs(626) <= (layer0_outputs(8566)) xor (layer0_outputs(6080));
    outputs(627) <= not(layer0_outputs(7791)) or (layer0_outputs(1923));
    outputs(628) <= (layer0_outputs(4389)) xor (layer0_outputs(12644));
    outputs(629) <= layer0_outputs(5493);
    outputs(630) <= not((layer0_outputs(1247)) xor (layer0_outputs(9035)));
    outputs(631) <= layer0_outputs(1725);
    outputs(632) <= layer0_outputs(1913);
    outputs(633) <= (layer0_outputs(1526)) xor (layer0_outputs(12703));
    outputs(634) <= (layer0_outputs(9603)) or (layer0_outputs(10002));
    outputs(635) <= (layer0_outputs(10738)) xor (layer0_outputs(3320));
    outputs(636) <= (layer0_outputs(8504)) xor (layer0_outputs(8910));
    outputs(637) <= not((layer0_outputs(12142)) and (layer0_outputs(7186)));
    outputs(638) <= not((layer0_outputs(11185)) xor (layer0_outputs(931)));
    outputs(639) <= not(layer0_outputs(2563));
    outputs(640) <= not(layer0_outputs(7394));
    outputs(641) <= (layer0_outputs(5108)) and (layer0_outputs(10991));
    outputs(642) <= (layer0_outputs(5816)) and not (layer0_outputs(8235));
    outputs(643) <= layer0_outputs(5354);
    outputs(644) <= not(layer0_outputs(1354));
    outputs(645) <= not((layer0_outputs(8320)) xor (layer0_outputs(692)));
    outputs(646) <= layer0_outputs(8921);
    outputs(647) <= not((layer0_outputs(12405)) and (layer0_outputs(8783)));
    outputs(648) <= not(layer0_outputs(2446));
    outputs(649) <= layer0_outputs(7856);
    outputs(650) <= not((layer0_outputs(10059)) and (layer0_outputs(1400)));
    outputs(651) <= layer0_outputs(3219);
    outputs(652) <= not(layer0_outputs(1920));
    outputs(653) <= not(layer0_outputs(5526)) or (layer0_outputs(4499));
    outputs(654) <= not(layer0_outputs(3894));
    outputs(655) <= layer0_outputs(7211);
    outputs(656) <= layer0_outputs(10701);
    outputs(657) <= (layer0_outputs(3088)) xor (layer0_outputs(7610));
    outputs(658) <= not(layer0_outputs(1611)) or (layer0_outputs(1146));
    outputs(659) <= (layer0_outputs(1972)) xor (layer0_outputs(6210));
    outputs(660) <= (layer0_outputs(2736)) and not (layer0_outputs(5660));
    outputs(661) <= layer0_outputs(4190);
    outputs(662) <= (layer0_outputs(6211)) xor (layer0_outputs(8921));
    outputs(663) <= layer0_outputs(2397);
    outputs(664) <= not(layer0_outputs(1791)) or (layer0_outputs(4368));
    outputs(665) <= not(layer0_outputs(12791));
    outputs(666) <= layer0_outputs(5859);
    outputs(667) <= layer0_outputs(7692);
    outputs(668) <= layer0_outputs(8987);
    outputs(669) <= not(layer0_outputs(3295));
    outputs(670) <= not(layer0_outputs(2454)) or (layer0_outputs(12565));
    outputs(671) <= layer0_outputs(2028);
    outputs(672) <= not((layer0_outputs(1804)) or (layer0_outputs(10287)));
    outputs(673) <= (layer0_outputs(8735)) xor (layer0_outputs(2178));
    outputs(674) <= not(layer0_outputs(9354));
    outputs(675) <= layer0_outputs(4851);
    outputs(676) <= layer0_outputs(7040);
    outputs(677) <= not(layer0_outputs(3540));
    outputs(678) <= not((layer0_outputs(7988)) and (layer0_outputs(9566)));
    outputs(679) <= not((layer0_outputs(372)) xor (layer0_outputs(2364)));
    outputs(680) <= not((layer0_outputs(917)) and (layer0_outputs(11493)));
    outputs(681) <= layer0_outputs(3668);
    outputs(682) <= (layer0_outputs(7563)) and not (layer0_outputs(10667));
    outputs(683) <= not((layer0_outputs(6733)) or (layer0_outputs(6419)));
    outputs(684) <= not(layer0_outputs(2814));
    outputs(685) <= not((layer0_outputs(7087)) or (layer0_outputs(5596)));
    outputs(686) <= not(layer0_outputs(11250));
    outputs(687) <= not((layer0_outputs(11707)) xor (layer0_outputs(3062)));
    outputs(688) <= (layer0_outputs(6528)) and (layer0_outputs(10343));
    outputs(689) <= not((layer0_outputs(6961)) xor (layer0_outputs(11149)));
    outputs(690) <= layer0_outputs(11527);
    outputs(691) <= not((layer0_outputs(8482)) xor (layer0_outputs(4053)));
    outputs(692) <= not((layer0_outputs(10642)) or (layer0_outputs(10952)));
    outputs(693) <= not(layer0_outputs(12489));
    outputs(694) <= not(layer0_outputs(6946)) or (layer0_outputs(9981));
    outputs(695) <= layer0_outputs(2026);
    outputs(696) <= not((layer0_outputs(11915)) xor (layer0_outputs(1145)));
    outputs(697) <= not((layer0_outputs(9478)) or (layer0_outputs(10623)));
    outputs(698) <= layer0_outputs(11427);
    outputs(699) <= not(layer0_outputs(4888));
    outputs(700) <= layer0_outputs(9509);
    outputs(701) <= not(layer0_outputs(3013));
    outputs(702) <= not((layer0_outputs(3271)) and (layer0_outputs(5630)));
    outputs(703) <= (layer0_outputs(4046)) xor (layer0_outputs(9762));
    outputs(704) <= layer0_outputs(7674);
    outputs(705) <= not((layer0_outputs(7236)) xor (layer0_outputs(8519)));
    outputs(706) <= (layer0_outputs(6397)) xor (layer0_outputs(8335));
    outputs(707) <= (layer0_outputs(2548)) and (layer0_outputs(8952));
    outputs(708) <= not((layer0_outputs(9771)) or (layer0_outputs(6170)));
    outputs(709) <= (layer0_outputs(10853)) xor (layer0_outputs(10013));
    outputs(710) <= not(layer0_outputs(2021)) or (layer0_outputs(1519));
    outputs(711) <= not((layer0_outputs(8168)) xor (layer0_outputs(11986)));
    outputs(712) <= (layer0_outputs(492)) and not (layer0_outputs(3498));
    outputs(713) <= not(layer0_outputs(953));
    outputs(714) <= (layer0_outputs(1698)) or (layer0_outputs(4785));
    outputs(715) <= not(layer0_outputs(5417)) or (layer0_outputs(913));
    outputs(716) <= layer0_outputs(9496);
    outputs(717) <= not((layer0_outputs(2387)) and (layer0_outputs(1261)));
    outputs(718) <= (layer0_outputs(6180)) and not (layer0_outputs(966));
    outputs(719) <= layer0_outputs(10281);
    outputs(720) <= not((layer0_outputs(10918)) xor (layer0_outputs(9747)));
    outputs(721) <= (layer0_outputs(10320)) xor (layer0_outputs(6176));
    outputs(722) <= not(layer0_outputs(2648)) or (layer0_outputs(522));
    outputs(723) <= not(layer0_outputs(11028));
    outputs(724) <= not(layer0_outputs(10845));
    outputs(725) <= not(layer0_outputs(1908));
    outputs(726) <= layer0_outputs(7184);
    outputs(727) <= not((layer0_outputs(6953)) xor (layer0_outputs(4777)));
    outputs(728) <= (layer0_outputs(6590)) and not (layer0_outputs(7676));
    outputs(729) <= (layer0_outputs(11377)) xor (layer0_outputs(10780));
    outputs(730) <= not(layer0_outputs(11795));
    outputs(731) <= layer0_outputs(6228);
    outputs(732) <= not((layer0_outputs(1583)) and (layer0_outputs(2651)));
    outputs(733) <= not((layer0_outputs(7454)) xor (layer0_outputs(516)));
    outputs(734) <= (layer0_outputs(495)) and not (layer0_outputs(9567));
    outputs(735) <= not(layer0_outputs(6643)) or (layer0_outputs(8965));
    outputs(736) <= not((layer0_outputs(4294)) or (layer0_outputs(5337)));
    outputs(737) <= (layer0_outputs(11235)) and (layer0_outputs(1114));
    outputs(738) <= not((layer0_outputs(9728)) and (layer0_outputs(6596)));
    outputs(739) <= (layer0_outputs(1229)) and (layer0_outputs(6389));
    outputs(740) <= (layer0_outputs(9541)) and not (layer0_outputs(1131));
    outputs(741) <= not(layer0_outputs(2620)) or (layer0_outputs(10702));
    outputs(742) <= layer0_outputs(2553);
    outputs(743) <= (layer0_outputs(12060)) xor (layer0_outputs(939));
    outputs(744) <= (layer0_outputs(4300)) and (layer0_outputs(3426));
    outputs(745) <= not(layer0_outputs(7686));
    outputs(746) <= layer0_outputs(1596);
    outputs(747) <= not(layer0_outputs(4847));
    outputs(748) <= not((layer0_outputs(12097)) xor (layer0_outputs(10715)));
    outputs(749) <= not(layer0_outputs(3296));
    outputs(750) <= not((layer0_outputs(12603)) or (layer0_outputs(9092)));
    outputs(751) <= (layer0_outputs(10259)) xor (layer0_outputs(5771));
    outputs(752) <= not(layer0_outputs(855));
    outputs(753) <= not(layer0_outputs(9168));
    outputs(754) <= not((layer0_outputs(10153)) xor (layer0_outputs(12571)));
    outputs(755) <= layer0_outputs(10094);
    outputs(756) <= (layer0_outputs(3641)) or (layer0_outputs(62));
    outputs(757) <= not((layer0_outputs(10499)) xor (layer0_outputs(1219)));
    outputs(758) <= not((layer0_outputs(12211)) or (layer0_outputs(2378)));
    outputs(759) <= not((layer0_outputs(8653)) xor (layer0_outputs(9751)));
    outputs(760) <= not(layer0_outputs(6000));
    outputs(761) <= not((layer0_outputs(5416)) and (layer0_outputs(8832)));
    outputs(762) <= (layer0_outputs(10015)) xor (layer0_outputs(7615));
    outputs(763) <= layer0_outputs(5112);
    outputs(764) <= (layer0_outputs(6265)) and (layer0_outputs(5094));
    outputs(765) <= layer0_outputs(9487);
    outputs(766) <= not((layer0_outputs(723)) xor (layer0_outputs(2200)));
    outputs(767) <= layer0_outputs(1654);
    outputs(768) <= layer0_outputs(11698);
    outputs(769) <= not(layer0_outputs(47));
    outputs(770) <= (layer0_outputs(11016)) xor (layer0_outputs(1994));
    outputs(771) <= (layer0_outputs(10383)) or (layer0_outputs(9577));
    outputs(772) <= not(layer0_outputs(11044));
    outputs(773) <= not(layer0_outputs(3644));
    outputs(774) <= not((layer0_outputs(7118)) xor (layer0_outputs(10934)));
    outputs(775) <= not(layer0_outputs(3833));
    outputs(776) <= (layer0_outputs(3423)) xor (layer0_outputs(10584));
    outputs(777) <= not(layer0_outputs(12142)) or (layer0_outputs(11141));
    outputs(778) <= not(layer0_outputs(7766)) or (layer0_outputs(11391));
    outputs(779) <= layer0_outputs(5777);
    outputs(780) <= not(layer0_outputs(6141));
    outputs(781) <= not((layer0_outputs(5118)) xor (layer0_outputs(3857)));
    outputs(782) <= (layer0_outputs(1870)) and (layer0_outputs(6270));
    outputs(783) <= not((layer0_outputs(11766)) and (layer0_outputs(2897)));
    outputs(784) <= not((layer0_outputs(9296)) and (layer0_outputs(299)));
    outputs(785) <= not(layer0_outputs(8943));
    outputs(786) <= not((layer0_outputs(9953)) xor (layer0_outputs(12610)));
    outputs(787) <= not((layer0_outputs(9149)) xor (layer0_outputs(10130)));
    outputs(788) <= (layer0_outputs(153)) xor (layer0_outputs(2640));
    outputs(789) <= not(layer0_outputs(2187));
    outputs(790) <= not((layer0_outputs(4495)) and (layer0_outputs(6987)));
    outputs(791) <= layer0_outputs(7857);
    outputs(792) <= layer0_outputs(12463);
    outputs(793) <= not(layer0_outputs(8576)) or (layer0_outputs(11287));
    outputs(794) <= (layer0_outputs(3236)) and not (layer0_outputs(372));
    outputs(795) <= (layer0_outputs(11552)) and not (layer0_outputs(5639));
    outputs(796) <= not(layer0_outputs(2092));
    outputs(797) <= not(layer0_outputs(2489));
    outputs(798) <= layer0_outputs(3569);
    outputs(799) <= not(layer0_outputs(2904));
    outputs(800) <= layer0_outputs(3007);
    outputs(801) <= layer0_outputs(9239);
    outputs(802) <= not(layer0_outputs(3133));
    outputs(803) <= layer0_outputs(4128);
    outputs(804) <= not(layer0_outputs(9246));
    outputs(805) <= not((layer0_outputs(8513)) xor (layer0_outputs(3708)));
    outputs(806) <= not(layer0_outputs(9027));
    outputs(807) <= layer0_outputs(9382);
    outputs(808) <= (layer0_outputs(1647)) and (layer0_outputs(2342));
    outputs(809) <= (layer0_outputs(7661)) and not (layer0_outputs(2433));
    outputs(810) <= (layer0_outputs(10784)) and (layer0_outputs(2769));
    outputs(811) <= layer0_outputs(8730);
    outputs(812) <= not(layer0_outputs(1511));
    outputs(813) <= (layer0_outputs(7948)) xor (layer0_outputs(1774));
    outputs(814) <= not(layer0_outputs(746));
    outputs(815) <= layer0_outputs(12253);
    outputs(816) <= (layer0_outputs(7193)) xor (layer0_outputs(166));
    outputs(817) <= (layer0_outputs(6257)) and not (layer0_outputs(6861));
    outputs(818) <= not((layer0_outputs(8075)) xor (layer0_outputs(5365)));
    outputs(819) <= layer0_outputs(1722);
    outputs(820) <= not((layer0_outputs(1441)) and (layer0_outputs(403)));
    outputs(821) <= (layer0_outputs(9509)) and (layer0_outputs(10731));
    outputs(822) <= not(layer0_outputs(11799));
    outputs(823) <= not((layer0_outputs(2951)) xor (layer0_outputs(5227)));
    outputs(824) <= not((layer0_outputs(1296)) and (layer0_outputs(1665)));
    outputs(825) <= layer0_outputs(12067);
    outputs(826) <= not((layer0_outputs(2288)) xor (layer0_outputs(5870)));
    outputs(827) <= (layer0_outputs(4865)) xor (layer0_outputs(3975));
    outputs(828) <= (layer0_outputs(3094)) xor (layer0_outputs(8654));
    outputs(829) <= (layer0_outputs(2047)) xor (layer0_outputs(6821));
    outputs(830) <= (layer0_outputs(6631)) xor (layer0_outputs(10314));
    outputs(831) <= not(layer0_outputs(1164));
    outputs(832) <= not((layer0_outputs(11506)) xor (layer0_outputs(5220)));
    outputs(833) <= not(layer0_outputs(5298));
    outputs(834) <= (layer0_outputs(11555)) xor (layer0_outputs(3083));
    outputs(835) <= not((layer0_outputs(1159)) xor (layer0_outputs(2491)));
    outputs(836) <= not(layer0_outputs(12106));
    outputs(837) <= layer0_outputs(6296);
    outputs(838) <= (layer0_outputs(1570)) xor (layer0_outputs(10758));
    outputs(839) <= not((layer0_outputs(5194)) xor (layer0_outputs(2966)));
    outputs(840) <= not((layer0_outputs(11742)) xor (layer0_outputs(2429)));
    outputs(841) <= (layer0_outputs(10121)) xor (layer0_outputs(12247));
    outputs(842) <= '1';
    outputs(843) <= layer0_outputs(7289);
    outputs(844) <= layer0_outputs(2802);
    outputs(845) <= not((layer0_outputs(9182)) xor (layer0_outputs(2044)));
    outputs(846) <= layer0_outputs(10472);
    outputs(847) <= layer0_outputs(8835);
    outputs(848) <= (layer0_outputs(7238)) and (layer0_outputs(7905));
    outputs(849) <= not(layer0_outputs(552));
    outputs(850) <= (layer0_outputs(7438)) or (layer0_outputs(11863));
    outputs(851) <= not(layer0_outputs(6834));
    outputs(852) <= not(layer0_outputs(233));
    outputs(853) <= (layer0_outputs(1160)) xor (layer0_outputs(6597));
    outputs(854) <= layer0_outputs(11703);
    outputs(855) <= not(layer0_outputs(9276));
    outputs(856) <= not(layer0_outputs(5535)) or (layer0_outputs(7929));
    outputs(857) <= layer0_outputs(12233);
    outputs(858) <= layer0_outputs(5052);
    outputs(859) <= layer0_outputs(9948);
    outputs(860) <= layer0_outputs(1030);
    outputs(861) <= (layer0_outputs(10773)) xor (layer0_outputs(10082));
    outputs(862) <= not(layer0_outputs(4102));
    outputs(863) <= (layer0_outputs(6838)) xor (layer0_outputs(3561));
    outputs(864) <= (layer0_outputs(3543)) xor (layer0_outputs(511));
    outputs(865) <= not(layer0_outputs(3006));
    outputs(866) <= (layer0_outputs(6639)) and not (layer0_outputs(97));
    outputs(867) <= not(layer0_outputs(10659));
    outputs(868) <= (layer0_outputs(2861)) or (layer0_outputs(7253));
    outputs(869) <= layer0_outputs(5570);
    outputs(870) <= not(layer0_outputs(1091)) or (layer0_outputs(1793));
    outputs(871) <= not(layer0_outputs(2070));
    outputs(872) <= not(layer0_outputs(5492)) or (layer0_outputs(295));
    outputs(873) <= layer0_outputs(4306);
    outputs(874) <= not(layer0_outputs(3322));
    outputs(875) <= not((layer0_outputs(2708)) xor (layer0_outputs(2364)));
    outputs(876) <= (layer0_outputs(12579)) and not (layer0_outputs(10182));
    outputs(877) <= not(layer0_outputs(631)) or (layer0_outputs(4303));
    outputs(878) <= layer0_outputs(10488);
    outputs(879) <= (layer0_outputs(11852)) xor (layer0_outputs(9667));
    outputs(880) <= layer0_outputs(7831);
    outputs(881) <= layer0_outputs(1331);
    outputs(882) <= not(layer0_outputs(1991)) or (layer0_outputs(9700));
    outputs(883) <= layer0_outputs(7530);
    outputs(884) <= not(layer0_outputs(7932));
    outputs(885) <= not(layer0_outputs(4382)) or (layer0_outputs(10576));
    outputs(886) <= not((layer0_outputs(7824)) xor (layer0_outputs(1696)));
    outputs(887) <= not((layer0_outputs(5384)) xor (layer0_outputs(6626)));
    outputs(888) <= not(layer0_outputs(9221));
    outputs(889) <= not((layer0_outputs(4806)) xor (layer0_outputs(4739)));
    outputs(890) <= not((layer0_outputs(7246)) xor (layer0_outputs(5693)));
    outputs(891) <= layer0_outputs(1736);
    outputs(892) <= (layer0_outputs(3010)) and not (layer0_outputs(6443));
    outputs(893) <= not(layer0_outputs(8681));
    outputs(894) <= layer0_outputs(6731);
    outputs(895) <= not(layer0_outputs(10900)) or (layer0_outputs(3065));
    outputs(896) <= (layer0_outputs(2557)) xor (layer0_outputs(11648));
    outputs(897) <= layer0_outputs(9059);
    outputs(898) <= layer0_outputs(3803);
    outputs(899) <= (layer0_outputs(9488)) and not (layer0_outputs(12399));
    outputs(900) <= not(layer0_outputs(1953));
    outputs(901) <= not(layer0_outputs(8958));
    outputs(902) <= not(layer0_outputs(8042));
    outputs(903) <= not((layer0_outputs(11701)) and (layer0_outputs(12561)));
    outputs(904) <= layer0_outputs(9992);
    outputs(905) <= layer0_outputs(2848);
    outputs(906) <= not((layer0_outputs(4464)) xor (layer0_outputs(1456)));
    outputs(907) <= layer0_outputs(12428);
    outputs(908) <= not(layer0_outputs(1284));
    outputs(909) <= layer0_outputs(3238);
    outputs(910) <= layer0_outputs(10995);
    outputs(911) <= not((layer0_outputs(10682)) xor (layer0_outputs(417)));
    outputs(912) <= not(layer0_outputs(12195)) or (layer0_outputs(9650));
    outputs(913) <= not((layer0_outputs(790)) xor (layer0_outputs(7874)));
    outputs(914) <= layer0_outputs(3567);
    outputs(915) <= not(layer0_outputs(3133)) or (layer0_outputs(10116));
    outputs(916) <= not(layer0_outputs(7001));
    outputs(917) <= (layer0_outputs(3111)) and not (layer0_outputs(10324));
    outputs(918) <= (layer0_outputs(3675)) xor (layer0_outputs(7827));
    outputs(919) <= layer0_outputs(7230);
    outputs(920) <= not(layer0_outputs(6184));
    outputs(921) <= (layer0_outputs(4697)) xor (layer0_outputs(5608));
    outputs(922) <= (layer0_outputs(9320)) xor (layer0_outputs(4599));
    outputs(923) <= not(layer0_outputs(11807)) or (layer0_outputs(10762));
    outputs(924) <= layer0_outputs(3159);
    outputs(925) <= not(layer0_outputs(5670));
    outputs(926) <= not((layer0_outputs(12292)) xor (layer0_outputs(590)));
    outputs(927) <= not((layer0_outputs(4805)) xor (layer0_outputs(3278)));
    outputs(928) <= not((layer0_outputs(5439)) xor (layer0_outputs(4720)));
    outputs(929) <= (layer0_outputs(12091)) xor (layer0_outputs(3770));
    outputs(930) <= layer0_outputs(4997);
    outputs(931) <= (layer0_outputs(2998)) xor (layer0_outputs(748));
    outputs(932) <= (layer0_outputs(3578)) and not (layer0_outputs(938));
    outputs(933) <= (layer0_outputs(9823)) and not (layer0_outputs(11027));
    outputs(934) <= (layer0_outputs(8066)) xor (layer0_outputs(12719));
    outputs(935) <= not(layer0_outputs(11392));
    outputs(936) <= layer0_outputs(8474);
    outputs(937) <= not((layer0_outputs(7832)) or (layer0_outputs(3469)));
    outputs(938) <= layer0_outputs(6517);
    outputs(939) <= (layer0_outputs(6471)) xor (layer0_outputs(3953));
    outputs(940) <= not((layer0_outputs(3822)) xor (layer0_outputs(11139)));
    outputs(941) <= not(layer0_outputs(4632));
    outputs(942) <= (layer0_outputs(10602)) xor (layer0_outputs(7444));
    outputs(943) <= not(layer0_outputs(10254));
    outputs(944) <= not(layer0_outputs(4264)) or (layer0_outputs(1968));
    outputs(945) <= not((layer0_outputs(660)) xor (layer0_outputs(3464)));
    outputs(946) <= not((layer0_outputs(11974)) xor (layer0_outputs(4094)));
    outputs(947) <= not(layer0_outputs(10837));
    outputs(948) <= not(layer0_outputs(1143)) or (layer0_outputs(10072));
    outputs(949) <= not(layer0_outputs(6606)) or (layer0_outputs(12088));
    outputs(950) <= layer0_outputs(10965);
    outputs(951) <= not((layer0_outputs(6601)) or (layer0_outputs(862)));
    outputs(952) <= not(layer0_outputs(63));
    outputs(953) <= (layer0_outputs(11082)) xor (layer0_outputs(497));
    outputs(954) <= (layer0_outputs(1015)) xor (layer0_outputs(3669));
    outputs(955) <= layer0_outputs(9390);
    outputs(956) <= not((layer0_outputs(3811)) xor (layer0_outputs(12516)));
    outputs(957) <= not((layer0_outputs(7840)) xor (layer0_outputs(5224)));
    outputs(958) <= layer0_outputs(10696);
    outputs(959) <= (layer0_outputs(3425)) xor (layer0_outputs(11534));
    outputs(960) <= (layer0_outputs(6425)) and not (layer0_outputs(2371));
    outputs(961) <= (layer0_outputs(201)) xor (layer0_outputs(3881));
    outputs(962) <= (layer0_outputs(9803)) and not (layer0_outputs(11266));
    outputs(963) <= (layer0_outputs(12239)) xor (layer0_outputs(2217));
    outputs(964) <= (layer0_outputs(1926)) and not (layer0_outputs(2729));
    outputs(965) <= not(layer0_outputs(3554)) or (layer0_outputs(10087));
    outputs(966) <= layer0_outputs(12436);
    outputs(967) <= (layer0_outputs(12373)) and (layer0_outputs(185));
    outputs(968) <= not((layer0_outputs(7566)) xor (layer0_outputs(4770)));
    outputs(969) <= not((layer0_outputs(4819)) xor (layer0_outputs(1758)));
    outputs(970) <= not(layer0_outputs(879));
    outputs(971) <= not(layer0_outputs(1986));
    outputs(972) <= not((layer0_outputs(12494)) xor (layer0_outputs(6578)));
    outputs(973) <= not((layer0_outputs(335)) and (layer0_outputs(10474)));
    outputs(974) <= not(layer0_outputs(1393));
    outputs(975) <= (layer0_outputs(7096)) xor (layer0_outputs(3194));
    outputs(976) <= layer0_outputs(10398);
    outputs(977) <= not(layer0_outputs(11004));
    outputs(978) <= layer0_outputs(11870);
    outputs(979) <= not((layer0_outputs(7542)) and (layer0_outputs(3862)));
    outputs(980) <= (layer0_outputs(12544)) xor (layer0_outputs(3968));
    outputs(981) <= (layer0_outputs(4507)) or (layer0_outputs(8400));
    outputs(982) <= layer0_outputs(7670);
    outputs(983) <= layer0_outputs(726);
    outputs(984) <= not((layer0_outputs(7721)) and (layer0_outputs(2037)));
    outputs(985) <= not(layer0_outputs(12519)) or (layer0_outputs(7811));
    outputs(986) <= (layer0_outputs(5368)) xor (layer0_outputs(8464));
    outputs(987) <= not(layer0_outputs(765)) or (layer0_outputs(4842));
    outputs(988) <= not(layer0_outputs(1492));
    outputs(989) <= not(layer0_outputs(3740));
    outputs(990) <= not(layer0_outputs(10712));
    outputs(991) <= not(layer0_outputs(12027));
    outputs(992) <= not(layer0_outputs(92)) or (layer0_outputs(7333));
    outputs(993) <= not(layer0_outputs(1056)) or (layer0_outputs(5162));
    outputs(994) <= (layer0_outputs(815)) xor (layer0_outputs(9434));
    outputs(995) <= not(layer0_outputs(5444));
    outputs(996) <= layer0_outputs(6317);
    outputs(997) <= (layer0_outputs(1117)) xor (layer0_outputs(10270));
    outputs(998) <= layer0_outputs(6156);
    outputs(999) <= not(layer0_outputs(12493)) or (layer0_outputs(2524));
    outputs(1000) <= not((layer0_outputs(12728)) and (layer0_outputs(3457)));
    outputs(1001) <= layer0_outputs(5827);
    outputs(1002) <= (layer0_outputs(2013)) xor (layer0_outputs(5761));
    outputs(1003) <= (layer0_outputs(3390)) xor (layer0_outputs(8571));
    outputs(1004) <= (layer0_outputs(7998)) and not (layer0_outputs(5772));
    outputs(1005) <= not(layer0_outputs(2439));
    outputs(1006) <= (layer0_outputs(9388)) and (layer0_outputs(12049));
    outputs(1007) <= layer0_outputs(10421);
    outputs(1008) <= not((layer0_outputs(37)) xor (layer0_outputs(5156)));
    outputs(1009) <= layer0_outputs(12538);
    outputs(1010) <= not(layer0_outputs(3396));
    outputs(1011) <= layer0_outputs(4189);
    outputs(1012) <= not(layer0_outputs(249)) or (layer0_outputs(5583));
    outputs(1013) <= (layer0_outputs(83)) xor (layer0_outputs(4562));
    outputs(1014) <= layer0_outputs(12781);
    outputs(1015) <= (layer0_outputs(11783)) or (layer0_outputs(1662));
    outputs(1016) <= layer0_outputs(12487);
    outputs(1017) <= not(layer0_outputs(2264));
    outputs(1018) <= (layer0_outputs(12013)) and (layer0_outputs(9327));
    outputs(1019) <= (layer0_outputs(841)) xor (layer0_outputs(7336));
    outputs(1020) <= not((layer0_outputs(6009)) and (layer0_outputs(4740)));
    outputs(1021) <= (layer0_outputs(10483)) xor (layer0_outputs(1827));
    outputs(1022) <= (layer0_outputs(3251)) xor (layer0_outputs(8896));
    outputs(1023) <= (layer0_outputs(1241)) xor (layer0_outputs(11726));
    outputs(1024) <= (layer0_outputs(1984)) and not (layer0_outputs(7495));
    outputs(1025) <= (layer0_outputs(10778)) xor (layer0_outputs(8396));
    outputs(1026) <= layer0_outputs(8854);
    outputs(1027) <= not((layer0_outputs(658)) xor (layer0_outputs(7237)));
    outputs(1028) <= not(layer0_outputs(4539));
    outputs(1029) <= layer0_outputs(8710);
    outputs(1030) <= (layer0_outputs(7261)) xor (layer0_outputs(5192));
    outputs(1031) <= not(layer0_outputs(455));
    outputs(1032) <= not((layer0_outputs(3799)) or (layer0_outputs(532)));
    outputs(1033) <= not(layer0_outputs(2334));
    outputs(1034) <= (layer0_outputs(12094)) and not (layer0_outputs(6684));
    outputs(1035) <= layer0_outputs(8531);
    outputs(1036) <= layer0_outputs(4473);
    outputs(1037) <= (layer0_outputs(2819)) xor (layer0_outputs(9314));
    outputs(1038) <= not((layer0_outputs(643)) and (layer0_outputs(9557)));
    outputs(1039) <= not(layer0_outputs(11473));
    outputs(1040) <= (layer0_outputs(4694)) and not (layer0_outputs(8210));
    outputs(1041) <= (layer0_outputs(5205)) xor (layer0_outputs(3186));
    outputs(1042) <= (layer0_outputs(11108)) xor (layer0_outputs(4964));
    outputs(1043) <= (layer0_outputs(4273)) and not (layer0_outputs(3854));
    outputs(1044) <= not(layer0_outputs(10347));
    outputs(1045) <= not((layer0_outputs(1081)) and (layer0_outputs(10891)));
    outputs(1046) <= not((layer0_outputs(12459)) xor (layer0_outputs(7058)));
    outputs(1047) <= (layer0_outputs(504)) and not (layer0_outputs(6599));
    outputs(1048) <= layer0_outputs(1523);
    outputs(1049) <= not((layer0_outputs(11691)) xor (layer0_outputs(6624)));
    outputs(1050) <= layer0_outputs(6182);
    outputs(1051) <= not(layer0_outputs(8964));
    outputs(1052) <= not((layer0_outputs(7486)) xor (layer0_outputs(3999)));
    outputs(1053) <= layer0_outputs(2103);
    outputs(1054) <= not(layer0_outputs(2171));
    outputs(1055) <= not((layer0_outputs(9099)) xor (layer0_outputs(4126)));
    outputs(1056) <= (layer0_outputs(8680)) and (layer0_outputs(10605));
    outputs(1057) <= not(layer0_outputs(12556));
    outputs(1058) <= not((layer0_outputs(3613)) xor (layer0_outputs(2398)));
    outputs(1059) <= not(layer0_outputs(4627));
    outputs(1060) <= (layer0_outputs(5704)) and not (layer0_outputs(2266));
    outputs(1061) <= layer0_outputs(1306);
    outputs(1062) <= (layer0_outputs(2251)) xor (layer0_outputs(9724));
    outputs(1063) <= (layer0_outputs(6622)) xor (layer0_outputs(8659));
    outputs(1064) <= not((layer0_outputs(2261)) and (layer0_outputs(11082)));
    outputs(1065) <= layer0_outputs(10604);
    outputs(1066) <= (layer0_outputs(9179)) or (layer0_outputs(5169));
    outputs(1067) <= not(layer0_outputs(749));
    outputs(1068) <= layer0_outputs(7378);
    outputs(1069) <= (layer0_outputs(6963)) xor (layer0_outputs(722));
    outputs(1070) <= not((layer0_outputs(5674)) xor (layer0_outputs(10839)));
    outputs(1071) <= not((layer0_outputs(9776)) xor (layer0_outputs(4302)));
    outputs(1072) <= (layer0_outputs(279)) and not (layer0_outputs(5950));
    outputs(1073) <= (layer0_outputs(7601)) and not (layer0_outputs(6340));
    outputs(1074) <= not((layer0_outputs(10664)) xor (layer0_outputs(2922)));
    outputs(1075) <= not(layer0_outputs(8039));
    outputs(1076) <= not(layer0_outputs(2171));
    outputs(1077) <= layer0_outputs(8842);
    outputs(1078) <= layer0_outputs(5474);
    outputs(1079) <= layer0_outputs(11679);
    outputs(1080) <= (layer0_outputs(7955)) or (layer0_outputs(8241));
    outputs(1081) <= not(layer0_outputs(7224));
    outputs(1082) <= not(layer0_outputs(10136)) or (layer0_outputs(2283));
    outputs(1083) <= (layer0_outputs(6706)) xor (layer0_outputs(3376));
    outputs(1084) <= (layer0_outputs(10577)) xor (layer0_outputs(11098));
    outputs(1085) <= not(layer0_outputs(10660));
    outputs(1086) <= not((layer0_outputs(6522)) xor (layer0_outputs(12477)));
    outputs(1087) <= layer0_outputs(1690);
    outputs(1088) <= (layer0_outputs(3432)) xor (layer0_outputs(626));
    outputs(1089) <= layer0_outputs(8195);
    outputs(1090) <= (layer0_outputs(4318)) and (layer0_outputs(5568));
    outputs(1091) <= layer0_outputs(1222);
    outputs(1092) <= not((layer0_outputs(7425)) and (layer0_outputs(3415)));
    outputs(1093) <= (layer0_outputs(12749)) and not (layer0_outputs(4446));
    outputs(1094) <= layer0_outputs(10167);
    outputs(1095) <= not((layer0_outputs(7729)) xor (layer0_outputs(3921)));
    outputs(1096) <= not((layer0_outputs(1800)) xor (layer0_outputs(1288)));
    outputs(1097) <= (layer0_outputs(6222)) and (layer0_outputs(2767));
    outputs(1098) <= not(layer0_outputs(8563));
    outputs(1099) <= not((layer0_outputs(10901)) and (layer0_outputs(5457)));
    outputs(1100) <= not((layer0_outputs(8480)) or (layer0_outputs(7302)));
    outputs(1101) <= not((layer0_outputs(644)) xor (layer0_outputs(6714)));
    outputs(1102) <= (layer0_outputs(5237)) xor (layer0_outputs(11938));
    outputs(1103) <= (layer0_outputs(8369)) xor (layer0_outputs(10035));
    outputs(1104) <= (layer0_outputs(12422)) or (layer0_outputs(10640));
    outputs(1105) <= not((layer0_outputs(5802)) or (layer0_outputs(7672)));
    outputs(1106) <= layer0_outputs(5083);
    outputs(1107) <= layer0_outputs(6022);
    outputs(1108) <= not(layer0_outputs(5561)) or (layer0_outputs(11323));
    outputs(1109) <= not(layer0_outputs(2393)) or (layer0_outputs(1234));
    outputs(1110) <= layer0_outputs(12013);
    outputs(1111) <= (layer0_outputs(4806)) xor (layer0_outputs(9652));
    outputs(1112) <= not(layer0_outputs(8440));
    outputs(1113) <= not((layer0_outputs(8187)) xor (layer0_outputs(6378)));
    outputs(1114) <= not(layer0_outputs(2927));
    outputs(1115) <= (layer0_outputs(6348)) xor (layer0_outputs(3222));
    outputs(1116) <= not(layer0_outputs(4525));
    outputs(1117) <= (layer0_outputs(9548)) xor (layer0_outputs(9394));
    outputs(1118) <= layer0_outputs(2273);
    outputs(1119) <= (layer0_outputs(9577)) xor (layer0_outputs(1675));
    outputs(1120) <= not(layer0_outputs(5960));
    outputs(1121) <= (layer0_outputs(518)) xor (layer0_outputs(8161));
    outputs(1122) <= not(layer0_outputs(12158));
    outputs(1123) <= layer0_outputs(3976);
    outputs(1124) <= layer0_outputs(12075);
    outputs(1125) <= not(layer0_outputs(4551));
    outputs(1126) <= not(layer0_outputs(6112));
    outputs(1127) <= not(layer0_outputs(2961));
    outputs(1128) <= not((layer0_outputs(5625)) xor (layer0_outputs(7132)));
    outputs(1129) <= not(layer0_outputs(10810));
    outputs(1130) <= not(layer0_outputs(4478));
    outputs(1131) <= layer0_outputs(1683);
    outputs(1132) <= layer0_outputs(9071);
    outputs(1133) <= layer0_outputs(4117);
    outputs(1134) <= layer0_outputs(4173);
    outputs(1135) <= not(layer0_outputs(12038));
    outputs(1136) <= not(layer0_outputs(6133));
    outputs(1137) <= not(layer0_outputs(3440)) or (layer0_outputs(2032));
    outputs(1138) <= not((layer0_outputs(4388)) or (layer0_outputs(9118)));
    outputs(1139) <= not(layer0_outputs(4048));
    outputs(1140) <= (layer0_outputs(362)) xor (layer0_outputs(12708));
    outputs(1141) <= layer0_outputs(2572);
    outputs(1142) <= not(layer0_outputs(75));
    outputs(1143) <= not(layer0_outputs(11288));
    outputs(1144) <= not(layer0_outputs(12712));
    outputs(1145) <= not(layer0_outputs(7122));
    outputs(1146) <= layer0_outputs(12428);
    outputs(1147) <= not(layer0_outputs(9303));
    outputs(1148) <= (layer0_outputs(8323)) xor (layer0_outputs(9990));
    outputs(1149) <= not((layer0_outputs(10797)) xor (layer0_outputs(5760)));
    outputs(1150) <= (layer0_outputs(8945)) and not (layer0_outputs(10511));
    outputs(1151) <= not(layer0_outputs(3137));
    outputs(1152) <= (layer0_outputs(333)) xor (layer0_outputs(9558));
    outputs(1153) <= (layer0_outputs(9135)) and not (layer0_outputs(3309));
    outputs(1154) <= not(layer0_outputs(8651));
    outputs(1155) <= layer0_outputs(6802);
    outputs(1156) <= layer0_outputs(5943);
    outputs(1157) <= layer0_outputs(3353);
    outputs(1158) <= (layer0_outputs(6058)) and (layer0_outputs(9605));
    outputs(1159) <= not(layer0_outputs(10373));
    outputs(1160) <= layer0_outputs(1722);
    outputs(1161) <= not(layer0_outputs(9014));
    outputs(1162) <= not(layer0_outputs(11373));
    outputs(1163) <= layer0_outputs(8671);
    outputs(1164) <= layer0_outputs(11764);
    outputs(1165) <= (layer0_outputs(4067)) xor (layer0_outputs(10532));
    outputs(1166) <= not(layer0_outputs(10033));
    outputs(1167) <= layer0_outputs(7609);
    outputs(1168) <= (layer0_outputs(1956)) xor (layer0_outputs(4545));
    outputs(1169) <= (layer0_outputs(8300)) xor (layer0_outputs(3169));
    outputs(1170) <= layer0_outputs(62);
    outputs(1171) <= not(layer0_outputs(11683)) or (layer0_outputs(1733));
    outputs(1172) <= (layer0_outputs(4096)) or (layer0_outputs(5906));
    outputs(1173) <= not((layer0_outputs(5916)) xor (layer0_outputs(5470)));
    outputs(1174) <= not((layer0_outputs(2382)) xor (layer0_outputs(9486)));
    outputs(1175) <= layer0_outputs(12151);
    outputs(1176) <= layer0_outputs(8775);
    outputs(1177) <= not(layer0_outputs(11112));
    outputs(1178) <= not(layer0_outputs(118));
    outputs(1179) <= not(layer0_outputs(6097));
    outputs(1180) <= not(layer0_outputs(462));
    outputs(1181) <= layer0_outputs(2689);
    outputs(1182) <= (layer0_outputs(6168)) and not (layer0_outputs(6861));
    outputs(1183) <= not(layer0_outputs(8316)) or (layer0_outputs(4781));
    outputs(1184) <= layer0_outputs(9239);
    outputs(1185) <= not(layer0_outputs(7974)) or (layer0_outputs(12552));
    outputs(1186) <= layer0_outputs(10416);
    outputs(1187) <= layer0_outputs(3539);
    outputs(1188) <= not(layer0_outputs(868));
    outputs(1189) <= not(layer0_outputs(5314));
    outputs(1190) <= (layer0_outputs(9770)) xor (layer0_outputs(10310));
    outputs(1191) <= (layer0_outputs(4972)) and not (layer0_outputs(3507));
    outputs(1192) <= (layer0_outputs(6054)) xor (layer0_outputs(5528));
    outputs(1193) <= not(layer0_outputs(3312));
    outputs(1194) <= not(layer0_outputs(3696));
    outputs(1195) <= layer0_outputs(6918);
    outputs(1196) <= not((layer0_outputs(10393)) xor (layer0_outputs(11268)));
    outputs(1197) <= not((layer0_outputs(9540)) or (layer0_outputs(12095)));
    outputs(1198) <= not((layer0_outputs(8840)) xor (layer0_outputs(8192)));
    outputs(1199) <= not(layer0_outputs(10034)) or (layer0_outputs(11150));
    outputs(1200) <= (layer0_outputs(5942)) or (layer0_outputs(4126));
    outputs(1201) <= not((layer0_outputs(5003)) xor (layer0_outputs(5498)));
    outputs(1202) <= layer0_outputs(181);
    outputs(1203) <= not(layer0_outputs(687)) or (layer0_outputs(9974));
    outputs(1204) <= (layer0_outputs(10844)) xor (layer0_outputs(617));
    outputs(1205) <= not((layer0_outputs(10258)) xor (layer0_outputs(4593)));
    outputs(1206) <= not(layer0_outputs(3178));
    outputs(1207) <= not((layer0_outputs(5754)) xor (layer0_outputs(7481)));
    outputs(1208) <= not(layer0_outputs(2007));
    outputs(1209) <= not(layer0_outputs(4858)) or (layer0_outputs(4984));
    outputs(1210) <= not(layer0_outputs(12395));
    outputs(1211) <= (layer0_outputs(6479)) and (layer0_outputs(1708));
    outputs(1212) <= layer0_outputs(6791);
    outputs(1213) <= layer0_outputs(3683);
    outputs(1214) <= not(layer0_outputs(3102)) or (layer0_outputs(8420));
    outputs(1215) <= not(layer0_outputs(996));
    outputs(1216) <= (layer0_outputs(2408)) xor (layer0_outputs(4495));
    outputs(1217) <= (layer0_outputs(7158)) xor (layer0_outputs(11297));
    outputs(1218) <= (layer0_outputs(1510)) and not (layer0_outputs(42));
    outputs(1219) <= (layer0_outputs(6111)) and not (layer0_outputs(6122));
    outputs(1220) <= layer0_outputs(7221);
    outputs(1221) <= layer0_outputs(10192);
    outputs(1222) <= not(layer0_outputs(7349));
    outputs(1223) <= layer0_outputs(9482);
    outputs(1224) <= not(layer0_outputs(11685));
    outputs(1225) <= (layer0_outputs(957)) xor (layer0_outputs(8858));
    outputs(1226) <= (layer0_outputs(7244)) or (layer0_outputs(10255));
    outputs(1227) <= layer0_outputs(1577);
    outputs(1228) <= layer0_outputs(2628);
    outputs(1229) <= not((layer0_outputs(12156)) xor (layer0_outputs(9060)));
    outputs(1230) <= layer0_outputs(8608);
    outputs(1231) <= not(layer0_outputs(7143));
    outputs(1232) <= (layer0_outputs(10799)) xor (layer0_outputs(8560));
    outputs(1233) <= (layer0_outputs(11325)) xor (layer0_outputs(11575));
    outputs(1234) <= not(layer0_outputs(7356));
    outputs(1235) <= (layer0_outputs(4644)) and (layer0_outputs(7316));
    outputs(1236) <= (layer0_outputs(1979)) xor (layer0_outputs(10597));
    outputs(1237) <= layer0_outputs(128);
    outputs(1238) <= not(layer0_outputs(9191)) or (layer0_outputs(2673));
    outputs(1239) <= not(layer0_outputs(11904));
    outputs(1240) <= (layer0_outputs(8896)) xor (layer0_outputs(4606));
    outputs(1241) <= (layer0_outputs(4576)) and not (layer0_outputs(10030));
    outputs(1242) <= not((layer0_outputs(9054)) xor (layer0_outputs(10396)));
    outputs(1243) <= not(layer0_outputs(5389)) or (layer0_outputs(3743));
    outputs(1244) <= not((layer0_outputs(2207)) or (layer0_outputs(6923)));
    outputs(1245) <= not(layer0_outputs(11713));
    outputs(1246) <= (layer0_outputs(1246)) xor (layer0_outputs(11739));
    outputs(1247) <= layer0_outputs(8470);
    outputs(1248) <= (layer0_outputs(12354)) and (layer0_outputs(2015));
    outputs(1249) <= (layer0_outputs(2868)) and not (layer0_outputs(3851));
    outputs(1250) <= not((layer0_outputs(2677)) or (layer0_outputs(2936)));
    outputs(1251) <= layer0_outputs(431);
    outputs(1252) <= not((layer0_outputs(2567)) xor (layer0_outputs(10319)));
    outputs(1253) <= not(layer0_outputs(2021));
    outputs(1254) <= not(layer0_outputs(6188));
    outputs(1255) <= layer0_outputs(6609);
    outputs(1256) <= layer0_outputs(4895);
    outputs(1257) <= (layer0_outputs(8914)) or (layer0_outputs(7602));
    outputs(1258) <= not((layer0_outputs(2836)) xor (layer0_outputs(4021)));
    outputs(1259) <= layer0_outputs(7119);
    outputs(1260) <= not((layer0_outputs(1707)) xor (layer0_outputs(3756)));
    outputs(1261) <= not((layer0_outputs(9020)) xor (layer0_outputs(11940)));
    outputs(1262) <= not((layer0_outputs(7919)) xor (layer0_outputs(7207)));
    outputs(1263) <= not((layer0_outputs(7309)) xor (layer0_outputs(8995)));
    outputs(1264) <= (layer0_outputs(6919)) xor (layer0_outputs(8730));
    outputs(1265) <= not((layer0_outputs(8309)) xor (layer0_outputs(5886)));
    outputs(1266) <= (layer0_outputs(4334)) xor (layer0_outputs(4043));
    outputs(1267) <= not(layer0_outputs(7920));
    outputs(1268) <= layer0_outputs(4196);
    outputs(1269) <= layer0_outputs(4832);
    outputs(1270) <= layer0_outputs(12692);
    outputs(1271) <= (layer0_outputs(2023)) xor (layer0_outputs(1509));
    outputs(1272) <= not((layer0_outputs(4181)) and (layer0_outputs(12555)));
    outputs(1273) <= (layer0_outputs(560)) and not (layer0_outputs(5276));
    outputs(1274) <= not(layer0_outputs(5927));
    outputs(1275) <= not(layer0_outputs(12002));
    outputs(1276) <= not(layer0_outputs(2275));
    outputs(1277) <= not(layer0_outputs(8180)) or (layer0_outputs(5638));
    outputs(1278) <= layer0_outputs(5717);
    outputs(1279) <= (layer0_outputs(2211)) xor (layer0_outputs(9531));
    outputs(1280) <= layer0_outputs(5463);
    outputs(1281) <= not(layer0_outputs(9280));
    outputs(1282) <= not((layer0_outputs(7899)) or (layer0_outputs(10351)));
    outputs(1283) <= (layer0_outputs(10221)) and (layer0_outputs(9640));
    outputs(1284) <= layer0_outputs(9979);
    outputs(1285) <= not((layer0_outputs(7531)) or (layer0_outputs(872)));
    outputs(1286) <= layer0_outputs(1966);
    outputs(1287) <= (layer0_outputs(10943)) and not (layer0_outputs(11727));
    outputs(1288) <= not(layer0_outputs(10230));
    outputs(1289) <= (layer0_outputs(9875)) and not (layer0_outputs(7926));
    outputs(1290) <= (layer0_outputs(9066)) and (layer0_outputs(636));
    outputs(1291) <= (layer0_outputs(7009)) xor (layer0_outputs(12105));
    outputs(1292) <= (layer0_outputs(377)) and (layer0_outputs(2466));
    outputs(1293) <= (layer0_outputs(10427)) and (layer0_outputs(12030));
    outputs(1294) <= (layer0_outputs(3801)) and (layer0_outputs(8128));
    outputs(1295) <= not((layer0_outputs(11723)) or (layer0_outputs(2220)));
    outputs(1296) <= (layer0_outputs(10006)) and (layer0_outputs(12597));
    outputs(1297) <= not((layer0_outputs(9498)) xor (layer0_outputs(11992)));
    outputs(1298) <= not((layer0_outputs(8518)) xor (layer0_outputs(482)));
    outputs(1299) <= layer0_outputs(9056);
    outputs(1300) <= layer0_outputs(5289);
    outputs(1301) <= (layer0_outputs(4815)) and not (layer0_outputs(9548));
    outputs(1302) <= (layer0_outputs(6429)) and not (layer0_outputs(10534));
    outputs(1303) <= (layer0_outputs(8876)) xor (layer0_outputs(284));
    outputs(1304) <= (layer0_outputs(6077)) and not (layer0_outputs(2637));
    outputs(1305) <= (layer0_outputs(6249)) xor (layer0_outputs(7120));
    outputs(1306) <= (layer0_outputs(1266)) xor (layer0_outputs(9598));
    outputs(1307) <= not((layer0_outputs(2222)) xor (layer0_outputs(11172)));
    outputs(1308) <= layer0_outputs(11645);
    outputs(1309) <= layer0_outputs(4187);
    outputs(1310) <= not((layer0_outputs(4805)) or (layer0_outputs(333)));
    outputs(1311) <= (layer0_outputs(5922)) and not (layer0_outputs(9919));
    outputs(1312) <= (layer0_outputs(2589)) xor (layer0_outputs(10306));
    outputs(1313) <= (layer0_outputs(1937)) and not (layer0_outputs(6790));
    outputs(1314) <= (layer0_outputs(6781)) xor (layer0_outputs(7622));
    outputs(1315) <= (layer0_outputs(11831)) and (layer0_outputs(1592));
    outputs(1316) <= not(layer0_outputs(3928));
    outputs(1317) <= (layer0_outputs(12779)) and not (layer0_outputs(3301));
    outputs(1318) <= not((layer0_outputs(3290)) xor (layer0_outputs(4531)));
    outputs(1319) <= (layer0_outputs(5276)) xor (layer0_outputs(7940));
    outputs(1320) <= (layer0_outputs(1835)) and not (layer0_outputs(3751));
    outputs(1321) <= (layer0_outputs(1993)) xor (layer0_outputs(7789));
    outputs(1322) <= (layer0_outputs(3081)) xor (layer0_outputs(2265));
    outputs(1323) <= not((layer0_outputs(8610)) xor (layer0_outputs(1026)));
    outputs(1324) <= (layer0_outputs(11165)) and not (layer0_outputs(8914));
    outputs(1325) <= layer0_outputs(530);
    outputs(1326) <= not((layer0_outputs(9198)) or (layer0_outputs(6546)));
    outputs(1327) <= (layer0_outputs(1402)) xor (layer0_outputs(5392));
    outputs(1328) <= (layer0_outputs(451)) and not (layer0_outputs(8203));
    outputs(1329) <= (layer0_outputs(3634)) and (layer0_outputs(6489));
    outputs(1330) <= (layer0_outputs(9806)) and not (layer0_outputs(2738));
    outputs(1331) <= (layer0_outputs(2418)) and not (layer0_outputs(2336));
    outputs(1332) <= (layer0_outputs(7633)) xor (layer0_outputs(2319));
    outputs(1333) <= not(layer0_outputs(6360));
    outputs(1334) <= (layer0_outputs(8367)) and not (layer0_outputs(5462));
    outputs(1335) <= layer0_outputs(1655);
    outputs(1336) <= layer0_outputs(4962);
    outputs(1337) <= layer0_outputs(5987);
    outputs(1338) <= not(layer0_outputs(7258));
    outputs(1339) <= layer0_outputs(5849);
    outputs(1340) <= not((layer0_outputs(4818)) or (layer0_outputs(5575)));
    outputs(1341) <= (layer0_outputs(7966)) and (layer0_outputs(12265));
    outputs(1342) <= (layer0_outputs(11939)) and not (layer0_outputs(11583));
    outputs(1343) <= layer0_outputs(6031);
    outputs(1344) <= (layer0_outputs(7573)) and not (layer0_outputs(12204));
    outputs(1345) <= not((layer0_outputs(8473)) or (layer0_outputs(1535)));
    outputs(1346) <= (layer0_outputs(5215)) xor (layer0_outputs(4625));
    outputs(1347) <= layer0_outputs(2798);
    outputs(1348) <= not((layer0_outputs(3179)) or (layer0_outputs(7366)));
    outputs(1349) <= not(layer0_outputs(5941));
    outputs(1350) <= not((layer0_outputs(4023)) xor (layer0_outputs(11265)));
    outputs(1351) <= (layer0_outputs(3834)) and not (layer0_outputs(7799));
    outputs(1352) <= not(layer0_outputs(8001));
    outputs(1353) <= not(layer0_outputs(11038));
    outputs(1354) <= not((layer0_outputs(11705)) xor (layer0_outputs(3038)));
    outputs(1355) <= (layer0_outputs(7425)) and (layer0_outputs(183));
    outputs(1356) <= not(layer0_outputs(4513)) or (layer0_outputs(11930));
    outputs(1357) <= (layer0_outputs(6967)) xor (layer0_outputs(12560));
    outputs(1358) <= (layer0_outputs(12773)) xor (layer0_outputs(12688));
    outputs(1359) <= layer0_outputs(9352);
    outputs(1360) <= layer0_outputs(64);
    outputs(1361) <= (layer0_outputs(6084)) and (layer0_outputs(11247));
    outputs(1362) <= (layer0_outputs(8664)) xor (layer0_outputs(7596));
    outputs(1363) <= (layer0_outputs(12602)) and not (layer0_outputs(8353));
    outputs(1364) <= not((layer0_outputs(1297)) xor (layer0_outputs(11014)));
    outputs(1365) <= (layer0_outputs(3307)) and (layer0_outputs(11825));
    outputs(1366) <= (layer0_outputs(11333)) and not (layer0_outputs(9093));
    outputs(1367) <= not((layer0_outputs(9887)) xor (layer0_outputs(11599)));
    outputs(1368) <= not((layer0_outputs(590)) xor (layer0_outputs(8785)));
    outputs(1369) <= (layer0_outputs(10401)) xor (layer0_outputs(7672));
    outputs(1370) <= (layer0_outputs(7548)) and (layer0_outputs(10101));
    outputs(1371) <= not(layer0_outputs(7332));
    outputs(1372) <= (layer0_outputs(7901)) and not (layer0_outputs(6611));
    outputs(1373) <= (layer0_outputs(9621)) and not (layer0_outputs(8888));
    outputs(1374) <= (layer0_outputs(6311)) and not (layer0_outputs(3584));
    outputs(1375) <= (layer0_outputs(4671)) xor (layer0_outputs(2519));
    outputs(1376) <= layer0_outputs(4302);
    outputs(1377) <= layer0_outputs(4472);
    outputs(1378) <= (layer0_outputs(10322)) xor (layer0_outputs(6716));
    outputs(1379) <= not(layer0_outputs(9311));
    outputs(1380) <= not(layer0_outputs(2742));
    outputs(1381) <= (layer0_outputs(12108)) xor (layer0_outputs(1249));
    outputs(1382) <= (layer0_outputs(2409)) and not (layer0_outputs(3292));
    outputs(1383) <= (layer0_outputs(4558)) xor (layer0_outputs(10637));
    outputs(1384) <= layer0_outputs(1700);
    outputs(1385) <= not((layer0_outputs(11153)) xor (layer0_outputs(10740)));
    outputs(1386) <= layer0_outputs(847);
    outputs(1387) <= not((layer0_outputs(5360)) xor (layer0_outputs(9938)));
    outputs(1388) <= (layer0_outputs(7612)) and not (layer0_outputs(5165));
    outputs(1389) <= layer0_outputs(9574);
    outputs(1390) <= not((layer0_outputs(3591)) xor (layer0_outputs(2240)));
    outputs(1391) <= not((layer0_outputs(6943)) xor (layer0_outputs(7039)));
    outputs(1392) <= (layer0_outputs(11648)) xor (layer0_outputs(8196));
    outputs(1393) <= layer0_outputs(8883);
    outputs(1394) <= (layer0_outputs(392)) xor (layer0_outputs(11833));
    outputs(1395) <= (layer0_outputs(7388)) and (layer0_outputs(9713));
    outputs(1396) <= (layer0_outputs(1035)) and not (layer0_outputs(5883));
    outputs(1397) <= not(layer0_outputs(2525));
    outputs(1398) <= (layer0_outputs(7154)) xor (layer0_outputs(4483));
    outputs(1399) <= (layer0_outputs(198)) and not (layer0_outputs(877));
    outputs(1400) <= not(layer0_outputs(10811));
    outputs(1401) <= (layer0_outputs(2324)) and not (layer0_outputs(9459));
    outputs(1402) <= not((layer0_outputs(1974)) xor (layer0_outputs(9420)));
    outputs(1403) <= not(layer0_outputs(8035));
    outputs(1404) <= (layer0_outputs(11425)) xor (layer0_outputs(2387));
    outputs(1405) <= not((layer0_outputs(194)) xor (layer0_outputs(8652)));
    outputs(1406) <= (layer0_outputs(2202)) xor (layer0_outputs(6530));
    outputs(1407) <= (layer0_outputs(3096)) xor (layer0_outputs(12008));
    outputs(1408) <= (layer0_outputs(11823)) xor (layer0_outputs(7896));
    outputs(1409) <= not((layer0_outputs(8131)) or (layer0_outputs(11132)));
    outputs(1410) <= layer0_outputs(883);
    outputs(1411) <= (layer0_outputs(12042)) xor (layer0_outputs(7954));
    outputs(1412) <= not(layer0_outputs(7724));
    outputs(1413) <= not(layer0_outputs(568));
    outputs(1414) <= not(layer0_outputs(45));
    outputs(1415) <= (layer0_outputs(1780)) xor (layer0_outputs(11910));
    outputs(1416) <= (layer0_outputs(5545)) xor (layer0_outputs(9665));
    outputs(1417) <= not(layer0_outputs(9313));
    outputs(1418) <= (layer0_outputs(734)) and not (layer0_outputs(11477));
    outputs(1419) <= (layer0_outputs(1519)) xor (layer0_outputs(1350));
    outputs(1420) <= (layer0_outputs(5619)) and not (layer0_outputs(9601));
    outputs(1421) <= (layer0_outputs(9497)) and (layer0_outputs(11306));
    outputs(1422) <= layer0_outputs(6142);
    outputs(1423) <= not((layer0_outputs(12444)) xor (layer0_outputs(2392)));
    outputs(1424) <= (layer0_outputs(9413)) xor (layer0_outputs(7073));
    outputs(1425) <= (layer0_outputs(11842)) xor (layer0_outputs(11804));
    outputs(1426) <= (layer0_outputs(7345)) xor (layer0_outputs(5473));
    outputs(1427) <= (layer0_outputs(1077)) xor (layer0_outputs(8675));
    outputs(1428) <= (layer0_outputs(12122)) and not (layer0_outputs(1087));
    outputs(1429) <= not(layer0_outputs(5114));
    outputs(1430) <= not((layer0_outputs(2259)) xor (layer0_outputs(88)));
    outputs(1431) <= (layer0_outputs(2407)) and not (layer0_outputs(6966));
    outputs(1432) <= not(layer0_outputs(11470));
    outputs(1433) <= layer0_outputs(5554);
    outputs(1434) <= (layer0_outputs(12294)) xor (layer0_outputs(9082));
    outputs(1435) <= (layer0_outputs(11372)) and not (layer0_outputs(9949));
    outputs(1436) <= (layer0_outputs(10308)) xor (layer0_outputs(10567));
    outputs(1437) <= not((layer0_outputs(7611)) xor (layer0_outputs(6163)));
    outputs(1438) <= not((layer0_outputs(3127)) xor (layer0_outputs(9283)));
    outputs(1439) <= not((layer0_outputs(7492)) xor (layer0_outputs(9888)));
    outputs(1440) <= (layer0_outputs(8650)) and (layer0_outputs(2980));
    outputs(1441) <= (layer0_outputs(11823)) xor (layer0_outputs(7175));
    outputs(1442) <= layer0_outputs(942);
    outputs(1443) <= not((layer0_outputs(11761)) or (layer0_outputs(11311)));
    outputs(1444) <= not((layer0_outputs(7153)) or (layer0_outputs(8163)));
    outputs(1445) <= (layer0_outputs(3654)) xor (layer0_outputs(10893));
    outputs(1446) <= (layer0_outputs(3406)) and not (layer0_outputs(12209));
    outputs(1447) <= (layer0_outputs(7614)) xor (layer0_outputs(192));
    outputs(1448) <= not((layer0_outputs(2133)) xor (layer0_outputs(10119)));
    outputs(1449) <= not(layer0_outputs(9));
    outputs(1450) <= (layer0_outputs(12302)) and not (layer0_outputs(3471));
    outputs(1451) <= not((layer0_outputs(6913)) or (layer0_outputs(12296)));
    outputs(1452) <= (layer0_outputs(6318)) and not (layer0_outputs(9049));
    outputs(1453) <= not((layer0_outputs(12634)) xor (layer0_outputs(1546)));
    outputs(1454) <= (layer0_outputs(10234)) and not (layer0_outputs(12348));
    outputs(1455) <= (layer0_outputs(5961)) and not (layer0_outputs(12348));
    outputs(1456) <= (layer0_outputs(6883)) xor (layer0_outputs(4885));
    outputs(1457) <= not(layer0_outputs(9491));
    outputs(1458) <= '0';
    outputs(1459) <= layer0_outputs(10458);
    outputs(1460) <= '0';
    outputs(1461) <= (layer0_outputs(10279)) and not (layer0_outputs(4915));
    outputs(1462) <= (layer0_outputs(6049)) xor (layer0_outputs(7849));
    outputs(1463) <= (layer0_outputs(11193)) xor (layer0_outputs(9631));
    outputs(1464) <= (layer0_outputs(2686)) and not (layer0_outputs(2764));
    outputs(1465) <= layer0_outputs(5383);
    outputs(1466) <= not((layer0_outputs(1786)) or (layer0_outputs(2188)));
    outputs(1467) <= (layer0_outputs(5852)) and (layer0_outputs(2604));
    outputs(1468) <= (layer0_outputs(3520)) and not (layer0_outputs(2539));
    outputs(1469) <= (layer0_outputs(8944)) and (layer0_outputs(2363));
    outputs(1470) <= (layer0_outputs(1411)) and not (layer0_outputs(10313));
    outputs(1471) <= (layer0_outputs(9897)) and not (layer0_outputs(3097));
    outputs(1472) <= (layer0_outputs(7414)) and (layer0_outputs(10440));
    outputs(1473) <= (layer0_outputs(12284)) and not (layer0_outputs(1646));
    outputs(1474) <= (layer0_outputs(6356)) and not (layer0_outputs(2050));
    outputs(1475) <= not((layer0_outputs(2682)) or (layer0_outputs(11668)));
    outputs(1476) <= (layer0_outputs(9205)) and not (layer0_outputs(3938));
    outputs(1477) <= not((layer0_outputs(450)) or (layer0_outputs(4814)));
    outputs(1478) <= not((layer0_outputs(4991)) or (layer0_outputs(12075)));
    outputs(1479) <= not((layer0_outputs(10301)) or (layer0_outputs(11478)));
    outputs(1480) <= (layer0_outputs(5097)) and not (layer0_outputs(6111));
    outputs(1481) <= (layer0_outputs(8831)) xor (layer0_outputs(6682));
    outputs(1482) <= (layer0_outputs(1716)) and (layer0_outputs(12103));
    outputs(1483) <= layer0_outputs(5697);
    outputs(1484) <= layer0_outputs(11464);
    outputs(1485) <= layer0_outputs(11364);
    outputs(1486) <= (layer0_outputs(2406)) and not (layer0_outputs(1279));
    outputs(1487) <= layer0_outputs(2318);
    outputs(1488) <= layer0_outputs(4580);
    outputs(1489) <= (layer0_outputs(11997)) xor (layer0_outputs(7822));
    outputs(1490) <= not(layer0_outputs(7171));
    outputs(1491) <= (layer0_outputs(8432)) and not (layer0_outputs(11548));
    outputs(1492) <= not(layer0_outputs(1195));
    outputs(1493) <= layer0_outputs(10989);
    outputs(1494) <= (layer0_outputs(7032)) xor (layer0_outputs(11095));
    outputs(1495) <= not(layer0_outputs(2755));
    outputs(1496) <= (layer0_outputs(8402)) xor (layer0_outputs(4454));
    outputs(1497) <= (layer0_outputs(9945)) and (layer0_outputs(5030));
    outputs(1498) <= not(layer0_outputs(2305));
    outputs(1499) <= not((layer0_outputs(7871)) xor (layer0_outputs(6467)));
    outputs(1500) <= not((layer0_outputs(8417)) xor (layer0_outputs(11363)));
    outputs(1501) <= not((layer0_outputs(4047)) or (layer0_outputs(11168)));
    outputs(1502) <= (layer0_outputs(9808)) and (layer0_outputs(5659));
    outputs(1503) <= (layer0_outputs(10279)) and (layer0_outputs(9932));
    outputs(1504) <= (layer0_outputs(7585)) and not (layer0_outputs(10551));
    outputs(1505) <= (layer0_outputs(4691)) and (layer0_outputs(8862));
    outputs(1506) <= not(layer0_outputs(10538));
    outputs(1507) <= (layer0_outputs(823)) and (layer0_outputs(11633));
    outputs(1508) <= layer0_outputs(11578);
    outputs(1509) <= (layer0_outputs(5901)) xor (layer0_outputs(7915));
    outputs(1510) <= not((layer0_outputs(4288)) xor (layer0_outputs(12059)));
    outputs(1511) <= layer0_outputs(8376);
    outputs(1512) <= not(layer0_outputs(10788));
    outputs(1513) <= (layer0_outputs(4903)) and not (layer0_outputs(1288));
    outputs(1514) <= not(layer0_outputs(2338));
    outputs(1515) <= not(layer0_outputs(7591));
    outputs(1516) <= not(layer0_outputs(10339));
    outputs(1517) <= (layer0_outputs(318)) and not (layer0_outputs(3531));
    outputs(1518) <= not(layer0_outputs(2201));
    outputs(1519) <= layer0_outputs(1875);
    outputs(1520) <= (layer0_outputs(4310)) xor (layer0_outputs(11519));
    outputs(1521) <= (layer0_outputs(2701)) and (layer0_outputs(3284));
    outputs(1522) <= (layer0_outputs(6817)) xor (layer0_outputs(10989));
    outputs(1523) <= not((layer0_outputs(10244)) or (layer0_outputs(8698)));
    outputs(1524) <= not((layer0_outputs(9128)) or (layer0_outputs(3660)));
    outputs(1525) <= (layer0_outputs(2349)) and (layer0_outputs(4400));
    outputs(1526) <= (layer0_outputs(71)) xor (layer0_outputs(10523));
    outputs(1527) <= not(layer0_outputs(7753));
    outputs(1528) <= (layer0_outputs(381)) and (layer0_outputs(289));
    outputs(1529) <= (layer0_outputs(1244)) and not (layer0_outputs(8612));
    outputs(1530) <= not(layer0_outputs(2443));
    outputs(1531) <= (layer0_outputs(11471)) and not (layer0_outputs(11352));
    outputs(1532) <= (layer0_outputs(11002)) and not (layer0_outputs(2465));
    outputs(1533) <= not((layer0_outputs(2709)) xor (layer0_outputs(407)));
    outputs(1534) <= not(layer0_outputs(478));
    outputs(1535) <= not((layer0_outputs(4846)) xor (layer0_outputs(8797)));
    outputs(1536) <= layer0_outputs(11138);
    outputs(1537) <= layer0_outputs(3501);
    outputs(1538) <= (layer0_outputs(2154)) and not (layer0_outputs(10194));
    outputs(1539) <= not(layer0_outputs(7895));
    outputs(1540) <= (layer0_outputs(1632)) and (layer0_outputs(4894));
    outputs(1541) <= not((layer0_outputs(5609)) or (layer0_outputs(5481)));
    outputs(1542) <= not((layer0_outputs(389)) xor (layer0_outputs(2124)));
    outputs(1543) <= not(layer0_outputs(8638));
    outputs(1544) <= (layer0_outputs(7471)) and (layer0_outputs(12390));
    outputs(1545) <= (layer0_outputs(12623)) and not (layer0_outputs(4838));
    outputs(1546) <= not((layer0_outputs(11339)) xor (layer0_outputs(4183)));
    outputs(1547) <= layer0_outputs(6671);
    outputs(1548) <= not(layer0_outputs(9462));
    outputs(1549) <= not((layer0_outputs(1102)) xor (layer0_outputs(9775)));
    outputs(1550) <= layer0_outputs(3445);
    outputs(1551) <= (layer0_outputs(3514)) and not (layer0_outputs(3085));
    outputs(1552) <= not((layer0_outputs(2402)) or (layer0_outputs(2335)));
    outputs(1553) <= not((layer0_outputs(864)) xor (layer0_outputs(2204)));
    outputs(1554) <= not((layer0_outputs(6067)) or (layer0_outputs(2471)));
    outputs(1555) <= not((layer0_outputs(10540)) xor (layer0_outputs(1458)));
    outputs(1556) <= layer0_outputs(11686);
    outputs(1557) <= not(layer0_outputs(10184));
    outputs(1558) <= (layer0_outputs(12551)) and not (layer0_outputs(6220));
    outputs(1559) <= layer0_outputs(6042);
    outputs(1560) <= (layer0_outputs(12760)) and not (layer0_outputs(10986));
    outputs(1561) <= not(layer0_outputs(8292));
    outputs(1562) <= (layer0_outputs(8633)) and (layer0_outputs(10141));
    outputs(1563) <= (layer0_outputs(4737)) xor (layer0_outputs(2799));
    outputs(1564) <= (layer0_outputs(10405)) and not (layer0_outputs(8801));
    outputs(1565) <= not(layer0_outputs(10058));
    outputs(1566) <= not((layer0_outputs(514)) or (layer0_outputs(6913)));
    outputs(1567) <= not((layer0_outputs(7817)) xor (layer0_outputs(12124)));
    outputs(1568) <= not(layer0_outputs(1242));
    outputs(1569) <= (layer0_outputs(8359)) and not (layer0_outputs(8099));
    outputs(1570) <= (layer0_outputs(11243)) and not (layer0_outputs(2084));
    outputs(1571) <= not(layer0_outputs(4515));
    outputs(1572) <= layer0_outputs(8439);
    outputs(1573) <= not(layer0_outputs(5390));
    outputs(1574) <= (layer0_outputs(7394)) and not (layer0_outputs(5235));
    outputs(1575) <= (layer0_outputs(163)) and (layer0_outputs(6897));
    outputs(1576) <= (layer0_outputs(1593)) and not (layer0_outputs(7462));
    outputs(1577) <= not(layer0_outputs(4999));
    outputs(1578) <= layer0_outputs(6073);
    outputs(1579) <= (layer0_outputs(10372)) xor (layer0_outputs(2941));
    outputs(1580) <= not((layer0_outputs(4898)) or (layer0_outputs(5690)));
    outputs(1581) <= not((layer0_outputs(2987)) xor (layer0_outputs(3165)));
    outputs(1582) <= not(layer0_outputs(11696)) or (layer0_outputs(4412));
    outputs(1583) <= not((layer0_outputs(10884)) or (layer0_outputs(10687)));
    outputs(1584) <= not((layer0_outputs(11967)) xor (layer0_outputs(8046)));
    outputs(1585) <= not((layer0_outputs(6502)) and (layer0_outputs(399)));
    outputs(1586) <= not((layer0_outputs(1854)) or (layer0_outputs(7902)));
    outputs(1587) <= (layer0_outputs(9398)) and (layer0_outputs(11733));
    outputs(1588) <= (layer0_outputs(11537)) and (layer0_outputs(10402));
    outputs(1589) <= (layer0_outputs(6551)) xor (layer0_outputs(4174));
    outputs(1590) <= (layer0_outputs(12314)) and (layer0_outputs(8505));
    outputs(1591) <= (layer0_outputs(11810)) and (layer0_outputs(10539));
    outputs(1592) <= (layer0_outputs(6760)) xor (layer0_outputs(7534));
    outputs(1593) <= not((layer0_outputs(4877)) or (layer0_outputs(11968)));
    outputs(1594) <= not((layer0_outputs(1635)) or (layer0_outputs(9755)));
    outputs(1595) <= not((layer0_outputs(623)) xor (layer0_outputs(9617)));
    outputs(1596) <= (layer0_outputs(5248)) xor (layer0_outputs(2480));
    outputs(1597) <= (layer0_outputs(8804)) and not (layer0_outputs(7935));
    outputs(1598) <= (layer0_outputs(12558)) xor (layer0_outputs(11624));
    outputs(1599) <= (layer0_outputs(2538)) and not (layer0_outputs(12386));
    outputs(1600) <= (layer0_outputs(122)) and not (layer0_outputs(6090));
    outputs(1601) <= (layer0_outputs(5465)) and (layer0_outputs(3692));
    outputs(1602) <= '0';
    outputs(1603) <= not((layer0_outputs(3495)) xor (layer0_outputs(6242)));
    outputs(1604) <= layer0_outputs(1002);
    outputs(1605) <= (layer0_outputs(1368)) and (layer0_outputs(11229));
    outputs(1606) <= (layer0_outputs(4904)) and not (layer0_outputs(1650));
    outputs(1607) <= (layer0_outputs(11263)) and (layer0_outputs(4849));
    outputs(1608) <= layer0_outputs(5050);
    outputs(1609) <= (layer0_outputs(10105)) xor (layer0_outputs(6023));
    outputs(1610) <= not(layer0_outputs(3992));
    outputs(1611) <= (layer0_outputs(10986)) xor (layer0_outputs(7939));
    outputs(1612) <= not((layer0_outputs(155)) xor (layer0_outputs(4859)));
    outputs(1613) <= not((layer0_outputs(4656)) xor (layer0_outputs(10169)));
    outputs(1614) <= not((layer0_outputs(9247)) xor (layer0_outputs(6252)));
    outputs(1615) <= not((layer0_outputs(8970)) xor (layer0_outputs(6098)));
    outputs(1616) <= not(layer0_outputs(9369));
    outputs(1617) <= not((layer0_outputs(11213)) xor (layer0_outputs(3851)));
    outputs(1618) <= (layer0_outputs(9130)) and not (layer0_outputs(472));
    outputs(1619) <= not((layer0_outputs(679)) xor (layer0_outputs(6317)));
    outputs(1620) <= (layer0_outputs(5831)) and (layer0_outputs(12619));
    outputs(1621) <= layer0_outputs(2399);
    outputs(1622) <= '0';
    outputs(1623) <= (layer0_outputs(5494)) and not (layer0_outputs(6053));
    outputs(1624) <= layer0_outputs(1602);
    outputs(1625) <= (layer0_outputs(4998)) and (layer0_outputs(8495));
    outputs(1626) <= (layer0_outputs(420)) xor (layer0_outputs(5273));
    outputs(1627) <= not(layer0_outputs(6547));
    outputs(1628) <= (layer0_outputs(8325)) and not (layer0_outputs(4831));
    outputs(1629) <= (layer0_outputs(125)) and not (layer0_outputs(3129));
    outputs(1630) <= (layer0_outputs(54)) and not (layer0_outputs(8532));
    outputs(1631) <= (layer0_outputs(8660)) and not (layer0_outputs(9311));
    outputs(1632) <= not((layer0_outputs(2648)) xor (layer0_outputs(8847)));
    outputs(1633) <= not(layer0_outputs(2731));
    outputs(1634) <= (layer0_outputs(5412)) and (layer0_outputs(9338));
    outputs(1635) <= (layer0_outputs(4800)) and (layer0_outputs(6011));
    outputs(1636) <= (layer0_outputs(1941)) and not (layer0_outputs(12215));
    outputs(1637) <= (layer0_outputs(5799)) and not (layer0_outputs(1459));
    outputs(1638) <= '0';
    outputs(1639) <= not((layer0_outputs(5692)) or (layer0_outputs(4269)));
    outputs(1640) <= not((layer0_outputs(11746)) xor (layer0_outputs(12758)));
    outputs(1641) <= not((layer0_outputs(6790)) or (layer0_outputs(6513)));
    outputs(1642) <= (layer0_outputs(11884)) and not (layer0_outputs(5450));
    outputs(1643) <= (layer0_outputs(9472)) and (layer0_outputs(7045));
    outputs(1644) <= (layer0_outputs(3350)) xor (layer0_outputs(3645));
    outputs(1645) <= (layer0_outputs(11206)) and not (layer0_outputs(4189));
    outputs(1646) <= layer0_outputs(3257);
    outputs(1647) <= layer0_outputs(1430);
    outputs(1648) <= (layer0_outputs(8174)) and (layer0_outputs(3383));
    outputs(1649) <= not((layer0_outputs(2987)) xor (layer0_outputs(8092)));
    outputs(1650) <= (layer0_outputs(1115)) xor (layer0_outputs(5188));
    outputs(1651) <= layer0_outputs(7099);
    outputs(1652) <= (layer0_outputs(3028)) and not (layer0_outputs(5440));
    outputs(1653) <= (layer0_outputs(9667)) xor (layer0_outputs(12574));
    outputs(1654) <= not((layer0_outputs(1311)) xor (layer0_outputs(9584)));
    outputs(1655) <= (layer0_outputs(11260)) xor (layer0_outputs(5100));
    outputs(1656) <= not((layer0_outputs(3639)) xor (layer0_outputs(11424)));
    outputs(1657) <= (layer0_outputs(1611)) and not (layer0_outputs(4821));
    outputs(1658) <= not(layer0_outputs(473));
    outputs(1659) <= layer0_outputs(2935);
    outputs(1660) <= (layer0_outputs(2919)) and (layer0_outputs(5201));
    outputs(1661) <= (layer0_outputs(5543)) and not (layer0_outputs(6134));
    outputs(1662) <= (layer0_outputs(3174)) and not (layer0_outputs(6540));
    outputs(1663) <= layer0_outputs(5178);
    outputs(1664) <= not((layer0_outputs(12649)) or (layer0_outputs(6256)));
    outputs(1665) <= not((layer0_outputs(5371)) xor (layer0_outputs(7327)));
    outputs(1666) <= (layer0_outputs(9793)) xor (layer0_outputs(3534));
    outputs(1667) <= (layer0_outputs(12727)) and not (layer0_outputs(1715));
    outputs(1668) <= (layer0_outputs(11181)) xor (layer0_outputs(7897));
    outputs(1669) <= (layer0_outputs(11543)) and not (layer0_outputs(5563));
    outputs(1670) <= not(layer0_outputs(5585));
    outputs(1671) <= (layer0_outputs(3951)) and not (layer0_outputs(10530));
    outputs(1672) <= not(layer0_outputs(4124));
    outputs(1673) <= (layer0_outputs(11462)) and not (layer0_outputs(3859));
    outputs(1674) <= (layer0_outputs(6614)) and not (layer0_outputs(7266));
    outputs(1675) <= not((layer0_outputs(5310)) xor (layer0_outputs(10399)));
    outputs(1676) <= not(layer0_outputs(10538));
    outputs(1677) <= (layer0_outputs(10641)) xor (layer0_outputs(6752));
    outputs(1678) <= not((layer0_outputs(4705)) xor (layer0_outputs(2603)));
    outputs(1679) <= not((layer0_outputs(2735)) xor (layer0_outputs(4025)));
    outputs(1680) <= layer0_outputs(3155);
    outputs(1681) <= (layer0_outputs(10227)) xor (layer0_outputs(7564));
    outputs(1682) <= not((layer0_outputs(2215)) xor (layer0_outputs(12090)));
    outputs(1683) <= (layer0_outputs(6114)) and not (layer0_outputs(8120));
    outputs(1684) <= not(layer0_outputs(1142));
    outputs(1685) <= (layer0_outputs(6455)) and not (layer0_outputs(12323));
    outputs(1686) <= (layer0_outputs(9020)) and (layer0_outputs(29));
    outputs(1687) <= (layer0_outputs(462)) xor (layer0_outputs(1624));
    outputs(1688) <= (layer0_outputs(10525)) and (layer0_outputs(10217));
    outputs(1689) <= (layer0_outputs(10112)) and not (layer0_outputs(4024));
    outputs(1690) <= (layer0_outputs(7440)) xor (layer0_outputs(12042));
    outputs(1691) <= (layer0_outputs(8187)) xor (layer0_outputs(1070));
    outputs(1692) <= (layer0_outputs(12510)) and (layer0_outputs(4646));
    outputs(1693) <= (layer0_outputs(4896)) and not (layer0_outputs(3593));
    outputs(1694) <= (layer0_outputs(4162)) and (layer0_outputs(12293));
    outputs(1695) <= not(layer0_outputs(2827));
    outputs(1696) <= not((layer0_outputs(12416)) xor (layer0_outputs(1041)));
    outputs(1697) <= not(layer0_outputs(4979)) or (layer0_outputs(9620));
    outputs(1698) <= (layer0_outputs(9537)) xor (layer0_outputs(7140));
    outputs(1699) <= not((layer0_outputs(6309)) xor (layer0_outputs(8159)));
    outputs(1700) <= not((layer0_outputs(2773)) xor (layer0_outputs(9609)));
    outputs(1701) <= layer0_outputs(1768);
    outputs(1702) <= (layer0_outputs(6816)) xor (layer0_outputs(9863));
    outputs(1703) <= layer0_outputs(4075);
    outputs(1704) <= layer0_outputs(5320);
    outputs(1705) <= not(layer0_outputs(6971));
    outputs(1706) <= (layer0_outputs(5369)) and (layer0_outputs(5554));
    outputs(1707) <= not((layer0_outputs(8269)) xor (layer0_outputs(11360)));
    outputs(1708) <= (layer0_outputs(2405)) and not (layer0_outputs(7671));
    outputs(1709) <= (layer0_outputs(270)) and not (layer0_outputs(7341));
    outputs(1710) <= not((layer0_outputs(6362)) xor (layer0_outputs(6126)));
    outputs(1711) <= not((layer0_outputs(6592)) xor (layer0_outputs(1709)));
    outputs(1712) <= (layer0_outputs(658)) and not (layer0_outputs(5028));
    outputs(1713) <= (layer0_outputs(8113)) and not (layer0_outputs(10863));
    outputs(1714) <= not((layer0_outputs(10828)) or (layer0_outputs(12527)));
    outputs(1715) <= not((layer0_outputs(6730)) or (layer0_outputs(7940)));
    outputs(1716) <= not(layer0_outputs(2089));
    outputs(1717) <= (layer0_outputs(8728)) and (layer0_outputs(2449));
    outputs(1718) <= not(layer0_outputs(12328));
    outputs(1719) <= not((layer0_outputs(12730)) xor (layer0_outputs(10875)));
    outputs(1720) <= (layer0_outputs(8229)) xor (layer0_outputs(10555));
    outputs(1721) <= (layer0_outputs(12220)) and (layer0_outputs(7944));
    outputs(1722) <= not(layer0_outputs(9735));
    outputs(1723) <= '0';
    outputs(1724) <= not(layer0_outputs(10895));
    outputs(1725) <= not((layer0_outputs(8513)) xor (layer0_outputs(3945)));
    outputs(1726) <= not((layer0_outputs(3926)) xor (layer0_outputs(10222)));
    outputs(1727) <= not((layer0_outputs(4086)) or (layer0_outputs(1560)));
    outputs(1728) <= (layer0_outputs(10191)) and (layer0_outputs(10321));
    outputs(1729) <= (layer0_outputs(3056)) xor (layer0_outputs(11352));
    outputs(1730) <= not(layer0_outputs(7130));
    outputs(1731) <= not((layer0_outputs(12270)) xor (layer0_outputs(10213)));
    outputs(1732) <= not(layer0_outputs(4303));
    outputs(1733) <= (layer0_outputs(6438)) and not (layer0_outputs(3795));
    outputs(1734) <= (layer0_outputs(10532)) and not (layer0_outputs(9031));
    outputs(1735) <= (layer0_outputs(9204)) and not (layer0_outputs(8490));
    outputs(1736) <= (layer0_outputs(10501)) and not (layer0_outputs(6275));
    outputs(1737) <= (layer0_outputs(4619)) xor (layer0_outputs(9308));
    outputs(1738) <= (layer0_outputs(1420)) xor (layer0_outputs(2470));
    outputs(1739) <= not((layer0_outputs(3238)) or (layer0_outputs(2237)));
    outputs(1740) <= not(layer0_outputs(2133));
    outputs(1741) <= (layer0_outputs(10137)) and not (layer0_outputs(365));
    outputs(1742) <= not((layer0_outputs(3761)) or (layer0_outputs(11052)));
    outputs(1743) <= not((layer0_outputs(5754)) xor (layer0_outputs(5491)));
    outputs(1744) <= not(layer0_outputs(12446));
    outputs(1745) <= (layer0_outputs(2784)) xor (layer0_outputs(8146));
    outputs(1746) <= (layer0_outputs(6007)) xor (layer0_outputs(8492));
    outputs(1747) <= not(layer0_outputs(5877));
    outputs(1748) <= not(layer0_outputs(12685));
    outputs(1749) <= (layer0_outputs(2544)) xor (layer0_outputs(5483));
    outputs(1750) <= not(layer0_outputs(10550));
    outputs(1751) <= not((layer0_outputs(4668)) xor (layer0_outputs(12055)));
    outputs(1752) <= (layer0_outputs(10102)) and not (layer0_outputs(3138));
    outputs(1753) <= (layer0_outputs(11646)) and (layer0_outputs(6553));
    outputs(1754) <= (layer0_outputs(6028)) and not (layer0_outputs(8399));
    outputs(1755) <= (layer0_outputs(10537)) and not (layer0_outputs(2799));
    outputs(1756) <= not((layer0_outputs(4680)) xor (layer0_outputs(2761)));
    outputs(1757) <= not((layer0_outputs(807)) or (layer0_outputs(7619)));
    outputs(1758) <= (layer0_outputs(500)) xor (layer0_outputs(3863));
    outputs(1759) <= layer0_outputs(2502);
    outputs(1760) <= (layer0_outputs(3466)) and (layer0_outputs(11144));
    outputs(1761) <= (layer0_outputs(4144)) and not (layer0_outputs(1633));
    outputs(1762) <= not(layer0_outputs(10591));
    outputs(1763) <= (layer0_outputs(3888)) and not (layer0_outputs(2270));
    outputs(1764) <= (layer0_outputs(9260)) and not (layer0_outputs(11702));
    outputs(1765) <= not(layer0_outputs(9679));
    outputs(1766) <= not((layer0_outputs(10683)) or (layer0_outputs(3918)));
    outputs(1767) <= (layer0_outputs(694)) and (layer0_outputs(2238));
    outputs(1768) <= (layer0_outputs(9556)) and not (layer0_outputs(6385));
    outputs(1769) <= not(layer0_outputs(1310));
    outputs(1770) <= not((layer0_outputs(6952)) or (layer0_outputs(12188)));
    outputs(1771) <= layer0_outputs(2588);
    outputs(1772) <= not(layer0_outputs(1501)) or (layer0_outputs(2408));
    outputs(1773) <= not((layer0_outputs(3326)) or (layer0_outputs(3588)));
    outputs(1774) <= not((layer0_outputs(7797)) or (layer0_outputs(3640)));
    outputs(1775) <= not((layer0_outputs(9790)) xor (layer0_outputs(165)));
    outputs(1776) <= layer0_outputs(6336);
    outputs(1777) <= not((layer0_outputs(9411)) or (layer0_outputs(6378)));
    outputs(1778) <= not(layer0_outputs(10353));
    outputs(1779) <= not((layer0_outputs(356)) xor (layer0_outputs(3152)));
    outputs(1780) <= (layer0_outputs(11831)) and not (layer0_outputs(5186));
    outputs(1781) <= (layer0_outputs(3099)) xor (layer0_outputs(4920));
    outputs(1782) <= (layer0_outputs(2147)) xor (layer0_outputs(11072));
    outputs(1783) <= (layer0_outputs(9169)) and (layer0_outputs(10588));
    outputs(1784) <= (layer0_outputs(2138)) and not (layer0_outputs(1181));
    outputs(1785) <= layer0_outputs(2152);
    outputs(1786) <= (layer0_outputs(4812)) and not (layer0_outputs(11369));
    outputs(1787) <= (layer0_outputs(11664)) and not (layer0_outputs(9147));
    outputs(1788) <= (layer0_outputs(9371)) and not (layer0_outputs(2781));
    outputs(1789) <= not((layer0_outputs(10677)) xor (layer0_outputs(307)));
    outputs(1790) <= (layer0_outputs(2038)) xor (layer0_outputs(924));
    outputs(1791) <= (layer0_outputs(1360)) and (layer0_outputs(7961));
    outputs(1792) <= layer0_outputs(8224);
    outputs(1793) <= layer0_outputs(6785);
    outputs(1794) <= layer0_outputs(9331);
    outputs(1795) <= not((layer0_outputs(1948)) or (layer0_outputs(9079)));
    outputs(1796) <= layer0_outputs(9569);
    outputs(1797) <= not(layer0_outputs(7420));
    outputs(1798) <= (layer0_outputs(9504)) xor (layer0_outputs(6370));
    outputs(1799) <= not((layer0_outputs(4150)) xor (layer0_outputs(2847)));
    outputs(1800) <= (layer0_outputs(10104)) and not (layer0_outputs(6953));
    outputs(1801) <= (layer0_outputs(6793)) and not (layer0_outputs(8887));
    outputs(1802) <= not((layer0_outputs(7325)) xor (layer0_outputs(5084)));
    outputs(1803) <= (layer0_outputs(11645)) and (layer0_outputs(7109));
    outputs(1804) <= not((layer0_outputs(10081)) xor (layer0_outputs(7669)));
    outputs(1805) <= not((layer0_outputs(6046)) xor (layer0_outputs(1242)));
    outputs(1806) <= not((layer0_outputs(9587)) xor (layer0_outputs(11523)));
    outputs(1807) <= (layer0_outputs(7848)) xor (layer0_outputs(5454));
    outputs(1808) <= not((layer0_outputs(8057)) xor (layer0_outputs(5850)));
    outputs(1809) <= not(layer0_outputs(4876));
    outputs(1810) <= (layer0_outputs(3354)) and not (layer0_outputs(6134));
    outputs(1811) <= (layer0_outputs(693)) and not (layer0_outputs(6427));
    outputs(1812) <= (layer0_outputs(5979)) and not (layer0_outputs(7070));
    outputs(1813) <= '0';
    outputs(1814) <= not((layer0_outputs(7514)) xor (layer0_outputs(4514)));
    outputs(1815) <= not(layer0_outputs(8160));
    outputs(1816) <= not(layer0_outputs(5621));
    outputs(1817) <= (layer0_outputs(4958)) and not (layer0_outputs(2028));
    outputs(1818) <= (layer0_outputs(3602)) xor (layer0_outputs(12344));
    outputs(1819) <= (layer0_outputs(7369)) xor (layer0_outputs(8301));
    outputs(1820) <= (layer0_outputs(6006)) and (layer0_outputs(1826));
    outputs(1821) <= not((layer0_outputs(4360)) xor (layer0_outputs(755)));
    outputs(1822) <= not(layer0_outputs(8419));
    outputs(1823) <= (layer0_outputs(11060)) xor (layer0_outputs(12741));
    outputs(1824) <= not((layer0_outputs(12731)) or (layer0_outputs(2749)));
    outputs(1825) <= not(layer0_outputs(5574));
    outputs(1826) <= (layer0_outputs(5355)) and not (layer0_outputs(6436));
    outputs(1827) <= not((layer0_outputs(1061)) xor (layer0_outputs(5042)));
    outputs(1828) <= layer0_outputs(10237);
    outputs(1829) <= (layer0_outputs(7026)) and not (layer0_outputs(12523));
    outputs(1830) <= '0';
    outputs(1831) <= not((layer0_outputs(10065)) or (layer0_outputs(4319)));
    outputs(1832) <= (layer0_outputs(2005)) xor (layer0_outputs(2839));
    outputs(1833) <= not((layer0_outputs(2801)) or (layer0_outputs(12713)));
    outputs(1834) <= (layer0_outputs(2820)) and not (layer0_outputs(2065));
    outputs(1835) <= (layer0_outputs(3615)) and not (layer0_outputs(472));
    outputs(1836) <= not((layer0_outputs(7209)) or (layer0_outputs(9285)));
    outputs(1837) <= (layer0_outputs(892)) xor (layer0_outputs(3675));
    outputs(1838) <= (layer0_outputs(11508)) xor (layer0_outputs(2665));
    outputs(1839) <= layer0_outputs(1039);
    outputs(1840) <= (layer0_outputs(10905)) xor (layer0_outputs(350));
    outputs(1841) <= not((layer0_outputs(7728)) or (layer0_outputs(9646)));
    outputs(1842) <= layer0_outputs(11995);
    outputs(1843) <= not(layer0_outputs(8023));
    outputs(1844) <= (layer0_outputs(6202)) and not (layer0_outputs(4820));
    outputs(1845) <= not((layer0_outputs(2942)) or (layer0_outputs(10301)));
    outputs(1846) <= (layer0_outputs(538)) xor (layer0_outputs(9372));
    outputs(1847) <= not((layer0_outputs(450)) or (layer0_outputs(8173)));
    outputs(1848) <= (layer0_outputs(7986)) xor (layer0_outputs(3778));
    outputs(1849) <= (layer0_outputs(2979)) and (layer0_outputs(10763));
    outputs(1850) <= layer0_outputs(6746);
    outputs(1851) <= (layer0_outputs(7553)) xor (layer0_outputs(336));
    outputs(1852) <= (layer0_outputs(9461)) xor (layer0_outputs(2916));
    outputs(1853) <= (layer0_outputs(1161)) and (layer0_outputs(1105));
    outputs(1854) <= (layer0_outputs(6085)) and not (layer0_outputs(11784));
    outputs(1855) <= (layer0_outputs(103)) and (layer0_outputs(11793));
    outputs(1856) <= not(layer0_outputs(9651));
    outputs(1857) <= not(layer0_outputs(150));
    outputs(1858) <= not((layer0_outputs(8308)) or (layer0_outputs(6819)));
    outputs(1859) <= '0';
    outputs(1860) <= (layer0_outputs(9430)) and not (layer0_outputs(12678));
    outputs(1861) <= layer0_outputs(6416);
    outputs(1862) <= '0';
    outputs(1863) <= not((layer0_outputs(3752)) or (layer0_outputs(67)));
    outputs(1864) <= layer0_outputs(4912);
    outputs(1865) <= not(layer0_outputs(8409));
    outputs(1866) <= not((layer0_outputs(2972)) xor (layer0_outputs(6588)));
    outputs(1867) <= not(layer0_outputs(4103));
    outputs(1868) <= (layer0_outputs(7006)) and not (layer0_outputs(4145));
    outputs(1869) <= not(layer0_outputs(10429));
    outputs(1870) <= (layer0_outputs(10960)) xor (layer0_outputs(9374));
    outputs(1871) <= layer0_outputs(2483);
    outputs(1872) <= not(layer0_outputs(9795));
    outputs(1873) <= layer0_outputs(6692);
    outputs(1874) <= not((layer0_outputs(7120)) xor (layer0_outputs(10418)));
    outputs(1875) <= (layer0_outputs(7958)) and not (layer0_outputs(3590));
    outputs(1876) <= (layer0_outputs(946)) xor (layer0_outputs(3235));
    outputs(1877) <= not((layer0_outputs(12363)) xor (layer0_outputs(3768)));
    outputs(1878) <= (layer0_outputs(6992)) xor (layer0_outputs(5101));
    outputs(1879) <= layer0_outputs(7314);
    outputs(1880) <= (layer0_outputs(2362)) and (layer0_outputs(7071));
    outputs(1881) <= (layer0_outputs(5468)) xor (layer0_outputs(5668));
    outputs(1882) <= (layer0_outputs(12234)) and not (layer0_outputs(9287));
    outputs(1883) <= (layer0_outputs(4082)) and not (layer0_outputs(351));
    outputs(1884) <= not((layer0_outputs(9106)) xor (layer0_outputs(1359)));
    outputs(1885) <= (layer0_outputs(5388)) and (layer0_outputs(1677));
    outputs(1886) <= (layer0_outputs(1863)) and (layer0_outputs(2719));
    outputs(1887) <= not((layer0_outputs(5350)) xor (layer0_outputs(11054)));
    outputs(1888) <= (layer0_outputs(7453)) and not (layer0_outputs(7836));
    outputs(1889) <= (layer0_outputs(247)) xor (layer0_outputs(664));
    outputs(1890) <= (layer0_outputs(9164)) xor (layer0_outputs(402));
    outputs(1891) <= not(layer0_outputs(6945));
    outputs(1892) <= (layer0_outputs(7274)) xor (layer0_outputs(10819));
    outputs(1893) <= not((layer0_outputs(137)) xor (layer0_outputs(3788)));
    outputs(1894) <= (layer0_outputs(10569)) and not (layer0_outputs(11714));
    outputs(1895) <= layer0_outputs(11799);
    outputs(1896) <= not(layer0_outputs(9457));
    outputs(1897) <= (layer0_outputs(12098)) xor (layer0_outputs(11608));
    outputs(1898) <= (layer0_outputs(8296)) and (layer0_outputs(317));
    outputs(1899) <= (layer0_outputs(1889)) and not (layer0_outputs(10049));
    outputs(1900) <= not((layer0_outputs(1094)) xor (layer0_outputs(1642)));
    outputs(1901) <= (layer0_outputs(2348)) xor (layer0_outputs(834));
    outputs(1902) <= not(layer0_outputs(1298));
    outputs(1903) <= (layer0_outputs(4852)) and (layer0_outputs(1227));
    outputs(1904) <= not((layer0_outputs(6342)) or (layer0_outputs(10061)));
    outputs(1905) <= (layer0_outputs(8645)) and not (layer0_outputs(5969));
    outputs(1906) <= (layer0_outputs(4275)) and not (layer0_outputs(4327));
    outputs(1907) <= (layer0_outputs(1713)) xor (layer0_outputs(10939));
    outputs(1908) <= layer0_outputs(11683);
    outputs(1909) <= (layer0_outputs(6988)) and not (layer0_outputs(5879));
    outputs(1910) <= (layer0_outputs(8711)) and not (layer0_outputs(6198));
    outputs(1911) <= not(layer0_outputs(10364));
    outputs(1912) <= '0';
    outputs(1913) <= (layer0_outputs(11056)) and not (layer0_outputs(6381));
    outputs(1914) <= (layer0_outputs(12505)) and (layer0_outputs(6100));
    outputs(1915) <= (layer0_outputs(6191)) xor (layer0_outputs(6689));
    outputs(1916) <= (layer0_outputs(10838)) and not (layer0_outputs(6866));
    outputs(1917) <= layer0_outputs(6329);
    outputs(1918) <= (layer0_outputs(12695)) and (layer0_outputs(10547));
    outputs(1919) <= (layer0_outputs(1485)) xor (layer0_outputs(10791));
    outputs(1920) <= not((layer0_outputs(116)) or (layer0_outputs(11978)));
    outputs(1921) <= layer0_outputs(9162);
    outputs(1922) <= not((layer0_outputs(8602)) or (layer0_outputs(11819)));
    outputs(1923) <= (layer0_outputs(5928)) and not (layer0_outputs(4838));
    outputs(1924) <= layer0_outputs(4665);
    outputs(1925) <= not((layer0_outputs(2613)) xor (layer0_outputs(5279)));
    outputs(1926) <= layer0_outputs(11155);
    outputs(1927) <= layer0_outputs(2564);
    outputs(1928) <= (layer0_outputs(3574)) xor (layer0_outputs(9861));
    outputs(1929) <= (layer0_outputs(5810)) and not (layer0_outputs(12613));
    outputs(1930) <= (layer0_outputs(7019)) and not (layer0_outputs(9267));
    outputs(1931) <= (layer0_outputs(9164)) xor (layer0_outputs(4134));
    outputs(1932) <= not(layer0_outputs(10921)) or (layer0_outputs(9620));
    outputs(1933) <= not((layer0_outputs(3541)) xor (layer0_outputs(6193)));
    outputs(1934) <= (layer0_outputs(2727)) and not (layer0_outputs(268));
    outputs(1935) <= (layer0_outputs(11390)) and (layer0_outputs(12502));
    outputs(1936) <= not((layer0_outputs(2788)) xor (layer0_outputs(8575)));
    outputs(1937) <= not((layer0_outputs(937)) xor (layer0_outputs(3157)));
    outputs(1938) <= not((layer0_outputs(3214)) or (layer0_outputs(11005)));
    outputs(1939) <= (layer0_outputs(3263)) and not (layer0_outputs(1735));
    outputs(1940) <= not((layer0_outputs(7496)) xor (layer0_outputs(2674)));
    outputs(1941) <= not((layer0_outputs(11173)) xor (layer0_outputs(2474)));
    outputs(1942) <= not((layer0_outputs(7814)) or (layer0_outputs(6776)));
    outputs(1943) <= (layer0_outputs(8647)) and (layer0_outputs(3689));
    outputs(1944) <= not(layer0_outputs(6424));
    outputs(1945) <= (layer0_outputs(5978)) xor (layer0_outputs(11536));
    outputs(1946) <= not(layer0_outputs(9160));
    outputs(1947) <= layer0_outputs(9497);
    outputs(1948) <= not((layer0_outputs(11142)) or (layer0_outputs(2693)));
    outputs(1949) <= (layer0_outputs(11264)) and not (layer0_outputs(9886));
    outputs(1950) <= layer0_outputs(11030);
    outputs(1951) <= (layer0_outputs(12381)) xor (layer0_outputs(5265));
    outputs(1952) <= (layer0_outputs(2873)) and not (layer0_outputs(2145));
    outputs(1953) <= (layer0_outputs(785)) xor (layer0_outputs(9287));
    outputs(1954) <= not((layer0_outputs(2774)) xor (layer0_outputs(7641)));
    outputs(1955) <= (layer0_outputs(1650)) xor (layer0_outputs(11558));
    outputs(1956) <= not(layer0_outputs(11923));
    outputs(1957) <= (layer0_outputs(227)) and not (layer0_outputs(7616));
    outputs(1958) <= (layer0_outputs(10602)) and not (layer0_outputs(11983));
    outputs(1959) <= not((layer0_outputs(2828)) xor (layer0_outputs(1786)));
    outputs(1960) <= not(layer0_outputs(9608));
    outputs(1961) <= (layer0_outputs(12412)) and not (layer0_outputs(3108));
    outputs(1962) <= (layer0_outputs(2164)) and (layer0_outputs(2974));
    outputs(1963) <= (layer0_outputs(2562)) and not (layer0_outputs(11855));
    outputs(1964) <= (layer0_outputs(9005)) and (layer0_outputs(8660));
    outputs(1965) <= not(layer0_outputs(2747));
    outputs(1966) <= (layer0_outputs(2372)) and not (layer0_outputs(10764));
    outputs(1967) <= layer0_outputs(7496);
    outputs(1968) <= not((layer0_outputs(8348)) xor (layer0_outputs(7449)));
    outputs(1969) <= '0';
    outputs(1970) <= (layer0_outputs(12262)) and not (layer0_outputs(12758));
    outputs(1971) <= not(layer0_outputs(4379));
    outputs(1972) <= (layer0_outputs(12623)) and not (layer0_outputs(6859));
    outputs(1973) <= '0';
    outputs(1974) <= not((layer0_outputs(3091)) xor (layer0_outputs(1514)));
    outputs(1975) <= not((layer0_outputs(2432)) xor (layer0_outputs(3814)));
    outputs(1976) <= not((layer0_outputs(7679)) xor (layer0_outputs(10636)));
    outputs(1977) <= not((layer0_outputs(11714)) or (layer0_outputs(6541)));
    outputs(1978) <= (layer0_outputs(4003)) and (layer0_outputs(412));
    outputs(1979) <= not(layer0_outputs(12146)) or (layer0_outputs(12404));
    outputs(1980) <= (layer0_outputs(8841)) and not (layer0_outputs(8831));
    outputs(1981) <= not((layer0_outputs(8230)) and (layer0_outputs(9876)));
    outputs(1982) <= layer0_outputs(5632);
    outputs(1983) <= not(layer0_outputs(1657));
    outputs(1984) <= not((layer0_outputs(10929)) or (layer0_outputs(708)));
    outputs(1985) <= not(layer0_outputs(3941));
    outputs(1986) <= not((layer0_outputs(1103)) xor (layer0_outputs(12098)));
    outputs(1987) <= not((layer0_outputs(12773)) xor (layer0_outputs(10613)));
    outputs(1988) <= not(layer0_outputs(9866));
    outputs(1989) <= layer0_outputs(6560);
    outputs(1990) <= (layer0_outputs(7128)) and not (layer0_outputs(1668));
    outputs(1991) <= not((layer0_outputs(5499)) xor (layer0_outputs(8076)));
    outputs(1992) <= not((layer0_outputs(5583)) xor (layer0_outputs(7136)));
    outputs(1993) <= (layer0_outputs(4394)) and not (layer0_outputs(5168));
    outputs(1994) <= layer0_outputs(787);
    outputs(1995) <= (layer0_outputs(4366)) xor (layer0_outputs(4857));
    outputs(1996) <= not((layer0_outputs(5387)) xor (layer0_outputs(6995)));
    outputs(1997) <= not((layer0_outputs(1498)) xor (layer0_outputs(10916)));
    outputs(1998) <= not((layer0_outputs(7479)) xor (layer0_outputs(8745)));
    outputs(1999) <= not((layer0_outputs(6934)) xor (layer0_outputs(7625)));
    outputs(2000) <= (layer0_outputs(10695)) xor (layer0_outputs(6212));
    outputs(2001) <= (layer0_outputs(8838)) and (layer0_outputs(4617));
    outputs(2002) <= not((layer0_outputs(4091)) xor (layer0_outputs(3574)));
    outputs(2003) <= layer0_outputs(10171);
    outputs(2004) <= (layer0_outputs(9402)) xor (layer0_outputs(447));
    outputs(2005) <= (layer0_outputs(3930)) and (layer0_outputs(11597));
    outputs(2006) <= not(layer0_outputs(990));
    outputs(2007) <= not(layer0_outputs(10747));
    outputs(2008) <= not((layer0_outputs(2649)) or (layer0_outputs(1638)));
    outputs(2009) <= not((layer0_outputs(6005)) or (layer0_outputs(2397)));
    outputs(2010) <= (layer0_outputs(10093)) xor (layer0_outputs(1143));
    outputs(2011) <= (layer0_outputs(8645)) and not (layer0_outputs(3800));
    outputs(2012) <= (layer0_outputs(10935)) and (layer0_outputs(7010));
    outputs(2013) <= not(layer0_outputs(4971));
    outputs(2014) <= (layer0_outputs(4689)) xor (layer0_outputs(10308));
    outputs(2015) <= layer0_outputs(3915);
    outputs(2016) <= (layer0_outputs(3162)) and not (layer0_outputs(8074));
    outputs(2017) <= (layer0_outputs(370)) and not (layer0_outputs(3690));
    outputs(2018) <= (layer0_outputs(10078)) and not (layer0_outputs(11908));
    outputs(2019) <= (layer0_outputs(4746)) or (layer0_outputs(1004));
    outputs(2020) <= (layer0_outputs(9665)) and not (layer0_outputs(8963));
    outputs(2021) <= (layer0_outputs(8450)) and not (layer0_outputs(5067));
    outputs(2022) <= layer0_outputs(5463);
    outputs(2023) <= (layer0_outputs(7933)) xor (layer0_outputs(5173));
    outputs(2024) <= (layer0_outputs(4639)) and (layer0_outputs(4626));
    outputs(2025) <= not((layer0_outputs(1748)) xor (layer0_outputs(11021)));
    outputs(2026) <= not((layer0_outputs(5396)) or (layer0_outputs(870)));
    outputs(2027) <= not((layer0_outputs(109)) or (layer0_outputs(11684)));
    outputs(2028) <= not(layer0_outputs(9092));
    outputs(2029) <= not(layer0_outputs(7141));
    outputs(2030) <= (layer0_outputs(6956)) and not (layer0_outputs(12596));
    outputs(2031) <= (layer0_outputs(10457)) and not (layer0_outputs(6263));
    outputs(2032) <= (layer0_outputs(6233)) and (layer0_outputs(7275));
    outputs(2033) <= not((layer0_outputs(10751)) or (layer0_outputs(12589)));
    outputs(2034) <= not(layer0_outputs(209));
    outputs(2035) <= not((layer0_outputs(9815)) xor (layer0_outputs(7656)));
    outputs(2036) <= not((layer0_outputs(1381)) or (layer0_outputs(9561)));
    outputs(2037) <= (layer0_outputs(8098)) and not (layer0_outputs(5930));
    outputs(2038) <= (layer0_outputs(4031)) and (layer0_outputs(2157));
    outputs(2039) <= not((layer0_outputs(6239)) xor (layer0_outputs(11342)));
    outputs(2040) <= (layer0_outputs(5961)) xor (layer0_outputs(3272));
    outputs(2041) <= not(layer0_outputs(7859));
    outputs(2042) <= (layer0_outputs(6511)) xor (layer0_outputs(7690));
    outputs(2043) <= '0';
    outputs(2044) <= layer0_outputs(7863);
    outputs(2045) <= (layer0_outputs(4320)) and (layer0_outputs(6826));
    outputs(2046) <= not((layer0_outputs(2214)) xor (layer0_outputs(6593)));
    outputs(2047) <= (layer0_outputs(8097)) and not (layer0_outputs(11811));
    outputs(2048) <= not(layer0_outputs(6096));
    outputs(2049) <= not(layer0_outputs(4594)) or (layer0_outputs(7737));
    outputs(2050) <= not((layer0_outputs(8182)) xor (layer0_outputs(6245)));
    outputs(2051) <= (layer0_outputs(5452)) and (layer0_outputs(2033));
    outputs(2052) <= (layer0_outputs(10727)) and not (layer0_outputs(2702));
    outputs(2053) <= (layer0_outputs(1444)) and (layer0_outputs(12047));
    outputs(2054) <= (layer0_outputs(8249)) and not (layer0_outputs(310));
    outputs(2055) <= (layer0_outputs(10481)) xor (layer0_outputs(2212));
    outputs(2056) <= (layer0_outputs(781)) and (layer0_outputs(12576));
    outputs(2057) <= (layer0_outputs(12490)) and (layer0_outputs(12416));
    outputs(2058) <= not(layer0_outputs(4823));
    outputs(2059) <= layer0_outputs(8737);
    outputs(2060) <= (layer0_outputs(1253)) and (layer0_outputs(10114));
    outputs(2061) <= layer0_outputs(8747);
    outputs(2062) <= (layer0_outputs(11148)) xor (layer0_outputs(7609));
    outputs(2063) <= layer0_outputs(11146);
    outputs(2064) <= not(layer0_outputs(7273));
    outputs(2065) <= not(layer0_outputs(2845));
    outputs(2066) <= not((layer0_outputs(314)) xor (layer0_outputs(6825)));
    outputs(2067) <= not((layer0_outputs(11397)) or (layer0_outputs(7549)));
    outputs(2068) <= (layer0_outputs(4206)) and not (layer0_outputs(1913));
    outputs(2069) <= (layer0_outputs(8673)) and (layer0_outputs(529));
    outputs(2070) <= layer0_outputs(1304);
    outputs(2071) <= not(layer0_outputs(7445));
    outputs(2072) <= (layer0_outputs(6586)) and not (layer0_outputs(2585));
    outputs(2073) <= not(layer0_outputs(1775));
    outputs(2074) <= not((layer0_outputs(1977)) or (layer0_outputs(11795)));
    outputs(2075) <= (layer0_outputs(12044)) xor (layer0_outputs(2958));
    outputs(2076) <= not((layer0_outputs(8988)) xor (layer0_outputs(9182)));
    outputs(2077) <= not((layer0_outputs(8421)) or (layer0_outputs(2684)));
    outputs(2078) <= not((layer0_outputs(8428)) xor (layer0_outputs(8265)));
    outputs(2079) <= (layer0_outputs(2151)) xor (layer0_outputs(4611));
    outputs(2080) <= not(layer0_outputs(873));
    outputs(2081) <= not((layer0_outputs(8452)) or (layer0_outputs(12725)));
    outputs(2082) <= not(layer0_outputs(2034));
    outputs(2083) <= (layer0_outputs(5)) and (layer0_outputs(9344));
    outputs(2084) <= layer0_outputs(3549);
    outputs(2085) <= (layer0_outputs(3117)) and not (layer0_outputs(10358));
    outputs(2086) <= layer0_outputs(3306);
    outputs(2087) <= layer0_outputs(9923);
    outputs(2088) <= (layer0_outputs(613)) and not (layer0_outputs(9677));
    outputs(2089) <= (layer0_outputs(3260)) and not (layer0_outputs(11809));
    outputs(2090) <= (layer0_outputs(2671)) xor (layer0_outputs(4786));
    outputs(2091) <= (layer0_outputs(5785)) and not (layer0_outputs(1096));
    outputs(2092) <= not((layer0_outputs(11449)) xor (layer0_outputs(254)));
    outputs(2093) <= layer0_outputs(4129);
    outputs(2094) <= not((layer0_outputs(2180)) or (layer0_outputs(8271)));
    outputs(2095) <= (layer0_outputs(6712)) xor (layer0_outputs(10070));
    outputs(2096) <= (layer0_outputs(9415)) xor (layer0_outputs(5128));
    outputs(2097) <= not((layer0_outputs(137)) or (layer0_outputs(7293)));
    outputs(2098) <= not(layer0_outputs(9159));
    outputs(2099) <= (layer0_outputs(10739)) xor (layer0_outputs(1281));
    outputs(2100) <= (layer0_outputs(4638)) xor (layer0_outputs(7693));
    outputs(2101) <= (layer0_outputs(10886)) and (layer0_outputs(4763));
    outputs(2102) <= (layer0_outputs(9377)) xor (layer0_outputs(8592));
    outputs(2103) <= (layer0_outputs(5512)) and not (layer0_outputs(821));
    outputs(2104) <= not((layer0_outputs(8964)) xor (layer0_outputs(5236)));
    outputs(2105) <= not((layer0_outputs(2573)) xor (layer0_outputs(4696)));
    outputs(2106) <= not((layer0_outputs(5602)) xor (layer0_outputs(2522)));
    outputs(2107) <= (layer0_outputs(8535)) and not (layer0_outputs(1494));
    outputs(2108) <= not(layer0_outputs(11605));
    outputs(2109) <= layer0_outputs(5253);
    outputs(2110) <= not(layer0_outputs(8334));
    outputs(2111) <= (layer0_outputs(7911)) and (layer0_outputs(8959));
    outputs(2112) <= not(layer0_outputs(4231)) or (layer0_outputs(1859));
    outputs(2113) <= (layer0_outputs(3874)) and (layer0_outputs(11514));
    outputs(2114) <= not((layer0_outputs(7076)) xor (layer0_outputs(2064)));
    outputs(2115) <= not((layer0_outputs(10467)) xor (layer0_outputs(4710)));
    outputs(2116) <= not((layer0_outputs(3337)) or (layer0_outputs(10858)));
    outputs(2117) <= layer0_outputs(3142);
    outputs(2118) <= not((layer0_outputs(2479)) xor (layer0_outputs(11367)));
    outputs(2119) <= (layer0_outputs(458)) xor (layer0_outputs(5700));
    outputs(2120) <= (layer0_outputs(10957)) xor (layer0_outputs(4859));
    outputs(2121) <= not((layer0_outputs(9137)) xor (layer0_outputs(6742)));
    outputs(2122) <= not((layer0_outputs(10031)) xor (layer0_outputs(5023)));
    outputs(2123) <= not((layer0_outputs(1466)) or (layer0_outputs(1172)));
    outputs(2124) <= (layer0_outputs(6323)) xor (layer0_outputs(1542));
    outputs(2125) <= (layer0_outputs(3860)) and not (layer0_outputs(4874));
    outputs(2126) <= (layer0_outputs(3482)) and not (layer0_outputs(2678));
    outputs(2127) <= not((layer0_outputs(9962)) xor (layer0_outputs(2169)));
    outputs(2128) <= not(layer0_outputs(4274)) or (layer0_outputs(1707));
    outputs(2129) <= (layer0_outputs(12407)) xor (layer0_outputs(5775));
    outputs(2130) <= not((layer0_outputs(11092)) xor (layer0_outputs(12393)));
    outputs(2131) <= (layer0_outputs(3529)) and not (layer0_outputs(10095));
    outputs(2132) <= '0';
    outputs(2133) <= (layer0_outputs(12683)) and (layer0_outputs(8375));
    outputs(2134) <= (layer0_outputs(9782)) and not (layer0_outputs(11415));
    outputs(2135) <= not((layer0_outputs(240)) xor (layer0_outputs(10587)));
    outputs(2136) <= not(layer0_outputs(8760));
    outputs(2137) <= (layer0_outputs(876)) and (layer0_outputs(4595));
    outputs(2138) <= (layer0_outputs(2368)) and not (layer0_outputs(671));
    outputs(2139) <= not((layer0_outputs(2640)) xor (layer0_outputs(1942)));
    outputs(2140) <= (layer0_outputs(687)) xor (layer0_outputs(12026));
    outputs(2141) <= not(layer0_outputs(5540));
    outputs(2142) <= (layer0_outputs(5442)) and (layer0_outputs(3207));
    outputs(2143) <= (layer0_outputs(1141)) xor (layer0_outputs(5006));
    outputs(2144) <= not((layer0_outputs(12777)) xor (layer0_outputs(9999)));
    outputs(2145) <= (layer0_outputs(10970)) and (layer0_outputs(4033));
    outputs(2146) <= (layer0_outputs(3979)) or (layer0_outputs(3957));
    outputs(2147) <= not(layer0_outputs(293));
    outputs(2148) <= (layer0_outputs(3638)) and (layer0_outputs(11005));
    outputs(2149) <= not(layer0_outputs(11076));
    outputs(2150) <= (layer0_outputs(11739)) and not (layer0_outputs(3512));
    outputs(2151) <= (layer0_outputs(5326)) xor (layer0_outputs(4858));
    outputs(2152) <= (layer0_outputs(7043)) xor (layer0_outputs(9582));
    outputs(2153) <= not((layer0_outputs(10900)) xor (layer0_outputs(10641)));
    outputs(2154) <= not((layer0_outputs(1194)) xor (layer0_outputs(4211)));
    outputs(2155) <= layer0_outputs(56);
    outputs(2156) <= not((layer0_outputs(9669)) xor (layer0_outputs(10731)));
    outputs(2157) <= (layer0_outputs(7031)) and not (layer0_outputs(9085));
    outputs(2158) <= not((layer0_outputs(4557)) xor (layer0_outputs(4287)));
    outputs(2159) <= not((layer0_outputs(9705)) xor (layer0_outputs(3033)));
    outputs(2160) <= (layer0_outputs(9282)) and not (layer0_outputs(2113));
    outputs(2161) <= not((layer0_outputs(10917)) or (layer0_outputs(11892)));
    outputs(2162) <= not((layer0_outputs(12165)) xor (layer0_outputs(9028)));
    outputs(2163) <= (layer0_outputs(9448)) and (layer0_outputs(10264));
    outputs(2164) <= not(layer0_outputs(12349));
    outputs(2165) <= (layer0_outputs(8032)) and (layer0_outputs(7927));
    outputs(2166) <= (layer0_outputs(126)) and (layer0_outputs(10947));
    outputs(2167) <= (layer0_outputs(10901)) and (layer0_outputs(1398));
    outputs(2168) <= not((layer0_outputs(3264)) xor (layer0_outputs(1387)));
    outputs(2169) <= not((layer0_outputs(7583)) xor (layer0_outputs(3683)));
    outputs(2170) <= not((layer0_outputs(3177)) xor (layer0_outputs(4006)));
    outputs(2171) <= (layer0_outputs(6089)) and not (layer0_outputs(8710));
    outputs(2172) <= (layer0_outputs(5895)) and (layer0_outputs(3454));
    outputs(2173) <= not(layer0_outputs(10142));
    outputs(2174) <= not((layer0_outputs(4499)) xor (layer0_outputs(7448)));
    outputs(2175) <= (layer0_outputs(2543)) xor (layer0_outputs(2879));
    outputs(2176) <= (layer0_outputs(8200)) and not (layer0_outputs(7135));
    outputs(2177) <= not((layer0_outputs(11391)) xor (layer0_outputs(10896)));
    outputs(2178) <= (layer0_outputs(9272)) and not (layer0_outputs(5150));
    outputs(2179) <= (layer0_outputs(5264)) and not (layer0_outputs(10441));
    outputs(2180) <= (layer0_outputs(2293)) and not (layer0_outputs(10349));
    outputs(2181) <= (layer0_outputs(7025)) and not (layer0_outputs(10499));
    outputs(2182) <= (layer0_outputs(3894)) and not (layer0_outputs(6413));
    outputs(2183) <= layer0_outputs(8756);
    outputs(2184) <= (layer0_outputs(5030)) and not (layer0_outputs(8121));
    outputs(2185) <= (layer0_outputs(11065)) xor (layer0_outputs(11011));
    outputs(2186) <= '0';
    outputs(2187) <= (layer0_outputs(6308)) and (layer0_outputs(5294));
    outputs(2188) <= layer0_outputs(1855);
    outputs(2189) <= not(layer0_outputs(1723));
    outputs(2190) <= (layer0_outputs(8002)) xor (layer0_outputs(1666));
    outputs(2191) <= layer0_outputs(3446);
    outputs(2192) <= not(layer0_outputs(3588));
    outputs(2193) <= not(layer0_outputs(11474));
    outputs(2194) <= not(layer0_outputs(12488));
    outputs(2195) <= layer0_outputs(9820);
    outputs(2196) <= (layer0_outputs(9545)) and (layer0_outputs(1781));
    outputs(2197) <= not((layer0_outputs(3923)) xor (layer0_outputs(10022)));
    outputs(2198) <= not((layer0_outputs(12388)) or (layer0_outputs(793)));
    outputs(2199) <= (layer0_outputs(7548)) xor (layer0_outputs(6801));
    outputs(2200) <= not((layer0_outputs(4353)) xor (layer0_outputs(8027)));
    outputs(2201) <= (layer0_outputs(8648)) and (layer0_outputs(11837));
    outputs(2202) <= (layer0_outputs(8705)) and not (layer0_outputs(9053));
    outputs(2203) <= '0';
    outputs(2204) <= (layer0_outputs(11392)) or (layer0_outputs(3799));
    outputs(2205) <= not((layer0_outputs(3630)) xor (layer0_outputs(3213)));
    outputs(2206) <= not((layer0_outputs(5502)) or (layer0_outputs(12313)));
    outputs(2207) <= not((layer0_outputs(1682)) xor (layer0_outputs(5839)));
    outputs(2208) <= (layer0_outputs(1327)) and not (layer0_outputs(10091));
    outputs(2209) <= (layer0_outputs(1599)) and not (layer0_outputs(5724));
    outputs(2210) <= not(layer0_outputs(7757));
    outputs(2211) <= not((layer0_outputs(1962)) xor (layer0_outputs(11341)));
    outputs(2212) <= not(layer0_outputs(2420)) or (layer0_outputs(7630));
    outputs(2213) <= not((layer0_outputs(11881)) xor (layer0_outputs(1754)));
    outputs(2214) <= layer0_outputs(7411);
    outputs(2215) <= not(layer0_outputs(11010));
    outputs(2216) <= layer0_outputs(3990);
    outputs(2217) <= (layer0_outputs(9762)) and (layer0_outputs(5632));
    outputs(2218) <= not((layer0_outputs(416)) or (layer0_outputs(4780)));
    outputs(2219) <= not(layer0_outputs(4358));
    outputs(2220) <= not(layer0_outputs(11834));
    outputs(2221) <= not(layer0_outputs(8870));
    outputs(2222) <= (layer0_outputs(10090)) and (layer0_outputs(156));
    outputs(2223) <= layer0_outputs(9173);
    outputs(2224) <= (layer0_outputs(1930)) and (layer0_outputs(9129));
    outputs(2225) <= not((layer0_outputs(10433)) xor (layer0_outputs(76)));
    outputs(2226) <= not((layer0_outputs(11019)) or (layer0_outputs(2241)));
    outputs(2227) <= (layer0_outputs(11888)) xor (layer0_outputs(12022));
    outputs(2228) <= layer0_outputs(5188);
    outputs(2229) <= (layer0_outputs(7862)) and not (layer0_outputs(5210));
    outputs(2230) <= (layer0_outputs(8581)) xor (layer0_outputs(3617));
    outputs(2231) <= not((layer0_outputs(8253)) or (layer0_outputs(12079)));
    outputs(2232) <= not((layer0_outputs(6068)) or (layer0_outputs(9612)));
    outputs(2233) <= layer0_outputs(12199);
    outputs(2234) <= (layer0_outputs(4459)) and (layer0_outputs(5324));
    outputs(2235) <= (layer0_outputs(10054)) and not (layer0_outputs(9789));
    outputs(2236) <= (layer0_outputs(4952)) xor (layer0_outputs(9799));
    outputs(2237) <= (layer0_outputs(10874)) and not (layer0_outputs(4399));
    outputs(2238) <= not((layer0_outputs(8948)) xor (layer0_outputs(8366)));
    outputs(2239) <= layer0_outputs(11578);
    outputs(2240) <= not(layer0_outputs(6412));
    outputs(2241) <= (layer0_outputs(9811)) and not (layer0_outputs(5667));
    outputs(2242) <= (layer0_outputs(2141)) and not (layer0_outputs(7864));
    outputs(2243) <= not(layer0_outputs(5135));
    outputs(2244) <= (layer0_outputs(12701)) xor (layer0_outputs(2657));
    outputs(2245) <= not((layer0_outputs(10552)) or (layer0_outputs(6510)));
    outputs(2246) <= not((layer0_outputs(5185)) xor (layer0_outputs(523)));
    outputs(2247) <= (layer0_outputs(4633)) xor (layer0_outputs(8631));
    outputs(2248) <= layer0_outputs(9345);
    outputs(2249) <= (layer0_outputs(7735)) and (layer0_outputs(3708));
    outputs(2250) <= not((layer0_outputs(12089)) xor (layer0_outputs(6778)));
    outputs(2251) <= (layer0_outputs(8176)) and (layer0_outputs(5513));
    outputs(2252) <= (layer0_outputs(9004)) and not (layer0_outputs(6063));
    outputs(2253) <= (layer0_outputs(4222)) xor (layer0_outputs(11883));
    outputs(2254) <= (layer0_outputs(7062)) and not (layer0_outputs(3213));
    outputs(2255) <= not(layer0_outputs(10978));
    outputs(2256) <= not((layer0_outputs(1369)) or (layer0_outputs(8303)));
    outputs(2257) <= layer0_outputs(5336);
    outputs(2258) <= not((layer0_outputs(2572)) or (layer0_outputs(10775)));
    outputs(2259) <= not((layer0_outputs(5018)) xor (layer0_outputs(1531)));
    outputs(2260) <= not((layer0_outputs(11131)) xor (layer0_outputs(12514)));
    outputs(2261) <= not(layer0_outputs(8453));
    outputs(2262) <= (layer0_outputs(9397)) and (layer0_outputs(9339));
    outputs(2263) <= (layer0_outputs(4446)) xor (layer0_outputs(12772));
    outputs(2264) <= (layer0_outputs(10776)) and (layer0_outputs(6267));
    outputs(2265) <= not((layer0_outputs(5665)) or (layer0_outputs(8445)));
    outputs(2266) <= (layer0_outputs(9668)) and not (layer0_outputs(9125));
    outputs(2267) <= (layer0_outputs(962)) and not (layer0_outputs(4380));
    outputs(2268) <= not(layer0_outputs(8726)) or (layer0_outputs(12180));
    outputs(2269) <= not(layer0_outputs(2520));
    outputs(2270) <= (layer0_outputs(1267)) and not (layer0_outputs(4895));
    outputs(2271) <= not((layer0_outputs(10274)) xor (layer0_outputs(11926)));
    outputs(2272) <= not((layer0_outputs(11620)) xor (layer0_outputs(5776)));
    outputs(2273) <= '0';
    outputs(2274) <= not(layer0_outputs(3912));
    outputs(2275) <= not(layer0_outputs(9722));
    outputs(2276) <= (layer0_outputs(6485)) xor (layer0_outputs(7283));
    outputs(2277) <= '0';
    outputs(2278) <= not((layer0_outputs(6960)) or (layer0_outputs(12236)));
    outputs(2279) <= (layer0_outputs(11240)) xor (layer0_outputs(10754));
    outputs(2280) <= (layer0_outputs(11981)) and not (layer0_outputs(106));
    outputs(2281) <= not((layer0_outputs(7962)) or (layer0_outputs(6769)));
    outputs(2282) <= not((layer0_outputs(7904)) xor (layer0_outputs(7004)));
    outputs(2283) <= '0';
    outputs(2284) <= not(layer0_outputs(12131));
    outputs(2285) <= not((layer0_outputs(2498)) xor (layer0_outputs(4081)));
    outputs(2286) <= not((layer0_outputs(6214)) xor (layer0_outputs(11197)));
    outputs(2287) <= not((layer0_outputs(8315)) or (layer0_outputs(8950)));
    outputs(2288) <= not(layer0_outputs(6890));
    outputs(2289) <= (layer0_outputs(1449)) xor (layer0_outputs(4237));
    outputs(2290) <= (layer0_outputs(905)) xor (layer0_outputs(3035));
    outputs(2291) <= (layer0_outputs(954)) and not (layer0_outputs(12256));
    outputs(2292) <= not((layer0_outputs(1929)) or (layer0_outputs(8541)));
    outputs(2293) <= (layer0_outputs(3774)) and not (layer0_outputs(10209));
    outputs(2294) <= (layer0_outputs(1518)) and not (layer0_outputs(7356));
    outputs(2295) <= layer0_outputs(12202);
    outputs(2296) <= (layer0_outputs(12412)) and not (layer0_outputs(9839));
    outputs(2297) <= (layer0_outputs(5645)) and not (layer0_outputs(5854));
    outputs(2298) <= (layer0_outputs(9855)) xor (layer0_outputs(9823));
    outputs(2299) <= not((layer0_outputs(1920)) xor (layer0_outputs(9968)));
    outputs(2300) <= not((layer0_outputs(7893)) xor (layer0_outputs(6677)));
    outputs(2301) <= (layer0_outputs(5167)) and (layer0_outputs(981));
    outputs(2302) <= layer0_outputs(4878);
    outputs(2303) <= not((layer0_outputs(7295)) or (layer0_outputs(6129)));
    outputs(2304) <= (layer0_outputs(6500)) xor (layer0_outputs(7061));
    outputs(2305) <= not((layer0_outputs(7421)) xor (layer0_outputs(4278)));
    outputs(2306) <= (layer0_outputs(11414)) xor (layer0_outputs(164));
    outputs(2307) <= (layer0_outputs(11843)) xor (layer0_outputs(1052));
    outputs(2308) <= (layer0_outputs(10945)) and not (layer0_outputs(34));
    outputs(2309) <= (layer0_outputs(11224)) and not (layer0_outputs(7187));
    outputs(2310) <= (layer0_outputs(3391)) and not (layer0_outputs(7647));
    outputs(2311) <= not((layer0_outputs(2294)) or (layer0_outputs(9931)));
    outputs(2312) <= not((layer0_outputs(8184)) or (layer0_outputs(3642)));
    outputs(2313) <= (layer0_outputs(6371)) and not (layer0_outputs(11029));
    outputs(2314) <= not(layer0_outputs(2058));
    outputs(2315) <= not(layer0_outputs(6936));
    outputs(2316) <= not((layer0_outputs(8529)) xor (layer0_outputs(4892)));
    outputs(2317) <= (layer0_outputs(21)) and (layer0_outputs(8878));
    outputs(2318) <= not((layer0_outputs(9502)) xor (layer0_outputs(781)));
    outputs(2319) <= layer0_outputs(4845);
    outputs(2320) <= not((layer0_outputs(2086)) and (layer0_outputs(8551)));
    outputs(2321) <= not((layer0_outputs(3937)) xor (layer0_outputs(10236)));
    outputs(2322) <= (layer0_outputs(2872)) xor (layer0_outputs(2834));
    outputs(2323) <= (layer0_outputs(5861)) and not (layer0_outputs(2815));
    outputs(2324) <= (layer0_outputs(5504)) and (layer0_outputs(5741));
    outputs(2325) <= (layer0_outputs(2250)) xor (layer0_outputs(7429));
    outputs(2326) <= layer0_outputs(7106);
    outputs(2327) <= (layer0_outputs(9697)) xor (layer0_outputs(9869));
    outputs(2328) <= not((layer0_outputs(2510)) or (layer0_outputs(3969)));
    outputs(2329) <= not(layer0_outputs(9998));
    outputs(2330) <= (layer0_outputs(7145)) and not (layer0_outputs(8916));
    outputs(2331) <= (layer0_outputs(6876)) xor (layer0_outputs(8641));
    outputs(2332) <= (layer0_outputs(11907)) and not (layer0_outputs(9717));
    outputs(2333) <= (layer0_outputs(11526)) xor (layer0_outputs(7960));
    outputs(2334) <= (layer0_outputs(7228)) and (layer0_outputs(5113));
    outputs(2335) <= (layer0_outputs(542)) and (layer0_outputs(4242));
    outputs(2336) <= not((layer0_outputs(11712)) or (layer0_outputs(9322)));
    outputs(2337) <= not((layer0_outputs(3195)) xor (layer0_outputs(6898)));
    outputs(2338) <= not((layer0_outputs(2074)) xor (layer0_outputs(10114)));
    outputs(2339) <= layer0_outputs(2002);
    outputs(2340) <= not((layer0_outputs(1177)) xor (layer0_outputs(12746)));
    outputs(2341) <= layer0_outputs(1826);
    outputs(2342) <= not((layer0_outputs(7908)) or (layer0_outputs(8233)));
    outputs(2343) <= (layer0_outputs(1539)) and not (layer0_outputs(653));
    outputs(2344) <= (layer0_outputs(8594)) and not (layer0_outputs(8084));
    outputs(2345) <= (layer0_outputs(2121)) xor (layer0_outputs(3927));
    outputs(2346) <= not((layer0_outputs(7839)) or (layer0_outputs(4158)));
    outputs(2347) <= layer0_outputs(3306);
    outputs(2348) <= (layer0_outputs(2127)) and (layer0_outputs(8823));
    outputs(2349) <= (layer0_outputs(8503)) xor (layer0_outputs(1819));
    outputs(2350) <= not(layer0_outputs(4401));
    outputs(2351) <= not((layer0_outputs(1088)) or (layer0_outputs(803)));
    outputs(2352) <= not(layer0_outputs(10471));
    outputs(2353) <= not((layer0_outputs(11669)) xor (layer0_outputs(7605)));
    outputs(2354) <= not(layer0_outputs(11863));
    outputs(2355) <= not((layer0_outputs(6894)) xor (layer0_outputs(3663)));
    outputs(2356) <= (layer0_outputs(10464)) xor (layer0_outputs(2378));
    outputs(2357) <= (layer0_outputs(10621)) xor (layer0_outputs(7343));
    outputs(2358) <= (layer0_outputs(11598)) xor (layer0_outputs(221));
    outputs(2359) <= not((layer0_outputs(6224)) and (layer0_outputs(3523)));
    outputs(2360) <= (layer0_outputs(8614)) and not (layer0_outputs(9543));
    outputs(2361) <= layer0_outputs(9734);
    outputs(2362) <= layer0_outputs(160);
    outputs(2363) <= not(layer0_outputs(10796));
    outputs(2364) <= (layer0_outputs(4773)) and not (layer0_outputs(978));
    outputs(2365) <= (layer0_outputs(4397)) xor (layer0_outputs(9047));
    outputs(2366) <= (layer0_outputs(353)) and not (layer0_outputs(12518));
    outputs(2367) <= not((layer0_outputs(6788)) or (layer0_outputs(6577)));
    outputs(2368) <= not((layer0_outputs(1263)) or (layer0_outputs(1958)));
    outputs(2369) <= not(layer0_outputs(8054));
    outputs(2370) <= not(layer0_outputs(3649));
    outputs(2371) <= (layer0_outputs(2372)) and not (layer0_outputs(4842));
    outputs(2372) <= (layer0_outputs(10846)) xor (layer0_outputs(8678));
    outputs(2373) <= not(layer0_outputs(2025));
    outputs(2374) <= (layer0_outputs(9086)) and (layer0_outputs(2186));
    outputs(2375) <= (layer0_outputs(4811)) and not (layer0_outputs(5330));
    outputs(2376) <= not((layer0_outputs(4157)) or (layer0_outputs(7131)));
    outputs(2377) <= (layer0_outputs(3368)) and not (layer0_outputs(645));
    outputs(2378) <= not((layer0_outputs(3932)) and (layer0_outputs(12682)));
    outputs(2379) <= not((layer0_outputs(2429)) or (layer0_outputs(11673)));
    outputs(2380) <= (layer0_outputs(961)) and not (layer0_outputs(2717));
    outputs(2381) <= (layer0_outputs(8249)) xor (layer0_outputs(8069));
    outputs(2382) <= layer0_outputs(11745);
    outputs(2383) <= not((layer0_outputs(4490)) or (layer0_outputs(9845)));
    outputs(2384) <= (layer0_outputs(1423)) xor (layer0_outputs(108));
    outputs(2385) <= (layer0_outputs(3798)) and not (layer0_outputs(7096));
    outputs(2386) <= (layer0_outputs(8297)) and not (layer0_outputs(9131));
    outputs(2387) <= (layer0_outputs(11850)) and (layer0_outputs(3257));
    outputs(2388) <= layer0_outputs(10127);
    outputs(2389) <= (layer0_outputs(1889)) and not (layer0_outputs(2388));
    outputs(2390) <= (layer0_outputs(2385)) xor (layer0_outputs(9756));
    outputs(2391) <= not((layer0_outputs(5719)) or (layer0_outputs(9302)));
    outputs(2392) <= not((layer0_outputs(9146)) xor (layer0_outputs(6941)));
    outputs(2393) <= not((layer0_outputs(3129)) xor (layer0_outputs(1882)));
    outputs(2394) <= not((layer0_outputs(8866)) or (layer0_outputs(10297)));
    outputs(2395) <= not((layer0_outputs(11787)) or (layer0_outputs(9530)));
    outputs(2396) <= (layer0_outputs(8812)) and (layer0_outputs(90));
    outputs(2397) <= (layer0_outputs(726)) and (layer0_outputs(2854));
    outputs(2398) <= not(layer0_outputs(8556));
    outputs(2399) <= not((layer0_outputs(9699)) or (layer0_outputs(10936)));
    outputs(2400) <= (layer0_outputs(2285)) and not (layer0_outputs(3595));
    outputs(2401) <= (layer0_outputs(2428)) xor (layer0_outputs(5960));
    outputs(2402) <= not(layer0_outputs(507));
    outputs(2403) <= not(layer0_outputs(1830));
    outputs(2404) <= (layer0_outputs(5025)) and not (layer0_outputs(9285));
    outputs(2405) <= (layer0_outputs(8181)) xor (layer0_outputs(10735));
    outputs(2406) <= not(layer0_outputs(11983)) or (layer0_outputs(3687));
    outputs(2407) <= not(layer0_outputs(319));
    outputs(2408) <= (layer0_outputs(7994)) and not (layer0_outputs(676));
    outputs(2409) <= not((layer0_outputs(2891)) or (layer0_outputs(3827)));
    outputs(2410) <= not((layer0_outputs(3741)) or (layer0_outputs(11729)));
    outputs(2411) <= layer0_outputs(6709);
    outputs(2412) <= not(layer0_outputs(1610));
    outputs(2413) <= (layer0_outputs(5007)) and (layer0_outputs(2170));
    outputs(2414) <= not(layer0_outputs(2131));
    outputs(2415) <= not(layer0_outputs(8994));
    outputs(2416) <= (layer0_outputs(8901)) and not (layer0_outputs(4209));
    outputs(2417) <= not((layer0_outputs(8510)) or (layer0_outputs(11452)));
    outputs(2418) <= (layer0_outputs(3175)) xor (layer0_outputs(6272));
    outputs(2419) <= layer0_outputs(11191);
    outputs(2420) <= (layer0_outputs(4079)) and not (layer0_outputs(11955));
    outputs(2421) <= layer0_outputs(6432);
    outputs(2422) <= (layer0_outputs(3946)) xor (layer0_outputs(4916));
    outputs(2423) <= layer0_outputs(4817);
    outputs(2424) <= (layer0_outputs(12251)) and not (layer0_outputs(1555));
    outputs(2425) <= not(layer0_outputs(11560));
    outputs(2426) <= layer0_outputs(12470);
    outputs(2427) <= not((layer0_outputs(12187)) xor (layer0_outputs(9642)));
    outputs(2428) <= not((layer0_outputs(7509)) or (layer0_outputs(8290)));
    outputs(2429) <= (layer0_outputs(1544)) and not (layer0_outputs(3023));
    outputs(2430) <= (layer0_outputs(9909)) xor (layer0_outputs(7409));
    outputs(2431) <= (layer0_outputs(12204)) xor (layer0_outputs(7487));
    outputs(2432) <= (layer0_outputs(6989)) and not (layer0_outputs(1580));
    outputs(2433) <= (layer0_outputs(2783)) and (layer0_outputs(2373));
    outputs(2434) <= not((layer0_outputs(266)) or (layer0_outputs(5518)));
    outputs(2435) <= not(layer0_outputs(8193));
    outputs(2436) <= (layer0_outputs(8129)) and (layer0_outputs(5086));
    outputs(2437) <= not((layer0_outputs(1319)) xor (layer0_outputs(6355)));
    outputs(2438) <= layer0_outputs(1528);
    outputs(2439) <= not((layer0_outputs(8153)) xor (layer0_outputs(11118)));
    outputs(2440) <= (layer0_outputs(165)) xor (layer0_outputs(5918));
    outputs(2441) <= (layer0_outputs(1131)) xor (layer0_outputs(403));
    outputs(2442) <= (layer0_outputs(363)) xor (layer0_outputs(6711));
    outputs(2443) <= not(layer0_outputs(10768));
    outputs(2444) <= not((layer0_outputs(8246)) xor (layer0_outputs(7882)));
    outputs(2445) <= (layer0_outputs(532)) xor (layer0_outputs(618));
    outputs(2446) <= (layer0_outputs(9121)) xor (layer0_outputs(8308));
    outputs(2447) <= (layer0_outputs(7852)) xor (layer0_outputs(1151));
    outputs(2448) <= layer0_outputs(12671);
    outputs(2449) <= (layer0_outputs(2195)) and not (layer0_outputs(1310));
    outputs(2450) <= not((layer0_outputs(12279)) or (layer0_outputs(6901)));
    outputs(2451) <= layer0_outputs(7525);
    outputs(2452) <= (layer0_outputs(1820)) and (layer0_outputs(8448));
    outputs(2453) <= (layer0_outputs(6579)) and (layer0_outputs(9127));
    outputs(2454) <= (layer0_outputs(4393)) xor (layer0_outputs(10287));
    outputs(2455) <= (layer0_outputs(4198)) and not (layer0_outputs(7173));
    outputs(2456) <= (layer0_outputs(6223)) and not (layer0_outputs(9062));
    outputs(2457) <= layer0_outputs(2495);
    outputs(2458) <= layer0_outputs(6031);
    outputs(2459) <= (layer0_outputs(677)) and (layer0_outputs(9108));
    outputs(2460) <= not(layer0_outputs(5399));
    outputs(2461) <= not((layer0_outputs(12077)) xor (layer0_outputs(425)));
    outputs(2462) <= not(layer0_outputs(4338));
    outputs(2463) <= not(layer0_outputs(1491));
    outputs(2464) <= (layer0_outputs(1915)) and not (layer0_outputs(12449));
    outputs(2465) <= (layer0_outputs(9348)) xor (layer0_outputs(5424));
    outputs(2466) <= layer0_outputs(3778);
    outputs(2467) <= not(layer0_outputs(662));
    outputs(2468) <= (layer0_outputs(5731)) and not (layer0_outputs(3889));
    outputs(2469) <= (layer0_outputs(8625)) and not (layer0_outputs(7928));
    outputs(2470) <= not(layer0_outputs(10605));
    outputs(2471) <= (layer0_outputs(1364)) and not (layer0_outputs(10670));
    outputs(2472) <= not((layer0_outputs(1987)) xor (layer0_outputs(728)));
    outputs(2473) <= not(layer0_outputs(7660));
    outputs(2474) <= not((layer0_outputs(8410)) xor (layer0_outputs(4227)));
    outputs(2475) <= (layer0_outputs(12053)) xor (layer0_outputs(1495));
    outputs(2476) <= (layer0_outputs(6274)) and not (layer0_outputs(11660));
    outputs(2477) <= not((layer0_outputs(120)) xor (layer0_outputs(12046)));
    outputs(2478) <= layer0_outputs(7335);
    outputs(2479) <= not(layer0_outputs(1847));
    outputs(2480) <= (layer0_outputs(3994)) and (layer0_outputs(6628));
    outputs(2481) <= layer0_outputs(5006);
    outputs(2482) <= (layer0_outputs(3340)) and not (layer0_outputs(8335));
    outputs(2483) <= not(layer0_outputs(10794));
    outputs(2484) <= not((layer0_outputs(9115)) or (layer0_outputs(7515)));
    outputs(2485) <= (layer0_outputs(3621)) and (layer0_outputs(4293));
    outputs(2486) <= layer0_outputs(1214);
    outputs(2487) <= layer0_outputs(1701);
    outputs(2488) <= not((layer0_outputs(4553)) xor (layer0_outputs(5847)));
    outputs(2489) <= (layer0_outputs(12335)) and not (layer0_outputs(3232));
    outputs(2490) <= layer0_outputs(10355);
    outputs(2491) <= not((layer0_outputs(1804)) xor (layer0_outputs(6404)));
    outputs(2492) <= (layer0_outputs(1964)) and (layer0_outputs(11215));
    outputs(2493) <= (layer0_outputs(4332)) xor (layer0_outputs(7163));
    outputs(2494) <= (layer0_outputs(8869)) and not (layer0_outputs(7032));
    outputs(2495) <= (layer0_outputs(9770)) and (layer0_outputs(10100));
    outputs(2496) <= (layer0_outputs(11507)) and not (layer0_outputs(4230));
    outputs(2497) <= (layer0_outputs(1078)) xor (layer0_outputs(1940));
    outputs(2498) <= not(layer0_outputs(5905));
    outputs(2499) <= (layer0_outputs(7457)) and not (layer0_outputs(12229));
    outputs(2500) <= not(layer0_outputs(7264)) or (layer0_outputs(10229));
    outputs(2501) <= not((layer0_outputs(7667)) xor (layer0_outputs(3283)));
    outputs(2502) <= (layer0_outputs(11242)) and not (layer0_outputs(3595));
    outputs(2503) <= not((layer0_outputs(10201)) xor (layer0_outputs(4579)));
    outputs(2504) <= (layer0_outputs(12116)) xor (layer0_outputs(6459));
    outputs(2505) <= (layer0_outputs(2949)) and (layer0_outputs(6924));
    outputs(2506) <= (layer0_outputs(506)) xor (layer0_outputs(4959));
    outputs(2507) <= (layer0_outputs(1898)) and (layer0_outputs(12200));
    outputs(2508) <= not(layer0_outputs(7156));
    outputs(2509) <= (layer0_outputs(3951)) and (layer0_outputs(2657));
    outputs(2510) <= (layer0_outputs(11328)) and not (layer0_outputs(853));
    outputs(2511) <= (layer0_outputs(10059)) and not (layer0_outputs(708));
    outputs(2512) <= (layer0_outputs(6453)) and not (layer0_outputs(6507));
    outputs(2513) <= '0';
    outputs(2514) <= (layer0_outputs(6116)) xor (layer0_outputs(9009));
    outputs(2515) <= (layer0_outputs(10073)) xor (layer0_outputs(2652));
    outputs(2516) <= (layer0_outputs(5446)) and not (layer0_outputs(6862));
    outputs(2517) <= not((layer0_outputs(10565)) xor (layer0_outputs(7656)));
    outputs(2518) <= not((layer0_outputs(7299)) xor (layer0_outputs(9445)));
    outputs(2519) <= not(layer0_outputs(7450));
    outputs(2520) <= layer0_outputs(8119);
    outputs(2521) <= '0';
    outputs(2522) <= (layer0_outputs(7411)) and (layer0_outputs(3762));
    outputs(2523) <= layer0_outputs(12375);
    outputs(2524) <= not((layer0_outputs(9156)) xor (layer0_outputs(4923)));
    outputs(2525) <= not((layer0_outputs(8299)) xor (layer0_outputs(10713)));
    outputs(2526) <= not((layer0_outputs(8358)) or (layer0_outputs(1402)));
    outputs(2527) <= layer0_outputs(12768);
    outputs(2528) <= not((layer0_outputs(7014)) xor (layer0_outputs(5102)));
    outputs(2529) <= (layer0_outputs(12333)) and not (layer0_outputs(343));
    outputs(2530) <= (layer0_outputs(7654)) and not (layer0_outputs(5781));
    outputs(2531) <= not((layer0_outputs(11651)) xor (layer0_outputs(2943)));
    outputs(2532) <= (layer0_outputs(4956)) and (layer0_outputs(6673));
    outputs(2533) <= (layer0_outputs(4091)) xor (layer0_outputs(2294));
    outputs(2534) <= (layer0_outputs(7519)) and not (layer0_outputs(3125));
    outputs(2535) <= not((layer0_outputs(8227)) xor (layer0_outputs(4862)));
    outputs(2536) <= (layer0_outputs(6217)) and not (layer0_outputs(1067));
    outputs(2537) <= (layer0_outputs(815)) and not (layer0_outputs(11794));
    outputs(2538) <= layer0_outputs(3876);
    outputs(2539) <= (layer0_outputs(11023)) xor (layer0_outputs(12701));
    outputs(2540) <= layer0_outputs(4637);
    outputs(2541) <= (layer0_outputs(10441)) xor (layer0_outputs(3197));
    outputs(2542) <= not(layer0_outputs(5347));
    outputs(2543) <= not(layer0_outputs(5733));
    outputs(2544) <= (layer0_outputs(11884)) and not (layer0_outputs(3134));
    outputs(2545) <= not((layer0_outputs(150)) or (layer0_outputs(10828)));
    outputs(2546) <= (layer0_outputs(2350)) xor (layer0_outputs(11026));
    outputs(2547) <= not((layer0_outputs(7108)) xor (layer0_outputs(5166)));
    outputs(2548) <= layer0_outputs(6675);
    outputs(2549) <= not(layer0_outputs(2670)) or (layer0_outputs(4521));
    outputs(2550) <= not((layer0_outputs(9204)) xor (layer0_outputs(4846)));
    outputs(2551) <= not(layer0_outputs(12765));
    outputs(2552) <= (layer0_outputs(1425)) and not (layer0_outputs(3468));
    outputs(2553) <= layer0_outputs(411);
    outputs(2554) <= (layer0_outputs(5973)) xor (layer0_outputs(198));
    outputs(2555) <= not((layer0_outputs(11206)) xor (layer0_outputs(1918)));
    outputs(2556) <= not((layer0_outputs(12662)) or (layer0_outputs(8055)));
    outputs(2557) <= layer0_outputs(10629);
    outputs(2558) <= (layer0_outputs(9733)) xor (layer0_outputs(7623));
    outputs(2559) <= not(layer0_outputs(57));
    outputs(2560) <= not(layer0_outputs(146));
    outputs(2561) <= layer0_outputs(9319);
    outputs(2562) <= not((layer0_outputs(8928)) xor (layer0_outputs(1687)));
    outputs(2563) <= not(layer0_outputs(10686)) or (layer0_outputs(1199));
    outputs(2564) <= layer0_outputs(4654);
    outputs(2565) <= not((layer0_outputs(5841)) xor (layer0_outputs(8287)));
    outputs(2566) <= not(layer0_outputs(8894));
    outputs(2567) <= not((layer0_outputs(810)) and (layer0_outputs(4314)));
    outputs(2568) <= not(layer0_outputs(12435));
    outputs(2569) <= layer0_outputs(3987);
    outputs(2570) <= not(layer0_outputs(5396));
    outputs(2571) <= (layer0_outputs(3015)) and not (layer0_outputs(2278));
    outputs(2572) <= not(layer0_outputs(11744));
    outputs(2573) <= not(layer0_outputs(910));
    outputs(2574) <= not((layer0_outputs(301)) and (layer0_outputs(6104)));
    outputs(2575) <= (layer0_outputs(11493)) xor (layer0_outputs(9165));
    outputs(2576) <= layer0_outputs(5116);
    outputs(2577) <= layer0_outputs(12565);
    outputs(2578) <= layer0_outputs(11742);
    outputs(2579) <= not((layer0_outputs(1832)) xor (layer0_outputs(6075)));
    outputs(2580) <= (layer0_outputs(4012)) and (layer0_outputs(3886));
    outputs(2581) <= (layer0_outputs(186)) xor (layer0_outputs(6963));
    outputs(2582) <= (layer0_outputs(8010)) and not (layer0_outputs(7189));
    outputs(2583) <= layer0_outputs(10099);
    outputs(2584) <= layer0_outputs(12101);
    outputs(2585) <= not((layer0_outputs(8483)) or (layer0_outputs(5034)));
    outputs(2586) <= not(layer0_outputs(3353));
    outputs(2587) <= (layer0_outputs(9070)) xor (layer0_outputs(725));
    outputs(2588) <= not(layer0_outputs(611));
    outputs(2589) <= (layer0_outputs(8809)) and not (layer0_outputs(4694));
    outputs(2590) <= layer0_outputs(6544);
    outputs(2591) <= not(layer0_outputs(9265)) or (layer0_outputs(11001));
    outputs(2592) <= not(layer0_outputs(7738)) or (layer0_outputs(6306));
    outputs(2593) <= (layer0_outputs(11794)) or (layer0_outputs(347));
    outputs(2594) <= layer0_outputs(10414);
    outputs(2595) <= layer0_outputs(5716);
    outputs(2596) <= not((layer0_outputs(1538)) or (layer0_outputs(8871)));
    outputs(2597) <= (layer0_outputs(11945)) xor (layer0_outputs(10649));
    outputs(2598) <= not((layer0_outputs(10530)) xor (layer0_outputs(6361)));
    outputs(2599) <= (layer0_outputs(947)) or (layer0_outputs(2689));
    outputs(2600) <= not(layer0_outputs(11315));
    outputs(2601) <= not(layer0_outputs(5825));
    outputs(2602) <= not(layer0_outputs(4871));
    outputs(2603) <= not(layer0_outputs(8988));
    outputs(2604) <= not((layer0_outputs(4669)) and (layer0_outputs(11822)));
    outputs(2605) <= (layer0_outputs(11458)) and not (layer0_outputs(711));
    outputs(2606) <= not(layer0_outputs(8346));
    outputs(2607) <= layer0_outputs(2896);
    outputs(2608) <= layer0_outputs(5902);
    outputs(2609) <= (layer0_outputs(8051)) or (layer0_outputs(4854));
    outputs(2610) <= not(layer0_outputs(7452));
    outputs(2611) <= not(layer0_outputs(2609)) or (layer0_outputs(10289));
    outputs(2612) <= layer0_outputs(7849);
    outputs(2613) <= layer0_outputs(1477);
    outputs(2614) <= layer0_outputs(7048);
    outputs(2615) <= not(layer0_outputs(4258)) or (layer0_outputs(3647));
    outputs(2616) <= layer0_outputs(2101);
    outputs(2617) <= not((layer0_outputs(8663)) xor (layer0_outputs(11728)));
    outputs(2618) <= not((layer0_outputs(8960)) xor (layer0_outputs(2740)));
    outputs(2619) <= not((layer0_outputs(3492)) xor (layer0_outputs(12422)));
    outputs(2620) <= layer0_outputs(8553);
    outputs(2621) <= not(layer0_outputs(224));
    outputs(2622) <= not(layer0_outputs(816));
    outputs(2623) <= not((layer0_outputs(2864)) or (layer0_outputs(4437)));
    outputs(2624) <= not((layer0_outputs(5968)) xor (layer0_outputs(8830)));
    outputs(2625) <= not((layer0_outputs(2887)) xor (layer0_outputs(10628)));
    outputs(2626) <= (layer0_outputs(11951)) or (layer0_outputs(9169));
    outputs(2627) <= not(layer0_outputs(5372)) or (layer0_outputs(5066));
    outputs(2628) <= layer0_outputs(4354);
    outputs(2629) <= (layer0_outputs(12237)) or (layer0_outputs(8882));
    outputs(2630) <= layer0_outputs(10034);
    outputs(2631) <= layer0_outputs(5857);
    outputs(2632) <= (layer0_outputs(808)) and (layer0_outputs(3511));
    outputs(2633) <= layer0_outputs(7643);
    outputs(2634) <= not(layer0_outputs(1454));
    outputs(2635) <= not((layer0_outputs(2488)) xor (layer0_outputs(10128)));
    outputs(2636) <= not(layer0_outputs(5485));
    outputs(2637) <= (layer0_outputs(11516)) xor (layer0_outputs(739));
    outputs(2638) <= (layer0_outputs(1577)) or (layer0_outputs(2077));
    outputs(2639) <= (layer0_outputs(9306)) or (layer0_outputs(9090));
    outputs(2640) <= layer0_outputs(12656);
    outputs(2641) <= (layer0_outputs(8934)) or (layer0_outputs(12569));
    outputs(2642) <= not((layer0_outputs(11448)) xor (layer0_outputs(8055)));
    outputs(2643) <= (layer0_outputs(18)) xor (layer0_outputs(558));
    outputs(2644) <= not((layer0_outputs(2156)) xor (layer0_outputs(8287)));
    outputs(2645) <= not(layer0_outputs(8929));
    outputs(2646) <= not((layer0_outputs(9862)) or (layer0_outputs(1409)));
    outputs(2647) <= not((layer0_outputs(370)) or (layer0_outputs(8618)));
    outputs(2648) <= not((layer0_outputs(6798)) or (layer0_outputs(3620)));
    outputs(2649) <= not(layer0_outputs(3270)) or (layer0_outputs(10283));
    outputs(2650) <= (layer0_outputs(11929)) xor (layer0_outputs(10815));
    outputs(2651) <= layer0_outputs(3185);
    outputs(2652) <= not((layer0_outputs(3856)) xor (layer0_outputs(369)));
    outputs(2653) <= layer0_outputs(9236);
    outputs(2654) <= (layer0_outputs(3453)) and not (layer0_outputs(8206));
    outputs(2655) <= not(layer0_outputs(2742));
    outputs(2656) <= not(layer0_outputs(6730));
    outputs(2657) <= layer0_outputs(8739);
    outputs(2658) <= not(layer0_outputs(365));
    outputs(2659) <= layer0_outputs(9605);
    outputs(2660) <= (layer0_outputs(4450)) xor (layer0_outputs(9828));
    outputs(2661) <= (layer0_outputs(942)) and not (layer0_outputs(7447));
    outputs(2662) <= not(layer0_outputs(2624));
    outputs(2663) <= layer0_outputs(2423);
    outputs(2664) <= not((layer0_outputs(8460)) and (layer0_outputs(2614)));
    outputs(2665) <= layer0_outputs(10668);
    outputs(2666) <= not((layer0_outputs(9952)) xor (layer0_outputs(7956)));
    outputs(2667) <= not(layer0_outputs(1515)) or (layer0_outputs(8166));
    outputs(2668) <= (layer0_outputs(9841)) and not (layer0_outputs(8695));
    outputs(2669) <= layer0_outputs(10619);
    outputs(2670) <= layer0_outputs(6719);
    outputs(2671) <= (layer0_outputs(5061)) or (layer0_outputs(6630));
    outputs(2672) <= not((layer0_outputs(7442)) or (layer0_outputs(6125)));
    outputs(2673) <= not(layer0_outputs(10482));
    outputs(2674) <= not(layer0_outputs(1910));
    outputs(2675) <= (layer0_outputs(12480)) xor (layer0_outputs(6589));
    outputs(2676) <= not((layer0_outputs(8807)) or (layer0_outputs(5177)));
    outputs(2677) <= (layer0_outputs(10490)) or (layer0_outputs(11899));
    outputs(2678) <= layer0_outputs(4558);
    outputs(2679) <= not((layer0_outputs(8565)) and (layer0_outputs(8751)));
    outputs(2680) <= not((layer0_outputs(921)) xor (layer0_outputs(5686)));
    outputs(2681) <= (layer0_outputs(2109)) and not (layer0_outputs(5580));
    outputs(2682) <= not(layer0_outputs(7701));
    outputs(2683) <= (layer0_outputs(7337)) xor (layer0_outputs(1431));
    outputs(2684) <= layer0_outputs(8108);
    outputs(2685) <= layer0_outputs(3453);
    outputs(2686) <= not((layer0_outputs(9378)) xor (layer0_outputs(5277)));
    outputs(2687) <= not(layer0_outputs(4352));
    outputs(2688) <= layer0_outputs(9686);
    outputs(2689) <= not(layer0_outputs(3046));
    outputs(2690) <= not(layer0_outputs(6889));
    outputs(2691) <= layer0_outputs(3540);
    outputs(2692) <= not((layer0_outputs(5213)) xor (layer0_outputs(4344)));
    outputs(2693) <= not(layer0_outputs(2545));
    outputs(2694) <= layer0_outputs(3729);
    outputs(2695) <= layer0_outputs(3490);
    outputs(2696) <= (layer0_outputs(99)) and not (layer0_outputs(4215));
    outputs(2697) <= (layer0_outputs(232)) or (layer0_outputs(2608));
    outputs(2698) <= (layer0_outputs(10657)) xor (layer0_outputs(4102));
    outputs(2699) <= (layer0_outputs(2813)) xor (layer0_outputs(11676));
    outputs(2700) <= (layer0_outputs(906)) and not (layer0_outputs(715));
    outputs(2701) <= not((layer0_outputs(2773)) and (layer0_outputs(6729)));
    outputs(2702) <= not(layer0_outputs(11736));
    outputs(2703) <= (layer0_outputs(12093)) or (layer0_outputs(6229));
    outputs(2704) <= not(layer0_outputs(960));
    outputs(2705) <= layer0_outputs(5502);
    outputs(2706) <= (layer0_outputs(3634)) and (layer0_outputs(1285));
    outputs(2707) <= layer0_outputs(3700);
    outputs(2708) <= not((layer0_outputs(11767)) xor (layer0_outputs(1219)));
    outputs(2709) <= not((layer0_outputs(1972)) and (layer0_outputs(310)));
    outputs(2710) <= not(layer0_outputs(8431)) or (layer0_outputs(5416));
    outputs(2711) <= not((layer0_outputs(8925)) xor (layer0_outputs(6659)));
    outputs(2712) <= (layer0_outputs(1931)) and not (layer0_outputs(12028));
    outputs(2713) <= not((layer0_outputs(2396)) or (layer0_outputs(2688)));
    outputs(2714) <= not((layer0_outputs(12230)) xor (layer0_outputs(220)));
    outputs(2715) <= layer0_outputs(11778);
    outputs(2716) <= not((layer0_outputs(4192)) or (layer0_outputs(10429)));
    outputs(2717) <= (layer0_outputs(5605)) and (layer0_outputs(6583));
    outputs(2718) <= not((layer0_outputs(2006)) and (layer0_outputs(2592)));
    outputs(2719) <= not(layer0_outputs(4873));
    outputs(2720) <= (layer0_outputs(2840)) xor (layer0_outputs(7289));
    outputs(2721) <= not((layer0_outputs(7866)) xor (layer0_outputs(748)));
    outputs(2722) <= layer0_outputs(4683);
    outputs(2723) <= layer0_outputs(1960);
    outputs(2724) <= layer0_outputs(4097);
    outputs(2725) <= (layer0_outputs(7733)) and not (layer0_outputs(5700));
    outputs(2726) <= (layer0_outputs(1252)) and not (layer0_outputs(12614));
    outputs(2727) <= not((layer0_outputs(9380)) xor (layer0_outputs(3065)));
    outputs(2728) <= not((layer0_outputs(8721)) and (layer0_outputs(6802)));
    outputs(2729) <= layer0_outputs(1951);
    outputs(2730) <= not(layer0_outputs(11920));
    outputs(2731) <= (layer0_outputs(3215)) xor (layer0_outputs(5462));
    outputs(2732) <= not(layer0_outputs(4640));
    outputs(2733) <= (layer0_outputs(4929)) xor (layer0_outputs(9270));
    outputs(2734) <= layer0_outputs(9719);
    outputs(2735) <= (layer0_outputs(7473)) xor (layer0_outputs(7918));
    outputs(2736) <= (layer0_outputs(1965)) xor (layer0_outputs(11237));
    outputs(2737) <= (layer0_outputs(7949)) and not (layer0_outputs(673));
    outputs(2738) <= not(layer0_outputs(3072));
    outputs(2739) <= (layer0_outputs(6878)) and (layer0_outputs(4939));
    outputs(2740) <= layer0_outputs(3126);
    outputs(2741) <= not(layer0_outputs(2679)) or (layer0_outputs(3979));
    outputs(2742) <= (layer0_outputs(9323)) or (layer0_outputs(4151));
    outputs(2743) <= not(layer0_outputs(7270)) or (layer0_outputs(12048));
    outputs(2744) <= layer0_outputs(11806);
    outputs(2745) <= not(layer0_outputs(11534));
    outputs(2746) <= not(layer0_outputs(1376));
    outputs(2747) <= (layer0_outputs(259)) xor (layer0_outputs(12272));
    outputs(2748) <= (layer0_outputs(1881)) or (layer0_outputs(4460));
    outputs(2749) <= layer0_outputs(11917);
    outputs(2750) <= not((layer0_outputs(5913)) xor (layer0_outputs(6355)));
    outputs(2751) <= layer0_outputs(5257);
    outputs(2752) <= not(layer0_outputs(9005));
    outputs(2753) <= not(layer0_outputs(4768)) or (layer0_outputs(10812));
    outputs(2754) <= (layer0_outputs(9378)) xor (layer0_outputs(8808));
    outputs(2755) <= not((layer0_outputs(7823)) xor (layer0_outputs(7232)));
    outputs(2756) <= not(layer0_outputs(6372));
    outputs(2757) <= not(layer0_outputs(11528));
    outputs(2758) <= (layer0_outputs(8792)) and not (layer0_outputs(7890));
    outputs(2759) <= (layer0_outputs(11525)) and not (layer0_outputs(2560));
    outputs(2760) <= not(layer0_outputs(12192));
    outputs(2761) <= (layer0_outputs(1183)) or (layer0_outputs(9201));
    outputs(2762) <= (layer0_outputs(12562)) xor (layer0_outputs(5663));
    outputs(2763) <= not(layer0_outputs(11207));
    outputs(2764) <= (layer0_outputs(6827)) xor (layer0_outputs(3345));
    outputs(2765) <= (layer0_outputs(11579)) and not (layer0_outputs(9582));
    outputs(2766) <= layer0_outputs(4367);
    outputs(2767) <= not(layer0_outputs(215)) or (layer0_outputs(8820));
    outputs(2768) <= layer0_outputs(11841);
    outputs(2769) <= not((layer0_outputs(7200)) xor (layer0_outputs(6930)));
    outputs(2770) <= not(layer0_outputs(4920));
    outputs(2771) <= not((layer0_outputs(2287)) xor (layer0_outputs(427)));
    outputs(2772) <= not(layer0_outputs(6810)) or (layer0_outputs(182));
    outputs(2773) <= (layer0_outputs(6341)) and not (layer0_outputs(2505));
    outputs(2774) <= not(layer0_outputs(7132));
    outputs(2775) <= layer0_outputs(5814);
    outputs(2776) <= not(layer0_outputs(12319));
    outputs(2777) <= (layer0_outputs(10771)) and not (layer0_outputs(3908));
    outputs(2778) <= (layer0_outputs(9083)) and not (layer0_outputs(11208));
    outputs(2779) <= (layer0_outputs(1549)) and (layer0_outputs(8641));
    outputs(2780) <= not(layer0_outputs(4988)) or (layer0_outputs(12620));
    outputs(2781) <= not(layer0_outputs(7313));
    outputs(2782) <= not(layer0_outputs(4165));
    outputs(2783) <= not(layer0_outputs(8393)) or (layer0_outputs(4612));
    outputs(2784) <= not(layer0_outputs(6094)) or (layer0_outputs(4892));
    outputs(2785) <= not((layer0_outputs(6226)) xor (layer0_outputs(4514)));
    outputs(2786) <= layer0_outputs(9585);
    outputs(2787) <= not((layer0_outputs(763)) or (layer0_outputs(4501)));
    outputs(2788) <= (layer0_outputs(3614)) and not (layer0_outputs(6909));
    outputs(2789) <= not((layer0_outputs(2229)) and (layer0_outputs(8729)));
    outputs(2790) <= not((layer0_outputs(5348)) and (layer0_outputs(8679)));
    outputs(2791) <= not(layer0_outputs(7768));
    outputs(2792) <= (layer0_outputs(11401)) xor (layer0_outputs(12503));
    outputs(2793) <= (layer0_outputs(9616)) and not (layer0_outputs(4032));
    outputs(2794) <= layer0_outputs(6032);
    outputs(2795) <= layer0_outputs(6565);
    outputs(2796) <= not((layer0_outputs(12304)) xor (layer0_outputs(7080)));
    outputs(2797) <= not(layer0_outputs(399));
    outputs(2798) <= not(layer0_outputs(2233)) or (layer0_outputs(9698));
    outputs(2799) <= layer0_outputs(3575);
    outputs(2800) <= not((layer0_outputs(5259)) xor (layer0_outputs(7644)));
    outputs(2801) <= not(layer0_outputs(5622));
    outputs(2802) <= (layer0_outputs(11400)) and not (layer0_outputs(1872));
    outputs(2803) <= not((layer0_outputs(8625)) xor (layer0_outputs(7268)));
    outputs(2804) <= not((layer0_outputs(1613)) or (layer0_outputs(11289)));
    outputs(2805) <= layer0_outputs(4975);
    outputs(2806) <= not(layer0_outputs(1176));
    outputs(2807) <= (layer0_outputs(12577)) and (layer0_outputs(10969));
    outputs(2808) <= not(layer0_outputs(7263)) or (layer0_outputs(9666));
    outputs(2809) <= (layer0_outputs(12788)) or (layer0_outputs(4545));
    outputs(2810) <= (layer0_outputs(12003)) or (layer0_outputs(545));
    outputs(2811) <= not((layer0_outputs(2219)) and (layer0_outputs(10167)));
    outputs(2812) <= layer0_outputs(4809);
    outputs(2813) <= not(layer0_outputs(550));
    outputs(2814) <= not((layer0_outputs(5206)) and (layer0_outputs(9110)));
    outputs(2815) <= not(layer0_outputs(2591));
    outputs(2816) <= not((layer0_outputs(3573)) xor (layer0_outputs(11367)));
    outputs(2817) <= not(layer0_outputs(281));
    outputs(2818) <= layer0_outputs(4153);
    outputs(2819) <= (layer0_outputs(9538)) xor (layer0_outputs(6337));
    outputs(2820) <= not(layer0_outputs(486)) or (layer0_outputs(12551));
    outputs(2821) <= not(layer0_outputs(11031));
    outputs(2822) <= not(layer0_outputs(6218));
    outputs(2823) <= (layer0_outputs(6641)) xor (layer0_outputs(4528));
    outputs(2824) <= not((layer0_outputs(8049)) xor (layer0_outputs(4040)));
    outputs(2825) <= not(layer0_outputs(7256)) or (layer0_outputs(7996));
    outputs(2826) <= (layer0_outputs(6680)) and not (layer0_outputs(479));
    outputs(2827) <= not(layer0_outputs(2247)) or (layer0_outputs(10424));
    outputs(2828) <= not((layer0_outputs(33)) xor (layer0_outputs(4601)));
    outputs(2829) <= not(layer0_outputs(7283));
    outputs(2830) <= not(layer0_outputs(571));
    outputs(2831) <= not(layer0_outputs(3855)) or (layer0_outputs(466));
    outputs(2832) <= not(layer0_outputs(5919)) or (layer0_outputs(8264));
    outputs(2833) <= layer0_outputs(12580);
    outputs(2834) <= not(layer0_outputs(2686));
    outputs(2835) <= not(layer0_outputs(3025)) or (layer0_outputs(8926));
    outputs(2836) <= not((layer0_outputs(7286)) xor (layer0_outputs(303)));
    outputs(2837) <= not(layer0_outputs(3899));
    outputs(2838) <= not(layer0_outputs(4325)) or (layer0_outputs(469));
    outputs(2839) <= (layer0_outputs(11067)) and not (layer0_outputs(8403));
    outputs(2840) <= not(layer0_outputs(7780));
    outputs(2841) <= (layer0_outputs(10698)) xor (layer0_outputs(127));
    outputs(2842) <= layer0_outputs(8681);
    outputs(2843) <= not(layer0_outputs(3107));
    outputs(2844) <= (layer0_outputs(3530)) xor (layer0_outputs(10775));
    outputs(2845) <= layer0_outputs(4734);
    outputs(2846) <= not(layer0_outputs(10387));
    outputs(2847) <= not(layer0_outputs(11200));
    outputs(2848) <= layer0_outputs(12167);
    outputs(2849) <= not(layer0_outputs(3032));
    outputs(2850) <= not((layer0_outputs(1892)) xor (layer0_outputs(5409)));
    outputs(2851) <= layer0_outputs(12341);
    outputs(2852) <= not(layer0_outputs(9360));
    outputs(2853) <= (layer0_outputs(1362)) xor (layer0_outputs(4772));
    outputs(2854) <= (layer0_outputs(10748)) xor (layer0_outputs(9318));
    outputs(2855) <= not(layer0_outputs(9526)) or (layer0_outputs(9733));
    outputs(2856) <= (layer0_outputs(12534)) xor (layer0_outputs(7352));
    outputs(2857) <= not(layer0_outputs(9475));
    outputs(2858) <= (layer0_outputs(409)) xor (layer0_outputs(5091));
    outputs(2859) <= not(layer0_outputs(9186)) or (layer0_outputs(7017));
    outputs(2860) <= (layer0_outputs(5551)) or (layer0_outputs(11183));
    outputs(2861) <= (layer0_outputs(7095)) and (layer0_outputs(2063));
    outputs(2862) <= not((layer0_outputs(10325)) xor (layer0_outputs(7777)));
    outputs(2863) <= not((layer0_outputs(5874)) xor (layer0_outputs(8245)));
    outputs(2864) <= (layer0_outputs(7211)) or (layer0_outputs(459));
    outputs(2865) <= not(layer0_outputs(6043));
    outputs(2866) <= not((layer0_outputs(12526)) and (layer0_outputs(1710)));
    outputs(2867) <= (layer0_outputs(2192)) or (layer0_outputs(3537));
    outputs(2868) <= not((layer0_outputs(888)) xor (layer0_outputs(4256)));
    outputs(2869) <= (layer0_outputs(607)) xor (layer0_outputs(5402));
    outputs(2870) <= not(layer0_outputs(4537));
    outputs(2871) <= not(layer0_outputs(5869));
    outputs(2872) <= not((layer0_outputs(6407)) and (layer0_outputs(5277)));
    outputs(2873) <= layer0_outputs(7761);
    outputs(2874) <= not(layer0_outputs(2476)) or (layer0_outputs(10656));
    outputs(2875) <= not(layer0_outputs(4732));
    outputs(2876) <= '1';
    outputs(2877) <= not((layer0_outputs(9163)) xor (layer0_outputs(3395)));
    outputs(2878) <= (layer0_outputs(10023)) and not (layer0_outputs(4216));
    outputs(2879) <= not((layer0_outputs(7819)) xor (layer0_outputs(7338)));
    outputs(2880) <= (layer0_outputs(3483)) and not (layer0_outputs(4505));
    outputs(2881) <= not(layer0_outputs(2982));
    outputs(2882) <= not((layer0_outputs(1693)) or (layer0_outputs(11229)));
    outputs(2883) <= (layer0_outputs(7415)) xor (layer0_outputs(11489));
    outputs(2884) <= not((layer0_outputs(9532)) xor (layer0_outputs(6173)));
    outputs(2885) <= layer0_outputs(2858);
    outputs(2886) <= not((layer0_outputs(4156)) xor (layer0_outputs(8643)));
    outputs(2887) <= not(layer0_outputs(10088));
    outputs(2888) <= (layer0_outputs(4046)) and not (layer0_outputs(7023));
    outputs(2889) <= layer0_outputs(9444);
    outputs(2890) <= not(layer0_outputs(284)) or (layer0_outputs(10076));
    outputs(2891) <= not((layer0_outputs(7381)) or (layer0_outputs(4876)));
    outputs(2892) <= not(layer0_outputs(5458)) or (layer0_outputs(12577));
    outputs(2893) <= (layer0_outputs(5301)) and not (layer0_outputs(5262));
    outputs(2894) <= (layer0_outputs(4084)) and not (layer0_outputs(4908));
    outputs(2895) <= not(layer0_outputs(6144));
    outputs(2896) <= not(layer0_outputs(10959));
    outputs(2897) <= layer0_outputs(10278);
    outputs(2898) <= layer0_outputs(10124);
    outputs(2899) <= (layer0_outputs(9818)) xor (layer0_outputs(10879));
    outputs(2900) <= not((layer0_outputs(195)) xor (layer0_outputs(6468)));
    outputs(2901) <= not(layer0_outputs(7841)) or (layer0_outputs(6070));
    outputs(2902) <= not(layer0_outputs(4448)) or (layer0_outputs(12208));
    outputs(2903) <= not(layer0_outputs(6839)) or (layer0_outputs(1163));
    outputs(2904) <= not((layer0_outputs(5658)) xor (layer0_outputs(10970)));
    outputs(2905) <= not((layer0_outputs(6218)) or (layer0_outputs(1767)));
    outputs(2906) <= layer0_outputs(4659);
    outputs(2907) <= (layer0_outputs(6490)) xor (layer0_outputs(10753));
    outputs(2908) <= (layer0_outputs(9687)) or (layer0_outputs(1602));
    outputs(2909) <= not((layer0_outputs(9036)) xor (layer0_outputs(2239)));
    outputs(2910) <= not((layer0_outputs(7805)) xor (layer0_outputs(6195)));
    outputs(2911) <= not(layer0_outputs(10080)) or (layer0_outputs(1446));
    outputs(2912) <= not(layer0_outputs(8701)) or (layer0_outputs(751));
    outputs(2913) <= (layer0_outputs(10302)) and not (layer0_outputs(6490));
    outputs(2914) <= (layer0_outputs(4449)) or (layer0_outputs(5495));
    outputs(2915) <= not((layer0_outputs(2518)) and (layer0_outputs(6498)));
    outputs(2916) <= not((layer0_outputs(2662)) xor (layer0_outputs(10479)));
    outputs(2917) <= not((layer0_outputs(12640)) xor (layer0_outputs(960)));
    outputs(2918) <= not(layer0_outputs(11556));
    outputs(2919) <= (layer0_outputs(2277)) and (layer0_outputs(1526));
    outputs(2920) <= not((layer0_outputs(10759)) xor (layer0_outputs(6367)));
    outputs(2921) <= not(layer0_outputs(12233));
    outputs(2922) <= layer0_outputs(10225);
    outputs(2923) <= not(layer0_outputs(7595)) or (layer0_outputs(6708));
    outputs(2924) <= not(layer0_outputs(11675));
    outputs(2925) <= not((layer0_outputs(4489)) or (layer0_outputs(3607)));
    outputs(2926) <= not(layer0_outputs(1050));
    outputs(2927) <= (layer0_outputs(6117)) xor (layer0_outputs(4714));
    outputs(2928) <= not(layer0_outputs(1484));
    outputs(2929) <= layer0_outputs(5012);
    outputs(2930) <= not(layer0_outputs(4873));
    outputs(2931) <= not(layer0_outputs(7780));
    outputs(2932) <= not(layer0_outputs(1692));
    outputs(2933) <= (layer0_outputs(4244)) or (layer0_outputs(9593));
    outputs(2934) <= (layer0_outputs(8407)) or (layer0_outputs(519));
    outputs(2935) <= not((layer0_outputs(9095)) xor (layer0_outputs(11145)));
    outputs(2936) <= not(layer0_outputs(9078));
    outputs(2937) <= not((layer0_outputs(1291)) or (layer0_outputs(713)));
    outputs(2938) <= not(layer0_outputs(2276));
    outputs(2939) <= not(layer0_outputs(9154)) or (layer0_outputs(12504));
    outputs(2940) <= not((layer0_outputs(8778)) or (layer0_outputs(7438)));
    outputs(2941) <= (layer0_outputs(10688)) or (layer0_outputs(11301));
    outputs(2942) <= layer0_outputs(11768);
    outputs(2943) <= layer0_outputs(12057);
    outputs(2944) <= (layer0_outputs(7769)) xor (layer0_outputs(4673));
    outputs(2945) <= (layer0_outputs(9850)) or (layer0_outputs(9300));
    outputs(2946) <= layer0_outputs(10600);
    outputs(2947) <= not(layer0_outputs(3090)) or (layer0_outputs(3406));
    outputs(2948) <= not(layer0_outputs(3989));
    outputs(2949) <= not(layer0_outputs(2017));
    outputs(2950) <= layer0_outputs(9178);
    outputs(2951) <= layer0_outputs(5423);
    outputs(2952) <= not(layer0_outputs(513)) or (layer0_outputs(10941));
    outputs(2953) <= (layer0_outputs(3225)) xor (layer0_outputs(6383));
    outputs(2954) <= layer0_outputs(8481);
    outputs(2955) <= not((layer0_outputs(12265)) and (layer0_outputs(860)));
    outputs(2956) <= not((layer0_outputs(8332)) and (layer0_outputs(8586)));
    outputs(2957) <= (layer0_outputs(7480)) and not (layer0_outputs(11886));
    outputs(2958) <= not((layer0_outputs(3485)) xor (layer0_outputs(3455)));
    outputs(2959) <= (layer0_outputs(8371)) or (layer0_outputs(11573));
    outputs(2960) <= (layer0_outputs(3600)) or (layer0_outputs(7787));
    outputs(2961) <= layer0_outputs(6308);
    outputs(2962) <= not((layer0_outputs(11382)) xor (layer0_outputs(4128)));
    outputs(2963) <= not(layer0_outputs(11541));
    outputs(2964) <= not((layer0_outputs(167)) or (layer0_outputs(9191)));
    outputs(2965) <= not(layer0_outputs(792));
    outputs(2966) <= (layer0_outputs(758)) or (layer0_outputs(8573));
    outputs(2967) <= not(layer0_outputs(5292)) or (layer0_outputs(1453));
    outputs(2968) <= (layer0_outputs(4245)) xor (layer0_outputs(3478));
    outputs(2969) <= (layer0_outputs(1290)) and not (layer0_outputs(11957));
    outputs(2970) <= not((layer0_outputs(11853)) xor (layer0_outputs(172)));
    outputs(2971) <= (layer0_outputs(564)) xor (layer0_outputs(10068));
    outputs(2972) <= (layer0_outputs(2760)) or (layer0_outputs(6811));
    outputs(2973) <= not((layer0_outputs(9253)) xor (layer0_outputs(10811)));
    outputs(2974) <= not(layer0_outputs(5395)) or (layer0_outputs(9227));
    outputs(2975) <= not((layer0_outputs(6281)) xor (layer0_outputs(12682)));
    outputs(2976) <= not(layer0_outputs(9221));
    outputs(2977) <= not((layer0_outputs(11936)) or (layer0_outputs(8140)));
    outputs(2978) <= layer0_outputs(3567);
    outputs(2979) <= layer0_outputs(11500);
    outputs(2980) <= layer0_outputs(1843);
    outputs(2981) <= not(layer0_outputs(12799));
    outputs(2982) <= (layer0_outputs(6095)) xor (layer0_outputs(12063));
    outputs(2983) <= layer0_outputs(2886);
    outputs(2984) <= (layer0_outputs(467)) and not (layer0_outputs(8385));
    outputs(2985) <= (layer0_outputs(10813)) or (layer0_outputs(11399));
    outputs(2986) <= (layer0_outputs(12051)) xor (layer0_outputs(10920));
    outputs(2987) <= not((layer0_outputs(12757)) and (layer0_outputs(8637)));
    outputs(2988) <= (layer0_outputs(2279)) or (layer0_outputs(10438));
    outputs(2989) <= not(layer0_outputs(6660)) or (layer0_outputs(3830));
    outputs(2990) <= not((layer0_outputs(4246)) xor (layer0_outputs(10768)));
    outputs(2991) <= (layer0_outputs(1617)) xor (layer0_outputs(4419));
    outputs(2992) <= not(layer0_outputs(7755));
    outputs(2993) <= not((layer0_outputs(9363)) xor (layer0_outputs(2861)));
    outputs(2994) <= not((layer0_outputs(7065)) xor (layer0_outputs(2940)));
    outputs(2995) <= not(layer0_outputs(3889)) or (layer0_outputs(5559));
    outputs(2996) <= layer0_outputs(12300);
    outputs(2997) <= (layer0_outputs(7195)) and not (layer0_outputs(7273));
    outputs(2998) <= layer0_outputs(11292);
    outputs(2999) <= (layer0_outputs(2782)) or (layer0_outputs(6512));
    outputs(3000) <= not(layer0_outputs(7512));
    outputs(3001) <= (layer0_outputs(7971)) and not (layer0_outputs(3910));
    outputs(3002) <= not((layer0_outputs(6498)) and (layer0_outputs(882)));
    outputs(3003) <= not(layer0_outputs(4185));
    outputs(3004) <= not((layer0_outputs(5245)) and (layer0_outputs(8748)));
    outputs(3005) <= layer0_outputs(11592);
    outputs(3006) <= not(layer0_outputs(585));
    outputs(3007) <= not(layer0_outputs(214));
    outputs(3008) <= not((layer0_outputs(8665)) xor (layer0_outputs(5395)));
    outputs(3009) <= not((layer0_outputs(3693)) xor (layer0_outputs(11946)));
    outputs(3010) <= not(layer0_outputs(5400));
    outputs(3011) <= not((layer0_outputs(4680)) and (layer0_outputs(8974)));
    outputs(3012) <= not((layer0_outputs(5216)) xor (layer0_outputs(9192)));
    outputs(3013) <= not(layer0_outputs(11344));
    outputs(3014) <= not(layer0_outputs(6489)) or (layer0_outputs(12138));
    outputs(3015) <= layer0_outputs(1322);
    outputs(3016) <= layer0_outputs(5863);
    outputs(3017) <= not((layer0_outputs(5069)) xor (layer0_outputs(1792)));
    outputs(3018) <= not(layer0_outputs(9661));
    outputs(3019) <= (layer0_outputs(10253)) or (layer0_outputs(12467));
    outputs(3020) <= (layer0_outputs(1036)) and not (layer0_outputs(4649));
    outputs(3021) <= (layer0_outputs(9846)) or (layer0_outputs(3509));
    outputs(3022) <= (layer0_outputs(2176)) and (layer0_outputs(5809));
    outputs(3023) <= layer0_outputs(10749);
    outputs(3024) <= not(layer0_outputs(2743));
    outputs(3025) <= (layer0_outputs(10235)) and not (layer0_outputs(5862));
    outputs(3026) <= (layer0_outputs(10189)) and (layer0_outputs(7278));
    outputs(3027) <= not(layer0_outputs(2865)) or (layer0_outputs(3460));
    outputs(3028) <= not(layer0_outputs(7896)) or (layer0_outputs(5316));
    outputs(3029) <= not((layer0_outputs(12774)) xor (layer0_outputs(9783)));
    outputs(3030) <= (layer0_outputs(6332)) and not (layer0_outputs(6887));
    outputs(3031) <= not(layer0_outputs(3797)) or (layer0_outputs(283));
    outputs(3032) <= not((layer0_outputs(4897)) xor (layer0_outputs(9629)));
    outputs(3033) <= not(layer0_outputs(2685)) or (layer0_outputs(4086));
    outputs(3034) <= not((layer0_outputs(8)) and (layer0_outputs(10857)));
    outputs(3035) <= (layer0_outputs(11297)) xor (layer0_outputs(8902));
    outputs(3036) <= (layer0_outputs(2703)) xor (layer0_outputs(10634));
    outputs(3037) <= (layer0_outputs(7476)) xor (layer0_outputs(4317));
    outputs(3038) <= (layer0_outputs(12154)) and not (layer0_outputs(1370));
    outputs(3039) <= layer0_outputs(11402);
    outputs(3040) <= not(layer0_outputs(1169));
    outputs(3041) <= not(layer0_outputs(6251));
    outputs(3042) <= not(layer0_outputs(2281));
    outputs(3043) <= (layer0_outputs(12120)) or (layer0_outputs(620));
    outputs(3044) <= not(layer0_outputs(4872));
    outputs(3045) <= (layer0_outputs(7937)) and not (layer0_outputs(848));
    outputs(3046) <= layer0_outputs(6951);
    outputs(3047) <= not(layer0_outputs(11541));
    outputs(3048) <= not(layer0_outputs(9642));
    outputs(3049) <= layer0_outputs(11652);
    outputs(3050) <= layer0_outputs(2960);
    outputs(3051) <= (layer0_outputs(6309)) xor (layer0_outputs(5241));
    outputs(3052) <= (layer0_outputs(5373)) xor (layer0_outputs(10999));
    outputs(3053) <= not((layer0_outputs(7910)) xor (layer0_outputs(7105)));
    outputs(3054) <= not(layer0_outputs(8)) or (layer0_outputs(12249));
    outputs(3055) <= not((layer0_outputs(6075)) and (layer0_outputs(9428)));
    outputs(3056) <= not(layer0_outputs(1050));
    outputs(3057) <= not(layer0_outputs(7714));
    outputs(3058) <= not(layer0_outputs(1311)) or (layer0_outputs(7147));
    outputs(3059) <= (layer0_outputs(5726)) xor (layer0_outputs(6892));
    outputs(3060) <= (layer0_outputs(2358)) xor (layer0_outputs(11033));
    outputs(3061) <= layer0_outputs(2423);
    outputs(3062) <= not(layer0_outputs(5062));
    outputs(3063) <= not((layer0_outputs(9434)) and (layer0_outputs(12431)));
    outputs(3064) <= layer0_outputs(12672);
    outputs(3065) <= not((layer0_outputs(6947)) xor (layer0_outputs(25)));
    outputs(3066) <= layer0_outputs(8089);
    outputs(3067) <= (layer0_outputs(5818)) xor (layer0_outputs(11057));
    outputs(3068) <= not(layer0_outputs(8397));
    outputs(3069) <= not(layer0_outputs(3804)) or (layer0_outputs(10151));
    outputs(3070) <= not((layer0_outputs(12679)) and (layer0_outputs(11186)));
    outputs(3071) <= (layer0_outputs(12122)) or (layer0_outputs(4749));
    outputs(3072) <= not(layer0_outputs(4442));
    outputs(3073) <= not((layer0_outputs(4913)) or (layer0_outputs(9241)));
    outputs(3074) <= not((layer0_outputs(5820)) xor (layer0_outputs(2089)));
    outputs(3075) <= layer0_outputs(11081);
    outputs(3076) <= not(layer0_outputs(12235));
    outputs(3077) <= not((layer0_outputs(4964)) or (layer0_outputs(151)));
    outputs(3078) <= not(layer0_outputs(7706));
    outputs(3079) <= not((layer0_outputs(1484)) or (layer0_outputs(11522)));
    outputs(3080) <= (layer0_outputs(6554)) and (layer0_outputs(4243));
    outputs(3081) <= not(layer0_outputs(1921));
    outputs(3082) <= not((layer0_outputs(1147)) xor (layer0_outputs(10922)));
    outputs(3083) <= (layer0_outputs(2946)) or (layer0_outputs(4541));
    outputs(3084) <= (layer0_outputs(12564)) xor (layer0_outputs(8043));
    outputs(3085) <= not(layer0_outputs(6567));
    outputs(3086) <= (layer0_outputs(8753)) and not (layer0_outputs(12794));
    outputs(3087) <= layer0_outputs(5823);
    outputs(3088) <= not(layer0_outputs(3863));
    outputs(3089) <= not((layer0_outputs(4583)) xor (layer0_outputs(12710)));
    outputs(3090) <= not((layer0_outputs(4918)) or (layer0_outputs(6325)));
    outputs(3091) <= layer0_outputs(7741);
    outputs(3092) <= not(layer0_outputs(8823));
    outputs(3093) <= not(layer0_outputs(7809));
    outputs(3094) <= not(layer0_outputs(11596)) or (layer0_outputs(8143));
    outputs(3095) <= not(layer0_outputs(1784));
    outputs(3096) <= (layer0_outputs(5573)) or (layer0_outputs(8398));
    outputs(3097) <= not(layer0_outputs(6938)) or (layer0_outputs(9861));
    outputs(3098) <= not(layer0_outputs(9551));
    outputs(3099) <= (layer0_outputs(1645)) and not (layer0_outputs(5432));
    outputs(3100) <= (layer0_outputs(7198)) or (layer0_outputs(4370));
    outputs(3101) <= not(layer0_outputs(12418));
    outputs(3102) <= layer0_outputs(8769);
    outputs(3103) <= not((layer0_outputs(10924)) xor (layer0_outputs(6691)));
    outputs(3104) <= not(layer0_outputs(11527));
    outputs(3105) <= not((layer0_outputs(8485)) and (layer0_outputs(117)));
    outputs(3106) <= layer0_outputs(3409);
    outputs(3107) <= layer0_outputs(1778);
    outputs(3108) <= layer0_outputs(12694);
    outputs(3109) <= (layer0_outputs(7710)) or (layer0_outputs(10212));
    outputs(3110) <= (layer0_outputs(260)) xor (layer0_outputs(499));
    outputs(3111) <= not((layer0_outputs(6851)) and (layer0_outputs(682)));
    outputs(3112) <= layer0_outputs(6228);
    outputs(3113) <= not(layer0_outputs(1601)) or (layer0_outputs(2913));
    outputs(3114) <= not((layer0_outputs(7152)) or (layer0_outputs(8209)));
    outputs(3115) <= not(layer0_outputs(4386)) or (layer0_outputs(3502));
    outputs(3116) <= not((layer0_outputs(1396)) xor (layer0_outputs(8154)));
    outputs(3117) <= not((layer0_outputs(7839)) xor (layer0_outputs(4233)));
    outputs(3118) <= layer0_outputs(3071);
    outputs(3119) <= not((layer0_outputs(9225)) and (layer0_outputs(4967)));
    outputs(3120) <= (layer0_outputs(6431)) and not (layer0_outputs(4726));
    outputs(3121) <= layer0_outputs(12025);
    outputs(3122) <= (layer0_outputs(833)) or (layer0_outputs(9746));
    outputs(3123) <= (layer0_outputs(6773)) xor (layer0_outputs(382));
    outputs(3124) <= not(layer0_outputs(11902));
    outputs(3125) <= layer0_outputs(12370);
    outputs(3126) <= not((layer0_outputs(5278)) or (layer0_outputs(6402)));
    outputs(3127) <= layer0_outputs(3869);
    outputs(3128) <= (layer0_outputs(10298)) xor (layer0_outputs(1189));
    outputs(3129) <= layer0_outputs(2983);
    outputs(3130) <= layer0_outputs(8884);
    outputs(3131) <= layer0_outputs(5148);
    outputs(3132) <= (layer0_outputs(5789)) or (layer0_outputs(824));
    outputs(3133) <= (layer0_outputs(10047)) xor (layer0_outputs(139));
    outputs(3134) <= layer0_outputs(8656);
    outputs(3135) <= (layer0_outputs(10203)) and not (layer0_outputs(4763));
    outputs(3136) <= not(layer0_outputs(9194));
    outputs(3137) <= not((layer0_outputs(7772)) xor (layer0_outputs(5555)));
    outputs(3138) <= not(layer0_outputs(10317)) or (layer0_outputs(12336));
    outputs(3139) <= (layer0_outputs(5466)) and (layer0_outputs(12732));
    outputs(3140) <= layer0_outputs(1300);
    outputs(3141) <= not(layer0_outputs(11926)) or (layer0_outputs(5805));
    outputs(3142) <= layer0_outputs(2537);
    outputs(3143) <= layer0_outputs(7188);
    outputs(3144) <= not(layer0_outputs(11066)) or (layer0_outputs(7317));
    outputs(3145) <= (layer0_outputs(5615)) xor (layer0_outputs(11268));
    outputs(3146) <= not((layer0_outputs(11381)) xor (layer0_outputs(8058)));
    outputs(3147) <= (layer0_outputs(5742)) and (layer0_outputs(7925));
    outputs(3148) <= layer0_outputs(10700);
    outputs(3149) <= not(layer0_outputs(8401));
    outputs(3150) <= not(layer0_outputs(3402));
    outputs(3151) <= (layer0_outputs(10803)) xor (layer0_outputs(5296));
    outputs(3152) <= not(layer0_outputs(12411)) or (layer0_outputs(2932));
    outputs(3153) <= layer0_outputs(6719);
    outputs(3154) <= not((layer0_outputs(11546)) or (layer0_outputs(12667)));
    outputs(3155) <= (layer0_outputs(7516)) xor (layer0_outputs(5061));
    outputs(3156) <= not(layer0_outputs(2838));
    outputs(3157) <= (layer0_outputs(9676)) xor (layer0_outputs(10671));
    outputs(3158) <= layer0_outputs(7539);
    outputs(3159) <= (layer0_outputs(6193)) xor (layer0_outputs(8230));
    outputs(3160) <= not(layer0_outputs(10646));
    outputs(3161) <= (layer0_outputs(8030)) xor (layer0_outputs(7082));
    outputs(3162) <= (layer0_outputs(2654)) or (layer0_outputs(6079));
    outputs(3163) <= layer0_outputs(8561);
    outputs(3164) <= (layer0_outputs(3319)) and (layer0_outputs(5464));
    outputs(3165) <= not(layer0_outputs(4330));
    outputs(3166) <= layer0_outputs(6782);
    outputs(3167) <= not(layer0_outputs(7743));
    outputs(3168) <= not(layer0_outputs(1023));
    outputs(3169) <= not(layer0_outputs(897));
    outputs(3170) <= not(layer0_outputs(6780));
    outputs(3171) <= not(layer0_outputs(6461));
    outputs(3172) <= layer0_outputs(7585);
    outputs(3173) <= not(layer0_outputs(7727));
    outputs(3174) <= not(layer0_outputs(1186));
    outputs(3175) <= not((layer0_outputs(8740)) xor (layer0_outputs(7631)));
    outputs(3176) <= (layer0_outputs(5346)) and (layer0_outputs(10690));
    outputs(3177) <= not(layer0_outputs(9723));
    outputs(3178) <= (layer0_outputs(5419)) and not (layer0_outputs(10178));
    outputs(3179) <= (layer0_outputs(9921)) and not (layer0_outputs(6783));
    outputs(3180) <= not(layer0_outputs(11359)) or (layer0_outputs(10913));
    outputs(3181) <= (layer0_outputs(5735)) xor (layer0_outputs(5894));
    outputs(3182) <= not(layer0_outputs(12041));
    outputs(3183) <= layer0_outputs(485);
    outputs(3184) <= (layer0_outputs(6156)) xor (layer0_outputs(11464));
    outputs(3185) <= (layer0_outputs(2840)) xor (layer0_outputs(4010));
    outputs(3186) <= layer0_outputs(10498);
    outputs(3187) <= not((layer0_outputs(627)) or (layer0_outputs(6681)));
    outputs(3188) <= (layer0_outputs(6768)) xor (layer0_outputs(10477));
    outputs(3189) <= layer0_outputs(6639);
    outputs(3190) <= (layer0_outputs(9817)) and not (layer0_outputs(4312));
    outputs(3191) <= not(layer0_outputs(10856));
    outputs(3192) <= layer0_outputs(3171);
    outputs(3193) <= (layer0_outputs(872)) and not (layer0_outputs(5518));
    outputs(3194) <= not(layer0_outputs(6088)) or (layer0_outputs(2876));
    outputs(3195) <= not(layer0_outputs(100));
    outputs(3196) <= layer0_outputs(5673);
    outputs(3197) <= layer0_outputs(11010);
    outputs(3198) <= not(layer0_outputs(9342)) or (layer0_outputs(9541));
    outputs(3199) <= (layer0_outputs(11634)) and (layer0_outputs(8500));
    outputs(3200) <= (layer0_outputs(4236)) and (layer0_outputs(1107));
    outputs(3201) <= not(layer0_outputs(3908));
    outputs(3202) <= (layer0_outputs(2748)) xor (layer0_outputs(7406));
    outputs(3203) <= not(layer0_outputs(7854));
    outputs(3204) <= (layer0_outputs(9052)) or (layer0_outputs(3466));
    outputs(3205) <= not(layer0_outputs(10854));
    outputs(3206) <= not((layer0_outputs(6896)) xor (layer0_outputs(5317)));
    outputs(3207) <= not(layer0_outputs(61));
    outputs(3208) <= (layer0_outputs(980)) xor (layer0_outputs(11185));
    outputs(3209) <= not((layer0_outputs(2219)) xor (layer0_outputs(7502)));
    outputs(3210) <= (layer0_outputs(5232)) xor (layer0_outputs(1975));
    outputs(3211) <= layer0_outputs(7503);
    outputs(3212) <= not(layer0_outputs(9051)) or (layer0_outputs(6207));
    outputs(3213) <= (layer0_outputs(90)) and not (layer0_outputs(11447));
    outputs(3214) <= not(layer0_outputs(10962));
    outputs(3215) <= not(layer0_outputs(9706));
    outputs(3216) <= (layer0_outputs(6347)) xor (layer0_outputs(679));
    outputs(3217) <= (layer0_outputs(330)) or (layer0_outputs(2804));
    outputs(3218) <= not(layer0_outputs(929));
    outputs(3219) <= not((layer0_outputs(5141)) and (layer0_outputs(12570)));
    outputs(3220) <= not((layer0_outputs(5458)) and (layer0_outputs(11985)));
    outputs(3221) <= not(layer0_outputs(1816));
    outputs(3222) <= layer0_outputs(4125);
    outputs(3223) <= (layer0_outputs(12483)) and not (layer0_outputs(7742));
    outputs(3224) <= not((layer0_outputs(11050)) xor (layer0_outputs(8970)));
    outputs(3225) <= not((layer0_outputs(7974)) and (layer0_outputs(1902)));
    outputs(3226) <= layer0_outputs(4420);
    outputs(3227) <= layer0_outputs(5636);
    outputs(3228) <= (layer0_outputs(4548)) xor (layer0_outputs(3861));
    outputs(3229) <= layer0_outputs(5769);
    outputs(3230) <= layer0_outputs(50);
    outputs(3231) <= layer0_outputs(353);
    outputs(3232) <= (layer0_outputs(1753)) xor (layer0_outputs(2361));
    outputs(3233) <= not((layer0_outputs(1011)) xor (layer0_outputs(3465)));
    outputs(3234) <= not((layer0_outputs(108)) xor (layer0_outputs(3598)));
    outputs(3235) <= layer0_outputs(1947);
    outputs(3236) <= (layer0_outputs(4222)) and not (layer0_outputs(10027));
    outputs(3237) <= not(layer0_outputs(10513)) or (layer0_outputs(3382));
    outputs(3238) <= not(layer0_outputs(1414));
    outputs(3239) <= not((layer0_outputs(12023)) or (layer0_outputs(131)));
    outputs(3240) <= layer0_outputs(6017);
    outputs(3241) <= (layer0_outputs(11481)) xor (layer0_outputs(94));
    outputs(3242) <= not(layer0_outputs(705));
    outputs(3243) <= (layer0_outputs(6613)) xor (layer0_outputs(2363));
    outputs(3244) <= not(layer0_outputs(8963));
    outputs(3245) <= (layer0_outputs(11518)) and not (layer0_outputs(10489));
    outputs(3246) <= (layer0_outputs(3488)) and not (layer0_outputs(5033));
    outputs(3247) <= (layer0_outputs(11849)) or (layer0_outputs(11701));
    outputs(3248) <= layer0_outputs(4194);
    outputs(3249) <= layer0_outputs(10341);
    outputs(3250) <= not((layer0_outputs(1566)) xor (layer0_outputs(7552)));
    outputs(3251) <= not(layer0_outputs(8279)) or (layer0_outputs(7177));
    outputs(3252) <= (layer0_outputs(9809)) or (layer0_outputs(9575));
    outputs(3253) <= (layer0_outputs(10861)) xor (layer0_outputs(8549));
    outputs(3254) <= (layer0_outputs(11477)) xor (layer0_outputs(9487));
    outputs(3255) <= layer0_outputs(6789);
    outputs(3256) <= layer0_outputs(2313);
    outputs(3257) <= (layer0_outputs(10036)) or (layer0_outputs(10436));
    outputs(3258) <= not((layer0_outputs(10458)) xor (layer0_outputs(10550)));
    outputs(3259) <= not(layer0_outputs(11466)) or (layer0_outputs(11112));
    outputs(3260) <= (layer0_outputs(7129)) or (layer0_outputs(12415));
    outputs(3261) <= not(layer0_outputs(2666));
    outputs(3262) <= not((layer0_outputs(12622)) xor (layer0_outputs(599)));
    outputs(3263) <= not(layer0_outputs(5690));
    outputs(3264) <= not(layer0_outputs(10231));
    outputs(3265) <= not((layer0_outputs(546)) xor (layer0_outputs(11423)));
    outputs(3266) <= not((layer0_outputs(1938)) and (layer0_outputs(2380)));
    outputs(3267) <= (layer0_outputs(4635)) or (layer0_outputs(5681));
    outputs(3268) <= (layer0_outputs(12274)) and (layer0_outputs(6817));
    outputs(3269) <= not(layer0_outputs(7461));
    outputs(3270) <= (layer0_outputs(3100)) and not (layer0_outputs(1876));
    outputs(3271) <= (layer0_outputs(7914)) and not (layer0_outputs(5229));
    outputs(3272) <= layer0_outputs(7678);
    outputs(3273) <= (layer0_outputs(7451)) xor (layer0_outputs(5921));
    outputs(3274) <= not(layer0_outputs(11181));
    outputs(3275) <= (layer0_outputs(4801)) or (layer0_outputs(5790));
    outputs(3276) <= (layer0_outputs(5524)) xor (layer0_outputs(5224));
    outputs(3277) <= layer0_outputs(9809);
    outputs(3278) <= (layer0_outputs(6899)) or (layer0_outputs(9685));
    outputs(3279) <= (layer0_outputs(6955)) xor (layer0_outputs(9401));
    outputs(3280) <= not((layer0_outputs(9441)) xor (layer0_outputs(1783)));
    outputs(3281) <= not(layer0_outputs(10522)) or (layer0_outputs(9843));
    outputs(3282) <= not(layer0_outputs(12709));
    outputs(3283) <= (layer0_outputs(5657)) and not (layer0_outputs(4467));
    outputs(3284) <= not(layer0_outputs(10200));
    outputs(3285) <= not(layer0_outputs(1590)) or (layer0_outputs(10098));
    outputs(3286) <= not(layer0_outputs(4850));
    outputs(3287) <= not(layer0_outputs(3555));
    outputs(3288) <= layer0_outputs(1837);
    outputs(3289) <= not(layer0_outputs(5757));
    outputs(3290) <= (layer0_outputs(11440)) and not (layer0_outputs(10802));
    outputs(3291) <= (layer0_outputs(1236)) xor (layer0_outputs(9348));
    outputs(3292) <= not(layer0_outputs(2875)) or (layer0_outputs(8728));
    outputs(3293) <= (layer0_outputs(1807)) or (layer0_outputs(3753));
    outputs(3294) <= (layer0_outputs(9651)) or (layer0_outputs(5923));
    outputs(3295) <= (layer0_outputs(2933)) xor (layer0_outputs(6644));
    outputs(3296) <= (layer0_outputs(8888)) xor (layer0_outputs(11708));
    outputs(3297) <= not(layer0_outputs(9933)) or (layer0_outputs(11870));
    outputs(3298) <= not((layer0_outputs(2639)) xor (layer0_outputs(6744)));
    outputs(3299) <= (layer0_outputs(8390)) and not (layer0_outputs(736));
    outputs(3300) <= (layer0_outputs(1565)) xor (layer0_outputs(4822));
    outputs(3301) <= (layer0_outputs(7363)) and not (layer0_outputs(4748));
    outputs(3302) <= not(layer0_outputs(1034));
    outputs(3303) <= layer0_outputs(5868);
    outputs(3304) <= not(layer0_outputs(8214));
    outputs(3305) <= not((layer0_outputs(1032)) xor (layer0_outputs(11330)));
    outputs(3306) <= layer0_outputs(9734);
    outputs(3307) <= not((layer0_outputs(2599)) or (layer0_outputs(1744)));
    outputs(3308) <= not(layer0_outputs(5707));
    outputs(3309) <= (layer0_outputs(2191)) or (layer0_outputs(6524));
    outputs(3310) <= layer0_outputs(3241);
    outputs(3311) <= not((layer0_outputs(6331)) xor (layer0_outputs(11909)));
    outputs(3312) <= layer0_outputs(2249);
    outputs(3313) <= not((layer0_outputs(7191)) xor (layer0_outputs(1694)));
    outputs(3314) <= (layer0_outputs(6131)) xor (layer0_outputs(5983));
    outputs(3315) <= not(layer0_outputs(2221));
    outputs(3316) <= layer0_outputs(9750);
    outputs(3317) <= (layer0_outputs(8143)) and (layer0_outputs(4159));
    outputs(3318) <= not((layer0_outputs(11678)) and (layer0_outputs(9429)));
    outputs(3319) <= not((layer0_outputs(5651)) and (layer0_outputs(7089)));
    outputs(3320) <= layer0_outputs(495);
    outputs(3321) <= (layer0_outputs(8013)) or (layer0_outputs(9338));
    outputs(3322) <= not((layer0_outputs(400)) and (layer0_outputs(4039)));
    outputs(3323) <= (layer0_outputs(5085)) and (layer0_outputs(11236));
    outputs(3324) <= not((layer0_outputs(2042)) xor (layer0_outputs(816)));
    outputs(3325) <= layer0_outputs(9392);
    outputs(3326) <= layer0_outputs(2990);
    outputs(3327) <= not(layer0_outputs(3597));
    outputs(3328) <= layer0_outputs(1820);
    outputs(3329) <= layer0_outputs(8852);
    outputs(3330) <= (layer0_outputs(4517)) xor (layer0_outputs(11809));
    outputs(3331) <= layer0_outputs(2190);
    outputs(3332) <= not((layer0_outputs(7463)) xor (layer0_outputs(208)));
    outputs(3333) <= not((layer0_outputs(10853)) and (layer0_outputs(5977)));
    outputs(3334) <= (layer0_outputs(2244)) xor (layer0_outputs(4365));
    outputs(3335) <= (layer0_outputs(5215)) xor (layer0_outputs(5586));
    outputs(3336) <= layer0_outputs(6739);
    outputs(3337) <= layer0_outputs(12149);
    outputs(3338) <= not(layer0_outputs(836)) or (layer0_outputs(2490));
    outputs(3339) <= not(layer0_outputs(3530));
    outputs(3340) <= (layer0_outputs(786)) xor (layer0_outputs(298));
    outputs(3341) <= (layer0_outputs(11577)) xor (layer0_outputs(2358));
    outputs(3342) <= not((layer0_outputs(2638)) xor (layer0_outputs(5606)));
    outputs(3343) <= not((layer0_outputs(8493)) and (layer0_outputs(1479)));
    outputs(3344) <= not((layer0_outputs(3424)) xor (layer0_outputs(8644)));
    outputs(3345) <= not((layer0_outputs(11497)) and (layer0_outputs(11407)));
    outputs(3346) <= not((layer0_outputs(2568)) xor (layer0_outputs(6307)));
    outputs(3347) <= (layer0_outputs(4953)) xor (layer0_outputs(2867));
    outputs(3348) <= layer0_outputs(2833);
    outputs(3349) <= (layer0_outputs(7621)) xor (layer0_outputs(379));
    outputs(3350) <= (layer0_outputs(10348)) xor (layer0_outputs(5526));
    outputs(3351) <= (layer0_outputs(10426)) or (layer0_outputs(9373));
    outputs(3352) <= '1';
    outputs(3353) <= layer0_outputs(4084);
    outputs(3354) <= not(layer0_outputs(12761));
    outputs(3355) <= not((layer0_outputs(7740)) and (layer0_outputs(338)));
    outputs(3356) <= layer0_outputs(9993);
    outputs(3357) <= not(layer0_outputs(4101)) or (layer0_outputs(7169));
    outputs(3358) <= not((layer0_outputs(12636)) and (layer0_outputs(1326)));
    outputs(3359) <= (layer0_outputs(492)) and (layer0_outputs(8746));
    outputs(3360) <= (layer0_outputs(12346)) xor (layer0_outputs(3097));
    outputs(3361) <= (layer0_outputs(11198)) and not (layer0_outputs(5054));
    outputs(3362) <= layer0_outputs(9019);
    outputs(3363) <= (layer0_outputs(10120)) xor (layer0_outputs(7879));
    outputs(3364) <= not(layer0_outputs(8356)) or (layer0_outputs(10340));
    outputs(3365) <= not((layer0_outputs(3727)) xor (layer0_outputs(5719)));
    outputs(3366) <= (layer0_outputs(11719)) or (layer0_outputs(9011));
    outputs(3367) <= not(layer0_outputs(6887));
    outputs(3368) <= layer0_outputs(4940);
    outputs(3369) <= not(layer0_outputs(3039));
    outputs(3370) <= layer0_outputs(9956);
    outputs(3371) <= not((layer0_outputs(9042)) and (layer0_outputs(3463)));
    outputs(3372) <= not(layer0_outputs(4415));
    outputs(3373) <= not((layer0_outputs(3726)) xor (layer0_outputs(104)));
    outputs(3374) <= not(layer0_outputs(12368)) or (layer0_outputs(12183));
    outputs(3375) <= (layer0_outputs(4975)) xor (layer0_outputs(6395));
    outputs(3376) <= layer0_outputs(1985);
    outputs(3377) <= (layer0_outputs(10679)) xor (layer0_outputs(4823));
    outputs(3378) <= not(layer0_outputs(1651)) or (layer0_outputs(8911));
    outputs(3379) <= (layer0_outputs(6264)) or (layer0_outputs(168));
    outputs(3380) <= layer0_outputs(4434);
    outputs(3381) <= layer0_outputs(493);
    outputs(3382) <= not((layer0_outputs(7730)) xor (layer0_outputs(3162)));
    outputs(3383) <= not((layer0_outputs(6964)) xor (layer0_outputs(457)));
    outputs(3384) <= layer0_outputs(3168);
    outputs(3385) <= (layer0_outputs(12568)) and not (layer0_outputs(7400));
    outputs(3386) <= not(layer0_outputs(2152));
    outputs(3387) <= layer0_outputs(5081);
    outputs(3388) <= not((layer0_outputs(2345)) or (layer0_outputs(7399)));
    outputs(3389) <= not(layer0_outputs(5527));
    outputs(3390) <= (layer0_outputs(211)) and not (layer0_outputs(5055));
    outputs(3391) <= layer0_outputs(2975);
    outputs(3392) <= not((layer0_outputs(8145)) and (layer0_outputs(12693)));
    outputs(3393) <= layer0_outputs(12231);
    outputs(3394) <= not(layer0_outputs(1089));
    outputs(3395) <= layer0_outputs(9329);
    outputs(3396) <= (layer0_outputs(10135)) and (layer0_outputs(10969));
    outputs(3397) <= not(layer0_outputs(9141)) or (layer0_outputs(3742));
    outputs(3398) <= not((layer0_outputs(3832)) and (layer0_outputs(1863)));
    outputs(3399) <= not(layer0_outputs(2361));
    outputs(3400) <= not(layer0_outputs(3680));
    outputs(3401) <= (layer0_outputs(11238)) xor (layer0_outputs(10277));
    outputs(3402) <= not((layer0_outputs(5772)) xor (layer0_outputs(1887)));
    outputs(3403) <= not((layer0_outputs(8584)) and (layer0_outputs(488)));
    outputs(3404) <= not(layer0_outputs(1697));
    outputs(3405) <= not(layer0_outputs(4549));
    outputs(3406) <= (layer0_outputs(2194)) xor (layer0_outputs(10773));
    outputs(3407) <= not((layer0_outputs(6373)) xor (layer0_outputs(7987)));
    outputs(3408) <= not((layer0_outputs(9522)) xor (layer0_outputs(8870)));
    outputs(3409) <= layer0_outputs(3396);
    outputs(3410) <= (layer0_outputs(9067)) xor (layer0_outputs(10363));
    outputs(3411) <= not((layer0_outputs(3886)) and (layer0_outputs(2095)));
    outputs(3412) <= not((layer0_outputs(1753)) xor (layer0_outputs(3143)));
    outputs(3413) <= (layer0_outputs(1128)) and (layer0_outputs(302));
    outputs(3414) <= (layer0_outputs(8500)) xor (layer0_outputs(2046));
    outputs(3415) <= (layer0_outputs(4095)) and not (layer0_outputs(9040));
    outputs(3416) <= layer0_outputs(12399);
    outputs(3417) <= not(layer0_outputs(3568)) or (layer0_outputs(6650));
    outputs(3418) <= not((layer0_outputs(6025)) and (layer0_outputs(11162)));
    outputs(3419) <= not(layer0_outputs(4982)) or (layer0_outputs(3414));
    outputs(3420) <= not(layer0_outputs(7660));
    outputs(3421) <= '1';
    outputs(3422) <= not((layer0_outputs(7077)) and (layer0_outputs(4220)));
    outputs(3423) <= (layer0_outputs(2073)) or (layer0_outputs(754));
    outputs(3424) <= layer0_outputs(2826);
    outputs(3425) <= not((layer0_outputs(5247)) xor (layer0_outputs(2959)));
    outputs(3426) <= (layer0_outputs(6529)) xor (layer0_outputs(10276));
    outputs(3427) <= not((layer0_outputs(9751)) xor (layer0_outputs(5054)));
    outputs(3428) <= layer0_outputs(6863);
    outputs(3429) <= layer0_outputs(4789);
    outputs(3430) <= (layer0_outputs(7352)) and not (layer0_outputs(10469));
    outputs(3431) <= not(layer0_outputs(10883)) or (layer0_outputs(9641));
    outputs(3432) <= layer0_outputs(1435);
    outputs(3433) <= layer0_outputs(4878);
    outputs(3434) <= not(layer0_outputs(1439)) or (layer0_outputs(680));
    outputs(3435) <= not(layer0_outputs(7435));
    outputs(3436) <= layer0_outputs(11828);
    outputs(3437) <= not(layer0_outputs(8477));
    outputs(3438) <= not((layer0_outputs(10882)) or (layer0_outputs(8072)));
    outputs(3439) <= not(layer0_outputs(9635)) or (layer0_outputs(8035));
    outputs(3440) <= not((layer0_outputs(7887)) xor (layer0_outputs(9763)));
    outputs(3441) <= (layer0_outputs(6707)) and (layer0_outputs(7046));
    outputs(3442) <= (layer0_outputs(3218)) or (layer0_outputs(7149));
    outputs(3443) <= (layer0_outputs(10855)) and (layer0_outputs(1728));
    outputs(3444) <= not((layer0_outputs(7472)) xor (layer0_outputs(7304)));
    outputs(3445) <= layer0_outputs(1289);
    outputs(3446) <= (layer0_outputs(3776)) and (layer0_outputs(10043));
    outputs(3447) <= layer0_outputs(5184);
    outputs(3448) <= not((layer0_outputs(2842)) xor (layer0_outputs(380)));
    outputs(3449) <= not(layer0_outputs(1652)) or (layer0_outputs(4426));
    outputs(3450) <= not(layer0_outputs(1307)) or (layer0_outputs(11482));
    outputs(3451) <= not(layer0_outputs(1031));
    outputs(3452) <= not(layer0_outputs(11245));
    outputs(3453) <= not(layer0_outputs(1497));
    outputs(3454) <= not(layer0_outputs(4686)) or (layer0_outputs(433));
    outputs(3455) <= not((layer0_outputs(5736)) xor (layer0_outputs(423)));
    outputs(3456) <= not(layer0_outputs(11093));
    outputs(3457) <= not((layer0_outputs(9926)) or (layer0_outputs(5362)));
    outputs(3458) <= (layer0_outputs(8940)) and (layer0_outputs(5152));
    outputs(3459) <= layer0_outputs(12657);
    outputs(3460) <= not((layer0_outputs(2964)) and (layer0_outputs(6380)));
    outputs(3461) <= not(layer0_outputs(12160));
    outputs(3462) <= layer0_outputs(3670);
    outputs(3463) <= not((layer0_outputs(4969)) xor (layer0_outputs(5709)));
    outputs(3464) <= not(layer0_outputs(825));
    outputs(3465) <= (layer0_outputs(10612)) or (layer0_outputs(3304));
    outputs(3466) <= layer0_outputs(6032);
    outputs(3467) <= (layer0_outputs(4177)) xor (layer0_outputs(11891));
    outputs(3468) <= not((layer0_outputs(1598)) and (layer0_outputs(487)));
    outputs(3469) <= (layer0_outputs(1345)) xor (layer0_outputs(2329));
    outputs(3470) <= not((layer0_outputs(12171)) and (layer0_outputs(4213)));
    outputs(3471) <= not((layer0_outputs(5937)) and (layer0_outputs(7071)));
    outputs(3472) <= not((layer0_outputs(8618)) xor (layer0_outputs(6361)));
    outputs(3473) <= layer0_outputs(5987);
    outputs(3474) <= layer0_outputs(3174);
    outputs(3475) <= (layer0_outputs(465)) xor (layer0_outputs(2051));
    outputs(3476) <= not(layer0_outputs(8763));
    outputs(3477) <= (layer0_outputs(12760)) xor (layer0_outputs(8936));
    outputs(3478) <= layer0_outputs(1688);
    outputs(3479) <= layer0_outputs(8796);
    outputs(3480) <= layer0_outputs(1431);
    outputs(3481) <= not((layer0_outputs(7021)) xor (layer0_outputs(9614)));
    outputs(3482) <= layer0_outputs(11838);
    outputs(3483) <= (layer0_outputs(4756)) xor (layer0_outputs(11453));
    outputs(3484) <= layer0_outputs(3080);
    outputs(3485) <= (layer0_outputs(5688)) xor (layer0_outputs(5646));
    outputs(3486) <= layer0_outputs(684);
    outputs(3487) <= layer0_outputs(6740);
    outputs(3488) <= not((layer0_outputs(6081)) and (layer0_outputs(4405)));
    outputs(3489) <= not((layer0_outputs(9149)) and (layer0_outputs(1229)));
    outputs(3490) <= layer0_outputs(12539);
    outputs(3491) <= not((layer0_outputs(1666)) or (layer0_outputs(6257)));
    outputs(3492) <= not((layer0_outputs(9763)) and (layer0_outputs(10338)));
    outputs(3493) <= (layer0_outputs(3550)) xor (layer0_outputs(12264));
    outputs(3494) <= layer0_outputs(6726);
    outputs(3495) <= not(layer0_outputs(10580)) or (layer0_outputs(7157));
    outputs(3496) <= not((layer0_outputs(10110)) and (layer0_outputs(12411)));
    outputs(3497) <= not((layer0_outputs(2285)) and (layer0_outputs(8974)));
    outputs(3498) <= (layer0_outputs(9120)) xor (layer0_outputs(7074));
    outputs(3499) <= layer0_outputs(11227);
    outputs(3500) <= not(layer0_outputs(6119)) or (layer0_outputs(9143));
    outputs(3501) <= layer0_outputs(6544);
    outputs(3502) <= (layer0_outputs(8609)) xor (layer0_outputs(2265));
    outputs(3503) <= not(layer0_outputs(12111));
    outputs(3504) <= (layer0_outputs(4131)) xor (layer0_outputs(10629));
    outputs(3505) <= not(layer0_outputs(9782)) or (layer0_outputs(7979));
    outputs(3506) <= not((layer0_outputs(5145)) xor (layer0_outputs(6081)));
    outputs(3507) <= layer0_outputs(1678);
    outputs(3508) <= (layer0_outputs(12093)) and not (layer0_outputs(6759));
    outputs(3509) <= not((layer0_outputs(2621)) xor (layer0_outputs(11647)));
    outputs(3510) <= not((layer0_outputs(5021)) xor (layer0_outputs(9211)));
    outputs(3511) <= (layer0_outputs(11446)) and not (layer0_outputs(12322));
    outputs(3512) <= (layer0_outputs(2094)) xor (layer0_outputs(6594));
    outputs(3513) <= layer0_outputs(3433);
    outputs(3514) <= not((layer0_outputs(10170)) xor (layer0_outputs(4374)));
    outputs(3515) <= not((layer0_outputs(5540)) xor (layer0_outputs(3518)));
    outputs(3516) <= not((layer0_outputs(5226)) xor (layer0_outputs(11046)));
    outputs(3517) <= not((layer0_outputs(175)) and (layer0_outputs(10894)));
    outputs(3518) <= layer0_outputs(3765);
    outputs(3519) <= (layer0_outputs(4144)) and (layer0_outputs(7758));
    outputs(3520) <= (layer0_outputs(6599)) or (layer0_outputs(8310));
    outputs(3521) <= (layer0_outputs(5044)) and not (layer0_outputs(5680));
    outputs(3522) <= not(layer0_outputs(10569));
    outputs(3523) <= (layer0_outputs(2726)) xor (layer0_outputs(11656));
    outputs(3524) <= layer0_outputs(11417);
    outputs(3525) <= (layer0_outputs(11900)) xor (layer0_outputs(2600));
    outputs(3526) <= not(layer0_outputs(12608));
    outputs(3527) <= not(layer0_outputs(6277)) or (layer0_outputs(1533));
    outputs(3528) <= layer0_outputs(3149);
    outputs(3529) <= (layer0_outputs(7137)) and not (layer0_outputs(3735));
    outputs(3530) <= (layer0_outputs(10925)) xor (layer0_outputs(6720));
    outputs(3531) <= not(layer0_outputs(132));
    outputs(3532) <= not(layer0_outputs(11988));
    outputs(3533) <= not((layer0_outputs(2116)) xor (layer0_outputs(3400)));
    outputs(3534) <= layer0_outputs(11588);
    outputs(3535) <= not((layer0_outputs(5926)) xor (layer0_outputs(12214)));
    outputs(3536) <= (layer0_outputs(3265)) or (layer0_outputs(4830));
    outputs(3537) <= not((layer0_outputs(7888)) xor (layer0_outputs(12528)));
    outputs(3538) <= not(layer0_outputs(1406)) or (layer0_outputs(9757));
    outputs(3539) <= not((layer0_outputs(3528)) and (layer0_outputs(6666)));
    outputs(3540) <= (layer0_outputs(10707)) xor (layer0_outputs(439));
    outputs(3541) <= not(layer0_outputs(2132));
    outputs(3542) <= (layer0_outputs(8567)) and (layer0_outputs(2094));
    outputs(3543) <= layer0_outputs(6935);
    outputs(3544) <= (layer0_outputs(9386)) and not (layer0_outputs(5768));
    outputs(3545) <= not(layer0_outputs(4868)) or (layer0_outputs(12092));
    outputs(3546) <= (layer0_outputs(11178)) and not (layer0_outputs(7786));
    outputs(3547) <= (layer0_outputs(5561)) xor (layer0_outputs(5938));
    outputs(3548) <= not(layer0_outputs(11680)) or (layer0_outputs(1071));
    outputs(3549) <= not((layer0_outputs(11674)) xor (layer0_outputs(1916)));
    outputs(3550) <= not(layer0_outputs(11562));
    outputs(3551) <= (layer0_outputs(11836)) and (layer0_outputs(12394));
    outputs(3552) <= not((layer0_outputs(7212)) xor (layer0_outputs(7773)));
    outputs(3553) <= (layer0_outputs(5340)) or (layer0_outputs(3662));
    outputs(3554) <= not(layer0_outputs(12720)) or (layer0_outputs(2038));
    outputs(3555) <= layer0_outputs(8005);
    outputs(3556) <= layer0_outputs(10377);
    outputs(3557) <= (layer0_outputs(9256)) or (layer0_outputs(3524));
    outputs(3558) <= not((layer0_outputs(447)) xor (layer0_outputs(4197)));
    outputs(3559) <= not(layer0_outputs(1028)) or (layer0_outputs(9037));
    outputs(3560) <= not(layer0_outputs(9245)) or (layer0_outputs(2710));
    outputs(3561) <= not(layer0_outputs(10926));
    outputs(3562) <= (layer0_outputs(10083)) xor (layer0_outputs(1130));
    outputs(3563) <= (layer0_outputs(9074)) xor (layer0_outputs(8307));
    outputs(3564) <= layer0_outputs(10253);
    outputs(3565) <= not(layer0_outputs(1671));
    outputs(3566) <= (layer0_outputs(2752)) or (layer0_outputs(3044));
    outputs(3567) <= layer0_outputs(10241);
    outputs(3568) <= (layer0_outputs(5095)) xor (layer0_outputs(8326));
    outputs(3569) <= layer0_outputs(4361);
    outputs(3570) <= not((layer0_outputs(6463)) xor (layer0_outputs(4803)));
    outputs(3571) <= not(layer0_outputs(1162)) or (layer0_outputs(7513));
    outputs(3572) <= not((layer0_outputs(11928)) xor (layer0_outputs(4342)));
    outputs(3573) <= not((layer0_outputs(488)) xor (layer0_outputs(4511)));
    outputs(3574) <= not(layer0_outputs(3325));
    outputs(3575) <= not((layer0_outputs(5109)) or (layer0_outputs(7622)));
    outputs(3576) <= (layer0_outputs(6594)) xor (layer0_outputs(563));
    outputs(3577) <= not((layer0_outputs(395)) xor (layer0_outputs(3632)));
    outputs(3578) <= not(layer0_outputs(7307));
    outputs(3579) <= (layer0_outputs(1346)) or (layer0_outputs(4287));
    outputs(3580) <= (layer0_outputs(6737)) xor (layer0_outputs(7816));
    outputs(3581) <= not(layer0_outputs(12066));
    outputs(3582) <= (layer0_outputs(9769)) xor (layer0_outputs(2030));
    outputs(3583) <= (layer0_outputs(2022)) and not (layer0_outputs(9824));
    outputs(3584) <= (layer0_outputs(4385)) xor (layer0_outputs(922));
    outputs(3585) <= layer0_outputs(10313);
    outputs(3586) <= not(layer0_outputs(8024));
    outputs(3587) <= not((layer0_outputs(8220)) or (layer0_outputs(6299)));
    outputs(3588) <= layer0_outputs(6020);
    outputs(3589) <= not(layer0_outputs(4580));
    outputs(3590) <= not((layer0_outputs(7451)) xor (layer0_outputs(5345)));
    outputs(3591) <= layer0_outputs(7787);
    outputs(3592) <= (layer0_outputs(6999)) xor (layer0_outputs(7337));
    outputs(3593) <= not((layer0_outputs(7371)) xor (layer0_outputs(6575)));
    outputs(3594) <= (layer0_outputs(34)) xor (layer0_outputs(11992));
    outputs(3595) <= not(layer0_outputs(11790));
    outputs(3596) <= (layer0_outputs(3927)) xor (layer0_outputs(6423));
    outputs(3597) <= not((layer0_outputs(5155)) xor (layer0_outputs(11713)));
    outputs(3598) <= (layer0_outputs(9778)) xor (layer0_outputs(9341));
    outputs(3599) <= not(layer0_outputs(6187));
    outputs(3600) <= layer0_outputs(7649);
    outputs(3601) <= layer0_outputs(2310);
    outputs(3602) <= (layer0_outputs(9575)) and not (layer0_outputs(8535));
    outputs(3603) <= not(layer0_outputs(4799)) or (layer0_outputs(2137));
    outputs(3604) <= not(layer0_outputs(7998));
    outputs(3605) <= not((layer0_outputs(5328)) xor (layer0_outputs(718)));
    outputs(3606) <= (layer0_outputs(9421)) xor (layer0_outputs(8475));
    outputs(3607) <= (layer0_outputs(1124)) xor (layer0_outputs(4956));
    outputs(3608) <= not((layer0_outputs(3964)) or (layer0_outputs(5129)));
    outputs(3609) <= layer0_outputs(12409);
    outputs(3610) <= not(layer0_outputs(11163)) or (layer0_outputs(3151));
    outputs(3611) <= not(layer0_outputs(639)) or (layer0_outputs(686));
    outputs(3612) <= not(layer0_outputs(9024));
    outputs(3613) <= layer0_outputs(7694);
    outputs(3614) <= not(layer0_outputs(6428));
    outputs(3615) <= layer0_outputs(5086);
    outputs(3616) <= layer0_outputs(6867);
    outputs(3617) <= layer0_outputs(846);
    outputs(3618) <= not(layer0_outputs(10131)) or (layer0_outputs(1247));
    outputs(3619) <= (layer0_outputs(12491)) or (layer0_outputs(8224));
    outputs(3620) <= not(layer0_outputs(5374));
    outputs(3621) <= not(layer0_outputs(7941));
    outputs(3622) <= (layer0_outputs(11191)) xor (layer0_outputs(2011));
    outputs(3623) <= not(layer0_outputs(8361)) or (layer0_outputs(5959));
    outputs(3624) <= (layer0_outputs(12010)) xor (layer0_outputs(3873));
    outputs(3625) <= (layer0_outputs(5824)) xor (layer0_outputs(4552));
    outputs(3626) <= not((layer0_outputs(3416)) xor (layer0_outputs(9851)));
    outputs(3627) <= (layer0_outputs(10252)) and (layer0_outputs(1785));
    outputs(3628) <= not((layer0_outputs(2863)) and (layer0_outputs(5079)));
    outputs(3629) <= not(layer0_outputs(225)) or (layer0_outputs(12369));
    outputs(3630) <= layer0_outputs(1265);
    outputs(3631) <= not(layer0_outputs(6329));
    outputs(3632) <= not(layer0_outputs(1905)) or (layer0_outputs(7951));
    outputs(3633) <= not(layer0_outputs(12436));
    outputs(3634) <= not(layer0_outputs(12585));
    outputs(3635) <= (layer0_outputs(11623)) xor (layer0_outputs(5457));
    outputs(3636) <= (layer0_outputs(10973)) and (layer0_outputs(2473));
    outputs(3637) <= not((layer0_outputs(2341)) or (layer0_outputs(11216)));
    outputs(3638) <= (layer0_outputs(296)) xor (layer0_outputs(12137));
    outputs(3639) <= not(layer0_outputs(301));
    outputs(3640) <= not((layer0_outputs(8673)) xor (layer0_outputs(3941)));
    outputs(3641) <= (layer0_outputs(7101)) xor (layer0_outputs(4395));
    outputs(3642) <= not(layer0_outputs(1400));
    outputs(3643) <= not(layer0_outputs(4518));
    outputs(3644) <= (layer0_outputs(10431)) or (layer0_outputs(9098));
    outputs(3645) <= not(layer0_outputs(858)) or (layer0_outputs(5967));
    outputs(3646) <= not(layer0_outputs(7959));
    outputs(3647) <= not(layer0_outputs(508));
    outputs(3648) <= (layer0_outputs(5740)) and not (layer0_outputs(3363));
    outputs(3649) <= (layer0_outputs(9162)) and not (layer0_outputs(285));
    outputs(3650) <= (layer0_outputs(8424)) xor (layer0_outputs(11639));
    outputs(3651) <= not(layer0_outputs(10673));
    outputs(3652) <= not((layer0_outputs(8171)) and (layer0_outputs(7013)));
    outputs(3653) <= layer0_outputs(373);
    outputs(3654) <= not(layer0_outputs(6566));
    outputs(3655) <= not((layer0_outputs(9814)) and (layer0_outputs(3747)));
    outputs(3656) <= not((layer0_outputs(8073)) xor (layer0_outputs(6147)));
    outputs(3657) <= not(layer0_outputs(6160));
    outputs(3658) <= (layer0_outputs(1397)) xor (layer0_outputs(329));
    outputs(3659) <= layer0_outputs(2724);
    outputs(3660) <= (layer0_outputs(6045)) and (layer0_outputs(12517));
    outputs(3661) <= (layer0_outputs(12021)) or (layer0_outputs(4993));
    outputs(3662) <= not(layer0_outputs(6206));
    outputs(3663) <= not(layer0_outputs(11079)) or (layer0_outputs(686));
    outputs(3664) <= (layer0_outputs(9674)) and (layer0_outputs(3285));
    outputs(3665) <= not((layer0_outputs(12400)) and (layer0_outputs(4861)));
    outputs(3666) <= not(layer0_outputs(10910)) or (layer0_outputs(526));
    outputs(3667) <= not(layer0_outputs(10568));
    outputs(3668) <= not(layer0_outputs(3184)) or (layer0_outputs(280));
    outputs(3669) <= not(layer0_outputs(10352));
    outputs(3670) <= layer0_outputs(5881);
    outputs(3671) <= not(layer0_outputs(11640));
    outputs(3672) <= not((layer0_outputs(7900)) and (layer0_outputs(8217)));
    outputs(3673) <= not(layer0_outputs(2847)) or (layer0_outputs(10955));
    outputs(3674) <= not(layer0_outputs(180)) or (layer0_outputs(6301));
    outputs(3675) <= not((layer0_outputs(7707)) and (layer0_outputs(498)));
    outputs(3676) <= not(layer0_outputs(6105)) or (layer0_outputs(2707));
    outputs(3677) <= layer0_outputs(3852);
    outputs(3678) <= not(layer0_outputs(11801));
    outputs(3679) <= not((layer0_outputs(669)) xor (layer0_outputs(9443)));
    outputs(3680) <= not((layer0_outputs(169)) and (layer0_outputs(4863)));
    outputs(3681) <= not((layer0_outputs(9452)) xor (layer0_outputs(9525)));
    outputs(3682) <= (layer0_outputs(11140)) and not (layer0_outputs(2457));
    outputs(3683) <= not((layer0_outputs(5021)) xor (layer0_outputs(5326)));
    outputs(3684) <= not((layer0_outputs(1726)) xor (layer0_outputs(6988)));
    outputs(3685) <= not((layer0_outputs(5810)) xor (layer0_outputs(2836)));
    outputs(3686) <= not(layer0_outputs(12017));
    outputs(3687) <= not(layer0_outputs(6942));
    outputs(3688) <= not(layer0_outputs(4729));
    outputs(3689) <= not((layer0_outputs(12556)) xor (layer0_outputs(1000)));
    outputs(3690) <= (layer0_outputs(2777)) xor (layer0_outputs(4987));
    outputs(3691) <= not(layer0_outputs(11018)) or (layer0_outputs(4789));
    outputs(3692) <= (layer0_outputs(7778)) and (layer0_outputs(9349));
    outputs(3693) <= not((layer0_outputs(11162)) and (layer0_outputs(10591)));
    outputs(3694) <= not((layer0_outputs(9768)) xor (layer0_outputs(4707)));
    outputs(3695) <= not(layer0_outputs(12473));
    outputs(3696) <= (layer0_outputs(6250)) and not (layer0_outputs(8276));
    outputs(3697) <= not((layer0_outputs(1770)) or (layer0_outputs(1287)));
    outputs(3698) <= not(layer0_outputs(6835));
    outputs(3699) <= not(layer0_outputs(4936)) or (layer0_outputs(8968));
    outputs(3700) <= not((layer0_outputs(9152)) and (layer0_outputs(3725)));
    outputs(3701) <= not(layer0_outputs(4897));
    outputs(3702) <= layer0_outputs(6010);
    outputs(3703) <= (layer0_outputs(8510)) and not (layer0_outputs(9212));
    outputs(3704) <= not((layer0_outputs(3593)) xor (layer0_outputs(657)));
    outputs(3705) <= layer0_outputs(4916);
    outputs(3706) <= not(layer0_outputs(3285)) or (layer0_outputs(758));
    outputs(3707) <= not(layer0_outputs(5118));
    outputs(3708) <= layer0_outputs(9459);
    outputs(3709) <= (layer0_outputs(5203)) or (layer0_outputs(1446));
    outputs(3710) <= layer0_outputs(2176);
    outputs(3711) <= not((layer0_outputs(1072)) and (layer0_outputs(144)));
    outputs(3712) <= (layer0_outputs(731)) xor (layer0_outputs(9719));
    outputs(3713) <= not(layer0_outputs(2937));
    outputs(3714) <= layer0_outputs(9989);
    outputs(3715) <= (layer0_outputs(103)) xor (layer0_outputs(1266));
    outputs(3716) <= not(layer0_outputs(2559)) or (layer0_outputs(7147));
    outputs(3717) <= not(layer0_outputs(9477));
    outputs(3718) <= not(layer0_outputs(2903));
    outputs(3719) <= layer0_outputs(10156);
    outputs(3720) <= layer0_outputs(8013);
    outputs(3721) <= (layer0_outputs(8893)) xor (layer0_outputs(3958));
    outputs(3722) <= (layer0_outputs(2354)) or (layer0_outputs(616));
    outputs(3723) <= (layer0_outputs(3340)) and not (layer0_outputs(792));
    outputs(3724) <= not(layer0_outputs(1747)) or (layer0_outputs(5737));
    outputs(3725) <= not((layer0_outputs(6738)) xor (layer0_outputs(1751)));
    outputs(3726) <= not(layer0_outputs(3552));
    outputs(3727) <= (layer0_outputs(7683)) xor (layer0_outputs(12129));
    outputs(3728) <= layer0_outputs(12573);
    outputs(3729) <= layer0_outputs(1037);
    outputs(3730) <= (layer0_outputs(3739)) and (layer0_outputs(5984));
    outputs(3731) <= not(layer0_outputs(4906));
    outputs(3732) <= not(layer0_outputs(7529));
    outputs(3733) <= (layer0_outputs(11379)) or (layer0_outputs(1765));
    outputs(3734) <= not(layer0_outputs(2442));
    outputs(3735) <= not(layer0_outputs(4198)) or (layer0_outputs(4508));
    outputs(3736) <= not(layer0_outputs(5321)) or (layer0_outputs(9958));
    outputs(3737) <= (layer0_outputs(7008)) or (layer0_outputs(8754));
    outputs(3738) <= not((layer0_outputs(5303)) xor (layer0_outputs(8937)));
    outputs(3739) <= (layer0_outputs(4355)) and (layer0_outputs(6190));
    outputs(3740) <= not((layer0_outputs(10334)) xor (layer0_outputs(3130)));
    outputs(3741) <= layer0_outputs(3584);
    outputs(3742) <= not((layer0_outputs(10459)) xor (layer0_outputs(9580)));
    outputs(3743) <= (layer0_outputs(6244)) or (layer0_outputs(2433));
    outputs(3744) <= not((layer0_outputs(3427)) xor (layer0_outputs(1137)));
    outputs(3745) <= (layer0_outputs(9566)) and (layer0_outputs(2975));
    outputs(3746) <= not(layer0_outputs(6318));
    outputs(3747) <= (layer0_outputs(959)) and not (layer0_outputs(9006));
    outputs(3748) <= not((layer0_outputs(4312)) or (layer0_outputs(4115)));
    outputs(3749) <= layer0_outputs(6435);
    outputs(3750) <= not(layer0_outputs(12145));
    outputs(3751) <= (layer0_outputs(11915)) or (layer0_outputs(1012));
    outputs(3752) <= not(layer0_outputs(8257)) or (layer0_outputs(157));
    outputs(3753) <= not(layer0_outputs(12775));
    outputs(3754) <= not((layer0_outputs(9598)) xor (layer0_outputs(6621)));
    outputs(3755) <= not(layer0_outputs(3087));
    outputs(3756) <= not((layer0_outputs(9351)) xor (layer0_outputs(2712)));
    outputs(3757) <= layer0_outputs(3164);
    outputs(3758) <= (layer0_outputs(1329)) and not (layer0_outputs(7002));
    outputs(3759) <= layer0_outputs(3078);
    outputs(3760) <= not((layer0_outputs(2348)) xor (layer0_outputs(7095)));
    outputs(3761) <= (layer0_outputs(8511)) and not (layer0_outputs(4894));
    outputs(3762) <= not(layer0_outputs(4027));
    outputs(3763) <= (layer0_outputs(8182)) and not (layer0_outputs(9950));
    outputs(3764) <= (layer0_outputs(10744)) and not (layer0_outputs(2227));
    outputs(3765) <= layer0_outputs(2232);
    outputs(3766) <= not(layer0_outputs(6765));
    outputs(3767) <= not((layer0_outputs(6793)) xor (layer0_outputs(11035)));
    outputs(3768) <= layer0_outputs(10414);
    outputs(3769) <= (layer0_outputs(6188)) and not (layer0_outputs(5182));
    outputs(3770) <= not(layer0_outputs(11116));
    outputs(3771) <= (layer0_outputs(7392)) and (layer0_outputs(12414));
    outputs(3772) <= (layer0_outputs(8940)) and not (layer0_outputs(4259));
    outputs(3773) <= (layer0_outputs(6860)) or (layer0_outputs(1059));
    outputs(3774) <= not(layer0_outputs(240));
    outputs(3775) <= layer0_outputs(3204);
    outputs(3776) <= (layer0_outputs(16)) xor (layer0_outputs(6014));
    outputs(3777) <= (layer0_outputs(10053)) xor (layer0_outputs(5531));
    outputs(3778) <= (layer0_outputs(2980)) xor (layer0_outputs(7215));
    outputs(3779) <= not(layer0_outputs(6048)) or (layer0_outputs(3791));
    outputs(3780) <= not(layer0_outputs(11459));
    outputs(3781) <= (layer0_outputs(12004)) xor (layer0_outputs(3192));
    outputs(3782) <= not(layer0_outputs(720));
    outputs(3783) <= not(layer0_outputs(5743)) or (layer0_outputs(1723));
    outputs(3784) <= (layer0_outputs(7493)) or (layer0_outputs(11609));
    outputs(3785) <= layer0_outputs(9119);
    outputs(3786) <= not((layer0_outputs(2381)) xor (layer0_outputs(10726)));
    outputs(3787) <= not((layer0_outputs(7367)) or (layer0_outputs(136)));
    outputs(3788) <= layer0_outputs(2401);
    outputs(3789) <= (layer0_outputs(5221)) and not (layer0_outputs(8123));
    outputs(3790) <= (layer0_outputs(1773)) xor (layer0_outputs(7536));
    outputs(3791) <= not(layer0_outputs(4218));
    outputs(3792) <= (layer0_outputs(2618)) or (layer0_outputs(2036));
    outputs(3793) <= layer0_outputs(463);
    outputs(3794) <= not((layer0_outputs(9819)) xor (layer0_outputs(6320)));
    outputs(3795) <= layer0_outputs(7597);
    outputs(3796) <= not(layer0_outputs(11111)) or (layer0_outputs(9880));
    outputs(3797) <= (layer0_outputs(3833)) xor (layer0_outputs(10000));
    outputs(3798) <= not((layer0_outputs(11751)) xor (layer0_outputs(261)));
    outputs(3799) <= not(layer0_outputs(1399));
    outputs(3800) <= not(layer0_outputs(4116));
    outputs(3801) <= layer0_outputs(8235);
    outputs(3802) <= (layer0_outputs(2052)) and (layer0_outputs(5346));
    outputs(3803) <= not((layer0_outputs(11934)) and (layer0_outputs(1627)));
    outputs(3804) <= not((layer0_outputs(1771)) and (layer0_outputs(10309)));
    outputs(3805) <= not(layer0_outputs(5187));
    outputs(3806) <= not((layer0_outputs(6911)) xor (layer0_outputs(2775)));
    outputs(3807) <= (layer0_outputs(12157)) or (layer0_outputs(4957));
    outputs(3808) <= (layer0_outputs(2699)) or (layer0_outputs(3977));
    outputs(3809) <= not(layer0_outputs(5519));
    outputs(3810) <= (layer0_outputs(8578)) xor (layer0_outputs(2368));
    outputs(3811) <= not(layer0_outputs(8106));
    outputs(3812) <= not(layer0_outputs(8998)) or (layer0_outputs(4130));
    outputs(3813) <= (layer0_outputs(2380)) and not (layer0_outputs(2988));
    outputs(3814) <= not((layer0_outputs(4116)) or (layer0_outputs(12327)));
    outputs(3815) <= layer0_outputs(3255);
    outputs(3816) <= not((layer0_outputs(1924)) xor (layer0_outputs(11365)));
    outputs(3817) <= (layer0_outputs(8423)) or (layer0_outputs(9235));
    outputs(3818) <= layer0_outputs(3709);
    outputs(3819) <= not((layer0_outputs(3815)) xor (layer0_outputs(2597)));
    outputs(3820) <= not((layer0_outputs(3323)) xor (layer0_outputs(8339)));
    outputs(3821) <= not(layer0_outputs(5035));
    outputs(3822) <= layer0_outputs(4891);
    outputs(3823) <= not(layer0_outputs(11763)) or (layer0_outputs(10836));
    outputs(3824) <= (layer0_outputs(9686)) and (layer0_outputs(10891));
    outputs(3825) <= (layer0_outputs(10581)) xor (layer0_outputs(12036));
    outputs(3826) <= '1';
    outputs(3827) <= (layer0_outputs(9072)) or (layer0_outputs(11440));
    outputs(3828) <= (layer0_outputs(6042)) xor (layer0_outputs(1223));
    outputs(3829) <= (layer0_outputs(6274)) xor (layer0_outputs(9929));
    outputs(3830) <= layer0_outputs(1187);
    outputs(3831) <= not(layer0_outputs(11315));
    outputs(3832) <= not(layer0_outputs(3650)) or (layer0_outputs(11961));
    outputs(3833) <= not(layer0_outputs(3202)) or (layer0_outputs(2508));
    outputs(3834) <= (layer0_outputs(6086)) xor (layer0_outputs(11458));
    outputs(3835) <= not((layer0_outputs(2086)) or (layer0_outputs(2781)));
    outputs(3836) <= (layer0_outputs(12568)) and not (layer0_outputs(10650));
    outputs(3837) <= not(layer0_outputs(8802));
    outputs(3838) <= (layer0_outputs(4591)) xor (layer0_outputs(7683));
    outputs(3839) <= layer0_outputs(10427);
    outputs(3840) <= not(layer0_outputs(5873));
    outputs(3841) <= (layer0_outputs(9246)) or (layer0_outputs(11467));
    outputs(3842) <= (layer0_outputs(10700)) xor (layer0_outputs(11966));
    outputs(3843) <= layer0_outputs(7039);
    outputs(3844) <= (layer0_outputs(859)) and not (layer0_outputs(5627));
    outputs(3845) <= not(layer0_outputs(936));
    outputs(3846) <= layer0_outputs(593);
    outputs(3847) <= (layer0_outputs(1065)) xor (layer0_outputs(89));
    outputs(3848) <= not((layer0_outputs(3205)) or (layer0_outputs(7136)));
    outputs(3849) <= not(layer0_outputs(4423));
    outputs(3850) <= layer0_outputs(405);
    outputs(3851) <= (layer0_outputs(7657)) and (layer0_outputs(948));
    outputs(3852) <= not((layer0_outputs(1436)) xor (layer0_outputs(10011)));
    outputs(3853) <= not((layer0_outputs(7831)) xor (layer0_outputs(11480)));
    outputs(3854) <= layer0_outputs(3410);
    outputs(3855) <= (layer0_outputs(6491)) and (layer0_outputs(10562));
    outputs(3856) <= not(layer0_outputs(2880));
    outputs(3857) <= (layer0_outputs(12784)) xor (layer0_outputs(2582));
    outputs(3858) <= (layer0_outputs(4827)) xor (layer0_outputs(9222));
    outputs(3859) <= not(layer0_outputs(2466));
    outputs(3860) <= layer0_outputs(4320);
    outputs(3861) <= (layer0_outputs(5422)) xor (layer0_outputs(12437));
    outputs(3862) <= layer0_outputs(1436);
    outputs(3863) <= (layer0_outputs(10575)) xor (layer0_outputs(9611));
    outputs(3864) <= not(layer0_outputs(3159));
    outputs(3865) <= not(layer0_outputs(2413)) or (layer0_outputs(537));
    outputs(3866) <= not((layer0_outputs(55)) or (layer0_outputs(269)));
    outputs(3867) <= not(layer0_outputs(7430));
    outputs(3868) <= not(layer0_outputs(1198));
    outputs(3869) <= (layer0_outputs(6879)) xor (layer0_outputs(9720));
    outputs(3870) <= (layer0_outputs(1970)) xor (layer0_outputs(9586));
    outputs(3871) <= not(layer0_outputs(784));
    outputs(3872) <= not(layer0_outputs(7319));
    outputs(3873) <= layer0_outputs(8412);
    outputs(3874) <= not(layer0_outputs(9662));
    outputs(3875) <= layer0_outputs(4898);
    outputs(3876) <= not(layer0_outputs(8800));
    outputs(3877) <= (layer0_outputs(3073)) xor (layer0_outputs(892));
    outputs(3878) <= layer0_outputs(6025);
    outputs(3879) <= layer0_outputs(10161);
    outputs(3880) <= layer0_outputs(9941);
    outputs(3881) <= (layer0_outputs(8310)) xor (layer0_outputs(7100));
    outputs(3882) <= not(layer0_outputs(10235));
    outputs(3883) <= layer0_outputs(7197);
    outputs(3884) <= layer0_outputs(7151);
    outputs(3885) <= layer0_outputs(12080);
    outputs(3886) <= not(layer0_outputs(5051));
    outputs(3887) <= (layer0_outputs(239)) and not (layer0_outputs(7615));
    outputs(3888) <= layer0_outputs(11472);
    outputs(3889) <= not((layer0_outputs(6752)) or (layer0_outputs(12467)));
    outputs(3890) <= not(layer0_outputs(1224));
    outputs(3891) <= not(layer0_outputs(3781));
    outputs(3892) <= layer0_outputs(8081);
    outputs(3893) <= layer0_outputs(9140);
    outputs(3894) <= (layer0_outputs(11412)) or (layer0_outputs(8075));
    outputs(3895) <= layer0_outputs(6238);
    outputs(3896) <= not(layer0_outputs(671)) or (layer0_outputs(147));
    outputs(3897) <= layer0_outputs(4425);
    outputs(3898) <= (layer0_outputs(2927)) xor (layer0_outputs(7803));
    outputs(3899) <= (layer0_outputs(4685)) xor (layer0_outputs(7447));
    outputs(3900) <= (layer0_outputs(8776)) and (layer0_outputs(2307));
    outputs(3901) <= not(layer0_outputs(43));
    outputs(3902) <= not((layer0_outputs(10642)) xor (layer0_outputs(4093)));
    outputs(3903) <= not(layer0_outputs(4757));
    outputs(3904) <= not((layer0_outputs(8159)) xor (layer0_outputs(5765)));
    outputs(3905) <= (layer0_outputs(2762)) or (layer0_outputs(9739));
    outputs(3906) <= layer0_outputs(9085);
    outputs(3907) <= layer0_outputs(6785);
    outputs(3908) <= (layer0_outputs(5016)) and not (layer0_outputs(11747));
    outputs(3909) <= not(layer0_outputs(4665));
    outputs(3910) <= not((layer0_outputs(11726)) xor (layer0_outputs(119)));
    outputs(3911) <= layer0_outputs(8118);
    outputs(3912) <= not((layer0_outputs(4955)) or (layer0_outputs(4589)));
    outputs(3913) <= (layer0_outputs(987)) xor (layer0_outputs(719));
    outputs(3914) <= not(layer0_outputs(7617));
    outputs(3915) <= layer0_outputs(4623);
    outputs(3916) <= (layer0_outputs(2438)) and (layer0_outputs(10448));
    outputs(3917) <= layer0_outputs(5447);
    outputs(3918) <= (layer0_outputs(7706)) xor (layer0_outputs(3875));
    outputs(3919) <= layer0_outputs(11998);
    outputs(3920) <= (layer0_outputs(9599)) xor (layer0_outputs(11378));
    outputs(3921) <= not(layer0_outputs(8588));
    outputs(3922) <= (layer0_outputs(2078)) and not (layer0_outputs(255));
    outputs(3923) <= (layer0_outputs(6847)) and not (layer0_outputs(2488));
    outputs(3924) <= (layer0_outputs(9382)) and not (layer0_outputs(11655));
    outputs(3925) <= (layer0_outputs(571)) and (layer0_outputs(6150));
    outputs(3926) <= not(layer0_outputs(9850)) or (layer0_outputs(10061));
    outputs(3927) <= not(layer0_outputs(777));
    outputs(3928) <= not((layer0_outputs(964)) or (layer0_outputs(2714)));
    outputs(3929) <= not(layer0_outputs(2173));
    outputs(3930) <= (layer0_outputs(1204)) and not (layer0_outputs(430));
    outputs(3931) <= (layer0_outputs(5445)) and not (layer0_outputs(10783));
    outputs(3932) <= not(layer0_outputs(1196)) or (layer0_outputs(3008));
    outputs(3933) <= not(layer0_outputs(106));
    outputs(3934) <= (layer0_outputs(750)) xor (layer0_outputs(471));
    outputs(3935) <= (layer0_outputs(2356)) xor (layer0_outputs(9109));
    outputs(3936) <= layer0_outputs(9716);
    outputs(3937) <= not(layer0_outputs(6432));
    outputs(3938) <= not(layer0_outputs(1738));
    outputs(3939) <= not(layer0_outputs(5303));
    outputs(3940) <= not(layer0_outputs(12286)) or (layer0_outputs(2448));
    outputs(3941) <= not((layer0_outputs(9516)) xor (layer0_outputs(277)));
    outputs(3942) <= (layer0_outputs(1784)) xor (layer0_outputs(5675));
    outputs(3943) <= not((layer0_outputs(9223)) or (layer0_outputs(9174)));
    outputs(3944) <= not(layer0_outputs(11272)) or (layer0_outputs(11719));
    outputs(3945) <= not(layer0_outputs(1911)) or (layer0_outputs(4597));
    outputs(3946) <= not((layer0_outputs(3392)) xor (layer0_outputs(6565)));
    outputs(3947) <= layer0_outputs(8494);
    outputs(3948) <= not(layer0_outputs(5788)) or (layer0_outputs(8468));
    outputs(3949) <= not(layer0_outputs(9417));
    outputs(3950) <= layer0_outputs(6718);
    outputs(3951) <= (layer0_outputs(2695)) or (layer0_outputs(7259));
    outputs(3952) <= not(layer0_outputs(9446));
    outputs(3953) <= layer0_outputs(1798);
    outputs(3954) <= not((layer0_outputs(4288)) xor (layer0_outputs(1824)));
    outputs(3955) <= layer0_outputs(10350);
    outputs(3956) <= layer0_outputs(6815);
    outputs(3957) <= not(layer0_outputs(9892)) or (layer0_outputs(3690));
    outputs(3958) <= (layer0_outputs(10148)) xor (layer0_outputs(9519));
    outputs(3959) <= not(layer0_outputs(5821));
    outputs(3960) <= (layer0_outputs(7909)) xor (layer0_outputs(6715));
    outputs(3961) <= not(layer0_outputs(9853)) or (layer0_outputs(8153));
    outputs(3962) <= not((layer0_outputs(929)) xor (layer0_outputs(9208)));
    outputs(3963) <= (layer0_outputs(12639)) and not (layer0_outputs(12650));
    outputs(3964) <= layer0_outputs(6533);
    outputs(3965) <= not(layer0_outputs(1903));
    outputs(3966) <= not(layer0_outputs(2486));
    outputs(3967) <= not(layer0_outputs(9424));
    outputs(3968) <= not((layer0_outputs(4508)) xor (layer0_outputs(10008)));
    outputs(3969) <= layer0_outputs(475);
    outputs(3970) <= layer0_outputs(3290);
    outputs(3971) <= not(layer0_outputs(841)) or (layer0_outputs(28));
    outputs(3972) <= (layer0_outputs(7962)) and (layer0_outputs(11059));
    outputs(3973) <= not(layer0_outputs(5190)) or (layer0_outputs(10566));
    outputs(3974) <= not((layer0_outputs(11343)) xor (layer0_outputs(2622)));
    outputs(3975) <= not(layer0_outputs(4332));
    outputs(3976) <= (layer0_outputs(4054)) and not (layer0_outputs(1989));
    outputs(3977) <= layer0_outputs(453);
    outputs(3978) <= not(layer0_outputs(10024));
    outputs(3979) <= (layer0_outputs(9579)) xor (layer0_outputs(6051));
    outputs(3980) <= not((layer0_outputs(11129)) xor (layer0_outputs(11846)));
    outputs(3981) <= not(layer0_outputs(7620));
    outputs(3982) <= not((layer0_outputs(5921)) xor (layer0_outputs(68)));
    outputs(3983) <= not(layer0_outputs(4106));
    outputs(3984) <= (layer0_outputs(8612)) or (layer0_outputs(9187));
    outputs(3985) <= not((layer0_outputs(12059)) or (layer0_outputs(20)));
    outputs(3986) <= not(layer0_outputs(10504));
    outputs(3987) <= not((layer0_outputs(4088)) xor (layer0_outputs(7765)));
    outputs(3988) <= not(layer0_outputs(3616));
    outputs(3989) <= not((layer0_outputs(9431)) and (layer0_outputs(12748)));
    outputs(3990) <= not(layer0_outputs(10408)) or (layer0_outputs(3844));
    outputs(3991) <= layer0_outputs(11729);
    outputs(3992) <= (layer0_outputs(681)) and (layer0_outputs(12721));
    outputs(3993) <= layer0_outputs(6393);
    outputs(3994) <= (layer0_outputs(12037)) and not (layer0_outputs(5012));
    outputs(3995) <= not(layer0_outputs(12460));
    outputs(3996) <= layer0_outputs(871);
    outputs(3997) <= layer0_outputs(9269);
    outputs(3998) <= (layer0_outputs(550)) and (layer0_outputs(11340));
    outputs(3999) <= not(layer0_outputs(26)) or (layer0_outputs(3116));
    outputs(4000) <= layer0_outputs(5150);
    outputs(4001) <= not(layer0_outputs(6998));
    outputs(4002) <= layer0_outputs(9554);
    outputs(4003) <= layer0_outputs(8849);
    outputs(4004) <= layer0_outputs(984);
    outputs(4005) <= (layer0_outputs(4245)) xor (layer0_outputs(7910));
    outputs(4006) <= not(layer0_outputs(5305));
    outputs(4007) <= not((layer0_outputs(2277)) xor (layer0_outputs(6461)));
    outputs(4008) <= not((layer0_outputs(10633)) or (layer0_outputs(8954)));
    outputs(4009) <= (layer0_outputs(12432)) xor (layer0_outputs(7893));
    outputs(4010) <= (layer0_outputs(12319)) and not (layer0_outputs(5317));
    outputs(4011) <= layer0_outputs(11000);
    outputs(4012) <= (layer0_outputs(4149)) or (layer0_outputs(10254));
    outputs(4013) <= not(layer0_outputs(2566));
    outputs(4014) <= not((layer0_outputs(2879)) xor (layer0_outputs(6222)));
    outputs(4015) <= layer0_outputs(5282);
    outputs(4016) <= not((layer0_outputs(6534)) xor (layer0_outputs(4972)));
    outputs(4017) <= not(layer0_outputs(7214)) or (layer0_outputs(5986));
    outputs(4018) <= not((layer0_outputs(2605)) or (layer0_outputs(9067)));
    outputs(4019) <= not(layer0_outputs(12158));
    outputs(4020) <= not(layer0_outputs(9923));
    outputs(4021) <= not((layer0_outputs(5522)) xor (layer0_outputs(2595)));
    outputs(4022) <= not((layer0_outputs(4712)) and (layer0_outputs(7474)));
    outputs(4023) <= (layer0_outputs(11642)) and (layer0_outputs(3173));
    outputs(4024) <= not((layer0_outputs(1832)) xor (layer0_outputs(3274)));
    outputs(4025) <= not(layer0_outputs(10143));
    outputs(4026) <= (layer0_outputs(6726)) or (layer0_outputs(5613));
    outputs(4027) <= (layer0_outputs(12001)) xor (layer0_outputs(5323));
    outputs(4028) <= (layer0_outputs(573)) and not (layer0_outputs(11937));
    outputs(4029) <= (layer0_outputs(12583)) and not (layer0_outputs(5005));
    outputs(4030) <= (layer0_outputs(4122)) xor (layer0_outputs(4026));
    outputs(4031) <= layer0_outputs(3673);
    outputs(4032) <= not(layer0_outputs(5914));
    outputs(4033) <= not((layer0_outputs(5437)) or (layer0_outputs(943)));
    outputs(4034) <= not(layer0_outputs(5919));
    outputs(4035) <= (layer0_outputs(1399)) or (layer0_outputs(9150));
    outputs(4036) <= not(layer0_outputs(4813));
    outputs(4037) <= (layer0_outputs(12590)) xor (layer0_outputs(11686));
    outputs(4038) <= not((layer0_outputs(12181)) and (layer0_outputs(6005)));
    outputs(4039) <= (layer0_outputs(5230)) xor (layer0_outputs(7783));
    outputs(4040) <= layer0_outputs(4966);
    outputs(4041) <= (layer0_outputs(7382)) or (layer0_outputs(9991));
    outputs(4042) <= (layer0_outputs(7035)) and not (layer0_outputs(2208));
    outputs(4043) <= not(layer0_outputs(4094)) or (layer0_outputs(1127));
    outputs(4044) <= not(layer0_outputs(9355));
    outputs(4045) <= not((layer0_outputs(9864)) xor (layer0_outputs(11708)));
    outputs(4046) <= layer0_outputs(10719);
    outputs(4047) <= not((layer0_outputs(1153)) and (layer0_outputs(10174)));
    outputs(4048) <= not((layer0_outputs(9277)) xor (layer0_outputs(10145)));
    outputs(4049) <= not(layer0_outputs(7023)) or (layer0_outputs(1346));
    outputs(4050) <= layer0_outputs(10107);
    outputs(4051) <= not(layer0_outputs(8860));
    outputs(4052) <= (layer0_outputs(6772)) xor (layer0_outputs(10583));
    outputs(4053) <= (layer0_outputs(6424)) xor (layer0_outputs(9277));
    outputs(4054) <= (layer0_outputs(9533)) and not (layer0_outputs(3286));
    outputs(4055) <= not(layer0_outputs(7703));
    outputs(4056) <= not((layer0_outputs(1721)) and (layer0_outputs(9429)));
    outputs(4057) <= not((layer0_outputs(633)) and (layer0_outputs(1569)));
    outputs(4058) <= (layer0_outputs(12071)) xor (layer0_outputs(8691));
    outputs(4059) <= layer0_outputs(2823);
    outputs(4060) <= (layer0_outputs(1697)) and not (layer0_outputs(10269));
    outputs(4061) <= layer0_outputs(10428);
    outputs(4062) <= (layer0_outputs(4267)) xor (layer0_outputs(7518));
    outputs(4063) <= (layer0_outputs(3533)) and (layer0_outputs(2485));
    outputs(4064) <= (layer0_outputs(10847)) and not (layer0_outputs(3847));
    outputs(4065) <= not(layer0_outputs(10126));
    outputs(4066) <= (layer0_outputs(11815)) and not (layer0_outputs(7134));
    outputs(4067) <= not((layer0_outputs(4362)) or (layer0_outputs(6620)));
    outputs(4068) <= layer0_outputs(7277);
    outputs(4069) <= not(layer0_outputs(6298));
    outputs(4070) <= not(layer0_outputs(456));
    outputs(4071) <= not((layer0_outputs(11343)) xor (layer0_outputs(6845)));
    outputs(4072) <= (layer0_outputs(4519)) xor (layer0_outputs(9623));
    outputs(4073) <= not(layer0_outputs(9518)) or (layer0_outputs(10337));
    outputs(4074) <= (layer0_outputs(615)) xor (layer0_outputs(10820));
    outputs(4075) <= layer0_outputs(2292);
    outputs(4076) <= not(layer0_outputs(575));
    outputs(4077) <= not((layer0_outputs(7368)) xor (layer0_outputs(1864)));
    outputs(4078) <= not((layer0_outputs(11296)) or (layer0_outputs(656)));
    outputs(4079) <= layer0_outputs(4492);
    outputs(4080) <= not((layer0_outputs(2764)) xor (layer0_outputs(6246)));
    outputs(4081) <= not(layer0_outputs(5688));
    outputs(4082) <= layer0_outputs(448);
    outputs(4083) <= (layer0_outputs(11703)) xor (layer0_outputs(9029));
    outputs(4084) <= (layer0_outputs(7398)) and not (layer0_outputs(691));
    outputs(4085) <= not(layer0_outputs(11196));
    outputs(4086) <= not(layer0_outputs(4761)) or (layer0_outputs(6550));
    outputs(4087) <= (layer0_outputs(2067)) xor (layer0_outputs(9600));
    outputs(4088) <= not((layer0_outputs(12759)) xor (layer0_outputs(11666)));
    outputs(4089) <= layer0_outputs(1750);
    outputs(4090) <= not((layer0_outputs(727)) xor (layer0_outputs(7537)));
    outputs(4091) <= (layer0_outputs(7066)) xor (layer0_outputs(2821));
    outputs(4092) <= not((layer0_outputs(1755)) and (layer0_outputs(9096)));
    outputs(4093) <= not(layer0_outputs(527)) or (layer0_outputs(8167));
    outputs(4094) <= (layer0_outputs(9813)) and not (layer0_outputs(1089));
    outputs(4095) <= not((layer0_outputs(12640)) or (layer0_outputs(4707)));
    outputs(4096) <= not(layer0_outputs(2083));
    outputs(4097) <= not(layer0_outputs(6060)) or (layer0_outputs(3233));
    outputs(4098) <= not(layer0_outputs(10282));
    outputs(4099) <= not((layer0_outputs(1264)) or (layer0_outputs(4047)));
    outputs(4100) <= (layer0_outputs(12083)) and not (layer0_outputs(5057));
    outputs(4101) <= (layer0_outputs(4526)) and (layer0_outputs(6849));
    outputs(4102) <= not(layer0_outputs(11090));
    outputs(4103) <= (layer0_outputs(8319)) xor (layer0_outputs(2373));
    outputs(4104) <= not(layer0_outputs(6770));
    outputs(4105) <= (layer0_outputs(10767)) or (layer0_outputs(3193));
    outputs(4106) <= not((layer0_outputs(6816)) xor (layer0_outputs(8933)));
    outputs(4107) <= layer0_outputs(8118);
    outputs(4108) <= not((layer0_outputs(11395)) xor (layer0_outputs(4057)));
    outputs(4109) <= not(layer0_outputs(12126));
    outputs(4110) <= not(layer0_outputs(2984));
    outputs(4111) <= (layer0_outputs(753)) xor (layer0_outputs(9390));
    outputs(4112) <= (layer0_outputs(4160)) and not (layer0_outputs(7708));
    outputs(4113) <= not(layer0_outputs(112));
    outputs(4114) <= layer0_outputs(8907);
    outputs(4115) <= not((layer0_outputs(8295)) and (layer0_outputs(10729)));
    outputs(4116) <= (layer0_outputs(3419)) xor (layer0_outputs(1207));
    outputs(4117) <= layer0_outputs(2445);
    outputs(4118) <= not((layer0_outputs(645)) xor (layer0_outputs(5017)));
    outputs(4119) <= layer0_outputs(3197);
    outputs(4120) <= layer0_outputs(8463);
    outputs(4121) <= not(layer0_outputs(1766));
    outputs(4122) <= (layer0_outputs(5934)) and (layer0_outputs(477));
    outputs(4123) <= not(layer0_outputs(12536)) or (layer0_outputs(2832));
    outputs(4124) <= layer0_outputs(3024);
    outputs(4125) <= not(layer0_outputs(866));
    outputs(4126) <= not(layer0_outputs(6483)) or (layer0_outputs(10790));
    outputs(4127) <= (layer0_outputs(10622)) xor (layer0_outputs(6139));
    outputs(4128) <= not(layer0_outputs(5254));
    outputs(4129) <= not((layer0_outputs(9129)) xor (layer0_outputs(8377)));
    outputs(4130) <= not(layer0_outputs(7680));
    outputs(4131) <= (layer0_outputs(7367)) xor (layer0_outputs(2565));
    outputs(4132) <= layer0_outputs(11049);
    outputs(4133) <= (layer0_outputs(11488)) and not (layer0_outputs(138));
    outputs(4134) <= not((layer0_outputs(10063)) xor (layer0_outputs(10961)));
    outputs(4135) <= layer0_outputs(10071);
    outputs(4136) <= (layer0_outputs(6477)) xor (layer0_outputs(3807));
    outputs(4137) <= not(layer0_outputs(11496));
    outputs(4138) <= layer0_outputs(801);
    outputs(4139) <= not((layer0_outputs(2630)) xor (layer0_outputs(12248)));
    outputs(4140) <= not((layer0_outputs(1395)) xor (layer0_outputs(10388)));
    outputs(4141) <= not((layer0_outputs(3976)) and (layer0_outputs(6030)));
    outputs(4142) <= not((layer0_outputs(9768)) xor (layer0_outputs(8649)));
    outputs(4143) <= not(layer0_outputs(6282)) or (layer0_outputs(11316));
    outputs(4144) <= not(layer0_outputs(9391));
    outputs(4145) <= (layer0_outputs(6485)) and not (layer0_outputs(8435));
    outputs(4146) <= (layer0_outputs(8329)) xor (layer0_outputs(2985));
    outputs(4147) <= not((layer0_outputs(2839)) xor (layer0_outputs(4849)));
    outputs(4148) <= (layer0_outputs(11577)) or (layer0_outputs(2255));
    outputs(4149) <= layer0_outputs(8271);
    outputs(4150) <= (layer0_outputs(11590)) xor (layer0_outputs(696));
    outputs(4151) <= (layer0_outputs(8523)) and not (layer0_outputs(2072));
    outputs(4152) <= not((layer0_outputs(1756)) or (layer0_outputs(1380)));
    outputs(4153) <= (layer0_outputs(6474)) xor (layer0_outputs(6362));
    outputs(4154) <= (layer0_outputs(8179)) and not (layer0_outputs(6689));
    outputs(4155) <= layer0_outputs(6473);
    outputs(4156) <= (layer0_outputs(5013)) xor (layer0_outputs(11629));
    outputs(4157) <= (layer0_outputs(12498)) or (layer0_outputs(11650));
    outputs(4158) <= not(layer0_outputs(9029)) or (layer0_outputs(4089));
    outputs(4159) <= not(layer0_outputs(3548));
    outputs(4160) <= not(layer0_outputs(9306));
    outputs(4161) <= (layer0_outputs(2877)) and not (layer0_outputs(1894));
    outputs(4162) <= (layer0_outputs(3929)) xor (layer0_outputs(12054));
    outputs(4163) <= (layer0_outputs(5978)) xor (layer0_outputs(9727));
    outputs(4164) <= (layer0_outputs(10531)) xor (layer0_outputs(10070));
    outputs(4165) <= not(layer0_outputs(10950));
    outputs(4166) <= (layer0_outputs(12115)) xor (layer0_outputs(5425));
    outputs(4167) <= layer0_outputs(9060);
    outputs(4168) <= not(layer0_outputs(7312));
    outputs(4169) <= not(layer0_outputs(4355)) or (layer0_outputs(906));
    outputs(4170) <= not(layer0_outputs(9559));
    outputs(4171) <= (layer0_outputs(7739)) xor (layer0_outputs(3151));
    outputs(4172) <= (layer0_outputs(4754)) and not (layer0_outputs(4944));
    outputs(4173) <= layer0_outputs(4867);
    outputs(4174) <= not(layer0_outputs(12657));
    outputs(4175) <= layer0_outputs(3748);
    outputs(4176) <= not((layer0_outputs(8281)) xor (layer0_outputs(9992)));
    outputs(4177) <= not(layer0_outputs(4520));
    outputs(4178) <= layer0_outputs(4476);
    outputs(4179) <= (layer0_outputs(8348)) xor (layer0_outputs(4798));
    outputs(4180) <= (layer0_outputs(11932)) or (layer0_outputs(9757));
    outputs(4181) <= not(layer0_outputs(12144)) or (layer0_outputs(9960));
    outputs(4182) <= not(layer0_outputs(9209)) or (layer0_outputs(4914));
    outputs(4183) <= not(layer0_outputs(1847));
    outputs(4184) <= not((layer0_outputs(2948)) xor (layer0_outputs(6776)));
    outputs(4185) <= not((layer0_outputs(7185)) or (layer0_outputs(11730)));
    outputs(4186) <= not(layer0_outputs(2880));
    outputs(4187) <= not(layer0_outputs(12496));
    outputs(4188) <= layer0_outputs(3857);
    outputs(4189) <= not(layer0_outputs(3092)) or (layer0_outputs(5822));
    outputs(4190) <= not(layer0_outputs(5530));
    outputs(4191) <= layer0_outputs(2493);
    outputs(4192) <= (layer0_outputs(7865)) and not (layer0_outputs(3841));
    outputs(4193) <= not(layer0_outputs(8955));
    outputs(4194) <= not((layer0_outputs(3823)) xor (layer0_outputs(5131)));
    outputs(4195) <= layer0_outputs(3020);
    outputs(4196) <= not((layer0_outputs(12352)) xor (layer0_outputs(907)));
    outputs(4197) <= layer0_outputs(7041);
    outputs(4198) <= (layer0_outputs(891)) and not (layer0_outputs(11937));
    outputs(4199) <= layer0_outputs(2536);
    outputs(4200) <= not((layer0_outputs(3067)) xor (layer0_outputs(7921)));
    outputs(4201) <= layer0_outputs(11803);
    outputs(4202) <= layer0_outputs(6928);
    outputs(4203) <= not(layer0_outputs(3307));
    outputs(4204) <= not(layer0_outputs(6041));
    outputs(4205) <= not(layer0_outputs(12398));
    outputs(4206) <= not(layer0_outputs(9594));
    outputs(4207) <= layer0_outputs(6596);
    outputs(4208) <= (layer0_outputs(9357)) and (layer0_outputs(12574));
    outputs(4209) <= layer0_outputs(536);
    outputs(4210) <= not((layer0_outputs(10792)) xor (layer0_outputs(6612)));
    outputs(4211) <= not((layer0_outputs(11369)) xor (layer0_outputs(40)));
    outputs(4212) <= (layer0_outputs(2515)) and (layer0_outputs(4403));
    outputs(4213) <= layer0_outputs(10671);
    outputs(4214) <= not((layer0_outputs(2646)) or (layer0_outputs(7474)));
    outputs(4215) <= layer0_outputs(8037);
    outputs(4216) <= (layer0_outputs(5132)) and (layer0_outputs(4203));
    outputs(4217) <= (layer0_outputs(64)) and not (layer0_outputs(2));
    outputs(4218) <= (layer0_outputs(10169)) and (layer0_outputs(4363));
    outputs(4219) <= layer0_outputs(2078);
    outputs(4220) <= not(layer0_outputs(5233));
    outputs(4221) <= (layer0_outputs(10348)) xor (layer0_outputs(4315));
    outputs(4222) <= not(layer0_outputs(444));
    outputs(4223) <= (layer0_outputs(9272)) xor (layer0_outputs(1042));
    outputs(4224) <= (layer0_outputs(8426)) and not (layer0_outputs(9341));
    outputs(4225) <= not((layer0_outputs(4059)) or (layer0_outputs(3967)));
    outputs(4226) <= (layer0_outputs(11847)) xor (layer0_outputs(3438));
    outputs(4227) <= (layer0_outputs(1060)) xor (layer0_outputs(3516));
    outputs(4228) <= layer0_outputs(3069);
    outputs(4229) <= not((layer0_outputs(7594)) or (layer0_outputs(7409)));
    outputs(4230) <= not(layer0_outputs(5341));
    outputs(4231) <= layer0_outputs(5426);
    outputs(4232) <= not((layer0_outputs(4019)) and (layer0_outputs(9601)));
    outputs(4233) <= not((layer0_outputs(3134)) or (layer0_outputs(1845)));
    outputs(4234) <= layer0_outputs(11832);
    outputs(4235) <= (layer0_outputs(7716)) xor (layer0_outputs(9456));
    outputs(4236) <= (layer0_outputs(1093)) and (layer0_outputs(9499));
    outputs(4237) <= layer0_outputs(1630);
    outputs(4238) <= not((layer0_outputs(5495)) or (layer0_outputs(626)));
    outputs(4239) <= (layer0_outputs(2535)) xor (layer0_outputs(1909));
    outputs(4240) <= (layer0_outputs(9508)) and (layer0_outputs(3394));
    outputs(4241) <= not((layer0_outputs(3646)) xor (layer0_outputs(6349)));
    outputs(4242) <= not(layer0_outputs(6368)) or (layer0_outputs(1132));
    outputs(4243) <= (layer0_outputs(5289)) and (layer0_outputs(2347));
    outputs(4244) <= (layer0_outputs(5619)) xor (layer0_outputs(5304));
    outputs(4245) <= (layer0_outputs(11570)) and (layer0_outputs(11973));
    outputs(4246) <= layer0_outputs(3916);
    outputs(4247) <= not(layer0_outputs(3852));
    outputs(4248) <= not((layer0_outputs(5796)) xor (layer0_outputs(454)));
    outputs(4249) <= not((layer0_outputs(3015)) xor (layer0_outputs(2260)));
    outputs(4250) <= not((layer0_outputs(5885)) or (layer0_outputs(7464)));
    outputs(4251) <= not((layer0_outputs(9013)) and (layer0_outputs(1841)));
    outputs(4252) <= (layer0_outputs(1489)) xor (layer0_outputs(1434));
    outputs(4253) <= layer0_outputs(5889);
    outputs(4254) <= (layer0_outputs(11964)) xor (layer0_outputs(713));
    outputs(4255) <= layer0_outputs(6607);
    outputs(4256) <= not((layer0_outputs(10093)) or (layer0_outputs(12190)));
    outputs(4257) <= not(layer0_outputs(5000));
    outputs(4258) <= (layer0_outputs(7511)) and not (layer0_outputs(6518));
    outputs(4259) <= (layer0_outputs(3494)) xor (layer0_outputs(5288));
    outputs(4260) <= layer0_outputs(5541);
    outputs(4261) <= layer0_outputs(4800);
    outputs(4262) <= layer0_outputs(258);
    outputs(4263) <= not((layer0_outputs(364)) and (layer0_outputs(5049)));
    outputs(4264) <= layer0_outputs(12240);
    outputs(4265) <= layer0_outputs(9883);
    outputs(4266) <= (layer0_outputs(4631)) and (layer0_outputs(272));
    outputs(4267) <= (layer0_outputs(6520)) and (layer0_outputs(1961));
    outputs(4268) <= (layer0_outputs(9914)) and not (layer0_outputs(8398));
    outputs(4269) <= not(layer0_outputs(8338));
    outputs(4270) <= not(layer0_outputs(893));
    outputs(4271) <= not(layer0_outputs(5572));
    outputs(4272) <= layer0_outputs(5911);
    outputs(4273) <= (layer0_outputs(3397)) xor (layer0_outputs(4609));
    outputs(4274) <= not((layer0_outputs(4059)) or (layer0_outputs(4674)));
    outputs(4275) <= (layer0_outputs(2469)) xor (layer0_outputs(9683));
    outputs(4276) <= (layer0_outputs(226)) xor (layer0_outputs(7745));
    outputs(4277) <= layer0_outputs(7408);
    outputs(4278) <= layer0_outputs(8422);
    outputs(4279) <= (layer0_outputs(12742)) xor (layer0_outputs(9430));
    outputs(4280) <= not(layer0_outputs(9077));
    outputs(4281) <= (layer0_outputs(2862)) and (layer0_outputs(3846));
    outputs(4282) <= (layer0_outputs(1757)) and not (layer0_outputs(3837));
    outputs(4283) <= not(layer0_outputs(2904));
    outputs(4284) <= not((layer0_outputs(8166)) xor (layer0_outputs(4829)));
    outputs(4285) <= (layer0_outputs(5448)) and not (layer0_outputs(7632));
    outputs(4286) <= not(layer0_outputs(10772));
    outputs(4287) <= not(layer0_outputs(2731));
    outputs(4288) <= not(layer0_outputs(6420)) or (layer0_outputs(4948));
    outputs(4289) <= (layer0_outputs(3947)) xor (layer0_outputs(914));
    outputs(4290) <= not(layer0_outputs(9249));
    outputs(4291) <= not((layer0_outputs(5787)) and (layer0_outputs(1137)));
    outputs(4292) <= (layer0_outputs(623)) or (layer0_outputs(6278));
    outputs(4293) <= not((layer0_outputs(5361)) xor (layer0_outputs(4173)));
    outputs(4294) <= not(layer0_outputs(5965));
    outputs(4295) <= (layer0_outputs(10690)) and not (layer0_outputs(11677));
    outputs(4296) <= (layer0_outputs(7842)) or (layer0_outputs(6026));
    outputs(4297) <= (layer0_outputs(9064)) xor (layer0_outputs(918));
    outputs(4298) <= (layer0_outputs(24)) xor (layer0_outputs(7704));
    outputs(4299) <= not(layer0_outputs(8121));
    outputs(4300) <= (layer0_outputs(10067)) or (layer0_outputs(11603));
    outputs(4301) <= not(layer0_outputs(2900));
    outputs(4302) <= not(layer0_outputs(935));
    outputs(4303) <= (layer0_outputs(7917)) xor (layer0_outputs(1681));
    outputs(4304) <= not((layer0_outputs(11164)) xor (layer0_outputs(11893)));
    outputs(4305) <= not(layer0_outputs(1317));
    outputs(4306) <= (layer0_outputs(3948)) and (layer0_outputs(5794));
    outputs(4307) <= not(layer0_outputs(7300));
    outputs(4308) <= (layer0_outputs(4978)) xor (layer0_outputs(1607));
    outputs(4309) <= not((layer0_outputs(7168)) or (layer0_outputs(1120)));
    outputs(4310) <= not(layer0_outputs(12191)) or (layer0_outputs(5647));
    outputs(4311) <= not((layer0_outputs(1348)) xor (layer0_outputs(3499)));
    outputs(4312) <= (layer0_outputs(12222)) xor (layer0_outputs(9175));
    outputs(4313) <= (layer0_outputs(12011)) xor (layer0_outputs(10609));
    outputs(4314) <= not((layer0_outputs(8108)) and (layer0_outputs(8583)));
    outputs(4315) <= (layer0_outputs(8354)) and not (layer0_outputs(3664));
    outputs(4316) <= not(layer0_outputs(12439)) or (layer0_outputs(9472));
    outputs(4317) <= layer0_outputs(8916);
    outputs(4318) <= layer0_outputs(8863);
    outputs(4319) <= layer0_outputs(4370);
    outputs(4320) <= not((layer0_outputs(10568)) xor (layer0_outputs(7795)));
    outputs(4321) <= (layer0_outputs(10721)) and (layer0_outputs(5923));
    outputs(4322) <= (layer0_outputs(8250)) and (layer0_outputs(12236));
    outputs(4323) <= (layer0_outputs(2389)) and not (layer0_outputs(6366));
    outputs(4324) <= (layer0_outputs(2697)) xor (layer0_outputs(507));
    outputs(4325) <= not((layer0_outputs(579)) xor (layer0_outputs(10001)));
    outputs(4326) <= (layer0_outputs(3676)) xor (layer0_outputs(8387));
    outputs(4327) <= not((layer0_outputs(12474)) xor (layer0_outputs(7573)));
    outputs(4328) <= not(layer0_outputs(3569)) or (layer0_outputs(945));
    outputs(4329) <= not((layer0_outputs(5750)) xor (layer0_outputs(9166)));
    outputs(4330) <= not((layer0_outputs(1248)) and (layer0_outputs(11326)));
    outputs(4331) <= not((layer0_outputs(10884)) xor (layer0_outputs(2989)));
    outputs(4332) <= layer0_outputs(11593);
    outputs(4333) <= layer0_outputs(1275);
    outputs(4334) <= not(layer0_outputs(3136)) or (layer0_outputs(8561));
    outputs(4335) <= (layer0_outputs(10074)) xor (layer0_outputs(3758));
    outputs(4336) <= not(layer0_outputs(6369));
    outputs(4337) <= layer0_outputs(4171);
    outputs(4338) <= not(layer0_outputs(4604)) or (layer0_outputs(7053));
    outputs(4339) <= layer0_outputs(1584);
    outputs(4340) <= not(layer0_outputs(2540));
    outputs(4341) <= (layer0_outputs(11762)) and (layer0_outputs(8748));
    outputs(4342) <= (layer0_outputs(7574)) and not (layer0_outputs(10413));
    outputs(4343) <= (layer0_outputs(8347)) and (layer0_outputs(237));
    outputs(4344) <= not(layer0_outputs(7572));
    outputs(4345) <= not((layer0_outputs(2104)) or (layer0_outputs(596)));
    outputs(4346) <= not((layer0_outputs(11789)) xor (layer0_outputs(6165)));
    outputs(4347) <= layer0_outputs(7335);
    outputs(4348) <= not((layer0_outputs(9253)) xor (layer0_outputs(649)));
    outputs(4349) <= not(layer0_outputs(9510)) or (layer0_outputs(1899));
    outputs(4350) <= (layer0_outputs(5081)) and not (layer0_outputs(6819));
    outputs(4351) <= not((layer0_outputs(4652)) xor (layer0_outputs(4932)));
    outputs(4352) <= not((layer0_outputs(4548)) xor (layer0_outputs(3624)));
    outputs(4353) <= (layer0_outputs(8471)) xor (layer0_outputs(7547));
    outputs(4354) <= not(layer0_outputs(3910));
    outputs(4355) <= layer0_outputs(5794);
    outputs(4356) <= (layer0_outputs(9563)) xor (layer0_outputs(10410));
    outputs(4357) <= layer0_outputs(10858);
    outputs(4358) <= layer0_outputs(6280);
    outputs(4359) <= (layer0_outputs(7736)) and not (layer0_outputs(11405));
    outputs(4360) <= not(layer0_outputs(11631));
    outputs(4361) <= (layer0_outputs(3671)) and not (layer0_outputs(4179));
    outputs(4362) <= not((layer0_outputs(8156)) and (layer0_outputs(12351)));
    outputs(4363) <= layer0_outputs(7029);
    outputs(4364) <= (layer0_outputs(4120)) and (layer0_outputs(1640));
    outputs(4365) <= not(layer0_outputs(12618));
    outputs(4366) <= layer0_outputs(4573);
    outputs(4367) <= not((layer0_outputs(5409)) xor (layer0_outputs(10662)));
    outputs(4368) <= (layer0_outputs(5180)) and (layer0_outputs(9393));
    outputs(4369) <= not((layer0_outputs(9238)) xor (layer0_outputs(6501)));
    outputs(4370) <= layer0_outputs(11547);
    outputs(4371) <= not(layer0_outputs(5036)) or (layer0_outputs(1935));
    outputs(4372) <= (layer0_outputs(3401)) and (layer0_outputs(3719));
    outputs(4373) <= not(layer0_outputs(10239));
    outputs(4374) <= layer0_outputs(9796);
    outputs(4375) <= layer0_outputs(1069);
    outputs(4376) <= not(layer0_outputs(5479));
    outputs(4377) <= not(layer0_outputs(9739)) or (layer0_outputs(1424));
    outputs(4378) <= not((layer0_outputs(2878)) xor (layer0_outputs(5433)));
    outputs(4379) <= not((layer0_outputs(12593)) xor (layer0_outputs(2172)));
    outputs(4380) <= not(layer0_outputs(7181));
    outputs(4381) <= not(layer0_outputs(908)) or (layer0_outputs(391));
    outputs(4382) <= not((layer0_outputs(7719)) or (layer0_outputs(3167)));
    outputs(4383) <= not(layer0_outputs(2504));
    outputs(4384) <= (layer0_outputs(987)) xor (layer0_outputs(10426));
    outputs(4385) <= (layer0_outputs(7530)) or (layer0_outputs(9293));
    outputs(4386) <= not((layer0_outputs(10862)) xor (layer0_outputs(2331)));
    outputs(4387) <= not((layer0_outputs(1408)) or (layer0_outputs(7219)));
    outputs(4388) <= not((layer0_outputs(10368)) xor (layer0_outputs(10273)));
    outputs(4389) <= layer0_outputs(891);
    outputs(4390) <= not(layer0_outputs(1268));
    outputs(4391) <= not((layer0_outputs(5842)) xor (layer0_outputs(9199)));
    outputs(4392) <= layer0_outputs(11048);
    outputs(4393) <= layer0_outputs(11220);
    outputs(4394) <= not(layer0_outputs(5795));
    outputs(4395) <= not(layer0_outputs(9318));
    outputs(4396) <= layer0_outputs(991);
    outputs(4397) <= (layer0_outputs(172)) or (layer0_outputs(5112));
    outputs(4398) <= not(layer0_outputs(8152)) or (layer0_outputs(3448));
    outputs(4399) <= layer0_outputs(6557);
    outputs(4400) <= layer0_outputs(6467);
    outputs(4401) <= not(layer0_outputs(7231));
    outputs(4402) <= not(layer0_outputs(5878)) or (layer0_outputs(12066));
    outputs(4403) <= not((layer0_outputs(10658)) xor (layer0_outputs(6235)));
    outputs(4404) <= not((layer0_outputs(3170)) xor (layer0_outputs(3611)));
    outputs(4405) <= layer0_outputs(5294);
    outputs(4406) <= not(layer0_outputs(390));
    outputs(4407) <= not(layer0_outputs(2395));
    outputs(4408) <= (layer0_outputs(3256)) or (layer0_outputs(4391));
    outputs(4409) <= (layer0_outputs(7946)) xor (layer0_outputs(6314));
    outputs(4410) <= not(layer0_outputs(2841));
    outputs(4411) <= layer0_outputs(8177);
    outputs(4412) <= (layer0_outputs(1883)) xor (layer0_outputs(6204));
    outputs(4413) <= not(layer0_outputs(10985));
    outputs(4414) <= layer0_outputs(3741);
    outputs(4415) <= (layer0_outputs(4321)) and not (layer0_outputs(2410));
    outputs(4416) <= (layer0_outputs(11037)) and not (layer0_outputs(6376));
    outputs(4417) <= not(layer0_outputs(7531));
    outputs(4418) <= not(layer0_outputs(4121));
    outputs(4419) <= not(layer0_outputs(8216));
    outputs(4420) <= (layer0_outputs(226)) xor (layer0_outputs(4592));
    outputs(4421) <= not((layer0_outputs(12153)) and (layer0_outputs(6688)));
    outputs(4422) <= not((layer0_outputs(8602)) or (layer0_outputs(6574)));
    outputs(4423) <= layer0_outputs(6280);
    outputs(4424) <= (layer0_outputs(2957)) xor (layer0_outputs(5997));
    outputs(4425) <= not((layer0_outputs(10041)) and (layer0_outputs(6727)));
    outputs(4426) <= (layer0_outputs(971)) and not (layer0_outputs(9206));
    outputs(4427) <= (layer0_outputs(3192)) xor (layer0_outputs(431));
    outputs(4428) <= (layer0_outputs(10265)) xor (layer0_outputs(10123));
    outputs(4429) <= not((layer0_outputs(2441)) xor (layer0_outputs(8453)));
    outputs(4430) <= (layer0_outputs(4734)) and (layer0_outputs(9560));
    outputs(4431) <= not(layer0_outputs(9595));
    outputs(4432) <= (layer0_outputs(6552)) and not (layer0_outputs(10653));
    outputs(4433) <= not((layer0_outputs(4157)) xor (layer0_outputs(812)));
    outputs(4434) <= not((layer0_outputs(555)) xor (layer0_outputs(7461)));
    outputs(4435) <= (layer0_outputs(12537)) and not (layer0_outputs(7459));
    outputs(4436) <= layer0_outputs(7936);
    outputs(4437) <= (layer0_outputs(8541)) xor (layer0_outputs(11290));
    outputs(4438) <= layer0_outputs(2193);
    outputs(4439) <= not((layer0_outputs(11003)) or (layer0_outputs(6648)));
    outputs(4440) <= (layer0_outputs(10346)) xor (layer0_outputs(10367));
    outputs(4441) <= not(layer0_outputs(8294));
    outputs(4442) <= layer0_outputs(1901);
    outputs(4443) <= layer0_outputs(11519);
    outputs(4444) <= (layer0_outputs(8895)) xor (layer0_outputs(6837));
    outputs(4445) <= (layer0_outputs(9393)) xor (layer0_outputs(6071));
    outputs(4446) <= layer0_outputs(666);
    outputs(4447) <= not((layer0_outputs(2262)) or (layer0_outputs(12660)));
    outputs(4448) <= (layer0_outputs(4371)) xor (layer0_outputs(10209));
    outputs(4449) <= (layer0_outputs(8497)) and (layer0_outputs(8666));
    outputs(4450) <= (layer0_outputs(12484)) and not (layer0_outputs(11062));
    outputs(4451) <= not(layer0_outputs(8750));
    outputs(4452) <= (layer0_outputs(2500)) and (layer0_outputs(2105));
    outputs(4453) <= not((layer0_outputs(5411)) or (layer0_outputs(4946)));
    outputs(4454) <= layer0_outputs(388);
    outputs(4455) <= not(layer0_outputs(9797));
    outputs(4456) <= not(layer0_outputs(6321));
    outputs(4457) <= (layer0_outputs(8989)) and not (layer0_outputs(5843));
    outputs(4458) <= layer0_outputs(9586);
    outputs(4459) <= not((layer0_outputs(11248)) and (layer0_outputs(8256)));
    outputs(4460) <= (layer0_outputs(10506)) xor (layer0_outputs(10395));
    outputs(4461) <= not(layer0_outputs(12677));
    outputs(4462) <= (layer0_outputs(10907)) and not (layer0_outputs(8197));
    outputs(4463) <= (layer0_outputs(7638)) and not (layer0_outputs(11598));
    outputs(4464) <= (layer0_outputs(7261)) and not (layer0_outputs(8406));
    outputs(4465) <= not(layer0_outputs(7869));
    outputs(4466) <= not((layer0_outputs(752)) xor (layer0_outputs(10732)));
    outputs(4467) <= layer0_outputs(12271);
    outputs(4468) <= (layer0_outputs(12652)) and not (layer0_outputs(1339));
    outputs(4469) <= layer0_outputs(3189);
    outputs(4470) <= not(layer0_outputs(1616)) or (layer0_outputs(5491));
    outputs(4471) <= (layer0_outputs(10331)) xor (layer0_outputs(210));
    outputs(4472) <= not(layer0_outputs(966));
    outputs(4473) <= not(layer0_outputs(2841));
    outputs(4474) <= not((layer0_outputs(2915)) xor (layer0_outputs(474)));
    outputs(4475) <= (layer0_outputs(1663)) and not (layer0_outputs(8387));
    outputs(4476) <= layer0_outputs(5146);
    outputs(4477) <= (layer0_outputs(10385)) and not (layer0_outputs(3076));
    outputs(4478) <= (layer0_outputs(8190)) xor (layer0_outputs(12628));
    outputs(4479) <= not((layer0_outputs(8703)) or (layer0_outputs(11757)));
    outputs(4480) <= not((layer0_outputs(11740)) xor (layer0_outputs(314)));
    outputs(4481) <= layer0_outputs(11110);
    outputs(4482) <= (layer0_outputs(3635)) and (layer0_outputs(9296));
    outputs(4483) <= (layer0_outputs(7332)) and not (layer0_outputs(9248));
    outputs(4484) <= layer0_outputs(7676);
    outputs(4485) <= (layer0_outputs(8085)) and not (layer0_outputs(6452));
    outputs(4486) <= not((layer0_outputs(12392)) xor (layer0_outputs(4469)));
    outputs(4487) <= layer0_outputs(8054);
    outputs(4488) <= not(layer0_outputs(11338)) or (layer0_outputs(10300));
    outputs(4489) <= not(layer0_outputs(4456));
    outputs(4490) <= (layer0_outputs(5508)) and (layer0_outputs(7315));
    outputs(4491) <= layer0_outputs(11606);
    outputs(4492) <= layer0_outputs(1353);
    outputs(4493) <= not((layer0_outputs(5499)) and (layer0_outputs(6590)));
    outputs(4494) <= not(layer0_outputs(6586)) or (layer0_outputs(10052));
    outputs(4495) <= not(layer0_outputs(582));
    outputs(4496) <= not(layer0_outputs(2552)) or (layer0_outputs(1478));
    outputs(4497) <= layer0_outputs(973);
    outputs(4498) <= not(layer0_outputs(4788));
    outputs(4499) <= layer0_outputs(8222);
    outputs(4500) <= not(layer0_outputs(5099));
    outputs(4501) <= (layer0_outputs(3845)) and (layer0_outputs(8534));
    outputs(4502) <= not((layer0_outputs(276)) and (layer0_outputs(6358)));
    outputs(4503) <= not(layer0_outputs(216)) or (layer0_outputs(8139));
    outputs(4504) <= not(layer0_outputs(2076));
    outputs(4505) <= not(layer0_outputs(10609));
    outputs(4506) <= not(layer0_outputs(98));
    outputs(4507) <= layer0_outputs(6569);
    outputs(4508) <= not(layer0_outputs(3018));
    outputs(4509) <= not((layer0_outputs(6652)) xor (layer0_outputs(7938)));
    outputs(4510) <= not((layer0_outputs(6642)) xor (layer0_outputs(7198)));
    outputs(4511) <= not(layer0_outputs(4180));
    outputs(4512) <= (layer0_outputs(7391)) and (layer0_outputs(8497));
    outputs(4513) <= not((layer0_outputs(6647)) and (layer0_outputs(12163)));
    outputs(4514) <= layer0_outputs(6231);
    outputs(4515) <= (layer0_outputs(12705)) xor (layer0_outputs(636));
    outputs(4516) <= (layer0_outputs(880)) xor (layer0_outputs(11901));
    outputs(4517) <= (layer0_outputs(9918)) xor (layer0_outputs(12518));
    outputs(4518) <= not(layer0_outputs(3074)) or (layer0_outputs(5285));
    outputs(4519) <= (layer0_outputs(8738)) and not (layer0_outputs(12283));
    outputs(4520) <= not(layer0_outputs(5684));
    outputs(4521) <= not(layer0_outputs(8022));
    outputs(4522) <= not(layer0_outputs(9520));
    outputs(4523) <= (layer0_outputs(7814)) xor (layer0_outputs(12778));
    outputs(4524) <= not((layer0_outputs(6108)) xor (layer0_outputs(11828)));
    outputs(4525) <= not(layer0_outputs(4357));
    outputs(4526) <= layer0_outputs(9319);
    outputs(4527) <= not((layer0_outputs(926)) or (layer0_outputs(9049)));
    outputs(4528) <= not(layer0_outputs(8436));
    outputs(4529) <= not(layer0_outputs(11953));
    outputs(4530) <= not((layer0_outputs(6430)) and (layer0_outputs(7210)));
    outputs(4531) <= not((layer0_outputs(1008)) xor (layer0_outputs(12321)));
    outputs(4532) <= (layer0_outputs(6659)) and not (layer0_outputs(10378));
    outputs(4533) <= not(layer0_outputs(6837));
    outputs(4534) <= not((layer0_outputs(6910)) xor (layer0_outputs(8058)));
    outputs(4535) <= not((layer0_outputs(4060)) and (layer0_outputs(1048)));
    outputs(4536) <= (layer0_outputs(2422)) xor (layer0_outputs(8286));
    outputs(4537) <= layer0_outputs(7583);
    outputs(4538) <= not(layer0_outputs(10667));
    outputs(4539) <= (layer0_outputs(12414)) xor (layer0_outputs(3282));
    outputs(4540) <= not((layer0_outputs(7532)) xor (layer0_outputs(7752)));
    outputs(4541) <= layer0_outputs(8461);
    outputs(4542) <= (layer0_outputs(11355)) and not (layer0_outputs(11478));
    outputs(4543) <= not((layer0_outputs(9660)) or (layer0_outputs(1684)));
    outputs(4544) <= (layer0_outputs(12775)) xor (layer0_outputs(12052));
    outputs(4545) <= not(layer0_outputs(4106));
    outputs(4546) <= (layer0_outputs(2189)) and not (layer0_outputs(6638));
    outputs(4547) <= not(layer0_outputs(9024));
    outputs(4548) <= (layer0_outputs(12043)) and not (layer0_outputs(7390));
    outputs(4549) <= not((layer0_outputs(7210)) xor (layer0_outputs(3154)));
    outputs(4550) <= layer0_outputs(453);
    outputs(4551) <= not((layer0_outputs(2918)) and (layer0_outputs(10343)));
    outputs(4552) <= not(layer0_outputs(5753));
    outputs(4553) <= not((layer0_outputs(4021)) xor (layer0_outputs(8147)));
    outputs(4554) <= not(layer0_outputs(364));
    outputs(4555) <= layer0_outputs(3900);
    outputs(4556) <= layer0_outputs(11044);
    outputs(4557) <= (layer0_outputs(3342)) and not (layer0_outputs(4395));
    outputs(4558) <= not((layer0_outputs(8202)) xor (layer0_outputs(7272)));
    outputs(4559) <= (layer0_outputs(3706)) and (layer0_outputs(10781));
    outputs(4560) <= (layer0_outputs(7779)) xor (layer0_outputs(1542));
    outputs(4561) <= not(layer0_outputs(5838)) or (layer0_outputs(5002));
    outputs(4562) <= layer0_outputs(1945);
    outputs(4563) <= (layer0_outputs(6745)) and not (layer0_outputs(5166));
    outputs(4564) <= (layer0_outputs(7485)) and not (layer0_outputs(10521));
    outputs(4565) <= (layer0_outputs(3699)) or (layer0_outputs(4844));
    outputs(4566) <= not(layer0_outputs(10883));
    outputs(4567) <= (layer0_outputs(3094)) xor (layer0_outputs(4110));
    outputs(4568) <= (layer0_outputs(7112)) and not (layer0_outputs(5162));
    outputs(4569) <= not(layer0_outputs(1302));
    outputs(4570) <= not((layer0_outputs(1473)) and (layer0_outputs(5953)));
    outputs(4571) <= not(layer0_outputs(1977));
    outputs(4572) <= layer0_outputs(6857);
    outputs(4573) <= not(layer0_outputs(7508));
    outputs(4574) <= (layer0_outputs(11300)) xor (layer0_outputs(4675));
    outputs(4575) <= not(layer0_outputs(1683));
    outputs(4576) <= not(layer0_outputs(9884)) or (layer0_outputs(4073));
    outputs(4577) <= not((layer0_outputs(10336)) xor (layer0_outputs(7833)));
    outputs(4578) <= (layer0_outputs(3801)) and not (layer0_outputs(10442));
    outputs(4579) <= (layer0_outputs(3755)) xor (layer0_outputs(725));
    outputs(4580) <= (layer0_outputs(6612)) and not (layer0_outputs(838));
    outputs(4581) <= not((layer0_outputs(4968)) or (layer0_outputs(10799)));
    outputs(4582) <= (layer0_outputs(327)) and (layer0_outputs(4417));
    outputs(4583) <= not(layer0_outputs(3273));
    outputs(4584) <= (layer0_outputs(8056)) and (layer0_outputs(11227));
    outputs(4585) <= not(layer0_outputs(401));
    outputs(4586) <= not((layer0_outputs(5028)) or (layer0_outputs(12735)));
    outputs(4587) <= (layer0_outputs(3754)) and not (layer0_outputs(1396));
    outputs(4588) <= layer0_outputs(3944);
    outputs(4589) <= not(layer0_outputs(1606));
    outputs(4590) <= (layer0_outputs(1214)) and not (layer0_outputs(2546));
    outputs(4591) <= (layer0_outputs(6859)) xor (layer0_outputs(3653));
    outputs(4592) <= layer0_outputs(9265);
    outputs(4593) <= not((layer0_outputs(3737)) xor (layer0_outputs(12375)));
    outputs(4594) <= not((layer0_outputs(10856)) xor (layer0_outputs(2382)));
    outputs(4595) <= not(layer0_outputs(5261));
    outputs(4596) <= (layer0_outputs(10115)) xor (layer0_outputs(1667));
    outputs(4597) <= layer0_outputs(9294);
    outputs(4598) <= (layer0_outputs(12424)) xor (layer0_outputs(1619));
    outputs(4599) <= (layer0_outputs(11158)) and not (layer0_outputs(10926));
    outputs(4600) <= (layer0_outputs(3973)) and (layer0_outputs(8845));
    outputs(4601) <= not((layer0_outputs(9666)) xor (layer0_outputs(4172)));
    outputs(4602) <= layer0_outputs(4863);
    outputs(4603) <= not((layer0_outputs(11275)) xor (layer0_outputs(12753)));
    outputs(4604) <= not(layer0_outputs(8364));
    outputs(4605) <= layer0_outputs(3858);
    outputs(4606) <= (layer0_outputs(7593)) and not (layer0_outputs(2230));
    outputs(4607) <= not(layer0_outputs(9679));
    outputs(4608) <= not(layer0_outputs(10762));
    outputs(4609) <= not((layer0_outputs(9607)) xor (layer0_outputs(1868)));
    outputs(4610) <= (layer0_outputs(12415)) xor (layer0_outputs(903));
    outputs(4611) <= (layer0_outputs(6846)) and (layer0_outputs(9373));
    outputs(4612) <= layer0_outputs(486);
    outputs(4613) <= not((layer0_outputs(4802)) or (layer0_outputs(1975)));
    outputs(4614) <= not(layer0_outputs(12653));
    outputs(4615) <= not(layer0_outputs(2106));
    outputs(4616) <= (layer0_outputs(9380)) xor (layer0_outputs(8368));
    outputs(4617) <= layer0_outputs(7774);
    outputs(4618) <= layer0_outputs(11050);
    outputs(4619) <= (layer0_outputs(6854)) and not (layer0_outputs(12324));
    outputs(4620) <= (layer0_outputs(8145)) xor (layer0_outputs(7537));
    outputs(4621) <= not((layer0_outputs(7007)) xor (layer0_outputs(4971)));
    outputs(4622) <= not(layer0_outputs(2314));
    outputs(4623) <= (layer0_outputs(362)) and not (layer0_outputs(562));
    outputs(4624) <= not((layer0_outputs(11428)) or (layer0_outputs(4529)));
    outputs(4625) <= layer0_outputs(10161);
    outputs(4626) <= layer0_outputs(10864);
    outputs(4627) <= not(layer0_outputs(421));
    outputs(4628) <= (layer0_outputs(8986)) or (layer0_outputs(6908));
    outputs(4629) <= not(layer0_outputs(4457)) or (layer0_outputs(12447));
    outputs(4630) <= (layer0_outputs(3859)) xor (layer0_outputs(720));
    outputs(4631) <= not(layer0_outputs(12162)) or (layer0_outputs(8682));
    outputs(4632) <= (layer0_outputs(2824)) and not (layer0_outputs(7748));
    outputs(4633) <= not(layer0_outputs(224));
    outputs(4634) <= not((layer0_outputs(8038)) and (layer0_outputs(3491)));
    outputs(4635) <= not((layer0_outputs(10867)) xor (layer0_outputs(2480)));
    outputs(4636) <= layer0_outputs(11654);
    outputs(4637) <= not((layer0_outputs(10389)) xor (layer0_outputs(2695)));
    outputs(4638) <= (layer0_outputs(5991)) or (layer0_outputs(632));
    outputs(4639) <= (layer0_outputs(11615)) xor (layer0_outputs(10263));
    outputs(4640) <= layer0_outputs(7505);
    outputs(4641) <= (layer0_outputs(9946)) and not (layer0_outputs(2497));
    outputs(4642) <= not((layer0_outputs(5804)) xor (layer0_outputs(10946)));
    outputs(4643) <= (layer0_outputs(2186)) and (layer0_outputs(1836));
    outputs(4644) <= not((layer0_outputs(4242)) xor (layer0_outputs(2327)));
    outputs(4645) <= (layer0_outputs(11858)) and (layer0_outputs(5336));
    outputs(4646) <= not((layer0_outputs(4549)) xor (layer0_outputs(2995)));
    outputs(4647) <= (layer0_outputs(10906)) or (layer0_outputs(6782));
    outputs(4648) <= layer0_outputs(5820);
    outputs(4649) <= (layer0_outputs(11659)) and (layer0_outputs(3610));
    outputs(4650) <= layer0_outputs(12141);
    outputs(4651) <= not((layer0_outputs(5306)) xor (layer0_outputs(9180)));
    outputs(4652) <= not(layer0_outputs(8634));
    outputs(4653) <= layer0_outputs(5542);
    outputs(4654) <= layer0_outputs(1128);
    outputs(4655) <= (layer0_outputs(2341)) xor (layer0_outputs(7022));
    outputs(4656) <= not(layer0_outputs(10228));
    outputs(4657) <= layer0_outputs(7299);
    outputs(4658) <= layer0_outputs(11329);
    outputs(4659) <= not(layer0_outputs(5170)) or (layer0_outputs(9543));
    outputs(4660) <= not(layer0_outputs(4887));
    outputs(4661) <= not(layer0_outputs(9706));
    outputs(4662) <= layer0_outputs(8028);
    outputs(4663) <= not(layer0_outputs(11890));
    outputs(4664) <= not((layer0_outputs(624)) xor (layer0_outputs(8158)));
    outputs(4665) <= not(layer0_outputs(5202));
    outputs(4666) <= not((layer0_outputs(7424)) xor (layer0_outputs(9701)));
    outputs(4667) <= not(layer0_outputs(9317));
    outputs(4668) <= not(layer0_outputs(141));
    outputs(4669) <= not(layer0_outputs(2407));
    outputs(4670) <= (layer0_outputs(11423)) xor (layer0_outputs(7189));
    outputs(4671) <= layer0_outputs(8767);
    outputs(4672) <= (layer0_outputs(4942)) xor (layer0_outputs(5441));
    outputs(4673) <= layer0_outputs(1828);
    outputs(4674) <= not(layer0_outputs(1507));
    outputs(4675) <= not((layer0_outputs(10876)) xor (layer0_outputs(10264)));
    outputs(4676) <= (layer0_outputs(6581)) and not (layer0_outputs(12615));
    outputs(4677) <= (layer0_outputs(8972)) and not (layer0_outputs(3332));
    outputs(4678) <= not(layer0_outputs(11592));
    outputs(4679) <= not((layer0_outputs(10284)) xor (layer0_outputs(9141)));
    outputs(4680) <= (layer0_outputs(11209)) and (layer0_outputs(8779));
    outputs(4681) <= layer0_outputs(12345);
    outputs(4682) <= (layer0_outputs(79)) and (layer0_outputs(148));
    outputs(4683) <= not(layer0_outputs(9268));
    outputs(4684) <= (layer0_outputs(6203)) and not (layer0_outputs(12535));
    outputs(4685) <= not((layer0_outputs(6500)) xor (layer0_outputs(3224)));
    outputs(4686) <= layer0_outputs(9236);
    outputs(4687) <= (layer0_outputs(6697)) and not (layer0_outputs(641));
    outputs(4688) <= layer0_outputs(2055);
    outputs(4689) <= not((layer0_outputs(2115)) xor (layer0_outputs(9025)));
    outputs(4690) <= not(layer0_outputs(1544));
    outputs(4691) <= not(layer0_outputs(849)) or (layer0_outputs(8659));
    outputs(4692) <= not(layer0_outputs(9994));
    outputs(4693) <= (layer0_outputs(1817)) and (layer0_outputs(9884));
    outputs(4694) <= not(layer0_outputs(7308));
    outputs(4695) <= not(layer0_outputs(7877));
    outputs(4696) <= not(layer0_outputs(4459)) or (layer0_outputs(8201));
    outputs(4697) <= (layer0_outputs(10468)) xor (layer0_outputs(3276));
    outputs(4698) <= (layer0_outputs(1113)) xor (layer0_outputs(6124));
    outputs(4699) <= (layer0_outputs(5446)) xor (layer0_outputs(7965));
    outputs(4700) <= not(layer0_outputs(5930));
    outputs(4701) <= not((layer0_outputs(1661)) or (layer0_outputs(2314)));
    outputs(4702) <= not((layer0_outputs(5211)) xor (layer0_outputs(11654)));
    outputs(4703) <= not(layer0_outputs(2819)) or (layer0_outputs(3747));
    outputs(4704) <= (layer0_outputs(11971)) and not (layer0_outputs(10425));
    outputs(4705) <= (layer0_outputs(1070)) xor (layer0_outputs(8499));
    outputs(4706) <= not((layer0_outputs(5403)) and (layer0_outputs(8707)));
    outputs(4707) <= layer0_outputs(8177);
    outputs(4708) <= not((layer0_outputs(7905)) and (layer0_outputs(8408)));
    outputs(4709) <= (layer0_outputs(369)) and (layer0_outputs(3121));
    outputs(4710) <= not(layer0_outputs(8554)) or (layer0_outputs(4556));
    outputs(4711) <= (layer0_outputs(2037)) and (layer0_outputs(1643));
    outputs(4712) <= layer0_outputs(4777);
    outputs(4713) <= not(layer0_outputs(8842));
    outputs(4714) <= (layer0_outputs(7012)) xor (layer0_outputs(5470));
    outputs(4715) <= layer0_outputs(10051);
    outputs(4716) <= (layer0_outputs(3355)) or (layer0_outputs(8905));
    outputs(4717) <= (layer0_outputs(4491)) and not (layer0_outputs(2431));
    outputs(4718) <= (layer0_outputs(12269)) and not (layer0_outputs(3506));
    outputs(4719) <= not(layer0_outputs(2352));
    outputs(4720) <= not(layer0_outputs(8279));
    outputs(4721) <= not((layer0_outputs(12761)) and (layer0_outputs(1949)));
    outputs(4722) <= layer0_outputs(9539);
    outputs(4723) <= not(layer0_outputs(596));
    outputs(4724) <= not((layer0_outputs(10784)) xor (layer0_outputs(6375)));
    outputs(4725) <= (layer0_outputs(8479)) xor (layer0_outputs(5687));
    outputs(4726) <= not((layer0_outputs(9376)) xor (layer0_outputs(5214)));
    outputs(4727) <= (layer0_outputs(10554)) or (layer0_outputs(9670));
    outputs(4728) <= not((layer0_outputs(9139)) or (layer0_outputs(648)));
    outputs(4729) <= (layer0_outputs(8794)) and (layer0_outputs(11885));
    outputs(4730) <= layer0_outputs(9290);
    outputs(4731) <= not(layer0_outputs(11282));
    outputs(4732) <= (layer0_outputs(1893)) or (layer0_outputs(783));
    outputs(4733) <= not(layer0_outputs(1269));
    outputs(4734) <= (layer0_outputs(1752)) xor (layer0_outputs(3389));
    outputs(4735) <= layer0_outputs(6991);
    outputs(4736) <= not(layer0_outputs(2959));
    outputs(4737) <= not((layer0_outputs(135)) and (layer0_outputs(7600)));
    outputs(4738) <= (layer0_outputs(185)) xor (layer0_outputs(9791));
    outputs(4739) <= not((layer0_outputs(6737)) xor (layer0_outputs(2914)));
    outputs(4740) <= not(layer0_outputs(8053));
    outputs(4741) <= (layer0_outputs(6695)) and not (layer0_outputs(8754));
    outputs(4742) <= not(layer0_outputs(8082));
    outputs(4743) <= (layer0_outputs(9507)) xor (layer0_outputs(10622));
    outputs(4744) <= not(layer0_outputs(4136));
    outputs(4745) <= not(layer0_outputs(3934));
    outputs(4746) <= (layer0_outputs(2564)) xor (layer0_outputs(602));
    outputs(4747) <= layer0_outputs(3061);
    outputs(4748) <= (layer0_outputs(11593)) and (layer0_outputs(12757));
    outputs(4749) <= (layer0_outputs(1679)) xor (layer0_outputs(6576));
    outputs(4750) <= (layer0_outputs(3408)) and (layer0_outputs(4640));
    outputs(4751) <= not(layer0_outputs(10705)) or (layer0_outputs(11750));
    outputs(4752) <= (layer0_outputs(7817)) and not (layer0_outputs(12420));
    outputs(4753) <= not(layer0_outputs(7558));
    outputs(4754) <= (layer0_outputs(7576)) xor (layer0_outputs(3228));
    outputs(4755) <= not((layer0_outputs(11147)) xor (layer0_outputs(2068)));
    outputs(4756) <= layer0_outputs(12295);
    outputs(4757) <= (layer0_outputs(7515)) and not (layer0_outputs(5290));
    outputs(4758) <= not(layer0_outputs(10446));
    outputs(4759) <= (layer0_outputs(829)) xor (layer0_outputs(2311));
    outputs(4760) <= layer0_outputs(502);
    outputs(4761) <= layer0_outputs(5117);
    outputs(4762) <= not(layer0_outputs(764)) or (layer0_outputs(4015));
    outputs(4763) <= not((layer0_outputs(11256)) xor (layer0_outputs(4762)));
    outputs(4764) <= not(layer0_outputs(12621));
    outputs(4765) <= (layer0_outputs(5866)) xor (layer0_outputs(1983));
    outputs(4766) <= layer0_outputs(8378);
    outputs(4767) <= layer0_outputs(8700);
    outputs(4768) <= layer0_outputs(1336);
    outputs(4769) <= not(layer0_outputs(9039));
    outputs(4770) <= (layer0_outputs(11487)) and not (layer0_outputs(311));
    outputs(4771) <= not(layer0_outputs(3631));
    outputs(4772) <= not(layer0_outputs(3289)) or (layer0_outputs(9064));
    outputs(4773) <= (layer0_outputs(5993)) and (layer0_outputs(2551));
    outputs(4774) <= not(layer0_outputs(7426));
    outputs(4775) <= not(layer0_outputs(11953));
    outputs(4776) <= layer0_outputs(12751);
    outputs(4777) <= not(layer0_outputs(10290));
    outputs(4778) <= not((layer0_outputs(5405)) xor (layer0_outputs(11987)));
    outputs(4779) <= not((layer0_outputs(7951)) xor (layer0_outputs(8080)));
    outputs(4780) <= (layer0_outputs(12531)) and not (layer0_outputs(7046));
    outputs(4781) <= layer0_outputs(9554);
    outputs(4782) <= not((layer0_outputs(2720)) xor (layer0_outputs(5888)));
    outputs(4783) <= layer0_outputs(11980);
    outputs(4784) <= not(layer0_outputs(8670)) or (layer0_outputs(11765));
    outputs(4785) <= not(layer0_outputs(5621));
    outputs(4786) <= not(layer0_outputs(3117));
    outputs(4787) <= layer0_outputs(4981);
    outputs(4788) <= not(layer0_outputs(10285));
    outputs(4789) <= (layer0_outputs(9481)) and (layer0_outputs(7301));
    outputs(4790) <= not(layer0_outputs(4630)) or (layer0_outputs(2308));
    outputs(4791) <= not(layer0_outputs(3517));
    outputs(4792) <= not(layer0_outputs(7083));
    outputs(4793) <= (layer0_outputs(2510)) or (layer0_outputs(7144));
    outputs(4794) <= not(layer0_outputs(4570));
    outputs(4795) <= not(layer0_outputs(9184)) or (layer0_outputs(1324));
    outputs(4796) <= (layer0_outputs(6854)) or (layer0_outputs(12130));
    outputs(4797) <= not(layer0_outputs(3686));
    outputs(4798) <= layer0_outputs(419);
    outputs(4799) <= (layer0_outputs(1122)) and not (layer0_outputs(9869));
    outputs(4800) <= layer0_outputs(10200);
    outputs(4801) <= not((layer0_outputs(3264)) and (layer0_outputs(4307)));
    outputs(4802) <= not(layer0_outputs(9317));
    outputs(4803) <= (layer0_outputs(11445)) xor (layer0_outputs(1463));
    outputs(4804) <= not((layer0_outputs(451)) or (layer0_outputs(10204)));
    outputs(4805) <= (layer0_outputs(3424)) xor (layer0_outputs(6002));
    outputs(4806) <= not(layer0_outputs(1660));
    outputs(4807) <= (layer0_outputs(4080)) xor (layer0_outputs(6684));
    outputs(4808) <= not((layer0_outputs(3016)) xor (layer0_outputs(2789)));
    outputs(4809) <= not(layer0_outputs(5607)) or (layer0_outputs(2692));
    outputs(4810) <= layer0_outputs(3532);
    outputs(4811) <= (layer0_outputs(2785)) xor (layer0_outputs(3475));
    outputs(4812) <= not(layer0_outputs(2005)) or (layer0_outputs(3991));
    outputs(4813) <= not(layer0_outputs(2435));
    outputs(4814) <= not(layer0_outputs(2790)) or (layer0_outputs(3266));
    outputs(4815) <= (layer0_outputs(10983)) xor (layer0_outputs(1810));
    outputs(4816) <= not(layer0_outputs(912));
    outputs(4817) <= not(layer0_outputs(1907));
    outputs(4818) <= not(layer0_outputs(2398));
    outputs(4819) <= not(layer0_outputs(8920));
    outputs(4820) <= not((layer0_outputs(8434)) xor (layer0_outputs(5152)));
    outputs(4821) <= (layer0_outputs(8025)) or (layer0_outputs(7504));
    outputs(4822) <= layer0_outputs(8600);
    outputs(4823) <= layer0_outputs(1779);
    outputs(4824) <= not((layer0_outputs(10029)) xor (layer0_outputs(9410)));
    outputs(4825) <= not((layer0_outputs(7187)) xor (layer0_outputs(1286)));
    outputs(4826) <= not(layer0_outputs(9856)) or (layer0_outputs(1095));
    outputs(4827) <= layer0_outputs(7051);
    outputs(4828) <= not((layer0_outputs(6579)) and (layer0_outputs(9235)));
    outputs(4829) <= layer0_outputs(8614);
    outputs(4830) <= (layer0_outputs(1083)) and not (layer0_outputs(9631));
    outputs(4831) <= layer0_outputs(7894);
    outputs(4832) <= not((layer0_outputs(8006)) and (layer0_outputs(2854)));
    outputs(4833) <= (layer0_outputs(2343)) and not (layer0_outputs(4738));
    outputs(4834) <= layer0_outputs(2754);
    outputs(4835) <= layer0_outputs(4961);
    outputs(4836) <= not(layer0_outputs(10454));
    outputs(4837) <= not(layer0_outputs(4223)) or (layer0_outputs(7876));
    outputs(4838) <= not(layer0_outputs(7173));
    outputs(4839) <= (layer0_outputs(12672)) and not (layer0_outputs(3163));
    outputs(4840) <= (layer0_outputs(8302)) and not (layer0_outputs(5988));
    outputs(4841) <= layer0_outputs(8086);
    outputs(4842) <= (layer0_outputs(8859)) and (layer0_outputs(10075));
    outputs(4843) <= (layer0_outputs(10574)) xor (layer0_outputs(5897));
    outputs(4844) <= (layer0_outputs(8017)) and not (layer0_outputs(1091));
    outputs(4845) <= layer0_outputs(4108);
    outputs(4846) <= not((layer0_outputs(2594)) xor (layer0_outputs(10956)));
    outputs(4847) <= not(layer0_outputs(10680));
    outputs(4848) <= layer0_outputs(11589);
    outputs(4849) <= (layer0_outputs(2268)) xor (layer0_outputs(11461));
    outputs(4850) <= not((layer0_outputs(11318)) xor (layer0_outputs(10865)));
    outputs(4851) <= not(layer0_outputs(7726));
    outputs(4852) <= not(layer0_outputs(8204));
    outputs(4853) <= not((layer0_outputs(7099)) xor (layer0_outputs(6954)));
    outputs(4854) <= not((layer0_outputs(8886)) xor (layer0_outputs(8985)));
    outputs(4855) <= not((layer0_outputs(8699)) or (layer0_outputs(672)));
    outputs(4856) <= layer0_outputs(161);
    outputs(4857) <= (layer0_outputs(2870)) and not (layer0_outputs(4932));
    outputs(4858) <= layer0_outputs(12147);
    outputs(4859) <= not(layer0_outputs(4487));
    outputs(4860) <= not(layer0_outputs(8173));
    outputs(4861) <= (layer0_outputs(10787)) xor (layer0_outputs(2356));
    outputs(4862) <= (layer0_outputs(3172)) xor (layer0_outputs(11961));
    outputs(4863) <= layer0_outputs(8124);
    outputs(4864) <= (layer0_outputs(5853)) or (layer0_outputs(5200));
    outputs(4865) <= not((layer0_outputs(11483)) and (layer0_outputs(5792)));
    outputs(4866) <= (layer0_outputs(5375)) and not (layer0_outputs(3820));
    outputs(4867) <= not(layer0_outputs(8478)) or (layer0_outputs(7607));
    outputs(4868) <= (layer0_outputs(7794)) and not (layer0_outputs(607));
    outputs(4869) <= layer0_outputs(2592);
    outputs(4870) <= (layer0_outputs(840)) and (layer0_outputs(10886));
    outputs(4871) <= not((layer0_outputs(10655)) xor (layer0_outputs(5895)));
    outputs(4872) <= layer0_outputs(10748);
    outputs(4873) <= not((layer0_outputs(10592)) xor (layer0_outputs(3650)));
    outputs(4874) <= not((layer0_outputs(3155)) xor (layer0_outputs(10014)));
    outputs(4875) <= not(layer0_outputs(9639));
    outputs(4876) <= (layer0_outputs(1829)) xor (layer0_outputs(6462));
    outputs(4877) <= not(layer0_outputs(4364));
    outputs(4878) <= layer0_outputs(10542);
    outputs(4879) <= layer0_outputs(3342);
    outputs(4880) <= not((layer0_outputs(12581)) xor (layer0_outputs(2156)));
    outputs(4881) <= not(layer0_outputs(5515));
    outputs(4882) <= layer0_outputs(1782);
    outputs(4883) <= (layer0_outputs(3108)) xor (layer0_outputs(4298));
    outputs(4884) <= (layer0_outputs(3121)) or (layer0_outputs(4079));
    outputs(4885) <= (layer0_outputs(2231)) xor (layer0_outputs(10438));
    outputs(4886) <= not(layer0_outputs(4729));
    outputs(4887) <= not(layer0_outputs(8219));
    outputs(4888) <= not((layer0_outputs(9288)) xor (layer0_outputs(9320)));
    outputs(4889) <= not(layer0_outputs(2838));
    outputs(4890) <= layer0_outputs(11735);
    outputs(4891) <= not((layer0_outputs(11060)) xor (layer0_outputs(12134)));
    outputs(4892) <= not((layer0_outputs(803)) xor (layer0_outputs(9308)));
    outputs(4893) <= not(layer0_outputs(5160));
    outputs(4894) <= (layer0_outputs(9806)) xor (layer0_outputs(4629));
    outputs(4895) <= not((layer0_outputs(878)) xor (layer0_outputs(9417)));
    outputs(4896) <= not((layer0_outputs(534)) xor (layer0_outputs(6066)));
    outputs(4897) <= (layer0_outputs(5681)) or (layer0_outputs(637));
    outputs(4898) <= not((layer0_outputs(8101)) xor (layer0_outputs(3812)));
    outputs(4899) <= not(layer0_outputs(2934));
    outputs(4900) <= (layer0_outputs(2359)) xor (layer0_outputs(1090));
    outputs(4901) <= not((layer0_outputs(2414)) xor (layer0_outputs(1157)));
    outputs(4902) <= (layer0_outputs(1559)) xor (layer0_outputs(10288));
    outputs(4903) <= not(layer0_outputs(196)) or (layer0_outputs(688));
    outputs(4904) <= not(layer0_outputs(3655));
    outputs(4905) <= (layer0_outputs(8489)) and (layer0_outputs(1151));
    outputs(4906) <= '1';
    outputs(4907) <= (layer0_outputs(10548)) xor (layer0_outputs(8766));
    outputs(4908) <= not((layer0_outputs(11499)) xor (layer0_outputs(7140)));
    outputs(4909) <= not(layer0_outputs(3101));
    outputs(4910) <= (layer0_outputs(11728)) and not (layer0_outputs(9640));
    outputs(4911) <= (layer0_outputs(5723)) and not (layer0_outputs(11632));
    outputs(4912) <= not((layer0_outputs(10765)) or (layer0_outputs(3767)));
    outputs(4913) <= not(layer0_outputs(5845));
    outputs(4914) <= (layer0_outputs(4479)) and (layer0_outputs(8437));
    outputs(4915) <= not(layer0_outputs(10544));
    outputs(4916) <= layer0_outputs(4225);
    outputs(4917) <= not(layer0_outputs(5851));
    outputs(4918) <= (layer0_outputs(10189)) and not (layer0_outputs(12315));
    outputs(4919) <= not(layer0_outputs(1047)) or (layer0_outputs(3586));
    outputs(4920) <= layer0_outputs(59);
    outputs(4921) <= not((layer0_outputs(7196)) xor (layer0_outputs(6721)));
    outputs(4922) <= not((layer0_outputs(2416)) xor (layer0_outputs(5163)));
    outputs(4923) <= layer0_outputs(2252);
    outputs(4924) <= not(layer0_outputs(11416));
    outputs(4925) <= (layer0_outputs(12091)) and (layer0_outputs(7008));
    outputs(4926) <= not((layer0_outputs(1085)) and (layer0_outputs(5650)));
    outputs(4927) <= (layer0_outputs(3047)) xor (layer0_outputs(1677));
    outputs(4928) <= (layer0_outputs(11038)) and not (layer0_outputs(9496));
    outputs(4929) <= layer0_outputs(2532);
    outputs(4930) <= not((layer0_outputs(7822)) xor (layer0_outputs(4485)));
    outputs(4931) <= not(layer0_outputs(2894)) or (layer0_outputs(12300));
    outputs(4932) <= (layer0_outputs(10520)) xor (layer0_outputs(7243));
    outputs(4933) <= (layer0_outputs(9138)) xor (layer0_outputs(3057));
    outputs(4934) <= (layer0_outputs(4917)) or (layer0_outputs(2043));
    outputs(4935) <= not(layer0_outputs(10024)) or (layer0_outputs(6654));
    outputs(4936) <= (layer0_outputs(4741)) xor (layer0_outputs(12780));
    outputs(4937) <= not(layer0_outputs(9077));
    outputs(4938) <= not((layer0_outputs(6945)) or (layer0_outputs(10232)));
    outputs(4939) <= layer0_outputs(10058);
    outputs(4940) <= not((layer0_outputs(6704)) xor (layer0_outputs(913)));
    outputs(4941) <= (layer0_outputs(5418)) xor (layer0_outputs(7314));
    outputs(4942) <= not((layer0_outputs(991)) xor (layer0_outputs(1990)));
    outputs(4943) <= (layer0_outputs(12687)) xor (layer0_outputs(11235));
    outputs(4944) <= (layer0_outputs(12572)) and (layer0_outputs(5453));
    outputs(4945) <= (layer0_outputs(5893)) xor (layer0_outputs(4637));
    outputs(4946) <= layer0_outputs(4501);
    outputs(4947) <= (layer0_outputs(12364)) xor (layer0_outputs(8433));
    outputs(4948) <= not((layer0_outputs(8951)) or (layer0_outputs(4559)));
    outputs(4949) <= layer0_outputs(8422);
    outputs(4950) <= not((layer0_outputs(2918)) xor (layer0_outputs(5559)));
    outputs(4951) <= (layer0_outputs(10029)) xor (layer0_outputs(2936));
    outputs(4952) <= (layer0_outputs(11280)) xor (layer0_outputs(11434));
    outputs(4953) <= layer0_outputs(2607);
    outputs(4954) <= not((layer0_outputs(8414)) or (layer0_outputs(2569)));
    outputs(4955) <= not(layer0_outputs(3336));
    outputs(4956) <= (layer0_outputs(3958)) xor (layer0_outputs(23));
    outputs(4957) <= (layer0_outputs(7084)) and not (layer0_outputs(3328));
    outputs(4958) <= (layer0_outputs(12177)) and not (layer0_outputs(4475));
    outputs(4959) <= (layer0_outputs(12087)) xor (layer0_outputs(4561));
    outputs(4960) <= layer0_outputs(4739);
    outputs(4961) <= layer0_outputs(5708);
    outputs(4962) <= layer0_outputs(1882);
    outputs(4963) <= not((layer0_outputs(8188)) xor (layer0_outputs(7730)));
    outputs(4964) <= (layer0_outputs(12164)) xor (layer0_outputs(8832));
    outputs(4965) <= not((layer0_outputs(2542)) xor (layer0_outputs(1790)));
    outputs(4966) <= layer0_outputs(9234);
    outputs(4967) <= not((layer0_outputs(5172)) xor (layer0_outputs(5640)));
    outputs(4968) <= not((layer0_outputs(757)) and (layer0_outputs(10243)));
    outputs(4969) <= (layer0_outputs(12627)) and (layer0_outputs(574));
    outputs(4970) <= layer0_outputs(11971);
    outputs(4971) <= layer0_outputs(4117);
    outputs(4972) <= (layer0_outputs(8774)) and not (layer0_outputs(8068));
    outputs(4973) <= not(layer0_outputs(1632)) or (layer0_outputs(4700));
    outputs(4974) <= (layer0_outputs(5509)) xor (layer0_outputs(5406));
    outputs(4975) <= not(layer0_outputs(10485));
    outputs(4976) <= layer0_outputs(5661);
    outputs(4977) <= (layer0_outputs(11893)) xor (layer0_outputs(2367));
    outputs(4978) <= not(layer0_outputs(11457)) or (layer0_outputs(6063));
    outputs(4979) <= not(layer0_outputs(10329)) or (layer0_outputs(2973));
    outputs(4980) <= layer0_outputs(5587);
    outputs(4981) <= not(layer0_outputs(6109));
    outputs(4982) <= (layer0_outputs(9291)) xor (layer0_outputs(12254));
    outputs(4983) <= (layer0_outputs(9197)) xor (layer0_outputs(3458));
    outputs(4984) <= (layer0_outputs(1462)) and (layer0_outputs(3917));
    outputs(4985) <= layer0_outputs(7259);
    outputs(4986) <= not(layer0_outputs(5059));
    outputs(4987) <= not(layer0_outputs(3705));
    outputs(4988) <= not(layer0_outputs(1412));
    outputs(4989) <= layer0_outputs(10789);
    outputs(4990) <= not(layer0_outputs(8952)) or (layer0_outputs(9001));
    outputs(4991) <= (layer0_outputs(5789)) and not (layer0_outputs(8270));
    outputs(4992) <= layer0_outputs(7651);
    outputs(4993) <= not((layer0_outputs(7488)) xor (layer0_outputs(6543)));
    outputs(4994) <= not(layer0_outputs(2641));
    outputs(4995) <= (layer0_outputs(10511)) and not (layer0_outputs(6975));
    outputs(4996) <= not(layer0_outputs(617));
    outputs(4997) <= layer0_outputs(5856);
    outputs(4998) <= (layer0_outputs(10889)) and not (layer0_outputs(5456));
    outputs(4999) <= layer0_outputs(6168);
    outputs(5000) <= not((layer0_outputs(712)) xor (layer0_outputs(12148)));
    outputs(5001) <= not(layer0_outputs(8861)) or (layer0_outputs(2979));
    outputs(5002) <= layer0_outputs(782);
    outputs(5003) <= not(layer0_outputs(171));
    outputs(5004) <= layer0_outputs(3819);
    outputs(5005) <= not(layer0_outputs(8128)) or (layer0_outputs(796));
    outputs(5006) <= not(layer0_outputs(5296));
    outputs(5007) <= (layer0_outputs(1201)) or (layer0_outputs(367));
    outputs(5008) <= not((layer0_outputs(2917)) xor (layer0_outputs(11684)));
    outputs(5009) <= not((layer0_outputs(4698)) xor (layer0_outputs(3302)));
    outputs(5010) <= (layer0_outputs(11681)) xor (layer0_outputs(2622));
    outputs(5011) <= layer0_outputs(4265);
    outputs(5012) <= layer0_outputs(6069);
    outputs(5013) <= layer0_outputs(1052);
    outputs(5014) <= layer0_outputs(1837);
    outputs(5015) <= not(layer0_outputs(3053));
    outputs(5016) <= not(layer0_outputs(11313));
    outputs(5017) <= (layer0_outputs(2182)) xor (layer0_outputs(4590));
    outputs(5018) <= not(layer0_outputs(10561)) or (layer0_outputs(12061));
    outputs(5019) <= not(layer0_outputs(6698)) or (layer0_outputs(5864));
    outputs(5020) <= not((layer0_outputs(7254)) xor (layer0_outputs(1525)));
    outputs(5021) <= not(layer0_outputs(8954));
    outputs(5022) <= not((layer0_outputs(2499)) or (layer0_outputs(5196)));
    outputs(5023) <= not((layer0_outputs(638)) xor (layer0_outputs(1152)));
    outputs(5024) <= layer0_outputs(8562);
    outputs(5025) <= layer0_outputs(502);
    outputs(5026) <= not(layer0_outputs(11150));
    outputs(5027) <= layer0_outputs(6760);
    outputs(5028) <= layer0_outputs(1212);
    outputs(5029) <= not(layer0_outputs(11568));
    outputs(5030) <= (layer0_outputs(6475)) xor (layer0_outputs(3935));
    outputs(5031) <= not(layer0_outputs(12754));
    outputs(5032) <= not(layer0_outputs(4036));
    outputs(5033) <= (layer0_outputs(8158)) xor (layer0_outputs(4950));
    outputs(5034) <= not(layer0_outputs(1911)) or (layer0_outputs(6440));
    outputs(5035) <= not(layer0_outputs(10581)) or (layer0_outputs(12345));
    outputs(5036) <= not(layer0_outputs(7436)) or (layer0_outputs(11535));
    outputs(5037) <= layer0_outputs(9340);
    outputs(5038) <= (layer0_outputs(2409)) and (layer0_outputs(8080));
    outputs(5039) <= not((layer0_outputs(2645)) or (layer0_outputs(10466)));
    outputs(5040) <= layer0_outputs(5633);
    outputs(5041) <= not((layer0_outputs(8591)) or (layer0_outputs(1734)));
    outputs(5042) <= layer0_outputs(11033);
    outputs(5043) <= layer0_outputs(5728);
    outputs(5044) <= not(layer0_outputs(11084));
    outputs(5045) <= layer0_outputs(7728);
    outputs(5046) <= layer0_outputs(10821);
    outputs(5047) <= not(layer0_outputs(3955));
    outputs(5048) <= (layer0_outputs(2908)) or (layer0_outputs(250));
    outputs(5049) <= layer0_outputs(1133);
    outputs(5050) <= (layer0_outputs(10510)) and (layer0_outputs(1621));
    outputs(5051) <= layer0_outputs(12295);
    outputs(5052) <= not((layer0_outputs(908)) xor (layer0_outputs(5852)));
    outputs(5053) <= layer0_outputs(12430);
    outputs(5054) <= layer0_outputs(1099);
    outputs(5055) <= not(layer0_outputs(10917));
    outputs(5056) <= (layer0_outputs(445)) xor (layer0_outputs(5635));
    outputs(5057) <= not(layer0_outputs(7264));
    outputs(5058) <= layer0_outputs(11851);
    outputs(5059) <= (layer0_outputs(8579)) xor (layer0_outputs(11457));
    outputs(5060) <= not(layer0_outputs(9112)) or (layer0_outputs(3709));
    outputs(5061) <= not(layer0_outputs(9002));
    outputs(5062) <= not(layer0_outputs(7246));
    outputs(5063) <= (layer0_outputs(1222)) xor (layer0_outputs(11919));
    outputs(5064) <= not((layer0_outputs(4900)) xor (layer0_outputs(3759)));
    outputs(5065) <= not(layer0_outputs(11274));
    outputs(5066) <= not((layer0_outputs(767)) xor (layer0_outputs(1851)));
    outputs(5067) <= not((layer0_outputs(1631)) xor (layer0_outputs(2988)));
    outputs(5068) <= (layer0_outputs(8007)) xor (layer0_outputs(5140));
    outputs(5069) <= not((layer0_outputs(7796)) xor (layer0_outputs(4184)));
    outputs(5070) <= not(layer0_outputs(6363));
    outputs(5071) <= (layer0_outputs(3581)) xor (layer0_outputs(8680));
    outputs(5072) <= not(layer0_outputs(1321));
    outputs(5073) <= not((layer0_outputs(6519)) xor (layer0_outputs(2254)));
    outputs(5074) <= layer0_outputs(10781);
    outputs(5075) <= (layer0_outputs(11560)) xor (layer0_outputs(4438));
    outputs(5076) <= (layer0_outputs(5064)) and (layer0_outputs(10104));
    outputs(5077) <= (layer0_outputs(515)) xor (layer0_outputs(6322));
    outputs(5078) <= not((layer0_outputs(10594)) or (layer0_outputs(5523)));
    outputs(5079) <= (layer0_outputs(2451)) xor (layer0_outputs(6797));
    outputs(5080) <= (layer0_outputs(3518)) xor (layer0_outputs(9452));
    outputs(5081) <= not(layer0_outputs(6682));
    outputs(5082) <= (layer0_outputs(11854)) xor (layer0_outputs(8377));
    outputs(5083) <= not((layer0_outputs(1712)) xor (layer0_outputs(9895)));
    outputs(5084) <= layer0_outputs(3107);
    outputs(5085) <= not(layer0_outputs(3432));
    outputs(5086) <= (layer0_outputs(8518)) and not (layer0_outputs(11610));
    outputs(5087) <= not(layer0_outputs(11984));
    outputs(5088) <= layer0_outputs(3058);
    outputs(5089) <= not((layer0_outputs(1732)) xor (layer0_outputs(6635)));
    outputs(5090) <= layer0_outputs(1326);
    outputs(5091) <= layer0_outputs(1180);
    outputs(5092) <= not(layer0_outputs(2386));
    outputs(5093) <= layer0_outputs(7330);
    outputs(5094) <= (layer0_outputs(1609)) xor (layer0_outputs(7017));
    outputs(5095) <= layer0_outputs(1554);
    outputs(5096) <= layer0_outputs(9753);
    outputs(5097) <= (layer0_outputs(6976)) and not (layer0_outputs(3101));
    outputs(5098) <= (layer0_outputs(2118)) xor (layer0_outputs(11386));
    outputs(5099) <= not((layer0_outputs(5060)) and (layer0_outputs(4462)));
    outputs(5100) <= layer0_outputs(914);
    outputs(5101) <= (layer0_outputs(6629)) and not (layer0_outputs(9145));
    outputs(5102) <= not(layer0_outputs(1235));
    outputs(5103) <= not(layer0_outputs(766)) or (layer0_outputs(5808));
    outputs(5104) <= (layer0_outputs(3083)) and not (layer0_outputs(3093));
    outputs(5105) <= not(layer0_outputs(6514));
    outputs(5106) <= not(layer0_outputs(3331)) or (layer0_outputs(11455));
    outputs(5107) <= (layer0_outputs(7972)) and not (layer0_outputs(3779));
    outputs(5108) <= not(layer0_outputs(9937));
    outputs(5109) <= not(layer0_outputs(6906));
    outputs(5110) <= (layer0_outputs(394)) xor (layer0_outputs(6677));
    outputs(5111) <= (layer0_outputs(11040)) and not (layer0_outputs(7100));
    outputs(5112) <= not((layer0_outputs(6373)) xor (layer0_outputs(10291)));
    outputs(5113) <= not(layer0_outputs(9731));
    outputs(5114) <= layer0_outputs(12340);
    outputs(5115) <= (layer0_outputs(5222)) xor (layer0_outputs(3949));
    outputs(5116) <= layer0_outputs(7613);
    outputs(5117) <= not((layer0_outputs(3463)) xor (layer0_outputs(2525)));
    outputs(5118) <= not(layer0_outputs(5712));
    outputs(5119) <= not(layer0_outputs(3450));
    outputs(5120) <= not(layer0_outputs(4953)) or (layer0_outputs(2475));
    outputs(5121) <= (layer0_outputs(7306)) xor (layer0_outputs(3830));
    outputs(5122) <= layer0_outputs(3751);
    outputs(5123) <= (layer0_outputs(9563)) and (layer0_outputs(11653));
    outputs(5124) <= not(layer0_outputs(9375));
    outputs(5125) <= not((layer0_outputs(8596)) xor (layer0_outputs(664)));
    outputs(5126) <= not(layer0_outputs(581));
    outputs(5127) <= (layer0_outputs(5138)) and (layer0_outputs(9040));
    outputs(5128) <= not((layer0_outputs(10316)) xor (layer0_outputs(8734)));
    outputs(5129) <= (layer0_outputs(4141)) and (layer0_outputs(8909));
    outputs(5130) <= not((layer0_outputs(8107)) xor (layer0_outputs(9213)));
    outputs(5131) <= not((layer0_outputs(59)) xor (layer0_outputs(6636)));
    outputs(5132) <= (layer0_outputs(3000)) xor (layer0_outputs(3363));
    outputs(5133) <= layer0_outputs(861);
    outputs(5134) <= (layer0_outputs(12250)) xor (layer0_outputs(4488));
    outputs(5135) <= layer0_outputs(12224);
    outputs(5136) <= (layer0_outputs(2399)) and not (layer0_outputs(12363));
    outputs(5137) <= layer0_outputs(3458);
    outputs(5138) <= not(layer0_outputs(7842));
    outputs(5139) <= (layer0_outputs(2084)) xor (layer0_outputs(10755));
    outputs(5140) <= not(layer0_outputs(6090));
    outputs(5141) <= not(layer0_outputs(3359));
    outputs(5142) <= (layer0_outputs(9671)) xor (layer0_outputs(3913));
    outputs(5143) <= layer0_outputs(10361);
    outputs(5144) <= (layer0_outputs(560)) and not (layer0_outputs(6241));
    outputs(5145) <= layer0_outputs(12045);
    outputs(5146) <= not((layer0_outputs(4282)) xor (layer0_outputs(553)));
    outputs(5147) <= (layer0_outputs(7592)) and (layer0_outputs(8042));
    outputs(5148) <= not(layer0_outputs(10806)) or (layer0_outputs(315));
    outputs(5149) <= layer0_outputs(41);
    outputs(5150) <= not((layer0_outputs(498)) and (layer0_outputs(3723)));
    outputs(5151) <= not(layer0_outputs(10360));
    outputs(5152) <= (layer0_outputs(2969)) xor (layer0_outputs(5560));
    outputs(5153) <= not((layer0_outputs(1766)) xor (layer0_outputs(10042)));
    outputs(5154) <= (layer0_outputs(9732)) xor (layer0_outputs(11055));
    outputs(5155) <= (layer0_outputs(7825)) and not (layer0_outputs(6542));
    outputs(5156) <= layer0_outputs(5799);
    outputs(5157) <= not(layer0_outputs(6151));
    outputs(5158) <= not(layer0_outputs(3628));
    outputs(5159) <= not((layer0_outputs(4026)) or (layer0_outputs(8620)));
    outputs(5160) <= (layer0_outputs(1064)) xor (layer0_outputs(1072));
    outputs(5161) <= not((layer0_outputs(5009)) or (layer0_outputs(1197)));
    outputs(5162) <= not(layer0_outputs(3384));
    outputs(5163) <= layer0_outputs(8850);
    outputs(5164) <= (layer0_outputs(22)) xor (layer0_outputs(7125));
    outputs(5165) <= not(layer0_outputs(10384));
    outputs(5166) <= (layer0_outputs(11711)) xor (layer0_outputs(10812));
    outputs(5167) <= not(layer0_outputs(6969));
    outputs(5168) <= (layer0_outputs(8210)) xor (layer0_outputs(8076));
    outputs(5169) <= (layer0_outputs(5253)) xor (layer0_outputs(12533));
    outputs(5170) <= layer0_outputs(9994);
    outputs(5171) <= (layer0_outputs(3170)) and not (layer0_outputs(8047));
    outputs(5172) <= layer0_outputs(8395);
    outputs(5173) <= not(layer0_outputs(9663));
    outputs(5174) <= not(layer0_outputs(12337));
    outputs(5175) <= not((layer0_outputs(11100)) xor (layer0_outputs(8031)));
    outputs(5176) <= (layer0_outputs(9948)) and not (layer0_outputs(12168));
    outputs(5177) <= not(layer0_outputs(10327));
    outputs(5178) <= not((layer0_outputs(1988)) or (layer0_outputs(10597)));
    outputs(5179) <= layer0_outputs(1376);
    outputs(5180) <= layer0_outputs(2843);
    outputs(5181) <= not((layer0_outputs(4474)) xor (layer0_outputs(3433)));
    outputs(5182) <= not(layer0_outputs(4966)) or (layer0_outputs(885));
    outputs(5183) <= (layer0_outputs(1655)) and not (layer0_outputs(1407));
    outputs(5184) <= (layer0_outputs(8836)) xor (layer0_outputs(8384));
    outputs(5185) <= (layer0_outputs(10198)) and not (layer0_outputs(1329));
    outputs(5186) <= not((layer0_outputs(3237)) xor (layer0_outputs(6668)));
    outputs(5187) <= not(layer0_outputs(3144));
    outputs(5188) <= not(layer0_outputs(7567));
    outputs(5189) <= not((layer0_outputs(2877)) xor (layer0_outputs(1645)));
    outputs(5190) <= not(layer0_outputs(5896));
    outputs(5191) <= layer0_outputs(9922);
    outputs(5192) <= (layer0_outputs(970)) xor (layer0_outputs(2191));
    outputs(5193) <= layer0_outputs(3378);
    outputs(5194) <= layer0_outputs(7880);
    outputs(5195) <= not((layer0_outputs(3089)) xor (layer0_outputs(3880)));
    outputs(5196) <= not((layer0_outputs(8191)) xor (layer0_outputs(6503)));
    outputs(5197) <= (layer0_outputs(855)) or (layer0_outputs(9867));
    outputs(5198) <= layer0_outputs(5098);
    outputs(5199) <= not((layer0_outputs(8547)) and (layer0_outputs(9705)));
    outputs(5200) <= (layer0_outputs(8022)) xor (layer0_outputs(5041));
    outputs(5201) <= (layer0_outputs(7490)) and (layer0_outputs(3391));
    outputs(5202) <= not((layer0_outputs(3212)) xor (layer0_outputs(9148)));
    outputs(5203) <= (layer0_outputs(9567)) and not (layer0_outputs(10112));
    outputs(5204) <= not(layer0_outputs(651));
    outputs(5205) <= not((layer0_outputs(7561)) xor (layer0_outputs(8031)));
    outputs(5206) <= (layer0_outputs(10505)) and not (layer0_outputs(6487));
    outputs(5207) <= not((layer0_outputs(5534)) xor (layer0_outputs(11702)));
    outputs(5208) <= not((layer0_outputs(2805)) xor (layer0_outputs(10242)));
    outputs(5209) <= not(layer0_outputs(4851));
    outputs(5210) <= (layer0_outputs(5144)) or (layer0_outputs(5273));
    outputs(5211) <= layer0_outputs(3757);
    outputs(5212) <= (layer0_outputs(7939)) xor (layer0_outputs(7752));
    outputs(5213) <= not((layer0_outputs(10100)) xor (layer0_outputs(2512)));
    outputs(5214) <= (layer0_outputs(10549)) xor (layer0_outputs(2254));
    outputs(5215) <= (layer0_outputs(11327)) and (layer0_outputs(11039));
    outputs(5216) <= (layer0_outputs(3535)) xor (layer0_outputs(9592));
    outputs(5217) <= not((layer0_outputs(6213)) and (layer0_outputs(2035)));
    outputs(5218) <= not((layer0_outputs(12135)) xor (layer0_outputs(4678)));
    outputs(5219) <= not((layer0_outputs(3423)) or (layer0_outputs(4598)));
    outputs(5220) <= (layer0_outputs(4435)) xor (layer0_outputs(5940));
    outputs(5221) <= (layer0_outputs(8247)) and not (layer0_outputs(11820));
    outputs(5222) <= layer0_outputs(1308);
    outputs(5223) <= not((layer0_outputs(71)) xor (layer0_outputs(5714)));
    outputs(5224) <= not((layer0_outputs(9081)) xor (layer0_outputs(2991)));
    outputs(5225) <= not(layer0_outputs(2728));
    outputs(5226) <= layer0_outputs(6472);
    outputs(5227) <= (layer0_outputs(3120)) or (layer0_outputs(10187));
    outputs(5228) <= layer0_outputs(11419);
    outputs(5229) <= not(layer0_outputs(1517));
    outputs(5230) <= not(layer0_outputs(9368));
    outputs(5231) <= not((layer0_outputs(6452)) xor (layer0_outputs(7834)));
    outputs(5232) <= (layer0_outputs(8690)) or (layer0_outputs(5419));
    outputs(5233) <= not(layer0_outputs(10474));
    outputs(5234) <= not((layer0_outputs(4110)) or (layer0_outputs(3783)));
    outputs(5235) <= layer0_outputs(12308);
    outputs(5236) <= not((layer0_outputs(7176)) xor (layer0_outputs(2164)));
    outputs(5237) <= (layer0_outputs(5601)) xor (layer0_outputs(10091));
    outputs(5238) <= layer0_outputs(4752);
    outputs(5239) <= layer0_outputs(8962);
    outputs(5240) <= (layer0_outputs(10946)) xor (layer0_outputs(6347));
    outputs(5241) <= (layer0_outputs(11745)) and not (layer0_outputs(9565));
    outputs(5242) <= not(layer0_outputs(1432));
    outputs(5243) <= (layer0_outputs(7744)) xor (layer0_outputs(2741));
    outputs(5244) <= (layer0_outputs(8521)) or (layer0_outputs(11107));
    outputs(5245) <= layer0_outputs(5274);
    outputs(5246) <= (layer0_outputs(7373)) xor (layer0_outputs(5585));
    outputs(5247) <= not((layer0_outputs(11933)) or (layer0_outputs(2256)));
    outputs(5248) <= not(layer0_outputs(896)) or (layer0_outputs(8795));
    outputs(5249) <= not(layer0_outputs(5359));
    outputs(5250) <= not(layer0_outputs(2453));
    outputs(5251) <= (layer0_outputs(10578)) and (layer0_outputs(3303));
    outputs(5252) <= (layer0_outputs(3691)) xor (layer0_outputs(6400));
    outputs(5253) <= layer0_outputs(10072);
    outputs(5254) <= (layer0_outputs(7647)) xor (layer0_outputs(3560));
    outputs(5255) <= not(layer0_outputs(6375));
    outputs(5256) <= not((layer0_outputs(12186)) and (layer0_outputs(10631)));
    outputs(5257) <= not((layer0_outputs(5105)) or (layer0_outputs(7005)));
    outputs(5258) <= (layer0_outputs(361)) or (layer0_outputs(12051));
    outputs(5259) <= not(layer0_outputs(921));
    outputs(5260) <= layer0_outputs(2269);
    outputs(5261) <= (layer0_outputs(10869)) xor (layer0_outputs(4432));
    outputs(5262) <= (layer0_outputs(8098)) and not (layer0_outputs(12718));
    outputs(5263) <= (layer0_outputs(3689)) xor (layer0_outputs(10366));
    outputs(5264) <= (layer0_outputs(5756)) or (layer0_outputs(11664));
    outputs(5265) <= layer0_outputs(8611);
    outputs(5266) <= layer0_outputs(12322);
    outputs(5267) <= layer0_outputs(12309);
    outputs(5268) <= not(layer0_outputs(4151));
    outputs(5269) <= not((layer0_outputs(114)) and (layer0_outputs(269)));
    outputs(5270) <= not(layer0_outputs(8569));
    outputs(5271) <= (layer0_outputs(4429)) and not (layer0_outputs(6582));
    outputs(5272) <= (layer0_outputs(4650)) and (layer0_outputs(7044));
    outputs(5273) <= not(layer0_outputs(5160));
    outputs(5274) <= not(layer0_outputs(400));
    outputs(5275) <= not((layer0_outputs(7526)) xor (layer0_outputs(2483)));
    outputs(5276) <= (layer0_outputs(238)) and not (layer0_outputs(8677));
    outputs(5277) <= (layer0_outputs(3755)) and (layer0_outputs(4335));
    outputs(5278) <= (layer0_outputs(11638)) and (layer0_outputs(10043));
    outputs(5279) <= not((layer0_outputs(4191)) xor (layer0_outputs(3452)));
    outputs(5280) <= layer0_outputs(1545);
    outputs(5281) <= not((layer0_outputs(9383)) and (layer0_outputs(206)));
    outputs(5282) <= not(layer0_outputs(5779));
    outputs(5283) <= layer0_outputs(2611);
    outputs(5284) <= not(layer0_outputs(8183)) or (layer0_outputs(6938));
    outputs(5285) <= not(layer0_outputs(9224));
    outputs(5286) <= not(layer0_outputs(7876));
    outputs(5287) <= not(layer0_outputs(217));
    outputs(5288) <= layer0_outputs(3293);
    outputs(5289) <= (layer0_outputs(4530)) and (layer0_outputs(5469));
    outputs(5290) <= (layer0_outputs(674)) and not (layer0_outputs(7844));
    outputs(5291) <= not(layer0_outputs(10847));
    outputs(5292) <= not((layer0_outputs(9176)) or (layer0_outputs(7179)));
    outputs(5293) <= not(layer0_outputs(201));
    outputs(5294) <= (layer0_outputs(10423)) or (layer0_outputs(130));
    outputs(5295) <= not(layer0_outputs(1018));
    outputs(5296) <= (layer0_outputs(5306)) xor (layer0_outputs(8116));
    outputs(5297) <= layer0_outputs(1471);
    outputs(5298) <= not(layer0_outputs(11293));
    outputs(5299) <= not(layer0_outputs(145));
    outputs(5300) <= not((layer0_outputs(8211)) or (layer0_outputs(11385)));
    outputs(5301) <= not(layer0_outputs(9231));
    outputs(5302) <= (layer0_outputs(8776)) xor (layer0_outputs(4661));
    outputs(5303) <= not((layer0_outputs(3227)) or (layer0_outputs(11065)));
    outputs(5304) <= layer0_outputs(8941);
    outputs(5305) <= (layer0_outputs(9523)) and not (layer0_outputs(6985));
    outputs(5306) <= (layer0_outputs(1401)) or (layer0_outputs(7002));
    outputs(5307) <= (layer0_outputs(12218)) xor (layer0_outputs(8514));
    outputs(5308) <= not(layer0_outputs(9155));
    outputs(5309) <= layer0_outputs(1739);
    outputs(5310) <= not((layer0_outputs(7206)) xor (layer0_outputs(11317)));
    outputs(5311) <= layer0_outputs(9821);
    outputs(5312) <= not(layer0_outputs(12601));
    outputs(5313) <= (layer0_outputs(5525)) xor (layer0_outputs(4254));
    outputs(5314) <= (layer0_outputs(4504)) and not (layer0_outputs(3526));
    outputs(5315) <= not(layer0_outputs(4653));
    outputs(5316) <= (layer0_outputs(318)) xor (layer0_outputs(12698));
    outputs(5317) <= not((layer0_outputs(3309)) xor (layer0_outputs(3084)));
    outputs(5318) <= not((layer0_outputs(2153)) xor (layer0_outputs(9381)));
    outputs(5319) <= not(layer0_outputs(4879));
    outputs(5320) <= (layer0_outputs(3460)) xor (layer0_outputs(11408));
    outputs(5321) <= layer0_outputs(1954);
    outputs(5322) <= layer0_outputs(2475);
    outputs(5323) <= not((layer0_outputs(11498)) or (layer0_outputs(9544)));
    outputs(5324) <= not((layer0_outputs(6086)) xor (layer0_outputs(3991)));
    outputs(5325) <= (layer0_outputs(5807)) and not (layer0_outputs(6836));
    outputs(5326) <= not((layer0_outputs(10708)) or (layer0_outputs(9356)));
    outputs(5327) <= (layer0_outputs(4444)) xor (layer0_outputs(8306));
    outputs(5328) <= not((layer0_outputs(2338)) and (layer0_outputs(10885)));
    outputs(5329) <= not((layer0_outputs(9353)) or (layer0_outputs(3754)));
    outputs(5330) <= not(layer0_outputs(2058));
    outputs(5331) <= layer0_outputs(287);
    outputs(5332) <= (layer0_outputs(1575)) and (layer0_outputs(10730));
    outputs(5333) <= not((layer0_outputs(10122)) xor (layer0_outputs(4291)));
    outputs(5334) <= not(layer0_outputs(2579));
    outputs(5335) <= (layer0_outputs(566)) and not (layer0_outputs(8418));
    outputs(5336) <= not(layer0_outputs(2749));
    outputs(5337) <= not(layer0_outputs(11694));
    outputs(5338) <= layer0_outputs(1969);
    outputs(5339) <= layer0_outputs(2732);
    outputs(5340) <= layer0_outputs(8791);
    outputs(5341) <= not(layer0_outputs(407)) or (layer0_outputs(5113));
    outputs(5342) <= not(layer0_outputs(9713));
    outputs(5343) <= not(layer0_outputs(769)) or (layer0_outputs(8906));
    outputs(5344) <= layer0_outputs(10691);
    outputs(5345) <= not((layer0_outputs(5363)) and (layer0_outputs(11095)));
    outputs(5346) <= not((layer0_outputs(4622)) xor (layer0_outputs(5793)));
    outputs(5347) <= not(layer0_outputs(11532));
    outputs(5348) <= not(layer0_outputs(904));
    outputs(5349) <= not((layer0_outputs(2337)) xor (layer0_outputs(3883)));
    outputs(5350) <= not((layer0_outputs(8067)) xor (layer0_outputs(9698)));
    outputs(5351) <= (layer0_outputs(978)) xor (layer0_outputs(8152));
    outputs(5352) <= not((layer0_outputs(6679)) xor (layer0_outputs(1033)));
    outputs(5353) <= not(layer0_outputs(4417));
    outputs(5354) <= not((layer0_outputs(9464)) xor (layer0_outputs(5548)));
    outputs(5355) <= not((layer0_outputs(12457)) or (layer0_outputs(10512)));
    outputs(5356) <= layer0_outputs(89);
    outputs(5357) <= not(layer0_outputs(525));
    outputs(5358) <= not(layer0_outputs(4111));
    outputs(5359) <= not(layer0_outputs(3673));
    outputs(5360) <= not((layer0_outputs(5699)) xor (layer0_outputs(3764)));
    outputs(5361) <= (layer0_outputs(8405)) xor (layer0_outputs(3538));
    outputs(5362) <= (layer0_outputs(2030)) xor (layer0_outputs(5957));
    outputs(5363) <= layer0_outputs(3172);
    outputs(5364) <= not(layer0_outputs(5345));
    outputs(5365) <= not((layer0_outputs(1818)) and (layer0_outputs(7011)));
    outputs(5366) <= not(layer0_outputs(5422)) or (layer0_outputs(2901));
    outputs(5367) <= not(layer0_outputs(11491));
    outputs(5368) <= not(layer0_outputs(3645));
    outputs(5369) <= (layer0_outputs(3354)) and not (layer0_outputs(4290));
    outputs(5370) <= not(layer0_outputs(6591));
    outputs(5371) <= not((layer0_outputs(835)) xor (layer0_outputs(4831)));
    outputs(5372) <= layer0_outputs(12182);
    outputs(5373) <= not((layer0_outputs(5085)) and (layer0_outputs(11663)));
    outputs(5374) <= layer0_outputs(4064);
    outputs(5375) <= not(layer0_outputs(1728));
    outputs(5376) <= not((layer0_outputs(3331)) xor (layer0_outputs(9069)));
    outputs(5377) <= layer0_outputs(6230);
    outputs(5378) <= (layer0_outputs(2855)) xor (layer0_outputs(241));
    outputs(5379) <= not(layer0_outputs(1858));
    outputs(5380) <= not((layer0_outputs(12251)) and (layer0_outputs(12371)));
    outputs(5381) <= (layer0_outputs(180)) xor (layer0_outputs(7480));
    outputs(5382) <= not(layer0_outputs(6860));
    outputs(5383) <= (layer0_outputs(10003)) xor (layer0_outputs(3745));
    outputs(5384) <= not((layer0_outputs(9565)) xor (layer0_outputs(10705)));
    outputs(5385) <= not((layer0_outputs(10060)) xor (layer0_outputs(11608)));
    outputs(5386) <= not((layer0_outputs(2282)) xor (layer0_outputs(3721)));
    outputs(5387) <= (layer0_outputs(4713)) or (layer0_outputs(4167));
    outputs(5388) <= not((layer0_outputs(4119)) xor (layer0_outputs(5218)));
    outputs(5389) <= not((layer0_outputs(487)) or (layer0_outputs(11266)));
    outputs(5390) <= not((layer0_outputs(3366)) xor (layer0_outputs(11375)));
    outputs(5391) <= layer0_outputs(1528);
    outputs(5392) <= (layer0_outputs(11239)) and not (layer0_outputs(11677));
    outputs(5393) <= not((layer0_outputs(5427)) xor (layer0_outputs(257)));
    outputs(5394) <= (layer0_outputs(10903)) and not (layer0_outputs(5805));
    outputs(5395) <= (layer0_outputs(7870)) and (layer0_outputs(4718));
    outputs(5396) <= not((layer0_outputs(972)) xor (layer0_outputs(9300)));
    outputs(5397) <= not((layer0_outputs(4500)) and (layer0_outputs(4309)));
    outputs(5398) <= layer0_outputs(2907);
    outputs(5399) <= (layer0_outputs(8186)) and (layer0_outputs(5850));
    outputs(5400) <= (layer0_outputs(3063)) xor (layer0_outputs(5660));
    outputs(5401) <= (layer0_outputs(4331)) xor (layer0_outputs(11083));
    outputs(5402) <= layer0_outputs(1308);
    outputs(5403) <= layer0_outputs(3629);
    outputs(5404) <= layer0_outputs(6781);
    outputs(5405) <= (layer0_outputs(9527)) and (layer0_outputs(10048));
    outputs(5406) <= not(layer0_outputs(1323));
    outputs(5407) <= (layer0_outputs(6572)) and not (layer0_outputs(244));
    outputs(5408) <= (layer0_outputs(3891)) and not (layer0_outputs(11707));
    outputs(5409) <= not((layer0_outputs(11938)) xor (layer0_outputs(7588)));
    outputs(5410) <= not((layer0_outputs(12481)) or (layer0_outputs(4004)));
    outputs(5411) <= layer0_outputs(999);
    outputs(5412) <= not(layer0_outputs(4044));
    outputs(5413) <= not(layer0_outputs(10494));
    outputs(5414) <= (layer0_outputs(434)) xor (layer0_outputs(2379));
    outputs(5415) <= not(layer0_outputs(4439));
    outputs(5416) <= layer0_outputs(2134);
    outputs(5417) <= not((layer0_outputs(7117)) xor (layer0_outputs(4717)));
    outputs(5418) <= (layer0_outputs(2752)) or (layer0_outputs(5523));
    outputs(5419) <= not((layer0_outputs(5445)) and (layer0_outputs(1410)));
    outputs(5420) <= (layer0_outputs(11459)) and not (layer0_outputs(2676));
    outputs(5421) <= layer0_outputs(10014);
    outputs(5422) <= (layer0_outputs(11001)) xor (layer0_outputs(5578));
    outputs(5423) <= not((layer0_outputs(9905)) xor (layer0_outputs(1103)));
    outputs(5424) <= (layer0_outputs(876)) xor (layer0_outputs(11533));
    outputs(5425) <= (layer0_outputs(7994)) xor (layer0_outputs(1933));
    outputs(5426) <= (layer0_outputs(6393)) xor (layer0_outputs(12792));
    outputs(5427) <= not(layer0_outputs(1362));
    outputs(5428) <= (layer0_outputs(9316)) and not (layer0_outputs(8289));
    outputs(5429) <= (layer0_outputs(8234)) and not (layer0_outputs(8344));
    outputs(5430) <= layer0_outputs(4607);
    outputs(5431) <= layer0_outputs(11244);
    outputs(5432) <= layer0_outputs(11489);
    outputs(5433) <= not(layer0_outputs(7977));
    outputs(5434) <= not(layer0_outputs(6304));
    outputs(5435) <= not((layer0_outputs(9102)) or (layer0_outputs(11383)));
    outputs(5436) <= (layer0_outputs(8922)) xor (layer0_outputs(10063));
    outputs(5437) <= (layer0_outputs(7151)) and (layer0_outputs(2551));
    outputs(5438) <= layer0_outputs(12599);
    outputs(5439) <= not(layer0_outputs(3358));
    outputs(5440) <= (layer0_outputs(10923)) xor (layer0_outputs(436));
    outputs(5441) <= not(layer0_outputs(1496));
    outputs(5442) <= not((layer0_outputs(3393)) and (layer0_outputs(6870)));
    outputs(5443) <= not((layer0_outputs(1101)) xor (layer0_outputs(10032)));
    outputs(5444) <= layer0_outputs(8819);
    outputs(5445) <= (layer0_outputs(7662)) xor (layer0_outputs(12494));
    outputs(5446) <= layer0_outputs(12616);
    outputs(5447) <= (layer0_outputs(12543)) and not (layer0_outputs(1182));
    outputs(5448) <= not((layer0_outputs(396)) or (layer0_outputs(6656)));
    outputs(5449) <= not(layer0_outputs(6243));
    outputs(5450) <= layer0_outputs(2039);
    outputs(5451) <= not(layer0_outputs(2501));
    outputs(5452) <= (layer0_outputs(1705)) xor (layer0_outputs(10127));
    outputs(5453) <= layer0_outputs(10928);
    outputs(5454) <= (layer0_outputs(6717)) xor (layer0_outputs(336));
    outputs(5455) <= (layer0_outputs(2999)) and not (layer0_outputs(4512));
    outputs(5456) <= layer0_outputs(5322);
    outputs(5457) <= layer0_outputs(176);
    outputs(5458) <= not(layer0_outputs(6939));
    outputs(5459) <= layer0_outputs(11800);
    outputs(5460) <= layer0_outputs(6536);
    outputs(5461) <= not(layer0_outputs(11034));
    outputs(5462) <= not((layer0_outputs(8107)) xor (layer0_outputs(4533)));
    outputs(5463) <= layer0_outputs(9331);
    outputs(5464) <= layer0_outputs(4341);
    outputs(5465) <= not((layer0_outputs(6523)) xor (layer0_outputs(357)));
    outputs(5466) <= (layer0_outputs(10440)) and not (layer0_outputs(2627));
    outputs(5467) <= not(layer0_outputs(8229));
    outputs(5468) <= layer0_outputs(12007);
    outputs(5469) <= not((layer0_outputs(476)) xor (layer0_outputs(2309)));
    outputs(5470) <= layer0_outputs(3596);
    outputs(5471) <= not((layer0_outputs(3049)) xor (layer0_outputs(4098)));
    outputs(5472) <= not((layer0_outputs(7721)) and (layer0_outputs(9968)));
    outputs(5473) <= not((layer0_outputs(665)) xor (layer0_outputs(833)));
    outputs(5474) <= (layer0_outputs(10743)) and not (layer0_outputs(12168));
    outputs(5475) <= layer0_outputs(10362);
    outputs(5476) <= not(layer0_outputs(6528));
    outputs(5477) <= (layer0_outputs(10251)) and (layer0_outputs(7749));
    outputs(5478) <= not((layer0_outputs(1796)) xor (layer0_outputs(8787)));
    outputs(5479) <= not(layer0_outputs(7142));
    outputs(5480) <= layer0_outputs(7880);
    outputs(5481) <= layer0_outputs(1630);
    outputs(5482) <= not(layer0_outputs(4528));
    outputs(5483) <= layer0_outputs(762);
    outputs(5484) <= (layer0_outputs(7815)) and (layer0_outputs(6558));
    outputs(5485) <= (layer0_outputs(9104)) or (layer0_outputs(12511));
    outputs(5486) <= not(layer0_outputs(4406));
    outputs(5487) <= (layer0_outputs(11948)) and not (layer0_outputs(4385));
    outputs(5488) <= (layer0_outputs(7260)) xor (layer0_outputs(12173));
    outputs(5489) <= (layer0_outputs(3750)) xor (layer0_outputs(11271));
    outputs(5490) <= layer0_outputs(2336);
    outputs(5491) <= not(layer0_outputs(7318));
    outputs(5492) <= layer0_outputs(4850);
    outputs(5493) <= (layer0_outputs(7507)) xor (layer0_outputs(1195));
    outputs(5494) <= not((layer0_outputs(11956)) or (layer0_outputs(1859)));
    outputs(5495) <= not(layer0_outputs(11017));
    outputs(5496) <= layer0_outputs(6102);
    outputs(5497) <= not((layer0_outputs(7930)) and (layer0_outputs(9898)));
    outputs(5498) <= not(layer0_outputs(12626));
    outputs(5499) <= not(layer0_outputs(72));
    outputs(5500) <= layer0_outputs(11447);
    outputs(5501) <= (layer0_outputs(11754)) and not (layer0_outputs(12479));
    outputs(5502) <= layer0_outputs(2106);
    outputs(5503) <= not(layer0_outputs(5569));
    outputs(5504) <= layer0_outputs(1730);
    outputs(5505) <= (layer0_outputs(5952)) xor (layer0_outputs(5840));
    outputs(5506) <= not((layer0_outputs(10857)) xor (layer0_outputs(4922)));
    outputs(5507) <= (layer0_outputs(2093)) xor (layer0_outputs(3597));
    outputs(5508) <= not(layer0_outputs(1352));
    outputs(5509) <= not((layer0_outputs(7341)) xor (layer0_outputs(2753)));
    outputs(5510) <= not(layer0_outputs(9950));
    outputs(5511) <= layer0_outputs(1298);
    outputs(5512) <= layer0_outputs(10647);
    outputs(5513) <= layer0_outputs(4380);
    outputs(5514) <= (layer0_outputs(1637)) xor (layer0_outputs(7523));
    outputs(5515) <= (layer0_outputs(2635)) and (layer0_outputs(818));
    outputs(5516) <= layer0_outputs(7807);
    outputs(5517) <= (layer0_outputs(6288)) and not (layer0_outputs(6980));
    outputs(5518) <= not((layer0_outputs(7287)) or (layer0_outputs(7718)));
    outputs(5519) <= (layer0_outputs(12631)) xor (layer0_outputs(6283));
    outputs(5520) <= not(layer0_outputs(8788)) or (layer0_outputs(7351));
    outputs(5521) <= not((layer0_outputs(11366)) and (layer0_outputs(5631)));
    outputs(5522) <= layer0_outputs(7152);
    outputs(5523) <= not((layer0_outputs(6749)) xor (layer0_outputs(1925)));
    outputs(5524) <= (layer0_outputs(7802)) xor (layer0_outputs(4215));
    outputs(5525) <= (layer0_outputs(1120)) xor (layer0_outputs(2543));
    outputs(5526) <= (layer0_outputs(3017)) and not (layer0_outputs(2796));
    outputs(5527) <= layer0_outputs(8100);
    outputs(5528) <= not(layer0_outputs(10220));
    outputs(5529) <= not((layer0_outputs(9028)) xor (layer0_outputs(10704)));
    outputs(5530) <= (layer0_outputs(1565)) and not (layer0_outputs(6660));
    outputs(5531) <= not(layer0_outputs(11896));
    outputs(5532) <= not(layer0_outputs(5909));
    outputs(5533) <= not(layer0_outputs(3612));
    outputs(5534) <= (layer0_outputs(8757)) and (layer0_outputs(9532));
    outputs(5535) <= not(layer0_outputs(3479));
    outputs(5536) <= (layer0_outputs(11288)) xor (layer0_outputs(11103));
    outputs(5537) <= layer0_outputs(6403);
    outputs(5538) <= not((layer0_outputs(12600)) xor (layer0_outputs(5855)));
    outputs(5539) <= not(layer0_outputs(8753));
    outputs(5540) <= not(layer0_outputs(9710));
    outputs(5541) <= not((layer0_outputs(2670)) and (layer0_outputs(11614)));
    outputs(5542) <= (layer0_outputs(4982)) and not (layer0_outputs(2976));
    outputs(5543) <= layer0_outputs(9314);
    outputs(5544) <= (layer0_outputs(8116)) or (layer0_outputs(9470));
    outputs(5545) <= not(layer0_outputs(5713));
    outputs(5546) <= not(layer0_outputs(5521));
    outputs(5547) <= layer0_outputs(541);
    outputs(5548) <= (layer0_outputs(5074)) and (layer0_outputs(11833));
    outputs(5549) <= not((layer0_outputs(10804)) xor (layer0_outputs(11814)));
    outputs(5550) <= not(layer0_outputs(11630));
    outputs(5551) <= (layer0_outputs(5811)) and not (layer0_outputs(8865));
    outputs(5552) <= not(layer0_outputs(4512));
    outputs(5553) <= not(layer0_outputs(11764));
    outputs(5554) <= not(layer0_outputs(7602));
    outputs(5555) <= not((layer0_outputs(9083)) xor (layer0_outputs(7001)));
    outputs(5556) <= not((layer0_outputs(10463)) xor (layer0_outputs(3503)));
    outputs(5557) <= not(layer0_outputs(3658)) or (layer0_outputs(8012));
    outputs(5558) <= not((layer0_outputs(9914)) or (layer0_outputs(4889)));
    outputs(5559) <= not(layer0_outputs(4681)) or (layer0_outputs(1589));
    outputs(5560) <= (layer0_outputs(6354)) xor (layer0_outputs(1452));
    outputs(5561) <= (layer0_outputs(830)) xor (layer0_outputs(6582));
    outputs(5562) <= not(layer0_outputs(282));
    outputs(5563) <= layer0_outputs(1468);
    outputs(5564) <= (layer0_outputs(10304)) xor (layer0_outputs(4040));
    outputs(5565) <= layer0_outputs(7570);
    outputs(5566) <= (layer0_outputs(8976)) xor (layer0_outputs(12630));
    outputs(5567) <= not((layer0_outputs(12651)) xor (layer0_outputs(10658)));
    outputs(5568) <= not((layer0_outputs(2020)) or (layer0_outputs(537)));
    outputs(5569) <= not(layer0_outputs(2108));
    outputs(5570) <= not(layer0_outputs(5002));
    outputs(5571) <= not((layer0_outputs(10148)) or (layer0_outputs(8101)));
    outputs(5572) <= layer0_outputs(3899);
    outputs(5573) <= (layer0_outputs(7043)) xor (layer0_outputs(4326));
    outputs(5574) <= (layer0_outputs(5187)) and (layer0_outputs(11099));
    outputs(5575) <= layer0_outputs(10559);
    outputs(5576) <= not(layer0_outputs(6799));
    outputs(5577) <= layer0_outputs(12680);
    outputs(5578) <= not((layer0_outputs(8355)) xor (layer0_outputs(4226)));
    outputs(5579) <= (layer0_outputs(9307)) xor (layer0_outputs(10012));
    outputs(5580) <= layer0_outputs(12482);
    outputs(5581) <= (layer0_outputs(7144)) xor (layer0_outputs(11350));
    outputs(5582) <= not((layer0_outputs(11845)) or (layer0_outputs(4275)));
    outputs(5583) <= not(layer0_outputs(2258));
    outputs(5584) <= (layer0_outputs(5391)) xor (layer0_outputs(5656));
    outputs(5585) <= not((layer0_outputs(5868)) or (layer0_outputs(814)));
    outputs(5586) <= not((layer0_outputs(12350)) or (layer0_outputs(1943)));
    outputs(5587) <= not(layer0_outputs(2324));
    outputs(5588) <= layer0_outputs(5082);
    outputs(5589) <= layer0_outputs(4065);
    outputs(5590) <= not((layer0_outputs(11115)) xor (layer0_outputs(5729)));
    outputs(5591) <= not(layer0_outputs(5141));
    outputs(5592) <= layer0_outputs(10095);
    outputs(5593) <= layer0_outputs(1185);
    outputs(5594) <= (layer0_outputs(4190)) xor (layer0_outputs(8040));
    outputs(5595) <= layer0_outputs(9445);
    outputs(5596) <= not((layer0_outputs(11)) or (layer0_outputs(9264)));
    outputs(5597) <= layer0_outputs(6704);
    outputs(5598) <= not(layer0_outputs(5139));
    outputs(5599) <= not(layer0_outputs(10553));
    outputs(5600) <= not((layer0_outputs(5907)) xor (layer0_outputs(11944)));
    outputs(5601) <= not((layer0_outputs(2415)) or (layer0_outputs(2082)));
    outputs(5602) <= (layer0_outputs(12099)) and not (layer0_outputs(10397));
    outputs(5603) <= not((layer0_outputs(12538)) xor (layer0_outputs(8786)));
    outputs(5604) <= not((layer0_outputs(1554)) xor (layer0_outputs(3188)));
    outputs(5605) <= (layer0_outputs(735)) and not (layer0_outputs(6019));
    outputs(5606) <= not((layer0_outputs(12037)) xor (layer0_outputs(4801)));
    outputs(5607) <= (layer0_outputs(10624)) xor (layer0_outputs(2422));
    outputs(5608) <= not((layer0_outputs(323)) xor (layer0_outputs(7861)));
    outputs(5609) <= not((layer0_outputs(5469)) xor (layer0_outputs(3114)));
    outputs(5610) <= (layer0_outputs(4741)) and (layer0_outputs(288));
    outputs(5611) <= not(layer0_outputs(440));
    outputs(5612) <= not(layer0_outputs(12729));
    outputs(5613) <= (layer0_outputs(9805)) and not (layer0_outputs(12110));
    outputs(5614) <= layer0_outputs(9643);
    outputs(5615) <= (layer0_outputs(327)) or (layer0_outputs(3710));
    outputs(5616) <= layer0_outputs(9939);
    outputs(5617) <= (layer0_outputs(5269)) and not (layer0_outputs(4547));
    outputs(5618) <= not(layer0_outputs(5056));
    outputs(5619) <= not(layer0_outputs(8919));
    outputs(5620) <= layer0_outputs(4674);
    outputs(5621) <= not((layer0_outputs(9500)) xor (layer0_outputs(10839)));
    outputs(5622) <= not((layer0_outputs(7134)) or (layer0_outputs(11094)));
    outputs(5623) <= (layer0_outputs(9595)) or (layer0_outputs(6552));
    outputs(5624) <= not(layer0_outputs(12594));
    outputs(5625) <= not(layer0_outputs(11427));
    outputs(5626) <= not((layer0_outputs(11463)) and (layer0_outputs(7505)));
    outputs(5627) <= layer0_outputs(10533);
    outputs(5628) <= layer0_outputs(3665);
    outputs(5629) <= layer0_outputs(2834);
    outputs(5630) <= not((layer0_outputs(8548)) and (layer0_outputs(3831)));
    outputs(5631) <= not((layer0_outputs(9693)) xor (layer0_outputs(1097)));
    outputs(5632) <= not(layer0_outputs(3940));
    outputs(5633) <= not(layer0_outputs(1386));
    outputs(5634) <= (layer0_outputs(11557)) xor (layer0_outputs(630));
    outputs(5635) <= layer0_outputs(5552);
    outputs(5636) <= layer0_outputs(12563);
    outputs(5637) <= not((layer0_outputs(9958)) xor (layer0_outputs(2025)));
    outputs(5638) <= (layer0_outputs(6533)) xor (layer0_outputs(4310));
    outputs(5639) <= not(layer0_outputs(397));
    outputs(5640) <= not((layer0_outputs(10625)) and (layer0_outputs(2485)));
    outputs(5641) <= layer0_outputs(2681);
    outputs(5642) <= not(layer0_outputs(9627));
    outputs(5643) <= layer0_outputs(10595);
    outputs(5644) <= layer0_outputs(11773);
    outputs(5645) <= layer0_outputs(11195);
    outputs(5646) <= layer0_outputs(11586);
    outputs(5647) <= (layer0_outputs(8687)) xor (layer0_outputs(878));
    outputs(5648) <= (layer0_outputs(9887)) xor (layer0_outputs(5108));
    outputs(5649) <= not((layer0_outputs(8060)) and (layer0_outputs(6761)));
    outputs(5650) <= layer0_outputs(12292);
    outputs(5651) <= not(layer0_outputs(2108));
    outputs(5652) <= not((layer0_outputs(3149)) or (layer0_outputs(4723)));
    outputs(5653) <= not((layer0_outputs(3176)) xor (layer0_outputs(10541)));
    outputs(5654) <= not((layer0_outputs(7041)) and (layer0_outputs(503)));
    outputs(5655) <= not(layer0_outputs(12497));
    outputs(5656) <= not(layer0_outputs(6602));
    outputs(5657) <= not(layer0_outputs(6029)) or (layer0_outputs(10164));
    outputs(5658) <= (layer0_outputs(7861)) xor (layer0_outputs(12346));
    outputs(5659) <= (layer0_outputs(1795)) or (layer0_outputs(4041));
    outputs(5660) <= layer0_outputs(10352);
    outputs(5661) <= not(layer0_outputs(4124));
    outputs(5662) <= (layer0_outputs(6899)) xor (layer0_outputs(12741));
    outputs(5663) <= not(layer0_outputs(1643));
    outputs(5664) <= layer0_outputs(5749);
    outputs(5665) <= layer0_outputs(11972);
    outputs(5666) <= layer0_outputs(8800);
    outputs(5667) <= not((layer0_outputs(3901)) xor (layer0_outputs(7606)));
    outputs(5668) <= not((layer0_outputs(10694)) xor (layer0_outputs(11869)));
    outputs(5669) <= not((layer0_outputs(2117)) and (layer0_outputs(12243)));
    outputs(5670) <= (layer0_outputs(4554)) and (layer0_outputs(4888));
    outputs(5671) <= not(layer0_outputs(1748));
    outputs(5672) <= not(layer0_outputs(6480));
    outputs(5673) <= not(layer0_outputs(3854));
    outputs(5674) <= not(layer0_outputs(5426)) or (layer0_outputs(3548));
    outputs(5675) <= (layer0_outputs(2198)) xor (layer0_outputs(7800));
    outputs(5676) <= not((layer0_outputs(10606)) xor (layer0_outputs(12645)));
    outputs(5677) <= not((layer0_outputs(9546)) and (layer0_outputs(12039)));
    outputs(5678) <= (layer0_outputs(4543)) xor (layer0_outputs(8640));
    outputs(5679) <= (layer0_outputs(1919)) xor (layer0_outputs(4639));
    outputs(5680) <= (layer0_outputs(2807)) xor (layer0_outputs(4715));
    outputs(5681) <= (layer0_outputs(392)) or (layer0_outputs(4742));
    outputs(5682) <= not(layer0_outputs(9796));
    outputs(5683) <= not(layer0_outputs(12070)) or (layer0_outputs(12005));
    outputs(5684) <= (layer0_outputs(5255)) xor (layer0_outputs(2006));
    outputs(5685) <= (layer0_outputs(1461)) and (layer0_outputs(8405));
    outputs(5686) <= not(layer0_outputs(6423));
    outputs(5687) <= layer0_outputs(11337);
    outputs(5688) <= not((layer0_outputs(11439)) or (layer0_outputs(7296)));
    outputs(5689) <= not(layer0_outputs(194)) or (layer0_outputs(822));
    outputs(5690) <= not((layer0_outputs(7183)) xor (layer0_outputs(10994)));
    outputs(5691) <= layer0_outputs(2645);
    outputs(5692) <= not((layer0_outputs(6299)) xor (layer0_outputs(5075)));
    outputs(5693) <= layer0_outputs(9772);
    outputs(5694) <= (layer0_outputs(5527)) xor (layer0_outputs(12404));
    outputs(5695) <= layer0_outputs(12342);
    outputs(5696) <= (layer0_outputs(7212)) and not (layer0_outputs(7528));
    outputs(5697) <= layer0_outputs(10473);
    outputs(5698) <= layer0_outputs(10037);
    outputs(5699) <= not((layer0_outputs(70)) or (layer0_outputs(5358)));
    outputs(5700) <= layer0_outputs(2096);
    outputs(5701) <= not(layer0_outputs(9053)) or (layer0_outputs(521));
    outputs(5702) <= (layer0_outputs(690)) xor (layer0_outputs(8736));
    outputs(5703) <= (layer0_outputs(3872)) and not (layer0_outputs(7790));
    outputs(5704) <= (layer0_outputs(744)) xor (layer0_outputs(11595));
    outputs(5705) <= layer0_outputs(4960);
    outputs(5706) <= not((layer0_outputs(8204)) xor (layer0_outputs(557)));
    outputs(5707) <= not(layer0_outputs(10562));
    outputs(5708) <= not(layer0_outputs(10915));
    outputs(5709) <= not((layer0_outputs(4441)) xor (layer0_outputs(2508)));
    outputs(5710) <= layer0_outputs(7148);
    outputs(5711) <= (layer0_outputs(8093)) xor (layer0_outputs(9340));
    outputs(5712) <= not(layer0_outputs(9744));
    outputs(5713) <= not(layer0_outputs(2726));
    outputs(5714) <= not((layer0_outputs(2859)) xor (layer0_outputs(12676)));
    outputs(5715) <= layer0_outputs(7434);
    outputs(5716) <= not(layer0_outputs(11417));
    outputs(5717) <= not(layer0_outputs(11198));
    outputs(5718) <= (layer0_outputs(1158)) and (layer0_outputs(5562));
    outputs(5719) <= not(layer0_outputs(4942)) or (layer0_outputs(4503));
    outputs(5720) <= not((layer0_outputs(2177)) and (layer0_outputs(4161)));
    outputs(5721) <= not(layer0_outputs(6360));
    outputs(5722) <= (layer0_outputs(10654)) and not (layer0_outputs(10443));
    outputs(5723) <= not((layer0_outputs(6808)) xor (layer0_outputs(8744)));
    outputs(5724) <= (layer0_outputs(5671)) xor (layer0_outputs(2098));
    outputs(5725) <= not((layer0_outputs(1949)) xor (layer0_outputs(12112)));
    outputs(5726) <= not((layer0_outputs(4840)) or (layer0_outputs(8672)));
    outputs(5727) <= layer0_outputs(4787);
    outputs(5728) <= (layer0_outputs(3946)) and not (layer0_outputs(11960));
    outputs(5729) <= not(layer0_outputs(6807));
    outputs(5730) <= not(layer0_outputs(1232));
    outputs(5731) <= (layer0_outputs(10837)) and (layer0_outputs(4764));
    outputs(5732) <= not(layer0_outputs(3510));
    outputs(5733) <= not((layer0_outputs(12743)) or (layer0_outputs(6822)));
    outputs(5734) <= layer0_outputs(11706);
    outputs(5735) <= not(layer0_outputs(3716));
    outputs(5736) <= not((layer0_outputs(1343)) xor (layer0_outputs(4055)));
    outputs(5737) <= layer0_outputs(4584);
    outputs(5738) <= (layer0_outputs(39)) or (layer0_outputs(129));
    outputs(5739) <= (layer0_outputs(3773)) and (layer0_outputs(11280));
    outputs(5740) <= (layer0_outputs(1018)) xor (layer0_outputs(40));
    outputs(5741) <= not((layer0_outputs(11204)) xor (layer0_outputs(5945)));
    outputs(5742) <= (layer0_outputs(12185)) and (layer0_outputs(2955));
    outputs(5743) <= not(layer0_outputs(4977));
    outputs(5744) <= layer0_outputs(9942);
    outputs(5745) <= not(layer0_outputs(2902)) or (layer0_outputs(4337));
    outputs(5746) <= not(layer0_outputs(5354));
    outputs(5747) <= layer0_outputs(9972);
    outputs(5748) <= not(layer0_outputs(2456));
    outputs(5749) <= (layer0_outputs(175)) and (layer0_outputs(9576));
    outputs(5750) <= not((layer0_outputs(11345)) xor (layer0_outputs(12707)));
    outputs(5751) <= not(layer0_outputs(7677));
    outputs(5752) <= not(layer0_outputs(5312)) or (layer0_outputs(11691));
    outputs(5753) <= (layer0_outputs(4961)) xor (layer0_outputs(9193));
    outputs(5754) <= not((layer0_outputs(11730)) xor (layer0_outputs(7021)));
    outputs(5755) <= not((layer0_outputs(4967)) xor (layer0_outputs(12339)));
    outputs(5756) <= not(layer0_outputs(11348));
    outputs(5757) <= (layer0_outputs(171)) xor (layer0_outputs(5603));
    outputs(5758) <= not((layer0_outputs(3782)) xor (layer0_outputs(7364)));
    outputs(5759) <= not((layer0_outputs(11547)) or (layer0_outputs(7375)));
    outputs(5760) <= not((layer0_outputs(2430)) xor (layer0_outputs(8127)));
    outputs(5761) <= (layer0_outputs(6421)) xor (layer0_outputs(9278));
    outputs(5762) <= (layer0_outputs(3811)) xor (layer0_outputs(9542));
    outputs(5763) <= not((layer0_outputs(12707)) or (layer0_outputs(9377)));
    outputs(5764) <= not(layer0_outputs(839));
    outputs(5765) <= (layer0_outputs(1500)) and not (layer0_outputs(6137));
    outputs(5766) <= not(layer0_outputs(9349)) or (layer0_outputs(4757));
    outputs(5767) <= (layer0_outputs(11370)) or (layer0_outputs(920));
    outputs(5768) <= (layer0_outputs(8037)) and (layer0_outputs(6240));
    outputs(5769) <= layer0_outputs(7617);
    outputs(5770) <= layer0_outputs(3386);
    outputs(5771) <= (layer0_outputs(12418)) and not (layer0_outputs(2660));
    outputs(5772) <= (layer0_outputs(3559)) xor (layer0_outputs(10507));
    outputs(5773) <= (layer0_outputs(1113)) xor (layer0_outputs(11557));
    outputs(5774) <= not((layer0_outputs(4195)) xor (layer0_outputs(9252)));
    outputs(5775) <= not((layer0_outputs(11199)) xor (layer0_outputs(10589)));
    outputs(5776) <= (layer0_outputs(9905)) and (layer0_outputs(8411));
    outputs(5777) <= layer0_outputs(11035);
    outputs(5778) <= not((layer0_outputs(995)) xor (layer0_outputs(7082)));
    outputs(5779) <= not(layer0_outputs(77));
    outputs(5780) <= (layer0_outputs(1740)) xor (layer0_outputs(9344));
    outputs(5781) <= layer0_outputs(6773);
    outputs(5782) <= layer0_outputs(3295);
    outputs(5783) <= not(layer0_outputs(3499));
    outputs(5784) <= (layer0_outputs(121)) and not (layer0_outputs(2168));
    outputs(5785) <= not(layer0_outputs(6352));
    outputs(5786) <= not(layer0_outputs(504));
    outputs(5787) <= layer0_outputs(1315);
    outputs(5788) <= layer0_outputs(11952);
    outputs(5789) <= (layer0_outputs(11682)) and not (layer0_outputs(7747));
    outputs(5790) <= layer0_outputs(11410);
    outputs(5791) <= layer0_outputs(3175);
    outputs(5792) <= not((layer0_outputs(9957)) xor (layer0_outputs(3299)));
    outputs(5793) <= (layer0_outputs(143)) xor (layer0_outputs(5595));
    outputs(5794) <= not((layer0_outputs(3026)) xor (layer0_outputs(8593)));
    outputs(5795) <= (layer0_outputs(9302)) and not (layer0_outputs(9926));
    outputs(5796) <= layer0_outputs(5730);
    outputs(5797) <= not((layer0_outputs(10559)) xor (layer0_outputs(7319)));
    outputs(5798) <= layer0_outputs(7141);
    outputs(5799) <= (layer0_outputs(7844)) xor (layer0_outputs(650));
    outputs(5800) <= (layer0_outputs(12024)) and not (layer0_outputs(4824));
    outputs(5801) <= not(layer0_outputs(780));
    outputs(5802) <= layer0_outputs(8925);
    outputs(5803) <= not((layer0_outputs(11820)) or (layer0_outputs(4219)));
    outputs(5804) <= not(layer0_outputs(4096));
    outputs(5805) <= not(layer0_outputs(11660));
    outputs(5806) <= not(layer0_outputs(3016));
    outputs(5807) <= (layer0_outputs(9822)) and not (layer0_outputs(5343));
    outputs(5808) <= not(layer0_outputs(10503));
    outputs(5809) <= layer0_outputs(12786);
    outputs(5810) <= layer0_outputs(5329);
    outputs(5811) <= not((layer0_outputs(9648)) or (layer0_outputs(2969)));
    outputs(5812) <= (layer0_outputs(4494)) xor (layer0_outputs(6199));
    outputs(5813) <= not((layer0_outputs(9273)) and (layer0_outputs(7937)));
    outputs(5814) <= (layer0_outputs(10215)) xor (layer0_outputs(9086));
    outputs(5815) <= (layer0_outputs(1703)) and not (layer0_outputs(9920));
    outputs(5816) <= not(layer0_outputs(2565));
    outputs(5817) <= (layer0_outputs(3513)) xor (layer0_outputs(3399));
    outputs(5818) <= layer0_outputs(7557);
    outputs(5819) <= not(layer0_outputs(12003));
    outputs(5820) <= layer0_outputs(1617);
    outputs(5821) <= not(layer0_outputs(12434)) or (layer0_outputs(509));
    outputs(5822) <= layer0_outputs(6291);
    outputs(5823) <= not((layer0_outputs(5667)) or (layer0_outputs(154)));
    outputs(5824) <= layer0_outputs(5648);
    outputs(5825) <= layer0_outputs(11410);
    outputs(5826) <= layer0_outputs(10332);
    outputs(5827) <= (layer0_outputs(11269)) and not (layer0_outputs(10683));
    outputs(5828) <= not(layer0_outputs(6127)) or (layer0_outputs(12493));
    outputs(5829) <= not((layer0_outputs(9396)) or (layer0_outputs(12610)));
    outputs(5830) <= (layer0_outputs(6703)) xor (layer0_outputs(1338));
    outputs(5831) <= (layer0_outputs(2791)) and not (layer0_outputs(4225));
    outputs(5832) <= not(layer0_outputs(285));
    outputs(5833) <= not((layer0_outputs(8407)) or (layer0_outputs(10616)));
    outputs(5834) <= not(layer0_outputs(1472));
    outputs(5835) <= not((layer0_outputs(1900)) xor (layer0_outputs(7903)));
    outputs(5836) <= layer0_outputs(3158);
    outputs(5837) <= not(layer0_outputs(2708)) or (layer0_outputs(9839));
    outputs(5838) <= not(layer0_outputs(7068));
    outputs(5839) <= not((layer0_outputs(6828)) xor (layer0_outputs(6094)));
    outputs(5840) <= (layer0_outputs(11479)) and (layer0_outputs(12353));
    outputs(5841) <= (layer0_outputs(3967)) xor (layer0_outputs(363));
    outputs(5842) <= (layer0_outputs(1116)) or (layer0_outputs(5377));
    outputs(5843) <= not((layer0_outputs(8795)) xor (layer0_outputs(7501)));
    outputs(5844) <= layer0_outputs(784);
    outputs(5845) <= not(layer0_outputs(135));
    outputs(5846) <= (layer0_outputs(11018)) and not (layer0_outputs(940));
    outputs(5847) <= (layer0_outputs(7389)) and (layer0_outputs(2439));
    outputs(5848) <= (layer0_outputs(12420)) and not (layer0_outputs(12549));
    outputs(5849) <= not((layer0_outputs(8236)) xor (layer0_outputs(6311)));
    outputs(5850) <= (layer0_outputs(8802)) and (layer0_outputs(5206));
    outputs(5851) <= (layer0_outputs(2079)) and not (layer0_outputs(2513));
    outputs(5852) <= layer0_outputs(3076);
    outputs(5853) <= not(layer0_outputs(7639));
    outputs(5854) <= layer0_outputs(595);
    outputs(5855) <= layer0_outputs(6572);
    outputs(5856) <= not((layer0_outputs(8887)) xor (layer0_outputs(9969)));
    outputs(5857) <= not(layer0_outputs(7450));
    outputs(5858) <= layer0_outputs(9606);
    outputs(5859) <= layer0_outputs(12327);
    outputs(5860) <= not(layer0_outputs(8393)) or (layer0_outputs(5567));
    outputs(5861) <= (layer0_outputs(3124)) and not (layer0_outputs(4600));
    outputs(5862) <= (layer0_outputs(8213)) xor (layer0_outputs(2874));
    outputs(5863) <= not((layer0_outputs(3095)) or (layer0_outputs(5008)));
    outputs(5864) <= not(layer0_outputs(4979));
    outputs(5865) <= (layer0_outputs(7089)) xor (layer0_outputs(10795));
    outputs(5866) <= (layer0_outputs(812)) xor (layer0_outputs(6863));
    outputs(5867) <= not((layer0_outputs(9037)) or (layer0_outputs(7750)));
    outputs(5868) <= not((layer0_outputs(11901)) xor (layer0_outputs(2620)));
    outputs(5869) <= (layer0_outputs(8785)) xor (layer0_outputs(8372));
    outputs(5870) <= layer0_outputs(11717);
    outputs(5871) <= not((layer0_outputs(4272)) or (layer0_outputs(12069)));
    outputs(5872) <= not(layer0_outputs(305));
    outputs(5873) <= (layer0_outputs(2552)) xor (layer0_outputs(2884));
    outputs(5874) <= layer0_outputs(7108);
    outputs(5875) <= layer0_outputs(7988);
    outputs(5876) <= (layer0_outputs(8468)) xor (layer0_outputs(8729));
    outputs(5877) <= (layer0_outputs(2621)) or (layer0_outputs(4010));
    outputs(5878) <= (layer0_outputs(2931)) and not (layer0_outputs(615));
    outputs(5879) <= (layer0_outputs(12511)) xor (layer0_outputs(6570));
    outputs(5880) <= (layer0_outputs(359)) or (layer0_outputs(5288));
    outputs(5881) <= layer0_outputs(2067);
    outputs(5882) <= not(layer0_outputs(11772));
    outputs(5883) <= (layer0_outputs(2230)) xor (layer0_outputs(8593));
    outputs(5884) <= layer0_outputs(11737);
    outputs(5885) <= not(layer0_outputs(5989));
    outputs(5886) <= not(layer0_outputs(10699));
    outputs(5887) <= (layer0_outputs(3352)) and not (layer0_outputs(1300));
    outputs(5888) <= not(layer0_outputs(2347));
    outputs(5889) <= (layer0_outputs(1193)) xor (layer0_outputs(976));
    outputs(5890) <= layer0_outputs(2267);
    outputs(5891) <= not(layer0_outputs(5071));
    outputs(5892) <= (layer0_outputs(7595)) and (layer0_outputs(8819));
    outputs(5893) <= not(layer0_outputs(7590));
    outputs(5894) <= not(layer0_outputs(4127));
    outputs(5895) <= not(layer0_outputs(7113));
    outputs(5896) <= not((layer0_outputs(11101)) or (layer0_outputs(1200)));
    outputs(5897) <= not((layer0_outputs(1504)) xor (layer0_outputs(5189)));
    outputs(5898) <= layer0_outputs(5949);
    outputs(5899) <= not(layer0_outputs(7085));
    outputs(5900) <= layer0_outputs(4669);
    outputs(5901) <= not((layer0_outputs(5208)) or (layer0_outputs(4480)));
    outputs(5902) <= not((layer0_outputs(10899)) or (layer0_outputs(2220)));
    outputs(5903) <= (layer0_outputs(6109)) and not (layer0_outputs(5614));
    outputs(5904) <= (layer0_outputs(4115)) xor (layer0_outputs(10096));
    outputs(5905) <= (layer0_outputs(6765)) and (layer0_outputs(10728));
    outputs(5906) <= not((layer0_outputs(2876)) or (layer0_outputs(3470)));
    outputs(5907) <= (layer0_outputs(6020)) xor (layer0_outputs(6152));
    outputs(5908) <= not(layer0_outputs(4025));
    outputs(5909) <= (layer0_outputs(916)) and not (layer0_outputs(10515));
    outputs(5910) <= layer0_outputs(1610);
    outputs(5911) <= not((layer0_outputs(2208)) xor (layer0_outputs(9657)));
    outputs(5912) <= not(layer0_outputs(10679)) or (layer0_outputs(5620));
    outputs(5913) <= not((layer0_outputs(6339)) xor (layer0_outputs(82)));
    outputs(5914) <= (layer0_outputs(3255)) xor (layer0_outputs(11203));
    outputs(5915) <= (layer0_outputs(7280)) xor (layer0_outputs(6641));
    outputs(5916) <= (layer0_outputs(2857)) xor (layer0_outputs(265));
    outputs(5917) <= layer0_outputs(10957);
    outputs(5918) <= not(layer0_outputs(10685)) or (layer0_outputs(11867));
    outputs(5919) <= (layer0_outputs(6290)) and not (layer0_outputs(4708));
    outputs(5920) <= layer0_outputs(9772);
    outputs(5921) <= not((layer0_outputs(7092)) xor (layer0_outputs(3962)));
    outputs(5922) <= (layer0_outputs(435)) xor (layer0_outputs(3602));
    outputs(5923) <= (layer0_outputs(12541)) and (layer0_outputs(4297));
    outputs(5924) <= layer0_outputs(6030);
    outputs(5925) <= not(layer0_outputs(604));
    outputs(5926) <= not((layer0_outputs(7372)) or (layer0_outputs(11731)));
    outputs(5927) <= not(layer0_outputs(3687));
    outputs(5928) <= not((layer0_outputs(2699)) xor (layer0_outputs(9284)));
    outputs(5929) <= (layer0_outputs(8248)) or (layer0_outputs(1759));
    outputs(5930) <= not((layer0_outputs(11301)) or (layer0_outputs(10341)));
    outputs(5931) <= layer0_outputs(11779);
    outputs(5932) <= not((layer0_outputs(5567)) xor (layer0_outputs(9254)));
    outputs(5933) <= layer0_outputs(4280);
    outputs(5934) <= not((layer0_outputs(9808)) xor (layer0_outputs(4968)));
    outputs(5935) <= layer0_outputs(6227);
    outputs(5936) <= (layer0_outputs(1314)) xor (layer0_outputs(6792));
    outputs(5937) <= layer0_outputs(12597);
    outputs(5938) <= layer0_outputs(8877);
    outputs(5939) <= not(layer0_outputs(11758));
    outputs(5940) <= (layer0_outputs(3528)) xor (layer0_outputs(9859));
    outputs(5941) <= not((layer0_outputs(5991)) or (layer0_outputs(718)));
    outputs(5942) <= not((layer0_outputs(12034)) or (layer0_outputs(9137)));
    outputs(5943) <= layer0_outputs(2270);
    outputs(5944) <= (layer0_outputs(4468)) xor (layer0_outputs(12182));
    outputs(5945) <= layer0_outputs(1284);
    outputs(5946) <= (layer0_outputs(10710)) xor (layer0_outputs(4200));
    outputs(5947) <= not(layer0_outputs(7059));
    outputs(5948) <= layer0_outputs(1096);
    outputs(5949) <= not((layer0_outputs(12614)) xor (layer0_outputs(9433)));
    outputs(5950) <= not(layer0_outputs(8440)) or (layer0_outputs(8676));
    outputs(5951) <= not((layer0_outputs(8720)) xor (layer0_outputs(826)));
    outputs(5952) <= not(layer0_outputs(8264)) or (layer0_outputs(9151));
    outputs(5953) <= not((layer0_outputs(12016)) or (layer0_outputs(3486)));
    outputs(5954) <= not(layer0_outputs(11659));
    outputs(5955) <= (layer0_outputs(10533)) and not (layer0_outputs(1846));
    outputs(5956) <= not(layer0_outputs(1946));
    outputs(5957) <= not(layer0_outputs(4056));
    outputs(5958) <= (layer0_outputs(3318)) xor (layer0_outputs(2360));
    outputs(5959) <= not(layer0_outputs(1573));
    outputs(5960) <= (layer0_outputs(7733)) and not (layer0_outputs(5259));
    outputs(5961) <= not(layer0_outputs(3405));
    outputs(5962) <= not(layer0_outputs(2801));
    outputs(5963) <= layer0_outputs(765);
    outputs(5964) <= not(layer0_outputs(4420));
    outputs(5965) <= not((layer0_outputs(10543)) xor (layer0_outputs(1976)));
    outputs(5966) <= layer0_outputs(9980);
    outputs(5967) <= not(layer0_outputs(5695)) or (layer0_outputs(7980));
    outputs(5968) <= (layer0_outputs(120)) xor (layer0_outputs(2777));
    outputs(5969) <= not((layer0_outputs(355)) xor (layer0_outputs(4518)));
    outputs(5970) <= (layer0_outputs(3484)) xor (layer0_outputs(2136));
    outputs(5971) <= layer0_outputs(8605);
    outputs(5972) <= (layer0_outputs(3904)) and not (layer0_outputs(4006));
    outputs(5973) <= not(layer0_outputs(3724)) or (layer0_outputs(11958));
    outputs(5974) <= not(layer0_outputs(8852));
    outputs(5975) <= not(layer0_outputs(5603));
    outputs(5976) <= not(layer0_outputs(4793));
    outputs(5977) <= (layer0_outputs(2684)) xor (layer0_outputs(1585));
    outputs(5978) <= (layer0_outputs(857)) xor (layer0_outputs(3787));
    outputs(5979) <= (layer0_outputs(2201)) and not (layer0_outputs(7790));
    outputs(5980) <= (layer0_outputs(2549)) and not (layer0_outputs(5835));
    outputs(5981) <= layer0_outputs(1659);
    outputs(5982) <= layer0_outputs(5844);
    outputs(5983) <= (layer0_outputs(5783)) and (layer0_outputs(8411));
    outputs(5984) <= not(layer0_outputs(11009));
    outputs(5985) <= (layer0_outputs(3605)) xor (layer0_outputs(1433));
    outputs(5986) <= (layer0_outputs(10750)) or (layer0_outputs(11003));
    outputs(5987) <= layer0_outputs(8281);
    outputs(5988) <= (layer0_outputs(441)) xor (layer0_outputs(11776));
    outputs(5989) <= not((layer0_outputs(9229)) xor (layer0_outputs(3774)));
    outputs(5990) <= (layer0_outputs(12612)) and not (layer0_outputs(3599));
    outputs(5991) <= not((layer0_outputs(12731)) xor (layer0_outputs(7803)));
    outputs(5992) <= layer0_outputs(5718);
    outputs(5993) <= (layer0_outputs(99)) xor (layer0_outputs(11250));
    outputs(5994) <= (layer0_outputs(10048)) xor (layer0_outputs(9761));
    outputs(5995) <= (layer0_outputs(10257)) xor (layer0_outputs(12255));
    outputs(5996) <= not((layer0_outputs(3036)) or (layer0_outputs(3160)));
    outputs(5997) <= (layer0_outputs(954)) and not (layer0_outputs(8975));
    outputs(5998) <= (layer0_outputs(10317)) xor (layer0_outputs(5832));
    outputs(5999) <= layer0_outputs(2435);
    outputs(6000) <= layer0_outputs(8700);
    outputs(6001) <= not(layer0_outputs(6029)) or (layer0_outputs(9059));
    outputs(6002) <= not((layer0_outputs(4428)) and (layer0_outputs(3557)));
    outputs(6003) <= not(layer0_outputs(10152)) or (layer0_outputs(7902));
    outputs(6004) <= layer0_outputs(2822);
    outputs(6005) <= not(layer0_outputs(7643));
    outputs(6006) <= layer0_outputs(12558);
    outputs(6007) <= (layer0_outputs(4750)) and (layer0_outputs(7415));
    outputs(6008) <= not((layer0_outputs(6564)) xor (layer0_outputs(3267)));
    outputs(6009) <= not((layer0_outputs(6099)) xor (layer0_outputs(10866)));
    outputs(6010) <= not(layer0_outputs(1336));
    outputs(6011) <= layer0_outputs(9106);
    outputs(6012) <= layer0_outputs(734);
    outputs(6013) <= (layer0_outputs(9310)) xor (layer0_outputs(3840));
    outputs(6014) <= layer0_outputs(8273);
    outputs(6015) <= not(layer0_outputs(8847)) or (layer0_outputs(10385));
    outputs(6016) <= (layer0_outputs(5233)) or (layer0_outputs(27));
    outputs(6017) <= not((layer0_outputs(2487)) or (layer0_outputs(1460)));
    outputs(6018) <= layer0_outputs(14);
    outputs(6019) <= layer0_outputs(3733);
    outputs(6020) <= not(layer0_outputs(7886));
    outputs(6021) <= not(layer0_outputs(5867));
    outputs(6022) <= not((layer0_outputs(1521)) xor (layer0_outputs(8892)));
    outputs(6023) <= (layer0_outputs(4969)) xor (layer0_outputs(11237));
    outputs(6024) <= not(layer0_outputs(3724)) or (layer0_outputs(956));
    outputs(6025) <= (layer0_outputs(32)) xor (layer0_outputs(4163));
    outputs(6026) <= (layer0_outputs(10057)) and not (layer0_outputs(5695));
    outputs(6027) <= (layer0_outputs(6761)) xor (layer0_outputs(9422));
    outputs(6028) <= not((layer0_outputs(10997)) xor (layer0_outputs(9919)));
    outputs(6029) <= not(layer0_outputs(699));
    outputs(6030) <= not(layer0_outputs(6503));
    outputs(6031) <= (layer0_outputs(1357)) and not (layer0_outputs(385));
    outputs(6032) <= not(layer0_outputs(9955));
    outputs(6033) <= layer0_outputs(7592);
    outputs(6034) <= not(layer0_outputs(3225));
    outputs(6035) <= not((layer0_outputs(2240)) xor (layer0_outputs(5475)));
    outputs(6036) <= not(layer0_outputs(189)) or (layer0_outputs(12548));
    outputs(6037) <= not(layer0_outputs(11096));
    outputs(6038) <= (layer0_outputs(3909)) and not (layer0_outputs(11128));
    outputs(6039) <= (layer0_outputs(2574)) and (layer0_outputs(2321));
    outputs(6040) <= layer0_outputs(12559);
    outputs(6041) <= (layer0_outputs(12651)) xor (layer0_outputs(7166));
    outputs(6042) <= not(layer0_outputs(6959));
    outputs(6043) <= layer0_outputs(1158);
    outputs(6044) <= not(layer0_outputs(8813)) or (layer0_outputs(1710));
    outputs(6045) <= not((layer0_outputs(5020)) xor (layer0_outputs(377)));
    outputs(6046) <= (layer0_outputs(8130)) xor (layer0_outputs(4294));
    outputs(6047) <= layer0_outputs(2169);
    outputs(6048) <= layer0_outputs(53);
    outputs(6049) <= not(layer0_outputs(12214));
    outputs(6050) <= layer0_outputs(10756);
    outputs(6051) <= not((layer0_outputs(220)) xor (layer0_outputs(12632)));
    outputs(6052) <= layer0_outputs(7696);
    outputs(6053) <= not((layer0_outputs(12161)) xor (layer0_outputs(4575)));
    outputs(6054) <= not(layer0_outputs(7060));
    outputs(6055) <= (layer0_outputs(2561)) and not (layer0_outputs(5920));
    outputs(6056) <= not(layer0_outputs(1337));
    outputs(6057) <= layer0_outputs(8137);
    outputs(6058) <= layer0_outputs(2226);
    outputs(6059) <= layer0_outputs(4050);
    outputs(6060) <= not((layer0_outputs(5825)) xor (layer0_outputs(5009)));
    outputs(6061) <= not((layer0_outputs(5132)) xor (layer0_outputs(9215)));
    outputs(6062) <= not(layer0_outputs(4089));
    outputs(6063) <= (layer0_outputs(6977)) xor (layer0_outputs(10848));
    outputs(6064) <= not(layer0_outputs(6201));
    outputs(6065) <= not(layer0_outputs(11474)) or (layer0_outputs(9986));
    outputs(6066) <= not(layer0_outputs(6050));
    outputs(6067) <= not(layer0_outputs(11360));
    outputs(6068) <= layer0_outputs(2556);
    outputs(6069) <= not(layer0_outputs(6064));
    outputs(6070) <= not(layer0_outputs(570));
    outputs(6071) <= (layer0_outputs(11309)) and not (layer0_outputs(8904));
    outputs(6072) <= (layer0_outputs(11320)) and not (layer0_outputs(10035));
    outputs(6073) <= (layer0_outputs(8026)) xor (layer0_outputs(1771));
    outputs(6074) <= not((layer0_outputs(1652)) xor (layer0_outputs(8824)));
    outputs(6075) <= not((layer0_outputs(10062)) xor (layer0_outputs(7588)));
    outputs(6076) <= not((layer0_outputs(12461)) xor (layer0_outputs(6918)));
    outputs(6077) <= not(layer0_outputs(1030)) or (layer0_outputs(242));
    outputs(6078) <= not(layer0_outputs(6822));
    outputs(6079) <= not(layer0_outputs(3792));
    outputs(6080) <= layer0_outputs(4531);
    outputs(6081) <= layer0_outputs(6814);
    outputs(6082) <= (layer0_outputs(556)) and not (layer0_outputs(2315));
    outputs(6083) <= not(layer0_outputs(7363));
    outputs(6084) <= not((layer0_outputs(10703)) xor (layer0_outputs(439)));
    outputs(6085) <= (layer0_outputs(8288)) and (layer0_outputs(8309));
    outputs(6086) <= not((layer0_outputs(8327)) xor (layer0_outputs(278)));
    outputs(6087) <= layer0_outputs(1168);
    outputs(6088) <= layer0_outputs(4458);
    outputs(6089) <= layer0_outputs(7784);
    outputs(6090) <= not((layer0_outputs(2619)) and (layer0_outputs(5532)));
    outputs(6091) <= not(layer0_outputs(6728));
    outputs(6092) <= (layer0_outputs(30)) and not (layer0_outputs(11614));
    outputs(6093) <= (layer0_outputs(12402)) and not (layer0_outputs(7913));
    outputs(6094) <= not(layer0_outputs(7690)) or (layer0_outputs(697));
    outputs(6095) <= layer0_outputs(7343);
    outputs(6096) <= not((layer0_outputs(4935)) xor (layer0_outputs(10311)));
    outputs(6097) <= (layer0_outputs(11617)) xor (layer0_outputs(3684));
    outputs(6098) <= (layer0_outputs(8083)) and not (layer0_outputs(9219));
    outputs(6099) <= not(layer0_outputs(5958));
    outputs(6100) <= not(layer0_outputs(11087));
    outputs(6101) <= layer0_outputs(8630);
    outputs(6102) <= layer0_outputs(2734);
    outputs(6103) <= layer0_outputs(11554);
    outputs(6104) <= not(layer0_outputs(2257));
    outputs(6105) <= not(layer0_outputs(11442));
    outputs(6106) <= not((layer0_outputs(12339)) xor (layer0_outputs(4233)));
    outputs(6107) <= (layer0_outputs(10188)) and not (layer0_outputs(11374));
    outputs(6108) <= not(layer0_outputs(10585));
    outputs(6109) <= not((layer0_outputs(6387)) xor (layer0_outputs(10226)));
    outputs(6110) <= (layer0_outputs(547)) xor (layer0_outputs(9852));
    outputs(6111) <= (layer0_outputs(9833)) and not (layer0_outputs(1251));
    outputs(6112) <= not(layer0_outputs(3793));
    outputs(6113) <= not(layer0_outputs(7769)) or (layer0_outputs(7237));
    outputs(6114) <= not(layer0_outputs(988));
    outputs(6115) <= not((layer0_outputs(9910)) or (layer0_outputs(5692)));
    outputs(6116) <= layer0_outputs(4009);
    outputs(6117) <= (layer0_outputs(2498)) xor (layer0_outputs(9944));
    outputs(6118) <= layer0_outputs(11429);
    outputs(6119) <= (layer0_outputs(11070)) xor (layer0_outputs(36));
    outputs(6120) <= (layer0_outputs(7542)) and not (layer0_outputs(9740));
    outputs(6121) <= (layer0_outputs(3139)) xor (layer0_outputs(7348));
    outputs(6122) <= (layer0_outputs(6584)) xor (layer0_outputs(2454));
    outputs(6123) <= not((layer0_outputs(292)) xor (layer0_outputs(2251)));
    outputs(6124) <= layer0_outputs(10713);
    outputs(6125) <= (layer0_outputs(7216)) and (layer0_outputs(8913));
    outputs(6126) <= not((layer0_outputs(7065)) or (layer0_outputs(1839)));
    outputs(6127) <= layer0_outputs(11539);
    outputs(6128) <= (layer0_outputs(1054)) and not (layer0_outputs(1669));
    outputs(6129) <= not(layer0_outputs(2444));
    outputs(6130) <= not(layer0_outputs(12164));
    outputs(6131) <= not(layer0_outputs(12018));
    outputs(6132) <= (layer0_outputs(1123)) and not (layer0_outputs(10501));
    outputs(6133) <= not((layer0_outputs(10168)) xor (layer0_outputs(4044)));
    outputs(6134) <= not(layer0_outputs(1851));
    outputs(6135) <= (layer0_outputs(125)) and not (layer0_outputs(9874));
    outputs(6136) <= (layer0_outputs(11291)) xor (layer0_outputs(10809));
    outputs(6137) <= not(layer0_outputs(7522));
    outputs(6138) <= layer0_outputs(6336);
    outputs(6139) <= layer0_outputs(9408);
    outputs(6140) <= (layer0_outputs(2441)) or (layer0_outputs(7608));
    outputs(6141) <= not((layer0_outputs(8855)) or (layer0_outputs(12485)));
    outputs(6142) <= (layer0_outputs(2730)) xor (layer0_outputs(2308));
    outputs(6143) <= (layer0_outputs(6035)) and (layer0_outputs(12739));
    outputs(6144) <= (layer0_outputs(11432)) and (layer0_outputs(3124));
    outputs(6145) <= not(layer0_outputs(5497));
    outputs(6146) <= layer0_outputs(4299);
    outputs(6147) <= not((layer0_outputs(3037)) and (layer0_outputs(5120)));
    outputs(6148) <= not(layer0_outputs(775));
    outputs(6149) <= layer0_outputs(1119);
    outputs(6150) <= not(layer0_outputs(7538));
    outputs(6151) <= not(layer0_outputs(650));
    outputs(6152) <= (layer0_outputs(1879)) xor (layer0_outputs(11335));
    outputs(6153) <= (layer0_outputs(6340)) xor (layer0_outputs(10669));
    outputs(6154) <= (layer0_outputs(7912)) and not (layer0_outputs(7830));
    outputs(6155) <= (layer0_outputs(12503)) and not (layer0_outputs(6215));
    outputs(6156) <= (layer0_outputs(6539)) xor (layer0_outputs(4422));
    outputs(6157) <= layer0_outputs(2001);
    outputs(6158) <= (layer0_outputs(2206)) and not (layer0_outputs(530));
    outputs(6159) <= not(layer0_outputs(9172));
    outputs(6160) <= (layer0_outputs(3583)) and not (layer0_outputs(9181));
    outputs(6161) <= (layer0_outputs(2173)) and (layer0_outputs(10760));
    outputs(6162) <= not(layer0_outputs(1211));
    outputs(6163) <= not((layer0_outputs(4675)) xor (layer0_outputs(2856)));
    outputs(6164) <= (layer0_outputs(5267)) xor (layer0_outputs(2351));
    outputs(6165) <= layer0_outputs(6289);
    outputs(6166) <= not(layer0_outputs(4547));
    outputs(6167) <= not(layer0_outputs(12781));
    outputs(6168) <= (layer0_outputs(3084)) and (layer0_outputs(4976));
    outputs(6169) <= (layer0_outputs(10684)) xor (layer0_outputs(4614));
    outputs(6170) <= layer0_outputs(11721);
    outputs(6171) <= not((layer0_outputs(9825)) or (layer0_outputs(6958)));
    outputs(6172) <= not((layer0_outputs(3428)) xor (layer0_outputs(11077)));
    outputs(6173) <= layer0_outputs(8507);
    outputs(6174) <= (layer0_outputs(5858)) xor (layer0_outputs(3971));
    outputs(6175) <= (layer0_outputs(12624)) and (layer0_outputs(11166));
    outputs(6176) <= (layer0_outputs(2591)) and (layer0_outputs(5732));
    outputs(6177) <= layer0_outputs(10783);
    outputs(6178) <= (layer0_outputs(12370)) and not (layer0_outputs(354));
    outputs(6179) <= layer0_outputs(4373);
    outputs(6180) <= not(layer0_outputs(49));
    outputs(6181) <= not((layer0_outputs(4826)) xor (layer0_outputs(11635)));
    outputs(6182) <= not(layer0_outputs(5135)) or (layer0_outputs(1742));
    outputs(6183) <= not(layer0_outputs(8732)) or (layer0_outputs(3606));
    outputs(6184) <= layer0_outputs(10468);
    outputs(6185) <= (layer0_outputs(8756)) xor (layer0_outputs(5720));
    outputs(6186) <= not(layer0_outputs(11815));
    outputs(6187) <= layer0_outputs(2297);
    outputs(6188) <= layer0_outputs(969);
    outputs(6189) <= not(layer0_outputs(5159));
    outputs(6190) <= layer0_outputs(3325);
    outputs(6191) <= (layer0_outputs(5240)) xor (layer0_outputs(1330));
    outputs(6192) <= not((layer0_outputs(386)) xor (layer0_outputs(1465)));
    outputs(6193) <= (layer0_outputs(7204)) or (layer0_outputs(8999));
    outputs(6194) <= not(layer0_outputs(12749));
    outputs(6195) <= not(layer0_outputs(10216));
    outputs(6196) <= not((layer0_outputs(11160)) xor (layer0_outputs(3532)));
    outputs(6197) <= (layer0_outputs(8313)) and (layer0_outputs(8395));
    outputs(6198) <= (layer0_outputs(1245)) xor (layer0_outputs(2945));
    outputs(6199) <= not((layer0_outputs(11792)) xor (layer0_outputs(5900)));
    outputs(6200) <= not((layer0_outputs(10004)) and (layer0_outputs(5596)));
    outputs(6201) <= layer0_outputs(10480);
    outputs(6202) <= layer0_outputs(11895);
    outputs(6203) <= not(layer0_outputs(1037));
    outputs(6204) <= (layer0_outputs(4433)) xor (layer0_outputs(8194));
    outputs(6205) <= layer0_outputs(6374);
    outputs(6206) <= (layer0_outputs(415)) or (layer0_outputs(10320));
    outputs(6207) <= not(layer0_outputs(6271)) or (layer0_outputs(3681));
    outputs(6208) <= layer0_outputs(4362);
    outputs(6209) <= layer0_outputs(3278);
    outputs(6210) <= not((layer0_outputs(10766)) or (layer0_outputs(5070)));
    outputs(6211) <= not((layer0_outputs(1744)) xor (layer0_outputs(4890)));
    outputs(6212) <= not((layer0_outputs(11925)) or (layer0_outputs(1450)));
    outputs(6213) <= layer0_outputs(7340);
    outputs(6214) <= layer0_outputs(12210);
    outputs(6215) <= (layer0_outputs(2556)) or (layer0_outputs(7596));
    outputs(6216) <= not(layer0_outputs(9837)) or (layer0_outputs(646));
    outputs(6217) <= layer0_outputs(6260);
    outputs(6218) <= layer0_outputs(321);
    outputs(6219) <= not(layer0_outputs(3187));
    outputs(6220) <= not((layer0_outputs(5421)) xor (layer0_outputs(12796)));
    outputs(6221) <= not(layer0_outputs(12220)) or (layer0_outputs(4268));
    outputs(6222) <= (layer0_outputs(4586)) and not (layer0_outputs(11510));
    outputs(6223) <= (layer0_outputs(10740)) xor (layer0_outputs(8263));
    outputs(6224) <= not(layer0_outputs(2013));
    outputs(6225) <= not(layer0_outputs(2440));
    outputs(6226) <= layer0_outputs(149);
    outputs(6227) <= (layer0_outputs(6021)) and not (layer0_outputs(11342));
    outputs(6228) <= not((layer0_outputs(11357)) xor (layer0_outputs(3206)));
    outputs(6229) <= (layer0_outputs(5394)) xor (layer0_outputs(12752));
    outputs(6230) <= layer0_outputs(9243);
    outputs(6231) <= layer0_outputs(9217);
    outputs(6232) <= (layer0_outputs(5623)) or (layer0_outputs(1999));
    outputs(6233) <= layer0_outputs(9271);
    outputs(6234) <= (layer0_outputs(10624)) xor (layer0_outputs(6232));
    outputs(6235) <= not(layer0_outputs(9982));
    outputs(6236) <= not(layer0_outputs(10327));
    outputs(6237) <= (layer0_outputs(4383)) xor (layer0_outputs(1315));
    outputs(6238) <= not((layer0_outputs(10176)) or (layer0_outputs(10445)));
    outputs(6239) <= not(layer0_outputs(11214));
    outputs(6240) <= not(layer0_outputs(2437)) or (layer0_outputs(10718));
    outputs(6241) <= layer0_outputs(5098);
    outputs(6242) <= layer0_outputs(8360);
    outputs(6243) <= not(layer0_outputs(11102));
    outputs(6244) <= not((layer0_outputs(2616)) xor (layer0_outputs(2281)));
    outputs(6245) <= not(layer0_outputs(9925));
    outputs(6246) <= (layer0_outputs(3945)) and (layer0_outputs(7057));
    outputs(6247) <= not((layer0_outputs(2463)) xor (layer0_outputs(11067)));
    outputs(6248) <= (layer0_outputs(3001)) and not (layer0_outputs(1387));
    outputs(6249) <= not((layer0_outputs(4304)) xor (layer0_outputs(12058)));
    outputs(6250) <= not(layer0_outputs(378));
    outputs(6251) <= not((layer0_outputs(5101)) xor (layer0_outputs(3473)));
    outputs(6252) <= not((layer0_outputs(7240)) xor (layer0_outputs(1155)));
    outputs(6253) <= not((layer0_outputs(4463)) xor (layer0_outputs(1809)));
    outputs(6254) <= layer0_outputs(10564);
    outputs(6255) <= not((layer0_outputs(8675)) xor (layer0_outputs(1254)));
    outputs(6256) <= layer0_outputs(3275);
    outputs(6257) <= layer0_outputs(7726);
    outputs(6258) <= not((layer0_outputs(6867)) xor (layer0_outputs(4480)));
    outputs(6259) <= (layer0_outputs(7748)) and not (layer0_outputs(4324));
    outputs(6260) <= not(layer0_outputs(5299));
    outputs(6261) <= (layer0_outputs(9531)) xor (layer0_outputs(10761));
    outputs(6262) <= layer0_outputs(6653);
    outputs(6263) <= not(layer0_outputs(5974));
    outputs(6264) <= not(layer0_outputs(8968));
    outputs(6265) <= not((layer0_outputs(3445)) or (layer0_outputs(2044)));
    outputs(6266) <= not(layer0_outputs(2811));
    outputs(6267) <= not(layer0_outputs(10512));
    outputs(6268) <= layer0_outputs(2797);
    outputs(6269) <= layer0_outputs(9694);
    outputs(6270) <= layer0_outputs(2995);
    outputs(6271) <= layer0_outputs(9075);
    outputs(6272) <= not(layer0_outputs(3653));
    outputs(6273) <= layer0_outputs(8011);
    outputs(6274) <= not(layer0_outputs(1914));
    outputs(6275) <= not((layer0_outputs(2127)) xor (layer0_outputs(3288)));
    outputs(6276) <= not(layer0_outputs(9322));
    outputs(6277) <= (layer0_outputs(3968)) and not (layer0_outputs(9671));
    outputs(6278) <= not(layer0_outputs(10703));
    outputs(6279) <= not(layer0_outputs(7992)) or (layer0_outputs(2410));
    outputs(6280) <= layer0_outputs(12268);
    outputs(6281) <= layer0_outputs(10321);
    outputs(6282) <= not((layer0_outputs(802)) xor (layer0_outputs(11872)));
    outputs(6283) <= not((layer0_outputs(692)) xor (layer0_outputs(4353)));
    outputs(6284) <= not((layer0_outputs(1499)) or (layer0_outputs(2796)));
    outputs(6285) <= layer0_outputs(1379);
    outputs(6286) <= (layer0_outputs(10739)) xor (layer0_outputs(11716));
    outputs(6287) <= layer0_outputs(1340);
    outputs(6288) <= (layer0_outputs(4018)) xor (layer0_outputs(4363));
    outputs(6289) <= not((layer0_outputs(6161)) xor (layer0_outputs(6165)));
    outputs(6290) <= (layer0_outputs(11126)) xor (layer0_outputs(10399));
    outputs(6291) <= layer0_outputs(259);
    outputs(6292) <= not((layer0_outputs(3036)) xor (layer0_outputs(632)));
    outputs(6293) <= not((layer0_outputs(5972)) xor (layer0_outputs(6457)));
    outputs(6294) <= not((layer0_outputs(5862)) or (layer0_outputs(11565)));
    outputs(6295) <= not((layer0_outputs(11972)) xor (layer0_outputs(12755)));
    outputs(6296) <= not(layer0_outputs(11715));
    outputs(6297) <= (layer0_outputs(7229)) xor (layer0_outputs(1148));
    outputs(6298) <= (layer0_outputs(10860)) xor (layer0_outputs(6353));
    outputs(6299) <= (layer0_outputs(10001)) xor (layer0_outputs(8999));
    outputs(6300) <= layer0_outputs(12035);
    outputs(6301) <= not((layer0_outputs(5605)) or (layer0_outputs(2115)));
    outputs(6302) <= not(layer0_outputs(10688));
    outputs(6303) <= (layer0_outputs(2167)) and (layer0_outputs(11633));
    outputs(6304) <= (layer0_outputs(8874)) and (layer0_outputs(6483));
    outputs(6305) <= layer0_outputs(7720);
    outputs(6306) <= (layer0_outputs(11981)) xor (layer0_outputs(7771));
    outputs(6307) <= (layer0_outputs(789)) and (layer0_outputs(8790));
    outputs(6308) <= (layer0_outputs(8591)) and (layer0_outputs(12113));
    outputs(6309) <= layer0_outputs(8579);
    outputs(6310) <= not((layer0_outputs(2753)) xor (layer0_outputs(7395)));
    outputs(6311) <= not((layer0_outputs(9943)) xor (layer0_outputs(6714)));
    outputs(6312) <= not(layer0_outputs(1106)) or (layer0_outputs(12342));
    outputs(6313) <= (layer0_outputs(12426)) xor (layer0_outputs(6952));
    outputs(6314) <= layer0_outputs(7569);
    outputs(6315) <= (layer0_outputs(10191)) and not (layer0_outputs(7504));
    outputs(6316) <= not(layer0_outputs(9687));
    outputs(6317) <= not((layer0_outputs(8178)) xor (layer0_outputs(6139)));
    outputs(6318) <= not((layer0_outputs(10363)) xor (layer0_outputs(11164)));
    outputs(6319) <= not(layer0_outputs(2745));
    outputs(6320) <= (layer0_outputs(5618)) and not (layer0_outputs(10407));
    outputs(6321) <= not((layer0_outputs(1332)) xor (layer0_outputs(8165)));
    outputs(6322) <= layer0_outputs(3087);
    outputs(6323) <= not((layer0_outputs(5230)) or (layer0_outputs(1058)));
    outputs(6324) <= layer0_outputs(7427);
    outputs(6325) <= (layer0_outputs(4210)) and (layer0_outputs(1534));
    outputs(6326) <= (layer0_outputs(8509)) or (layer0_outputs(337));
    outputs(6327) <= (layer0_outputs(995)) xor (layer0_outputs(5891));
    outputs(6328) <= not((layer0_outputs(2381)) or (layer0_outputs(6279)));
    outputs(6329) <= (layer0_outputs(6060)) xor (layer0_outputs(5602));
    outputs(6330) <= not((layer0_outputs(729)) xor (layer0_outputs(8516)));
    outputs(6331) <= not((layer0_outputs(8134)) xor (layer0_outputs(1540)));
    outputs(6332) <= (layer0_outputs(12670)) or (layer0_outputs(5227));
    outputs(6333) <= not(layer0_outputs(9207));
    outputs(6334) <= layer0_outputs(11624);
    outputs(6335) <= not((layer0_outputs(9158)) xor (layer0_outputs(12104)));
    outputs(6336) <= (layer0_outputs(1735)) xor (layer0_outputs(6750));
    outputs(6337) <= not((layer0_outputs(323)) or (layer0_outputs(6969)));
    outputs(6338) <= (layer0_outputs(9225)) xor (layer0_outputs(3009));
    outputs(6339) <= not((layer0_outputs(12608)) xor (layer0_outputs(8112)));
    outputs(6340) <= not(layer0_outputs(6269));
    outputs(6341) <= not((layer0_outputs(3736)) xor (layer0_outputs(8040)));
    outputs(6342) <= (layer0_outputs(4949)) and not (layer0_outputs(12434));
    outputs(6343) <= not(layer0_outputs(10665));
    outputs(6344) <= not(layer0_outputs(406));
    outputs(6345) <= (layer0_outputs(11941)) xor (layer0_outputs(8538));
    outputs(6346) <= not(layer0_outputs(5683));
    outputs(6347) <= (layer0_outputs(12154)) xor (layer0_outputs(11267));
    outputs(6348) <= layer0_outputs(2920);
    outputs(6349) <= layer0_outputs(3516);
    outputs(6350) <= (layer0_outputs(10303)) xor (layer0_outputs(2944));
    outputs(6351) <= (layer0_outputs(5949)) xor (layer0_outputs(3093));
    outputs(6352) <= (layer0_outputs(582)) xor (layer0_outputs(3201));
    outputs(6353) <= layer0_outputs(4298);
    outputs(6354) <= (layer0_outputs(4951)) xor (layer0_outputs(9735));
    outputs(6355) <= layer0_outputs(11014);
    outputs(6356) <= not(layer0_outputs(170)) or (layer0_outputs(3570));
    outputs(6357) <= (layer0_outputs(8588)) and not (layer0_outputs(6447));
    outputs(6358) <= (layer0_outputs(3679)) xor (layer0_outputs(1560));
    outputs(6359) <= layer0_outputs(6536);
    outputs(6360) <= not(layer0_outputs(5482));
    outputs(6361) <= not(layer0_outputs(12573));
    outputs(6362) <= not((layer0_outputs(2940)) or (layer0_outputs(5202)));
    outputs(6363) <= not(layer0_outputs(7162));
    outputs(6364) <= (layer0_outputs(8336)) and not (layer0_outputs(11843));
    outputs(6365) <= layer0_outputs(12584);
    outputs(6366) <= not((layer0_outputs(3103)) xor (layer0_outputs(1721)));
    outputs(6367) <= layer0_outputs(6814);
    outputs(6368) <= not(layer0_outputs(12723));
    outputs(6369) <= (layer0_outputs(1794)) xor (layer0_outputs(4764));
    outputs(6370) <= layer0_outputs(5898);
    outputs(6371) <= (layer0_outputs(12662)) and (layer0_outputs(4755));
    outputs(6372) <= not((layer0_outputs(4510)) xor (layer0_outputs(11511)));
    outputs(6373) <= not(layer0_outputs(12));
    outputs(6374) <= not(layer0_outputs(3320));
    outputs(6375) <= (layer0_outputs(11622)) and not (layer0_outputs(4657));
    outputs(6376) <= not((layer0_outputs(4735)) xor (layer0_outputs(8657)));
    outputs(6377) <= not(layer0_outputs(38));
    outputs(6378) <= (layer0_outputs(625)) and not (layer0_outputs(5666));
    outputs(6379) <= not((layer0_outputs(880)) and (layer0_outputs(10020)));
    outputs(6380) <= (layer0_outputs(3216)) and (layer0_outputs(42));
    outputs(6381) <= layer0_outputs(1379);
    outputs(6382) <= not(layer0_outputs(12382));
    outputs(6383) <= not((layer0_outputs(3643)) or (layer0_outputs(10094)));
    outputs(6384) <= (layer0_outputs(9559)) or (layer0_outputs(5484));
    outputs(6385) <= not(layer0_outputs(12245));
    outputs(6386) <= not((layer0_outputs(1595)) xor (layer0_outputs(12266)));
    outputs(6387) <= layer0_outputs(1754);
    outputs(6388) <= layer0_outputs(10410);
    outputs(6389) <= (layer0_outputs(10306)) or (layer0_outputs(11904));
    outputs(6390) <= (layer0_outputs(9347)) and (layer0_outputs(10329));
    outputs(6391) <= not(layer0_outputs(4681));
    outputs(6392) <= not((layer0_outputs(10271)) xor (layer0_outputs(11724)));
    outputs(6393) <= (layer0_outputs(9412)) and not (layer0_outputs(11876));
    outputs(6394) <= (layer0_outputs(8008)) and not (layer0_outputs(414));
    outputs(6395) <= (layer0_outputs(2129)) xor (layer0_outputs(10769));
    outputs(6396) <= (layer0_outputs(5539)) xor (layer0_outputs(181));
    outputs(6397) <= not((layer0_outputs(6137)) xor (layer0_outputs(3831)));
    outputs(6398) <= not(layer0_outputs(3409));
    outputs(6399) <= not(layer0_outputs(905)) or (layer0_outputs(7789));
    outputs(6400) <= not((layer0_outputs(3393)) and (layer0_outputs(2771)));
    outputs(6401) <= (layer0_outputs(434)) xor (layer0_outputs(510));
    outputs(6402) <= not((layer0_outputs(614)) and (layer0_outputs(9270)));
    outputs(6403) <= layer0_outputs(1615);
    outputs(6404) <= layer0_outputs(11868);
    outputs(6405) <= layer0_outputs(3623);
    outputs(6406) <= not(layer0_outputs(4791));
    outputs(6407) <= not((layer0_outputs(540)) xor (layer0_outputs(1783)));
    outputs(6408) <= not((layer0_outputs(11673)) xor (layer0_outputs(8689)));
    outputs(6409) <= not(layer0_outputs(10233));
    outputs(6410) <= not(layer0_outputs(9893));
    outputs(6411) <= not(layer0_outputs(6259));
    outputs(6412) <= not((layer0_outputs(4258)) xor (layer0_outputs(12642)));
    outputs(6413) <= not(layer0_outputs(8009)) or (layer0_outputs(8427));
    outputs(6414) <= layer0_outputs(5947);
    outputs(6415) <= (layer0_outputs(8473)) xor (layer0_outputs(4468));
    outputs(6416) <= not(layer0_outputs(4497));
    outputs(6417) <= not((layer0_outputs(4843)) xor (layer0_outputs(7682)));
    outputs(6418) <= (layer0_outputs(4240)) xor (layer0_outputs(4062));
    outputs(6419) <= (layer0_outputs(11384)) and not (layer0_outputs(7688));
    outputs(6420) <= not(layer0_outputs(2976)) or (layer0_outputs(8156));
    outputs(6421) <= (layer0_outputs(8595)) xor (layer0_outputs(1017));
    outputs(6422) <= (layer0_outputs(5629)) or (layer0_outputs(2733));
    outputs(6423) <= layer0_outputs(11365);
    outputs(6424) <= (layer0_outputs(5370)) or (layer0_outputs(9787));
    outputs(6425) <= (layer0_outputs(2012)) or (layer0_outputs(3834));
    outputs(6426) <= (layer0_outputs(1016)) xor (layer0_outputs(5351));
    outputs(6427) <= (layer0_outputs(8637)) and (layer0_outputs(3725));
    outputs(6428) <= (layer0_outputs(12702)) and not (layer0_outputs(8540));
    outputs(6429) <= (layer0_outputs(1385)) xor (layer0_outputs(9482));
    outputs(6430) <= not(layer0_outputs(12560));
    outputs(6431) <= layer0_outputs(7456);
    outputs(6432) <= (layer0_outputs(12547)) xor (layer0_outputs(11241));
    outputs(6433) <= (layer0_outputs(12484)) xor (layer0_outputs(7201));
    outputs(6434) <= layer0_outputs(5924);
    outputs(6435) <= layer0_outputs(3580);
    outputs(6436) <= (layer0_outputs(11322)) xor (layer0_outputs(8064));
    outputs(6437) <= not((layer0_outputs(7466)) xor (layer0_outputs(7627)));
    outputs(6438) <= (layer0_outputs(1417)) or (layer0_outputs(7248));
    outputs(6439) <= (layer0_outputs(4221)) and (layer0_outputs(9569));
    outputs(6440) <= (layer0_outputs(11228)) xor (layer0_outputs(7458));
    outputs(6441) <= not((layer0_outputs(10600)) xor (layer0_outputs(9127)));
    outputs(6442) <= not((layer0_outputs(7687)) xor (layer0_outputs(11419)));
    outputs(6443) <= not(layer0_outputs(468));
    outputs(6444) <= not((layer0_outputs(11955)) xor (layer0_outputs(11356)));
    outputs(6445) <= (layer0_outputs(1182)) xor (layer0_outputs(5808));
    outputs(6446) <= layer0_outputs(11774);
    outputs(6447) <= not(layer0_outputs(2611));
    outputs(6448) <= (layer0_outputs(6364)) xor (layer0_outputs(10415));
    outputs(6449) <= (layer0_outputs(12226)) or (layer0_outputs(8218));
    outputs(6450) <= (layer0_outputs(5905)) xor (layer0_outputs(7219));
    outputs(6451) <= not(layer0_outputs(8109)) or (layer0_outputs(7304));
    outputs(6452) <= layer0_outputs(635);
    outputs(6453) <= not(layer0_outputs(10991));
    outputs(6454) <= layer0_outputs(105);
    outputs(6455) <= layer0_outputs(5292);
    outputs(6456) <= not(layer0_outputs(2712));
    outputs(6457) <= not(layer0_outputs(10150));
    outputs(6458) <= not((layer0_outputs(2529)) xor (layer0_outputs(12387)));
    outputs(6459) <= not((layer0_outputs(246)) xor (layer0_outputs(5572)));
    outputs(6460) <= not(layer0_outputs(10869));
    outputs(6461) <= not(layer0_outputs(2284)) or (layer0_outputs(11188));
    outputs(6462) <= layer0_outputs(1513);
    outputs(6463) <= not(layer0_outputs(11136));
    outputs(6464) <= not(layer0_outputs(1496));
    outputs(6465) <= (layer0_outputs(4747)) xor (layer0_outputs(11515));
    outputs(6466) <= (layer0_outputs(6523)) xor (layer0_outputs(3112));
    outputs(6467) <= layer0_outputs(7);
    outputs(6468) <= not((layer0_outputs(8880)) xor (layer0_outputs(5076)));
    outputs(6469) <= not(layer0_outputs(1907));
    outputs(6470) <= (layer0_outputs(8213)) xor (layer0_outputs(759));
    outputs(6471) <= (layer0_outputs(5848)) xor (layer0_outputs(8607));
    outputs(6472) <= not((layer0_outputs(3078)) xor (layer0_outputs(506)));
    outputs(6473) <= not(layer0_outputs(2022));
    outputs(6474) <= not(layer0_outputs(4529));
    outputs(6475) <= not((layer0_outputs(9114)) xor (layer0_outputs(4083)));
    outputs(6476) <= not((layer0_outputs(12592)) or (layer0_outputs(12454)));
    outputs(6477) <= (layer0_outputs(4771)) xor (layer0_outputs(9416));
    outputs(6478) <= (layer0_outputs(3029)) xor (layer0_outputs(8978));
    outputs(6479) <= (layer0_outputs(1634)) xor (layer0_outputs(5872));
    outputs(6480) <= not((layer0_outputs(11517)) and (layer0_outputs(5516)));
    outputs(6481) <= not((layer0_outputs(4286)) or (layer0_outputs(698)));
    outputs(6482) <= layer0_outputs(9474);
    outputs(6483) <= not((layer0_outputs(8254)) xor (layer0_outputs(2996)));
    outputs(6484) <= layer0_outputs(5996);
    outputs(6485) <= not((layer0_outputs(2824)) or (layer0_outputs(12078)));
    outputs(6486) <= not((layer0_outputs(10785)) xor (layer0_outputs(3866)));
    outputs(6487) <= not(layer0_outputs(2000));
    outputs(6488) <= not(layer0_outputs(8771));
    outputs(6489) <= (layer0_outputs(2334)) xor (layer0_outputs(8283));
    outputs(6490) <= not((layer0_outputs(735)) xor (layer0_outputs(7040)));
    outputs(6491) <= (layer0_outputs(12752)) xor (layer0_outputs(188));
    outputs(6492) <= (layer0_outputs(2405)) xor (layer0_outputs(7074));
    outputs(6493) <= (layer0_outputs(393)) or (layer0_outputs(7818));
    outputs(6494) <= not((layer0_outputs(6449)) xor (layer0_outputs(9252)));
    outputs(6495) <= layer0_outputs(6538);
    outputs(6496) <= not((layer0_outputs(6192)) xor (layer0_outputs(12595)));
    outputs(6497) <= (layer0_outputs(7407)) and not (layer0_outputs(1668));
    outputs(6498) <= not(layer0_outputs(10309));
    outputs(6499) <= (layer0_outputs(7296)) xor (layer0_outputs(9250));
    outputs(6500) <= not((layer0_outputs(7205)) and (layer0_outputs(8557)));
    outputs(6501) <= (layer0_outputs(6476)) xor (layer0_outputs(1432));
    outputs(6502) <= not(layer0_outputs(5955));
    outputs(6503) <= (layer0_outputs(5192)) and (layer0_outputs(7767));
    outputs(6504) <= not(layer0_outputs(8632)) or (layer0_outputs(11491));
    outputs(6505) <= not(layer0_outputs(3150));
    outputs(6506) <= (layer0_outputs(12453)) xor (layer0_outputs(2192));
    outputs(6507) <= (layer0_outputs(8498)) xor (layer0_outputs(4618));
    outputs(6508) <= not((layer0_outputs(826)) xor (layer0_outputs(4008)));
    outputs(6509) <= not((layer0_outputs(564)) xor (layer0_outputs(10219)));
    outputs(6510) <= not((layer0_outputs(8773)) xor (layer0_outputs(3784)));
    outputs(6511) <= (layer0_outputs(10486)) xor (layer0_outputs(10355));
    outputs(6512) <= not((layer0_outputs(8621)) xor (layer0_outputs(7665)));
    outputs(6513) <= (layer0_outputs(3980)) and not (layer0_outputs(7003));
    outputs(6514) <= not((layer0_outputs(1941)) xor (layer0_outputs(7393)));
    outputs(6515) <= not((layer0_outputs(4390)) or (layer0_outputs(5167)));
    outputs(6516) <= not((layer0_outputs(11924)) or (layer0_outputs(4005)));
    outputs(6517) <= (layer0_outputs(5653)) xor (layer0_outputs(10246));
    outputs(6518) <= not((layer0_outputs(6740)) and (layer0_outputs(4176)));
    outputs(6519) <= (layer0_outputs(4645)) and not (layer0_outputs(9443));
    outputs(6520) <= not(layer0_outputs(4066));
    outputs(6521) <= not(layer0_outputs(3489));
    outputs(6522) <= not((layer0_outputs(2284)) xor (layer0_outputs(4776)));
    outputs(6523) <= not(layer0_outputs(6897));
    outputs(6524) <= not(layer0_outputs(6076));
    outputs(6525) <= layer0_outputs(6892);
    outputs(6526) <= not((layer0_outputs(1586)) xor (layer0_outputs(572)));
    outputs(6527) <= layer0_outputs(6810);
    outputs(6528) <= not(layer0_outputs(1636)) or (layer0_outputs(9918));
    outputs(6529) <= not((layer0_outputs(7078)) xor (layer0_outputs(2688)));
    outputs(6530) <= not((layer0_outputs(4359)) or (layer0_outputs(9634)));
    outputs(6531) <= layer0_outputs(7806);
    outputs(6532) <= not((layer0_outputs(10849)) xor (layer0_outputs(2300)));
    outputs(6533) <= not(layer0_outputs(7347)) or (layer0_outputs(8484));
    outputs(6534) <= not((layer0_outputs(5843)) xor (layer0_outputs(12680)));
    outputs(6535) <= not((layer0_outputs(7064)) and (layer0_outputs(7038)));
    outputs(6536) <= layer0_outputs(5876);
    outputs(6537) <= (layer0_outputs(12648)) xor (layer0_outputs(4286));
    outputs(6538) <= not((layer0_outputs(6071)) xor (layer0_outputs(7562)));
    outputs(6539) <= (layer0_outputs(5151)) and not (layer0_outputs(300));
    outputs(6540) <= not((layer0_outputs(8866)) xor (layer0_outputs(6209)));
    outputs(6541) <= layer0_outputs(6791);
    outputs(6542) <= not((layer0_outputs(8255)) xor (layer0_outputs(9301)));
    outputs(6543) <= layer0_outputs(5760);
    outputs(6544) <= not((layer0_outputs(1751)) or (layer0_outputs(8167)));
    outputs(6545) <= not((layer0_outputs(3924)) or (layer0_outputs(9682)));
    outputs(6546) <= layer0_outputs(8115);
    outputs(6547) <= layer0_outputs(10702);
    outputs(6548) <= (layer0_outputs(10038)) xor (layer0_outputs(9499));
    outputs(6549) <= not((layer0_outputs(2493)) and (layer0_outputs(408)));
    outputs(6550) <= not(layer0_outputs(213));
    outputs(6551) <= not((layer0_outputs(6303)) xor (layer0_outputs(6247)));
    outputs(6552) <= (layer0_outputs(3202)) xor (layer0_outputs(11612));
    outputs(6553) <= layer0_outputs(11448);
    outputs(6554) <= (layer0_outputs(124)) xor (layer0_outputs(4610));
    outputs(6555) <= (layer0_outputs(6120)) and (layer0_outputs(9807));
    outputs(6556) <= not(layer0_outputs(7630));
    outputs(6557) <= layer0_outputs(3705);
    outputs(6558) <= not(layer0_outputs(828));
    outputs(6559) <= (layer0_outputs(11923)) or (layer0_outputs(294));
    outputs(6560) <= not((layer0_outputs(629)) xor (layer0_outputs(3986)));
    outputs(6561) <= (layer0_outputs(11226)) or (layer0_outputs(5639));
    outputs(6562) <= (layer0_outputs(9105)) xor (layer0_outputs(5878));
    outputs(6563) <= layer0_outputs(3182);
    outputs(6564) <= layer0_outputs(10497);
    outputs(6565) <= layer0_outputs(5604);
    outputs(6566) <= (layer0_outputs(2003)) and not (layer0_outputs(331));
    outputs(6567) <= not((layer0_outputs(12596)) xor (layer0_outputs(12764)));
    outputs(6568) <= not(layer0_outputs(9483));
    outputs(6569) <= (layer0_outputs(5407)) xor (layer0_outputs(1724));
    outputs(6570) <= not((layer0_outputs(552)) xor (layer0_outputs(12592)));
    outputs(6571) <= not((layer0_outputs(4517)) xor (layer0_outputs(5948)));
    outputs(6572) <= not((layer0_outputs(8111)) or (layer0_outputs(1173)));
    outputs(6573) <= layer0_outputs(8928);
    outputs(6574) <= not(layer0_outputs(3226));
    outputs(6575) <= (layer0_outputs(3210)) xor (layer0_outputs(6824));
    outputs(6576) <= not((layer0_outputs(1027)) xor (layer0_outputs(1608)));
    outputs(6577) <= not((layer0_outputs(10979)) xor (layer0_outputs(9068)));
    outputs(6578) <= (layer0_outputs(3782)) xor (layer0_outputs(4339));
    outputs(6579) <= (layer0_outputs(9740)) and not (layer0_outputs(8577));
    outputs(6580) <= layer0_outputs(6835);
    outputs(6581) <= layer0_outputs(3677);
    outputs(6582) <= not(layer0_outputs(3201)) or (layer0_outputs(1667));
    outputs(6583) <= (layer0_outputs(3643)) xor (layer0_outputs(1228));
    outputs(6584) <= not(layer0_outputs(10054)) or (layer0_outputs(10639));
    outputs(6585) <= not((layer0_outputs(2437)) xor (layer0_outputs(3324)));
    outputs(6586) <= layer0_outputs(5507);
    outputs(6587) <= not(layer0_outputs(3965)) or (layer0_outputs(12023));
    outputs(6588) <= not(layer0_outputs(6040)) or (layer0_outputs(3504));
    outputs(6589) <= not((layer0_outputs(12417)) xor (layer0_outputs(2723)));
    outputs(6590) <= layer0_outputs(11015);
    outputs(6591) <= not((layer0_outputs(2419)) and (layer0_outputs(5035)));
    outputs(6592) <= layer0_outputs(5123);
    outputs(6593) <= not((layer0_outputs(12297)) xor (layer0_outputs(12259)));
    outputs(6594) <= not(layer0_outputs(4214)) or (layer0_outputs(4695));
    outputs(6595) <= not((layer0_outputs(3624)) xor (layer0_outputs(9123)));
    outputs(6596) <= not((layer0_outputs(9534)) xor (layer0_outputs(6981)));
    outputs(6597) <= not(layer0_outputs(1640));
    outputs(6598) <= not((layer0_outputs(1595)) xor (layer0_outputs(11909)));
    outputs(6599) <= (layer0_outputs(6942)) xor (layer0_outputs(2567));
    outputs(6600) <= (layer0_outputs(4611)) xor (layer0_outputs(7155));
    outputs(6601) <= layer0_outputs(1558);
    outputs(6602) <= layer0_outputs(7380);
    outputs(6603) <= not((layer0_outputs(2185)) xor (layer0_outputs(11253)));
    outputs(6604) <= (layer0_outputs(4034)) xor (layer0_outputs(6849));
    outputs(6605) <= (layer0_outputs(6720)) xor (layer0_outputs(6662));
    outputs(6606) <= not(layer0_outputs(4011));
    outputs(6607) <= not((layer0_outputs(4164)) xor (layer0_outputs(11805)));
    outputs(6608) <= not((layer0_outputs(6091)) xor (layer0_outputs(3586)));
    outputs(6609) <= layer0_outputs(2204);
    outputs(6610) <= not(layer0_outputs(3936));
    outputs(6611) <= (layer0_outputs(4392)) and not (layer0_outputs(4579));
    outputs(6612) <= layer0_outputs(723);
    outputs(6613) <= not(layer0_outputs(12094));
    outputs(6614) <= not(layer0_outputs(9335));
    outputs(6615) <= not((layer0_outputs(8134)) xor (layer0_outputs(4555)));
    outputs(6616) <= (layer0_outputs(8142)) xor (layer0_outputs(11006));
    outputs(6617) <= (layer0_outputs(10942)) xor (layer0_outputs(11618));
    outputs(6618) <= not((layer0_outputs(2394)) xor (layer0_outputs(2205)));
    outputs(6619) <= not(layer0_outputs(7781));
    outputs(6620) <= not(layer0_outputs(6492));
    outputs(6621) <= not((layer0_outputs(4349)) or (layer0_outputs(11394)));
    outputs(6622) <= not(layer0_outputs(3701));
    outputs(6623) <= (layer0_outputs(11042)) xor (layer0_outputs(11607));
    outputs(6624) <= layer0_outputs(11274);
    outputs(6625) <= (layer0_outputs(4109)) and (layer0_outputs(12040));
    outputs(6626) <= not((layer0_outputs(11756)) xor (layer0_outputs(2977)));
    outputs(6627) <= not(layer0_outputs(10816));
    outputs(6628) <= (layer0_outputs(3533)) xor (layer0_outputs(9070));
    outputs(6629) <= (layer0_outputs(2578)) xor (layer0_outputs(9709));
    outputs(6630) <= not(layer0_outputs(6376));
    outputs(6631) <= (layer0_outputs(3911)) xor (layer0_outputs(10377));
    outputs(6632) <= (layer0_outputs(2937)) xor (layer0_outputs(6585));
    outputs(6633) <= not((layer0_outputs(256)) or (layer0_outputs(10473)));
    outputs(6634) <= not((layer0_outputs(5740)) xor (layer0_outputs(1998)));
    outputs(6635) <= layer0_outputs(5830);
    outputs(6636) <= not(layer0_outputs(2687));
    outputs(6637) <= not((layer0_outputs(9604)) xor (layer0_outputs(9590)));
    outputs(6638) <= (layer0_outputs(8865)) and not (layer0_outputs(3323));
    outputs(6639) <= not((layer0_outputs(1581)) and (layer0_outputs(11636)));
    outputs(6640) <= (layer0_outputs(8643)) xor (layer0_outputs(9080));
    outputs(6641) <= layer0_outputs(3356);
    outputs(6642) <= not(layer0_outputs(7234)) or (layer0_outputs(1221));
    outputs(6643) <= (layer0_outputs(4441)) xor (layer0_outputs(7282));
    outputs(6644) <= (layer0_outputs(5950)) xor (layer0_outputs(9222));
    outputs(6645) <= not(layer0_outputs(2892));
    outputs(6646) <= not((layer0_outputs(881)) xor (layer0_outputs(1746)));
    outputs(6647) <= layer0_outputs(5854);
    outputs(6648) <= not(layer0_outputs(1035));
    outputs(6649) <= not(layer0_outputs(10009));
    outputs(6650) <= (layer0_outputs(9909)) xor (layer0_outputs(4991));
    outputs(6651) <= not((layer0_outputs(4848)) xor (layer0_outputs(2529)));
    outputs(6652) <= not(layer0_outputs(10618));
    outputs(6653) <= layer0_outputs(9978);
    outputs(6654) <= (layer0_outputs(5806)) xor (layer0_outputs(1808));
    outputs(6655) <= (layer0_outputs(2035)) xor (layer0_outputs(12740));
    outputs(6656) <= layer0_outputs(11584);
    outputs(6657) <= not((layer0_outputs(3448)) xor (layer0_outputs(5284)));
    outputs(6658) <= not((layer0_outputs(9515)) and (layer0_outputs(427)));
    outputs(6659) <= not(layer0_outputs(3120));
    outputs(6660) <= not(layer0_outputs(4465));
    outputs(6661) <= not((layer0_outputs(10792)) xor (layer0_outputs(1793)));
    outputs(6662) <= not(layer0_outputs(11834)) or (layer0_outputs(10057));
    outputs(6663) <= not((layer0_outputs(6873)) or (layer0_outputs(1117)));
    outputs(6664) <= not((layer0_outputs(7907)) and (layer0_outputs(3398)));
    outputs(6665) <= layer0_outputs(9826);
    outputs(6666) <= (layer0_outputs(2464)) and (layer0_outputs(1673));
    outputs(6667) <= (layer0_outputs(828)) xor (layer0_outputs(8715));
    outputs(6668) <= not(layer0_outputs(11777)) or (layer0_outputs(7250));
    outputs(6669) <= (layer0_outputs(11403)) xor (layer0_outputs(10736));
    outputs(6670) <= (layer0_outputs(6548)) and not (layer0_outputs(10431));
    outputs(6671) <= layer0_outputs(6458);
    outputs(6672) <= not((layer0_outputs(7103)) xor (layer0_outputs(2403)));
    outputs(6673) <= not(layer0_outputs(6895));
    outputs(6674) <= not(layer0_outputs(6407));
    outputs(6675) <= not((layer0_outputs(5951)) xor (layer0_outputs(11694)));
    outputs(6676) <= not(layer0_outputs(8489));
    outputs(6677) <= layer0_outputs(3419);
    outputs(6678) <= not((layer0_outputs(8822)) or (layer0_outputs(4030)));
    outputs(6679) <= not(layer0_outputs(761));
    outputs(6680) <= not((layer0_outputs(1779)) xor (layer0_outputs(1512)));
    outputs(6681) <= not(layer0_outputs(7824));
    outputs(6682) <= (layer0_outputs(8064)) and (layer0_outputs(4092));
    outputs(6683) <= not(layer0_outputs(4828));
    outputs(6684) <= not(layer0_outputs(10395));
    outputs(6685) <= not(layer0_outputs(579)) or (layer0_outputs(1394));
    outputs(6686) <= not((layer0_outputs(1580)) or (layer0_outputs(11285)));
    outputs(6687) <= not((layer0_outputs(8883)) and (layer0_outputs(8967)));
    outputs(6688) <= not(layer0_outputs(4626));
    outputs(6689) <= (layer0_outputs(12228)) xor (layer0_outputs(9091));
    outputs(6690) <= not((layer0_outputs(9721)) xor (layer0_outputs(8302)));
    outputs(6691) <= (layer0_outputs(6890)) xor (layer0_outputs(7281));
    outputs(6692) <= layer0_outputs(4401);
    outputs(6693) <= layer0_outputs(6110);
    outputs(6694) <= not(layer0_outputs(11589));
    outputs(6695) <= not((layer0_outputs(8342)) xor (layer0_outputs(1457)));
    outputs(6696) <= not((layer0_outputs(10404)) xor (layer0_outputs(618)));
    outputs(6697) <= not((layer0_outputs(10477)) xor (layer0_outputs(3436)));
    outputs(6698) <= not(layer0_outputs(1918));
    outputs(6699) <= layer0_outputs(7606);
    outputs(6700) <= not((layer0_outputs(3743)) xor (layer0_outputs(2930)));
    outputs(6701) <= not(layer0_outputs(7945));
    outputs(6702) <= (layer0_outputs(11700)) xor (layer0_outputs(12004));
    outputs(6703) <= not((layer0_outputs(4630)) and (layer0_outputs(619)));
    outputs(6704) <= layer0_outputs(10085);
    outputs(6705) <= not((layer0_outputs(12419)) xor (layer0_outputs(11130)));
    outputs(6706) <= (layer0_outputs(1260)) xor (layer0_outputs(10461));
    outputs(6707) <= (layer0_outputs(9792)) or (layer0_outputs(894));
    outputs(6708) <= (layer0_outputs(6214)) xor (layer0_outputs(7945));
    outputs(6709) <= (layer0_outputs(2971)) and not (layer0_outputs(3840));
    outputs(6710) <= not(layer0_outputs(10056)) or (layer0_outputs(6181));
    outputs(6711) <= layer0_outputs(6994);
    outputs(6712) <= not((layer0_outputs(11454)) and (layer0_outputs(804)));
    outputs(6713) <= not(layer0_outputs(4043));
    outputs(6714) <= (layer0_outputs(11272)) or (layer0_outputs(9194));
    outputs(6715) <= (layer0_outputs(9702)) and not (layer0_outputs(5813));
    outputs(6716) <= not(layer0_outputs(2452));
    outputs(6717) <= not((layer0_outputs(72)) xor (layer0_outputs(5171)));
    outputs(6718) <= (layer0_outputs(12635)) xor (layer0_outputs(11193));
    outputs(6719) <= (layer0_outputs(12485)) and not (layer0_outputs(5094));
    outputs(6720) <= not(layer0_outputs(11927));
    outputs(6721) <= not((layer0_outputs(8752)) or (layer0_outputs(10240)));
    outputs(6722) <= not((layer0_outputs(4635)) xor (layer0_outputs(9929)));
    outputs(6723) <= not((layer0_outputs(6417)) xor (layer0_outputs(3767)));
    outputs(6724) <= not(layer0_outputs(1390)) or (layer0_outputs(2514));
    outputs(6725) <= layer0_outputs(5942);
    outputs(6726) <= (layer0_outputs(8525)) xor (layer0_outputs(1457));
    outputs(6727) <= (layer0_outputs(4973)) xor (layer0_outputs(10294));
    outputs(6728) <= (layer0_outputs(3713)) and (layer0_outputs(7139));
    outputs(6729) <= not(layer0_outputs(977));
    outputs(6730) <= not(layer0_outputs(5783));
    outputs(6731) <= (layer0_outputs(6987)) xor (layer0_outputs(11043));
    outputs(6732) <= not((layer0_outputs(11747)) xor (layer0_outputs(11658)));
    outputs(6733) <= (layer0_outputs(9682)) xor (layer0_outputs(9332));
    outputs(6734) <= (layer0_outputs(12443)) and not (layer0_outputs(3661));
    outputs(6735) <= not(layer0_outputs(9407));
    outputs(6736) <= not((layer0_outputs(4281)) xor (layer0_outputs(10563)));
    outputs(6737) <= not((layer0_outputs(6951)) xor (layer0_outputs(7426)));
    outputs(6738) <= layer0_outputs(2002);
    outputs(6739) <= (layer0_outputs(3647)) xor (layer0_outputs(11460));
    outputs(6740) <= (layer0_outputs(1394)) xor (layer0_outputs(9943));
    outputs(6741) <= not((layer0_outputs(10546)) xor (layer0_outputs(6971)));
    outputs(6742) <= not((layer0_outputs(3209)) and (layer0_outputs(7048)));
    outputs(6743) <= not(layer0_outputs(2790)) or (layer0_outputs(6078));
    outputs(6744) <= not((layer0_outputs(5933)) xor (layer0_outputs(2458)));
    outputs(6745) <= (layer0_outputs(7828)) xor (layer0_outputs(12390));
    outputs(6746) <= layer0_outputs(1138);
    outputs(6747) <= layer0_outputs(11816);
    outputs(6748) <= (layer0_outputs(5104)) and not (layer0_outputs(7133));
    outputs(6749) <= layer0_outputs(11845);
    outputs(6750) <= not((layer0_outputs(3341)) or (layer0_outputs(8102)));
    outputs(6751) <= not((layer0_outputs(7360)) xor (layer0_outputs(1202)));
    outputs(6752) <= not((layer0_outputs(9571)) xor (layer0_outputs(4721)));
    outputs(6753) <= not(layer0_outputs(7571));
    outputs(6754) <= not((layer0_outputs(12290)) xor (layer0_outputs(33)));
    outputs(6755) <= (layer0_outputs(2303)) xor (layer0_outputs(12722));
    outputs(6756) <= not(layer0_outputs(1465)) or (layer0_outputs(10866));
    outputs(6757) <= not((layer0_outputs(4077)) xor (layer0_outputs(3130)));
    outputs(6758) <= not((layer0_outputs(1094)) and (layer0_outputs(1967)));
    outputs(6759) <= layer0_outputs(8046);
    outputs(6760) <= layer0_outputs(704);
    outputs(6761) <= not(layer0_outputs(9146));
    outputs(6762) <= layer0_outputs(4292);
    outputs(6763) <= not(layer0_outputs(4725)) or (layer0_outputs(5946));
    outputs(6764) <= (layer0_outputs(497)) xor (layer0_outputs(9754));
    outputs(6765) <= (layer0_outputs(12586)) xor (layer0_outputs(10291));
    outputs(6766) <= (layer0_outputs(9489)) xor (layer0_outputs(12064));
    outputs(6767) <= not(layer0_outputs(10106));
    outputs(6768) <= (layer0_outputs(11871)) xor (layer0_outputs(9015));
    outputs(6769) <= layer0_outputs(10219);
    outputs(6770) <= (layer0_outputs(12086)) or (layer0_outputs(9428));
    outputs(6771) <= layer0_outputs(6998);
    outputs(6772) <= not((layer0_outputs(8342)) xor (layer0_outputs(7233)));
    outputs(6773) <= not(layer0_outputs(944));
    outputs(6774) <= layer0_outputs(11640);
    outputs(6775) <= not((layer0_outputs(5435)) xor (layer0_outputs(3841)));
    outputs(6776) <= layer0_outputs(11667);
    outputs(6777) <= layer0_outputs(580);
    outputs(6778) <= layer0_outputs(4523);
    outputs(6779) <= layer0_outputs(11751);
    outputs(6780) <= not((layer0_outputs(8170)) xor (layer0_outputs(6387)));
    outputs(6781) <= not((layer0_outputs(1522)) xor (layer0_outputs(5566)));
    outputs(6782) <= not((layer0_outputs(6551)) xor (layer0_outputs(10545)));
    outputs(6783) <= not((layer0_outputs(10505)) xor (layer0_outputs(4191)));
    outputs(6784) <= layer0_outputs(12647);
    outputs(6785) <= layer0_outputs(12006);
    outputs(6786) <= layer0_outputs(3989);
    outputs(6787) <= not((layer0_outputs(9157)) and (layer0_outputs(8760)));
    outputs(6788) <= layer0_outputs(5780);
    outputs(6789) <= not(layer0_outputs(11706));
    outputs(6790) <= not(layer0_outputs(17)) or (layer0_outputs(10411));
    outputs(6791) <= (layer0_outputs(4881)) and not (layer0_outputs(2214));
    outputs(6792) <= (layer0_outputs(12273)) xor (layer0_outputs(702));
    outputs(6793) <= (layer0_outputs(1054)) xor (layer0_outputs(6967));
    outputs(6794) <= (layer0_outputs(7258)) and not (layer0_outputs(8966));
    outputs(6795) <= layer0_outputs(4515);
    outputs(6796) <= (layer0_outputs(1421)) xor (layer0_outputs(8446));
    outputs(6797) <= layer0_outputs(11895);
    outputs(6798) <= layer0_outputs(11251);
    outputs(6799) <= not(layer0_outputs(6529)) or (layer0_outputs(7081));
    outputs(6800) <= not(layer0_outputs(4530));
    outputs(6801) <= not((layer0_outputs(6208)) and (layer0_outputs(9508)));
    outputs(6802) <= not(layer0_outputs(4431));
    outputs(6803) <= not(layer0_outputs(10534));
    outputs(6804) <= not((layer0_outputs(7389)) and (layer0_outputs(7126)));
    outputs(6805) <= not((layer0_outputs(9450)) and (layer0_outputs(11030)));
    outputs(6806) <= not((layer0_outputs(8958)) xor (layer0_outputs(904)));
    outputs(6807) <= not(layer0_outputs(2355));
    outputs(6808) <= (layer0_outputs(11263)) xor (layer0_outputs(722));
    outputs(6809) <= not((layer0_outputs(6568)) xor (layer0_outputs(9018)));
    outputs(6810) <= not(layer0_outputs(10402));
    outputs(6811) <= (layer0_outputs(4428)) and (layer0_outputs(6905));
    outputs(6812) <= not(layer0_outputs(8584)) or (layer0_outputs(4410));
    outputs(6813) <= not(layer0_outputs(8557));
    outputs(6814) <= not((layer0_outputs(8810)) xor (layer0_outputs(11264)));
    outputs(6815) <= (layer0_outputs(88)) xor (layer0_outputs(4458));
    outputs(6816) <= layer0_outputs(223);
    outputs(6817) <= not((layer0_outputs(5126)) or (layer0_outputs(7044)));
    outputs(6818) <= not((layer0_outputs(7465)) xor (layer0_outputs(8516)));
    outputs(6819) <= not((layer0_outputs(5593)) xor (layer0_outputs(86)));
    outputs(6820) <= (layer0_outputs(9148)) xor (layer0_outputs(9632));
    outputs(6821) <= not((layer0_outputs(9610)) xor (layer0_outputs(7318)));
    outputs(6822) <= (layer0_outputs(12)) xor (layer0_outputs(3970));
    outputs(6823) <= (layer0_outputs(6145)) and (layer0_outputs(5871));
    outputs(6824) <= not((layer0_outputs(545)) xor (layer0_outputs(11204)));
    outputs(6825) <= layer0_outputs(7601);
    outputs(6826) <= layer0_outputs(9063);
    outputs(6827) <= not((layer0_outputs(3814)) xor (layer0_outputs(1962)));
    outputs(6828) <= not((layer0_outputs(7460)) xor (layer0_outputs(6149)));
    outputs(6829) <= not(layer0_outputs(7285));
    outputs(6830) <= (layer0_outputs(11433)) xor (layer0_outputs(8562));
    outputs(6831) <= (layer0_outputs(1423)) xor (layer0_outputs(7298));
    outputs(6832) <= not(layer0_outputs(965));
    outputs(6833) <= layer0_outputs(4398);
    outputs(6834) <= not(layer0_outputs(11028));
    outputs(6835) <= not((layer0_outputs(6576)) and (layer0_outputs(5173)));
    outputs(6836) <= not(layer0_outputs(11100)) or (layer0_outputs(2243));
    outputs(6837) <= not((layer0_outputs(3652)) xor (layer0_outputs(12207)));
    outputs(6838) <= (layer0_outputs(11850)) xor (layer0_outputs(443));
    outputs(6839) <= layer0_outputs(4770);
    outputs(6840) <= layer0_outputs(11780);
    outputs(6841) <= (layer0_outputs(8251)) or (layer0_outputs(5311));
    outputs(6842) <= layer0_outputs(7541);
    outputs(6843) <= not(layer0_outputs(3039)) or (layer0_outputs(2081));
    outputs(6844) <= not(layer0_outputs(8572));
    outputs(6845) <= not(layer0_outputs(5246));
    outputs(6846) <= not(layer0_outputs(8544));
    outputs(6847) <= not((layer0_outputs(7305)) xor (layer0_outputs(9359)));
    outputs(6848) <= not((layer0_outputs(4802)) xor (layer0_outputs(8301)));
    outputs(6849) <= layer0_outputs(6540);
    outputs(6850) <= layer0_outputs(3020);
    outputs(6851) <= not((layer0_outputs(5041)) xor (layer0_outputs(7529)));
    outputs(6852) <= layer0_outputs(4292);
    outputs(6853) <= not(layer0_outputs(3794)) or (layer0_outputs(7762));
    outputs(6854) <= not((layer0_outputs(5097)) xor (layer0_outputs(3510)));
    outputs(6855) <= (layer0_outputs(8431)) xor (layer0_outputs(12217));
    outputs(6856) <= (layer0_outputs(11120)) xor (layer0_outputs(2964));
    outputs(6857) <= not((layer0_outputs(12114)) xor (layer0_outputs(6237)));
    outputs(6858) <= layer0_outputs(6354);
    outputs(6859) <= not(layer0_outputs(6326));
    outputs(6860) <= (layer0_outputs(8259)) and not (layer0_outputs(10893));
    outputs(6861) <= layer0_outputs(1216);
    outputs(6862) <= not(layer0_outputs(2495));
    outputs(6863) <= not((layer0_outputs(3826)) xor (layer0_outputs(9822)));
    outputs(6864) <= not(layer0_outputs(4989));
    outputs(6865) <= layer0_outputs(7829);
    outputs(6866) <= not((layer0_outputs(3167)) xor (layer0_outputs(9683)));
    outputs(6867) <= layer0_outputs(3183);
    outputs(6868) <= not(layer0_outputs(10158));
    outputs(6869) <= (layer0_outputs(7957)) or (layer0_outputs(5107));
    outputs(6870) <= not(layer0_outputs(2344));
    outputs(6871) <= not(layer0_outputs(1110)) or (layer0_outputs(10079));
    outputs(6872) <= (layer0_outputs(9889)) xor (layer0_outputs(2371));
    outputs(6873) <= not((layer0_outputs(2850)) xor (layer0_outputs(2554)));
    outputs(6874) <= (layer0_outputs(432)) and not (layer0_outputs(3372));
    outputs(6875) <= not((layer0_outputs(795)) xor (layer0_outputs(10192)));
    outputs(6876) <= not(layer0_outputs(2452));
    outputs(6877) <= not((layer0_outputs(621)) xor (layer0_outputs(10390)));
    outputs(6878) <= layer0_outputs(454);
    outputs(6879) <= layer0_outputs(7697);
    outputs(6880) <= layer0_outputs(843);
    outputs(6881) <= layer0_outputs(1238);
    outputs(6882) <= layer0_outputs(1663);
    outputs(6883) <= not((layer0_outputs(8239)) xor (layer0_outputs(6983)));
    outputs(6884) <= (layer0_outputs(1029)) and (layer0_outputs(1591));
    outputs(6885) <= not(layer0_outputs(7978));
    outputs(6886) <= layer0_outputs(9240);
    outputs(6887) <= not((layer0_outputs(3279)) xor (layer0_outputs(3123)));
    outputs(6888) <= not((layer0_outputs(10203)) xor (layer0_outputs(1024)));
    outputs(6889) <= (layer0_outputs(6748)) or (layer0_outputs(4466));
    outputs(6890) <= (layer0_outputs(4201)) xor (layer0_outputs(1871));
    outputs(6891) <= not(layer0_outputs(11190));
    outputs(6892) <= not(layer0_outputs(4199)) or (layer0_outputs(9801));
    outputs(6893) <= not((layer0_outputs(10027)) xor (layer0_outputs(4994)));
    outputs(6894) <= not(layer0_outputs(5371));
    outputs(6895) <= (layer0_outputs(1822)) and not (layer0_outputs(3983));
    outputs(6896) <= not((layer0_outputs(6965)) xor (layer0_outputs(9014)));
    outputs(6897) <= layer0_outputs(325);
    outputs(6898) <= (layer0_outputs(2990)) xor (layer0_outputs(8878));
    outputs(6899) <= not((layer0_outputs(10439)) xor (layer0_outputs(3641)));
    outputs(6900) <= (layer0_outputs(12072)) xor (layer0_outputs(5344));
    outputs(6901) <= (layer0_outputs(5379)) xor (layer0_outputs(11337));
    outputs(6902) <= layer0_outputs(2929);
    outputs(6903) <= not((layer0_outputs(2599)) or (layer0_outputs(10509)));
    outputs(6904) <= (layer0_outputs(711)) xor (layer0_outputs(153));
    outputs(6905) <= (layer0_outputs(11445)) xor (layer0_outputs(5616));
    outputs(6906) <= layer0_outputs(5932);
    outputs(6907) <= not((layer0_outputs(4203)) or (layer0_outputs(9791)));
    outputs(6908) <= not((layer0_outputs(9835)) and (layer0_outputs(11088)));
    outputs(6909) <= not((layer0_outputs(1243)) or (layer0_outputs(4769)));
    outputs(6910) <= layer0_outputs(3825);
    outputs(6911) <= not(layer0_outputs(3053));
    outputs(6912) <= not((layer0_outputs(11111)) xor (layer0_outputs(2384)));
    outputs(6913) <= (layer0_outputs(1730)) xor (layer0_outputs(12432));
    outputs(6914) <= not((layer0_outputs(2934)) xor (layer0_outputs(4455)));
    outputs(6915) <= not((layer0_outputs(9201)) and (layer0_outputs(4197)));
    outputs(6916) <= layer0_outputs(4382);
    outputs(6917) <= not(layer0_outputs(10466));
    outputs(6918) <= not(layer0_outputs(9628));
    outputs(6919) <= (layer0_outputs(7494)) xor (layer0_outputs(9271));
    outputs(6920) <= not((layer0_outputs(5209)) xor (layer0_outputs(3651)));
    outputs(6921) <= not((layer0_outputs(3420)) xor (layer0_outputs(12326)));
    outputs(6922) <= not((layer0_outputs(1547)) xor (layer0_outputs(10333)));
    outputs(6923) <= not(layer0_outputs(12302));
    outputs(6924) <= (layer0_outputs(3287)) or (layer0_outputs(9513));
    outputs(6925) <= (layer0_outputs(11996)) and (layer0_outputs(1729));
    outputs(6926) <= layer0_outputs(5171);
    outputs(6927) <= (layer0_outputs(1127)) xor (layer0_outputs(3105));
    outputs(6928) <= not((layer0_outputs(8822)) or (layer0_outputs(7060)));
    outputs(6929) <= (layer0_outputs(1644)) and not (layer0_outputs(4456));
    outputs(6930) <= not(layer0_outputs(9411));
    outputs(6931) <= not(layer0_outputs(3974));
    outputs(6932) <= not(layer0_outputs(12124));
    outputs(6933) <= (layer0_outputs(11246)) and (layer0_outputs(3085));
    outputs(6934) <= layer0_outputs(8078);
    outputs(6935) <= (layer0_outputs(11768)) and not (layer0_outputs(10250));
    outputs(6936) <= (layer0_outputs(3103)) xor (layer0_outputs(5571));
    outputs(6937) <= not((layer0_outputs(5486)) xor (layer0_outputs(7746)));
    outputs(6938) <= (layer0_outputs(5529)) xor (layer0_outputs(1693));
    outputs(6939) <= (layer0_outputs(7785)) xor (layer0_outputs(3230));
    outputs(6940) <= (layer0_outputs(12500)) xor (layer0_outputs(3503));
    outputs(6941) <= not((layer0_outputs(7247)) xor (layer0_outputs(1010)));
    outputs(6942) <= not((layer0_outputs(3413)) and (layer0_outputs(8931)));
    outputs(6943) <= (layer0_outputs(8139)) xor (layer0_outputs(5037));
    outputs(6944) <= not(layer0_outputs(1366));
    outputs(6945) <= not(layer0_outputs(4815));
    outputs(6946) <= not(layer0_outputs(4452));
    outputs(6947) <= not(layer0_outputs(9553));
    outputs(6948) <= not(layer0_outputs(10701)) or (layer0_outputs(9726));
    outputs(6949) <= not((layer0_outputs(10838)) xor (layer0_outputs(1574)));
    outputs(6950) <= not(layer0_outputs(7381));
    outputs(6951) <= (layer0_outputs(3720)) and not (layer0_outputs(3792));
    outputs(6952) <= not(layer0_outputs(8008));
    outputs(6953) <= (layer0_outputs(5617)) xor (layer0_outputs(9684));
    outputs(6954) <= not((layer0_outputs(3277)) xor (layer0_outputs(9790)));
    outputs(6955) <= not((layer0_outputs(12700)) xor (layer0_outputs(8552)));
    outputs(6956) <= layer0_outputs(10344);
    outputs(6957) <= (layer0_outputs(4090)) xor (layer0_outputs(5557));
    outputs(6958) <= not(layer0_outputs(3714)) or (layer0_outputs(2453));
    outputs(6959) <= not(layer0_outputs(9890)) or (layer0_outputs(382));
    outputs(6960) <= not((layer0_outputs(8251)) xor (layer0_outputs(8717)));
    outputs(6961) <= not(layer0_outputs(7659));
    outputs(6962) <= layer0_outputs(8223);
    outputs(6963) <= layer0_outputs(2907);
    outputs(6964) <= not((layer0_outputs(4150)) or (layer0_outputs(637)));
    outputs(6965) <= not(layer0_outputs(4063));
    outputs(6966) <= not((layer0_outputs(35)) xor (layer0_outputs(1381)));
    outputs(6967) <= layer0_outputs(10590);
    outputs(6968) <= not((layer0_outputs(12708)) xor (layer0_outputs(2667)));
    outputs(6969) <= not((layer0_outputs(6627)) xor (layer0_outputs(10432)));
    outputs(6970) <= not(layer0_outputs(12197));
    outputs(6971) <= layer0_outputs(12280);
    outputs(6972) <= not((layer0_outputs(5797)) xor (layer0_outputs(11404)));
    outputs(6973) <= not((layer0_outputs(3614)) xor (layer0_outputs(7620)));
    outputs(6974) <= not(layer0_outputs(2239));
    outputs(6975) <= (layer0_outputs(12086)) or (layer0_outputs(8957));
    outputs(6976) <= (layer0_outputs(2238)) xor (layer0_outputs(9972));
    outputs(6977) <= not(layer0_outputs(1531));
    outputs(6978) <= (layer0_outputs(11435)) xor (layer0_outputs(2079));
    outputs(6979) <= layer0_outputs(11364);
    outputs(6980) <= (layer0_outputs(4169)) and (layer0_outputs(1608));
    outputs(6981) <= layer0_outputs(1);
    outputs(6982) <= not(layer0_outputs(7062));
    outputs(6983) <= not((layer0_outputs(6144)) xor (layer0_outputs(12721)));
    outputs(6984) <= (layer0_outputs(10696)) xor (layer0_outputs(5691));
    outputs(6985) <= layer0_outputs(1906);
    outputs(6986) <= not((layer0_outputs(6087)) xor (layer0_outputs(1438)));
    outputs(6987) <= not((layer0_outputs(4700)) xor (layer0_outputs(7402)));
    outputs(6988) <= not(layer0_outputs(9181));
    outputs(6989) <= not(layer0_outputs(3766));
    outputs(6990) <= (layer0_outputs(5068)) and (layer0_outputs(4623));
    outputs(6991) <= not(layer0_outputs(8755));
    outputs(6992) <= layer0_outputs(11685);
    outputs(6993) <= (layer0_outputs(5095)) xor (layer0_outputs(862));
    outputs(6994) <= (layer0_outputs(6777)) and not (layer0_outputs(7538));
    outputs(6995) <= not((layer0_outputs(8911)) xor (layer0_outputs(10817)));
    outputs(6996) <= (layer0_outputs(10131)) xor (layer0_outputs(8949));
    outputs(6997) <= not(layer0_outputs(7069));
    outputs(6998) <= (layer0_outputs(6064)) xor (layer0_outputs(8975));
    outputs(6999) <= not((layer0_outputs(9636)) xor (layer0_outputs(2018)));
    outputs(7000) <= not((layer0_outputs(11019)) xor (layer0_outputs(7868)));
    outputs(7001) <= (layer0_outputs(8352)) xor (layer0_outputs(8709));
    outputs(7002) <= layer0_outputs(6620);
    outputs(7003) <= layer0_outputs(11354);
    outputs(7004) <= (layer0_outputs(4740)) xor (layer0_outputs(3027));
    outputs(7005) <= not((layer0_outputs(6185)) and (layer0_outputs(7576)));
    outputs(7006) <= not(layer0_outputs(10502));
    outputs(7007) <= (layer0_outputs(721)) xor (layer0_outputs(1013));
    outputs(7008) <= not(layer0_outputs(12309));
    outputs(7009) <= not(layer0_outputs(12166));
    outputs(7010) <= not((layer0_outputs(4437)) or (layer0_outputs(5205)));
    outputs(7011) <= (layer0_outputs(11935)) xor (layer0_outputs(11582));
    outputs(7012) <= not(layer0_outputs(2702));
    outputs(7013) <= layer0_outputs(6990);
    outputs(7014) <= not(layer0_outputs(11542)) or (layer0_outputs(9815));
    outputs(7015) <= not((layer0_outputs(7598)) or (layer0_outputs(4918)));
    outputs(7016) <= not(layer0_outputs(548));
    outputs(7017) <= layer0_outputs(5195);
    outputs(7018) <= (layer0_outputs(11303)) and (layer0_outputs(5335));
    outputs(7019) <= not((layer0_outputs(1998)) xor (layer0_outputs(11307)));
    outputs(7020) <= (layer0_outputs(3750)) xor (layer0_outputs(1734));
    outputs(7021) <= layer0_outputs(3217);
    outputs(7022) <= layer0_outputs(2395);
    outputs(7023) <= not(layer0_outputs(8548));
    outputs(7024) <= not(layer0_outputs(4336));
    outputs(7025) <= not(layer0_outputs(9073)) or (layer0_outputs(1930));
    outputs(7026) <= (layer0_outputs(3512)) xor (layer0_outputs(1986));
    outputs(7027) <= not((layer0_outputs(4015)) xor (layer0_outputs(11430)));
    outputs(7028) <= (layer0_outputs(520)) and (layer0_outputs(11451));
    outputs(7029) <= layer0_outputs(11116);
    outputs(7030) <= not((layer0_outputs(1369)) xor (layer0_outputs(8402)));
    outputs(7031) <= layer0_outputs(12646);
    outputs(7032) <= not(layer0_outputs(11629));
    outputs(7033) <= layer0_outputs(5244);
    outputs(7034) <= not((layer0_outputs(2188)) xor (layer0_outputs(11175)));
    outputs(7035) <= (layer0_outputs(12787)) and (layer0_outputs(5330));
    outputs(7036) <= not((layer0_outputs(10786)) xor (layer0_outputs(7004)));
    outputs(7037) <= not(layer0_outputs(1392));
    outputs(7038) <= not((layer0_outputs(8063)) xor (layer0_outputs(2293)));
    outputs(7039) <= not(layer0_outputs(7543));
    outputs(7040) <= not(layer0_outputs(6359));
    outputs(7041) <= not(layer0_outputs(11332));
    outputs(7042) <= not((layer0_outputs(6564)) xor (layer0_outputs(5510)));
    outputs(7043) <= (layer0_outputs(5451)) xor (layer0_outputs(7855));
    outputs(7044) <= not((layer0_outputs(6732)) xor (layer0_outputs(697)));
    outputs(7045) <= layer0_outputs(5300);
    outputs(7046) <= layer0_outputs(2656);
    outputs(7047) <= (layer0_outputs(4778)) and not (layer0_outputs(5682));
    outputs(7048) <= layer0_outputs(2942);
    outputs(7049) <= not((layer0_outputs(7685)) xor (layer0_outputs(2249)));
    outputs(7050) <= not(layer0_outputs(12408));
    outputs(7051) <= layer0_outputs(12531);
    outputs(7052) <= not((layer0_outputs(11791)) xor (layer0_outputs(10432)));
    outputs(7053) <= (layer0_outputs(10932)) and (layer0_outputs(8825));
    outputs(7054) <= (layer0_outputs(6907)) xor (layer0_outputs(5563));
    outputs(7055) <= layer0_outputs(11061);
    outputs(7056) <= layer0_outputs(3609);
    outputs(7057) <= (layer0_outputs(5161)) and (layer0_outputs(9103));
    outputs(7058) <= not((layer0_outputs(8603)) xor (layer0_outputs(7413)));
    outputs(7059) <= layer0_outputs(9973);
    outputs(7060) <= layer0_outputs(7305);
    outputs(7061) <= not(layer0_outputs(12281));
    outputs(7062) <= (layer0_outputs(5510)) xor (layer0_outputs(6209));
    outputs(7063) <= not((layer0_outputs(7715)) xor (layer0_outputs(426)));
    outputs(7064) <= layer0_outputs(1364);
    outputs(7065) <= layer0_outputs(4758);
    outputs(7066) <= layer0_outputs(6120);
    outputs(7067) <= layer0_outputs(4556);
    outputs(7068) <= (layer0_outputs(1812)) and (layer0_outputs(438));
    outputs(7069) <= not(layer0_outputs(5815)) or (layer0_outputs(4291));
    outputs(7070) <= '1';
    outputs(7071) <= not(layer0_outputs(213)) or (layer0_outputs(7214));
    outputs(7072) <= not((layer0_outputs(805)) xor (layer0_outputs(2750)));
    outputs(7073) <= layer0_outputs(2150);
    outputs(7074) <= (layer0_outputs(6)) xor (layer0_outputs(9707));
    outputs(7075) <= layer0_outputs(12664);
    outputs(7076) <= (layer0_outputs(1412)) or (layer0_outputs(3843));
    outputs(7077) <= not(layer0_outputs(257));
    outputs(7078) <= not(layer0_outputs(3985));
    outputs(7079) <= not((layer0_outputs(5768)) or (layer0_outputs(12445)));
    outputs(7080) <= layer0_outputs(1126);
    outputs(7081) <= not((layer0_outputs(11979)) xor (layer0_outputs(8580)));
    outputs(7082) <= not((layer0_outputs(3332)) xor (layer0_outputs(5710)));
    outputs(7083) <= (layer0_outputs(4604)) xor (layer0_outputs(7784));
    outputs(7084) <= (layer0_outputs(515)) xor (layer0_outputs(652));
    outputs(7085) <= not(layer0_outputs(4959)) or (layer0_outputs(3390));
    outputs(7086) <= layer0_outputs(1505);
    outputs(7087) <= not(layer0_outputs(3259)) or (layer0_outputs(11533));
    outputs(7088) <= not(layer0_outputs(6211));
    outputs(7089) <= not((layer0_outputs(6812)) or (layer0_outputs(8863)));
    outputs(7090) <= not((layer0_outputs(902)) xor (layer0_outputs(5386)));
    outputs(7091) <= not(layer0_outputs(6009)) or (layer0_outputs(10120));
    outputs(7092) <= not((layer0_outputs(12401)) xor (layer0_outputs(6447)));
    outputs(7093) <= (layer0_outputs(8165)) and (layer0_outputs(2544));
    outputs(7094) <= (layer0_outputs(951)) xor (layer0_outputs(930));
    outputs(7095) <= not((layer0_outputs(1167)) or (layer0_outputs(6789)));
    outputs(7096) <= layer0_outputs(10513);
    outputs(7097) <= (layer0_outputs(1552)) xor (layer0_outputs(5556));
    outputs(7098) <= not(layer0_outputs(4343));
    outputs(7099) <= not((layer0_outputs(1498)) and (layer0_outputs(3422)));
    outputs(7100) <= not((layer0_outputs(8417)) xor (layer0_outputs(5664)));
    outputs(7101) <= layer0_outputs(6390);
    outputs(7102) <= (layer0_outputs(8366)) or (layer0_outputs(5533));
    outputs(7103) <= (layer0_outputs(11015)) and not (layer0_outputs(9323));
    outputs(7104) <= not(layer0_outputs(6312));
    outputs(7105) <= not((layer0_outputs(12361)) xor (layer0_outputs(6862)));
    outputs(7106) <= layer0_outputs(681);
    outputs(7107) <= not((layer0_outputs(10388)) xor (layer0_outputs(9986)));
    outputs(7108) <= not((layer0_outputs(9749)) xor (layer0_outputs(11012)));
    outputs(7109) <= (layer0_outputs(9801)) and not (layer0_outputs(10147));
    outputs(7110) <= (layer0_outputs(7865)) and (layer0_outputs(7269));
    outputs(7111) <= not((layer0_outputs(12453)) xor (layer0_outputs(1625)));
    outputs(7112) <= not(layer0_outputs(2042)) or (layer0_outputs(7828));
    outputs(7113) <= (layer0_outputs(12353)) xor (layer0_outputs(8282));
    outputs(7114) <= not(layer0_outputs(6292));
    outputs(7115) <= not((layer0_outputs(11565)) xor (layer0_outputs(2593)));
    outputs(7116) <= not((layer0_outputs(8747)) or (layer0_outputs(7853)));
    outputs(7117) <= (layer0_outputs(5570)) xor (layer0_outputs(2425));
    outputs(7118) <= (layer0_outputs(6597)) or (layer0_outputs(10286));
    outputs(7119) <= layer0_outputs(1084);
    outputs(7120) <= (layer0_outputs(712)) or (layer0_outputs(7836));
    outputs(7121) <= layer0_outputs(10322);
    outputs(7122) <= not((layer0_outputs(6052)) xor (layer0_outputs(628)));
    outputs(7123) <= (layer0_outputs(5390)) and (layer0_outputs(6319));
    outputs(7124) <= not((layer0_outputs(5031)) xor (layer0_outputs(1124)));
    outputs(7125) <= not(layer0_outputs(4249));
    outputs(7126) <= (layer0_outputs(9379)) or (layer0_outputs(4029));
    outputs(7127) <= not(layer0_outputs(6960)) or (layer0_outputs(1301));
    outputs(7128) <= layer0_outputs(1821);
    outputs(7129) <= layer0_outputs(12782);
    outputs(7130) <= (layer0_outputs(2031)) xor (layer0_outputs(4451));
    outputs(7131) <= layer0_outputs(8170);
    outputs(7132) <= not((layer0_outputs(4484)) xor (layer0_outputs(4188)));
    outputs(7133) <= (layer0_outputs(341)) xor (layer0_outputs(6306));
    outputs(7134) <= not((layer0_outputs(10245)) xor (layer0_outputs(8223)));
    outputs(7135) <= (layer0_outputs(4727)) xor (layer0_outputs(7170));
    outputs(7136) <= (layer0_outputs(12646)) xor (layer0_outputs(2282));
    outputs(7137) <= (layer0_outputs(9786)) xor (layer0_outputs(5840));
    outputs(7138) <= (layer0_outputs(1623)) xor (layer0_outputs(5813));
    outputs(7139) <= not(layer0_outputs(9820));
    outputs(7140) <= not((layer0_outputs(7840)) xor (layer0_outputs(1921)));
    outputs(7141) <= layer0_outputs(4636);
    outputs(7142) <= not(layer0_outputs(5953));
    outputs(7143) <= not(layer0_outputs(10987)) or (layer0_outputs(11806));
    outputs(7144) <= not(layer0_outputs(11103));
    outputs(7145) <= layer0_outputs(1772);
    outputs(7146) <= (layer0_outputs(1587)) and not (layer0_outputs(7979));
    outputs(7147) <= not((layer0_outputs(2460)) xor (layer0_outputs(864)));
    outputs(7148) <= (layer0_outputs(6574)) xor (layer0_outputs(9766));
    outputs(7149) <= not(layer0_outputs(700));
    outputs(7150) <= not(layer0_outputs(12739)) or (layer0_outputs(4603));
    outputs(7151) <= not(layer0_outputs(2743));
    outputs(7152) <= (layer0_outputs(6905)) xor (layer0_outputs(9876));
    outputs(7153) <= not((layer0_outputs(7997)) xor (layer0_outputs(7135)));
    outputs(7154) <= not(layer0_outputs(11203));
    outputs(7155) <= not((layer0_outputs(5293)) and (layer0_outputs(525)));
    outputs(7156) <= not(layer0_outputs(8376));
    outputs(7157) <= not((layer0_outputs(3796)) xor (layer0_outputs(1736)));
    outputs(7158) <= not((layer0_outputs(8857)) or (layer0_outputs(12096)));
    outputs(7159) <= layer0_outputs(512);
    outputs(7160) <= not(layer0_outputs(3250));
    outputs(7161) <= not(layer0_outputs(2417));
    outputs(7162) <= layer0_outputs(1745);
    outputs(7163) <= not((layer0_outputs(3002)) xor (layer0_outputs(6508)));
    outputs(7164) <= (layer0_outputs(11663)) xor (layer0_outputs(2518));
    outputs(7165) <= (layer0_outputs(433)) xor (layer0_outputs(948));
    outputs(7166) <= layer0_outputs(2143);
    outputs(7167) <= not((layer0_outputs(4123)) xor (layer0_outputs(3224)));
    outputs(7168) <= (layer0_outputs(9568)) and not (layer0_outputs(3254));
    outputs(7169) <= not((layer0_outputs(5380)) xor (layer0_outputs(8900)));
    outputs(7170) <= not((layer0_outputs(7564)) and (layer0_outputs(4726)));
    outputs(7171) <= (layer0_outputs(5669)) xor (layer0_outputs(11201));
    outputs(7172) <= (layer0_outputs(297)) and (layer0_outputs(5920));
    outputs(7173) <= not(layer0_outputs(5739));
    outputs(7174) <= not((layer0_outputs(12513)) xor (layer0_outputs(2304)));
    outputs(7175) <= not(layer0_outputs(28));
    outputs(7176) <= layer0_outputs(12380);
    outputs(7177) <= not((layer0_outputs(6666)) xor (layer0_outputs(4269)));
    outputs(7178) <= (layer0_outputs(12385)) xor (layer0_outputs(10805));
    outputs(7179) <= layer0_outputs(569);
    outputs(7180) <= (layer0_outputs(7510)) and (layer0_outputs(946));
    outputs(7181) <= layer0_outputs(2503);
    outputs(7182) <= not(layer0_outputs(11433));
    outputs(7183) <= layer0_outputs(11814);
    outputs(7184) <= layer0_outputs(5610);
    outputs(7185) <= not(layer0_outputs(7150));
    outputs(7186) <= layer0_outputs(7507);
    outputs(7187) <= (layer0_outputs(8864)) or (layer0_outputs(2680));
    outputs(7188) <= not((layer0_outputs(3954)) xor (layer0_outputs(10655)));
    outputs(7189) <= layer0_outputs(1463);
    outputs(7190) <= (layer0_outputs(1259)) xor (layer0_outputs(7466));
    outputs(7191) <= (layer0_outputs(2922)) and not (layer0_outputs(4722));
    outputs(7192) <= not(layer0_outputs(7887));
    outputs(7193) <= (layer0_outputs(4948)) xor (layer0_outputs(1944));
    outputs(7194) <= not((layer0_outputs(8766)) xor (layer0_outputs(6177)));
    outputs(7195) <= not((layer0_outputs(1413)) xor (layer0_outputs(5827)));
    outputs(7196) <= not((layer0_outputs(3276)) xor (layer0_outputs(10746)));
    outputs(7197) <= not((layer0_outputs(6138)) xor (layer0_outputs(8559)));
    outputs(7198) <= layer0_outputs(12100);
    outputs(7199) <= not((layer0_outputs(12668)) xor (layer0_outputs(7637)));
    outputs(7200) <= (layer0_outputs(2369)) xor (layer0_outputs(9218));
    outputs(7201) <= layer0_outputs(262);
    outputs(7202) <= layer0_outputs(6368);
    outputs(7203) <= not((layer0_outputs(7421)) xor (layer0_outputs(2145)));
    outputs(7204) <= not(layer0_outputs(10218)) or (layer0_outputs(9988));
    outputs(7205) <= (layer0_outputs(9011)) xor (layer0_outputs(5873));
    outputs(7206) <= not(layer0_outputs(2829));
    outputs(7207) <= (layer0_outputs(9357)) xor (layer0_outputs(10));
    outputs(7208) <= not(layer0_outputs(9897)) or (layer0_outputs(239));
    outputs(7209) <= not(layer0_outputs(4279)) or (layer0_outputs(1741));
    outputs(7210) <= (layer0_outputs(2386)) and not (layer0_outputs(4866));
    outputs(7211) <= (layer0_outputs(7234)) xor (layer0_outputs(12666));
    outputs(7212) <= (layer0_outputs(6562)) and (layer0_outputs(1696));
    outputs(7213) <= (layer0_outputs(6066)) and (layer0_outputs(6625));
    outputs(7214) <= not(layer0_outputs(12118));
    outputs(7215) <= layer0_outputs(1887);
    outputs(7216) <= layer0_outputs(5911);
    outputs(7217) <= (layer0_outputs(10134)) xor (layer0_outputs(10205));
    outputs(7218) <= not(layer0_outputs(5544));
    outputs(7219) <= layer0_outputs(11331);
    outputs(7220) <= layer0_outputs(2040);
    outputs(7221) <= (layer0_outputs(1606)) xor (layer0_outputs(5584));
    outputs(7222) <= not((layer0_outputs(11871)) xor (layer0_outputs(6583)));
    outputs(7223) <= (layer0_outputs(4101)) or (layer0_outputs(7883));
    outputs(7224) <= (layer0_outputs(5157)) xor (layer0_outputs(5275));
    outputs(7225) <= (layer0_outputs(1320)) and not (layer0_outputs(3978));
    outputs(7226) <= not((layer0_outputs(7112)) xor (layer0_outputs(7377)));
    outputs(7227) <= not((layer0_outputs(2826)) xor (layer0_outputs(836)));
    outputs(7228) <= not((layer0_outputs(8669)) xor (layer0_outputs(2711)));
    outputs(7229) <= (layer0_outputs(2312)) xor (layer0_outputs(10645));
    outputs(7230) <= layer0_outputs(7741);
    outputs(7231) <= layer0_outputs(1917);
    outputs(7232) <= layer0_outputs(1517);
    outputs(7233) <= (layer0_outputs(12325)) xor (layer0_outputs(10270));
    outputs(7234) <= layer0_outputs(6322);
    outputs(7235) <= not((layer0_outputs(1276)) xor (layer0_outputs(1190)));
    outputs(7236) <= (layer0_outputs(8231)) or (layer0_outputs(359));
    outputs(7237) <= not((layer0_outputs(8311)) xor (layer0_outputs(4927)));
    outputs(7238) <= not(layer0_outputs(8585));
    outputs(7239) <= layer0_outputs(3632);
    outputs(7240) <= (layer0_outputs(1719)) or (layer0_outputs(6751));
    outputs(7241) <= (layer0_outputs(7015)) xor (layer0_outputs(6212));
    outputs(7242) <= not((layer0_outputs(953)) and (layer0_outputs(2760)));
    outputs(7243) <= (layer0_outputs(5004)) and not (layer0_outputs(5617));
    outputs(7244) <= not((layer0_outputs(12507)) or (layer0_outputs(5158)));
    outputs(7245) <= (layer0_outputs(2905)) xor (layer0_outputs(7257));
    outputs(7246) <= not(layer0_outputs(6027));
    outputs(7247) <= not(layer0_outputs(1992));
    outputs(7248) <= (layer0_outputs(813)) xor (layer0_outputs(6683));
    outputs(7249) <= not((layer0_outputs(5341)) xor (layer0_outputs(11359)));
    outputs(7250) <= (layer0_outputs(7629)) xor (layer0_outputs(11504));
    outputs(7251) <= (layer0_outputs(6450)) or (layer0_outputs(4314));
    outputs(7252) <= (layer0_outputs(10172)) or (layer0_outputs(199));
    outputs(7253) <= (layer0_outputs(922)) xor (layer0_outputs(2260));
    outputs(7254) <= (layer0_outputs(12316)) xor (layer0_outputs(10479));
    outputs(7255) <= layer0_outputs(3054);
    outputs(7256) <= not((layer0_outputs(10439)) xor (layer0_outputs(9902)));
    outputs(7257) <= (layer0_outputs(8338)) xor (layer0_outputs(3698));
    outputs(7258) <= not(layer0_outputs(4989));
    outputs(7259) <= not((layer0_outputs(12014)) xor (layer0_outputs(2992)));
    outputs(7260) <= not((layer0_outputs(9638)) or (layer0_outputs(12733)));
    outputs(7261) <= layer0_outputs(782);
    outputs(7262) <= not((layer0_outputs(8240)) xor (layer0_outputs(7491)));
    outputs(7263) <= layer0_outputs(9753);
    outputs(7264) <= not((layer0_outputs(1064)) xor (layer0_outputs(3715)));
    outputs(7265) <= not(layer0_outputs(12767));
    outputs(7266) <= not((layer0_outputs(4154)) xor (layer0_outputs(10979)));
    outputs(7267) <= not((layer0_outputs(9643)) xor (layer0_outputs(10135)));
    outputs(7268) <= layer0_outputs(5698);
    outputs(7269) <= not(layer0_outputs(989));
    outputs(7270) <= not(layer0_outputs(10596));
    outputs(7271) <= (layer0_outputs(11218)) xor (layer0_outputs(5698));
    outputs(7272) <= not((layer0_outputs(1419)) or (layer0_outputs(4921)));
    outputs(7273) <= not((layer0_outputs(5856)) xor (layer0_outputs(10274)));
    outputs(7274) <= not(layer0_outputs(10996));
    outputs(7275) <= not((layer0_outputs(4811)) xor (layer0_outputs(6658)));
    outputs(7276) <= (layer0_outputs(5411)) and not (layer0_outputs(12159));
    outputs(7277) <= not(layer0_outputs(7272));
    outputs(7278) <= layer0_outputs(12664);
    outputs(7279) <= (layer0_outputs(12427)) xor (layer0_outputs(9454));
    outputs(7280) <= layer0_outputs(9022);
    outputs(7281) <= (layer0_outputs(9935)) and (layer0_outputs(3060));
    outputs(7282) <= layer0_outputs(7589);
    outputs(7283) <= layer0_outputs(2008);
    outputs(7284) <= not((layer0_outputs(246)) xor (layer0_outputs(3046)));
    outputs(7285) <= layer0_outputs(9941);
    outputs(7286) <= (layer0_outputs(8044)) and (layer0_outputs(7160));
    outputs(7287) <= (layer0_outputs(10406)) xor (layer0_outputs(1147));
    outputs(7288) <= (layer0_outputs(5350)) xor (layer0_outputs(6038));
    outputs(7289) <= (layer0_outputs(4341)) xor (layer0_outputs(1482));
    outputs(7290) <= not((layer0_outputs(4083)) xor (layer0_outputs(6138)));
    outputs(7291) <= layer0_outputs(3493);
    outputs(7292) <= not(layer0_outputs(1296));
    outputs(7293) <= not((layer0_outputs(8811)) xor (layer0_outputs(5656)));
    outputs(7294) <= (layer0_outputs(3603)) and not (layer0_outputs(9931));
    outputs(7295) <= layer0_outputs(863);
    outputs(7296) <= (layer0_outputs(8714)) or (layer0_outputs(6388));
    outputs(7297) <= not((layer0_outputs(2245)) xor (layer0_outputs(8278)));
    outputs(7298) <= not(layer0_outputs(6173));
    outputs(7299) <= not(layer0_outputs(568)) or (layer0_outputs(6039));
    outputs(7300) <= (layer0_outputs(73)) xor (layer0_outputs(6514));
    outputs(7301) <= not((layer0_outputs(12648)) xor (layer0_outputs(8381)));
    outputs(7302) <= not((layer0_outputs(8106)) and (layer0_outputs(3430)));
    outputs(7303) <= (layer0_outputs(5367)) xor (layer0_outputs(2370));
    outputs(7304) <= layer0_outputs(1849);
    outputs(7305) <= (layer0_outputs(4155)) xor (layer0_outputs(8986));
    outputs(7306) <= not(layer0_outputs(6624));
    outputs(7307) <= (layer0_outputs(1281)) or (layer0_outputs(3897));
    outputs(7308) <= (layer0_outputs(930)) and not (layer0_outputs(10836));
    outputs(7309) <= (layer0_outputs(264)) xor (layer0_outputs(6183));
    outputs(7310) <= layer0_outputs(3345);
    outputs(7311) <= not(layer0_outputs(10649));
    outputs(7312) <= (layer0_outputs(3443)) and not (layer0_outputs(684));
    outputs(7313) <= (layer0_outputs(5125)) xor (layer0_outputs(9503));
    outputs(7314) <= not((layer0_outputs(6866)) xor (layer0_outputs(6623)));
    outputs(7315) <= not((layer0_outputs(4277)) xor (layer0_outputs(1257)));
    outputs(7316) <= not(layer0_outputs(4954));
    outputs(7317) <= (layer0_outputs(7101)) xor (layer0_outputs(7995));
    outputs(7318) <= not(layer0_outputs(2587)) or (layer0_outputs(10961));
    outputs(7319) <= (layer0_outputs(7695)) xor (layer0_outputs(5064));
    outputs(7320) <= not((layer0_outputs(3656)) xor (layer0_outputs(1461)));
    outputs(7321) <= (layer0_outputs(10749)) xor (layer0_outputs(5781));
    outputs(7322) <= not(layer0_outputs(11089));
    outputs(7323) <= layer0_outputs(6667);
    outputs(7324) <= (layer0_outputs(7266)) xor (layer0_outputs(5925));
    outputs(7325) <= not((layer0_outputs(9549)) xor (layer0_outputs(3141)));
    outputs(7326) <= (layer0_outputs(7205)) xor (layer0_outputs(6492));
    outputs(7327) <= not((layer0_outputs(3912)) xor (layer0_outputs(11330)));
    outputs(7328) <= not((layer0_outputs(7058)) xor (layer0_outputs(9177)));
    outputs(7329) <= not(layer0_outputs(6877));
    outputs(7330) <= (layer0_outputs(5904)) or (layer0_outputs(2878));
    outputs(7331) <= (layer0_outputs(6972)) and (layer0_outputs(6334));
    outputs(7332) <= not((layer0_outputs(8392)) xor (layer0_outputs(11705)));
    outputs(7333) <= layer0_outputs(3180);
    outputs(7334) <= layer0_outputs(10342);
    outputs(7335) <= layer0_outputs(11958);
    outputs(7336) <= layer0_outputs(1642);
    outputs(7337) <= layer0_outputs(9041);
    outputs(7338) <= (layer0_outputs(9010)) and (layer0_outputs(5452));
    outputs(7339) <= not(layer0_outputs(8840));
    outputs(7340) <= layer0_outputs(4398);
    outputs(7341) <= not(layer0_outputs(10214));
    outputs(7342) <= (layer0_outputs(5102)) xor (layer0_outputs(12706));
    outputs(7343) <= not((layer0_outputs(4438)) xor (layer0_outputs(11179)));
    outputs(7344) <= (layer0_outputs(7111)) or (layer0_outputs(8133));
    outputs(7345) <= (layer0_outputs(2736)) or (layer0_outputs(12180));
    outputs(7346) <= not(layer0_outputs(9704));
    outputs(7347) <= layer0_outputs(7686);
    outputs(7348) <= (layer0_outputs(12034)) xor (layer0_outputs(12506));
    outputs(7349) <= not((layer0_outputs(10966)) xor (layer0_outputs(4055)));
    outputs(7350) <= not(layer0_outputs(5755));
    outputs(7351) <= (layer0_outputs(7518)) xor (layer0_outputs(8365));
    outputs(7352) <= layer0_outputs(10757);
    outputs(7353) <= not(layer0_outputs(3188));
    outputs(7354) <= not((layer0_outputs(8629)) xor (layer0_outputs(7307)));
    outputs(7355) <= not((layer0_outputs(11643)) xor (layer0_outputs(0)));
    outputs(7356) <= not((layer0_outputs(12152)) xor (layer0_outputs(1539)));
    outputs(7357) <= not((layer0_outputs(2309)) xor (layer0_outputs(12170)));
    outputs(7358) <= not((layer0_outputs(1737)) xor (layer0_outputs(1572)));
    outputs(7359) <= not((layer0_outputs(5620)) xor (layer0_outputs(11175)));
    outputs(7360) <= not(layer0_outputs(694));
    outputs(7361) <= (layer0_outputs(3953)) xor (layer0_outputs(104));
    outputs(7362) <= not((layer0_outputs(8206)) or (layer0_outputs(6154)));
    outputs(7363) <= not((layer0_outputs(8196)) xor (layer0_outputs(11306)));
    outputs(7364) <= layer0_outputs(1938);
    outputs(7365) <= not((layer0_outputs(1475)) and (layer0_outputs(3013)));
    outputs(7366) <= (layer0_outputs(12562)) xor (layer0_outputs(8936));
    outputs(7367) <= not(layer0_outputs(8330)) or (layer0_outputs(1107));
    outputs(7368) <= (layer0_outputs(12490)) xor (layer0_outputs(1626));
    outputs(7369) <= not((layer0_outputs(8590)) xor (layer0_outputs(8989)));
    outputs(7370) <= layer0_outputs(7920);
    outputs(7371) <= layer0_outputs(7714);
    outputs(7372) <= not((layer0_outputs(6107)) xor (layer0_outputs(11494)));
    outputs(7373) <= (layer0_outputs(5738)) xor (layer0_outputs(8391));
    outputs(7374) <= not(layer0_outputs(9125));
    outputs(7375) <= (layer0_outputs(4309)) xor (layer0_outputs(10554));
    outputs(7376) <= (layer0_outputs(8724)) xor (layer0_outputs(7050));
    outputs(7377) <= not((layer0_outputs(5874)) xor (layer0_outputs(3619)));
    outputs(7378) <= (layer0_outputs(4358)) and not (layer0_outputs(6118));
    outputs(7379) <= (layer0_outputs(12649)) xor (layer0_outputs(8502));
    outputs(7380) <= not((layer0_outputs(3311)) or (layer0_outputs(6172)));
    outputs(7381) <= not((layer0_outputs(6868)) xor (layer0_outputs(813)));
    outputs(7382) <= (layer0_outputs(5607)) xor (layer0_outputs(10233));
    outputs(7383) <= (layer0_outputs(6479)) xor (layer0_outputs(1939));
    outputs(7384) <= layer0_outputs(594);
    outputs(7385) <= not(layer0_outputs(2080));
    outputs(7386) <= (layer0_outputs(7806)) and not (layer0_outputs(11902));
    outputs(7387) <= not(layer0_outputs(3063));
    outputs(7388) <= not(layer0_outputs(1959));
    outputs(7389) <= not(layer0_outputs(12552)) or (layer0_outputs(5591));
    outputs(7390) <= (layer0_outputs(4118)) xor (layer0_outputs(3777));
    outputs(7391) <= not((layer0_outputs(12655)) xor (layer0_outputs(4253)));
    outputs(7392) <= (layer0_outputs(11486)) and not (layer0_outputs(4848));
    outputs(7393) <= not((layer0_outputs(4818)) or (layer0_outputs(10139)));
    outputs(7394) <= not((layer0_outputs(5541)) xor (layer0_outputs(9917)));
    outputs(7395) <= (layer0_outputs(10782)) xor (layer0_outputs(654));
    outputs(7396) <= not((layer0_outputs(2868)) xor (layer0_outputs(5803)));
    outputs(7397) <= (layer0_outputs(5092)) or (layer0_outputs(8773));
    outputs(7398) <= not((layer0_outputs(743)) xor (layer0_outputs(3598)));
    outputs(7399) <= (layer0_outputs(2224)) and not (layer0_outputs(12001));
    outputs(7400) <= (layer0_outputs(4381)) and (layer0_outputs(9542));
    outputs(7401) <= layer0_outputs(7516);
    outputs(7402) <= not((layer0_outputs(4221)) xor (layer0_outputs(12216)));
    outputs(7403) <= (layer0_outputs(9524)) xor (layer0_outputs(12575));
    outputs(7404) <= layer0_outputs(12535);
    outputs(7405) <= layer0_outputs(3775);
    outputs(7406) <= not((layer0_outputs(7281)) xor (layer0_outputs(10138)));
    outputs(7407) <= (layer0_outputs(141)) xor (layer0_outputs(12473));
    outputs(7408) <= layer0_outputs(8147);
    outputs(7409) <= not(layer0_outputs(1550));
    outputs(7410) <= not((layer0_outputs(12524)) and (layer0_outputs(6194)));
    outputs(7411) <= (layer0_outputs(5745)) xor (layer0_outputs(4527));
    outputs(7412) <= (layer0_outputs(10874)) xor (layer0_outputs(6874));
    outputs(7413) <= (layer0_outputs(6742)) xor (layer0_outputs(7054));
    outputs(7414) <= not(layer0_outputs(7087)) or (layer0_outputs(11692));
    outputs(7415) <= not((layer0_outputs(2)) and (layer0_outputs(3069)));
    outputs(7416) <= (layer0_outputs(9437)) and not (layer0_outputs(7037));
    outputs(7417) <= '0';
    outputs(7418) <= (layer0_outputs(6852)) xor (layer0_outputs(5773));
    outputs(7419) <= not((layer0_outputs(9350)) xor (layer0_outputs(6664)));
    outputs(7420) <= not(layer0_outputs(2060));
    outputs(7421) <= not(layer0_outputs(8867));
    outputs(7422) <= (layer0_outputs(4565)) and not (layer0_outputs(4497));
    outputs(7423) <= not(layer0_outputs(1363));
    outputs(7424) <= (layer0_outputs(4877)) and (layer0_outputs(8346));
    outputs(7425) <= (layer0_outputs(10744)) and not (layer0_outputs(5969));
    outputs(7426) <= (layer0_outputs(11465)) xor (layer0_outputs(8634));
    outputs(7427) <= not((layer0_outputs(8719)) xor (layer0_outputs(4522)));
    outputs(7428) <= layer0_outputs(7990);
    outputs(7429) <= not(layer0_outputs(10158));
    outputs(7430) <= (layer0_outputs(12143)) xor (layer0_outputs(8109));
    outputs(7431) <= not((layer0_outputs(853)) xor (layer0_outputs(932)));
    outputs(7432) <= layer0_outputs(794);
    outputs(7433) <= not((layer0_outputs(7416)) and (layer0_outputs(6613)));
    outputs(7434) <= layer0_outputs(9937);
    outputs(7435) <= (layer0_outputs(3031)) xor (layer0_outputs(11078));
    outputs(7436) <= not(layer0_outputs(8768));
    outputs(7437) <= not(layer0_outputs(5729)) or (layer0_outputs(10826));
    outputs(7438) <= (layer0_outputs(7370)) xor (layer0_outputs(11184));
    outputs(7439) <= layer0_outputs(2215);
    outputs(7440) <= (layer0_outputs(993)) and not (layer0_outputs(1825));
    outputs(7441) <= (layer0_outputs(2644)) xor (layer0_outputs(1557));
    outputs(7442) <= (layer0_outputs(355)) xor (layer0_outputs(6310));
    outputs(7443) <= layer0_outputs(9959);
    outputs(7444) <= not(layer0_outputs(2320));
    outputs(7445) <= layer0_outputs(5434);
    outputs(7446) <= not((layer0_outputs(5161)) xor (layer0_outputs(11495)));
    outputs(7447) <= layer0_outputs(1445);
    outputs(7448) <= layer0_outputs(10037);
    outputs(7449) <= (layer0_outputs(10988)) xor (layer0_outputs(8242));
    outputs(7450) <= not((layer0_outputs(2762)) xor (layer0_outputs(4540)));
    outputs(7451) <= (layer0_outputs(5906)) xor (layer0_outputs(4296));
    outputs(7452) <= not((layer0_outputs(8565)) xor (layer0_outputs(8274)));
    outputs(7453) <= (layer0_outputs(6441)) xor (layer0_outputs(6541));
    outputs(7454) <= (layer0_outputs(8074)) xor (layer0_outputs(663));
    outputs(7455) <= layer0_outputs(7691);
    outputs(7456) <= layer0_outputs(8017);
    outputs(7457) <= not((layer0_outputs(2981)) xor (layer0_outputs(3599)));
    outputs(7458) <= (layer0_outputs(6516)) and (layer0_outputs(8225));
    outputs(7459) <= not((layer0_outputs(12572)) xor (layer0_outputs(2807)));
    outputs(7460) <= not(layer0_outputs(6292));
    outputs(7461) <= layer0_outputs(11255);
    outputs(7462) <= layer0_outputs(6632);
    outputs(7463) <= not((layer0_outputs(11169)) xor (layer0_outputs(5137)));
    outputs(7464) <= not(layer0_outputs(12762));
    outputs(7465) <= (layer0_outputs(10177)) and not (layer0_outputs(1948));
    outputs(7466) <= not(layer0_outputs(10519));
    outputs(7467) <= (layer0_outputs(5447)) or (layer0_outputs(5829));
    outputs(7468) <= not((layer0_outputs(9663)) xor (layer0_outputs(8915)));
    outputs(7469) <= not((layer0_outputs(2647)) xor (layer0_outputs(3848)));
    outputs(7470) <= (layer0_outputs(701)) xor (layer0_outputs(591));
    outputs(7471) <= (layer0_outputs(6331)) xor (layer0_outputs(6649));
    outputs(7472) <= not((layer0_outputs(907)) xor (layer0_outputs(6685)));
    outputs(7473) <= not(layer0_outputs(9073));
    outputs(7474) <= not(layer0_outputs(8296));
    outputs(7475) <= not(layer0_outputs(12371));
    outputs(7476) <= not((layer0_outputs(4629)) and (layer0_outputs(7633)));
    outputs(7477) <= (layer0_outputs(10928)) xor (layer0_outputs(10368));
    outputs(7478) <= not((layer0_outputs(6325)) xor (layer0_outputs(7086)));
    outputs(7479) <= layer0_outputs(3404);
    outputs(7480) <= layer0_outputs(12367);
    outputs(7481) <= (layer0_outputs(6950)) xor (layer0_outputs(1504));
    outputs(7482) <= not((layer0_outputs(12636)) and (layer0_outputs(3242)));
    outputs(7483) <= not((layer0_outputs(2770)) xor (layer0_outputs(190)));
    outputs(7484) <= layer0_outputs(4899);
    outputs(7485) <= not(layer0_outputs(3622));
    outputs(7486) <= (layer0_outputs(2174)) xor (layer0_outputs(6585));
    outputs(7487) <= not((layer0_outputs(9315)) xor (layer0_outputs(936)));
    outputs(7488) <= not((layer0_outputs(11772)) and (layer0_outputs(839)));
    outputs(7489) <= (layer0_outputs(11368)) xor (layer0_outputs(1418));
    outputs(7490) <= layer0_outputs(12509);
    outputs(7491) <= not(layer0_outputs(12156));
    outputs(7492) <= not(layer0_outputs(3300)) or (layer0_outputs(8957));
    outputs(7493) <= not(layer0_outputs(11037)) or (layer0_outputs(5766));
    outputs(7494) <= layer0_outputs(3245);
    outputs(7495) <= not((layer0_outputs(10911)) and (layer0_outputs(6480)));
    outputs(7496) <= not(layer0_outputs(6465)) or (layer0_outputs(1815));
    outputs(7497) <= (layer0_outputs(10948)) xor (layer0_outputs(7344));
    outputs(7498) <= (layer0_outputs(5388)) xor (layer0_outputs(11106));
    outputs(7499) <= not((layer0_outputs(12230)) xor (layer0_outputs(6554)));
    outputs(7500) <= (layer0_outputs(6943)) or (layer0_outputs(8790));
    outputs(7501) <= (layer0_outputs(5096)) and not (layer0_outputs(67));
    outputs(7502) <= (layer0_outputs(4985)) and not (layer0_outputs(1133));
    outputs(7503) <= (layer0_outputs(10630)) xor (layer0_outputs(7628));
    outputs(7504) <= not((layer0_outputs(2527)) xor (layer0_outputs(12515)));
    outputs(7505) <= not((layer0_outputs(2947)) and (layer0_outputs(8890)));
    outputs(7506) <= (layer0_outputs(1074)) or (layer0_outputs(4502));
    outputs(7507) <= layer0_outputs(3546);
    outputs(7508) <= not(layer0_outputs(12578)) or (layer0_outputs(10682));
    outputs(7509) <= not((layer0_outputs(3417)) xor (layer0_outputs(4672)));
    outputs(7510) <= not(layer0_outputs(3127));
    outputs(7511) <= not((layer0_outputs(3996)) xor (layer0_outputs(2825)));
    outputs(7512) <= (layer0_outputs(4775)) xor (layer0_outputs(1926));
    outputs(7513) <= not(layer0_outputs(1383));
    outputs(7514) <= '1';
    outputs(7515) <= not(layer0_outputs(5935));
    outputs(7516) <= not((layer0_outputs(1760)) xor (layer0_outputs(7149)));
    outputs(7517) <= (layer0_outputs(4782)) xor (layer0_outputs(4706));
    outputs(7518) <= (layer0_outputs(6208)) xor (layer0_outputs(3900));
    outputs(7519) <= not(layer0_outputs(4538));
    outputs(7520) <= layer0_outputs(10052);
    outputs(7521) <= not((layer0_outputs(6940)) xor (layer0_outputs(5315)));
    outputs(7522) <= not((layer0_outputs(1144)) xor (layer0_outputs(5914)));
    outputs(7523) <= (layer0_outputs(830)) xor (layer0_outputs(2991));
    outputs(7524) <= not((layer0_outputs(3254)) or (layer0_outputs(8626)));
    outputs(7525) <= not(layer0_outputs(11259));
    outputs(7526) <= not(layer0_outputs(12619));
    outputs(7527) <= not((layer0_outputs(9720)) xor (layer0_outputs(7989)));
    outputs(7528) <= layer0_outputs(11553);
    outputs(7529) <= layer0_outputs(9288);
    outputs(7530) <= not(layer0_outputs(12466));
    outputs(7531) <= not(layer0_outputs(797));
    outputs(7532) <= (layer0_outputs(11603)) and (layer0_outputs(2617));
    outputs(7533) <= not((layer0_outputs(10918)) xor (layer0_outputs(8824)));
    outputs(7534) <= layer0_outputs(3677);
    outputs(7535) <= not(layer0_outputs(2651)) or (layer0_outputs(6236));
    outputs(7536) <= layer0_outputs(8016);
    outputs(7537) <= not(layer0_outputs(9956));
    outputs(7538) <= not((layer0_outputs(8392)) xor (layer0_outputs(11583)));
    outputs(7539) <= (layer0_outputs(6872)) xor (layer0_outputs(8011));
    outputs(7540) <= layer0_outputs(4536);
    outputs(7541) <= not(layer0_outputs(12716));
    outputs(7542) <= not((layer0_outputs(1809)) xor (layer0_outputs(12307)));
    outputs(7543) <= (layer0_outputs(10446)) and not (layer0_outputs(1958));
    outputs(7544) <= (layer0_outputs(7027)) xor (layer0_outputs(11024));
    outputs(7545) <= not(layer0_outputs(9473)) or (layer0_outputs(7165));
    outputs(7546) <= not(layer0_outputs(11484));
    outputs(7547) <= not(layer0_outputs(3842)) or (layer0_outputs(8781));
    outputs(7548) <= not(layer0_outputs(6545));
    outputs(7549) <= (layer0_outputs(8384)) xor (layer0_outputs(7875));
    outputs(7550) <= layer0_outputs(9545);
    outputs(7551) <= not(layer0_outputs(7241));
    outputs(7552) <= not((layer0_outputs(10227)) xor (layer0_outputs(6615)));
    outputs(7553) <= layer0_outputs(3964);
    outputs(7554) <= layer0_outputs(5519);
    outputs(7555) <= layer0_outputs(11549);
    outputs(7556) <= (layer0_outputs(12621)) xor (layer0_outputs(2187));
    outputs(7557) <= not(layer0_outputs(2071));
    outputs(7558) <= not((layer0_outputs(3373)) xor (layer0_outputs(11913)));
    outputs(7559) <= (layer0_outputs(2584)) xor (layer0_outputs(6611));
    outputs(7560) <= not((layer0_outputs(12654)) and (layer0_outputs(4071)));
    outputs(7561) <= layer0_outputs(4330);
    outputs(7562) <= not((layer0_outputs(1159)) xor (layer0_outputs(1790)));
    outputs(7563) <= layer0_outputs(8563);
    outputs(7564) <= not((layer0_outputs(685)) or (layer0_outputs(1857)));
    outputs(7565) <= not((layer0_outputs(6158)) xor (layer0_outputs(4907)));
    outputs(7566) <= not(layer0_outputs(7110));
    outputs(7567) <= (layer0_outputs(610)) xor (layer0_outputs(9161));
    outputs(7568) <= layer0_outputs(6608);
    outputs(7569) <= layer0_outputs(11860);
    outputs(7570) <= not(layer0_outputs(5357));
    outputs(7571) <= (layer0_outputs(11903)) or (layer0_outputs(7125));
    outputs(7572) <= not((layer0_outputs(9003)) xor (layer0_outputs(2809)));
    outputs(7573) <= layer0_outputs(2586);
    outputs(7574) <= not((layer0_outputs(4744)) and (layer0_outputs(2776)));
    outputs(7575) <= not((layer0_outputs(4678)) xor (layer0_outputs(11968)));
    outputs(7576) <= (layer0_outputs(9695)) or (layer0_outputs(5179));
    outputs(7577) <= not((layer0_outputs(7670)) xor (layer0_outputs(2033)));
    outputs(7578) <= not(layer0_outputs(11283));
    outputs(7579) <= not((layer0_outputs(167)) xor (layer0_outputs(9766)));
    outputs(7580) <= not(layer0_outputs(5731));
    outputs(7581) <= (layer0_outputs(9477)) or (layer0_outputs(10674));
    outputs(7582) <= not((layer0_outputs(2180)) xor (layer0_outputs(3258)));
    outputs(7583) <= not((layer0_outputs(1228)) xor (layer0_outputs(2479)));
    outputs(7584) <= not(layer0_outputs(6132));
    outputs(7585) <= not((layer0_outputs(2704)) xor (layer0_outputs(12705)));
    outputs(7586) <= layer0_outputs(6390);
    outputs(7587) <= not(layer0_outputs(2532)) or (layer0_outputs(10822));
    outputs(7588) <= not((layer0_outputs(577)) xor (layer0_outputs(789)));
    outputs(7589) <= (layer0_outputs(10625)) and not (layer0_outputs(11372));
    outputs(7590) <= layer0_outputs(1970);
    outputs(7591) <= not((layer0_outputs(3810)) xor (layer0_outputs(2183)));
    outputs(7592) <= (layer0_outputs(2748)) xor (layer0_outputs(10885));
    outputs(7593) <= layer0_outputs(6136);
    outputs(7594) <= layer0_outputs(7);
    outputs(7595) <= not((layer0_outputs(11924)) and (layer0_outputs(10023)));
    outputs(7596) <= layer0_outputs(1269);
    outputs(7597) <= (layer0_outputs(9281)) or (layer0_outputs(11290));
    outputs(7598) <= not(layer0_outputs(3529)) or (layer0_outputs(8188));
    outputs(7599) <= not((layer0_outputs(7976)) xor (layer0_outputs(3639)));
    outputs(7600) <= not((layer0_outputs(8339)) xor (layer0_outputs(9439)));
    outputs(7601) <= (layer0_outputs(7938)) and not (layer0_outputs(12783));
    outputs(7602) <= not(layer0_outputs(2860));
    outputs(7603) <= layer0_outputs(2102);
    outputs(7604) <= not(layer0_outputs(7870));
    outputs(7605) <= (layer0_outputs(6072)) and not (layer0_outputs(5242));
    outputs(7606) <= not((layer0_outputs(6143)) xor (layer0_outputs(7277)));
    outputs(7607) <= (layer0_outputs(4662)) xor (layer0_outputs(1172));
    outputs(7608) <= not((layer0_outputs(9375)) xor (layer0_outputs(9484)));
    outputs(7609) <= not(layer0_outputs(7026));
    outputs(7610) <= not((layer0_outputs(3026)) and (layer0_outputs(619)));
    outputs(7611) <= layer0_outputs(12243);
    outputs(7612) <= not(layer0_outputs(8373));
    outputs(7613) <= (layer0_outputs(12388)) or (layer0_outputs(418));
    outputs(7614) <= (layer0_outputs(9964)) and not (layer0_outputs(2530));
    outputs(7615) <= not((layer0_outputs(5826)) or (layer0_outputs(9143)));
    outputs(7616) <= not((layer0_outputs(6707)) and (layer0_outputs(5846)));
    outputs(7617) <= (layer0_outputs(6591)) or (layer0_outputs(11485));
    outputs(7618) <= (layer0_outputs(11508)) and (layer0_outputs(12563));
    outputs(7619) <= layer0_outputs(675);
    outputs(7620) <= not((layer0_outputs(1768)) or (layer0_outputs(8890)));
    outputs(7621) <= layer0_outputs(264);
    outputs(7622) <= not((layer0_outputs(281)) and (layer0_outputs(4374)));
    outputs(7623) <= not(layer0_outputs(11043)) or (layer0_outputs(5696));
    outputs(7624) <= layer0_outputs(10717);
    outputs(7625) <= not((layer0_outputs(12014)) xor (layer0_outputs(4166)));
    outputs(7626) <= not((layer0_outputs(12163)) and (layer0_outputs(5328)));
    outputs(7627) <= layer0_outputs(2199);
    outputs(7628) <= not((layer0_outputs(2250)) xor (layer0_outputs(2984)));
    outputs(7629) <= not((layer0_outputs(1635)) xor (layer0_outputs(12282)));
    outputs(7630) <= not((layer0_outputs(9215)) xor (layer0_outputs(6101)));
    outputs(7631) <= layer0_outputs(4840);
    outputs(7632) <= not(layer0_outputs(10508));
    outputs(7633) <= (layer0_outputs(8232)) and (layer0_outputs(2513));
    outputs(7634) <= layer0_outputs(9130);
    outputs(7635) <= (layer0_outputs(3035)) xor (layer0_outputs(10280));
    outputs(7636) <= layer0_outputs(3746);
    outputs(7637) <= (layer0_outputs(3853)) xor (layer0_outputs(1191));
    outputs(7638) <= (layer0_outputs(3600)) xor (layer0_outputs(5785));
    outputs(7639) <= not(layer0_outputs(12445));
    outputs(7640) <= (layer0_outputs(5866)) and (layer0_outputs(6048));
    outputs(7641) <= (layer0_outputs(6844)) and not (layer0_outputs(1437));
    outputs(7642) <= (layer0_outputs(4125)) xor (layer0_outputs(1654));
    outputs(7643) <= not(layer0_outputs(9901));
    outputs(7644) <= not((layer0_outputs(460)) xor (layer0_outputs(12770)));
    outputs(7645) <= (layer0_outputs(11451)) xor (layer0_outputs(10005));
    outputs(7646) <= layer0_outputs(12219);
    outputs(7647) <= not(layer0_outputs(5986));
    outputs(7648) <= (layer0_outputs(3480)) and (layer0_outputs(10465));
    outputs(7649) <= (layer0_outputs(3415)) and not (layer0_outputs(4035));
    outputs(7650) <= layer0_outputs(8587);
    outputs(7651) <= not((layer0_outputs(6112)) xor (layer0_outputs(10275)));
    outputs(7652) <= not((layer0_outputs(10976)) or (layer0_outputs(12641)));
    outputs(7653) <= not(layer0_outputs(9407));
    outputs(7654) <= layer0_outputs(9627);
    outputs(7655) <= not((layer0_outputs(8362)) xor (layer0_outputs(4104)));
    outputs(7656) <= (layer0_outputs(10855)) or (layer0_outputs(1419));
    outputs(7657) <= not((layer0_outputs(3482)) xor (layer0_outputs(540)));
    outputs(7658) <= not(layer0_outputs(7655));
    outputs(7659) <= not(layer0_outputs(2558));
    outputs(7660) <= (layer0_outputs(7797)) or (layer0_outputs(3535));
    outputs(7661) <= (layer0_outputs(3344)) xor (layer0_outputs(11442));
    outputs(7662) <= (layer0_outputs(10268)) xor (layer0_outputs(5703));
    outputs(7663) <= not((layer0_outputs(10876)) xor (layer0_outputs(4078)));
    outputs(7664) <= not((layer0_outputs(4069)) xor (layer0_outputs(8446)));
    outputs(7665) <= layer0_outputs(7263);
    outputs(7666) <= not((layer0_outputs(6028)) xor (layer0_outputs(9207)));
    outputs(7667) <= layer0_outputs(1256);
    outputs(7668) <= (layer0_outputs(11453)) xor (layer0_outputs(1824));
    outputs(7669) <= (layer0_outputs(10750)) xor (layer0_outputs(9283));
    outputs(7670) <= (layer0_outputs(5078)) xor (layer0_outputs(4324));
    outputs(7671) <= (layer0_outputs(7121)) xor (layer0_outputs(4170));
    outputs(7672) <= (layer0_outputs(11063)) and (layer0_outputs(1176));
    outputs(7673) <= layer0_outputs(9480);
    outputs(7674) <= layer0_outputs(7785);
    outputs(7675) <= not((layer0_outputs(8214)) xor (layer0_outputs(1934)));
    outputs(7676) <= layer0_outputs(4283);
    outputs(7677) <= layer0_outputs(11916);
    outputs(7678) <= layer0_outputs(3998);
    outputs(7679) <= not((layer0_outputs(10045)) xor (layer0_outputs(6711)));
    outputs(7680) <= layer0_outputs(10603);
    outputs(7681) <= layer0_outputs(9675);
    outputs(7682) <= not((layer0_outputs(10543)) xor (layer0_outputs(3858)));
    outputs(7683) <= (layer0_outputs(3609)) and (layer0_outputs(12357));
    outputs(7684) <= (layer0_outputs(11514)) and not (layer0_outputs(11522));
    outputs(7685) <= not((layer0_outputs(397)) or (layer0_outputs(5633)));
    outputs(7686) <= not((layer0_outputs(7354)) xor (layer0_outputs(6074)));
    outputs(7687) <= not((layer0_outputs(11808)) or (layer0_outputs(8626)));
    outputs(7688) <= layer0_outputs(11974);
    outputs(7689) <= (layer0_outputs(8595)) and not (layer0_outputs(11939));
    outputs(7690) <= not(layer0_outputs(1760));
    outputs(7691) <= not((layer0_outputs(12546)) xor (layer0_outputs(6428)));
    outputs(7692) <= layer0_outputs(2852);
    outputs(7693) <= not(layer0_outputs(8285));
    outputs(7694) <= not((layer0_outputs(3505)) and (layer0_outputs(12360)));
    outputs(7695) <= not(layer0_outputs(3321));
    outputs(7696) <= (layer0_outputs(2890)) xor (layer0_outputs(4251));
    outputs(7697) <= not(layer0_outputs(4349));
    outputs(7698) <= not((layer0_outputs(528)) or (layer0_outputs(12200)));
    outputs(7699) <= not(layer0_outputs(6993));
    outputs(7700) <= layer0_outputs(6438);
    outputs(7701) <= layer0_outputs(4760);
    outputs(7702) <= (layer0_outputs(3269)) and (layer0_outputs(10558));
    outputs(7703) <= not(layer0_outputs(4721));
    outputs(7704) <= not(layer0_outputs(11905));
    outputs(7705) <= (layer0_outputs(2393)) and not (layer0_outputs(5037));
    outputs(7706) <= (layer0_outputs(8956)) and not (layer0_outputs(8083));
    outputs(7707) <= not(layer0_outputs(11007)) or (layer0_outputs(1535));
    outputs(7708) <= (layer0_outputs(9748)) and not (layer0_outputs(8494));
    outputs(7709) <= (layer0_outputs(2994)) xor (layer0_outputs(8345));
    outputs(7710) <= (layer0_outputs(3697)) and not (layer0_outputs(6313));
    outputs(7711) <= not(layer0_outputs(7567)) or (layer0_outputs(4693));
    outputs(7712) <= not((layer0_outputs(2040)) xor (layer0_outputs(12334)));
    outputs(7713) <= layer0_outputs(1685);
    outputs(7714) <= not(layer0_outputs(3572));
    outputs(7715) <= layer0_outputs(10493);
    outputs(7716) <= (layer0_outputs(1118)) or (layer0_outputs(80));
    outputs(7717) <= not((layer0_outputs(1154)) xor (layer0_outputs(9386)));
    outputs(7718) <= not(layer0_outputs(11587));
    outputs(7719) <= layer0_outputs(3616);
    outputs(7720) <= layer0_outputs(6739);
    outputs(7721) <= not((layer0_outputs(8815)) xor (layer0_outputs(6598)));
    outputs(7722) <= not(layer0_outputs(9138));
    outputs(7723) <= not(layer0_outputs(6284)) or (layer0_outputs(12283));
    outputs(7724) <= not((layer0_outputs(6775)) or (layer0_outputs(1888)));
    outputs(7725) <= not(layer0_outputs(6865));
    outputs(7726) <= layer0_outputs(521);
    outputs(7727) <= (layer0_outputs(8559)) or (layer0_outputs(2339));
    outputs(7728) <= layer0_outputs(4781);
    outputs(7729) <= (layer0_outputs(12625)) xor (layer0_outputs(10240));
    outputs(7730) <= not(layer0_outputs(12652));
    outputs(7731) <= (layer0_outputs(580)) and not (layer0_outputs(10899));
    outputs(7732) <= not((layer0_outputs(12755)) and (layer0_outputs(4934)));
    outputs(7733) <= not(layer0_outputs(6603));
    outputs(7734) <= layer0_outputs(4164);
    outputs(7735) <= (layer0_outputs(6130)) xor (layer0_outputs(3765));
    outputs(7736) <= (layer0_outputs(351)) xor (layer0_outputs(11412));
    outputs(7737) <= layer0_outputs(6472);
    outputs(7738) <= not(layer0_outputs(7716));
    outputs(7739) <= (layer0_outputs(2992)) and not (layer0_outputs(5556));
    outputs(7740) <= (layer0_outputs(8267)) and not (layer0_outputs(12317));
    outputs(7741) <= not((layer0_outputs(1778)) xor (layer0_outputs(24)));
    outputs(7742) <= not((layer0_outputs(1659)) xor (layer0_outputs(10558)));
    outputs(7743) <= not(layer0_outputs(10984)) or (layer0_outputs(10777));
    outputs(7744) <= layer0_outputs(8765);
    outputs(7745) <= layer0_outputs(11665);
    outputs(7746) <= not(layer0_outputs(11258));
    outputs(7747) <= (layer0_outputs(4243)) and (layer0_outputs(376));
    outputs(7748) <= layer0_outputs(2010);
    outputs(7749) <= layer0_outputs(4796);
    outputs(7750) <= not(layer0_outputs(6818)) or (layer0_outputs(2588));
    outputs(7751) <= layer0_outputs(2765);
    outputs(7752) <= (layer0_outputs(3919)) and not (layer0_outputs(207));
    outputs(7753) <= not(layer0_outputs(688));
    outputs(7754) <= not((layer0_outputs(6494)) xor (layer0_outputs(7094)));
    outputs(7755) <= (layer0_outputs(8685)) and not (layer0_outputs(5010));
    outputs(7756) <= not(layer0_outputs(54));
    outputs(7757) <= not(layer0_outputs(979));
    outputs(7758) <= layer0_outputs(5472);
    outputs(7759) <= not(layer0_outputs(7249));
    outputs(7760) <= not((layer0_outputs(871)) or (layer0_outputs(6801)));
    outputs(7761) <= layer0_outputs(3565);
    outputs(7762) <= not(layer0_outputs(10808));
    outputs(7763) <= (layer0_outputs(1955)) or (layer0_outputs(10800));
    outputs(7764) <= not(layer0_outputs(2296));
    outputs(7765) <= (layer0_outputs(1639)) and not (layer0_outputs(6651));
    outputs(7766) <= not((layer0_outputs(6335)) xor (layer0_outputs(2817)));
    outputs(7767) <= (layer0_outputs(11539)) and not (layer0_outputs(10296));
    outputs(7768) <= layer0_outputs(5790);
    outputs(7769) <= not(layer0_outputs(11488));
    outputs(7770) <= (layer0_outputs(10138)) xor (layer0_outputs(7009));
    outputs(7771) <= (layer0_outputs(3145)) and not (layer0_outputs(11443));
    outputs(7772) <= layer0_outputs(9356);
    outputs(7773) <= not(layer0_outputs(7128));
    outputs(7774) <= not(layer0_outputs(11221));
    outputs(7775) <= not((layer0_outputs(2389)) and (layer0_outputs(9946)));
    outputs(7776) <= layer0_outputs(6961);
    outputs(7777) <= (layer0_outputs(5780)) xor (layer0_outputs(12320));
    outputs(7778) <= not(layer0_outputs(131));
    outputs(7779) <= not(layer0_outputs(2175));
    outputs(7780) <= not((layer0_outputs(10455)) and (layer0_outputs(9167)));
    outputs(7781) <= not((layer0_outputs(7276)) xor (layer0_outputs(8657)));
    outputs(7782) <= (layer0_outputs(10549)) and (layer0_outputs(5385));
    outputs(7783) <= layer0_outputs(7863);
    outputs(7784) <= layer0_outputs(12440);
    outputs(7785) <= not((layer0_outputs(5674)) and (layer0_outputs(12334)));
    outputs(7786) <= layer0_outputs(1904);
    outputs(7787) <= layer0_outputs(4138);
    outputs(7788) <= not((layer0_outputs(7102)) xor (layer0_outputs(11356)));
    outputs(7789) <= not(layer0_outputs(9462));
    outputs(7790) <= layer0_outputs(3153);
    outputs(7791) <= layer0_outputs(8751);
    outputs(7792) <= (layer0_outputs(2981)) and not (layer0_outputs(8351));
    outputs(7793) <= (layer0_outputs(788)) and not (layer0_outputs(8071));
    outputs(7794) <= not(layer0_outputs(7825));
    outputs(7795) <= layer0_outputs(3077);
    outputs(7796) <= not(layer0_outputs(8278));
    outputs(7797) <= layer0_outputs(8436);
    outputs(7798) <= layer0_outputs(5038);
    outputs(7799) <= not(layer0_outputs(9761));
    outputs(7800) <= layer0_outputs(6230);
    outputs(7801) <= layer0_outputs(6864);
    outputs(7802) <= (layer0_outputs(9507)) or (layer0_outputs(11749));
    outputs(7803) <= (layer0_outputs(6182)) xor (layer0_outputs(9388));
    outputs(7804) <= layer0_outputs(763);
    outputs(7805) <= (layer0_outputs(2207)) xor (layer0_outputs(6174));
    outputs(7806) <= (layer0_outputs(7449)) xor (layer0_outputs(12250));
    outputs(7807) <= (layer0_outputs(9881)) and not (layer0_outputs(5685));
    outputs(7808) <= layer0_outputs(8991);
    outputs(7809) <= layer0_outputs(7231);
    outputs(7810) <= not(layer0_outputs(8295));
    outputs(7811) <= not(layer0_outputs(95));
    outputs(7812) <= (layer0_outputs(1375)) xor (layer0_outputs(8713));
    outputs(7813) <= layer0_outputs(3471);
    outputs(7814) <= not((layer0_outputs(6595)) or (layer0_outputs(4408)));
    outputs(7815) <= not(layer0_outputs(2912));
    outputs(7816) <= not(layer0_outputs(7702));
    outputs(7817) <= not(layer0_outputs(4175));
    outputs(7818) <= (layer0_outputs(10746)) xor (layer0_outputs(11479));
    outputs(7819) <= layer0_outputs(8901);
    outputs(7820) <= not(layer0_outputs(5795)) or (layer0_outputs(7809));
    outputs(7821) <= layer0_outputs(5804);
    outputs(7822) <= layer0_outputs(2516);
    outputs(7823) <= layer0_outputs(4730);
    outputs(7824) <= not(layer0_outputs(4329)) or (layer0_outputs(2374));
    outputs(7825) <= not(layer0_outputs(2168));
    outputs(7826) <= (layer0_outputs(8027)) and not (layer0_outputs(2388));
    outputs(7827) <= layer0_outputs(9184);
    outputs(7828) <= layer0_outputs(3922);
    outputs(7829) <= not(layer0_outputs(1317));
    outputs(7830) <= layer0_outputs(12628);
    outputs(7831) <= not((layer0_outputs(6522)) xor (layer0_outputs(11967)));
    outputs(7832) <= not((layer0_outputs(4028)) xor (layer0_outputs(10733)));
    outputs(7833) <= (layer0_outputs(7232)) and not (layer0_outputs(5464));
    outputs(7834) <= layer0_outputs(2812);
    outputs(7835) <= (layer0_outputs(8930)) xor (layer0_outputs(12604));
    outputs(7836) <= not(layer0_outputs(1440));
    outputs(7837) <= layer0_outputs(6842);
    outputs(7838) <= (layer0_outputs(3558)) xor (layer0_outputs(1875));
    outputs(7839) <= not(layer0_outputs(8123));
    outputs(7840) <= not(layer0_outputs(9930));
    outputs(7841) <= layer0_outputs(8202);
    outputs(7842) <= layer0_outputs(12205);
    outputs(7843) <= not((layer0_outputs(11840)) xor (layer0_outputs(2306)));
    outputs(7844) <= not((layer0_outputs(11480)) or (layer0_outputs(5437)));
    outputs(7845) <= (layer0_outputs(10451)) xor (layer0_outputs(10948));
    outputs(7846) <= layer0_outputs(6297);
    outputs(7847) <= not(layer0_outputs(12546));
    outputs(7848) <= (layer0_outputs(1867)) and not (layer0_outputs(8515));
    outputs(7849) <= not(layer0_outputs(2159)) or (layer0_outputs(3876));
    outputs(7850) <= layer0_outputs(2596);
    outputs(7851) <= layer0_outputs(8307);
    outputs(7852) <= layer0_outputs(9183);
    outputs(7853) <= not(layer0_outputs(834));
    outputs(7854) <= (layer0_outputs(12510)) xor (layer0_outputs(2577));
    outputs(7855) <= not(layer0_outputs(6804));
    outputs(7856) <= not((layer0_outputs(4378)) xor (layer0_outputs(247)));
    outputs(7857) <= not((layer0_outputs(7194)) or (layer0_outputs(6416)));
    outputs(7858) <= not(layer0_outputs(5821));
    outputs(7859) <= not((layer0_outputs(8091)) or (layer0_outputs(7242)));
    outputs(7860) <= not((layer0_outputs(11627)) or (layer0_outputs(9220)));
    outputs(7861) <= not((layer0_outputs(11002)) xor (layer0_outputs(6475)));
    outputs(7862) <= not(layer0_outputs(2366));
    outputs(7863) <= (layer0_outputs(10787)) and (layer0_outputs(6349));
    outputs(7864) <= not((layer0_outputs(11069)) xor (layer0_outputs(704)));
    outputs(7865) <= not(layer0_outputs(186));
    outputs(7866) <= not(layer0_outputs(4492));
    outputs(7867) <= not(layer0_outputs(8457));
    outputs(7868) <= (layer0_outputs(12338)) and not (layer0_outputs(2560));
    outputs(7869) <= (layer0_outputs(2083)) or (layer0_outputs(2450));
    outputs(7870) <= not(layer0_outputs(831));
    outputs(7871) <= (layer0_outputs(11875)) xor (layer0_outputs(4929));
    outputs(7872) <= (layer0_outputs(4510)) xor (layer0_outputs(10674));
    outputs(7873) <= not(layer0_outputs(9126)) or (layer0_outputs(9597));
    outputs(7874) <= layer0_outputs(1220);
    outputs(7875) <= layer0_outputs(12525);
    outputs(7876) <= layer0_outputs(1134);
    outputs(7877) <= (layer0_outputs(4520)) xor (layer0_outputs(8834));
    outputs(7878) <= not((layer0_outputs(6495)) xor (layer0_outputs(1955)));
    outputs(7879) <= not(layer0_outputs(4038));
    outputs(7880) <= (layer0_outputs(8881)) xor (layer0_outputs(6110));
    outputs(7881) <= not((layer0_outputs(8057)) xor (layer0_outputs(3435)));
    outputs(7882) <= not(layer0_outputs(4454));
    outputs(7883) <= not(layer0_outputs(5590));
    outputs(7884) <= not((layer0_outputs(5193)) and (layer0_outputs(9788)));
    outputs(7885) <= not(layer0_outputs(10582));
    outputs(7886) <= layer0_outputs(7471);
    outputs(7887) <= not(layer0_outputs(5443));
    outputs(7888) <= (layer0_outputs(12087)) and not (layer0_outputs(919));
    outputs(7889) <= not(layer0_outputs(11989));
    outputs(7890) <= not((layer0_outputs(5398)) or (layer0_outputs(9714)));
    outputs(7891) <= not((layer0_outputs(4306)) xor (layer0_outputs(6108)));
    outputs(7892) <= not((layer0_outputs(9983)) xor (layer0_outputs(1758)));
    outputs(7893) <= layer0_outputs(8056);
    outputs(7894) <= not(layer0_outputs(3495));
    outputs(7895) <= (layer0_outputs(6542)) and (layer0_outputs(7665));
    outputs(7896) <= layer0_outputs(10715);
    outputs(7897) <= (layer0_outputs(2533)) xor (layer0_outputs(12343));
    outputs(7898) <= not(layer0_outputs(4875));
    outputs(7899) <= not(layer0_outputs(4983));
    outputs(7900) <= (layer0_outputs(6446)) or (layer0_outputs(11625));
    outputs(7901) <= layer0_outputs(6608);
    outputs(7902) <= not(layer0_outputs(5935));
    outputs(7903) <= (layer0_outputs(672)) and not (layer0_outputs(7942));
    outputs(7904) <= not(layer0_outputs(2853));
    outputs(7905) <= not((layer0_outputs(1989)) xor (layer0_outputs(10614)));
    outputs(7906) <= not((layer0_outputs(6893)) or (layer0_outputs(7756)));
    outputs(7907) <= not(layer0_outputs(3351));
    outputs(7908) <= layer0_outputs(1371);
    outputs(7909) <= layer0_outputs(1594);
    outputs(7910) <= not((layer0_outputs(7373)) and (layer0_outputs(5924)));
    outputs(7911) <= not(layer0_outputs(2691)) or (layer0_outputs(8951));
    outputs(7912) <= not(layer0_outputs(7961));
    outputs(7913) <= not(layer0_outputs(8362)) or (layer0_outputs(11437));
    outputs(7914) <= (layer0_outputs(1996)) and not (layer0_outputs(3871));
    outputs(7915) <= not((layer0_outputs(9233)) xor (layer0_outputs(9579)));
    outputs(7916) <= not((layer0_outputs(4146)) or (layer0_outputs(4411)));
    outputs(7917) <= not(layer0_outputs(4550));
    outputs(7918) <= layer0_outputs(5835);
    outputs(7919) <= not((layer0_outputs(4108)) xor (layer0_outputs(11034)));
    outputs(7920) <= not(layer0_outputs(12417));
    outputs(7921) <= not((layer0_outputs(4638)) xor (layer0_outputs(2639)));
    outputs(7922) <= layer0_outputs(11189);
    outputs(7923) <= not(layer0_outputs(12130));
    outputs(7924) <= not(layer0_outputs(2770));
    outputs(7925) <= (layer0_outputs(9628)) xor (layer0_outputs(12268));
    outputs(7926) <= layer0_outputs(11074);
    outputs(7927) <= not((layer0_outputs(252)) xor (layer0_outputs(6121)));
    outputs(7928) <= not(layer0_outputs(7311));
    outputs(7929) <= not(layer0_outputs(8466));
    outputs(7930) <= (layer0_outputs(12125)) and not (layer0_outputs(7284));
    outputs(7931) <= layer0_outputs(8722);
    outputs(7932) <= not((layer0_outputs(9857)) xor (layer0_outputs(9155)));
    outputs(7933) <= (layer0_outputs(965)) and not (layer0_outputs(2758));
    outputs(7934) <= not(layer0_outputs(7138));
    outputs(7935) <= layer0_outputs(1255);
    outputs(7936) <= not(layer0_outputs(11549));
    outputs(7937) <= (layer0_outputs(10607)) xor (layer0_outputs(860));
    outputs(7938) <= layer0_outputs(74);
    outputs(7939) <= (layer0_outputs(2625)) or (layer0_outputs(7116));
    outputs(7940) <= not(layer0_outputs(3845));
    outputs(7941) <= layer0_outputs(10243);
    outputs(7942) <= layer0_outputs(5203);
    outputs(7943) <= layer0_outputs(12441);
    outputs(7944) <= layer0_outputs(10572);
    outputs(7945) <= (layer0_outputs(356)) and not (layer0_outputs(11699));
    outputs(7946) <= layer0_outputs(6573);
    outputs(7947) <= not((layer0_outputs(8741)) or (layer0_outputs(4232)));
    outputs(7948) <= (layer0_outputs(258)) xor (layer0_outputs(12128));
    outputs(7949) <= not(layer0_outputs(8359));
    outputs(7950) <= not(layer0_outputs(10716));
    outputs(7951) <= not(layer0_outputs(7456));
    outputs(7952) <= not((layer0_outputs(7788)) or (layer0_outputs(7067)));
    outputs(7953) <= (layer0_outputs(1208)) xor (layer0_outputs(2763));
    outputs(7954) <= not(layer0_outputs(6984));
    outputs(7955) <= layer0_outputs(275);
    outputs(7956) <= not((layer0_outputs(3364)) xor (layer0_outputs(3914)));
    outputs(7957) <= layer0_outputs(2400);
    outputs(7958) <= not((layer0_outputs(1130)) xor (layer0_outputs(8099)));
    outputs(7959) <= (layer0_outputs(8844)) xor (layer0_outputs(7802));
    outputs(7960) <= not((layer0_outputs(6709)) xor (layer0_outputs(5928)));
    outputs(7961) <= not(layer0_outputs(3462)) or (layer0_outputs(8543));
    outputs(7962) <= not((layer0_outputs(2610)) xor (layer0_outputs(1623)));
    outputs(7963) <= not(layer0_outputs(8337));
    outputs(7964) <= (layer0_outputs(7170)) and not (layer0_outputs(4118));
    outputs(7965) <= (layer0_outputs(480)) and not (layer0_outputs(2178));
    outputs(7966) <= (layer0_outputs(5996)) xor (layer0_outputs(1382));
    outputs(7967) <= not((layer0_outputs(10827)) or (layer0_outputs(8805)));
    outputs(7968) <= not(layer0_outputs(12146));
    outputs(7969) <= not((layer0_outputs(11661)) or (layer0_outputs(3931)));
    outputs(7970) <= not(layer0_outputs(1483));
    outputs(7971) <= layer0_outputs(10693);
    outputs(7972) <= not(layer0_outputs(12438));
    outputs(7973) <= not(layer0_outputs(2738)) or (layer0_outputs(6470));
    outputs(7974) <= (layer0_outputs(11291)) and not (layer0_outputs(12629));
    outputs(7975) <= (layer0_outputs(10714)) or (layer0_outputs(5890));
    outputs(7976) <= not((layer0_outputs(9476)) xor (layer0_outputs(5614)));
    outputs(7977) <= not((layer0_outputs(5744)) or (layer0_outputs(8713)));
    outputs(7978) <= (layer0_outputs(3248)) and not (layer0_outputs(5746));
    outputs(7979) <= not(layer0_outputs(817)) or (layer0_outputs(9426));
    outputs(7980) <= not(layer0_outputs(3009));
    outputs(7981) <= not(layer0_outputs(4656));
    outputs(7982) <= not(layer0_outputs(11109)) or (layer0_outputs(9552));
    outputs(7983) <= layer0_outputs(7851);
    outputs(7984) <= layer0_outputs(8606);
    outputs(7985) <= not(layer0_outputs(193));
    outputs(7986) <= not((layer0_outputs(4608)) and (layer0_outputs(2845)));
    outputs(7987) <= (layer0_outputs(3161)) and not (layer0_outputs(10516));
    outputs(7988) <= not(layer0_outputs(3147)) or (layer0_outputs(12203));
    outputs(7989) <= not(layer0_outputs(5441));
    outputs(7990) <= layer0_outputs(3049);
    outputs(7991) <= not((layer0_outputs(868)) xor (layer0_outputs(7059)));
    outputs(7992) <= (layer0_outputs(11424)) xor (layer0_outputs(770));
    outputs(7993) <= layer0_outputs(12179);
    outputs(7994) <= layer0_outputs(7172);
    outputs(7995) <= (layer0_outputs(6838)) xor (layer0_outputs(5568));
    outputs(7996) <= layer0_outputs(11380);
    outputs(7997) <= (layer0_outputs(9688)) xor (layer0_outputs(5093));
    outputs(7998) <= layer0_outputs(5489);
    outputs(7999) <= not((layer0_outputs(11931)) xor (layer0_outputs(1374)));
    outputs(8000) <= layer0_outputs(11919);
    outputs(8001) <= (layer0_outputs(6679)) xor (layer0_outputs(5134));
    outputs(8002) <= layer0_outputs(3960);
    outputs(8003) <= (layer0_outputs(7171)) xor (layer0_outputs(9408));
    outputs(8004) <= not(layer0_outputs(6779));
    outputs(8005) <= (layer0_outputs(926)) and not (layer0_outputs(9107));
    outputs(8006) <= layer0_outputs(8374);
    outputs(8007) <= not(layer0_outputs(2484));
    outputs(8008) <= layer0_outputs(10175);
    outputs(8009) <= (layer0_outputs(925)) and (layer0_outputs(1230));
    outputs(8010) <= layer0_outputs(8619);
    outputs(8011) <= not((layer0_outputs(9116)) or (layer0_outputs(1618)));
    outputs(8012) <= (layer0_outputs(11284)) xor (layer0_outputs(4902));
    outputs(8013) <= not(layer0_outputs(3575));
    outputs(8014) <= not((layer0_outputs(292)) or (layer0_outputs(6330)));
    outputs(8015) <= layer0_outputs(7968);
    outputs(8016) <= not(layer0_outputs(9678)) or (layer0_outputs(1277));
    outputs(8017) <= not(layer0_outputs(12783));
    outputs(8018) <= not(layer0_outputs(7015)) or (layer0_outputs(471));
    outputs(8019) <= not(layer0_outputs(12589)) or (layer0_outputs(8851));
    outputs(8020) <= layer0_outputs(8685);
    outputs(8021) <= not(layer0_outputs(7734));
    outputs(8022) <= not(layer0_outputs(9033));
    outputs(8023) <= (layer0_outputs(11073)) xor (layer0_outputs(5137));
    outputs(8024) <= (layer0_outputs(6655)) xor (layer0_outputs(7107));
    outputs(8025) <= not(layer0_outputs(9190));
    outputs(8026) <= not(layer0_outputs(9389));
    outputs(8027) <= layer0_outputs(1082);
    outputs(8028) <= layer0_outputs(11748);
    outputs(8029) <= not(layer0_outputs(11579));
    outputs(8030) <= not((layer0_outputs(9591)) or (layer0_outputs(6512)));
    outputs(8031) <= not(layer0_outputs(3370));
    outputs(8032) <= not(layer0_outputs(8897));
    outputs(8033) <= not(layer0_outputs(12358));
    outputs(8034) <= not(layer0_outputs(1925));
    outputs(8035) <= not(layer0_outputs(12386));
    outputs(8036) <= layer0_outputs(6345);
    outputs(8037) <= layer0_outputs(5243);
    outputs(8038) <= (layer0_outputs(9241)) or (layer0_outputs(4039));
    outputs(8039) <= not(layer0_outputs(6294));
    outputs(8040) <= (layer0_outputs(10596)) and not (layer0_outputs(4308));
    outputs(8041) <= not(layer0_outputs(3536));
    outputs(8042) <= not((layer0_outputs(7217)) or (layer0_outputs(11483)));
    outputs(8043) <= not((layer0_outputs(10620)) or (layer0_outputs(1186)));
    outputs(8044) <= not(layer0_outputs(3283));
    outputs(8045) <= (layer0_outputs(8016)) xor (layer0_outputs(308));
    outputs(8046) <= (layer0_outputs(5110)) xor (layer0_outputs(9032));
    outputs(8047) <= not(layer0_outputs(2444)) or (layer0_outputs(9446));
    outputs(8048) <= not(layer0_outputs(4061)) or (layer0_outputs(3732));
    outputs(8049) <= (layer0_outputs(3203)) or (layer0_outputs(5983));
    outputs(8050) <= not(layer0_outputs(3305));
    outputs(8051) <= layer0_outputs(4839);
    outputs(8052) <= not(layer0_outputs(882));
    outputs(8053) <= layer0_outputs(12554);
    outputs(8054) <= (layer0_outputs(5460)) or (layer0_outputs(1058));
    outputs(8055) <= (layer0_outputs(741)) and not (layer0_outputs(3301));
    outputs(8056) <= not(layer0_outputs(2478));
    outputs(8057) <= not((layer0_outputs(6712)) xor (layer0_outputs(6930)));
    outputs(8058) <= layer0_outputs(11878);
    outputs(8059) <= (layer0_outputs(5480)) and (layer0_outputs(12576));
    outputs(8060) <= not(layer0_outputs(7709));
    outputs(8061) <= not(layer0_outputs(8856));
    outputs(8062) <= layer0_outputs(1016);
    outputs(8063) <= (layer0_outputs(5577)) and (layer0_outputs(11287));
    outputs(8064) <= not((layer0_outputs(8697)) or (layer0_outputs(1651)));
    outputs(8065) <= layer0_outputs(2553);
    outputs(8066) <= layer0_outputs(4052);
    outputs(8067) <= (layer0_outputs(5278)) and not (layer0_outputs(3338));
    outputs(8068) <= layer0_outputs(4019);
    outputs(8069) <= not(layer0_outputs(6413));
    outputs(8070) <= not(layer0_outputs(3897));
    outputs(8071) <= not(layer0_outputs(2547)) or (layer0_outputs(6012));
    outputs(8072) <= layer0_outputs(6326);
    outputs(8073) <= not(layer0_outputs(10258));
    outputs(8074) <= not(layer0_outputs(856));
    outputs(8075) <= (layer0_outputs(8234)) xor (layer0_outputs(6033));
    outputs(8076) <= not(layer0_outputs(3688));
    outputs(8077) <= not((layer0_outputs(7098)) or (layer0_outputs(107)));
    outputs(8078) <= layer0_outputs(1684);
    outputs(8079) <= layer0_outputs(8731);
    outputs(8080) <= not((layer0_outputs(3734)) xor (layer0_outputs(5490)));
    outputs(8081) <= not(layer0_outputs(1170)) or (layer0_outputs(702));
    outputs(8082) <= not(layer0_outputs(10125));
    outputs(8083) <= (layer0_outputs(9781)) and not (layer0_outputs(10880));
    outputs(8084) <= not(layer0_outputs(5372));
    outputs(8085) <= layer0_outputs(111);
    outputs(8086) <= layer0_outputs(47);
    outputs(8087) <= layer0_outputs(1803);
    outputs(8088) <= (layer0_outputs(1932)) xor (layer0_outputs(11780));
    outputs(8089) <= not((layer0_outputs(300)) or (layer0_outputs(975)));
    outputs(8090) <= not(layer0_outputs(9621));
    outputs(8091) <= (layer0_outputs(4670)) xor (layer0_outputs(1167));
    outputs(8092) <= layer0_outputs(11866);
    outputs(8093) <= (layer0_outputs(1512)) xor (layer0_outputs(2443));
    outputs(8094) <= (layer0_outputs(7354)) and not (layer0_outputs(4925));
    outputs(8095) <= layer0_outputs(10152);
    outputs(8096) <= layer0_outputs(4749);
    outputs(8097) <= layer0_outputs(4465);
    outputs(8098) <= not(layer0_outputs(4285));
    outputs(8099) <= layer0_outputs(9660);
    outputs(8100) <= not(layer0_outputs(11681));
    outputs(8101) <= not((layer0_outputs(7111)) or (layer0_outputs(7267)));
    outputs(8102) <= not(layer0_outputs(11510));
    outputs(8103) <= (layer0_outputs(10753)) and (layer0_outputs(8443));
    outputs(8104) <= not(layer0_outputs(7874));
    outputs(8105) <= layer0_outputs(1932);
    outputs(8106) <= layer0_outputs(7054);
    outputs(8107) <= not((layer0_outputs(11859)) or (layer0_outputs(9506)));
    outputs(8108) <= layer0_outputs(12542);
    outputs(8109) <= layer0_outputs(8942);
    outputs(8110) <= not((layer0_outputs(12266)) xor (layer0_outputs(8036)));
    outputs(8111) <= layer0_outputs(11344);
    outputs(8112) <= not((layer0_outputs(4301)) xor (layer0_outputs(4632)));
    outputs(8113) <= layer0_outputs(4361);
    outputs(8114) <= not((layer0_outputs(1189)) or (layer0_outputs(2573)));
    outputs(8115) <= layer0_outputs(6418);
    outputs(8116) <= (layer0_outputs(12109)) or (layer0_outputs(10727));
    outputs(8117) <= not((layer0_outputs(10457)) and (layer0_outputs(4273)));
    outputs(8118) <= not((layer0_outputs(5865)) and (layer0_outputs(1043)));
    outputs(8119) <= layer0_outputs(11906);
    outputs(8120) <= not((layer0_outputs(11331)) or (layer0_outputs(0)));
    outputs(8121) <= not(layer0_outputs(1068));
    outputs(8122) <= layer0_outputs(8333);
    outputs(8123) <= (layer0_outputs(2933)) xor (layer0_outputs(9564));
    outputs(8124) <= not((layer0_outputs(6673)) and (layer0_outputs(11040)));
    outputs(8125) <= (layer0_outputs(11575)) and (layer0_outputs(11749));
    outputs(8126) <= layer0_outputs(11750);
    outputs(8127) <= layer0_outputs(7858);
    outputs(8128) <= (layer0_outputs(10293)) or (layer0_outputs(12078));
    outputs(8129) <= not(layer0_outputs(2045)) or (layer0_outputs(10673));
    outputs(8130) <= layer0_outputs(6634);
    outputs(8131) <= layer0_outputs(11143);
    outputs(8132) <= not(layer0_outputs(4613));
    outputs(8133) <= layer0_outputs(7181);
    outputs(8134) <= not(layer0_outputs(5811));
    outputs(8135) <= not(layer0_outputs(7174));
    outputs(8136) <= not(layer0_outputs(6736));
    outputs(8137) <= not(layer0_outputs(10571));
    outputs(8138) <= (layer0_outputs(1366)) and not (layer0_outputs(3652));
    outputs(8139) <= not(layer0_outputs(11087));
    outputs(8140) <= (layer0_outputs(11173)) xor (layer0_outputs(79));
    outputs(8141) <= not((layer0_outputs(12006)) xor (layer0_outputs(6216)));
    outputs(8142) <= layer0_outputs(787);
    outputs(8143) <= layer0_outputs(9238);
    outputs(8144) <= not(layer0_outputs(1936));
    outputs(8145) <= not(layer0_outputs(7419)) or (layer0_outputs(8194));
    outputs(8146) <= not((layer0_outputs(4300)) and (layer0_outputs(9461)));
    outputs(8147) <= (layer0_outputs(4479)) xor (layer0_outputs(7746));
    outputs(8148) <= not((layer0_outputs(768)) or (layer0_outputs(6858)));
    outputs(8149) <= layer0_outputs(2887);
    outputs(8150) <= not((layer0_outputs(2782)) xor (layer0_outputs(10711)));
    outputs(8151) <= layer0_outputs(5573);
    outputs(8152) <= not((layer0_outputs(1013)) xor (layer0_outputs(11966)));
    outputs(8153) <= (layer0_outputs(1505)) xor (layer0_outputs(481));
    outputs(8154) <= (layer0_outputs(10580)) and (layer0_outputs(11244));
    outputs(8155) <= (layer0_outputs(6593)) and not (layer0_outputs(9072));
    outputs(8156) <= layer0_outputs(10211);
    outputs(8157) <= (layer0_outputs(5308)) and not (layer0_outputs(6405));
    outputs(8158) <= not(layer0_outputs(8653));
    outputs(8159) <= not(layer0_outputs(1579));
    outputs(8160) <= (layer0_outputs(8150)) and (layer0_outputs(10330));
    outputs(8161) <= layer0_outputs(11818);
    outputs(8162) <= (layer0_outputs(2225)) xor (layer0_outputs(11473));
    outputs(8163) <= not(layer0_outputs(7930));
    outputs(8164) <= (layer0_outputs(11261)) and (layer0_outputs(1063));
    outputs(8165) <= not((layer0_outputs(1514)) or (layer0_outputs(811)));
    outputs(8166) <= not(layer0_outputs(7077)) or (layer0_outputs(7631));
    outputs(8167) <= (layer0_outputs(7821)) or (layer0_outputs(4944));
    outputs(8168) <= layer0_outputs(7300);
    outputs(8169) <= layer0_outputs(7312);
    outputs(8170) <= not(layer0_outputs(11580));
    outputs(8171) <= layer0_outputs(4135);
    outputs(8172) <= layer0_outputs(4559);
    outputs(8173) <= not(layer0_outputs(8818));
    outputs(8174) <= not((layer0_outputs(6451)) xor (layer0_outputs(4175)));
    outputs(8175) <= layer0_outputs(7732);
    outputs(8176) <= not(layer0_outputs(8891));
    outputs(8177) <= not((layer0_outputs(386)) xor (layer0_outputs(158)));
    outputs(8178) <= not(layer0_outputs(11016));
    outputs(8179) <= layer0_outputs(43);
    outputs(8180) <= not(layer0_outputs(4941));
    outputs(8181) <= layer0_outputs(10406);
    outputs(8182) <= layer0_outputs(4450);
    outputs(8183) <= (layer0_outputs(10215)) and not (layer0_outputs(5793));
    outputs(8184) <= not((layer0_outputs(4731)) xor (layer0_outputs(12537)));
    outputs(8185) <= (layer0_outputs(4974)) and not (layer0_outputs(12756));
    outputs(8186) <= (layer0_outputs(9082)) and not (layer0_outputs(11013));
    outputs(8187) <= layer0_outputs(154);
    outputs(8188) <= (layer0_outputs(8061)) and not (layer0_outputs(5397));
    outputs(8189) <= (layer0_outputs(4372)) xor (layer0_outputs(7843));
    outputs(8190) <= not(layer0_outputs(2497));
    outputs(8191) <= not(layer0_outputs(7286));
    outputs(8192) <= (layer0_outputs(3379)) and (layer0_outputs(11348));
    outputs(8193) <= not(layer0_outputs(5624));
    outputs(8194) <= (layer0_outputs(12186)) xor (layer0_outputs(12155));
    outputs(8195) <= not((layer0_outputs(7442)) or (layer0_outputs(12055)));
    outputs(8196) <= not(layer0_outputs(1215));
    outputs(8197) <= not(layer0_outputs(2898));
    outputs(8198) <= (layer0_outputs(6538)) and not (layer0_outputs(5682));
    outputs(8199) <= (layer0_outputs(2818)) and (layer0_outputs(8529));
    outputs(8200) <= not((layer0_outputs(4196)) xor (layer0_outputs(1059)));
    outputs(8201) <= not(layer0_outputs(4845));
    outputs(8202) <= (layer0_outputs(7316)) and not (layer0_outputs(7063));
    outputs(8203) <= (layer0_outputs(10635)) and not (layer0_outputs(2658));
    outputs(8204) <= not((layer0_outputs(6983)) xor (layer0_outputs(5609)));
    outputs(8205) <= not(layer0_outputs(9749));
    outputs(8206) <= not((layer0_outputs(11940)) xor (layer0_outputs(12373)));
    outputs(8207) <= not((layer0_outputs(6708)) xor (layer0_outputs(8992)));
    outputs(8208) <= not(layer0_outputs(3738));
    outputs(8209) <= layer0_outputs(2223);
    outputs(8210) <= not(layer0_outputs(7889));
    outputs(8211) <= not(layer0_outputs(11869));
    outputs(8212) <= not(layer0_outputs(8598));
    outputs(8213) <= not((layer0_outputs(5236)) or (layer0_outputs(6496)));
    outputs(8214) <= not(layer0_outputs(7365));
    outputs(8215) <= layer0_outputs(8711);
    outputs(8216) <= not(layer0_outputs(1437));
    outputs(8217) <= layer0_outputs(5015);
    outputs(8218) <= not(layer0_outputs(5548));
    outputs(8219) <= not(layer0_outputs(3425));
    outputs(8220) <= layer0_outputs(2747);
    outputs(8221) <= not(layer0_outputs(9486));
    outputs(8222) <= layer0_outputs(1303);
    outputs(8223) <= not(layer0_outputs(10610));
    outputs(8224) <= not((layer0_outputs(3430)) xor (layer0_outputs(1689)));
    outputs(8225) <= layer0_outputs(11179);
    outputs(8226) <= not((layer0_outputs(10430)) xor (layer0_outputs(9419)));
    outputs(8227) <= (layer0_outputs(10295)) and (layer0_outputs(9794));
    outputs(8228) <= not((layer0_outputs(10021)) or (layer0_outputs(4779)));
    outputs(8229) <= not(layer0_outputs(12717)) or (layer0_outputs(11585));
    outputs(8230) <= not(layer0_outputs(2259)) or (layer0_outputs(11361));
    outputs(8231) <= not(layer0_outputs(5830));
    outputs(8232) <= (layer0_outputs(11159)) and (layer0_outputs(11617));
    outputs(8233) <= not(layer0_outputs(7963));
    outputs(8234) <= not(layer0_outputs(1215));
    outputs(8235) <= not(layer0_outputs(10545));
    outputs(8236) <= (layer0_outputs(2955)) or (layer0_outputs(1878));
    outputs(8237) <= (layer0_outputs(9812)) xor (layer0_outputs(1217));
    outputs(8238) <= not(layer0_outputs(9633));
    outputs(8239) <= not(layer0_outputs(3648));
    outputs(8240) <= not(layer0_outputs(890));
    outputs(8241) <= not((layer0_outputs(11637)) xor (layer0_outputs(8268)));
    outputs(8242) <= not(layer0_outputs(4068));
    outputs(8243) <= layer0_outputs(10774);
    outputs(8244) <= not(layer0_outputs(1553)) or (layer0_outputs(1335));
    outputs(8245) <= not((layer0_outputs(6195)) or (layer0_outputs(14)));
    outputs(8246) <= layer0_outputs(6265);
    outputs(8247) <= (layer0_outputs(9183)) xor (layer0_outputs(4384));
    outputs(8248) <= not((layer0_outputs(10271)) xor (layer0_outputs(2521)));
    outputs(8249) <= not((layer0_outputs(11470)) xor (layer0_outputs(9362)));
    outputs(8250) <= not(layer0_outputs(11249));
    outputs(8251) <= not((layer0_outputs(9188)) xor (layer0_outputs(761)));
    outputs(8252) <= (layer0_outputs(1537)) and (layer0_outputs(6587));
    outputs(8253) <= not(layer0_outputs(12714));
    outputs(8254) <= not(layer0_outputs(7161));
    outputs(8255) <= layer0_outputs(7203);
    outputs(8256) <= not((layer0_outputs(1777)) or (layer0_outputs(6589)));
    outputs(8257) <= (layer0_outputs(11914)) and (layer0_outputs(6314));
    outputs(8258) <= layer0_outputs(4521);
    outputs(8259) <= (layer0_outputs(491)) xor (layer0_outputs(2910));
    outputs(8260) <= layer0_outputs(10892);
    outputs(8261) <= not(layer0_outputs(7423));
    outputs(8262) <= (layer0_outputs(2643)) and (layer0_outputs(8015));
    outputs(8263) <= not((layer0_outputs(9399)) xor (layer0_outputs(384)));
    outputs(8264) <= not(layer0_outputs(7390));
    outputs(8265) <= layer0_outputs(8959);
    outputs(8266) <= not(layer0_outputs(184));
    outputs(8267) <= layer0_outputs(10734);
    outputs(8268) <= layer0_outputs(6469);
    outputs(8269) <= (layer0_outputs(11006)) xor (layer0_outputs(8162));
    outputs(8270) <= (layer0_outputs(10103)) and not (layer0_outputs(8636));
    outputs(8271) <= (layer0_outputs(8258)) and (layer0_outputs(2148));
    outputs(8272) <= not((layer0_outputs(8947)) or (layer0_outputs(5522)));
    outputs(8273) <= not((layer0_outputs(8624)) xor (layer0_outputs(8353)));
    outputs(8274) <= not(layer0_outputs(2203));
    outputs(8275) <= layer0_outputs(1473);
    outputs(8276) <= layer0_outputs(8104);
    outputs(8277) <= not((layer0_outputs(11492)) and (layer0_outputs(4748)));
    outputs(8278) <= layer0_outputs(12074);
    outputs(8279) <= layer0_outputs(10019);
    outputs(8280) <= layer0_outputs(8797);
    outputs(8281) <= layer0_outputs(8690);
    outputs(8282) <= layer0_outputs(10490);
    outputs(8283) <= not((layer0_outputs(7484)) or (layer0_outputs(10980)));
    outputs(8284) <= not(layer0_outputs(4525));
    outputs(8285) <= layer0_outputs(6931);
    outputs(8286) <= not((layer0_outputs(1936)) xor (layer0_outputs(3367)));
    outputs(8287) <= not(layer0_outputs(5739));
    outputs(8288) <= not(layer0_outputs(2213));
    outputs(8289) <= not((layer0_outputs(2212)) or (layer0_outputs(9523)));
    outputs(8290) <= not(layer0_outputs(9915));
    outputs(8291) <= (layer0_outputs(9061)) and (layer0_outputs(3236));
    outputs(8292) <= not((layer0_outputs(934)) xor (layer0_outputs(3644)));
    outputs(8293) <= (layer0_outputs(5022)) and (layer0_outputs(4671));
    outputs(8294) <= not(layer0_outputs(3221));
    outputs(8295) <= not(layer0_outputs(4103));
    outputs(8296) <= not(layer0_outputs(10187));
    outputs(8297) <= not(layer0_outputs(4613));
    outputs(8298) <= (layer0_outputs(1351)) xor (layer0_outputs(12356));
    outputs(8299) <= not(layer0_outputs(5612));
    outputs(8300) <= (layer0_outputs(2997)) and not (layer0_outputs(1479));
    outputs(8301) <= not(layer0_outputs(7494));
    outputs(8302) <= layer0_outputs(12725);
    outputs(8303) <= layer0_outputs(5589);
    outputs(8304) <= not(layer0_outputs(5219));
    outputs(8305) <= not(layer0_outputs(2844)) or (layer0_outputs(5319));
    outputs(8306) <= not(layer0_outputs(255));
    outputs(8307) <= not(layer0_outputs(11368));
    outputs(8308) <= layer0_outputs(1834);
    outputs(8309) <= not(layer0_outputs(10687));
    outputs(8310) <= not(layer0_outputs(464));
    outputs(8311) <= not(layer0_outputs(7174));
    outputs(8312) <= layer0_outputs(12654);
    outputs(8313) <= layer0_outputs(11950);
    outputs(8314) <= layer0_outputs(4725);
    outputs(8315) <= layer0_outputs(11160);
    outputs(8316) <= layer0_outputs(11085);
    outputs(8317) <= not(layer0_outputs(7712));
    outputs(8318) <= not(layer0_outputs(3824));
    outputs(8319) <= (layer0_outputs(9612)) or (layer0_outputs(11252));
    outputs(8320) <= layer0_outputs(248);
    outputs(8321) <= (layer0_outputs(2190)) and not (layer0_outputs(6494));
    outputs(8322) <= not((layer0_outputs(479)) or (layer0_outputs(4267)));
    outputs(8323) <= not(layer0_outputs(374));
    outputs(8324) <= not(layer0_outputs(10311));
    outputs(8325) <= (layer0_outputs(8388)) and not (layer0_outputs(6006));
    outputs(8326) <= (layer0_outputs(9442)) xor (layer0_outputs(1590));
    outputs(8327) <= (layer0_outputs(389)) and not (layer0_outputs(6103));
    outputs(8328) <= not(layer0_outputs(11943));
    outputs(8329) <= not(layer0_outputs(2679));
    outputs(8330) <= layer0_outputs(12100);
    outputs(8331) <= (layer0_outputs(5258)) and not (layer0_outputs(8853));
    outputs(8332) <= layer0_outputs(8814);
    outputs(8333) <= not((layer0_outputs(4910)) or (layer0_outputs(12277)));
    outputs(8334) <= layer0_outputs(1691);
    outputs(8335) <= not(layer0_outputs(5753)) or (layer0_outputs(2896));
    outputs(8336) <= (layer0_outputs(9405)) and (layer0_outputs(4397));
    outputs(8337) <= layer0_outputs(2136);
    outputs(8338) <= not(layer0_outputs(12579)) or (layer0_outputs(563));
    outputs(8339) <= not(layer0_outputs(190));
    outputs(8340) <= not(layer0_outputs(829));
    outputs(8341) <= (layer0_outputs(2654)) xor (layer0_outputs(3565));
    outputs(8342) <= layer0_outputs(1194);
    outputs(8343) <= not(layer0_outputs(644));
    outputs(8344) <= (layer0_outputs(10234)) xor (layer0_outputs(12631));
    outputs(8345) <= not((layer0_outputs(1180)) or (layer0_outputs(2527)));
    outputs(8346) <= not((layer0_outputs(6865)) or (layer0_outputs(10452)));
    outputs(8347) <= not((layer0_outputs(5680)) xor (layer0_outputs(5880)));
    outputs(8348) <= layer0_outputs(8938);
    outputs(8349) <= (layer0_outputs(6242)) xor (layer0_outputs(2812));
    outputs(8350) <= not((layer0_outputs(5241)) and (layer0_outputs(4794)));
    outputs(8351) <= not((layer0_outputs(429)) or (layer0_outputs(8450)));
    outputs(8352) <= not((layer0_outputs(503)) and (layer0_outputs(12578)));
    outputs(8353) <= not(layer0_outputs(8452));
    outputs(8354) <= layer0_outputs(2536);
    outputs(8355) <= not(layer0_outputs(4907));
    outputs(8356) <= layer0_outputs(766);
    outputs(8357) <= layer0_outputs(12032);
    outputs(8358) <= not((layer0_outputs(7892)) and (layer0_outputs(11058)));
    outputs(8359) <= layer0_outputs(8538);
    outputs(8360) <= not(layer0_outputs(1368));
    outputs(8361) <= not(layer0_outputs(1508)) or (layer0_outputs(1878));
    outputs(8362) <= (layer0_outputs(78)) and (layer0_outputs(8305));
    outputs(8363) <= not(layer0_outputs(4351));
    outputs(8364) <= (layer0_outputs(7857)) xor (layer0_outputs(11154));
    outputs(8365) <= not((layer0_outputs(5234)) xor (layer0_outputs(4523)));
    outputs(8366) <= not((layer0_outputs(9913)) xor (layer0_outputs(2538)));
    outputs(8367) <= not(layer0_outputs(7607));
    outputs(8368) <= not(layer0_outputs(768));
    outputs(8369) <= not(layer0_outputs(5016));
    outputs(8370) <= not((layer0_outputs(4786)) or (layer0_outputs(4427)));
    outputs(8371) <= layer0_outputs(11017);
    outputs(8372) <= not(layer0_outputs(6784));
    outputs(8373) <= not(layer0_outputs(1036));
    outputs(8374) <= (layer0_outputs(11528)) and (layer0_outputs(5514));
    outputs(8375) <= layer0_outputs(10019);
    outputs(8376) <= not(layer0_outputs(8574));
    outputs(8377) <= not(layer0_outputs(10782)) or (layer0_outputs(8642));
    outputs(8378) <= not(layer0_outputs(8351));
    outputs(8379) <= not((layer0_outputs(11123)) xor (layer0_outputs(129)));
    outputs(8380) <= not(layer0_outputs(3067));
    outputs(8381) <= not(layer0_outputs(10528));
    outputs(8382) <= not(layer0_outputs(986));
    outputs(8383) <= layer0_outputs(5589);
    outputs(8384) <= (layer0_outputs(8382)) xor (layer0_outputs(11157));
    outputs(8385) <= layer0_outputs(5143);
    outputs(8386) <= layer0_outputs(7650);
    outputs(8387) <= layer0_outputs(11425);
    outputs(8388) <= (layer0_outputs(3626)) and (layer0_outputs(9784));
    outputs(8389) <= not((layer0_outputs(11174)) xor (layer0_outputs(974)));
    outputs(8390) <= layer0_outputs(10564);
    outputs(8391) <= not(layer0_outputs(8520));
    outputs(8392) <= layer0_outputs(10360);
    outputs(8393) <= not(layer0_outputs(5468));
    outputs(8394) <= layer0_outputs(8474);
    outputs(8395) <= layer0_outputs(8023);
    outputs(8396) <= (layer0_outputs(2598)) xor (layer0_outputs(9413));
    outputs(8397) <= layer0_outputs(2096);
    outputs(8398) <= not((layer0_outputs(2248)) xor (layer0_outputs(2213)));
    outputs(8399) <= layer0_outputs(2144);
    outputs(8400) <= not(layer0_outputs(11122));
    outputs(8401) <= not((layer0_outputs(7366)) or (layer0_outputs(12728)));
    outputs(8402) <= (layer0_outputs(950)) xor (layer0_outputs(1506));
    outputs(8403) <= not(layer0_outputs(5492));
    outputs(8404) <= not((layer0_outputs(6948)) or (layer0_outputs(5263)));
    outputs(8405) <= not((layer0_outputs(11113)) xor (layer0_outputs(2714)));
    outputs(8406) <= layer0_outputs(6812);
    outputs(8407) <= (layer0_outputs(11838)) or (layer0_outputs(8656));
    outputs(8408) <= (layer0_outputs(9834)) and (layer0_outputs(6448));
    outputs(8409) <= layer0_outputs(6079);
    outputs(8410) <= not((layer0_outputs(12029)) xor (layer0_outputs(3756)));
    outputs(8411) <= not(layer0_outputs(9097));
    outputs(8412) <= (layer0_outputs(1450)) or (layer0_outputs(12242));
    outputs(8413) <= (layer0_outputs(1928)) xor (layer0_outputs(11487));
    outputs(8414) <= (layer0_outputs(10518)) and not (layer0_outputs(2390));
    outputs(8415) <= not(layer0_outputs(11611));
    outputs(8416) <= (layer0_outputs(12183)) xor (layer0_outputs(9934));
    outputs(8417) <= layer0_outputs(8458);
    outputs(8418) <= layer0_outputs(7377);
    outputs(8419) <= not(layer0_outputs(12419));
    outputs(8420) <= not(layer0_outputs(12147));
    outputs(8421) <= layer0_outputs(9947);
    outputs(8422) <= not(layer0_outputs(2343)) or (layer0_outputs(10536));
    outputs(8423) <= not((layer0_outputs(5032)) xor (layer0_outputs(4900)));
    outputs(8424) <= not(layer0_outputs(7753)) or (layer0_outputs(9036));
    outputs(8425) <= (layer0_outputs(6034)) and not (layer0_outputs(2065));
    outputs(8426) <= (layer0_outputs(9112)) xor (layer0_outputs(3601));
    outputs(8427) <= layer0_outputs(10805);
    outputs(8428) <= not((layer0_outputs(332)) xor (layer0_outputs(10875)));
    outputs(8429) <= not(layer0_outputs(5826));
    outputs(8430) <= layer0_outputs(11170);
    outputs(8431) <= layer0_outputs(7321);
    outputs(8432) <= (layer0_outputs(12377)) xor (layer0_outputs(4576));
    outputs(8433) <= (layer0_outputs(1670)) or (layer0_outputs(3474));
    outputs(8434) <= (layer0_outputs(11502)) xor (layer0_outputs(10492));
    outputs(8435) <= layer0_outputs(9068);
    outputs(8436) <= layer0_outputs(8793);
    outputs(8437) <= not(layer0_outputs(9900));
    outputs(8438) <= not(layer0_outputs(2218));
    outputs(8439) <= layer0_outputs(275);
    outputs(8440) <= not((layer0_outputs(6254)) xor (layer0_outputs(10524)));
    outputs(8441) <= not(layer0_outputs(8996));
    outputs(8442) <= not((layer0_outputs(8330)) or (layer0_outputs(11689)));
    outputs(8443) <= not((layer0_outputs(12442)) and (layer0_outputs(6307)));
    outputs(8444) <= not((layer0_outputs(9214)) and (layer0_outputs(4703)));
    outputs(8445) <= not((layer0_outputs(3988)) xor (layer0_outputs(4505)));
    outputs(8446) <= (layer0_outputs(5943)) and not (layer0_outputs(4874));
    outputs(8447) <= not((layer0_outputs(1340)) xor (layer0_outputs(10833)));
    outputs(8448) <= (layer0_outputs(12114)) xor (layer0_outputs(2644));
    outputs(8449) <= not(layer0_outputs(3907)) or (layer0_outputs(7711));
    outputs(8450) <= not((layer0_outputs(10050)) xor (layer0_outputs(11408)));
    outputs(8451) <= not(layer0_outputs(9911));
    outputs(8452) <= (layer0_outputs(9043)) or (layer0_outputs(12798));
    outputs(8453) <= not((layer0_outputs(1674)) and (layer0_outputs(9209)));
    outputs(8454) <= not((layer0_outputs(4751)) or (layer0_outputs(2253)));
    outputs(8455) <= not(layer0_outputs(6335));
    outputs(8456) <= (layer0_outputs(1413)) or (layer0_outputs(11665));
    outputs(8457) <= layer0_outputs(1584);
    outputs(8458) <= not((layer0_outputs(7453)) xor (layer0_outputs(3519)));
    outputs(8459) <= layer0_outputs(339);
    outputs(8460) <= not(layer0_outputs(10403));
    outputs(8461) <= not((layer0_outputs(3156)) xor (layer0_outputs(4819)));
    outputs(8462) <= layer0_outputs(5549);
    outputs(8463) <= not(layer0_outputs(2333));
    outputs(8464) <= layer0_outputs(5343);
    outputs(8465) <= (layer0_outputs(10742)) xor (layer0_outputs(5832));
    outputs(8466) <= (layer0_outputs(9255)) xor (layer0_outputs(4882));
    outputs(8467) <= not(layer0_outputs(4792));
    outputs(8468) <= not(layer0_outputs(4645)) or (layer0_outputs(11717));
    outputs(8469) <= not(layer0_outputs(127));
    outputs(8470) <= not(layer0_outputs(12291));
    outputs(8471) <= not(layer0_outputs(7090));
    outputs(8472) <= (layer0_outputs(5401)) and (layer0_outputs(3314));
    outputs(8473) <= (layer0_outputs(9404)) and not (layer0_outputs(5449));
    outputs(8474) <= layer0_outputs(4074);
    outputs(8475) <= not(layer0_outputs(798)) or (layer0_outputs(8261));
    outputs(8476) <= not(layer0_outputs(7621));
    outputs(8477) <= (layer0_outputs(6725)) and (layer0_outputs(6332));
    outputs(8478) <= layer0_outputs(1447);
    outputs(8479) <= layer0_outputs(736);
    outputs(8480) <= not(layer0_outputs(12212));
    outputs(8481) <= layer0_outputs(4328);
    outputs(8482) <= not(layer0_outputs(1524));
    outputs(8483) <= layer0_outputs(6809);
    outputs(8484) <= not(layer0_outputs(2344));
    outputs(8485) <= not((layer0_outputs(3456)) xor (layer0_outputs(6096)));
    outputs(8486) <= layer0_outputs(210);
    outputs(8487) <= layer0_outputs(5817);
    outputs(8488) <= not(layer0_outputs(5531));
    outputs(8489) <= not((layer0_outputs(5746)) or (layer0_outputs(3050)));
    outputs(8490) <= not(layer0_outputs(4724));
    outputs(8491) <= (layer0_outputs(5428)) xor (layer0_outputs(2097));
    outputs(8492) <= (layer0_outputs(8606)) and not (layer0_outputs(2600));
    outputs(8493) <= not(layer0_outputs(4007));
    outputs(8494) <= not(layer0_outputs(9865));
    outputs(8495) <= not(layer0_outputs(7845));
    outputs(8496) <= not(layer0_outputs(1858));
    outputs(8497) <= not(layer0_outputs(9930));
    outputs(8498) <= (layer0_outputs(5975)) and not (layer0_outputs(375));
    outputs(8499) <= (layer0_outputs(5204)) and not (layer0_outputs(8763));
    outputs(8500) <= not(layer0_outputs(3873));
    outputs(8501) <= (layer0_outputs(9645)) and not (layer0_outputs(2383));
    outputs(8502) <= not((layer0_outputs(9160)) and (layer0_outputs(10865)));
    outputs(8503) <= not(layer0_outputs(10868));
    outputs(8504) <= not(layer0_outputs(2985));
    outputs(8505) <= (layer0_outputs(9364)) or (layer0_outputs(12458));
    outputs(8506) <= not((layer0_outputs(10347)) xor (layer0_outputs(7501)));
    outputs(8507) <= not(layer0_outputs(12605));
    outputs(8508) <= not((layer0_outputs(6294)) or (layer0_outputs(7866)));
    outputs(8509) <= (layer0_outputs(740)) xor (layer0_outputs(3274));
    outputs(8510) <= layer0_outputs(9662);
    outputs(8511) <= not(layer0_outputs(2135)) or (layer0_outputs(1409));
    outputs(8512) <= (layer0_outputs(4112)) or (layer0_outputs(5440));
    outputs(8513) <= not((layer0_outputs(10053)) or (layer0_outputs(328)));
    outputs(8514) <= (layer0_outputs(11876)) and (layer0_outputs(5788));
    outputs(8515) <= not((layer0_outputs(2296)) and (layer0_outputs(8895)));
    outputs(8516) <= not(layer0_outputs(1520));
    outputs(8517) <= not(layer0_outputs(10678));
    outputs(8518) <= not(layer0_outputs(5275)) or (layer0_outputs(3369));
    outputs(8519) <= (layer0_outputs(12586)) xor (layer0_outputs(6652));
    outputs(8520) <= (layer0_outputs(716)) and (layer0_outputs(5618));
    outputs(8521) <= not((layer0_outputs(6717)) or (layer0_outputs(4007)));
    outputs(8522) <= (layer0_outputs(12132)) and (layer0_outputs(280));
    outputs(8523) <= (layer0_outputs(2287)) xor (layer0_outputs(7624));
    outputs(8524) <= (layer0_outputs(3745)) xor (layer0_outputs(8566));
    outputs(8525) <= layer0_outputs(7675);
    outputs(8526) <= not(layer0_outputs(3243));
    outputs(8527) <= not(layer0_outputs(5255));
    outputs(8528) <= layer0_outputs(10292);
    outputs(8529) <= (layer0_outputs(2256)) and (layer0_outputs(7342));
    outputs(8530) <= not(layer0_outputs(9153)) or (layer0_outputs(12175));
    outputs(8531) <= not(layer0_outputs(8391));
    outputs(8532) <= (layer0_outputs(9969)) and not (layer0_outputs(3816));
    outputs(8533) <= (layer0_outputs(271)) and not (layer0_outputs(11080));
    outputs(8534) <= (layer0_outputs(12331)) xor (layer0_outputs(6725));
    outputs(8535) <= layer0_outputs(4870);
    outputs(8536) <= (layer0_outputs(9284)) or (layer0_outputs(6515));
    outputs(8537) <= (layer0_outputs(219)) xor (layer0_outputs(4733));
    outputs(8538) <= not(layer0_outputs(2590));
    outputs(8539) <= not(layer0_outputs(5671));
    outputs(8540) <= layer0_outputs(6285);
    outputs(8541) <= not(layer0_outputs(8000));
    outputs(8542) <= layer0_outputs(8686);
    outputs(8543) <= not((layer0_outputs(542)) or (layer0_outputs(819)));
    outputs(8544) <= (layer0_outputs(9351)) xor (layer0_outputs(12335));
    outputs(8545) <= layer0_outputs(10694);
    outputs(8546) <= (layer0_outputs(1361)) and (layer0_outputs(2924));
    outputs(8547) <= not(layer0_outputs(3436)) or (layer0_outputs(11910));
    outputs(8548) <= not((layer0_outputs(8317)) xor (layer0_outputs(2901)));
    outputs(8549) <= layer0_outputs(6100);
    outputs(8550) <= not(layer0_outputs(8004));
    outputs(8551) <= not((layer0_outputs(6600)) xor (layer0_outputs(4568)));
    outputs(8552) <= (layer0_outputs(8220)) xor (layer0_outputs(8835));
    outputs(8553) <= (layer0_outputs(12073)) xor (layer0_outputs(10592));
    outputs(8554) <= not(layer0_outputs(12737)) or (layer0_outputs(9691));
    outputs(8555) <= not(layer0_outputs(6856)) or (layer0_outputs(10994));
    outputs(8556) <= not((layer0_outputs(10089)) xor (layer0_outputs(597)));
    outputs(8557) <= (layer0_outputs(12770)) and not (layer0_outputs(10055));
    outputs(8558) <= (layer0_outputs(3060)) xor (layer0_outputs(1439));
    outputs(8559) <= not(layer0_outputs(5908));
    outputs(8560) <= not((layer0_outputs(9870)) xor (layer0_outputs(817)));
    outputs(8561) <= not(layer0_outputs(1791));
    outputs(8562) <= not((layer0_outputs(11848)) and (layer0_outputs(5636)));
    outputs(8563) <= not(layer0_outputs(998));
    outputs(8564) <= layer0_outputs(1537);
    outputs(8565) <= (layer0_outputs(12121)) and (layer0_outputs(897));
    outputs(8566) <= not(layer0_outputs(9851));
    outputs(8567) <= not(layer0_outputs(4154));
    outputs(8568) <= (layer0_outputs(8739)) and not (layer0_outputs(6083));
    outputs(8569) <= layer0_outputs(9858);
    outputs(8570) <= (layer0_outputs(3294)) and not (layer0_outputs(9422));
    outputs(8571) <= not(layer0_outputs(11444));
    outputs(8572) <= not(layer0_outputs(1197));
    outputs(8573) <= (layer0_outputs(8236)) xor (layer0_outputs(4082));
    outputs(8574) <= layer0_outputs(11949);
    outputs(8575) <= not(layer0_outputs(5043));
    outputs(8576) <= layer0_outputs(10936);
    outputs(8577) <= layer0_outputs(177);
    outputs(8578) <= not(layer0_outputs(2482));
    outputs(8579) <= not(layer0_outputs(4235));
    outputs(8580) <= layer0_outputs(8590);
    outputs(8581) <= layer0_outputs(5106);
    outputs(8582) <= not((layer0_outputs(6436)) or (layer0_outputs(1527)));
    outputs(8583) <= not(layer0_outputs(2305));
    outputs(8584) <= not(layer0_outputs(1401)) or (layer0_outputs(423));
    outputs(8585) <= not((layer0_outputs(10031)) xor (layer0_outputs(11558)));
    outputs(8586) <= not((layer0_outputs(9460)) or (layer0_outputs(4254)));
    outputs(8587) <= not((layer0_outputs(12269)) xor (layer0_outputs(10379)));
    outputs(8588) <= layer0_outputs(4709);
    outputs(8589) <= layer0_outputs(4271);
    outputs(8590) <= not(layer0_outputs(138));
    outputs(8591) <= (layer0_outputs(3986)) and (layer0_outputs(4994));
    outputs(8592) <= (layer0_outputs(11388)) and (layer0_outputs(6239));
    outputs(8593) <= not(layer0_outputs(4239));
    outputs(8594) <= not((layer0_outputs(5855)) xor (layer0_outputs(9779)));
    outputs(8595) <= (layer0_outputs(9961)) and not (layer0_outputs(12442));
    outputs(8596) <= layer0_outputs(10825);
    outputs(8597) <= not((layer0_outputs(1895)) or (layer0_outputs(8298)));
    outputs(8598) <= (layer0_outputs(1006)) and not (layer0_outputs(1347));
    outputs(8599) <= (layer0_outputs(11027)) xor (layer0_outputs(2000));
    outputs(8600) <= not((layer0_outputs(1099)) xor (layer0_outputs(10859)));
    outputs(8601) <= not((layer0_outputs(11555)) xor (layer0_outputs(6)));
    outputs(8602) <= layer0_outputs(9672);
    outputs(8603) <= (layer0_outputs(8980)) xor (layer0_outputs(4035));
    outputs(8604) <= not((layer0_outputs(775)) xor (layer0_outputs(12314)));
    outputs(8605) <= not(layer0_outputs(3358)) or (layer0_outputs(3407));
    outputs(8606) <= not((layer0_outputs(1416)) or (layer0_outputs(7253)));
    outputs(8607) <= not(layer0_outputs(12747));
    outputs(8608) <= layer0_outputs(11591);
    outputs(8609) <= (layer0_outputs(11931)) xor (layer0_outputs(3545));
    outputs(8610) <= layer0_outputs(8543);
    outputs(8611) <= (layer0_outputs(12284)) and not (layer0_outputs(8745));
    outputs(8612) <= layer0_outputs(11202);
    outputs(8613) <= not(layer0_outputs(11253)) or (layer0_outputs(12459));
    outputs(8614) <= layer0_outputs(12704);
    outputs(8615) <= not((layer0_outputs(9959)) and (layer0_outputs(11389)));
    outputs(8616) <= (layer0_outputs(8613)) or (layer0_outputs(12525));
    outputs(8617) <= layer0_outputs(4105);
    outputs(8618) <= not(layer0_outputs(11323));
    outputs(8619) <= layer0_outputs(717);
    outputs(8620) <= not((layer0_outputs(6841)) xor (layer0_outputs(6065)));
    outputs(8621) <= not((layer0_outputs(6358)) xor (layer0_outputs(3623)));
    outputs(8622) <= not(layer0_outputs(205));
    outputs(8623) <= not(layer0_outputs(9113));
    outputs(8624) <= not(layer0_outputs(1555));
    outputs(8625) <= not((layer0_outputs(11526)) or (layer0_outputs(9830)));
    outputs(8626) <= layer0_outputs(8568);
    outputs(8627) <= (layer0_outputs(4709)) and (layer0_outputs(9483));
    outputs(8628) <= not((layer0_outputs(11305)) xor (layer0_outputs(6756)));
    outputs(8629) <= layer0_outputs(6366);
    outputs(8630) <= (layer0_outputs(6698)) xor (layer0_outputs(9501));
    outputs(8631) <= not((layer0_outputs(11962)) xor (layer0_outputs(4113)));
    outputs(8632) <= (layer0_outputs(633)) and not (layer0_outputs(10582));
    outputs(8633) <= (layer0_outputs(9358)) and not (layer0_outputs(8573));
    outputs(8634) <= layer0_outputs(733);
    outputs(8635) <= (layer0_outputs(6851)) and (layer0_outputs(2818));
    outputs(8636) <= (layer0_outputs(12021)) xor (layer0_outputs(6517));
    outputs(8637) <= not(layer0_outputs(4137));
    outputs(8638) <= not(layer0_outputs(8644));
    outputs(8639) <= not(layer0_outputs(1532));
    outputs(8640) <= layer0_outputs(5711);
    outputs(8641) <= (layer0_outputs(12133)) and (layer0_outputs(10672));
    outputs(8642) <= (layer0_outputs(3288)) xor (layer0_outputs(1573));
    outputs(8643) <= layer0_outputs(8175);
    outputs(8644) <= (layer0_outputs(7678)) and not (layer0_outputs(6420));
    outputs(8645) <= layer0_outputs(4914);
    outputs(8646) <= not(layer0_outputs(4498));
    outputs(8647) <= (layer0_outputs(7036)) and not (layer0_outputs(8834));
    outputs(8648) <= layer0_outputs(1844);
    outputs(8649) <= not((layer0_outputs(7928)) xor (layer0_outputs(7216)));
    outputs(8650) <= not(layer0_outputs(1282));
    outputs(8651) <= not(layer0_outputs(5641));
    outputs(8652) <= not((layer0_outputs(1378)) or (layer0_outputs(11561)));
    outputs(8653) <= not(layer0_outputs(3056));
    outputs(8654) <= not((layer0_outputs(2635)) xor (layer0_outputs(1351)));
    outputs(8655) <= not((layer0_outputs(11414)) xor (layer0_outputs(4687)));
    outputs(8656) <= (layer0_outputs(8086)) and not (layer0_outputs(12429));
    outputs(8657) <= layer0_outputs(10601);
    outputs(8658) <= not(layer0_outputs(4647)) or (layer0_outputs(1937));
    outputs(8659) <= (layer0_outputs(1538)) xor (layer0_outputs(6556));
    outputs(8660) <= layer0_outputs(11818);
    outputs(8661) <= (layer0_outputs(4224)) and (layer0_outputs(121));
    outputs(8662) <= layer0_outputs(11051);
    outputs(8663) <= (layer0_outputs(174)) and (layer0_outputs(2722));
    outputs(8664) <= not(layer0_outputs(11362));
    outputs(8665) <= not(layer0_outputs(3496));
    outputs(8666) <= layer0_outputs(11084);
    outputs(8667) <= not((layer0_outputs(635)) or (layer0_outputs(2531)));
    outputs(8668) <= not(layer0_outputs(3853));
    outputs(8669) <= (layer0_outputs(6442)) xor (layer0_outputs(2668));
    outputs(8670) <= not(layer0_outputs(229));
    outputs(8671) <= not(layer0_outputs(9045));
    outputs(8672) <= layer0_outputs(2182);
    outputs(8673) <= layer0_outputs(6166);
    outputs(8674) <= layer0_outputs(11844);
    outputs(8675) <= not(layer0_outputs(10795)) or (layer0_outputs(9079));
    outputs(8676) <= not((layer0_outputs(9553)) and (layer0_outputs(8718)));
    outputs(8677) <= (layer0_outputs(598)) xor (layer0_outputs(4279));
    outputs(8678) <= (layer0_outputs(7412)) xor (layer0_outputs(6928));
    outputs(8679) <= not(layer0_outputs(9153)) or (layer0_outputs(3820));
    outputs(8680) <= not(layer0_outputs(5512));
    outputs(8681) <= layer0_outputs(837);
    outputs(8682) <= not(layer0_outputs(4070));
    outputs(8683) <= not(layer0_outputs(11156));
    outputs(8684) <= not(layer0_outputs(8125)) or (layer0_outputs(7404));
    outputs(8685) <= not(layer0_outputs(6662));
    outputs(8686) <= (layer0_outputs(10608)) xor (layer0_outputs(2477));
    outputs(8687) <= (layer0_outputs(939)) and not (layer0_outputs(10462));
    outputs(8688) <= not((layer0_outputs(4389)) xor (layer0_outputs(12714)));
    outputs(8689) <= not(layer0_outputs(10841));
    outputs(8690) <= not(layer0_outputs(9291)) or (layer0_outputs(2609));
    outputs(8691) <= layer0_outputs(1964);
    outputs(8692) <= layer0_outputs(5067);
    outputs(8693) <= layer0_outputs(8192);
    outputs(8694) <= not(layer0_outputs(2411));
    outputs(8695) <= layer0_outputs(8314);
    outputs(8696) <= (layer0_outputs(1838)) or (layer0_outputs(345));
    outputs(8697) <= not((layer0_outputs(12172)) or (layer0_outputs(352)));
    outputs(8698) <= not(layer0_outputs(1226)) or (layer0_outputs(9916));
    outputs(8699) <= layer0_outputs(2490);
    outputs(8700) <= (layer0_outputs(7732)) or (layer0_outputs(7244));
    outputs(8701) <= not((layer0_outputs(1669)) or (layer0_outputs(10396)));
    outputs(8702) <= (layer0_outputs(1435)) and not (layer0_outputs(4522));
    outputs(8703) <= not(layer0_outputs(1628));
    outputs(8704) <= layer0_outputs(4829);
    outputs(8705) <= not(layer0_outputs(11389));
    outputs(8706) <= (layer0_outputs(3260)) and (layer0_outputs(1856));
    outputs(8707) <= not(layer0_outputs(8833));
    outputs(8708) <= not(layer0_outputs(1111));
    outputs(8709) <= layer0_outputs(7405);
    outputs(8710) <= layer0_outputs(10266);
    outputs(8711) <= not((layer0_outputs(7818)) or (layer0_outputs(9212)));
    outputs(8712) <= layer0_outputs(8798);
    outputs(8713) <= not(layer0_outputs(12043)) or (layer0_outputs(4283));
    outputs(8714) <= not(layer0_outputs(8897)) or (layer0_outputs(232));
    outputs(8715) <= (layer0_outputs(5967)) xor (layer0_outputs(9089));
    outputs(8716) <= not(layer0_outputs(10770));
    outputs(8717) <= not(layer0_outputs(4633)) or (layer0_outputs(1380));
    outputs(8718) <= (layer0_outputs(1335)) or (layer0_outputs(7725));
    outputs(8719) <= (layer0_outputs(5111)) xor (layer0_outputs(12479));
    outputs(8720) <= layer0_outputs(4131);
    outputs(8721) <= not(layer0_outputs(25));
    outputs(8722) <= not(layer0_outputs(1828));
    outputs(8723) <= layer0_outputs(1622);
    outputs(8724) <= not((layer0_outputs(7268)) or (layer0_outputs(11786)));
    outputs(8725) <= not(layer0_outputs(11581));
    outputs(8726) <= (layer0_outputs(4598)) and not (layer0_outputs(4922));
    outputs(8727) <= not((layer0_outputs(4263)) xor (layer0_outputs(7424)));
    outputs(8728) <= layer0_outputs(11945);
    outputs(8729) <= (layer0_outputs(326)) and not (layer0_outputs(3058));
    outputs(8730) <= not(layer0_outputs(8984));
    outputs(8731) <= (layer0_outputs(8881)) xor (layer0_outputs(2596));
    outputs(8732) <= not((layer0_outputs(1416)) xor (layer0_outputs(1227)));
    outputs(8733) <= layer0_outputs(6127);
    outputs(8734) <= not(layer0_outputs(6846));
    outputs(8735) <= not(layer0_outputs(10149)) or (layer0_outputs(2063));
    outputs(8736) <= (layer0_outputs(11985)) and not (layer0_outputs(4578));
    outputs(8737) <= not(layer0_outputs(3359)) or (layer0_outputs(11110));
    outputs(8738) <= (layer0_outputs(2391)) xor (layer0_outputs(7608));
    outputs(8739) <= not(layer0_outputs(404));
    outputs(8740) <= layer0_outputs(4229);
    outputs(8741) <= not((layer0_outputs(7248)) xor (layer0_outputs(6198)));
    outputs(8742) <= not((layer0_outputs(7795)) xor (layer0_outputs(7385)));
    outputs(8743) <= (layer0_outputs(4400)) xor (layer0_outputs(2759));
    outputs(8744) <= not(layer0_outputs(263)) or (layer0_outputs(7257));
    outputs(8745) <= not(layer0_outputs(485)) or (layer0_outputs(8289));
    outputs(8746) <= layer0_outputs(7422);
    outputs(8747) <= layer0_outputs(11766);
    outputs(8748) <= layer0_outputs(6327);
    outputs(8749) <= layer0_outputs(2662);
    outputs(8750) <= layer0_outputs(12262);
    outputs(8751) <= (layer0_outputs(10659)) and not (layer0_outputs(4241));
    outputs(8752) <= not((layer0_outputs(10724)) xor (layer0_outputs(12065)));
    outputs(8753) <= layer0_outputs(1285);
    outputs(8754) <= (layer0_outputs(9132)) and (layer0_outputs(10595));
    outputs(8755) <= (layer0_outputs(6275)) or (layer0_outputs(9696));
    outputs(8756) <= (layer0_outputs(8034)) xor (layer0_outputs(3330));
    outputs(8757) <= not(layer0_outputs(11639));
    outputs(8758) <= (layer0_outputs(10140)) xor (layer0_outputs(9610));
    outputs(8759) <= layer0_outputs(5382);
    outputs(8760) <= (layer0_outputs(9875)) and not (layer0_outputs(12559));
    outputs(8761) <= not(layer0_outputs(7709));
    outputs(8762) <= not(layer0_outputs(8636));
    outputs(8763) <= not((layer0_outputs(8284)) or (layer0_outputs(7522)));
    outputs(8764) <= (layer0_outputs(985)) and not (layer0_outputs(577));
    outputs(8765) <= not((layer0_outputs(7655)) xor (layer0_outputs(8383)));
    outputs(8766) <= not(layer0_outputs(10854));
    outputs(8767) <= layer0_outputs(7586);
    outputs(8768) <= layer0_outputs(2155);
    outputs(8769) <= layer0_outputs(11094);
    outputs(8770) <= not((layer0_outputs(2321)) and (layer0_outputs(5355)));
    outputs(8771) <= layer0_outputs(10017);
    outputs(8772) <= not(layer0_outputs(10102)) or (layer0_outputs(6518));
    outputs(8773) <= not((layer0_outputs(12285)) xor (layer0_outputs(4792)));
    outputs(8774) <= not((layer0_outputs(2245)) xor (layer0_outputs(4551)));
    outputs(8775) <= not(layer0_outputs(11373));
    outputs(8776) <= layer0_outputs(1384);
    outputs(8777) <= not(layer0_outputs(4855));
    outputs(8778) <= layer0_outputs(10927);
    outputs(8779) <= not(layer0_outputs(8617));
    outputs(8780) <= layer0_outputs(11984);
    outputs(8781) <= not(layer0_outputs(2088));
    outputs(8782) <= layer0_outputs(469);
    outputs(8783) <= (layer0_outputs(7260)) xor (layer0_outputs(2717));
    outputs(8784) <= (layer0_outputs(9784)) and (layer0_outputs(797));
    outputs(8785) <= not((layer0_outputs(5417)) or (layer0_outputs(9328)));
    outputs(8786) <= layer0_outputs(3631);
    outputs(8787) <= not(layer0_outputs(321));
    outputs(8788) <= not(layer0_outputs(12310)) or (layer0_outputs(1009));
    outputs(8789) <= layer0_outputs(11105);
    outputs(8790) <= not((layer0_outputs(10231)) or (layer0_outputs(10096)));
    outputs(8791) <= not((layer0_outputs(7297)) and (layer0_outputs(6493)));
    outputs(8792) <= not(layer0_outputs(6183));
    outputs(8793) <= layer0_outputs(11192);
    outputs(8794) <= not(layer0_outputs(4513));
    outputs(8795) <= (layer0_outputs(10437)) xor (layer0_outputs(1527));
    outputs(8796) <= not(layer0_outputs(11462));
    outputs(8797) <= not((layer0_outputs(9907)) or (layer0_outputs(8556)));
    outputs(8798) <= layer0_outputs(7376);
    outputs(8799) <= not((layer0_outputs(5333)) or (layer0_outputs(6741)));
    outputs(8800) <= (layer0_outputs(10796)) and not (layer0_outputs(7418));
    outputs(8801) <= not(layer0_outputs(176));
    outputs(8802) <= (layer0_outputs(8570)) xor (layer0_outputs(8620));
    outputs(8803) <= not(layer0_outputs(4524)) or (layer0_outputs(3549));
    outputs(8804) <= layer0_outputs(12040);
    outputs(8805) <= not((layer0_outputs(12025)) xor (layer0_outputs(8252)));
    outputs(8806) <= not(layer0_outputs(8333)) or (layer0_outputs(5892));
    outputs(8807) <= (layer0_outputs(10927)) and not (layer0_outputs(7441));
    outputs(8808) <= layer0_outputs(3915);
    outputs(8809) <= layer0_outputs(9888);
    outputs(8810) <= layer0_outputs(5536);
    outputs(8811) <= (layer0_outputs(7700)) and (layer0_outputs(8241));
    outputs(8812) <= layer0_outputs(10467);
    outputs(8813) <= not((layer0_outputs(6929)) xor (layer0_outputs(4394)));
    outputs(8814) <= layer0_outputs(5088);
    outputs(8815) <= (layer0_outputs(7804)) xor (layer0_outputs(401));
    outputs(8816) <= layer0_outputs(9021);
    outputs(8817) <= not((layer0_outputs(4624)) or (layer0_outputs(2962)));
    outputs(8818) <= not((layer0_outputs(3413)) xor (layer0_outputs(12709)));
    outputs(8819) <= layer0_outputs(2103);
    outputs(8820) <= not((layer0_outputs(10745)) xor (layer0_outputs(9847)));
    outputs(8821) <= not((layer0_outputs(8577)) xor (layer0_outputs(2559)));
    outputs(8822) <= not((layer0_outputs(10557)) and (layer0_outputs(8050)));
    outputs(8823) <= (layer0_outputs(9135)) and not (layer0_outputs(11897));
    outputs(8824) <= not((layer0_outputs(5543)) and (layer0_outputs(7473)));
    outputs(8825) <= (layer0_outputs(1079)) xor (layer0_outputs(11314));
    outputs(8826) <= not(layer0_outputs(10160));
    outputs(8827) <= layer0_outputs(8126);
    outputs(8828) <= (layer0_outputs(4837)) xor (layer0_outputs(7478));
    outputs(8829) <= (layer0_outputs(9128)) and not (layer0_outputs(11718));
    outputs(8830) <= layer0_outputs(11271);
    outputs(8831) <= not(layer0_outputs(2623));
    outputs(8832) <= (layer0_outputs(7735)) and (layer0_outputs(7584));
    outputs(8833) <= layer0_outputs(271);
    outputs(8834) <= not(layer0_outputs(7551));
    outputs(8835) <= not((layer0_outputs(12793)) xor (layer0_outputs(4377)));
    outputs(8836) <= layer0_outputs(6933);
    outputs(8837) <= (layer0_outputs(7560)) xor (layer0_outputs(4228));
    outputs(8838) <= not(layer0_outputs(4329));
    outputs(8839) <= layer0_outputs(7068);
    outputs(8840) <= (layer0_outputs(5213)) and not (layer0_outputs(8088));
    outputs(8841) <= layer0_outputs(3984);
    outputs(8842) <= layer0_outputs(4346);
    outputs(8843) <= not(layer0_outputs(7155));
    outputs(8844) <= not((layer0_outputs(2672)) and (layer0_outputs(9008)));
    outputs(8845) <= not(layer0_outputs(4937)) or (layer0_outputs(3361));
    outputs(8846) <= not(layer0_outputs(4794)) or (layer0_outputs(2375));
    outputs(8847) <= (layer0_outputs(6751)) or (layer0_outputs(1132));
    outputs(8848) <= not(layer0_outputs(1165));
    outputs(8849) <= not(layer0_outputs(8010));
    outputs(8850) <= not(layer0_outputs(7414));
    outputs(8851) <= layer0_outputs(6401);
    outputs(8852) <= layer0_outputs(1236);
    outputs(8853) <= (layer0_outputs(11482)) or (layer0_outputs(11636));
    outputs(8854) <= (layer0_outputs(493)) xor (layer0_outputs(1671));
    outputs(8855) <= layer0_outputs(9630);
    outputs(8856) <= (layer0_outputs(3190)) and not (layer0_outputs(9511));
    outputs(8857) <= layer0_outputs(1150);
    outputs(8858) <= (layer0_outputs(12191)) and not (layer0_outputs(5357));
    outputs(8859) <= (layer0_outputs(10944)) xor (layer0_outputs(228));
    outputs(8860) <= (layer0_outputs(6269)) or (layer0_outputs(1870));
    outputs(8861) <= not(layer0_outputs(11887));
    outputs(8862) <= not(layer0_outputs(12500));
    outputs(8863) <= not(layer0_outputs(3168));
    outputs(8864) <= not(layer0_outputs(5610));
    outputs(8865) <= not(layer0_outputs(1477));
    outputs(8866) <= layer0_outputs(10494);
    outputs(8867) <= (layer0_outputs(3594)) and (layer0_outputs(8945));
    outputs(8868) <= layer0_outputs(4105);
    outputs(8869) <= not(layer0_outputs(5956));
    outputs(8870) <= (layer0_outputs(6482)) xor (layer0_outputs(5331));
    outputs(8871) <= layer0_outputs(1209);
    outputs(8872) <= not(layer0_outputs(3937));
    outputs(8873) <= layer0_outputs(543);
    outputs(8874) <= not((layer0_outputs(1999)) or (layer0_outputs(1083)));
    outputs(8875) <= (layer0_outputs(12184)) xor (layer0_outputs(3000));
    outputs(8876) <= (layer0_outputs(10369)) xor (layer0_outputs(3272));
    outputs(8877) <= not((layer0_outputs(6993)) xor (layer0_outputs(5635)));
    outputs(8878) <= not(layer0_outputs(11653));
    outputs(8879) <= not(layer0_outputs(3334));
    outputs(8880) <= not(layer0_outputs(4386)) or (layer0_outputs(10491));
    outputs(8881) <= layer0_outputs(791);
    outputs(8882) <= not(layer0_outputs(7722));
    outputs(8883) <= not(layer0_outputs(11476));
    outputs(8884) <= layer0_outputs(5038);
    outputs(8885) <= not(layer0_outputs(11295));
    outputs(8886) <= (layer0_outputs(1815)) xor (layer0_outputs(9510));
    outputs(8887) <= not((layer0_outputs(102)) or (layer0_outputs(6061)));
    outputs(8888) <= not(layer0_outputs(3660));
    outputs(8889) <= (layer0_outputs(6827)) xor (layer0_outputs(5244));
    outputs(8890) <= not(layer0_outputs(9615));
    outputs(8891) <= not(layer0_outputs(8981));
    outputs(8892) <= layer0_outputs(7904);
    outputs(8893) <= not((layer0_outputs(3505)) or (layer0_outputs(7890)));
    outputs(8894) <= (layer0_outputs(8619)) and not (layer0_outputs(7165));
    outputs(8895) <= not((layer0_outputs(10524)) xor (layer0_outputs(6052)));
    outputs(8896) <= not(layer0_outputs(3924));
    outputs(8897) <= layer0_outputs(11824);
    outputs(8898) <= not((layer0_outputs(10611)) xor (layer0_outputs(3995)));
    outputs(8899) <= not((layer0_outputs(10133)) xor (layer0_outputs(3154)));
    outputs(8900) <= not(layer0_outputs(586)) or (layer0_outputs(9691));
    outputs(8901) <= (layer0_outputs(4333)) or (layer0_outputs(10382));
    outputs(8902) <= (layer0_outputs(6922)) and not (layer0_outputs(10060));
    outputs(8903) <= not(layer0_outputs(9647));
    outputs(8904) <= (layer0_outputs(6159)) or (layer0_outputs(12209));
    outputs(8905) <= not(layer0_outputs(2589));
    outputs(8906) <= not(layer0_outputs(6123));
    outputs(8907) <= not(layer0_outputs(6147)) or (layer0_outputs(12481));
    outputs(8908) <= layer0_outputs(10128);
    outputs(8909) <= (layer0_outputs(3437)) and not (layer0_outputs(11490));
    outputs(8910) <= not((layer0_outputs(5952)) xor (layer0_outputs(12734)));
    outputs(8911) <= not(layer0_outputs(11161));
    outputs(8912) <= layer0_outputs(10525);
    outputs(8913) <= (layer0_outputs(5243)) and not (layer0_outputs(10579));
    outputs(8914) <= (layer0_outputs(11278)) and (layer0_outputs(4504));
    outputs(8915) <= (layer0_outputs(10834)) xor (layer0_outputs(7859));
    outputs(8916) <= layer0_outputs(3405);
    outputs(8917) <= not((layer0_outputs(4356)) or (layer0_outputs(10119)));
    outputs(8918) <= layer0_outputs(304);
    outputs(8919) <= (layer0_outputs(7489)) and (layer0_outputs(12450));
    outputs(8920) <= layer0_outputs(569);
    outputs(8921) <= (layer0_outputs(1802)) and (layer0_outputs(4752));
    outputs(8922) <= not((layer0_outputs(7645)) or (layer0_outputs(1363)));
    outputs(8923) <= layer0_outputs(10464);
    outputs(8924) <= not((layer0_outputs(7635)) or (layer0_outputs(10634)));
    outputs(8925) <= not(layer0_outputs(3311));
    outputs(8926) <= not(layer0_outputs(3357));
    outputs(8927) <= layer0_outputs(2512);
    outputs(8928) <= (layer0_outputs(8794)) xor (layer0_outputs(6614));
    outputs(8929) <= not(layer0_outputs(8394));
    outputs(8930) <= not(layer0_outputs(4881));
    outputs(8931) <= layer0_outputs(8183);
    outputs(8932) <= not(layer0_outputs(299));
    outputs(8933) <= not((layer0_outputs(11490)) or (layer0_outputs(2440)));
    outputs(8934) <= (layer0_outputs(5992)) xor (layer0_outputs(8465));
    outputs(8935) <= not(layer0_outputs(5616));
    outputs(8936) <= (layer0_outputs(10449)) and not (layer0_outputs(6036));
    outputs(8937) <= not(layer0_outputs(8132));
    outputs(8938) <= layer0_outputs(5706);
    outputs(8939) <= not((layer0_outputs(7344)) xor (layer0_outputs(1313)));
    outputs(8940) <= (layer0_outputs(5181)) and not (layer0_outputs(8021));
    outputs(8941) <= layer0_outputs(1810);
    outputs(8942) <= not((layer0_outputs(8077)) xor (layer0_outputs(2426)));
    outputs(8943) <= not((layer0_outputs(3659)) xor (layer0_outputs(693)));
    outputs(8944) <= not((layer0_outputs(10669)) xor (layer0_outputs(937)));
    outputs(8945) <= layer0_outputs(6877);
    outputs(8946) <= not((layer0_outputs(4793)) xor (layer0_outputs(8600)));
    outputs(8947) <= (layer0_outputs(4136)) and not (layer0_outputs(11328));
    outputs(8948) <= not((layer0_outputs(5837)) or (layer0_outputs(4022)));
    outputs(8949) <= layer0_outputs(4219);
    outputs(8950) <= layer0_outputs(5363);
    outputs(8951) <= (layer0_outputs(4049)) or (layer0_outputs(3007));
    outputs(8952) <= not(layer0_outputs(1292)) or (layer0_outputs(11170));
    outputs(8953) <= not((layer0_outputs(1134)) xor (layer0_outputs(7867)));
    outputs(8954) <= (layer0_outputs(1700)) and not (layer0_outputs(9009));
    outputs(8955) <= not(layer0_outputs(595));
    outputs(8956) <= not(layer0_outputs(952));
    outputs(8957) <= layer0_outputs(11188);
    outputs(8958) <= layer0_outputs(7330);
    outputs(8959) <= (layer0_outputs(7725)) xor (layer0_outputs(2066));
    outputs(8960) <= (layer0_outputs(4682)) and (layer0_outputs(12406));
    outputs(8961) <= layer0_outputs(2957);
    outputs(8962) <= not(layer0_outputs(10084)) or (layer0_outputs(12486));
    outputs(8963) <= (layer0_outputs(10011)) and not (layer0_outputs(7632));
    outputs(8964) <= not(layer0_outputs(3930)) or (layer0_outputs(750));
    outputs(8965) <= layer0_outputs(2472);
    outputs(8966) <= not(layer0_outputs(2944));
    outputs(8967) <= not(layer0_outputs(11586));
    outputs(8968) <= (layer0_outputs(3621)) and not (layer0_outputs(771));
    outputs(8969) <= not(layer0_outputs(7884)) or (layer0_outputs(2153));
    outputs(8970) <= not(layer0_outputs(4169));
    outputs(8971) <= not((layer0_outputs(6315)) and (layer0_outputs(6900)));
    outputs(8972) <= not(layer0_outputs(6172));
    outputs(8973) <= not(layer0_outputs(2494));
    outputs(8974) <= layer0_outputs(3203);
    outputs(8975) <= layer0_outputs(3303);
    outputs(8976) <= (layer0_outputs(12488)) and not (layer0_outputs(306));
    outputs(8977) <= layer0_outputs(420);
    outputs(8978) <= not(layer0_outputs(3180));
    outputs(8979) <= (layer0_outputs(3315)) or (layer0_outputs(11689));
    outputs(8980) <= (layer0_outputs(3146)) and not (layer0_outputs(3521));
    outputs(8981) <= not(layer0_outputs(3659));
    outputs(8982) <= layer0_outputs(4836);
    outputs(8983) <= not((layer0_outputs(12742)) or (layer0_outputs(10134)));
    outputs(8984) <= not((layer0_outputs(11817)) or (layer0_outputs(5875)));
    outputs(8985) <= layer0_outputs(4348);
    outputs(8986) <= not(layer0_outputs(11993)) or (layer0_outputs(11752));
    outputs(8987) <= not(layer0_outputs(4904));
    outputs(8988) <= (layer0_outputs(12505)) and not (layer0_outputs(8555));
    outputs(8989) <= layer0_outputs(2261);
    outputs(8990) <= (layer0_outputs(7532)) xor (layer0_outputs(11377));
    outputs(8991) <= not((layer0_outputs(7497)) xor (layer0_outputs(3898)));
    outputs(8992) <= layer0_outputs(1664);
    outputs(8993) <= (layer0_outputs(716)) xor (layer0_outputs(6621));
    outputs(8994) <= not((layer0_outputs(7923)) xor (layer0_outputs(5351)));
    outputs(8995) <= (layer0_outputs(8693)) xor (layer0_outputs(7599));
    outputs(8996) <= layer0_outputs(7527);
    outputs(8997) <= layer0_outputs(6178);
    outputs(8998) <= not(layer0_outputs(603));
    outputs(8999) <= not((layer0_outputs(7190)) or (layer0_outputs(8574)));
    outputs(9000) <= not(layer0_outputs(10526)) or (layer0_outputs(9907));
    outputs(9001) <= not((layer0_outputs(4602)) or (layer0_outputs(10408)));
    outputs(9002) <= (layer0_outputs(3371)) and not (layer0_outputs(8904));
    outputs(9003) <= not(layer0_outputs(1179)) or (layer0_outputs(7995));
    outputs(9004) <= not(layer0_outputs(1231)) or (layer0_outputs(3249));
    outputs(9005) <= layer0_outputs(3763);
    outputs(9006) <= layer0_outputs(9673);
    outputs(9007) <= not((layer0_outputs(6091)) xor (layer0_outputs(7061)));
    outputs(9008) <= (layer0_outputs(4404)) and not (layer0_outputs(2335));
    outputs(9009) <= (layer0_outputs(4901)) xor (layer0_outputs(5225));
    outputs(9010) <= layer0_outputs(6298);
    outputs(9011) <= not(layer0_outputs(7503));
    outputs(9012) <= layer0_outputs(1491);
    outputs(9013) <= not((layer0_outputs(9057)) xor (layer0_outputs(6915)));
    outputs(9014) <= not((layer0_outputs(12465)) xor (layer0_outputs(5778)));
    outputs(9015) <= (layer0_outputs(11918)) and not (layer0_outputs(7925));
    outputs(9016) <= (layer0_outputs(7627)) and not (layer0_outputs(7663));
    outputs(9017) <= layer0_outputs(8905);
    outputs(9018) <= not((layer0_outputs(4319)) and (layer0_outputs(1225)));
    outputs(9019) <= (layer0_outputs(3684)) and not (layer0_outputs(4252));
    outputs(9020) <= layer0_outputs(3963);
    outputs(9021) <= not(layer0_outputs(3316));
    outputs(9022) <= (layer0_outputs(3444)) xor (layer0_outputs(9506));
    outputs(9023) <= layer0_outputs(8550);
    outputs(9024) <= layer0_outputs(7235);
    outputs(9025) <= (layer0_outputs(6982)) xor (layer0_outputs(7775));
    outputs(9026) <= (layer0_outputs(6694)) xor (layer0_outputs(1714));
    outputs(9027) <= layer0_outputs(2815);
    outputs(9028) <= (layer0_outputs(1952)) and not (layer0_outputs(5581));
    outputs(9029) <= layer0_outputs(2675);
    outputs(9030) <= layer0_outputs(4011);
    outputs(9031) <= layer0_outputs(11231);
    outputs(9032) <= not(layer0_outputs(1062));
    outputs(9033) <= not((layer0_outputs(12110)) xor (layer0_outputs(8261)));
    outputs(9034) <= not(layer0_outputs(2142));
    outputs(9035) <= not((layer0_outputs(3375)) xor (layer0_outputs(7792)));
    outputs(9036) <= not((layer0_outputs(474)) xor (layer0_outputs(11219)));
    outputs(9037) <= (layer0_outputs(5434)) xor (layer0_outputs(8846));
    outputs(9038) <= layer0_outputs(11999);
    outputs(9039) <= (layer0_outputs(4651)) xor (layer0_outputs(12047));
    outputs(9040) <= not(layer0_outputs(7397)) or (layer0_outputs(2132));
    outputs(9041) <= not(layer0_outputs(5773));
    outputs(9042) <= not(layer0_outputs(10677));
    outputs(9043) <= layer0_outputs(6896);
    outputs(9044) <= layer0_outputs(8688);
    outputs(9045) <= (layer0_outputs(6783)) and (layer0_outputs(12332));
    outputs(9046) <= not(layer0_outputs(4679));
    outputs(9047) <= not(layer0_outputs(6841));
    outputs(9048) <= (layer0_outputs(8663)) xor (layer0_outputs(9736));
    outputs(9049) <= not(layer0_outputs(7228));
    outputs(9050) <= not(layer0_outputs(3031));
    outputs(9051) <= layer0_outputs(12383);
    outputs(9052) <= not((layer0_outputs(10304)) and (layer0_outputs(2326)));
    outputs(9053) <= not(layer0_outputs(10232));
    outputs(9054) <= layer0_outputs(12149);
    outputs(9055) <= (layer0_outputs(1763)) xor (layer0_outputs(6806));
    outputs(9056) <= (layer0_outputs(3191)) xor (layer0_outputs(1960));
    outputs(9057) <= (layer0_outputs(3222)) and (layer0_outputs(10364));
    outputs(9058) <= layer0_outputs(1259);
    outputs(9059) <= not(layer0_outputs(10861)) or (layer0_outputs(10197));
    outputs(9060) <= (layer0_outputs(5413)) or (layer0_outputs(1495));
    outputs(9061) <= layer0_outputs(10068);
    outputs(9062) <= (layer0_outputs(2420)) xor (layer0_outputs(5538));
    outputs(9063) <= layer0_outputs(7138);
    outputs(9064) <= not(layer0_outputs(11032)) or (layer0_outputs(7291));
    outputs(9065) <= layer0_outputs(6955);
    outputs(9066) <= (layer0_outputs(11172)) and not (layer0_outputs(1983));
    outputs(9067) <= (layer0_outputs(9574)) and (layer0_outputs(981));
    outputs(9068) <= layer0_outputs(7329);
    outputs(9069) <= layer0_outputs(5606);
    outputs(9070) <= not(layer0_outputs(6004));
    outputs(9071) <= not((layer0_outputs(1048)) xor (layer0_outputs(5749)));
    outputs(9072) <= layer0_outputs(7929);
    outputs(9073) <= not(layer0_outputs(5534)) or (layer0_outputs(3443));
    outputs(9074) <= not((layer0_outputs(12754)) xor (layer0_outputs(1566)));
    outputs(9075) <= layer0_outputs(11529);
    outputs(9076) <= not((layer0_outputs(3473)) or (layer0_outputs(1472)));
    outputs(9077) <= (layer0_outputs(9132)) xor (layer0_outputs(8149));
    outputs(9078) <= layer0_outputs(3959);
    outputs(9079) <= (layer0_outputs(9289)) and (layer0_outputs(9017));
    outputs(9080) <= (layer0_outputs(231)) and not (layer0_outputs(9365));
    outputs(9081) <= not(layer0_outputs(306));
    outputs(9082) <= (layer0_outputs(5033)) xor (layer0_outputs(10173));
    outputs(9083) <= not(layer0_outputs(791));
    outputs(9084) <= not(layer0_outputs(5514));
    outputs(9085) <= layer0_outputs(5654);
    outputs(9086) <= (layer0_outputs(4211)) xor (layer0_outputs(9773));
    outputs(9087) <= not(layer0_outputs(4148));
    outputs(9088) <= (layer0_outputs(3920)) and not (layer0_outputs(1714));
    outputs(9089) <= not(layer0_outputs(6506));
    outputs(9090) <= (layer0_outputs(5802)) or (layer0_outputs(958));
    outputs(9091) <= (layer0_outputs(5724)) and not (layer0_outputs(6968));
    outputs(9092) <= not(layer0_outputs(5478)) or (layer0_outputs(96));
    outputs(9093) <= not(layer0_outputs(3191));
    outputs(9094) <= layer0_outputs(5408);
    outputs(9095) <= not(layer0_outputs(6537));
    outputs(9096) <= (layer0_outputs(7079)) xor (layer0_outputs(11097));
    outputs(9097) <= not(layer0_outputs(11987));
    outputs(9098) <= not((layer0_outputs(1251)) or (layer0_outputs(1393)));
    outputs(9099) <= not(layer0_outputs(4390));
    outputs(9100) <= not(layer0_outputs(10302));
    outputs(9101) <= (layer0_outputs(10663)) xor (layer0_outputs(11276));
    outputs(9102) <= not(layer0_outputs(449));
    outputs(9103) <= layer0_outputs(12089);
    outputs(9104) <= layer0_outputs(2950);
    outputs(9105) <= layer0_outputs(6383);
    outputs(9106) <= (layer0_outputs(12276)) xor (layer0_outputs(12583));
    outputs(9107) <= (layer0_outputs(2125)) and (layer0_outputs(2427));
    outputs(9108) <= not(layer0_outputs(7541));
    outputs(9109) <= layer0_outputs(4864);
    outputs(9110) <= not(layer0_outputs(10877));
    outputs(9111) <= not(layer0_outputs(2269)) or (layer0_outputs(11216));
    outputs(9112) <= (layer0_outputs(5029)) and (layer0_outputs(1053));
    outputs(9113) <= not(layer0_outputs(668));
    outputs(9114) <= (layer0_outputs(8858)) and not (layer0_outputs(10719));
    outputs(9115) <= (layer0_outputs(5732)) and not (layer0_outputs(11545));
    outputs(9116) <= (layer0_outputs(928)) and (layer0_outputs(6410));
    outputs(9117) <= layer0_outputs(1391);
    outputs(9118) <= not((layer0_outputs(11310)) xor (layer0_outputs(7220)));
    outputs(9119) <= (layer0_outputs(5912)) xor (layer0_outputs(11256));
    outputs(9120) <= (layer0_outputs(7535)) and (layer0_outputs(3872));
    outputs(9121) <= layer0_outputs(2243);
    outputs(9122) <= (layer0_outputs(11877)) and not (layer0_outputs(9715));
    outputs(9123) <= (layer0_outputs(39)) xor (layer0_outputs(5117));
    outputs(9124) <= (layer0_outputs(12117)) and (layer0_outputs(5678));
    outputs(9125) <= not((layer0_outputs(3620)) xor (layer0_outputs(12187)));
    outputs(9126) <= layer0_outputs(9289);
    outputs(9127) <= layer0_outputs(8085);
    outputs(9128) <= (layer0_outputs(7563)) and (layer0_outputs(9730));
    outputs(9129) <= not(layer0_outputs(4317));
    outputs(9130) <= (layer0_outputs(9454)) xor (layer0_outputs(3038));
    outputs(9131) <= layer0_outputs(5748);
    outputs(9132) <= layer0_outputs(9608);
    outputs(9133) <= not(layer0_outputs(741)) or (layer0_outputs(9150));
    outputs(9134) <= layer0_outputs(1125);
    outputs(9135) <= not(layer0_outputs(8793));
    outputs(9136) <= layer0_outputs(6957);
    outputs(9137) <= not(layer0_outputs(11553));
    outputs(9138) <= (layer0_outputs(7943)) xor (layer0_outputs(10129));
    outputs(9139) <= layer0_outputs(1205);
    outputs(9140) <= not(layer0_outputs(512));
    outputs(9141) <= not(layer0_outputs(9043)) or (layer0_outputs(1297));
    outputs(9142) <= not(layer0_outputs(4886));
    outputs(9143) <= (layer0_outputs(10330)) and (layer0_outputs(8141));
    outputs(9144) <= not(layer0_outputs(717));
    outputs(9145) <= layer0_outputs(6605);
    outputs(9146) <= layer0_outputs(5859);
    outputs(9147) <= not((layer0_outputs(8677)) and (layer0_outputs(10185)));
    outputs(9148) <= (layer0_outputs(6678)) and (layer0_outputs(10394));
    outputs(9149) <= not((layer0_outputs(10472)) xor (layer0_outputs(10225)));
    outputs(9150) <= (layer0_outputs(1857)) xor (layer0_outputs(6637));
    outputs(9151) <= (layer0_outputs(3994)) xor (layer0_outputs(1025));
    outputs(9152) <= not(layer0_outputs(9625));
    outputs(9153) <= not((layer0_outputs(10196)) xor (layer0_outputs(4373)));
    outputs(9154) <= not((layer0_outputs(4985)) and (layer0_outputs(3109)));
    outputs(9155) <= not((layer0_outputs(7423)) or (layer0_outputs(6055)));
    outputs(9156) <= not(layer0_outputs(11396));
    outputs(9157) <= not(layer0_outputs(1711)) or (layer0_outputs(6374));
    outputs(9158) <= layer0_outputs(2451);
    outputs(9159) <= not((layer0_outputs(11498)) or (layer0_outputs(8854)));
    outputs(9160) <= layer0_outputs(6705);
    outputs(9161) <= not(layer0_outputs(7024));
    outputs(9162) <= not(layer0_outputs(927));
    outputs(9163) <= (layer0_outputs(12566)) and (layer0_outputs(2785));
    outputs(9164) <= not((layer0_outputs(2505)) xor (layer0_outputs(11836)));
    outputs(9165) <= (layer0_outputs(8512)) xor (layer0_outputs(4232));
    outputs(9166) <= (layer0_outputs(6910)) xor (layer0_outputs(10085));
    outputs(9167) <= not(layer0_outputs(3843));
    outputs(9168) <= layer0_outputs(5119);
    outputs(9169) <= layer0_outputs(2655);
    outputs(9170) <= layer0_outputs(6792);
    outputs(9171) <= layer0_outputs(9202);
    outputs(9172) <= not((layer0_outputs(3981)) xor (layer0_outputs(5588)));
    outputs(9173) <= (layer0_outputs(7493)) xor (layer0_outputs(7437));
    outputs(9174) <= not(layer0_outputs(11310));
    outputs(9175) <= not(layer0_outputs(5909));
    outputs(9176) <= layer0_outputs(1171);
    outputs(9177) <= not(layer0_outputs(10319));
    outputs(9178) <= layer0_outputs(5334);
    outputs(9179) <= not(layer0_outputs(9654));
    outputs(9180) <= (layer0_outputs(11600)) xor (layer0_outputs(1890));
    outputs(9181) <= not((layer0_outputs(1139)) xor (layer0_outputs(5745)));
    outputs(9182) <= layer0_outputs(3366);
    outputs(9183) <= not((layer0_outputs(8597)) xor (layer0_outputs(6262)));
    outputs(9184) <= (layer0_outputs(7118)) and not (layer0_outputs(5093));
    outputs(9185) <= not((layer0_outputs(183)) xor (layer0_outputs(12637)));
    outputs(9186) <= not(layer0_outputs(1807));
    outputs(9187) <= (layer0_outputs(4596)) or (layer0_outputs(3702));
    outputs(9188) <= not((layer0_outputs(12482)) or (layer0_outputs(4919)));
    outputs(9189) <= (layer0_outputs(12062)) and (layer0_outputs(11270));
    outputs(9190) <= (layer0_outputs(3870)) and not (layer0_outputs(1090));
    outputs(9191) <= layer0_outputs(9878);
    outputs(9192) <= not(layer0_outputs(8705)) or (layer0_outputs(6888));
    outputs(9193) <= layer0_outputs(5124);
    outputs(9194) <= layer0_outputs(5699);
    outputs(9195) <= not((layer0_outputs(655)) or (layer0_outputs(2123)));
    outputs(9196) <= not((layer0_outputs(6324)) or (layer0_outputs(3606)));
    outputs(9197) <= layer0_outputs(627);
    outputs(9198) <= not(layer0_outputs(3878)) or (layer0_outputs(2913));
    outputs(9199) <= not(layer0_outputs(8047));
    outputs(9200) <= (layer0_outputs(7775)) and (layer0_outputs(970));
    outputs(9201) <= not(layer0_outputs(7776));
    outputs(9202) <= layer0_outputs(4765);
    outputs(9203) <= not((layer0_outputs(1191)) or (layer0_outputs(8539)));
    outputs(9204) <= not(layer0_outputs(4973));
    outputs(9205) <= (layer0_outputs(6339)) and not (layer0_outputs(9774));
    outputs(9206) <= (layer0_outputs(2650)) and (layer0_outputs(9275));
    outputs(9207) <= (layer0_outputs(8357)) and not (layer0_outputs(10344));
    outputs(9208) <= layer0_outputs(8172);
    outputs(9209) <= layer0_outputs(8476);
    outputs(9210) <= (layer0_outputs(10000)) and (layer0_outputs(11744));
    outputs(9211) <= not((layer0_outputs(1383)) and (layer0_outputs(6408)));
    outputs(9212) <= (layer0_outputs(8336)) xor (layer0_outputs(1834));
    outputs(9213) <= not((layer0_outputs(8604)) xor (layer0_outputs(9187)));
    outputs(9214) <= not((layer0_outputs(9147)) xor (layer0_outputs(3206)));
    outputs(9215) <= layer0_outputs(6735);
    outputs(9216) <= (layer0_outputs(368)) xor (layer0_outputs(4885));
    outputs(9217) <= (layer0_outputs(4591)) xor (layer0_outputs(7175));
    outputs(9218) <= (layer0_outputs(6724)) and (layer0_outputs(7982));
    outputs(9219) <= layer0_outputs(8004);
    outputs(9220) <= not(layer0_outputs(1139)) or (layer0_outputs(2802));
    outputs(9221) <= not(layer0_outputs(1781)) or (layer0_outputs(295));
    outputs(9222) <= (layer0_outputs(7443)) and (layer0_outputs(8826));
    outputs(9223) <= (layer0_outputs(6901)) and not (layer0_outputs(1648));
    outputs(9224) <= (layer0_outputs(5624)) and (layer0_outputs(3601));
    outputs(9225) <= not((layer0_outputs(3992)) xor (layer0_outputs(12244)));
    outputs(9226) <= layer0_outputs(2808);
    outputs(9227) <= (layer0_outputs(1661)) and not (layer0_outputs(12136));
    outputs(9228) <= not(layer0_outputs(111)) or (layer0_outputs(6644));
    outputs(9229) <= not(layer0_outputs(9892));
    outputs(9230) <= (layer0_outputs(8932)) and not (layer0_outputs(5833));
    outputs(9231) <= not((layer0_outputs(10016)) xor (layer0_outputs(11830)));
    outputs(9232) <= layer0_outputs(547);
    outputs(9233) <= not((layer0_outputs(6000)) or (layer0_outputs(10877)));
    outputs(9234) <= not(layer0_outputs(9163));
    outputs(9235) <= layer0_outputs(9097);
    outputs(9236) <= layer0_outputs(4835);
    outputs(9237) <= layer0_outputs(110);
    outputs(9238) <= layer0_outputs(10066);
    outputs(9239) <= not(layer0_outputs(5759));
    outputs(9240) <= layer0_outputs(9177);
    outputs(9241) <= (layer0_outputs(12529)) and not (layer0_outputs(3562));
    outputs(9242) <= (layer0_outputs(6437)) and not (layer0_outputs(8806));
    outputs(9243) <= not(layer0_outputs(7833));
    outputs(9244) <= layer0_outputs(9655);
    outputs(9245) <= not(layer0_outputs(4138));
    outputs(9246) <= not(layer0_outputs(1729));
    outputs(9247) <= not(layer0_outputs(11238));
    outputs(9248) <= not(layer0_outputs(52)) or (layer0_outputs(760));
    outputs(9249) <= not((layer0_outputs(659)) xor (layer0_outputs(7446)));
    outputs(9250) <= (layer0_outputs(707)) and not (layer0_outputs(609));
    outputs(9251) <= not((layer0_outputs(12112)) xor (layer0_outputs(9016)));
    outputs(9252) <= not(layer0_outputs(11692));
    outputs(9253) <= not(layer0_outputs(7654));
    outputs(9254) <= (layer0_outputs(109)) xor (layer0_outputs(5036));
    outputs(9255) <= (layer0_outputs(2555)) and (layer0_outputs(6495));
    outputs(9256) <= not((layer0_outputs(4778)) and (layer0_outputs(3048)));
    outputs(9257) <= not((layer0_outputs(9200)) xor (layer0_outputs(5436)));
    outputs(9258) <= not(layer0_outputs(2007));
    outputs(9259) <= (layer0_outputs(5176)) and not (layer0_outputs(9700));
    outputs(9260) <= not(layer0_outputs(5882)) or (layer0_outputs(1973));
    outputs(9261) <= layer0_outputs(10485);
    outputs(9262) <= (layer0_outputs(2681)) xor (layer0_outputs(9949));
    outputs(9263) <= not((layer0_outputs(9895)) and (layer0_outputs(3921)));
    outputs(9264) <= (layer0_outputs(4921)) xor (layer0_outputs(6527));
    outputs(9265) <= not(layer0_outputs(11873));
    outputs(9266) <= (layer0_outputs(8232)) xor (layer0_outputs(15));
    outputs(9267) <= (layer0_outputs(12199)) and (layer0_outputs(10689));
    outputs(9268) <= not(layer0_outputs(1670));
    outputs(9269) <= not(layer0_outputs(12263)) or (layer0_outputs(8939));
    outputs(9270) <= not(layer0_outputs(7092));
    outputs(9271) <= layer0_outputs(7284);
    outputs(9272) <= (layer0_outputs(10906)) xor (layer0_outputs(1954));
    outputs(9273) <= layer0_outputs(6184);
    outputs(9274) <= not(layer0_outputs(9000));
    outputs(9275) <= not(layer0_outputs(385));
    outputs(9276) <= layer0_outputs(6287);
    outputs(9277) <= (layer0_outputs(3508)) and not (layer0_outputs(6124));
    outputs(9278) <= (layer0_outputs(7642)) and not (layer0_outputs(4871));
    outputs(9279) <= not(layer0_outputs(12517)) or (layer0_outputs(1665));
    outputs(9280) <= layer0_outputs(3208);
    outputs(9281) <= not((layer0_outputs(9673)) xor (layer0_outputs(12794)));
    outputs(9282) <= not((layer0_outputs(3132)) or (layer0_outputs(4049)));
    outputs(9283) <= not(layer0_outputs(3869));
    outputs(9284) <= not((layer0_outputs(7477)) xor (layer0_outputs(3721)));
    outputs(9285) <= not((layer0_outputs(8169)) xor (layer0_outputs(11914)));
    outputs(9286) <= not(layer0_outputs(4612));
    outputs(9287) <= not((layer0_outputs(3294)) or (layer0_outputs(9580)));
    outputs(9288) <= (layer0_outputs(6839)) and not (layer0_outputs(4217));
    outputs(9289) <= not((layer0_outputs(3594)) and (layer0_outputs(5344)));
    outputs(9290) <= layer0_outputs(2458);
    outputs(9291) <= not(layer0_outputs(11405));
    outputs(9292) <= not(layer0_outputs(9210)) or (layer0_outputs(7794));
    outputs(9293) <= not((layer0_outputs(9303)) xor (layer0_outputs(11176)));
    outputs(9294) <= (layer0_outputs(10178)) xor (layer0_outputs(1104));
    outputs(9295) <= (layer0_outputs(5958)) and not (layer0_outputs(8803));
    outputs(9296) <= (layer0_outputs(10656)) and not (layer0_outputs(4471));
    outputs(9297) <= (layer0_outputs(11511)) and not (layer0_outputs(1605));
    outputs(9298) <= (layer0_outputs(10495)) and (layer0_outputs(5520));
    outputs(9299) <= not(layer0_outputs(2846));
    outputs(9300) <= not((layer0_outputs(2821)) xor (layer0_outputs(6622)));
    outputs(9301) <= (layer0_outputs(8061)) and not (layer0_outputs(5963));
    outputs(9302) <= layer0_outputs(11046);
    outputs(9303) <= not(layer0_outputs(4933));
    outputs(9304) <= (layer0_outputs(12162)) or (layer0_outputs(6330));
    outputs(9305) <= not(layer0_outputs(297));
    outputs(9306) <= layer0_outputs(12280);
    outputs(9307) <= (layer0_outputs(11644)) and (layer0_outputs(3024));
    outputs(9308) <= (layer0_outputs(7162)) xor (layer0_outputs(1470));
    outputs(9309) <= not((layer0_outputs(9274)) xor (layer0_outputs(11120)));
    outputs(9310) <= not((layer0_outputs(12278)) or (layer0_outputs(10819)));
    outputs(9311) <= (layer0_outputs(9885)) xor (layer0_outputs(8463));
    outputs(9312) <= (layer0_outputs(11822)) xor (layer0_outputs(10868));
    outputs(9313) <= layer0_outputs(1743);
    outputs(9314) <= (layer0_outputs(8503)) and (layer0_outputs(4563));
    outputs(9315) <= (layer0_outputs(9578)) and not (layer0_outputs(1405));
    outputs(9316) <= (layer0_outputs(12449)) and (layer0_outputs(5062));
    outputs(9317) <= not(layer0_outputs(6429));
    outputs(9318) <= layer0_outputs(5641);
    outputs(9319) <= layer0_outputs(2669);
    outputs(9320) <= layer0_outputs(1173);
    outputs(9321) <= layer0_outputs(9799);
    outputs(9322) <= (layer0_outputs(2073)) xor (layer0_outputs(7524));
    outputs(9323) <= (layer0_outputs(10803)) and not (layer0_outputs(10325));
    outputs(9324) <= not((layer0_outputs(3925)) xor (layer0_outputs(9119)));
    outputs(9325) <= not((layer0_outputs(8949)) or (layer0_outputs(10312)));
    outputs(9326) <= (layer0_outputs(7792)) and (layer0_outputs(3144));
    outputs(9327) <= (layer0_outputs(7455)) xor (layer0_outputs(10648));
    outputs(9328) <= layer0_outputs(6674);
    outputs(9329) <= not(layer0_outputs(9414)) or (layer0_outputs(1895));
    outputs(9330) <= not((layer0_outputs(10361)) xor (layer0_outputs(2049)));
    outputs(9331) <= (layer0_outputs(7580)) and not (layer0_outputs(9826));
    outputs(9332) <= not((layer0_outputs(10089)) or (layer0_outputs(8414)));
    outputs(9333) <= not(layer0_outputs(12443)) or (layer0_outputs(13));
    outputs(9334) <= (layer0_outputs(11861)) xor (layer0_outputs(11963));
    outputs(9335) <= layer0_outputs(1901);
    outputs(9336) <= layer0_outputs(2894);
    outputs(9337) <= (layer0_outputs(12301)) and not (layer0_outputs(2426));
    outputs(9338) <= (layer0_outputs(3347)) and (layer0_outputs(4009));
    outputs(9339) <= not(layer0_outputs(1961));
    outputs(9340) <= not((layer0_outputs(11114)) xor (layer0_outputs(3239)));
    outputs(9341) <= (layer0_outputs(11697)) and not (layer0_outputs(19));
    outputs(9342) <= layer0_outputs(6786);
    outputs(9343) <= not(layer0_outputs(8451));
    outputs(9344) <= not((layer0_outputs(9203)) xor (layer0_outputs(12787)));
    outputs(9345) <= not((layer0_outputs(3269)) or (layer0_outputs(243)));
    outputs(9346) <= not((layer0_outputs(7317)) xor (layer0_outputs(2124)));
    outputs(9347) <= not(layer0_outputs(9297));
    outputs(9348) <= layer0_outputs(12107);
    outputs(9349) <= layer0_outputs(6343);
    outputs(9350) <= not((layer0_outputs(2850)) xor (layer0_outputs(12048)));
    outputs(9351) <= (layer0_outputs(7898)) or (layer0_outputs(8172));
    outputs(9352) <= not(layer0_outputs(3313));
    outputs(9353) <= layer0_outputs(6261);
    outputs(9354) <= layer0_outputs(1370);
    outputs(9355) <= not(layer0_outputs(4797));
    outputs(9356) <= not(layer0_outputs(5079));
    outputs(9357) <= not(layer0_outputs(10561));
    outputs(9358) <= not((layer0_outputs(3933)) xor (layer0_outputs(8769)));
    outputs(9359) <= not(layer0_outputs(4868));
    outputs(9360) <= (layer0_outputs(179)) and not (layer0_outputs(3627));
    outputs(9361) <= not(layer0_outputs(6175));
    outputs(9362) <= (layer0_outputs(8997)) xor (layer0_outputs(805));
    outputs(9363) <= (layer0_outputs(1800)) xor (layer0_outputs(6140));
    outputs(9364) <= (layer0_outputs(3025)) xor (layer0_outputs(2471));
    outputs(9365) <= (layer0_outputs(10453)) xor (layer0_outputs(2623));
    outputs(9366) <= layer0_outputs(489);
    outputs(9367) <= not(layer0_outputs(9849));
    outputs(9368) <= layer0_outputs(3993);
    outputs(9369) <= not((layer0_outputs(7862)) xor (layer0_outputs(1502)));
    outputs(9370) <= (layer0_outputs(8948)) and not (layer0_outputs(7687));
    outputs(9371) <= layer0_outputs(12310);
    outputs(9372) <= (layer0_outputs(6045)) and (layer0_outputs(11294));
    outputs(9373) <= not((layer0_outputs(3181)) xor (layer0_outputs(1108)));
    outputs(9374) <= not((layer0_outputs(11219)) xor (layer0_outputs(9274)));
    outputs(9375) <= not(layer0_outputs(7011));
    outputs(9376) <= not(layer0_outputs(4761));
    outputs(9377) <= not(layer0_outputs(2503));
    outputs(9378) <= (layer0_outputs(6999)) and not (layer0_outputs(11891));
    outputs(9379) <= not(layer0_outputs(8694));
    outputs(9380) <= (layer0_outputs(11568)) and (layer0_outputs(2823));
    outputs(9381) <= layer0_outputs(8273);
    outputs(9382) <= (layer0_outputs(5300)) xor (layer0_outputs(10266));
    outputs(9383) <= layer0_outputs(12466);
    outputs(9384) <= not(layer0_outputs(11143)) or (layer0_outputs(7441));
    outputs(9385) <= not((layer0_outputs(2690)) or (layer0_outputs(6580)));
    outputs(9386) <= not(layer0_outputs(7121));
    outputs(9387) <= (layer0_outputs(11571)) and not (layer0_outputs(9738));
    outputs(9388) <= (layer0_outputs(7549)) xor (layer0_outputs(4949));
    outputs(9389) <= layer0_outputs(8087);
    outputs(9390) <= layer0_outputs(12750);
    outputs(9391) <= (layer0_outputs(11982)) and (layer0_outputs(4936));
    outputs(9392) <= not((layer0_outputs(8113)) and (layer0_outputs(10548)));
    outputs(9393) <= not(layer0_outputs(5298)) or (layer0_outputs(6169));
    outputs(9394) <= (layer0_outputs(7738)) and not (layer0_outputs(9157));
    outputs(9395) <= layer0_outputs(6300);
    outputs(9396) <= not(layer0_outputs(10798));
    outputs(9397) <= (layer0_outputs(5779)) and (layer0_outputs(10121));
    outputs(9398) <= (layer0_outputs(10873)) and not (layer0_outputs(3544));
    outputs(9399) <= (layer0_outputs(5798)) and not (layer0_outputs(1277));
    outputs(9400) <= (layer0_outputs(8066)) or (layer0_outputs(12064));
    outputs(9401) <= (layer0_outputs(1184)) and not (layer0_outputs(4145));
    outputs(9402) <= not(layer0_outputs(2476));
    outputs(9403) <= not((layer0_outputs(3504)) xor (layer0_outputs(927)));
    outputs(9404) <= not((layer0_outputs(10817)) xor (layer0_outputs(8576)));
    outputs(9405) <= (layer0_outputs(9145)) xor (layer0_outputs(3379));
    outputs(9406) <= not(layer0_outputs(11074));
    outputs(9407) <= (layer0_outputs(4605)) and not (layer0_outputs(8189));
    outputs(9408) <= not((layer0_outputs(5594)) xor (layer0_outputs(9729)));
    outputs(9409) <= not((layer0_outputs(4141)) or (layer0_outputs(11755)));
    outputs(9410) <= layer0_outputs(11411);
    outputs(9411) <= layer0_outputs(6690);
    outputs(9412) <= layer0_outputs(6264);
    outputs(9413) <= not((layer0_outputs(350)) xor (layer0_outputs(8935)));
    outputs(9414) <= not(layer0_outputs(5834)) or (layer0_outputs(426));
    outputs(9415) <= not((layer0_outputs(1179)) or (layer0_outputs(10461)));
    outputs(9416) <= layer0_outputs(320);
    outputs(9417) <= not(layer0_outputs(732));
    outputs(9418) <= not((layer0_outputs(4226)) xor (layer0_outputs(10190)));
    outputs(9419) <= not(layer0_outputs(11678)) or (layer0_outputs(4733));
    outputs(9420) <= not(layer0_outputs(12489));
    outputs(9421) <= not(layer0_outputs(2619));
    outputs(9422) <= layer0_outputs(1978);
    outputs(9423) <= layer0_outputs(10260);
    outputs(9424) <= not(layer0_outputs(11207));
    outputs(9425) <= layer0_outputs(10954);
    outputs(9426) <= (layer0_outputs(10873)) xor (layer0_outputs(5438));
    outputs(9427) <= not(layer0_outputs(12178)) or (layer0_outputs(2202));
    outputs(9428) <= not(layer0_outputs(3771));
    outputs(9429) <= not(layer0_outputs(11906));
    outputs(9430) <= (layer0_outputs(7921)) xor (layer0_outputs(11538));
    outputs(9431) <= not(layer0_outputs(10411));
    outputs(9432) <= (layer0_outputs(3104)) and (layer0_outputs(8589));
    outputs(9433) <= not((layer0_outputs(9924)) and (layer0_outputs(8587)));
    outputs(9434) <= (layer0_outputs(3098)) and not (layer0_outputs(340));
    outputs(9435) <= layer0_outputs(12711);
    outputs(9436) <= (layer0_outputs(376)) and not (layer0_outputs(7506));
    outputs(9437) <= (layer0_outputs(2578)) xor (layer0_outputs(3426));
    outputs(9438) <= not(layer0_outputs(7428));
    outputs(9439) <= layer0_outputs(7297);
    outputs(9440) <= layer0_outputs(1449);
    outputs(9441) <= not(layer0_outputs(10086));
    outputs(9442) <= layer0_outputs(5178);
    outputs(9443) <= (layer0_outputs(2412)) or (layer0_outputs(4676));
    outputs(9444) <= not(layer0_outputs(10333)) or (layer0_outputs(5407));
    outputs(9445) <= layer0_outputs(10386);
    outputs(9446) <= layer0_outputs(6186);
    outputs(9447) <= layer0_outputs(6422);
    outputs(9448) <= not((layer0_outputs(11309)) xor (layer0_outputs(195)));
    outputs(9449) <= (layer0_outputs(2746)) and not (layer0_outputs(4311));
    outputs(9450) <= not((layer0_outputs(12468)) xor (layer0_outputs(1418)));
    outputs(9451) <= not((layer0_outputs(11279)) or (layer0_outputs(11393)));
    outputs(9452) <= (layer0_outputs(6526)) and not (layer0_outputs(7987));
    outputs(9453) <= (layer0_outputs(11582)) and not (layer0_outputs(6632));
    outputs(9454) <= (layer0_outputs(12746)) and (layer0_outputs(12753));
    outputs(9455) <= (layer0_outputs(3333)) and not (layer0_outputs(10175));
    outputs(9456) <= not((layer0_outputs(1934)) xor (layer0_outputs(10151)));
    outputs(9457) <= layer0_outputs(11106);
    outputs(9458) <= layer0_outputs(2882);
    outputs(9459) <= (layer0_outputs(2786)) and (layer0_outputs(3638));
    outputs(9460) <= layer0_outputs(12140);
    outputs(9461) <= (layer0_outputs(3399)) xor (layer0_outputs(4519));
    outputs(9462) <= (layer0_outputs(8340)) and not (layer0_outputs(5302));
    outputs(9463) <= layer0_outputs(3731);
    outputs(9464) <= not(layer0_outputs(8305));
    outputs(9465) <= not(layer0_outputs(8806));
    outputs(9466) <= layer0_outputs(9527);
    outputs(9467) <= not((layer0_outputs(12189)) or (layer0_outputs(11769)));
    outputs(9468) <= not(layer0_outputs(1019));
    outputs(9469) <= not((layer0_outputs(12772)) xor (layer0_outputs(7619)));
    outputs(9470) <= not(layer0_outputs(7562)) or (layer0_outputs(8036));
    outputs(9471) <= (layer0_outputs(9326)) and (layer0_outputs(5420));
    outputs(9472) <= not((layer0_outputs(2114)) xor (layer0_outputs(3950)));
    outputs(9473) <= (layer0_outputs(5822)) or (layer0_outputs(9096));
    outputs(9474) <= not((layer0_outputs(11775)) xor (layer0_outputs(3960)));
    outputs(9475) <= (layer0_outputs(8455)) xor (layer0_outputs(3749));
    outputs(9476) <= (layer0_outputs(3867)) xor (layer0_outputs(11152));
    outputs(9477) <= layer0_outputs(6148);
    outputs(9478) <= (layer0_outputs(2390)) and (layer0_outputs(10760));
    outputs(9479) <= not(layer0_outputs(8189)) or (layer0_outputs(20));
    outputs(9480) <= (layer0_outputs(2391)) and not (layer0_outputs(1153));
    outputs(9481) <= (layer0_outputs(898)) and (layer0_outputs(7069));
    outputs(9482) <= not((layer0_outputs(5988)) xor (layer0_outputs(2210)));
    outputs(9483) <= layer0_outputs(4304);
    outputs(9484) <= not((layer0_outputs(1530)) xor (layer0_outputs(225)));
    outputs(9485) <= not((layer0_outputs(6545)) xor (layer0_outputs(8025)));
    outputs(9486) <= not((layer0_outputs(2494)) or (layer0_outputs(12474)));
    outputs(9487) <= (layer0_outputs(10224)) xor (layer0_outputs(9266));
    outputs(9488) <= layer0_outputs(7202);
    outputs(9489) <= not((layer0_outputs(8361)) xor (layer0_outputs(6844)));
    outputs(9490) <= not((layer0_outputs(12166)) xor (layer0_outputs(3711)));
    outputs(9491) <= not((layer0_outputs(8859)) xor (layer0_outputs(2139)));
    outputs(9492) <= (layer0_outputs(9701)) and (layer0_outputs(1761));
    outputs(9493) <= layer0_outputs(1524);
    outputs(9494) <= not((layer0_outputs(6283)) xor (layer0_outputs(6234)));
    outputs(9495) <= not(layer0_outputs(10350));
    outputs(9496) <= layer0_outputs(1043);
    outputs(9497) <= not(layer0_outputs(4854));
    outputs(9498) <= not((layer0_outputs(3259)) or (layer0_outputs(5430)));
    outputs(9499) <= not((layer0_outputs(12376)) or (layer0_outputs(10185)));
    outputs(9500) <= layer0_outputs(12123);
    outputs(9501) <= (layer0_outputs(1533)) or (layer0_outputs(2009));
    outputs(9502) <= layer0_outputs(10567);
    outputs(9503) <= not((layer0_outputs(1178)) xor (layer0_outputs(4986)));
    outputs(9504) <= not((layer0_outputs(934)) or (layer0_outputs(10514)));
    outputs(9505) <= not(layer0_outputs(8701)) or (layer0_outputs(9244));
    outputs(9506) <= not(layer0_outputs(4691)) or (layer0_outputs(6167));
    outputs(9507) <= (layer0_outputs(12144)) and not (layer0_outputs(8496));
    outputs(9508) <= not(layer0_outputs(5649));
    outputs(9509) <= layer0_outputs(9584);
    outputs(9510) <= not(layer0_outputs(2811));
    outputs(9511) <= (layer0_outputs(2134)) and not (layer0_outputs(342));
    outputs(9512) <= (layer0_outputs(6524)) and not (layer0_outputs(1066));
    outputs(9513) <= layer0_outputs(5228);
    outputs(9514) <= (layer0_outputs(11925)) or (layer0_outputs(5155));
    outputs(9515) <= layer0_outputs(7783);
    outputs(9516) <= (layer0_outputs(9765)) or (layer0_outputs(3215));
    outputs(9517) <= (layer0_outputs(4135)) xor (layer0_outputs(4112));
    outputs(9518) <= (layer0_outputs(11401)) and not (layer0_outputs(11824));
    outputs(9519) <= not((layer0_outputs(11810)) xor (layer0_outputs(9432)));
    outputs(9520) <= not(layer0_outputs(1325)) or (layer0_outputs(5590));
    outputs(9521) <= (layer0_outputs(4649)) and (layer0_outputs(1765));
    outputs(9522) <= not((layer0_outputs(4596)) xor (layer0_outputs(9853)));
    outputs(9523) <= not(layer0_outputs(80));
    outputs(9524) <= not((layer0_outputs(3047)) xor (layer0_outputs(11690)));
    outputs(9525) <= (layer0_outputs(309)) xor (layer0_outputs(452));
    outputs(9526) <= not(layer0_outputs(1770));
    outputs(9527) <= not(layer0_outputs(12520));
    outputs(9528) <= not((layer0_outputs(3005)) xor (layer0_outputs(731)));
    outputs(9529) <= layer0_outputs(9185);
    outputs(9530) <= not(layer0_outputs(11993));
    outputs(9531) <= (layer0_outputs(1358)) and (layer0_outputs(12557));
    outputs(9532) <= not(layer0_outputs(5479)) or (layer0_outputs(2301));
    outputs(9533) <= (layer0_outputs(404)) and not (layer0_outputs(8738));
    outputs(9534) <= layer0_outputs(5569);
    outputs(9535) <= not(layer0_outputs(5121));
    outputs(9536) <= (layer0_outputs(10971)) or (layer0_outputs(4810));
    outputs(9537) <= not((layer0_outputs(11292)) or (layer0_outputs(1301)));
    outputs(9538) <= not(layer0_outputs(1717));
    outputs(9539) <= not(layer0_outputs(8131));
    outputs(9540) <= not((layer0_outputs(5027)) xor (layer0_outputs(1727)));
    outputs(9541) <= not(layer0_outputs(5121));
    outputs(9542) <= not(layer0_outputs(5195));
    outputs(9543) <= not(layer0_outputs(7247));
    outputs(9544) <= (layer0_outputs(8913)) xor (layer0_outputs(7433));
    outputs(9545) <= (layer0_outputs(6293)) xor (layer0_outputs(4231));
    outputs(9546) <= not(layer0_outputs(10806));
    outputs(9547) <= not((layer0_outputs(12617)) or (layer0_outputs(7076)));
    outputs(9548) <= layer0_outputs(12711);
    outputs(9549) <= (layer0_outputs(1994)) xor (layer0_outputs(6970));
    outputs(9550) <= (layer0_outputs(1471)) and not (layer0_outputs(5080));
    outputs(9551) <= not(layer0_outputs(5164));
    outputs(9552) <= not(layer0_outputs(4566));
    outputs(9553) <= (layer0_outputs(5552)) xor (layer0_outputs(10261));
    outputs(9554) <= (layer0_outputs(8918)) and not (layer0_outputs(9775));
    outputs(9555) <= layer0_outputs(4532);
    outputs(9556) <= not((layer0_outputs(3336)) xor (layer0_outputs(8372)));
    outputs(9557) <= (layer0_outputs(10632)) xor (layer0_outputs(11761));
    outputs(9558) <= layer0_outputs(12033);
    outputs(9559) <= not((layer0_outputs(8427)) and (layer0_outputs(6832)));
    outputs(9560) <= (layer0_outputs(11852)) and not (layer0_outputs(6520));
    outputs(9561) <= not(layer0_outputs(5103)) or (layer0_outputs(9765));
    outputs(9562) <= layer0_outputs(7913);
    outputs(9563) <= layer0_outputs(3281);
    outputs(9564) <= not(layer0_outputs(9449)) or (layer0_outputs(3642));
    outputs(9565) <= layer0_outputs(821);
    outputs(9566) <= not((layer0_outputs(196)) and (layer0_outputs(6315)));
    outputs(9567) <= (layer0_outputs(9680)) xor (layer0_outputs(1164));
    outputs(9568) <= (layer0_outputs(6488)) and not (layer0_outputs(1452));
    outputs(9569) <= (layer0_outputs(9418)) xor (layer0_outputs(3043));
    outputs(9570) <= not(layer0_outputs(4714));
    outputs(9571) <= (layer0_outputs(10256)) xor (layer0_outputs(2906));
    outputs(9572) <= not(layer0_outputs(11223)) or (layer0_outputs(3070));
    outputs(9573) <= not((layer0_outputs(12647)) or (layer0_outputs(12028)));
    outputs(9574) <= (layer0_outputs(9062)) xor (layer0_outputs(7759));
    outputs(9575) <= not(layer0_outputs(11785));
    outputs(9576) <= not(layer0_outputs(710));
    outputs(9577) <= (layer0_outputs(6643)) and not (layer0_outputs(12020));
    outputs(9578) <= (layer0_outputs(5966)) and (layer0_outputs(8707));
    outputs(9579) <= (layer0_outputs(8631)) xor (layer0_outputs(12756));
    outputs(9580) <= not(layer0_outputs(7673));
    outputs(9581) <= (layer0_outputs(5104)) xor (layer0_outputs(5592));
    outputs(9582) <= layer0_outputs(3317);
    outputs(9583) <= not(layer0_outputs(4560));
    outputs(9584) <= not(layer0_outputs(5042));
    outputs(9585) <= not((layer0_outputs(2459)) or (layer0_outputs(2769)));
    outputs(9586) <= not((layer0_outputs(8262)) or (layer0_outputs(1451)));
    outputs(9587) <= not(layer0_outputs(8270));
    outputs(9588) <= layer0_outputs(2328);
    outputs(9589) <= not(layer0_outputs(10990));
    outputs(9590) <= (layer0_outputs(10752)) xor (layer0_outputs(1860));
    outputs(9591) <= (layer0_outputs(408)) or (layer0_outputs(7322));
    outputs(9592) <= not((layer0_outputs(9644)) xor (layer0_outputs(661)));
    outputs(9593) <= layer0_outputs(6099);
    outputs(9594) <= layer0_outputs(4442);
    outputs(9595) <= layer0_outputs(10897);
    outputs(9596) <= layer0_outputs(7835);
    outputs(9597) <= not((layer0_outputs(10623)) xor (layer0_outputs(4784)));
    outputs(9598) <= not(layer0_outputs(2385));
    outputs(9599) <= (layer0_outputs(8228)) and (layer0_outputs(6691));
    outputs(9600) <= not(layer0_outputs(5045)) or (layer0_outputs(7705));
    outputs(9601) <= layer0_outputs(11054);
    outputs(9602) <= layer0_outputs(1618);
    outputs(9603) <= not(layer0_outputs(9848));
    outputs(9604) <= not(layer0_outputs(2280));
    outputs(9605) <= not(layer0_outputs(6920));
    outputs(9606) <= (layer0_outputs(10338)) and (layer0_outputs(2020));
    outputs(9607) <= (layer0_outputs(9370)) xor (layer0_outputs(8331));
    outputs(9608) <= not((layer0_outputs(1303)) or (layer0_outputs(2920)));
    outputs(9609) <= layer0_outputs(9604);
    outputs(9610) <= not((layer0_outputs(134)) or (layer0_outputs(206)));
    outputs(9611) <= (layer0_outputs(4445)) and not (layer0_outputs(4662));
    outputs(9612) <= not(layer0_outputs(2267));
    outputs(9613) <= not(layer0_outputs(3218));
    outputs(9614) <= not(layer0_outputs(12455));
    outputs(9615) <= (layer0_outputs(776)) and not (layer0_outputs(7396));
    outputs(9616) <= (layer0_outputs(5331)) and (layer0_outputs(4753));
    outputs(9617) <= layer0_outputs(3723);
    outputs(9618) <= not(layer0_outputs(12385));
    outputs(9619) <= (layer0_outputs(11171)) and (layer0_outputs(5838));
    outputs(9620) <= (layer0_outputs(10553)) xor (layer0_outputs(11023));
    outputs(9621) <= layer0_outputs(9100);
    outputs(9622) <= not(layer0_outputs(1649));
    outputs(9623) <= (layer0_outputs(9188)) and (layer0_outputs(3527));
    outputs(9624) <= (layer0_outputs(7546)) and (layer0_outputs(8521));
    outputs(9625) <= layer0_outputs(133);
    outputs(9626) <= layer0_outputs(9583);
    outputs(9627) <= not((layer0_outputs(9292)) or (layer0_outputs(3196)));
    outputs(9628) <= (layer0_outputs(11057)) and not (layer0_outputs(11205));
    outputs(9629) <= (layer0_outputs(10459)) and (layer0_outputs(4348));
    outputs(9630) <= not((layer0_outputs(8927)) xor (layer0_outputs(8654)));
    outputs(9631) <= (layer0_outputs(3488)) and not (layer0_outputs(3563));
    outputs(9632) <= not((layer0_outputs(3577)) xor (layer0_outputs(6392)));
    outputs(9633) <= not(layer0_outputs(3906));
    outputs(9634) <= layer0_outputs(6092);
    outputs(9635) <= (layer0_outputs(10960)) and not (layer0_outputs(3771));
    outputs(9636) <= (layer0_outputs(1109)) and not (layer0_outputs(8596));
    outputs(9637) <= (layer0_outputs(7497)) and not (layer0_outputs(11880));
    outputs(9638) <= (layer0_outputs(12367)) xor (layer0_outputs(12497));
    outputs(9639) <= not((layer0_outputs(7458)) and (layer0_outputs(7514)));
    outputs(9640) <= (layer0_outputs(3223)) and not (layer0_outputs(2830));
    outputs(9641) <= not(layer0_outputs(6199)) or (layer0_outputs(2732));
    outputs(9642) <= not(layer0_outputs(9741));
    outputs(9643) <= layer0_outputs(2109);
    outputs(9644) <= layer0_outputs(9899);
    outputs(9645) <= not(layer0_outputs(203));
    outputs(9646) <= layer0_outputs(276);
    outputs(9647) <= (layer0_outputs(6443)) and not (layer0_outputs(4574));
    outputs(9648) <= (layer0_outputs(1550)) and not (layer0_outputs(6459));
    outputs(9649) <= (layer0_outputs(5493)) xor (layer0_outputs(1541));
    outputs(9650) <= (layer0_outputs(5168)) and not (layer0_outputs(4697));
    outputs(9651) <= not(layer0_outputs(10162));
    outputs(9652) <= layer0_outputs(8927);
    outputs(9653) <= not(layer0_outputs(1209));
    outputs(9654) <= (layer0_outputs(2504)) and not (layer0_outputs(1166));
    outputs(9655) <= (layer0_outputs(1170)) and (layer0_outputs(9581));
    outputs(9656) <= not(layer0_outputs(9685));
    outputs(9657) <= not((layer0_outputs(4828)) xor (layer0_outputs(2893)));
    outputs(9658) <= (layer0_outputs(338)) and not (layer0_outputs(348));
    outputs(9659) <= layer0_outputs(7369);
    outputs(9660) <= layer0_outputs(10079);
    outputs(9661) <= layer0_outputs(7262);
    outputs(9662) <= layer0_outputs(4165);
    outputs(9663) <= not(layer0_outputs(8687)) or (layer0_outputs(11475));
    outputs(9664) <= not(layer0_outputs(2209));
    outputs(9665) <= layer0_outputs(11905);
    outputs(9666) <= (layer0_outputs(3135)) xor (layer0_outputs(5784));
    outputs(9667) <= not((layer0_outputs(4564)) xor (layer0_outputs(8662)));
    outputs(9668) <= (layer0_outputs(12733)) and not (layer0_outputs(531));
    outputs(9669) <= (layer0_outputs(7331)) xor (layer0_outputs(7233));
    outputs(9670) <= (layer0_outputs(8487)) and not (layer0_outputs(1183));
    outputs(9671) <= (layer0_outputs(2236)) and not (layer0_outputs(12496));
    outputs(9672) <= (layer0_outputs(12566)) and not (layer0_outputs(215));
    outputs(9673) <= not((layer0_outputs(5631)) or (layer0_outputs(12244)));
    outputs(9674) <= layer0_outputs(4509);
    outputs(9675) <= not(layer0_outputs(9927));
    outputs(9676) <= layer0_outputs(6694);
    outputs(9677) <= (layer0_outputs(8429)) xor (layer0_outputs(6433));
    outputs(9678) <= not((layer0_outputs(8987)) xor (layer0_outputs(1548)));
    outputs(9679) <= not(layer0_outputs(11805));
    outputs(9680) <= not(layer0_outputs(10379));
    outputs(9681) <= not((layer0_outputs(289)) xor (layer0_outputs(9942)));
    outputs(9682) <= not(layer0_outputs(2290));
    outputs(9683) <= not((layer0_outputs(10328)) xor (layer0_outputs(3980)));
    outputs(9684) <= not((layer0_outputs(1706)) xor (layer0_outputs(10380)));
    outputs(9685) <= (layer0_outputs(12258)) or (layer0_outputs(6780));
    outputs(9686) <= not(layer0_outputs(12227));
    outputs(9687) <= not((layer0_outputs(9896)) xor (layer0_outputs(1097)));
    outputs(9688) <= layer0_outputs(6271);
    outputs(9689) <= not(layer0_outputs(6573));
    outputs(9690) <= (layer0_outputs(5156)) and not (layer0_outputs(10419));
    outputs(9691) <= not(layer0_outputs(5418));
    outputs(9692) <= (layer0_outputs(4655)) and (layer0_outputs(1024));
    outputs(9693) <= not((layer0_outputs(8536)) or (layer0_outputs(8526)));
    outputs(9694) <= not((layer0_outputs(1272)) xor (layer0_outputs(1861)));
    outputs(9695) <= (layer0_outputs(9916)) xor (layer0_outputs(2655));
    outputs(9696) <= not(layer0_outputs(12058));
    outputs(9697) <= (layer0_outputs(1805)) and not (layer0_outputs(2794));
    outputs(9698) <= layer0_outputs(10476);
    outputs(9699) <= layer0_outputs(173);
    outputs(9700) <= (layer0_outputs(12223)) xor (layer0_outputs(9995));
    outputs(9701) <= layer0_outputs(6468);
    outputs(9702) <= not(layer0_outputs(2929));
    outputs(9703) <= not((layer0_outputs(6425)) and (layer0_outputs(5164)));
    outputs(9704) <= (layer0_outputs(8423)) and (layer0_outputs(6488));
    outputs(9705) <= (layer0_outputs(5297)) and not (layer0_outputs(1848));
    outputs(9706) <= (layer0_outputs(8138)) xor (layer0_outputs(3234));
    outputs(9707) <= not(layer0_outputs(11251));
    outputs(9708) <= layer0_outputs(11651);
    outputs(9709) <= not(layer0_outputs(11041));
    outputs(9710) <= (layer0_outputs(4032)) and not (layer0_outputs(12263));
    outputs(9711) <= layer0_outputs(10424);
    outputs(9712) <= (layer0_outputs(7097)) xor (layer0_outputs(11008));
    outputs(9713) <= (layer0_outputs(5260)) and (layer0_outputs(2958));
    outputs(9714) <= layer0_outputs(2158);
    outputs(9715) <= (layer0_outputs(9008)) and not (layer0_outputs(12653));
    outputs(9716) <= not(layer0_outputs(8568));
    outputs(9717) <= (layer0_outputs(4689)) and (layer0_outputs(2947));
    outputs(9718) <= not(layer0_outputs(7520));
    outputs(9719) <= not(layer0_outputs(7342));
    outputs(9720) <= not(layer0_outputs(8864)) or (layer0_outputs(8429));
    outputs(9721) <= layer0_outputs(8598);
    outputs(9722) <= (layer0_outputs(2316)) and not (layer0_outputs(8294));
    outputs(9723) <= (layer0_outputs(1567)) and not (layer0_outputs(12550));
    outputs(9724) <= not(layer0_outputs(2046));
    outputs(9725) <= not(layer0_outputs(8613));
    outputs(9726) <= not(layer0_outputs(11912));
    outputs(9727) <= (layer0_outputs(7374)) and not (layer0_outputs(1614));
    outputs(9728) <= (layer0_outputs(6481)) and (layer0_outputs(798));
    outputs(9729) <= not(layer0_outputs(9500));
    outputs(9730) <= layer0_outputs(2489);
    outputs(9731) <= layer0_outputs(11688);
    outputs(9732) <= (layer0_outputs(5115)) and not (layer0_outputs(38));
    outputs(9733) <= (layer0_outputs(12019)) xor (layer0_outputs(8512));
    outputs(9734) <= not((layer0_outputs(6088)) and (layer0_outputs(9831)));
    outputs(9735) <= not((layer0_outputs(11731)) xor (layer0_outputs(55)));
    outputs(9736) <= (layer0_outputs(2983)) and not (layer0_outputs(10751));
    outputs(9737) <= not((layer0_outputs(8742)) xor (layer0_outputs(5412)));
    outputs(9738) <= layer0_outputs(11936);
    outputs(9739) <= not(layer0_outputs(3627));
    outputs(9740) <= layer0_outputs(9602);
    outputs(9741) <= not((layer0_outputs(3590)) xor (layer0_outputs(2118)));
    outputs(9742) <= (layer0_outputs(9033)) and not (layer0_outputs(3887));
    outputs(9743) <= not(layer0_outputs(9414)) or (layer0_outputs(8357));
    outputs(9744) <= layer0_outputs(48);
    outputs(9745) <= (layer0_outputs(12056)) xor (layer0_outputs(11907));
    outputs(9746) <= (layer0_outputs(6675)) xor (layer0_outputs(12513));
    outputs(9747) <= not(layer0_outputs(5718));
    outputs(9748) <= (layer0_outputs(7712)) and (layer0_outputs(12410));
    outputs(9749) <= (layer0_outputs(11736)) and (layer0_outputs(2557));
    outputs(9750) <= not((layer0_outputs(1338)) or (layer0_outputs(1027)));
    outputs(9751) <= (layer0_outputs(2271)) and (layer0_outputs(9330));
    outputs(9752) <= (layer0_outputs(1067)) and (layer0_outputs(10778));
    outputs(9753) <= (layer0_outputs(2833)) or (layer0_outputs(3973));
    outputs(9754) <= (layer0_outputs(10064)) xor (layer0_outputs(3744));
    outputs(9755) <= not((layer0_outputs(11048)) and (layer0_outputs(3773)));
    outputs(9756) <= (layer0_outputs(2555)) and not (layer0_outputs(10036));
    outputs(9757) <= not(layer0_outputs(5981));
    outputs(9758) <= layer0_outputs(7727);
    outputs(9759) <= layer0_outputs(6394);
    outputs(9760) <= not(layer0_outputs(4986));
    outputs(9761) <= not(layer0_outputs(8784));
    outputs(9762) <= layer0_outputs(4930);
    outputs(9763) <= not((layer0_outputs(4178)) or (layer0_outputs(12035)));
    outputs(9764) <= (layer0_outputs(6696)) xor (layer0_outputs(7600));
    outputs(9765) <= layer0_outputs(12627);
    outputs(9766) <= not(layer0_outputs(234));
    outputs(9767) <= layer0_outputs(11746);
    outputs(9768) <= layer0_outputs(2179);
    outputs(9769) <= (layer0_outputs(11197)) xor (layer0_outputs(413));
    outputs(9770) <= layer0_outputs(2888);
    outputs(9771) <= (layer0_outputs(2328)) and (layer0_outputs(852));
    outputs(9772) <= not(layer0_outputs(2056));
    outputs(9773) <= not(layer0_outputs(1328));
    outputs(9774) <= not((layer0_outputs(1098)) xor (layer0_outputs(168)));
    outputs(9775) <= not((layer0_outputs(4460)) or (layer0_outputs(2366)));
    outputs(9776) <= (layer0_outputs(6959)) and (layer0_outputs(8696));
    outputs(9777) <= not((layer0_outputs(4951)) xor (layer0_outputs(6279)));
    outputs(9778) <= (layer0_outputs(3314)) xor (layer0_outputs(11770));
    outputs(9779) <= not((layer0_outputs(10709)) xor (layer0_outputs(5926)));
    outputs(9780) <= layer0_outputs(9185);
    outputs(9781) <= (layer0_outputs(6128)) xor (layer0_outputs(5));
    outputs(9782) <= layer0_outputs(2291);
    outputs(9783) <= not(layer0_outputs(3617));
    outputs(9784) <= not((layer0_outputs(12323)) xor (layer0_outputs(11131)));
    outputs(9785) <= not(layer0_outputs(5907));
    outputs(9786) <= layer0_outputs(11437);
    outputs(9787) <= layer0_outputs(3737);
    outputs(9788) <= not((layer0_outputs(1782)) or (layer0_outputs(4947)));
    outputs(9789) <= layer0_outputs(6141);
    outputs(9790) <= (layer0_outputs(5163)) and not (layer0_outputs(424));
    outputs(9791) <= layer0_outputs(2181);
    outputs(9792) <= (layer0_outputs(10919)) xor (layer0_outputs(3950));
    outputs(9793) <= not((layer0_outputs(2727)) or (layer0_outputs(31)));
    outputs(9794) <= (layer0_outputs(12289)) xor (layer0_outputs(4350));
    outputs(9795) <= (layer0_outputs(12380)) and not (layer0_outputs(9474));
    outputs(9796) <= (layer0_outputs(4682)) and not (layer0_outputs(11208));
    outputs(9797) <= (layer0_outputs(8846)) and not (layer0_outputs(8049));
    outputs(9798) <= not((layer0_outputs(98)) and (layer0_outputs(5287)));
    outputs(9799) <= not(layer0_outputs(9741)) or (layer0_outputs(1116));
    outputs(9800) <= not(layer0_outputs(6226));
    outputs(9801) <= layer0_outputs(4264);
    outputs(9802) <= not((layer0_outputs(7837)) xor (layer0_outputs(11466)));
    outputs(9803) <= not(layer0_outputs(7959));
    outputs(9804) <= (layer0_outputs(7704)) and not (layer0_outputs(10196));
    outputs(9805) <= layer0_outputs(5142);
    outputs(9806) <= (layer0_outputs(11305)) xor (layer0_outputs(7702));
    outputs(9807) <= layer0_outputs(3233);
    outputs(9808) <= not(layer0_outputs(7685));
    outputs(9809) <= (layer0_outputs(3421)) xor (layer0_outputs(4482));
    outputs(9810) <= not(layer0_outputs(6069)) or (layer0_outputs(11864));
    outputs(9811) <= (layer0_outputs(1620)) or (layer0_outputs(10400));
    outputs(9812) <= not(layer0_outputs(11081));
    outputs(9813) <= layer0_outputs(9343);
    outputs(9814) <= layer0_outputs(2803);
    outputs(9815) <= (layer0_outputs(10583)) and not (layer0_outputs(3883));
    outputs(9816) <= (layer0_outputs(10845)) xor (layer0_outputs(6377));
    outputs(9817) <= not(layer0_outputs(3977));
    outputs(9818) <= (layer0_outputs(8879)) xor (layer0_outputs(3817));
    outputs(9819) <= layer0_outputs(5427);
    outputs(9820) <= not(layer0_outputs(11293));
    outputs(9821) <= (layer0_outputs(2478)) and (layer0_outputs(5364));
    outputs(9822) <= not(layer0_outputs(594));
    outputs(9823) <= (layer0_outputs(8181)) and (layer0_outputs(11088));
    outputs(9824) <= (layer0_outputs(6815)) xor (layer0_outputs(10914));
    outputs(9825) <= not((layer0_outputs(2931)) xor (layer0_outputs(4760)));
    outputs(9826) <= (layer0_outputs(8772)) and (layer0_outputs(9111));
    outputs(9827) <= layer0_outputs(9102);
    outputs(9828) <= (layer0_outputs(9475)) and (layer0_outputs(8894));
    outputs(9829) <= (layer0_outputs(7361)) and not (layer0_outputs(1295));
    outputs(9830) <= not(layer0_outputs(8484));
    outputs(9831) <= (layer0_outputs(9134)) and not (layer0_outputs(4277));
    outputs(9832) <= (layer0_outputs(1909)) xor (layer0_outputs(12431));
    outputs(9833) <= not((layer0_outputs(9000)) xor (layer0_outputs(11154)));
    outputs(9834) <= not(layer0_outputs(304));
    outputs(9835) <= not((layer0_outputs(9391)) xor (layer0_outputs(703)));
    outputs(9836) <= (layer0_outputs(6196)) and (layer0_outputs(1761));
    outputs(9837) <= layer0_outputs(1609);
    outputs(9838) <= not((layer0_outputs(5461)) or (layer0_outputs(1509)));
    outputs(9839) <= (layer0_outputs(12492)) xor (layer0_outputs(12745));
    outputs(9840) <= not(layer0_outputs(8537));
    outputs(9841) <= not(layer0_outputs(8148));
    outputs(9842) <= not(layer0_outputs(11670));
    outputs(9843) <= layer0_outputs(406);
    outputs(9844) <= not(layer0_outputs(5976));
    outputs(9845) <= (layer0_outputs(8135)) and not (layer0_outputs(3789));
    outputs(9846) <= not(layer0_outputs(10086));
    outputs(9847) <= layer0_outputs(10324);
    outputs(9848) <= not(layer0_outputs(6600));
    outputs(9849) <= (layer0_outputs(3372)) or (layer0_outputs(3128));
    outputs(9850) <= (layer0_outputs(10051)) and (layer0_outputs(3123));
    outputs(9851) <= not(layer0_outputs(2765));
    outputs(9852) <= not(layer0_outputs(4833)) or (layer0_outputs(5349));
    outputs(9853) <= layer0_outputs(3929);
    outputs(9854) <= (layer0_outputs(5545)) and not (layer0_outputs(1817));
    outputs(9855) <= (layer0_outputs(6249)) or (layer0_outputs(9231));
    outputs(9856) <= not(layer0_outputs(5932));
    outputs(9857) <= (layer0_outputs(11243)) xor (layer0_outputs(9744));
    outputs(9858) <= not((layer0_outputs(2436)) xor (layer0_outputs(7613)));
    outputs(9859) <= (layer0_outputs(5105)) xor (layer0_outputs(12524));
    outputs(9860) <= (layer0_outputs(2099)) and not (layer0_outputs(3021));
    outputs(9861) <= (layer0_outputs(4250)) and not (layer0_outputs(5307));
    outputs(9862) <= not((layer0_outputs(5340)) and (layer0_outputs(4333)));
    outputs(9863) <= not((layer0_outputs(4195)) xor (layer0_outputs(5186)));
    outputs(9864) <= not(layer0_outputs(3734)) or (layer0_outputs(2463));
    outputs(9865) <= not((layer0_outputs(11788)) or (layer0_outputs(4535)));
    outputs(9866) <= layer0_outputs(7098);
    outputs(9867) <= (layer0_outputs(6803)) or (layer0_outputs(10835));
    outputs(9868) <= layer0_outputs(9384);
    outputs(9869) <= not(layer0_outputs(3011));
    outputs(9870) <= (layer0_outputs(1850)) and not (layer0_outputs(1314));
    outputs(9871) <= layer0_outputs(3545);
    outputs(9872) <= not((layer0_outputs(3492)) xor (layer0_outputs(7338)));
    outputs(9873) <= not((layer0_outputs(463)) xor (layer0_outputs(3104)));
    outputs(9874) <= not(layer0_outputs(12368)) or (layer0_outputs(8328));
    outputs(9875) <= not((layer0_outputs(9293)) xor (layer0_outputs(1414)));
    outputs(9876) <= not(layer0_outputs(1129));
    outputs(9877) <= not((layer0_outputs(12407)) xor (layer0_outputs(2869)));
    outputs(9878) <= not(layer0_outputs(2221));
    outputs(9879) <= layer0_outputs(7975);
    outputs(9880) <= (layer0_outputs(9360)) or (layer0_outputs(10938));
    outputs(9881) <= not((layer0_outputs(6864)) xor (layer0_outputs(3914)));
    outputs(9882) <= not(layer0_outputs(9297));
    outputs(9883) <= not((layer0_outputs(5998)) or (layer0_outputs(8765)));
    outputs(9884) <= (layer0_outputs(7763)) xor (layer0_outputs(3713));
    outputs(9885) <= not((layer0_outputs(4364)) xor (layer0_outputs(785)));
    outputs(9886) <= layer0_outputs(2523);
    outputs(9887) <= (layer0_outputs(7413)) and (layer0_outputs(6344));
    outputs(9888) <= not(layer0_outputs(10213));
    outputs(9889) <= not(layer0_outputs(2474));
    outputs(9890) <= not((layer0_outputs(9831)) xor (layer0_outputs(12358)));
    outputs(9891) <= (layer0_outputs(307)) and not (layer0_outputs(113));
    outputs(9892) <= not(layer0_outputs(4323));
    outputs(9893) <= not((layer0_outputs(6105)) xor (layer0_outputs(9780)));
    outputs(9894) <= (layer0_outputs(6409)) and not (layer0_outputs(2450));
    outputs(9895) <= (layer0_outputs(3561)) xor (layer0_outputs(11525));
    outputs(9896) <= not(layer0_outputs(8829));
    outputs(9897) <= not((layer0_outputs(5282)) xor (layer0_outputs(8472)));
    outputs(9898) <= layer0_outputs(10272);
    outputs(9899) <= (layer0_outputs(6194)) or (layer0_outputs(6189));
    outputs(9900) <= layer0_outputs(8801);
    outputs(9901) <= layer0_outputs(11124);
    outputs(9902) <= not(layer0_outputs(8919));
    outputs(9903) <= (layer0_outputs(2315)) and (layer0_outputs(151));
    outputs(9904) <= not(layer0_outputs(7238));
    outputs(9905) <= (layer0_outputs(162)) and not (layer0_outputs(11886));
    outputs(9906) <= layer0_outputs(12675);
    outputs(9907) <= not(layer0_outputs(7020));
    outputs(9908) <= not((layer0_outputs(7533)) xor (layer0_outputs(4048)));
    outputs(9909) <= not((layer0_outputs(1444)) or (layer0_outputs(5048)));
    outputs(9910) <= layer0_outputs(8873);
    outputs(9911) <= (layer0_outputs(6391)) xor (layer0_outputs(2994));
    outputs(9912) <= (layer0_outputs(10633)) xor (layer0_outputs(9002));
    outputs(9913) <= not(layer0_outputs(11192));
    outputs(9914) <= layer0_outputs(9588);
    outputs(9915) <= not((layer0_outputs(5529)) xor (layer0_outputs(9537)));
    outputs(9916) <= not((layer0_outputs(6179)) xor (layer0_outputs(123)));
    outputs(9917) <= (layer0_outputs(8910)) xor (layer0_outputs(189));
    outputs(9918) <= (layer0_outputs(5267)) and (layer0_outputs(8524));
    outputs(9919) <= layer0_outputs(8045);
    outputs(9920) <= layer0_outputs(10083);
    outputs(9921) <= layer0_outputs(5148);
    outputs(9922) <= not((layer0_outputs(4119)) or (layer0_outputs(6721)));
    outputs(9923) <= layer0_outputs(3917);
    outputs(9924) <= not(layer0_outputs(3497));
    outputs(9925) <= not(layer0_outputs(7950));
    outputs(9926) <= layer0_outputs(12696);
    outputs(9927) <= not(layer0_outputs(1732));
    outputs(9928) <= not((layer0_outputs(10908)) or (layer0_outputs(11512)));
    outputs(9929) <= (layer0_outputs(11903)) xor (layer0_outputs(2713));
    outputs(9930) <= not(layer0_outputs(8416));
    outputs(9931) <= (layer0_outputs(4583)) and not (layer0_outputs(9249));
    outputs(9932) <= not((layer0_outputs(7016)) xor (layer0_outputs(9985)));
    outputs(9933) <= layer0_outputs(27);
    outputs(9934) <= (layer0_outputs(9658)) and not (layer0_outputs(2142));
    outputs(9935) <= not((layer0_outputs(10398)) xor (layer0_outputs(6016)));
    outputs(9936) <= not((layer0_outputs(11195)) xor (layer0_outputs(5404)));
    outputs(9937) <= (layer0_outputs(9431)) and not (layer0_outputs(2656));
    outputs(9938) <= (layer0_outputs(9964)) xor (layer0_outputs(7355));
    outputs(9939) <= not(layer0_outputs(2198)) or (layer0_outputs(5222));
    outputs(9940) <= not((layer0_outputs(2676)) xor (layer0_outputs(12642)));
    outputs(9941) <= not(layer0_outputs(12690));
    outputs(9942) <= layer0_outputs(11580);
    outputs(9943) <= not((layer0_outputs(4339)) xor (layer0_outputs(7328)));
    outputs(9944) <= (layer0_outputs(4698)) xor (layer0_outputs(1699));
    outputs(9945) <= not(layer0_outputs(3417));
    outputs(9946) <= (layer0_outputs(2647)) and (layer0_outputs(10552));
    outputs(9947) <= layer0_outputs(4478);
    outputs(9948) <= not((layer0_outputs(12584)) xor (layer0_outputs(484)));
    outputs(9949) <= layer0_outputs(4081);
    outputs(9950) <= not(layer0_outputs(12196)) or (layer0_outputs(3010));
    outputs(9951) <= layer0_outputs(3806);
    outputs(9952) <= not((layer0_outputs(9410)) and (layer0_outputs(9007)));
    outputs(9953) <= layer0_outputs(3547);
    outputs(9954) <= (layer0_outputs(1801)) xor (layer0_outputs(8433));
    outputs(9955) <= not((layer0_outputs(5588)) xor (layer0_outputs(3118)));
    outputs(9956) <= (layer0_outputs(2575)) and not (layer0_outputs(2705));
    outputs(9957) <= (layer0_outputs(2855)) and (layer0_outputs(12117));
    outputs(9958) <= (layer0_outputs(971)) and not (layer0_outputs(1141));
    outputs(9959) <= not(layer0_outputs(2561));
    outputs(9960) <= layer0_outputs(8992);
    outputs(9961) <= (layer0_outputs(6555)) xor (layer0_outputs(1006));
    outputs(9962) <= layer0_outputs(8466);
    outputs(9963) <= layer0_outputs(1001);
    outputs(9964) <= (layer0_outputs(245)) xor (layer0_outputs(10824));
    outputs(9965) <= (layer0_outputs(8552)) xor (layer0_outputs(9689));
    outputs(9966) <= not(layer0_outputs(3587)) or (layer0_outputs(10822));
    outputs(9967) <= not(layer0_outputs(4028));
    outputs(9968) <= not((layer0_outputs(1302)) or (layer0_outputs(7909)));
    outputs(9969) <= not(layer0_outputs(10237));
    outputs(9970) <= layer0_outputs(4174);
    outputs(9971) <= layer0_outputs(4256);
    outputs(9972) <= layer0_outputs(11536);
    outputs(9973) <= (layer0_outputs(1262)) and not (layer0_outputs(8480));
    outputs(9974) <= not(layer0_outputs(7334));
    outputs(9975) <= (layer0_outputs(11738)) and (layer0_outputs(4928));
    outputs(9976) <= not(layer0_outputs(8286));
    outputs(9977) <= not((layer0_outputs(5360)) xor (layer0_outputs(6926)));
    outputs(9978) <= not(layer0_outputs(10247));
    outputs(9979) <= (layer0_outputs(7922)) and not (layer0_outputs(7157));
    outputs(9980) <= not(layer0_outputs(440));
    outputs(9981) <= not((layer0_outputs(2242)) or (layer0_outputs(3082)));
    outputs(9982) <= not(layer0_outputs(5774));
    outputs(9983) <= layer0_outputs(7648);
    outputs(9984) <= not((layer0_outputs(2068)) or (layer0_outputs(6981)));
    outputs(9985) <= (layer0_outputs(9196)) and (layer0_outputs(211));
    outputs(9986) <= not((layer0_outputs(10523)) and (layer0_outputs(11676)));
    outputs(9987) <= (layer0_outputs(874)) and not (layer0_outputs(6267));
    outputs(9988) <= not(layer0_outputs(9437));
    outputs(9989) <= (layer0_outputs(9030)) xor (layer0_outputs(6400));
    outputs(9990) <= layer0_outputs(2593);
    outputs(9991) <= not((layer0_outputs(7614)) xor (layer0_outputs(11178)));
    outputs(9992) <= not(layer0_outputs(510));
    outputs(9993) <= not(layer0_outputs(11077));
    outputs(9994) <= not(layer0_outputs(8998));
    outputs(9995) <= (layer0_outputs(1487)) and (layer0_outputs(1125));
    outputs(9996) <= (layer0_outputs(12796)) xor (layer0_outputs(955));
    outputs(9997) <= (layer0_outputs(218)) or (layer0_outputs(11697));
    outputs(9998) <= not((layer0_outputs(696)) or (layer0_outputs(666)));
    outputs(9999) <= not(layer0_outputs(12355));
    outputs(10000) <= (layer0_outputs(2462)) and not (layer0_outputs(5702));
    outputs(10001) <= layer0_outputs(11604);
    outputs(10002) <= (layer0_outputs(8317)) and not (layer0_outputs(4077));
    outputs(10003) <= layer0_outputs(5017);
    outputs(10004) <= (layer0_outputs(7433)) and not (layer0_outputs(7290));
    outputs(10005) <= not(layer0_outputs(2122));
    outputs(10006) <= (layer0_outputs(1056)) and not (layer0_outputs(9006));
    outputs(10007) <= (layer0_outputs(12392)) and not (layer0_outputs(11524));
    outputs(10008) <= not((layer0_outputs(5637)) xor (layer0_outputs(10984)));
    outputs(10009) <= not(layer0_outputs(11743));
    outputs(10010) <= not(layer0_outputs(9805));
    outputs(10011) <= (layer0_outputs(3997)) and not (layer0_outputs(12103));
    outputs(10012) <= (layer0_outputs(7837)) xor (layer0_outputs(3766));
    outputs(10013) <= (layer0_outputs(10774)) xor (layer0_outputs(2384));
    outputs(10014) <= (layer0_outputs(4795)) and not (layer0_outputs(10741));
    outputs(10015) <= layer0_outputs(6807);
    outputs(10016) <= (layer0_outputs(1874)) and not (layer0_outputs(5970));
    outputs(10017) <= not((layer0_outputs(8667)) xor (layer0_outputs(3005)));
    outputs(10018) <= (layer0_outputs(10354)) xor (layer0_outputs(3014));
    outputs(10019) <= not((layer0_outputs(1295)) or (layer0_outputs(1756)));
    outputs(10020) <= not((layer0_outputs(8616)) xor (layer0_outputs(4496)));
    outputs(10021) <= layer0_outputs(851);
    outputs(10022) <= (layer0_outputs(10647)) and (layer0_outputs(499));
    outputs(10023) <= (layer0_outputs(657)) and not (layer0_outputs(5082));
    outputs(10024) <= not((layer0_outputs(3893)) or (layer0_outputs(8869)));
    outputs(10025) <= not((layer0_outputs(3693)) or (layer0_outputs(5003)));
    outputs(10026) <= (layer0_outputs(204)) xor (layer0_outputs(3489));
    outputs(10027) <= layer0_outputs(9626);
    outputs(10028) <= not((layer0_outputs(7521)) or (layer0_outputs(7084)));
    outputs(10029) <= layer0_outputs(10069);
    outputs(10030) <= (layer0_outputs(12305)) and not (layer0_outputs(11504));
    outputs(10031) <= not((layer0_outputs(877)) xor (layer0_outputs(11210)));
    outputs(10032) <= layer0_outputs(3691);
    outputs(10033) <= (layer0_outputs(6962)) and not (layer0_outputs(3564));
    outputs(10034) <= not((layer0_outputs(7782)) or (layer0_outputs(4824)));
    outputs(10035) <= layer0_outputs(3131);
    outputs(10036) <= (layer0_outputs(11066)) and (layer0_outputs(7691));
    outputs(10037) <= not(layer0_outputs(5359));
    outputs(10038) <= not((layer0_outputs(8364)) xor (layer0_outputs(12468)));
    outputs(10039) <= not(layer0_outputs(8207)) or (layer0_outputs(11812));
    outputs(10040) <= (layer0_outputs(911)) and not (layer0_outputs(12425));
    outputs(10041) <= not(layer0_outputs(4261));
    outputs(10042) <= not(layer0_outputs(2537));
    outputs(10043) <= not((layer0_outputs(7492)) xor (layer0_outputs(9178)));
    outputs(10044) <= (layer0_outputs(4657)) and not (layer0_outputs(5223));
    outputs(10045) <= layer0_outputs(9224);
    outputs(10046) <= not((layer0_outputs(6917)) xor (layer0_outputs(1945)));
    outputs(10047) <= layer0_outputs(11990);
    outputs(10048) <= (layer0_outputs(11400)) xor (layer0_outputs(484));
    outputs(10049) <= not((layer0_outputs(12039)) and (layer0_outputs(8827)));
    outputs(10050) <= not((layer0_outputs(11267)) or (layer0_outputs(7224)));
    outputs(10051) <= (layer0_outputs(5944)) xor (layer0_outputs(8885));
    outputs(10052) <= not((layer0_outputs(1248)) xor (layer0_outputs(7981)));
    outputs(10053) <= not(layer0_outputs(5216));
    outputs(10054) <= layer0_outputs(5722);
    outputs(10055) <= (layer0_outputs(9409)) and not (layer0_outputs(1547));
    outputs(10056) <= layer0_outputs(4321);
    outputs(10057) <= (layer0_outputs(5622)) xor (layer0_outputs(6114));
    outputs(10058) <= layer0_outputs(10988);
    outputs(10059) <= layer0_outputs(6949);
    outputs(10060) <= layer0_outputs(10882);
    outputs(10061) <= layer0_outputs(8490);
    outputs(10062) <= layer0_outputs(8400);
    outputs(10063) <= layer0_outputs(9547);
    outputs(10064) <= not((layer0_outputs(8530)) or (layer0_outputs(7907)));
    outputs(10065) <= layer0_outputs(5247);
    outputs(10066) <= not((layer0_outputs(11234)) or (layer0_outputs(1403)));
    outputs(10067) <= (layer0_outputs(10206)) xor (layer0_outputs(3472));
    outputs(10068) <= (layer0_outputs(7535)) and not (layer0_outputs(5546));
    outputs(10069) <= layer0_outputs(5456);
    outputs(10070) <= layer0_outputs(10619);
    outputs(10071) <= (layer0_outputs(1571)) or (layer0_outputs(345));
    outputs(10072) <= (layer0_outputs(12476)) and not (layer0_outputs(12120));
    outputs(10073) <= not(layer0_outputs(9282));
    outputs(10074) <= layer0_outputs(3140);
    outputs(10075) <= not(layer0_outputs(6059)) or (layer0_outputs(1061));
    outputs(10076) <= layer0_outputs(6115);
    outputs(10077) <= (layer0_outputs(896)) and not (layer0_outputs(6018));
    outputs(10078) <= layer0_outputs(11127);
    outputs(10079) <= layer0_outputs(12107);
    outputs(10080) <= not((layer0_outputs(3258)) xor (layer0_outputs(8839)));
    outputs(10081) <= (layer0_outputs(5828)) and (layer0_outputs(2509));
    outputs(10082) <= not(layer0_outputs(1305));
    outputs(10083) <= (layer0_outputs(7587)) xor (layer0_outputs(11200));
    outputs(10084) <= (layer0_outputs(2571)) xor (layer0_outputs(1695));
    outputs(10085) <= (layer0_outputs(3933)) and (layer0_outputs(9767));
    outputs(10086) <= (layer0_outputs(228)) and not (layer0_outputs(1371));
    outputs(10087) <= not(layer0_outputs(12354));
    outputs(10088) <= not((layer0_outputs(6474)) xor (layer0_outputs(4538)));
    outputs(10089) <= not((layer0_outputs(1038)) xor (layer0_outputs(8546)));
    outputs(10090) <= (layer0_outputs(1852)) and (layer0_outputs(1598));
    outputs(10091) <= layer0_outputs(2107);
    outputs(10092) <= not((layer0_outputs(10018)) xor (layer0_outputs(10968)));
    outputs(10093) <= layer0_outputs(3676);
    outputs(10094) <= layer0_outputs(367);
    outputs(10095) <= (layer0_outputs(12099)) and (layer0_outputs(8157));
    outputs(10096) <= not(layer0_outputs(10902));
    outputs(10097) <= not((layer0_outputs(4588)) or (layer0_outputs(9505)));
    outputs(10098) <= not((layer0_outputs(9680)) xor (layer0_outputs(8502)));
    outputs(10099) <= (layer0_outputs(1725)) xor (layer0_outputs(10985));
    outputs(10100) <= not((layer0_outputs(3726)) or (layer0_outputs(2312)));
    outputs(10101) <= not(layer0_outputs(4747));
    outputs(10102) <= (layer0_outputs(9798)) xor (layer0_outputs(7668));
    outputs(10103) <= layer0_outputs(3571);
    outputs(10104) <= layer0_outputs(6056);
    outputs(10105) <= not((layer0_outputs(11621)) xor (layer0_outputs(10848)));
    outputs(10106) <= layer0_outputs(4943);
    outputs(10107) <= (layer0_outputs(9970)) and not (layer0_outputs(4477));
    outputs(10108) <= (layer0_outputs(9690)) or (layer0_outputs(2461));
    outputs(10109) <= layer0_outputs(12464);
    outputs(10110) <= not(layer0_outputs(12441));
    outputs(10111) <= not(layer0_outputs(6809));
    outputs(10112) <= not(layer0_outputs(3011));
    outputs(10113) <= (layer0_outputs(4647)) and not (layer0_outputs(12092));
    outputs(10114) <= (layer0_outputs(6729)) and (layer0_outputs(2456));
    outputs(10115) <= layer0_outputs(11647);
    outputs(10116) <= not((layer0_outputs(7694)) or (layer0_outputs(4251)));
    outputs(10117) <= (layer0_outputs(5476)) xor (layer0_outputs(9438));
    outputs(10118) <= layer0_outputs(642);
    outputs(10119) <= (layer0_outputs(8260)) xor (layer0_outputs(11602));
    outputs(10120) <= (layer0_outputs(3999)) xor (layer0_outputs(5929));
    outputs(10121) <= (layer0_outputs(6651)) xor (layer0_outputs(10802));
    outputs(10122) <= layer0_outputs(3304);
    outputs(10123) <= not((layer0_outputs(10755)) xor (layer0_outputs(11696)));
    outputs(10124) <= not((layer0_outputs(7566)) or (layer0_outputs(9420)));
    outputs(10125) <= layer0_outputs(1892);
    outputs(10126) <= not((layer0_outputs(9266)) xor (layer0_outputs(4988)));
    outputs(10127) <= not(layer0_outputs(4980));
    outputs(10128) <= not(layer0_outputs(7430));
    outputs(10129) <= not(layer0_outputs(3878));
    outputs(10130) <= layer0_outputs(10420);
    outputs(10131) <= layer0_outputs(6251);
    outputs(10132) <= (layer0_outputs(334)) and not (layer0_outputs(446));
    outputs(10133) <= (layer0_outputs(9501)) and (layer0_outputs(11281));
    outputs(10134) <= (layer0_outputs(12223)) xor (layer0_outputs(9546));
    outputs(10135) <= not((layer0_outputs(2867)) xor (layer0_outputs(11970)));
    outputs(10136) <= (layer0_outputs(11441)) and not (layer0_outputs(4862));
    outputs(10137) <= layer0_outputs(218);
    outputs(10138) <= layer0_outputs(10541);
    outputs(10139) <= not((layer0_outputs(7554)) or (layer0_outputs(10145)));
    outputs(10140) <= (layer0_outputs(7569)) and (layer0_outputs(4107));
    outputs(10141) <= layer0_outputs(2472);
    outputs(10142) <= layer0_outputs(3004);
    outputs(10143) <= layer0_outputs(7164);
    outputs(10144) <= not(layer0_outputs(8843));
    outputs(10145) <= (layer0_outputs(12723)) and not (layer0_outputs(2634));
    outputs(10146) <= not((layer0_outputs(5106)) or (layer0_outputs(78)));
    outputs(10147) <= (layer0_outputs(3367)) and not (layer0_outputs(8712));
    outputs(10148) <= (layer0_outputs(6260)) xor (layer0_outputs(8960));
    outputs(10149) <= layer0_outputs(11194);
    outputs(10150) <= not(layer0_outputs(7479));
    outputs(10151) <= not((layer0_outputs(11625)) or (layer0_outputs(10710)));
    outputs(10152) <= (layer0_outputs(9745)) and not (layer0_outputs(3438));
    outputs(10153) <= layer0_outputs(6926);
    outputs(10154) <= not(layer0_outputs(11628));
    outputs(10155) <= layer0_outputs(11680);
    outputs(10156) <= not(layer0_outputs(2761));
    outputs(10157) <= not(layer0_outputs(12402)) or (layer0_outputs(963));
    outputs(10158) <= layer0_outputs(9764);
    outputs(10159) <= not(layer0_outputs(9904));
    outputs(10160) <= not(layer0_outputs(10894));
    outputs(10161) <= layer0_outputs(12352);
    outputs(10162) <= not(layer0_outputs(9294));
    outputs(10163) <= (layer0_outputs(11551)) xor (layer0_outputs(12341));
    outputs(10164) <= (layer0_outputs(6363)) or (layer0_outputs(6772));
    outputs(10165) <= (layer0_outputs(9858)) xor (layer0_outputs(5184));
    outputs(10166) <= layer0_outputs(9594);
    outputs(10167) <= (layer0_outputs(559)) xor (layer0_outputs(7252));
    outputs(10168) <= not((layer0_outputs(5655)) or (layer0_outputs(8496)));
    outputs(10169) <= not((layer0_outputs(9752)) or (layer0_outputs(2302)));
    outputs(10170) <= (layer0_outputs(4113)) xor (layer0_outputs(9591));
    outputs(10171) <= not((layer0_outputs(3401)) xor (layer0_outputs(6187)));
    outputs(10172) <= not(layer0_outputs(1493));
    outputs(10173) <= (layer0_outputs(2602)) xor (layer0_outputs(11380));
    outputs(10174) <= not(layer0_outputs(9385)) or (layer0_outputs(2235));
    outputs(10175) <= not(layer0_outputs(2370));
    outputs(10176) <= not(layer0_outputs(3211));
    outputs(10177) <= not((layer0_outputs(6743)) xor (layer0_outputs(3059)));
    outputs(10178) <= (layer0_outputs(5782)) xor (layer0_outputs(10390));
    outputs(10179) <= (layer0_outputs(11946)) and not (layer0_outputs(11024));
    outputs(10180) <= layer0_outputs(1620);
    outputs(10181) <= not((layer0_outputs(10143)) or (layer0_outputs(4771)));
    outputs(10182) <= layer0_outputs(6392);
    outputs(10183) <= not(layer0_outputs(612));
    outputs(10184) <= (layer0_outputs(8899)) or (layer0_outputs(231));
    outputs(10185) <= not(layer0_outputs(539));
    outputs(10186) <= (layer0_outputs(3795)) and not (layer0_outputs(4736));
    outputs(10187) <= not(layer0_outputs(6162));
    outputs(10188) <= (layer0_outputs(9562)) and (layer0_outputs(11407));
    outputs(10189) <= not(layer0_outputs(7475));
    outputs(10190) <= (layer0_outputs(11351)) and not (layer0_outputs(7454));
    outputs(10191) <= not(layer0_outputs(4683));
    outputs(10192) <= (layer0_outputs(12275)) and not (layer0_outputs(2716));
    outputs(10193) <= layer0_outputs(3373);
    outputs(10194) <= (layer0_outputs(9517)) and not (layer0_outputs(2533));
    outputs(10195) <= (layer0_outputs(2234)) and not (layer0_outputs(8048));
    outputs(10196) <= not(layer0_outputs(5074));
    outputs(10197) <= (layer0_outputs(3943)) xor (layer0_outputs(1203));
    outputs(10198) <= not(layer0_outputs(11991));
    outputs(10199) <= (layer0_outputs(7245)) and not (layer0_outputs(605));
    outputs(10200) <= not((layer0_outputs(130)) or (layer0_outputs(9026)));
    outputs(10201) <= layer0_outputs(3710);
    outputs(10202) <= not(layer0_outputs(6968));
    outputs(10203) <= layer0_outputs(9633);
    outputs(10204) <= not(layer0_outputs(8105));
    outputs(10205) <= (layer0_outputs(8110)) and not (layer0_outputs(9848));
    outputs(10206) <= (layer0_outputs(738)) xor (layer0_outputs(9136));
    outputs(10207) <= layer0_outputs(5432);
    outputs(10208) <= (layer0_outputs(573)) xor (layer0_outputs(4804));
    outputs(10209) <= (layer0_outputs(5612)) and (layer0_outputs(6259));
    outputs(10210) <= (layer0_outputs(4722)) and not (layer0_outputs(2673));
    outputs(10211) <= not((layer0_outputs(1963)) or (layer0_outputs(10488)));
    outputs(10212) <= not(layer0_outputs(155));
    outputs(10213) <= not(layer0_outputs(1275));
    outputs(10214) <= layer0_outputs(2711);
    outputs(10215) <= not((layer0_outputs(3704)) or (layer0_outputs(11867)));
    outputs(10216) <= not((layer0_outputs(5280)) xor (layer0_outputs(7737)));
    outputs(10217) <= not((layer0_outputs(3186)) xor (layer0_outputs(11090)));
    outputs(10218) <= not(layer0_outputs(11862));
    outputs(10219) <= layer0_outputs(3790);
    outputs(10220) <= layer0_outputs(11063);
    outputs(10221) <= (layer0_outputs(7653)) xor (layer0_outputs(4237));
    outputs(10222) <= (layer0_outputs(5676)) xor (layer0_outputs(5581));
    outputs(10223) <= layer0_outputs(10370);
    outputs(10224) <= not((layer0_outputs(6530)) or (layer0_outputs(4648)));
    outputs(10225) <= layer0_outputs(18);
    outputs(10226) <= layer0_outputs(1017);
    outputs(10227) <= layer0_outputs(8781);
    outputs(10228) <= not((layer0_outputs(8185)) or (layer0_outputs(1984)));
    outputs(10229) <= not((layer0_outputs(8555)) xor (layer0_outputs(6965)));
    outputs(10230) <= layer0_outputs(9814);
    outputs(10231) <= (layer0_outputs(6734)) and not (layer0_outputs(12704));
    outputs(10232) <= not((layer0_outputs(3802)) xor (layer0_outputs(4192)));
    outputs(10233) <= (layer0_outputs(8068)) xor (layer0_outputs(4308));
    outputs(10234) <= not((layer0_outputs(2209)) or (layer0_outputs(2024)));
    outputs(10235) <= not(layer0_outputs(10137)) or (layer0_outputs(7970));
    outputs(10236) <= not((layer0_outputs(9516)) xor (layer0_outputs(1749)));
    outputs(10237) <= (layer0_outputs(11569)) xor (layer0_outputs(625));
    outputs(10238) <= (layer0_outputs(1211)) and (layer0_outputs(5455));
    outputs(10239) <= not(layer0_outputs(1767));
    outputs(10240) <= (layer0_outputs(643)) and (layer0_outputs(10067));
    outputs(10241) <= not(layer0_outputs(6647));
    outputs(10242) <= (layer0_outputs(9711)) xor (layer0_outputs(3868));
    outputs(10243) <= (layer0_outputs(10832)) and not (layer0_outputs(3879));
    outputs(10244) <= (layer0_outputs(6637)) or (layer0_outputs(7226));
    outputs(10245) <= layer0_outputs(3871);
    outputs(10246) <= not(layer0_outputs(601));
    outputs(10247) <= not(layer0_outputs(9562));
    outputs(10248) <= '1';
    outputs(10249) <= not((layer0_outputs(7574)) xor (layer0_outputs(11626)));
    outputs(10250) <= (layer0_outputs(11413)) xor (layer0_outputs(11944));
    outputs(10251) <= layer0_outputs(1624);
    outputs(10252) <= (layer0_outputs(3297)) and not (layer0_outputs(12101));
    outputs(10253) <= (layer0_outputs(6980)) xor (layer0_outputs(10944));
    outputs(10254) <= (layer0_outputs(3898)) xor (layer0_outputs(7629));
    outputs(10255) <= layer0_outputs(5366);
    outputs(10256) <= layer0_outputs(7698);
    outputs(10257) <= not(layer0_outputs(3070)) or (layer0_outputs(8095));
    outputs(10258) <= not((layer0_outputs(1150)) xor (layer0_outputs(6775)));
    outputs(10259) <= not(layer0_outputs(2091)) or (layer0_outputs(10005));
    outputs(10260) <= layer0_outputs(3585);
    outputs(10261) <= not(layer0_outputs(12516));
    outputs(10262) <= not(layer0_outputs(11873));
    outputs(10263) <= (layer0_outputs(3106)) and not (layer0_outputs(9564));
    outputs(10264) <= not(layer0_outputs(126)) or (layer0_outputs(7475));
    outputs(10265) <= (layer0_outputs(1922)) and (layer0_outputs(1910));
    outputs(10266) <= not(layer0_outputs(12213)) or (layer0_outputs(11509));
    outputs(10267) <= layer0_outputs(10126);
    outputs(10268) <= layer0_outputs(6743);
    outputs(10269) <= not((layer0_outputs(10117)) and (layer0_outputs(7918)));
    outputs(10270) <= (layer0_outputs(3552)) or (layer0_outputs(8221));
    outputs(10271) <= (layer0_outputs(7603)) or (layer0_outputs(7570));
    outputs(10272) <= not(layer0_outputs(12291));
    outputs(10273) <= not(layer0_outputs(3462));
    outputs(10274) <= not(layer0_outputs(3371));
    outputs(10275) <= layer0_outputs(3173);
    outputs(10276) <= not((layer0_outputs(8804)) xor (layer0_outputs(11133)));
    outputs(10277) <= not(layer0_outputs(5250)) or (layer0_outputs(1007));
    outputs(10278) <= layer0_outputs(9890);
    outputs(10279) <= not(layer0_outputs(7723));
    outputs(10280) <= layer0_outputs(9394);
    outputs(10281) <= not((layer0_outputs(6268)) and (layer0_outputs(5049)));
    outputs(10282) <= not(layer0_outputs(4788));
    outputs(10283) <= (layer0_outputs(9321)) or (layer0_outputs(12738));
    outputs(10284) <= not((layer0_outputs(11801)) and (layer0_outputs(538)));
    outputs(10285) <= not(layer0_outputs(8860));
    outputs(10286) <= (layer0_outputs(1062)) xor (layer0_outputs(655));
    outputs(10287) <= layer0_outputs(9913);
    outputs(10288) <= not((layer0_outputs(9971)) xor (layer0_outputs(4684)));
    outputs(10289) <= not(layer0_outputs(7326));
    outputs(10290) <= not((layer0_outputs(6232)) xor (layer0_outputs(1629)));
    outputs(10291) <= not(layer0_outputs(11395));
    outputs(10292) <= not(layer0_outputs(1515)) or (layer0_outputs(10850));
    outputs(10293) <= not((layer0_outputs(1575)) xor (layer0_outputs(5705)));
    outputs(10294) <= not(layer0_outputs(4172));
    outputs(10295) <= not(layer0_outputs(7982));
    outputs(10296) <= (layer0_outputs(11349)) or (layer0_outputs(1966));
    outputs(10297) <= (layer0_outputs(738)) and not (layer0_outputs(6670));
    outputs(10298) <= (layer0_outputs(12514)) xor (layer0_outputs(2539));
    outputs(10299) <= layer0_outputs(4149);
    outputs(10300) <= not((layer0_outputs(1354)) xor (layer0_outputs(10681)));
    outputs(10301) <= not((layer0_outputs(6502)) and (layer0_outputs(4431)));
    outputs(10302) <= not(layer0_outputs(10040)) or (layer0_outputs(3612));
    outputs(10303) <= not((layer0_outputs(9061)) xor (layer0_outputs(11086)));
    outputs(10304) <= not((layer0_outputs(7552)) xor (layer0_outputs(7014)));
    outputs(10305) <= not(layer0_outputs(3733));
    outputs(10306) <= not((layer0_outputs(6989)) xor (layer0_outputs(4188)));
    outputs(10307) <= not(layer0_outputs(6878));
    outputs(10308) <= layer0_outputs(2303);
    outputs(10309) <= not((layer0_outputs(7468)) or (layer0_outputs(12171)));
    outputs(10310) <= (layer0_outputs(494)) and not (layer0_outputs(11894));
    outputs(10311) <= (layer0_outputs(2724)) xor (layer0_outputs(10725));
    outputs(10312) <= (layer0_outputs(11942)) xor (layer0_outputs(10764));
    outputs(10313) <= not(layer0_outputs(10780));
    outputs(10314) <= not((layer0_outputs(12450)) and (layer0_outputs(4865)));
    outputs(10315) <= layer0_outputs(8907);
    outputs(10316) <= not(layer0_outputs(501));
    outputs(10317) <= (layer0_outputs(5654)) or (layer0_outputs(8218));
    outputs(10318) <= not((layer0_outputs(475)) xor (layer0_outputs(8867)));
    outputs(10319) <= not(layer0_outputs(6748)) or (layer0_outputs(10726));
    outputs(10320) <= layer0_outputs(235);
    outputs(10321) <= not((layer0_outputs(5235)) xor (layer0_outputs(6403)));
    outputs(10322) <= not((layer0_outputs(2047)) xor (layer0_outputs(11402)));
    outputs(10323) <= not((layer0_outputs(4887)) or (layer0_outputs(9415)));
    outputs(10324) <= not(layer0_outputs(10147));
    outputs(10325) <= not((layer0_outputs(7900)) or (layer0_outputs(5040)));
    outputs(10326) <= (layer0_outputs(10611)) or (layer0_outputs(4340));
    outputs(10327) <= not(layer0_outputs(7278));
    outputs(10328) <= (layer0_outputs(9168)) and not (layer0_outputs(873));
    outputs(10329) <= layer0_outputs(10908);
    outputs(10330) <= not(layer0_outputs(4296));
    outputs(10331) <= not((layer0_outputs(1788)) xor (layer0_outputs(2081)));
    outputs(10332) <= not((layer0_outputs(3439)) xor (layer0_outputs(8615)));
    outputs(10333) <= not(layer0_outputs(5142)) or (layer0_outputs(11620));
    outputs(10334) <= not((layer0_outputs(638)) xor (layer0_outputs(857)));
    outputs(10335) <= not(layer0_outputs(11481));
    outputs(10336) <= not(layer0_outputs(10644));
    outputs(10337) <= layer0_outputs(7820);
    outputs(10338) <= not((layer0_outputs(11225)) xor (layer0_outputs(6680)));
    outputs(10339) <= layer0_outputs(8193);
    outputs(10340) <= layer0_outputs(12167);
    outputs(10341) <= layer0_outputs(5020);
    outputs(10342) <= not((layer0_outputs(4490)) xor (layer0_outputs(5709)));
    outputs(10343) <= not(layer0_outputs(10830));
    outputs(10344) <= (layer0_outputs(11007)) and not (layer0_outputs(1848));
    outputs(10345) <= (layer0_outputs(2101)) xor (layer0_outputs(8932));
    outputs(10346) <= not((layer0_outputs(9469)) xor (layer0_outputs(9298)));
    outputs(10347) <= (layer0_outputs(11494)) xor (layer0_outputs(1258));
    outputs(10348) <= (layer0_outputs(3387)) or (layer0_outputs(8225));
    outputs(10349) <= not((layer0_outputs(1493)) xor (layer0_outputs(9982)));
    outputs(10350) <= not((layer0_outputs(3392)) xor (layer0_outputs(2139)));
    outputs(10351) <= (layer0_outputs(10686)) or (layer0_outputs(12102));
    outputs(10352) <= not((layer0_outputs(5944)) xor (layer0_outputs(7864)));
    outputs(10353) <= layer0_outputs(3280);
    outputs(10354) <= (layer0_outputs(10601)) xor (layer0_outputs(1237));
    outputs(10355) <= not(layer0_outputs(10537));
    outputs(10356) <= not((layer0_outputs(4384)) xor (layer0_outputs(11371)));
    outputs(10357) <= not(layer0_outputs(10442));
    outputs(10358) <= layer0_outputs(272);
    outputs(10359) <= not(layer0_outputs(1312)) or (layer0_outputs(1240));
    outputs(10360) <= (layer0_outputs(2481)) xor (layer0_outputs(8592));
    outputs(10361) <= not((layer0_outputs(7559)) and (layer0_outputs(9727)));
    outputs(10362) <= not(layer0_outputs(7119));
    outputs(10363) <= not(layer0_outputs(1237)) or (layer0_outputs(10263));
    outputs(10364) <= (layer0_outputs(10028)) or (layer0_outputs(4947));
    outputs(10365) <= (layer0_outputs(10678)) xor (layer0_outputs(9358));
    outputs(10366) <= not((layer0_outputs(9492)) and (layer0_outputs(5791)));
    outputs(10367) <= not(layer0_outputs(7944)) or (layer0_outputs(5814));
    outputs(10368) <= (layer0_outputs(10653)) xor (layer0_outputs(866));
    outputs(10369) <= (layer0_outputs(312)) xor (layer0_outputs(3714));
    outputs(10370) <= not(layer0_outputs(7680));
    outputs(10371) <= not((layer0_outputs(2327)) xor (layer0_outputs(2595)));
    outputs(10372) <= (layer0_outputs(142)) xor (layer0_outputs(3707));
    outputs(10373) <= not((layer0_outputs(4241)) and (layer0_outputs(7469)));
    outputs(10374) <= not(layer0_outputs(4780));
    outputs(10375) <= layer0_outputs(10299);
    outputs(10376) <= not(layer0_outputs(1658));
    outputs(10377) <= not(layer0_outputs(6150)) or (layer0_outputs(5673));
    outputs(10378) <= not(layer0_outputs(9362));
    outputs(10379) <= (layer0_outputs(5501)) xor (layer0_outputs(11656));
    outputs(10380) <= not((layer0_outputs(4482)) xor (layer0_outputs(346)));
    outputs(10381) <= not(layer0_outputs(8087));
    outputs(10382) <= layer0_outputs(8737);
    outputs(10383) <= layer0_outputs(4127);
    outputs(10384) <= not(layer0_outputs(6388));
    outputs(10385) <= not((layer0_outputs(4408)) and (layer0_outputs(11141)));
    outputs(10386) <= (layer0_outputs(7989)) xor (layer0_outputs(243));
    outputs(10387) <= not(layer0_outputs(8045)) or (layer0_outputs(4435));
    outputs(10388) <= not((layer0_outputs(5899)) xor (layer0_outputs(7350)));
    outputs(10389) <= not(layer0_outputs(755)) or (layer0_outputs(11341));
    outputs(10390) <= layer0_outputs(10940);
    outputs(10391) <= not((layer0_outputs(8408)) or (layer0_outputs(7983)));
    outputs(10392) <= (layer0_outputs(7543)) and (layer0_outputs(3740));
    outputs(10393) <= not((layer0_outputs(6227)) or (layer0_outputs(279)));
    outputs(10394) <= not(layer0_outputs(3244));
    outputs(10395) <= not((layer0_outputs(2706)) xor (layer0_outputs(11604)));
    outputs(10396) <= not(layer0_outputs(6975)) or (layer0_outputs(10419));
    outputs(10397) <= (layer0_outputs(1375)) and not (layer0_outputs(8191));
    outputs(10398) <= (layer0_outputs(7498)) or (layer0_outputs(236));
    outputs(10399) <= not(layer0_outputs(12555));
    outputs(10400) <= layer0_outputs(739);
    outputs(10401) <= not(layer0_outputs(1699)) or (layer0_outputs(2678));
    outputs(10402) <= layer0_outputs(9133);
    outputs(10403) <= not(layer0_outputs(1327));
    outputs(10404) <= (layer0_outputs(3119)) xor (layer0_outputs(10435));
    outputs(10405) <= not(layer0_outputs(601));
    outputs(10406) <= (layer0_outputs(2468)) xor (layer0_outputs(5011));
    outputs(10407) <= not(layer0_outputs(10009)) or (layer0_outputs(2167));
    outputs(10408) <= not(layer0_outputs(1021)) or (layer0_outputs(5332));
    outputs(10409) <= layer0_outputs(1971);
    outputs(10410) <= (layer0_outputs(9038)) or (layer0_outputs(8693));
    outputs(10411) <= (layer0_outputs(807)) xor (layer0_outputs(9190));
    outputs(10412) <= (layer0_outputs(7658)) and not (layer0_outputs(483));
    outputs(10413) <= layer0_outputs(6710);
    outputs(10414) <= not(layer0_outputs(10776)) or (layer0_outputs(6405));
    outputs(10415) <= not(layer0_outputs(9493)) or (layer0_outputs(528));
    outputs(10416) <= (layer0_outputs(7310)) xor (layer0_outputs(5090));
    outputs(10417) <= not(layer0_outputs(7744));
    outputs(10418) <= not((layer0_outputs(3657)) xor (layer0_outputs(8325)));
    outputs(10419) <= not(layer0_outputs(2554));
    outputs(10420) <= not((layer0_outputs(5846)) xor (layer0_outputs(11119)));
    outputs(10421) <= (layer0_outputs(6384)) xor (layer0_outputs(701));
    outputs(10422) <= not((layer0_outputs(10146)) xor (layer0_outputs(1198)));
    outputs(10423) <= not(layer0_outputs(4812)) or (layer0_outputs(2011));
    outputs(10424) <= layer0_outputs(1352);
    outputs(10425) <= not((layer0_outputs(6755)) or (layer0_outputs(2045)));
    outputs(10426) <= layer0_outputs(1276);
    outputs(10427) <= not((layer0_outputs(6700)) xor (layer0_outputs(9844)));
    outputs(10428) <= layer0_outputs(2043);
    outputs(10429) <= not(layer0_outputs(10365)) or (layer0_outputs(7882));
    outputs(10430) <= layer0_outputs(7990);
    outputs(10431) <= layer0_outputs(11896);
    outputs(10432) <= not(layer0_outputs(8524));
    outputs(10433) <= not((layer0_outputs(9255)) or (layer0_outputs(7462)));
    outputs(10434) <= not((layer0_outputs(6281)) xor (layer0_outputs(12695)));
    outputs(10435) <= not(layer0_outputs(8628));
    outputs(10436) <= layer0_outputs(7681);
    outputs(10437) <= (layer0_outputs(10195)) xor (layer0_outputs(9993));
    outputs(10438) <= not((layer0_outputs(4711)) and (layer0_outputs(136)));
    outputs(10439) <= not(layer0_outputs(12406));
    outputs(10440) <= layer0_outputs(1641);
    outputs(10441) <= (layer0_outputs(2097)) or (layer0_outputs(6273));
    outputs(10442) <= not((layer0_outputs(3931)) xor (layer0_outputs(3657)));
    outputs(10443) <= not((layer0_outputs(418)) xor (layer0_outputs(2311)));
    outputs(10444) <= not((layer0_outputs(2064)) xor (layer0_outputs(10881)));
    outputs(10445) <= layer0_outputs(428);
    outputs(10446) <= not(layer0_outputs(2956));
    outputs(10447) <= not(layer0_outputs(9637));
    outputs(10448) <= layer0_outputs(585);
    outputs(10449) <= not((layer0_outputs(4067)) and (layer0_outputs(5601)));
    outputs(10450) <= not(layer0_outputs(10205)) or (layer0_outputs(3847));
    outputs(10451) <= layer0_outputs(294);
    outputs(10452) <= not((layer0_outputs(12594)) xor (layer0_outputs(8486)));
    outputs(10453) <= not((layer0_outputs(5318)) xor (layer0_outputs(12126)));
    outputs(10454) <= (layer0_outputs(4621)) and not (layer0_outputs(4996));
    outputs(10455) <= (layer0_outputs(11231)) xor (layer0_outputs(3944));
    outputs(10456) <= layer0_outputs(12217);
    outputs(10457) <= not(layer0_outputs(10924));
    outputs(10458) <= not((layer0_outputs(9525)) xor (layer0_outputs(986)));
    outputs(10459) <= not(layer0_outputs(9573));
    outputs(10460) <= not(layer0_outputs(9069)) or (layer0_outputs(4699));
    outputs(10461) <= not(layer0_outputs(3769)) or (layer0_outputs(1420));
    outputs(10462) <= not(layer0_outputs(6140));
    outputs(10463) <= not(layer0_outputs(10498)) or (layer0_outputs(2849));
    outputs(10464) <= not(layer0_outputs(5083)) or (layer0_outputs(10852));
    outputs(10465) <= not(layer0_outputs(91)) or (layer0_outputs(4473));
    outputs(10466) <= not(layer0_outputs(8599)) or (layer0_outputs(12303));
    outputs(10467) <= not(layer0_outputs(5044)) or (layer0_outputs(1162));
    outputs(10468) <= not(layer0_outputs(1294)) or (layer0_outputs(4366));
    outputs(10469) <= not((layer0_outputs(654)) and (layer0_outputs(4193)));
    outputs(10470) <= not((layer0_outputs(8814)) xor (layer0_outputs(11353)));
    outputs(10471) <= not(layer0_outputs(2664));
    outputs(10472) <= layer0_outputs(9521);
    outputs(10473) <= (layer0_outputs(4376)) xor (layer0_outputs(10923));
    outputs(10474) <= not(layer0_outputs(5748)) or (layer0_outputs(12509));
    outputs(10475) <= not(layer0_outputs(10305));
    outputs(10476) <= (layer0_outputs(12698)) or (layer0_outputs(432));
    outputs(10477) <= (layer0_outputs(4262)) and (layer0_outputs(11452));
    outputs(10478) <= not((layer0_outputs(11121)) xor (layer0_outputs(8120)));
    outputs(10479) <= not((layer0_outputs(9503)) and (layer0_outputs(142)));
    outputs(10480) <= (layer0_outputs(10808)) xor (layer0_outputs(7168));
    outputs(10481) <= not((layer0_outputs(219)) xor (layer0_outputs(3343)));
    outputs(10482) <= (layer0_outputs(3816)) or (layer0_outputs(9896));
    outputs(10483) <= not(layer0_outputs(10296));
    outputs(10484) <= layer0_outputs(7130);
    outputs(10485) <= layer0_outputs(1799);
    outputs(10486) <= (layer0_outputs(252)) xor (layer0_outputs(5869));
    outputs(10487) <= (layer0_outputs(9811)) xor (layer0_outputs(2264));
    outputs(10488) <= not((layer0_outputs(6655)) xor (layer0_outputs(6598)));
    outputs(10489) <= not(layer0_outputs(6076));
    outputs(10490) <= not(layer0_outputs(7220));
    outputs(10491) <= layer0_outputs(11047);
    outputs(10492) <= (layer0_outputs(2217)) xor (layer0_outputs(1407));
    outputs(10493) <= not((layer0_outputs(12201)) and (layer0_outputs(11396)));
    outputs(10494) <= (layer0_outputs(7699)) or (layer0_outputs(6778));
    outputs(10495) <= layer0_outputs(254);
    outputs(10496) <= (layer0_outputs(9210)) xor (layer0_outputs(6016));
    outputs(10497) <= not((layer0_outputs(7636)) and (layer0_outputs(12193)));
    outputs(10498) <= not((layer0_outputs(9151)) or (layer0_outputs(12512)));
    outputs(10499) <= not(layer0_outputs(5816)) or (layer0_outputs(10905));
    outputs(10500) <= not((layer0_outputs(9041)) xor (layer0_outputs(5210)));
    outputs(10501) <= (layer0_outputs(11041)) xor (layer0_outputs(9711));
    outputs(10502) <= (layer0_outputs(967)) xor (layer0_outputs(8725));
    outputs(10503) <= layer0_outputs(4571);
    outputs(10504) <= (layer0_outputs(11757)) xor (layer0_outputs(5977));
    outputs(10505) <= (layer0_outputs(10527)) xor (layer0_outputs(3728));
    outputs(10506) <= not(layer0_outputs(5058)) or (layer0_outputs(11957));
    outputs(10507) <= not((layer0_outputs(1331)) xor (layer0_outputs(8743)));
    outputs(10508) <= not(layer0_outputs(656));
    outputs(10509) <= (layer0_outputs(7999)) and (layer0_outputs(7405));
    outputs(10510) <= not(layer0_outputs(346));
    outputs(10511) <= not(layer0_outputs(8311));
    outputs(10512) <= (layer0_outputs(9983)) xor (layer0_outputs(1953));
    outputs(10513) <= (layer0_outputs(4710)) xor (layer0_outputs(7755));
    outputs(10514) <= not(layer0_outputs(10251)) or (layer0_outputs(10823));
    outputs(10515) <= not((layer0_outputs(11506)) and (layer0_outputs(4564)));
    outputs(10516) <= not(layer0_outputs(875));
    outputs(10517) <= not((layer0_outputs(7545)) xor (layer0_outputs(5696)));
    outputs(10518) <= (layer0_outputs(81)) or (layer0_outputs(4587));
    outputs(10519) <= not(layer0_outputs(12365));
    outputs(10520) <= layer0_outputs(8399);
    outputs(10521) <= (layer0_outputs(8006)) xor (layer0_outputs(8140));
    outputs(10522) <= layer0_outputs(12328);
    outputs(10523) <= not(layer0_outputs(9093));
    outputs(10524) <= not(layer0_outputs(661));
    outputs(10525) <= (layer0_outputs(3966)) or (layer0_outputs(7271));
    outputs(10526) <= (layer0_outputs(2446)) xor (layer0_outputs(4614));
    outputs(10527) <= not((layer0_outputs(2199)) and (layer0_outputs(3054)));
    outputs(10528) <= not(layer0_outputs(7759)) or (layer0_outputs(6937));
    outputs(10529) <= not(layer0_outputs(1389)) or (layer0_outputs(421));
    outputs(10530) <= not(layer0_outputs(11732)) or (layer0_outputs(10250));
    outputs(10531) <= not(layer0_outputs(10758));
    outputs(10532) <= not((layer0_outputs(3187)) xor (layer0_outputs(7554)));
    outputs(10533) <= not((layer0_outputs(9800)) xor (layer0_outputs(10903)));
    outputs(10534) <= layer0_outputs(9515);
    outputs(10535) <= (layer0_outputs(5151)) xor (layer0_outputs(11618));
    outputs(10536) <= not(layer0_outputs(6954));
    outputs(10537) <= not((layer0_outputs(11544)) xor (layer0_outputs(6995)));
    outputs(10538) <= (layer0_outputs(9894)) xor (layer0_outputs(9442));
    outputs(10539) <= (layer0_outputs(3297)) and (layer0_outputs(3633));
    outputs(10540) <= not((layer0_outputs(1687)) xor (layer0_outputs(7523)));
    outputs(10541) <= layer0_outputs(3126);
    outputs(10542) <= not((layer0_outputs(1051)) xor (layer0_outputs(7334)));
    outputs(10543) <= not((layer0_outputs(5669)) and (layer0_outputs(9063)));
    outputs(10544) <= not((layer0_outputs(1212)) xor (layer0_outputs(7850)));
    outputs(10545) <= not(layer0_outputs(2744)) or (layer0_outputs(2159));
    outputs(10546) <= (layer0_outputs(7997)) xor (layer0_outputs(8980));
    outputs(10547) <= (layer0_outputs(9325)) xor (layer0_outputs(9676));
    outputs(10548) <= not((layer0_outputs(9084)) and (layer0_outputs(6944)));
    outputs(10549) <= not(layer0_outputs(3596));
    outputs(10550) <= not((layer0_outputs(8424)) xor (layer0_outputs(9842)));
    outputs(10551) <= not(layer0_outputs(92)) or (layer0_outputs(11336));
    outputs(10552) <= not((layer0_outputs(12588)) xor (layer0_outputs(10193)));
    outputs(10553) <= not((layer0_outputs(5421)) xor (layer0_outputs(7897)));
    outputs(10554) <= not(layer0_outputs(854)) or (layer0_outputs(2150));
    outputs(10555) <= not((layer0_outputs(8454)) and (layer0_outputs(9625)));
    outputs(10556) <= layer0_outputs(7401);
    outputs(10557) <= not(layer0_outputs(7080));
    outputs(10558) <= (layer0_outputs(4000)) xor (layer0_outputs(11174));
    outputs(10559) <= (layer0_outputs(12550)) xor (layer0_outputs(6221));
    outputs(10560) <= not((layer0_outputs(1588)) xor (layer0_outputs(6916)));
    outputs(10561) <= (layer0_outputs(2360)) xor (layer0_outputs(3817));
    outputs(10562) <= not(layer0_outputs(6515));
    outputs(10563) <= (layer0_outputs(11634)) xor (layer0_outputs(6566));
    outputs(10564) <= not(layer0_outputs(12174));
    outputs(10565) <= not((layer0_outputs(12659)) xor (layer0_outputs(3068)));
    outputs(10566) <= not((layer0_outputs(4570)) xor (layer0_outputs(11085)));
    outputs(10567) <= (layer0_outputs(8371)) and not (layer0_outputs(4212));
    outputs(10568) <= layer0_outputs(7778);
    outputs(10569) <= not(layer0_outputs(496)) or (layer0_outputs(11393));
    outputs(10570) <= not((layer0_outputs(11187)) xor (layer0_outputs(2993)));
    outputs(10571) <= not(layer0_outputs(5334));
    outputs(10572) <= not(layer0_outputs(2131));
    outputs(10573) <= (layer0_outputs(524)) xor (layer0_outputs(6433));
    outputs(10574) <= (layer0_outputs(7801)) xor (layer0_outputs(4509));
    outputs(10575) <= layer0_outputs(4902);
    outputs(10576) <= (layer0_outputs(4679)) or (layer0_outputs(6676));
    outputs(10577) <= not(layer0_outputs(3592)) or (layer0_outputs(11879));
    outputs(10578) <= (layer0_outputs(1149)) xor (layer0_outputs(11225));
    outputs(10579) <= (layer0_outputs(7197)) or (layer0_outputs(648));
    outputs(10580) <= not(layer0_outputs(6978)) or (layer0_outputs(10692));
    outputs(10581) <= not(layer0_outputs(7767)) or (layer0_outputs(7208));
    outputs(10582) <= layer0_outputs(5900);
    outputs(10583) <= not(layer0_outputs(5145));
    outputs(10584) <= not((layer0_outputs(12189)) xor (layer0_outputs(205)));
    outputs(10585) <= not((layer0_outputs(7587)) and (layer0_outputs(1213)));
    outputs(10586) <= not((layer0_outputs(7209)) and (layer0_outputs(757)));
    outputs(10587) <= layer0_outputs(4703);
    outputs(10588) <= (layer0_outputs(2526)) or (layer0_outputs(12736));
    outputs(10589) <= (layer0_outputs(10939)) or (layer0_outputs(7634));
    outputs(10590) <= not((layer0_outputs(8347)) xor (layer0_outputs(6569)));
    outputs(10591) <= not(layer0_outputs(535));
    outputs(10592) <= not(layer0_outputs(959));
    outputs(10593) <= not((layer0_outputs(405)) and (layer0_outputs(11890)));
    outputs(10594) <= not((layer0_outputs(7577)) and (layer0_outputs(6505)));
    outputs(10595) <= not((layer0_outputs(7292)) and (layer0_outputs(2871)));
    outputs(10596) <= not((layer0_outputs(1119)) or (layer0_outputs(8578)));
    outputs(10597) <= (layer0_outputs(7025)) or (layer0_outputs(12000));
    outputs(10598) <= layer0_outputs(354);
    outputs(10599) <= layer0_outputs(4965);
    outputs(10600) <= not(layer0_outputs(9997)) or (layer0_outputs(4905));
    outputs(10601) <= (layer0_outputs(4625)) and (layer0_outputs(2650));
    outputs(10602) <= (layer0_outputs(11327)) xor (layer0_outputs(5261));
    outputs(10603) <= not((layer0_outputs(749)) xor (layer0_outputs(9080)));
    outputs(10604) <= not((layer0_outputs(10132)) xor (layer0_outputs(6763)));
    outputs(10605) <= not((layer0_outputs(11383)) xor (layer0_outputs(9345)));
    outputs(10606) <= layer0_outputs(8321);
    outputs(10607) <= (layer0_outputs(11544)) xor (layer0_outputs(3663));
    outputs(10608) <= (layer0_outputs(9842)) xor (layer0_outputs(11117));
    outputs(10609) <= layer0_outputs(9032);
    outputs(10610) <= (layer0_outputs(570)) xor (layer0_outputs(8077));
    outputs(10611) <= layer0_outputs(6723);
    outputs(10612) <= layer0_outputs(517);
    outputs(10613) <= not(layer0_outputs(93)) or (layer0_outputs(10628));
    outputs(10614) <= layer0_outputs(3515);
    outputs(10615) <= (layer0_outputs(4616)) xor (layer0_outputs(2584));
    outputs(10616) <= not((layer0_outputs(6062)) or (layer0_outputs(7034)));
    outputs(10617) <= layer0_outputs(10864);
    outputs(10618) <= (layer0_outputs(8195)) xor (layer0_outputs(11307));
    outputs(10619) <= not(layer0_outputs(12277));
    outputs(10620) <= not(layer0_outputs(3002));
    outputs(10621) <= layer0_outputs(5031);
    outputs(10622) <= not(layer0_outputs(9664));
    outputs(10623) <= not(layer0_outputs(6170));
    outputs(10624) <= layer0_outputs(7482);
    outputs(10625) <= not(layer0_outputs(3813));
    outputs(10626) <= not(layer0_outputs(12235));
    outputs(10627) <= not(layer0_outputs(1861)) or (layer0_outputs(12520));
    outputs(10628) <= (layer0_outputs(9492)) xor (layer0_outputs(3105));
    outputs(10629) <= not((layer0_outputs(11657)) xor (layer0_outputs(3198)));
    outputs(10630) <= not(layer0_outputs(9389));
    outputs(10631) <= not(layer0_outputs(10977)) or (layer0_outputs(8198));
    outputs(10632) <= not((layer0_outputs(12527)) xor (layer0_outputs(7422)));
    outputs(10633) <= not((layer0_outputs(7692)) and (layer0_outputs(4322)));
    outputs(10634) <= not(layer0_outputs(343)) or (layer0_outputs(9965));
    outputs(10635) <= (layer0_outputs(12732)) xor (layer0_outputs(7860));
    outputs(10636) <= not((layer0_outputs(11086)) xor (layer0_outputs(6023)));
    outputs(10637) <= (layer0_outputs(9732)) xor (layer0_outputs(8267));
    outputs(10638) <= not(layer0_outputs(3410));
    outputs(10639) <= layer0_outputs(5356);
    outputs(10640) <= not(layer0_outputs(819));
    outputs(10641) <= layer0_outputs(203);
    outputs(10642) <= not((layer0_outputs(9406)) or (layer0_outputs(11501)));
    outputs(10643) <= (layer0_outputs(2087)) or (layer0_outputs(5892));
    outputs(10644) <= layer0_outputs(2953);
    outputs(10645) <= not(layer0_outputs(7091));
    outputs(10646) <= not(layer0_outputs(8900));
    outputs(10647) <= not(layer0_outputs(5915)) or (layer0_outputs(12192));
    outputs(10648) <= (layer0_outputs(496)) xor (layer0_outputs(7715));
    outputs(10649) <= not((layer0_outputs(46)) xor (layer0_outputs(2729)));
    outputs(10650) <= layer0_outputs(5007);
    outputs(10651) <= (layer0_outputs(9007)) and not (layer0_outputs(2774));
    outputs(10652) <= layer0_outputs(2828);
    outputs(10653) <= (layer0_outputs(9039)) xor (layer0_outputs(2954));
    outputs(10654) <= not(layer0_outputs(12444));
    outputs(10655) <= (layer0_outputs(12369)) xor (layer0_outputs(2550));
    outputs(10656) <= not(layer0_outputs(4618)) or (layer0_outputs(8110));
    outputs(10657) <= not(layer0_outputs(12317));
    outputs(10658) <= not((layer0_outputs(9921)) xor (layer0_outputs(4597)));
    outputs(10659) <= (layer0_outputs(12155)) xor (layer0_outputs(4404));
    outputs(10660) <= layer0_outputs(8312);
    outputs(10661) <= layer0_outputs(5356);
    outputs(10662) <= layer0_outputs(8352);
    outputs(10663) <= not(layer0_outputs(5270));
    outputs(10664) <= (layer0_outputs(5954)) xor (layer0_outputs(5812));
    outputs(10665) <= not(layer0_outputs(8363));
    outputs(10666) <= not(layer0_outputs(7380)) or (layer0_outputs(5839));
    outputs(10667) <= not(layer0_outputs(8517));
    outputs(10668) <= not(layer0_outputs(4737)) or (layer0_outputs(5771));
    outputs(10669) <= (layer0_outputs(5800)) or (layer0_outputs(3184));
    outputs(10670) <= not(layer0_outputs(468));
    outputs(10671) <= (layer0_outputs(1612)) xor (layer0_outputs(12465));
    outputs(10672) <= not(layer0_outputs(1246)) or (layer0_outputs(9217));
    outputs(10673) <= not(layer0_outputs(3875));
    outputs(10674) <= not(layer0_outputs(589)) or (layer0_outputs(9596));
    outputs(10675) <= (layer0_outputs(5147)) or (layer0_outputs(3954));
    outputs(10676) <= (layer0_outputs(8097)) or (layer0_outputs(7798));
    outputs(10677) <= (layer0_outputs(10940)) xor (layer0_outputs(8094));
    outputs(10678) <= not(layer0_outputs(1546)) or (layer0_outputs(1014));
    outputs(10679) <= (layer0_outputs(2804)) xor (layer0_outputs(1750));
    outputs(10680) <= not(layer0_outputs(3790));
    outputs(10681) <= not((layer0_outputs(743)) xor (layer0_outputs(945)));
    outputs(10682) <= not(layer0_outputs(5777));
    outputs(10683) <= (layer0_outputs(10030)) xor (layer0_outputs(5312));
    outputs(10684) <= (layer0_outputs(4147)) xor (layer0_outputs(11209));
    outputs(10685) <= (layer0_outputs(11954)) xor (layer0_outputs(3343));
    outputs(10686) <= (layer0_outputs(6795)) xor (layer0_outputs(1051));
    outputs(10687) <= layer0_outputs(8052);
    outputs(10688) <= not(layer0_outputs(1333));
    outputs(10689) <= layer0_outputs(10720);
    outputs(10690) <= not((layer0_outputs(11917)) and (layer0_outputs(5521)));
    outputs(10691) <= not(layer0_outputs(5851));
    outputs(10692) <= (layer0_outputs(5770)) xor (layer0_outputs(7435));
    outputs(10693) <= not(layer0_outputs(3761));
    outputs(10694) <= layer0_outputs(9427);
    outputs(10695) <= not((layer0_outputs(11693)) and (layer0_outputs(12409)));
    outputs(10696) <= not((layer0_outputs(4425)) and (layer0_outputs(8067)));
    outputs(10697) <= not((layer0_outputs(2830)) and (layer0_outputs(265)));
    outputs(10698) <= (layer0_outputs(11709)) xor (layer0_outputs(8449));
    outputs(10699) <= not((layer0_outputs(9971)) xor (layer0_outputs(5916)));
    outputs(10700) <= layer0_outputs(3217);
    outputs(10701) <= not((layer0_outputs(8813)) and (layer0_outputs(10181)));
    outputs(10702) <= (layer0_outputs(10199)) or (layer0_outputs(12616));
    outputs(10703) <= not((layer0_outputs(202)) and (layer0_outputs(4452)));
    outputs(10704) <= not((layer0_outputs(5496)) xor (layer0_outputs(3536)));
    outputs(10705) <= not(layer0_outputs(806));
    outputs(10706) <= not(layer0_outputs(9568));
    outputs(10707) <= not((layer0_outputs(10356)) xor (layer0_outputs(886)));
    outputs(10708) <= not((layer0_outputs(3281)) xor (layer0_outputs(8103)));
    outputs(10709) <= (layer0_outputs(7073)) xor (layer0_outputs(608));
    outputs(10710) <= (layer0_outputs(5488)) xor (layer0_outputs(4295));
    outputs(10711) <= (layer0_outputs(12216)) xor (layer0_outputs(2092));
    outputs(10712) <= (layer0_outputs(4606)) and not (layer0_outputs(5598));
    outputs(10713) <= not(layer0_outputs(2289));
    outputs(10714) <= not(layer0_outputs(12486));
    outputs(10715) <= (layer0_outputs(10307)) or (layer0_outputs(4098));
    outputs(10716) <= (layer0_outputs(12501)) xor (layer0_outputs(6558));
    outputs(10717) <= (layer0_outputs(12362)) xor (layer0_outputs(6414));
    outputs(10718) <= not((layer0_outputs(8420)) xor (layer0_outputs(12645)));
    outputs(10719) <= not((layer0_outputs(2974)) xor (layer0_outputs(7555)));
    outputs(10720) <= not(layer0_outputs(5891)) or (layer0_outputs(8280));
    outputs(10721) <= layer0_outputs(1931);
    outputs(10722) <= not((layer0_outputs(6880)) xor (layer0_outputs(11098)));
    outputs(10723) <= not(layer0_outputs(12522));
    outputs(10724) <= (layer0_outputs(6312)) xor (layer0_outputs(349));
    outputs(10725) <= not(layer0_outputs(9330));
    outputs(10726) <= not(layer0_outputs(9232)) or (layer0_outputs(4347));
    outputs(10727) <= not((layer0_outputs(2197)) and (layer0_outputs(7167)));
    outputs(10728) <= not((layer0_outputs(5429)) and (layer0_outputs(6927)));
    outputs(10729) <= not((layer0_outputs(9908)) and (layer0_outputs(5863)));
    outputs(10730) <= not(layer0_outputs(10184)) or (layer0_outputs(3142));
    outputs(10731) <= layer0_outputs(3273);
    outputs(10732) <= layer0_outputs(3543);
    outputs(10733) <= not((layer0_outputs(10375)) xor (layer0_outputs(7107)));
    outputs(10734) <= not(layer0_outputs(901));
    outputs(10735) <= layer0_outputs(5917);
    outputs(10736) <= not((layer0_outputs(2914)) and (layer0_outputs(5010)));
    outputs(10737) <= layer0_outputs(6521);
    outputs(10738) <= not(layer0_outputs(332)) or (layer0_outputs(5066));
    outputs(10739) <= (layer0_outputs(11883)) and not (layer0_outputs(3442));
    outputs(10740) <= layer0_outputs(3697);
    outputs(10741) <= not(layer0_outputs(4601)) or (layer0_outputs(1184));
    outputs(10742) <= not(layer0_outputs(668)) or (layer0_outputs(7750));
    outputs(10743) <= layer0_outputs(1884);
    outputs(10744) <= not(layer0_outputs(4896));
    outputs(10745) <= not((layer0_outputs(4911)) or (layer0_outputs(4033)));
    outputs(10746) <= (layer0_outputs(7832)) or (layer0_outputs(11232));
    outputs(10747) <= (layer0_outputs(4627)) xor (layer0_outputs(7963));
    outputs(10748) <= not((layer0_outputs(2568)) xor (layer0_outputs(9476)));
    outputs(10749) <= (layer0_outputs(9536)) xor (layer0_outputs(3971));
    outputs(10750) <= (layer0_outputs(5759)) xor (layer0_outputs(2606));
    outputs(10751) <= (layer0_outputs(9760)) and not (layer0_outputs(9353));
    outputs(10752) <= not(layer0_outputs(6476));
    outputs(10753) <= (layer0_outputs(465)) or (layer0_outputs(361));
    outputs(10754) <= not(layer0_outputs(6344));
    outputs(10755) <= (layer0_outputs(5103)) or (layer0_outputs(2996));
    outputs(10756) <= not(layer0_outputs(6881)) or (layer0_outputs(4685));
    outputs(10757) <= not(layer0_outputs(10821));
    outputs(10758) <= not(layer0_outputs(12032));
    outputs(10759) <= not(layer0_outputs(9649)) or (layer0_outputs(7626));
    outputs(10760) <= not(layer0_outputs(8175)) or (layer0_outputs(1774));
    outputs(10761) <= (layer0_outputs(7764)) xor (layer0_outputs(5933));
    outputs(10762) <= not(layer0_outputs(482));
    outputs(10763) <= not(layer0_outputs(916)) or (layer0_outputs(5579));
    outputs(10764) <= not(layer0_outputs(8889)) or (layer0_outputs(7582));
    outputs(10765) <= not((layer0_outputs(5217)) and (layer0_outputs(6421)));
    outputs(10766) <= (layer0_outputs(3712)) xor (layer0_outputs(3478));
    outputs(10767) <= (layer0_outputs(10207)) or (layer0_outputs(3805));
    outputs(10768) <= not(layer0_outputs(5008));
    outputs(10769) <= (layer0_outputs(6044)) and not (layer0_outputs(3059));
    outputs(10770) <= (layer0_outputs(7467)) or (layer0_outputs(1403));
    outputs(10771) <= layer0_outputs(8374);
    outputs(10772) <= not((layer0_outputs(11083)) xor (layer0_outputs(12063)));
    outputs(10773) <= not((layer0_outputs(8627)) xor (layer0_outputs(5358)));
    outputs(10774) <= not(layer0_outputs(10342));
    outputs(10775) <= (layer0_outputs(9133)) or (layer0_outputs(5410));
    outputs(10776) <= (layer0_outputs(5444)) xor (layer0_outputs(5901));
    outputs(10777) <= layer0_outputs(6922);
    outputs(10778) <= not((layer0_outputs(10675)) xor (layer0_outputs(3848)));
    outputs(10779) <= not((layer0_outputs(8607)) and (layer0_outputs(976)));
    outputs(10780) <= (layer0_outputs(11564)) or (layer0_outputs(6731));
    outputs(10781) <= (layer0_outputs(3685)) xor (layer0_outputs(1055));
    outputs(10782) <= not((layer0_outputs(9055)) and (layer0_outputs(5801)));
    outputs(10783) <= layer0_outputs(2851);
    outputs(10784) <= not((layer0_outputs(12238)) xor (layer0_outputs(2691)));
    outputs(10785) <= not(layer0_outputs(549)) or (layer0_outputs(5992));
    outputs(10786) <= (layer0_outputs(2737)) or (layer0_outputs(8695));
    outputs(10787) <= not(layer0_outputs(11496)) or (layer0_outputs(5214));
    outputs(10788) <= not((layer0_outputs(5308)) and (layer0_outputs(3779)));
    outputs(10789) <= (layer0_outputs(8492)) xor (layer0_outputs(4677));
    outputs(10790) <= not(layer0_outputs(6426)) or (layer0_outputs(695));
    outputs(10791) <= not((layer0_outputs(5406)) xor (layer0_outputs(9750)));
    outputs(10792) <= not((layer0_outputs(901)) or (layer0_outputs(7793)));
    outputs(10793) <= not((layer0_outputs(2827)) xor (layer0_outputs(10480)));
    outputs(10794) <= not((layer0_outputs(6484)) xor (layer0_outputs(2325)));
    outputs(10795) <= not((layer0_outputs(1218)) xor (layer0_outputs(2971)));
    outputs(10796) <= not((layer0_outputs(9793)) xor (layer0_outputs(12629)));
    outputs(10797) <= not(layer0_outputs(9100));
    outputs(10798) <= layer0_outputs(9228);
    outputs(10799) <= not((layer0_outputs(8344)) or (layer0_outputs(689)));
    outputs(10800) <= (layer0_outputs(11378)) or (layer0_outputs(9882));
    outputs(10801) <= not(layer0_outputs(6454));
    outputs(10802) <= layer0_outputs(9689);
    outputs(10803) <= layer0_outputs(2892);
    outputs(10804) <= not(layer0_outputs(4706));
    outputs(10805) <= (layer0_outputs(1653)) and not (layer0_outputs(5319));
    outputs(10806) <= layer0_outputs(1835);
    outputs(10807) <= layer0_outputs(9891);
    outputs(10808) <= not((layer0_outputs(9812)) and (layer0_outputs(1985)));
    outputs(10809) <= (layer0_outputs(9889)) xor (layer0_outputs(5073));
    outputs(10810) <= not((layer0_outputs(7891)) xor (layer0_outputs(505)));
    outputs(10811) <= (layer0_outputs(3703)) xor (layer0_outputs(1349));
    outputs(10812) <= (layer0_outputs(6379)) xor (layer0_outputs(11716));
    outputs(10813) <= layer0_outputs(4659);
    outputs(10814) <= (layer0_outputs(9470)) or (layer0_outputs(8924));
    outputs(10815) <= not(layer0_outputs(7835)) or (layer0_outputs(5532));
    outputs(10816) <= not(layer0_outputs(9066)) or (layer0_outputs(5496));
    outputs(10817) <= not((layer0_outputs(609)) xor (layer0_outputs(3362)));
    outputs(10818) <= not((layer0_outputs(1020)) or (layer0_outputs(8247)));
    outputs(10819) <= (layer0_outputs(1160)) xor (layer0_outputs(4066));
    outputs(10820) <= not(layer0_outputs(4354));
    outputs(10821) <= (layer0_outputs(1583)) or (layer0_outputs(9829));
    outputs(10822) <= (layer0_outputs(3208)) or (layer0_outputs(9528));
    outputs(10823) <= (layer0_outputs(4447)) xor (layer0_outputs(8605));
    outputs(10824) <= (layer0_outputs(5339)) xor (layer0_outputs(3256));
    outputs(10825) <= not((layer0_outputs(3248)) xor (layer0_outputs(303)));
    outputs(10826) <= not((layer0_outputs(5564)) and (layer0_outputs(3784)));
    outputs(10827) <= not((layer0_outputs(12469)) and (layer0_outputs(7764)));
    outputs(10828) <= not((layer0_outputs(8821)) and (layer0_outputs(1529)));
    outputs(10829) <= not((layer0_outputs(3695)) xor (layer0_outputs(3919)));
    outputs(10830) <= not((layer0_outputs(5019)) xor (layer0_outputs(9122)));
    outputs(10831) <= not((layer0_outputs(8184)) xor (layer0_outputs(9927)));
    outputs(10832) <= (layer0_outputs(8350)) xor (layer0_outputs(4584));
    outputs(10833) <= (layer0_outputs(6690)) or (layer0_outputs(2306));
    outputs(10834) <= layer0_outputs(8646);
    outputs(10835) <= not((layer0_outputs(2626)) xor (layer0_outputs(5430)));
    outputs(10836) <= not(layer0_outputs(729)) or (layer0_outputs(6415));
    outputs(10837) <= (layer0_outputs(15)) or (layer0_outputs(10380));
    outputs(10838) <= (layer0_outputs(7050)) xor (layer0_outputs(1860));
    outputs(10839) <= not(layer0_outputs(8144)) or (layer0_outputs(9571));
    outputs(10840) <= not(layer0_outputs(4655));
    outputs(10841) <= not((layer0_outputs(6735)) xor (layer0_outputs(8456)));
    outputs(10842) <= layer0_outputs(4162);
    outputs(10843) <= layer0_outputs(12795);
    outputs(10844) <= not((layer0_outputs(3525)) xor (layer0_outputs(11609)));
    outputs(10845) <= (layer0_outputs(2362)) xor (layer0_outputs(12267));
    outputs(10846) <= not((layer0_outputs(4880)) or (layer0_outputs(11099)));
    outputs(10847) <= layer0_outputs(11858);
    outputs(10848) <= (layer0_outputs(3362)) and not (layer0_outputs(2725));
    outputs(10849) <= (layer0_outputs(5174)) xor (layer0_outputs(11449));
    outputs(10850) <= (layer0_outputs(4516)) xor (layer0_outputs(893));
    outputs(10851) <= (layer0_outputs(1239)) and not (layer0_outputs(10598));
    outputs(10852) <= not(layer0_outputs(974));
    outputs(10853) <= (layer0_outputs(2950)) xor (layer0_outputs(5381));
    outputs(10854) <= layer0_outputs(5985);
    outputs(10855) <= not(layer0_outputs(3326));
    outputs(10856) <= layer0_outputs(899);
    outputs(10857) <= (layer0_outputs(11205)) or (layer0_outputs(5476));
    outputs(10858) <= not(layer0_outputs(11260));
    outputs(10859) <= not(layer0_outputs(7952));
    outputs(10860) <= not((layer0_outputs(9933)) xor (layer0_outputs(9511)));
    outputs(10861) <= layer0_outputs(5124);
    outputs(10862) <= not(layer0_outputs(1601));
    outputs(10863) <= not((layer0_outputs(7984)) xor (layer0_outputs(6508)));
    outputs(10864) <= (layer0_outputs(10229)) xor (layer0_outputs(3972));
    outputs(10865) <= (layer0_outputs(10942)) xor (layer0_outputs(177));
    outputs(10866) <= (layer0_outputs(11887)) or (layer0_outputs(6919));
    outputs(10867) <= (layer0_outputs(2844)) and (layer0_outputs(5730));
    outputs(10868) <= (layer0_outputs(12478)) or (layer0_outputs(147));
    outputs(10869) <= not((layer0_outputs(9871)) xor (layer0_outputs(5801)));
    outputs(10870) <= layer0_outputs(12750);
    outputs(10871) <= not(layer0_outputs(11667)) or (layer0_outputs(2563));
    outputs(10872) <= (layer0_outputs(12519)) xor (layer0_outputs(6914));
    outputs(10873) <= not(layer0_outputs(9529));
    outputs(10874) <= (layer0_outputs(10216)) and not (layer0_outputs(12475));
    outputs(10875) <= layer0_outputs(6746);
    outputs(10876) <= not(layer0_outputs(915)) or (layer0_outputs(3383));
    outputs(10877) <= not(layer0_outputs(442));
    outputs(10878) <= not((layer0_outputs(4045)) xor (layer0_outputs(2659)));
    outputs(10879) <= not(layer0_outputs(11441));
    outputs(10880) <= layer0_outputs(6813);
    outputs(10881) <= not((layer0_outputs(6753)) xor (layer0_outputs(11921)));
    outputs(10882) <= layer0_outputs(12260);
    outputs(10883) <= (layer0_outputs(7618)) or (layer0_outputs(8862));
    outputs(10884) <= not((layer0_outputs(9387)) or (layer0_outputs(11021)));
    outputs(10885) <= not((layer0_outputs(11156)) xor (layer0_outputs(417)));
    outputs(10886) <= not(layer0_outputs(9248)) or (layer0_outputs(4532));
    outputs(10887) <= layer0_outputs(5917);
    outputs(10888) <= not((layer0_outputs(4620)) xor (layer0_outputs(3661)));
    outputs(10889) <= not(layer0_outputs(11965));
    outputs(10890) <= not((layer0_outputs(85)) xor (layer0_outputs(10544)));
    outputs(10891) <= not(layer0_outputs(737)) or (layer0_outputs(8303));
    outputs(10892) <= not((layer0_outputs(10392)) xor (layer0_outputs(2837)));
    outputs(10893) <= not(layer0_outputs(7624));
    outputs(10894) <= not((layer0_outputs(9418)) and (layer0_outputs(10238)));
    outputs(10895) <= not((layer0_outputs(9299)) xor (layer0_outputs(3335)));
    outputs(10896) <= (layer0_outputs(5530)) xor (layer0_outputs(5144));
    outputs(10897) <= (layer0_outputs(7879)) xor (layer0_outputs(2087));
    outputs(10898) <= (layer0_outputs(10871)) xor (layer0_outputs(7985));
    outputs(10899) <= (layer0_outputs(8658)) and (layer0_outputs(3210));
    outputs(10900) <= not(layer0_outputs(3692)) or (layer0_outputs(11469));
    outputs(10901) <= layer0_outputs(6510);
    outputs(10902) <= (layer0_outputs(5544)) xor (layer0_outputs(8079));
    outputs(10903) <= (layer0_outputs(6873)) and not (layer0_outputs(3558));
    outputs(10904) <= not(layer0_outputs(11394));
    outputs(10905) <= not(layer0_outputs(2140));
    outputs(10906) <= layer0_outputs(3825);
    outputs(10907) <= not((layer0_outputs(10797)) xor (layer0_outputs(4461)));
    outputs(10908) <= layer0_outputs(11559);
    outputs(10909) <= layer0_outputs(11248);
    outputs(10910) <= layer0_outputs(5509);
    outputs(10911) <= (layer0_outputs(11922)) or (layer0_outputs(773));
    outputs(10912) <= not(layer0_outputs(9573));
    outputs(10913) <= (layer0_outputs(9731)) and (layer0_outputs(11047));
    outputs(10914) <= (layer0_outputs(3808)) and (layer0_outputs(4414));
    outputs(10915) <= not(layer0_outputs(12088));
    outputs(10916) <= not(layer0_outputs(2447)) or (layer0_outputs(12194));
    outputs(10917) <= not((layer0_outputs(3051)) xor (layer0_outputs(5387)));
    outputs(10918) <= not(layer0_outputs(10444));
    outputs(10919) <= not(layer0_outputs(2181));
    outputs(10920) <= (layer0_outputs(11322)) xor (layer0_outputs(11695));
    outputs(10921) <= (layer0_outputs(7813)) xor (layer0_outputs(2923));
    outputs(10922) <= not(layer0_outputs(3152));
    outputs(10923) <= (layer0_outputs(7000)) xor (layer0_outputs(10676));
    outputs(10924) <= (layer0_outputs(6053)) xor (layer0_outputs(8501));
    outputs(10925) <= not(layer0_outputs(6667)) or (layer0_outputs(162));
    outputs(10926) <= layer0_outputs(11994);
    outputs(10927) <= not(layer0_outputs(9975)) or (layer0_outputs(9131));
    outputs(10928) <= not(layer0_outputs(8531)) or (layer0_outputs(11286));
    outputs(10929) <= (layer0_outputs(1731)) xor (layer0_outputs(1658));
    outputs(10930) <= (layer0_outputs(900)) xor (layer0_outputs(11455));
    outputs(10931) <= (layer0_outputs(3230)) xor (layer0_outputs(3467));
    outputs(10932) <= layer0_outputs(4546);
    outputs(10933) <= not((layer0_outputs(4326)) xor (layer0_outputs(8318)));
    outputs(10934) <= layer0_outputs(3111);
    outputs(10935) <= (layer0_outputs(1865)) and not (layer0_outputs(7517));
    outputs(10936) <= not(layer0_outputs(3397)) or (layer0_outputs(11465));
    outputs(10937) <= (layer0_outputs(11387)) xor (layer0_outputs(11885));
    outputs(10938) <= layer0_outputs(5436);
    outputs(10939) <= layer0_outputs(4886);
    outputs(10940) <= not((layer0_outputs(2649)) and (layer0_outputs(4746)));
    outputs(10941) <= not((layer0_outputs(10365)) xor (layer0_outputs(6563)));
    outputs(10942) <= (layer0_outputs(779)) xor (layer0_outputs(10471));
    outputs(10943) <= not(layer0_outputs(2809));
    outputs(10944) <= not((layer0_outputs(2778)) xor (layer0_outputs(6414)));
    outputs(10945) <= layer0_outputs(8298);
    outputs(10946) <= not((layer0_outputs(1252)) xor (layer0_outputs(11520)));
    outputs(10947) <= not((layer0_outputs(10323)) or (layer0_outputs(1912)));
    outputs(10948) <= not(layer0_outputs(5663));
    outputs(10949) <= not((layer0_outputs(10064)) xor (layer0_outputs(4334)));
    outputs(10950) <= not(layer0_outputs(2517));
    outputs(10951) <= not((layer0_outputs(6932)) xor (layer0_outputs(9857)));
    outputs(10952) <= layer0_outputs(8237);
    outputs(10953) <= (layer0_outputs(1386)) xor (layer0_outputs(2072));
    outputs(10954) <= not(layer0_outputs(4911));
    outputs(10955) <= not((layer0_outputs(7826)) xor (layer0_outputs(12065)));
    outputs(10956) <= (layer0_outputs(5397)) xor (layer0_outputs(2909));
    outputs(10957) <= (layer0_outputs(5291)) xor (layer0_outputs(9747));
    outputs(10958) <= not((layer0_outputs(10925)) xor (layer0_outputs(5333)));
    outputs(10959) <= not(layer0_outputs(12451));
    outputs(10960) <= not(layer0_outputs(12545));
    outputs(10961) <= (layer0_outputs(2713)) xor (layer0_outputs(9879));
    outputs(10962) <= not(layer0_outputs(1232));
    outputs(10963) <= not((layer0_outputs(7358)) xor (layer0_outputs(6397)));
    outputs(10964) <= (layer0_outputs(3449)) xor (layer0_outputs(5223));
    outputs(10965) <= (layer0_outputs(925)) or (layer0_outputs(12254));
    outputs(10966) <= not((layer0_outputs(3685)) xor (layer0_outputs(2112)));
    outputs(10967) <= not(layer0_outputs(867)) or (layer0_outputs(7582));
    outputs(10968) <= not((layer0_outputs(11879)) xor (layer0_outputs(10965)));
    outputs(10969) <= (layer0_outputs(973)) xor (layer0_outputs(6672));
    outputs(10970) <= not(layer0_outputs(1372));
    outputs(10971) <= not(layer0_outputs(2793)) or (layer0_outputs(2707));
    outputs(10972) <= not((layer0_outputs(5626)) xor (layer0_outputs(5744)));
    outputs(10973) <= not((layer0_outputs(6747)) xor (layer0_outputs(3235)));
    outputs(10974) <= not((layer0_outputs(11228)) xor (layer0_outputs(7408)));
    outputs(10975) <= (layer0_outputs(10648)) xor (layer0_outputs(10916));
    outputs(10976) <= not(layer0_outputs(7350)) or (layer0_outputs(309));
    outputs(10977) <= (layer0_outputs(8920)) xor (layer0_outputs(2664));
    outputs(10978) <= not((layer0_outputs(2614)) and (layer0_outputs(7899)));
    outputs(10979) <= not((layer0_outputs(159)) and (layer0_outputs(8379)));
    outputs(10980) <= not(layer0_outputs(9641));
    outputs(10981) <= not(layer0_outputs(1740));
    outputs(10982) <= (layer0_outputs(5040)) xor (layer0_outputs(7933));
    outputs(10983) <= (layer0_outputs(8457)) and not (layer0_outputs(8536));
    outputs(10984) <= not(layer0_outputs(7180)) or (layer0_outputs(11771));
    outputs(10985) <= not(layer0_outputs(7486));
    outputs(10986) <= (layer0_outputs(6430)) xor (layer0_outputs(12338));
    outputs(10987) <= not(layer0_outputs(11856));
    outputs(10988) <= layer0_outputs(286);
    outputs(10989) <= layer0_outputs(8841);
    outputs(10990) <= not(layer0_outputs(2524));
    outputs(10991) <= not((layer0_outputs(3052)) and (layer0_outputs(10478)));
    outputs(10992) <= layer0_outputs(5675);
    outputs(10993) <= (layer0_outputs(1510)) xor (layer0_outputs(249));
    outputs(10994) <= not((layer0_outputs(3112)) or (layer0_outputs(2258)));
    outputs(10995) <= layer0_outputs(1462);
    outputs(10996) <= not(layer0_outputs(12239)) or (layer0_outputs(1704));
    outputs(10997) <= not((layer0_outputs(11334)) xor (layer0_outputs(2968)));
    outputs(10998) <= not(layer0_outputs(3442)) or (layer0_outputs(4544));
    outputs(10999) <= not((layer0_outputs(4139)) xor (layer0_outputs(12000)));
    outputs(11000) <= (layer0_outputs(3266)) xor (layer0_outputs(10794));
    outputs(11001) <= not(layer0_outputs(6186));
    outputs(11002) <= not(layer0_outputs(1839));
    outputs(11003) <= layer0_outputs(11688);
    outputs(11004) <= not(layer0_outputs(6766));
    outputs(11005) <= (layer0_outputs(2721)) xor (layer0_outputs(8426));
    outputs(11006) <= (layer0_outputs(4262)) and (layer0_outputs(3446));
    outputs(11007) <= not(layer0_outputs(8740));
    outputs(11008) <= not(layer0_outputs(2346)) or (layer0_outputs(2864));
    outputs(11009) <= layer0_outputs(229);
    outputs(11010) <= not(layer0_outputs(3739)) or (layer0_outputs(11210));
    outputs(11011) <= layer0_outputs(5231);
    outputs(11012) <= not((layer0_outputs(10870)) xor (layer0_outputs(6176)));
    outputs(11013) <= not((layer0_outputs(7016)) xor (layer0_outputs(10496)));
    outputs(11014) <= not((layer0_outputs(6445)) xor (layer0_outputs(11821)));
    outputs(11015) <= (layer0_outputs(8929)) xor (layer0_outputs(11152));
    outputs(11016) <= not((layer0_outputs(3913)) or (layer0_outputs(10074)));
    outputs(11017) <= not((layer0_outputs(11829)) and (layer0_outputs(6365)));
    outputs(11018) <= not((layer0_outputs(10963)) xor (layer0_outputs(1599)));
    outputs(11019) <= (layer0_outputs(8585)) xor (layer0_outputs(715));
    outputs(11020) <= (layer0_outputs(4092)) xor (layer0_outputs(2768));
    outputs(11021) <= layer0_outputs(8168);
    outputs(11022) <= not(layer0_outputs(10049)) or (layer0_outputs(3147));
    outputs(11023) <= not((layer0_outputs(8692)) xor (layer0_outputs(9513)));
    outputs(11024) <= not(layer0_outputs(9441));
    outputs(11025) <= layer0_outputs(1592);
    outputs(11026) <= layer0_outputs(8671);
    outputs(11027) <= not((layer0_outputs(11982)) xor (layer0_outputs(3214)));
    outputs(11028) <= not((layer0_outputs(9198)) or (layer0_outputs(11988)));
    outputs(11029) <= (layer0_outputs(6357)) xor (layer0_outputs(759));
    outputs(11030) <= not((layer0_outputs(804)) or (layer0_outputs(3262)));
    outputs(11031) <= not(layer0_outputs(118)) or (layer0_outputs(10735));
    outputs(11032) <= (layer0_outputs(7820)) xor (layer0_outputs(8782));
    outputs(11033) <= not(layer0_outputs(7117)) or (layer0_outputs(5443));
    outputs(11034) <= not((layer0_outputs(1470)) xor (layer0_outputs(8893)));
    outputs(11035) <= layer0_outputs(6671);
    outputs(11036) <= not(layer0_outputs(9027));
    outputs(11037) <= not((layer0_outputs(75)) xor (layer0_outputs(371)));
    outputs(11038) <= not(layer0_outputs(6248));
    outputs(11039) <= layer0_outputs(7186);
    outputs(11040) <= layer0_outputs(1081);
    outputs(11041) <= not((layer0_outputs(2246)) xor (layer0_outputs(9976)));
    outputs(11042) <= not((layer0_outputs(12206)) xor (layer0_outputs(1104)));
    outputs(11043) <= not(layer0_outputs(3479));
    outputs(11044) <= layer0_outputs(7362);
    outputs(11045) <= (layer0_outputs(3033)) xor (layer0_outputs(3925));
    outputs(11046) <= not(layer0_outputs(4093)) or (layer0_outputs(1673));
    outputs(11047) <= not((layer0_outputs(574)) and (layer0_outputs(12683)));
    outputs(11048) <= not((layer0_outputs(2289)) xor (layer0_outputs(8150)));
    outputs(11049) <= (layer0_outputs(3551)) xor (layer0_outputs(7892));
    outputs(11050) <= not((layer0_outputs(8950)) xor (layer0_outputs(11812)));
    outputs(11051) <= not((layer0_outputs(2228)) xor (layer0_outputs(2874)));
    outputs(11052) <= (layer0_outputs(11492)) xor (layer0_outputs(12085));
    outputs(11053) <= not(layer0_outputs(9836));
    outputs(11054) <= layer0_outputs(1672);
    outputs(11055) <= not(layer0_outputs(8826));
    outputs(11056) <= not((layer0_outputs(6543)) xor (layer0_outputs(7586)));
    outputs(11057) <= not((layer0_outputs(4962)) and (layer0_outputs(641)));
    outputs(11058) <= not((layer0_outputs(3694)) xor (layer0_outputs(1563)));
    outputs(11059) <= not(layer0_outputs(6560));
    outputs(11060) <= not((layer0_outputs(8283)) xor (layer0_outputs(543)));
    outputs(11061) <= not((layer0_outputs(9332)) xor (layer0_outputs(7446)));
    outputs(11062) <= (layer0_outputs(7926)) or (layer0_outputs(9712));
    outputs(11063) <= not(layer0_outputs(8256));
    outputs(11064) <= (layer0_outputs(7971)) and not (layer0_outputs(1287));
    outputs(11065) <= not((layer0_outputs(6160)) xor (layer0_outputs(1278)));
    outputs(11066) <= (layer0_outputs(5011)) and not (layer0_outputs(4171));
    outputs(11067) <= not((layer0_outputs(12062)) xor (layer0_outputs(11564)));
    outputs(11068) <= not(layer0_outputs(9481));
    outputs(11069) <= (layer0_outputs(3008)) or (layer0_outputs(10026));
    outputs(11070) <= not((layer0_outputs(8696)) xor (layer0_outputs(2467)));
    outputs(11071) <= not(layer0_outputs(7966)) or (layer0_outputs(5897));
    outputs(11072) <= not(layer0_outputs(3240)) or (layer0_outputs(9278));
    outputs(11073) <= layer0_outputs(1002);
    outputs(11074) <= (layer0_outputs(1988)) and not (layer0_outputs(70));
    outputs(11075) <= (layer0_outputs(11898)) or (layer0_outputs(12015));
    outputs(11076) <= (layer0_outputs(4791)) xor (layer0_outputs(11277));
    outputs(11077) <= not((layer0_outputs(3603)) xor (layer0_outputs(3736)));
    outputs(11078) <= not((layer0_outputs(7360)) and (layer0_outputs(12495)));
    outputs(11079) <= not(layer0_outputs(1915)) or (layer0_outputs(4860));
    outputs(11080) <= not((layer0_outputs(2795)) xor (layer0_outputs(6577)));
    outputs(11081) <= (layer0_outputs(2571)) or (layer0_outputs(9369));
    outputs(11082) <= (layer0_outputs(5767)) xor (layer0_outputs(6404));
    outputs(11083) <= not(layer0_outputs(10007)) or (layer0_outputs(11548));
    outputs(11084) <= (layer0_outputs(1042)) xor (layer0_outputs(6104));
    outputs(11085) <= layer0_outputs(9855);
    outputs(11086) <= not(layer0_outputs(4774)) or (layer0_outputs(1068));
    outputs(11087) <= not(layer0_outputs(6912)) or (layer0_outputs(11138));
    outputs(11088) <= not((layer0_outputs(8564)) xor (layer0_outputs(5712)));
    outputs(11089) <= layer0_outputs(9335);
    outputs(11090) <= not((layer0_outputs(982)) xor (layer0_outputs(10565)));
    outputs(11091) <= layer0_outputs(10299);
    outputs(11092) <= layer0_outputs(6277);
    outputs(11093) <= not((layer0_outputs(1894)) xor (layer0_outputs(11797)));
    outputs(11094) <= not((layer0_outputs(9638)) or (layer0_outputs(12661)));
    outputs(11095) <= not((layer0_outputs(9785)) and (layer0_outputs(3418)));
    outputs(11096) <= layer0_outputs(4864);
    outputs(11097) <= not((layer0_outputs(9101)) xor (layer0_outputs(1187)));
    outputs(11098) <= not((layer0_outputs(8623)) xor (layer0_outputs(9576)));
    outputs(11099) <= (layer0_outputs(2206)) xor (layer0_outputs(1688));
    outputs(11100) <= (layer0_outputs(9440)) xor (layer0_outputs(7886));
    outputs(11101) <= (layer0_outputs(5090)) xor (layer0_outputs(12641));
    outputs(11102) <= not(layer0_outputs(2951));
    outputs(11103) <= not(layer0_outputs(3615)) or (layer0_outputs(12798));
    outputs(11104) <= not(layer0_outputs(9637));
    outputs(11105) <= not(layer0_outputs(5069));
    outputs(11106) <= layer0_outputs(11567);
    outputs(11107) <= not((layer0_outputs(11236)) xor (layer0_outputs(396)));
    outputs(11108) <= not((layer0_outputs(11856)) xor (layer0_outputs(3956)));
    outputs(11109) <= not(layer0_outputs(1486));
    outputs(11110) <= not(layer0_outputs(4268));
    outputs(11111) <= (layer0_outputs(6024)) xor (layer0_outputs(555));
    outputs(11112) <= not(layer0_outputs(9372));
    outputs(11113) <= (layer0_outputs(3327)) or (layer0_outputs(1406));
    outputs(11114) <= not((layer0_outputs(2530)) or (layer0_outputs(7967)));
    outputs(11115) <= not((layer0_outputs(1585)) and (layer0_outputs(9819)));
    outputs(11116) <= layer0_outputs(5941);
    outputs(11117) <= not(layer0_outputs(6979)) or (layer0_outputs(3229));
    outputs(11118) <= not((layer0_outputs(1255)) xor (layer0_outputs(6636)));
    outputs(11119) <= not((layer0_outputs(2730)) xor (layer0_outputs(983)));
    outputs(11120) <= not((layer0_outputs(6631)) and (layer0_outputs(1055)));
    outputs(11121) <= (layer0_outputs(7838)) and not (layer0_outputs(2883));
    outputs(11122) <= not((layer0_outputs(3604)) or (layer0_outputs(1377)));
    outputs(11123) <= not(layer0_outputs(5904));
    outputs(11124) <= not(layer0_outputs(9192)) or (layer0_outputs(1914));
    outputs(11125) <= not((layer0_outputs(1939)) xor (layer0_outputs(9952)));
    outputs(11126) <= not((layer0_outputs(1904)) and (layer0_outputs(9721)));
    outputs(11127) <= not((layer0_outputs(10958)) or (layer0_outputs(2745)));
    outputs(11128) <= (layer0_outputs(11911)) xor (layer0_outputs(9925));
    outputs(11129) <= not((layer0_outputs(9310)) xor (layer0_outputs(7679)));
    outputs(11130) <= layer0_outputs(187);
    outputs(11131) <= (layer0_outputs(6693)) xor (layer0_outputs(12658));
    outputs(11132) <= not((layer0_outputs(9987)) xor (layer0_outputs(6605)));
    outputs(11133) <= not((layer0_outputs(3411)) xor (layer0_outputs(3506)));
    outputs(11134) <= (layer0_outputs(8639)) xor (layer0_outputs(5269));
    outputs(11135) <= layer0_outputs(753);
    outputs(11136) <= not(layer0_outputs(1613));
    outputs(11137) <= not((layer0_outputs(11278)) and (layer0_outputs(5980)));
    outputs(11138) <= not(layer0_outputs(1129)) or (layer0_outputs(6409));
    outputs(11139) <= '1';
    outputs(11140) <= not(layer0_outputs(5677));
    outputs(11141) <= layer0_outputs(12767);
    outputs(11142) <= (layer0_outputs(8199)) or (layer0_outputs(11319));
    outputs(11143) <= layer0_outputs(7745);
    outputs(11144) <= (layer0_outputs(7668)) and not (layer0_outputs(12744));
    outputs(11145) <= (layer0_outputs(4121)) xor (layer0_outputs(2579));
    outputs(11146) <= not((layer0_outputs(1742)) or (layer0_outputs(2271)));
    outputs(11147) <= layer0_outputs(459);
    outputs(11148) <= layer0_outputs(10643);
    outputs(11149) <= not((layer0_outputs(10111)) and (layer0_outputs(4744)));
    outputs(11150) <= (layer0_outputs(1487)) xor (layer0_outputs(6456));
    outputs(11151) <= not((layer0_outputs(9829)) xor (layer0_outputs(10210)));
    outputs(11152) <= layer0_outputs(2885);
    outputs(11153) <= not(layer0_outputs(8938)) or (layer0_outputs(12285));
    outputs(11154) <= not(layer0_outputs(10452)) or (layer0_outputs(12012));
    outputs(11155) <= layer0_outputs(8438);
    outputs(11156) <= not(layer0_outputs(1391));
    outputs(11157) <= (layer0_outputs(3164)) xor (layer0_outputs(11217));
    outputs(11158) <= not((layer0_outputs(8242)) and (layer0_outputs(3160)));
    outputs(11159) <= not((layer0_outputs(10403)) xor (layer0_outputs(8743)));
    outputs(11160) <= layer0_outputs(984);
    outputs(11161) <= not(layer0_outputs(1121));
    outputs(11162) <= (layer0_outputs(1123)) xor (layer0_outputs(10652));
    outputs(11163) <= (layer0_outputs(1166)) xor (layer0_outputs(9668));
    outputs(11164) <= not(layer0_outputs(8668)) or (layer0_outputs(8702));
    outputs(11165) <= (layer0_outputs(11743)) xor (layer0_outputs(9618));
    outputs(11166) <= not(layer0_outputs(4208)) or (layer0_outputs(2509));
    outputs(11167) <= not(layer0_outputs(9366));
    outputs(11168) <= layer0_outputs(12799);
    outputs(11169) <= (layer0_outputs(4692)) xor (layer0_outputs(6087));
    outputs(11170) <= layer0_outputs(1425);
    outputs(11171) <= not(layer0_outputs(3374));
    outputs(11172) <= not(layer0_outputs(1262));
    outputs(11173) <= layer0_outputs(3183);
    outputs(11174) <= layer0_outputs(3566);
    outputs(11175) <= not(layer0_outputs(10445));
    outputs(11176) <= not(layer0_outputs(12073)) or (layer0_outputs(7386));
    outputs(11177) <= (layer0_outputs(12413)) xor (layer0_outputs(5550));
    outputs(11178) <= not(layer0_outputs(2696));
    outputs(11179) <= not((layer0_outputs(7156)) xor (layer0_outputs(5046)));
    outputs(11180) <= not((layer0_outputs(11760)) or (layer0_outputs(7556)));
    outputs(11181) <= not(layer0_outputs(2113));
    outputs(11182) <= layer0_outputs(6256);
    outputs(11183) <= (layer0_outputs(7072)) xor (layer0_outputs(3514));
    outputs(11184) <= (layer0_outputs(7227)) and not (layer0_outputs(3219));
    outputs(11185) <= not((layer0_outputs(4318)) and (layer0_outputs(1019)));
    outputs(11186) <= not((layer0_outputs(2613)) or (layer0_outputs(5240)));
    outputs(11187) <= not(layer0_outputs(4328));
    outputs(11188) <= (layer0_outputs(4424)) xor (layer0_outputs(17));
    outputs(11189) <= not((layer0_outputs(2779)) xor (layer0_outputs(8373)));
    outputs(11190) <= layer0_outputs(8117);
    outputs(11191) <= not(layer0_outputs(6464)) or (layer0_outputs(7782));
    outputs(11192) <= (layer0_outputs(1066)) or (layer0_outputs(11997));
    outputs(11193) <= not(layer0_outputs(5558));
    outputs(11194) <= not(layer0_outputs(4014)) or (layer0_outputs(1612));
    outputs(11195) <= (layer0_outputs(10194)) xor (layer0_outputs(9837));
    outputs(11196) <= layer0_outputs(1328);
    outputs(11197) <= not(layer0_outputs(9681));
    outputs(11198) <= not(layer0_outputs(1855));
    outputs(11199) <= (layer0_outputs(7487)) xor (layer0_outputs(6043));
    outputs(11200) <= not(layer0_outputs(3942)) or (layer0_outputs(8732));
    outputs(11201) <= layer0_outputs(6465);
    outputs(11202) <= (layer0_outputs(3487)) xor (layer0_outputs(490));
    outputs(11203) <= not(layer0_outputs(9834)) or (layer0_outputs(3832));
    outputs(11204) <= (layer0_outputs(7303)) and not (layer0_outputs(10956));
    outputs(11205) <= layer0_outputs(3962);
    outputs(11206) <= layer0_outputs(5198);
    outputs(11207) <= not((layer0_outputs(6284)) xor (layer0_outputs(5875)));
    outputs(11208) <= not(layer0_outputs(4610));
    outputs(11209) <= not((layer0_outputs(9216)) xor (layer0_outputs(3842)));
    outputs(11210) <= layer0_outputs(4631);
    outputs(11211) <= not(layer0_outputs(4915));
    outputs(11212) <= not((layer0_outputs(7546)) or (layer0_outputs(8821)));
    outputs(11213) <= (layer0_outputs(2574)) and (layer0_outputs(9171));
    outputs(11214) <= (layer0_outputs(1365)) xor (layer0_outputs(6562));
    outputs(11215) <= layer0_outputs(5477);
    outputs(11216) <= not((layer0_outputs(1100)) xor (layer0_outputs(12383)));
    outputs(11217) <= (layer0_outputs(2516)) or (layer0_outputs(12401));
    outputs(11218) <= layer0_outputs(77);
    outputs(11219) <= not((layer0_outputs(5023)) xor (layer0_outputs(3113)));
    outputs(11220) <= (layer0_outputs(1448)) xor (layer0_outputs(8875));
    outputs(11221) <= (layer0_outputs(10827)) xor (layer0_outputs(5383));
    outputs(11222) <= (layer0_outputs(10712)) or (layer0_outputs(2298));
    outputs(11223) <= not(layer0_outputs(2279));
    outputs(11224) <= not(layer0_outputs(4257));
    outputs(11225) <= not((layer0_outputs(10208)) xor (layer0_outputs(10579)));
    outputs(11226) <= not((layer0_outputs(11807)) xor (layer0_outputs(12540)));
    outputs(11227) <= not((layer0_outputs(445)) or (layer0_outputs(1076)));
    outputs(11228) <= layer0_outputs(2350);
    outputs(11229) <= not(layer0_outputs(6153));
    outputs(11230) <= layer0_outputs(11962);
    outputs(11231) <= (layer0_outputs(6462)) xor (layer0_outputs(6874));
    outputs(11232) <= not(layer0_outputs(1372));
    outputs(11233) <= (layer0_outputs(3019)) xor (layer0_outputs(6638));
    outputs(11234) <= not(layer0_outputs(6501));
    outputs(11235) <= layer0_outputs(9396);
    outputs(11236) <= (layer0_outputs(630)) xor (layer0_outputs(5679));
    outputs(11237) <= (layer0_outputs(7708)) or (layer0_outputs(11817));
    outputs(11238) <= not((layer0_outputs(9432)) xor (layer0_outputs(9479)));
    outputs(11239) <= not((layer0_outputs(2110)) xor (layer0_outputs(10262)));
    outputs(11240) <= not((layer0_outputs(6563)) xor (layer0_outputs(7235)));
    outputs(11241) <= not((layer0_outputs(6078)) xor (layer0_outputs(9195)));
    outputs(11242) <= not(layer0_outputs(4615));
    outputs(11243) <= not((layer0_outputs(8070)) xor (layer0_outputs(8246)));
    outputs(11244) <= not(layer0_outputs(5251));
    outputs(11245) <= not((layer0_outputs(3628)) xor (layer0_outputs(9998)));
    outputs(11246) <= not(layer0_outputs(7749));
    outputs(11247) <= layer0_outputs(5271);
    outputs(11248) <= (layer0_outputs(10708)) or (layer0_outputs(3807));
    outputs(11249) <= layer0_outputs(4352);
    outputs(11250) <= (layer0_outputs(10284)) or (layer0_outputs(8908));
    outputs(11251) <= not((layer0_outputs(11619)) xor (layer0_outputs(6068)));
    outputs(11252) <= layer0_outputs(6629);
    outputs(11253) <= not((layer0_outputs(5263)) and (layer0_outputs(1012)));
    outputs(11254) <= (layer0_outputs(5984)) and not (layer0_outputs(4628));
    outputs(11255) <= not((layer0_outputs(610)) and (layer0_outputs(10077)));
    outputs(11256) <= not((layer0_outputs(6125)) xor (layer0_outputs(2286)));
    outputs(11257) <= not((layer0_outputs(12240)) xor (layer0_outputs(5138)));
    outputs(11258) <= not((layer0_outputs(11070)) xor (layer0_outputs(9966)));
    outputs(11259) <= layer0_outputs(7671);
    outputs(11260) <= not(layer0_outputs(8525));
    outputs(11261) <= not((layer0_outputs(12638)) xor (layer0_outputs(115)));
    outputs(11262) <= (layer0_outputs(6640)) or (layer0_outputs(134));
    outputs(11263) <= not(layer0_outputs(4280));
    outputs(11264) <= (layer0_outputs(5487)) and not (layer0_outputs(1144));
    outputs(11265) <= layer0_outputs(3829);
    outputs(11266) <= (layer0_outputs(4668)) xor (layer0_outputs(11471));
    outputs(11267) <= not(layer0_outputs(4785));
    outputs(11268) <= not((layer0_outputs(8638)) and (layer0_outputs(10878)));
    outputs(11269) <= not(layer0_outputs(4041));
    outputs(11270) <= not(layer0_outputs(5597));
    outputs(11271) <= layer0_outputs(7386);
    outputs(11272) <= layer0_outputs(12601);
    outputs(11273) <= not(layer0_outputs(1084)) or (layer0_outputs(8976));
    outputs(11274) <= not(layer0_outputs(5763));
    outputs(11275) <= not(layer0_outputs(11314));
    outputs(11276) <= not((layer0_outputs(4235)) and (layer0_outputs(11398)));
    outputs(11277) <= (layer0_outputs(4207)) and not (layer0_outputs(320));
    outputs(11278) <= (layer0_outputs(11740)) and (layer0_outputs(10165));
    outputs(11279) <= layer0_outputs(3508);
    outputs(11280) <= (layer0_outputs(7192)) or (layer0_outputs(4042));
    outputs(11281) <= (layer0_outputs(11127)) and not (layer0_outputs(12267));
    outputs(11282) <= (layer0_outputs(10584)) and not (layer0_outputs(7808));
    outputs(11283) <= not(layer0_outputs(9743));
    outputs(11284) <= not((layer0_outputs(298)) and (layer0_outputs(5189)));
    outputs(11285) <= (layer0_outputs(7581)) and not (layer0_outputs(1521));
    outputs(11286) <= not((layer0_outputs(1701)) xor (layer0_outputs(779)));
    outputs(11287) <= not(layer0_outputs(11767)) or (layer0_outputs(381));
    outputs(11288) <= (layer0_outputs(11542)) xor (layer0_outputs(7239));
    outputs(11289) <= not((layer0_outputs(9022)) xor (layer0_outputs(10999)));
    outputs(11290) <= not(layer0_outputs(8254));
    outputs(11291) <= not((layer0_outputs(6627)) xor (layer0_outputs(119)));
    outputs(11292) <= layer0_outputs(12582);
    outputs(11293) <= layer0_outputs(1827);
    outputs(11294) <= (layer0_outputs(8341)) and not (layer0_outputs(8542));
    outputs(11295) <= not((layer0_outputs(7637)) or (layer0_outputs(1929)));
    outputs(11296) <= (layer0_outputs(1561)) and not (layer0_outputs(8642));
    outputs(11297) <= not((layer0_outputs(169)) xor (layer0_outputs(160)));
    outputs(11298) <= (layer0_outputs(7791)) xor (layer0_outputs(5143));
    outputs(11299) <= layer0_outputs(9458);
    outputs(11300) <= not(layer0_outputs(12279));
    outputs(11301) <= (layer0_outputs(5039)) and not (layer0_outputs(7208));
    outputs(11302) <= not(layer0_outputs(2709));
    outputs(11303) <= not(layer0_outputs(6716)) or (layer0_outputs(12689));
    outputs(11304) <= (layer0_outputs(10570)) xor (layer0_outputs(3895));
    outputs(11305) <= layer0_outputs(10967);
    outputs(11306) <= layer0_outputs(3542);
    outputs(11307) <= layer0_outputs(2601);
    outputs(11308) <= (layer0_outputs(4797)) xor (layer0_outputs(3671));
    outputs(11309) <= not(layer0_outputs(6439));
    outputs(11310) <= not((layer0_outputs(1)) xor (layer0_outputs(6911)));
    outputs(11311) <= layer0_outputs(4852);
    outputs(11312) <= layer0_outputs(2858);
    outputs(11313) <= (layer0_outputs(4087)) or (layer0_outputs(36));
    outputs(11314) <= not(layer0_outputs(1429)) or (layer0_outputs(7129));
    outputs(11315) <= (layer0_outputs(12452)) and not (layer0_outputs(5587));
    outputs(11316) <= layer0_outputs(1049);
    outputs(11317) <= not(layer0_outputs(12324));
    outputs(11318) <= not(layer0_outputs(12545));
    outputs(11319) <= not((layer0_outputs(9519)) xor (layer0_outputs(3664)));
    outputs(11320) <= not(layer0_outputs(10453)) or (layer0_outputs(8315));
    outputs(11321) <= not((layer0_outputs(4412)) xor (layer0_outputs(5507)));
    outputs(11322) <= not(layer0_outputs(7734));
    outputs(11323) <= (layer0_outputs(2547)) xor (layer0_outputs(3707));
    outputs(11324) <= (layer0_outputs(11721)) xor (layer0_outputs(5727));
    outputs(11325) <= not(layer0_outputs(516));
    outputs(11326) <= (layer0_outputs(5472)) and not (layer0_outputs(6455));
    outputs(11327) <= not((layer0_outputs(9423)) xor (layer0_outputs(4622)));
    outputs(11328) <= not((layer0_outputs(1156)) xor (layer0_outputs(2069)));
    outputs(11329) <= not((layer0_outputs(811)) xor (layer0_outputs(7302)));
    outputs(11330) <= not(layer0_outputs(5026)) or (layer0_outputs(10021));
    outputs(11331) <= (layer0_outputs(5989)) or (layer0_outputs(10585));
    outputs(11332) <= (layer0_outputs(6148)) xor (layer0_outputs(4837));
    outputs(11333) <= not((layer0_outputs(5997)) xor (layer0_outputs(859)));
    outputs(11334) <= layer0_outputs(10697);
    outputs(11335) <= not((layer0_outputs(11186)) xor (layer0_outputs(1664)));
    outputs(11336) <= not(layer0_outputs(9161));
    outputs(11337) <= not((layer0_outputs(11959)) and (layer0_outputs(2756)));
    outputs(11338) <= not(layer0_outputs(4146));
    outputs(11339) <= not(layer0_outputs(9384));
    outputs(11340) <= not((layer0_outputs(6587)) and (layer0_outputs(383)));
    outputs(11341) <= not(layer0_outputs(8505));
    outputs(11342) <= (layer0_outputs(11199)) or (layer0_outputs(5747));
    outputs(11343) <= (layer0_outputs(9458)) and not (layer0_outputs(2643));
    outputs(11344) <= not((layer0_outputs(8817)) and (layer0_outputs(8380)));
    outputs(11345) <= layer0_outputs(12446);
    outputs(11346) <= not(layer0_outputs(2111));
    outputs(11347) <= (layer0_outputs(1534)) and not (layer0_outputs(7339));
    outputs(11348) <= layer0_outputs(2759);
    outputs(11349) <= not(layer0_outputs(8432));
    outputs(11350) <= (layer0_outputs(8922)) or (layer0_outputs(10371));
    outputs(11351) <= not((layer0_outputs(3715)) xor (layer0_outputs(10046)));
    outputs(11352) <= layer0_outputs(1626);
    outputs(11353) <= not((layer0_outputs(1594)) xor (layer0_outputs(8683)));
    outputs(11354) <= not(layer0_outputs(1254));
    outputs(11355) <= layer0_outputs(209);
    outputs(11356) <= layer0_outputs(3220);
    outputs(11357) <= (layer0_outputs(8517)) xor (layer0_outputs(9653));
    outputs(11358) <= not(layer0_outputs(3939)) or (layer0_outputs(7736));
    outputs(11359) <= (layer0_outputs(6570)) xor (layer0_outputs(4369));
    outputs(11360) <= not((layer0_outputs(7812)) xor (layer0_outputs(348)));
    outputs(11361) <= not(layer0_outputs(9922));
    outputs(11362) <= not((layer0_outputs(5197)) xor (layer0_outputs(7203)));
    outputs(11363) <= '1';
    outputs(11364) <= not(layer0_outputs(7991));
    outputs(11365) <= (layer0_outputs(11710)) and not (layer0_outputs(11991));
    outputs(11366) <= not(layer0_outputs(3408));
    outputs(11367) <= layer0_outputs(5807);
    outputs(11368) <= layer0_outputs(4023);
    outputs(11369) <= (layer0_outputs(2119)) xor (layer0_outputs(4272));
    outputs(11370) <= not((layer0_outputs(5934)) xor (layer0_outputs(646)));
    outputs(11371) <= not((layer0_outputs(2415)) xor (layer0_outputs(11213)));
    outputs(11372) <= not(layer0_outputs(1475)) or (layer0_outputs(606));
    outputs(11373) <= not(layer0_outputs(3434));
    outputs(11374) <= not((layer0_outputs(620)) xor (layer0_outputs(3888)));
    outputs(11375) <= not((layer0_outputs(5565)) xor (layer0_outputs(10880)));
    outputs(11376) <= layer0_outputs(9427);
    outputs(11377) <= not(layer0_outputs(3075)) or (layer0_outputs(3480));
    outputs(11378) <= not((layer0_outputs(9324)) or (layer0_outputs(3572)));
    outputs(11379) <= not((layer0_outputs(10736)) xor (layer0_outputs(9004)));
    outputs(11380) <= layer0_outputs(11875);
    outputs(11381) <= not((layer0_outputs(5015)) and (layer0_outputs(2792)));
    outputs(11382) <= (layer0_outputs(11932)) xor (layer0_outputs(287));
    outputs(11383) <= layer0_outputs(4585);
    outputs(11384) <= not(layer0_outputs(1294));
    outputs(11385) <= (layer0_outputs(7000)) and not (layer0_outputs(2612));
    outputs(11386) <= not((layer0_outputs(6302)) and (layer0_outputs(541)));
    outputs(11387) <= (layer0_outputs(6592)) and not (layer0_outputs(10460));
    outputs(11388) <= not((layer0_outputs(1836)) or (layer0_outputs(7403)));
    outputs(11389) <= not(layer0_outputs(11965));
    outputs(11390) <= (layer0_outputs(4963)) xor (layer0_outputs(5293));
    outputs(11391) <= not((layer0_outputs(4903)) and (layer0_outputs(3221)));
    outputs(11392) <= layer0_outputs(61);
    outputs(11393) <= not((layer0_outputs(5836)) xor (layer0_outputs(4170)));
    outputs(11394) <= (layer0_outputs(122)) xor (layer0_outputs(2499));
    outputs(11395) <= not(layer0_outputs(56));
    outputs(11396) <= not(layer0_outputs(2570));
    outputs(11397) <= not((layer0_outputs(2288)) xor (layer0_outputs(9616)));
    outputs(11398) <= not(layer0_outputs(11));
    outputs(11399) <= not(layer0_outputs(2379)) or (layer0_outputs(7534));
    outputs(11400) <= (layer0_outputs(6891)) or (layer0_outputs(5381));
    outputs(11401) <= not(layer0_outputs(1843));
    outputs(11402) <= (layer0_outputs(11416)) xor (layer0_outputs(509));
    outputs(11403) <= layer0_outputs(8458);
    outputs(11404) <= layer0_outputs(4776);
    outputs(11405) <= layer0_outputs(9245);
    outputs(11406) <= not((layer0_outputs(10491)) and (layer0_outputs(6219)));
    outputs(11407) <= (layer0_outputs(1344)) xor (layer0_outputs(4313));
    outputs(11408) <= layer0_outputs(164);
    outputs(11409) <= not(layer0_outputs(3145)) or (layer0_outputs(11643));
    outputs(11410) <= (layer0_outputs(1250)) xor (layer0_outputs(558));
    outputs(11411) <= (layer0_outputs(10032)) or (layer0_outputs(8544));
    outputs(11412) <= not(layer0_outputs(11224)) or (layer0_outputs(5379));
    outputs(11413) <= not(layer0_outputs(2624)) or (layer0_outputs(143));
    outputs(11414) <= (layer0_outputs(3984)) xor (layer0_outputs(4335));
    outputs(11415) <= (layer0_outputs(10340)) xor (layer0_outputs(4323));
    outputs(11416) <= not((layer0_outputs(6382)) xor (layer0_outputs(11943)));
    outputs(11417) <= layer0_outputs(398);
    outputs(11418) <= not(layer0_outputs(6766));
    outputs(11419) <= not(layer0_outputs(2353));
    outputs(11420) <= not((layer0_outputs(920)) xor (layer0_outputs(12665)));
    outputs(11421) <= not(layer0_outputs(6609));
    outputs(11422) <= (layer0_outputs(12256)) or (layer0_outputs(4663));
    outputs(11423) <= (layer0_outputs(1762)) xor (layer0_outputs(12491));
    outputs(11424) <= not((layer0_outputs(7010)) and (layer0_outputs(5272)));
    outputs(11425) <= (layer0_outputs(1398)) xor (layer0_outputs(11601));
    outputs(11426) <= layer0_outputs(6561);
    outputs(11427) <= layer0_outputs(161);
    outputs(11428) <= layer0_outputs(6119);
    outputs(11429) <= not((layer0_outputs(2590)) xor (layer0_outputs(1995)));
    outputs(11430) <= not(layer0_outputs(2696));
    outputs(11431) <= layer0_outputs(4807);
    outputs(11432) <= not(layer0_outputs(308)) or (layer0_outputs(9613));
    outputs(11433) <= layer0_outputs(12643);
    outputs(11434) <= not((layer0_outputs(5716)) and (layer0_outputs(313)));
    outputs(11435) <= not((layer0_outputs(3522)) and (layer0_outputs(2263)));
    outputs(11436) <= not((layer0_outputs(11257)) or (layer0_outputs(4238)));
    outputs(11437) <= (layer0_outputs(3722)) xor (layer0_outputs(8084));
    outputs(11438) <= not((layer0_outputs(7577)) xor (layer0_outputs(3150)));
    outputs(11439) <= (layer0_outputs(6633)) or (layer0_outputs(6487));
    outputs(11440) <= (layer0_outputs(5393)) xor (layer0_outputs(2123));
    outputs(11441) <= layer0_outputs(5623);
    outputs(11442) <= not((layer0_outputs(11752)) xor (layer0_outputs(1844)));
    outputs(11443) <= layer0_outputs(8217);
    outputs(11444) <= layer0_outputs(12515);
    outputs(11445) <= not(layer0_outputs(4716));
    outputs(11446) <= layer0_outputs(6164);
    outputs(11447) <= (layer0_outputs(1990)) and not (layer0_outputs(8796));
    outputs(11448) <= layer0_outputs(6288);
    outputs(11449) <= (layer0_outputs(316)) and not (layer0_outputs(9944));
    outputs(11450) <= layer0_outputs(193);
    outputs(11451) <= (layer0_outputs(8498)) xor (layer0_outputs(9945));
    outputs(11452) <= (layer0_outputs(1799)) xor (layer0_outputs(1443));
    outputs(11453) <= not((layer0_outputs(12609)) xor (layer0_outputs(4496)));
    outputs(11454) <= layer0_outputs(8805);
    outputs(11455) <= not(layer0_outputs(1607));
    outputs(11456) <= not((layer0_outputs(3421)) xor (layer0_outputs(242)));
    outputs(11457) <= layer0_outputs(7917);
    outputs(11458) <= layer0_outputs(10910);
    outputs(11459) <= not((layer0_outputs(3952)) xor (layer0_outputs(8575)));
    outputs(11460) <= (layer0_outputs(9841)) xor (layer0_outputs(12020));
    outputs(11461) <= (layer0_outputs(994)) xor (layer0_outputs(10789));
    outputs(11462) <= (layer0_outputs(9409)) or (layer0_outputs(6882));
    outputs(11463) <= not(layer0_outputs(1073)) or (layer0_outputs(6159));
    outputs(11464) <= not(layer0_outputs(4816));
    outputs(11465) <= not(layer0_outputs(10018)) or (layer0_outputs(65));
    outputs(11466) <= not((layer0_outputs(5249)) xor (layer0_outputs(3055)));
    outputs(11467) <= not(layer0_outputs(1003));
    outputs(11468) <= not(layer0_outputs(52)) or (layer0_outputs(1047));
    outputs(11469) <= layer0_outputs(8569);
    outputs(11470) <= '1';
    outputs(11471) <= layer0_outputs(4939);
    outputs(11472) <= not((layer0_outputs(8034)) xor (layer0_outputs(6250)));
    outputs(11473) <= not((layer0_outputs(4247)) xor (layer0_outputs(9985)));
    outputs(11474) <= not((layer0_outputs(11324)) xor (layer0_outputs(6840)));
    outputs(11475) <= (layer0_outputs(12697)) xor (layer0_outputs(11857));
    outputs(11476) <= not((layer0_outputs(3554)) xor (layer0_outputs(4000)));
    outputs(11477) <= not((layer0_outputs(8873)) and (layer0_outputs(7323)));
    outputs(11478) <= not((layer0_outputs(241)) and (layer0_outputs(7223)));
    outputs(11479) <= layer0_outputs(1716);
    outputs(11480) <= not(layer0_outputs(7483));
    outputs(11481) <= not((layer0_outputs(11108)) and (layer0_outputs(7052)));
    outputs(11482) <= not(layer0_outputs(11404));
    outputs(11483) <= (layer0_outputs(69)) or (layer0_outputs(11089));
    outputs(11484) <= (layer0_outputs(3864)) xor (layer0_outputs(7579));
    outputs(11485) <= not(layer0_outputs(783)) or (layer0_outputs(5576));
    outputs(11486) <= not((layer0_outputs(3759)) and (layer0_outputs(3316)));
    outputs(11487) <= not((layer0_outputs(7371)) xor (layer0_outputs(6678)));
    outputs(11488) <= not(layer0_outputs(12076));
    outputs(11489) <= (layer0_outputs(9055)) and not (layer0_outputs(1299));
    outputs(11490) <= not(layer0_outputs(4311));
    outputs(11491) <= not(layer0_outputs(5207)) or (layer0_outputs(3523));
    outputs(11492) <= not((layer0_outputs(11426)) xor (layer0_outputs(3972)));
    outputs(11493) <= layer0_outputs(1405);
    outputs(11494) <= not(layer0_outputs(4360)) or (layer0_outputs(11183));
    outputs(11495) <= (layer0_outputs(12655)) xor (layer0_outputs(9795));
    outputs(11496) <= layer0_outputs(7821);
    outputs(11497) <= layer0_outputs(7772);
    outputs(11498) <= not(layer0_outputs(6755));
    outputs(11499) <= layer0_outputs(9652);
    outputs(11500) <= not(layer0_outputs(7873));
    outputs(11501) <= not((layer0_outputs(1993)) or (layer0_outputs(7604)));
    outputs(11502) <= not((layer0_outputs(10430)) xor (layer0_outputs(12134)));
    outputs(11503) <= not(layer0_outputs(6994));
    outputs(11504) <= not((layer0_outputs(10157)) xor (layer0_outputs(2636)));
    outputs(11505) <= (layer0_outputs(2162)) xor (layer0_outputs(8770));
    outputs(11506) <= not(layer0_outputs(8259)) or (layer0_outputs(4072));
    outputs(11507) <= not((layer0_outputs(5370)) or (layer0_outputs(1497)));
    outputs(11508) <= not(layer0_outputs(8985));
    outputs(11509) <= not(layer0_outputs(3411));
    outputs(11510) <= (layer0_outputs(2185)) xor (layer0_outputs(6350));
    outputs(11511) <= layer0_outputs(3061);
    outputs(11512) <= not(layer0_outputs(1733)) or (layer0_outputs(9352));
    outputs(11513) <= (layer0_outputs(8520)) and (layer0_outputs(12501));
    outputs(11514) <= not(layer0_outputs(7513));
    outputs(11515) <= (layer0_outputs(6001)) or (layer0_outputs(7006));
    outputs(11516) <= not((layer0_outputs(2881)) xor (layer0_outputs(2460)));
    outputs(11517) <= (layer0_outputs(6037)) xor (layer0_outputs(11628));
    outputs(11518) <= not((layer0_outputs(7236)) and (layer0_outputs(4931)));
    outputs(11519) <= (layer0_outputs(290)) and not (layer0_outputs(6618));
    outputs(11520) <= not(layer0_outputs(7434));
    outputs(11521) <= not(layer0_outputs(1830));
    outputs(11522) <= not((layer0_outputs(7605)) xor (layer0_outputs(8117)));
    outputs(11523) <= (layer0_outputs(1502)) and not (layer0_outputs(9928));
    outputs(11524) <= not(layer0_outputs(6821)) or (layer0_outputs(200));
    outputs(11525) <= not((layer0_outputs(3205)) xor (layer0_outputs(2800)));
    outputs(11526) <= layer0_outputs(8697);
    outputs(11527) <= layer0_outputs(3138);
    outputs(11528) <= (layer0_outputs(10975)) xor (layer0_outputs(9363));
    outputs(11529) <= not((layer0_outputs(4214)) and (layer0_outputs(1876)));
    outputs(11530) <= not(layer0_outputs(12311));
    outputs(11531) <= not((layer0_outputs(3866)) and (layer0_outputs(2174)));
    outputs(11532) <= not(layer0_outputs(12357));
    outputs(11533) <= layer0_outputs(11362);
    outputs(11534) <= (layer0_outputs(7757)) xor (layer0_outputs(2077));
    outputs(11535) <= (layer0_outputs(2070)) xor (layer0_outputs(6097));
    outputs(11536) <= layer0_outputs(3711);
    outputs(11537) <= not(layer0_outputs(670)) or (layer0_outputs(3896));
    outputs(11538) <= not((layer0_outputs(3237)) xor (layer0_outputs(10535)));
    outputs(11539) <= (layer0_outputs(4376)) xor (layer0_outputs(5879));
    outputs(11540) <= (layer0_outputs(11302)) xor (layer0_outputs(7267));
    outputs(11541) <= not((layer0_outputs(2438)) xor (layer0_outputs(6768)));
    outputs(11542) <= layer0_outputs(844);
    outputs(11543) <= (layer0_outputs(8698)) xor (layer0_outputs(8704));
    outputs(11544) <= not(layer0_outputs(7103));
    outputs(11545) <= not(layer0_outputs(6302));
    outputs(11546) <= not((layer0_outputs(9333)) xor (layer0_outputs(11848)));
    outputs(11547) <= not((layer0_outputs(9878)) xor (layer0_outputs(9016)));
    outputs(11548) <= not((layer0_outputs(7506)) xor (layer0_outputs(11960)));
    outputs(11549) <= not(layer0_outputs(1739));
    outputs(11550) <= layer0_outputs(2928);
    outputs(11551) <= (layer0_outputs(12554)) xor (layer0_outputs(7943));
    outputs(11552) <= not((layer0_outputs(3166)) xor (layer0_outputs(11053)));
    outputs(11553) <= (layer0_outputs(5513)) and not (layer0_outputs(8079));
    outputs(11554) <= layer0_outputs(8447);
    outputs(11555) <= not(layer0_outputs(2052));
    outputs(11556) <= not((layer0_outputs(1140)) xor (layer0_outputs(8533)));
    outputs(11557) <= (layer0_outputs(9802)) xor (layer0_outputs(9502));
    outputs(11558) <= not((layer0_outputs(4383)) xor (layer0_outputs(11854)));
    outputs(11559) <= (layer0_outputs(4754)) xor (layer0_outputs(10117));
    outputs(11560) <= (layer0_outputs(4608)) or (layer0_outputs(8982));
    outputs(11561) <= (layer0_outputs(3001)) and not (layer0_outputs(742));
    outputs(11562) <= not(layer0_outputs(536));
    outputs(11563) <= not(layer0_outputs(3291));
    outputs(11564) <= not(layer0_outputs(8771));
    outputs(11565) <= not(layer0_outputs(6046));
    outputs(11566) <= not((layer0_outputs(2820)) xor (layer0_outputs(6007)));
    outputs(11567) <= not((layer0_outputs(9560)) and (layer0_outputs(5071)));
    outputs(11568) <= layer0_outputs(2027);
    outputs(11569) <= not(layer0_outputs(511));
    outputs(11570) <= layer0_outputs(4909);
    outputs(11571) <= (layer0_outputs(5634)) or (layer0_outputs(6351));
    outputs(11572) <= not((layer0_outputs(9522)) xor (layer0_outputs(9932)));
    outputs(11573) <= not(layer0_outputs(6580));
    outputs(11574) <= (layer0_outputs(622)) xor (layer0_outputs(2465));
    outputs(11575) <= not(layer0_outputs(8784));
    outputs(11576) <= not((layer0_outputs(8481)) or (layer0_outputs(1536)));
    outputs(11577) <= (layer0_outputs(8272)) and not (layer0_outputs(12376));
    outputs(11578) <= not((layer0_outputs(4282)) xor (layer0_outputs(4068)));
    outputs(11579) <= not((layer0_outputs(10294)) xor (layer0_outputs(8530)));
    outputs(11580) <= layer0_outputs(3903);
    outputs(11581) <= (layer0_outputs(9860)) and not (layer0_outputs(778));
    outputs(11582) <= not((layer0_outputs(4160)) xor (layer0_outputs(9593)));
    outputs(11583) <= not(layer0_outputs(11532));
    outputs(11584) <= (layer0_outputs(5073)) xor (layer0_outputs(11835));
    outputs(11585) <= layer0_outputs(4167);
    outputs(11586) <= (layer0_outputs(9307)) xor (layer0_outputs(2694));
    outputs(11587) <= not((layer0_outputs(3727)) xor (layer0_outputs(1563)));
    outputs(11588) <= (layer0_outputs(5676)) and not (layer0_outputs(6811));
    outputs(11589) <= not(layer0_outputs(10238));
    outputs(11590) <= (layer0_outputs(2319)) xor (layer0_outputs(3637));
    outputs(11591) <= not((layer0_outputs(11808)) xor (layer0_outputs(8092)));
    outputs(11592) <= not((layer0_outputs(5792)) or (layer0_outputs(6055)));
    outputs(11593) <= (layer0_outputs(4038)) and (layer0_outputs(9013));
    outputs(11594) <= not((layer0_outputs(12246)) xor (layer0_outputs(6215)));
    outputs(11595) <= not(layer0_outputs(5683));
    outputs(11596) <= (layer0_outputs(2511)) or (layer0_outputs(6130));
    outputs(11597) <= not((layer0_outputs(3484)) xor (layer0_outputs(11900)));
    outputs(11598) <= layer0_outputs(1511);
    outputs(11599) <= layer0_outputs(6453);
    outputs(11600) <= layer0_outputs(3752);
    outputs(11601) <= not((layer0_outputs(9693)) xor (layer0_outputs(5139)));
    outputs(11602) <= (layer0_outputs(10224)) xor (layer0_outputs(8244));
    outputs(11603) <= layer0_outputs(4984);
    outputs(11604) <= (layer0_outputs(7303)) and (layer0_outputs(9337));
    outputs(11605) <= layer0_outputs(11031);
    outputs(11606) <= not(layer0_outputs(4377));
    outputs(11607) <= (layer0_outputs(5348)) xor (layer0_outputs(7279));
    outputs(11608) <= layer0_outputs(46);
    outputs(11609) <= layer0_outputs(5197);
    outputs(11610) <= (layer0_outputs(1625)) xor (layer0_outputs(6687));
    outputs(11611) <= (layer0_outputs(12463)) xor (layer0_outputs(12710));
    outputs(11612) <= (layer0_outputs(11672)) and not (layer0_outputs(10644));
    outputs(11613) <= (layer0_outputs(4937)) and not (layer0_outputs(9692));
    outputs(11614) <= not((layer0_outputs(3808)) xor (layer0_outputs(9597)));
    outputs(11615) <= layer0_outputs(5129);
    outputs(11616) <= not(layer0_outputs(11261)) or (layer0_outputs(5910));
    outputs(11617) <= not((layer0_outputs(5939)) xor (layer0_outputs(12176)));
    outputs(11618) <= not(layer0_outputs(4345));
    outputs(11619) <= not(layer0_outputs(11860));
    outputs(11620) <= not(layer0_outputs(3068));
    outputs(11621) <= not((layer0_outputs(7387)) xor (layer0_outputs(12196)));
    outputs(11622) <= (layer0_outputs(12227)) and not (layer0_outputs(1156));
    outputs(11623) <= (layer0_outputs(5670)) xor (layer0_outputs(3385));
    outputs(11624) <= layer0_outputs(429);
    outputs(11625) <= not((layer0_outputs(8197)) or (layer0_outputs(5796)));
    outputs(11626) <= not(layer0_outputs(2945));
    outputs(11627) <= layer0_outputs(5604);
    outputs(11628) <= not(layer0_outputs(12666));
    outputs(11629) <= (layer0_outputs(800)) xor (layer0_outputs(4152));
    outputs(11630) <= layer0_outputs(7274);
    outputs(11631) <= not(layer0_outputs(101));
    outputs(11632) <= (layer0_outputs(1155)) and not (layer0_outputs(3526));
    outputs(11633) <= not(layer0_outputs(7240));
    outputs(11634) <= not((layer0_outputs(3570)) xor (layer0_outputs(2608)));
    outputs(11635) <= not((layer0_outputs(7908)) or (layer0_outputs(347)));
    outputs(11636) <= (layer0_outputs(11406)) xor (layer0_outputs(2401));
    outputs(11637) <= (layer0_outputs(2292)) xor (layer0_outputs(8486));
    outputs(11638) <= not((layer0_outputs(1951)) xor (layer0_outputs(12077)));
    outputs(11639) <= not(layer0_outputs(9675)) or (layer0_outputs(3194));
    outputs(11640) <= (layer0_outputs(6083)) xor (layer0_outputs(4687));
    outputs(11641) <= not(layer0_outputs(1040));
    outputs(11642) <= not(layer0_outputs(578));
    outputs(11643) <= not(layer0_outputs(9088));
    outputs(11644) <= not(layer0_outputs(10078));
    outputs(11645) <= layer0_outputs(7159);
    outputs(11646) <= (layer0_outputs(12790)) or (layer0_outputs(5959));
    outputs(11647) <= not((layer0_outputs(1764)) xor (layer0_outputs(10256)));
    outputs(11648) <= layer0_outputs(3328);
    outputs(11649) <= not(layer0_outputs(8855));
    outputs(11650) <= layer0_outputs(8239);
    outputs(11651) <= (layer0_outputs(6364)) and not (layer0_outputs(6010));
    outputs(11652) <= not((layer0_outputs(7799)) xor (layer0_outputs(9810)));
    outputs(11653) <= layer0_outputs(9868);
    outputs(11654) <= (layer0_outputs(6102)) and (layer0_outputs(7315));
    outputs(11655) <= not(layer0_outputs(6246));
    outputs(11656) <= not((layer0_outputs(8148)) and (layer0_outputs(1278)));
    outputs(11657) <= (layer0_outputs(10087)) xor (layer0_outputs(7455));
    outputs(11658) <= (layer0_outputs(8669)) or (layer0_outputs(11601));
    outputs(11659) <= not((layer0_outputs(11336)) xor (layer0_outputs(1109)));
    outputs(11660) <= not((layer0_outputs(10218)) xor (layer0_outputs(649)));
    outputs(11661) <= (layer0_outputs(5927)) xor (layer0_outputs(5834));
    outputs(11662) <= not((layer0_outputs(9804)) or (layer0_outputs(6886)));
    outputs(11663) <= (layer0_outputs(12403)) xor (layer0_outputs(2973));
    outputs(11664) <= not(layer0_outputs(4143));
    outputs(11665) <= layer0_outputs(520);
    outputs(11666) <= (layer0_outputs(9995)) and not (layer0_outputs(7375));
    outputs(11667) <= (layer0_outputs(8124)) xor (layer0_outputs(10292));
    outputs(11668) <= not((layer0_outputs(10890)) xor (layer0_outputs(2935)));
    outputs(11669) <= (layer0_outputs(10818)) and (layer0_outputs(230));
    outputs(11670) <= not((layer0_outputs(11540)) and (layer0_outputs(11346)));
    outputs(11671) <= (layer0_outputs(2236)) and (layer0_outputs(10113));
    outputs(11672) <= not(layer0_outputs(8304));
    outputs(11673) <= layer0_outputs(3934);
    outputs(11674) <= layer0_outputs(10065);
    outputs(11675) <= layer0_outputs(5687);
    outputs(11676) <= (layer0_outputs(3386)) xor (layer0_outputs(549));
    outputs(11677) <= (layer0_outputs(10982)) xor (layer0_outputs(12439));
    outputs(11678) <= (layer0_outputs(6282)) xor (layer0_outputs(7729));
    outputs(11679) <= not((layer0_outputs(6826)) and (layer0_outputs(6253)));
    outputs(11680) <= not(layer0_outputs(11073)) or (layer0_outputs(1355));
    outputs(11681) <= (layer0_outputs(2088)) xor (layer0_outputs(9361));
    outputs(11682) <= (layer0_outputs(1426)) and not (layer0_outputs(9232));
    outputs(11683) <= layer0_outputs(8401);
    outputs(11684) <= (layer0_outputs(10105)) and not (layer0_outputs(12738));
    outputs(11685) <= (layer0_outputs(7508)) xor (layer0_outputs(10382));
    outputs(11686) <= layer0_outputs(11375);
    outputs(11687) <= not(layer0_outputs(3521));
    outputs(11688) <= (layer0_outputs(82)) and not (layer0_outputs(10050));
    outputs(11689) <= not((layer0_outputs(9456)) xor (layer0_outputs(1280)));
    outputs(11690) <= layer0_outputs(5248);
    outputs(11691) <= (layer0_outputs(11446)) xor (layer0_outputs(4152));
    outputs(11692) <= (layer0_outputs(2224)) and not (layer0_outputs(751));
    outputs(11693) <= not(layer0_outputs(7323));
    outputs(11694) <= (layer0_outputs(7916)) xor (layer0_outputs(2967));
    outputs(11695) <= layer0_outputs(3347);
    outputs(11696) <= layer0_outputs(1490);
    outputs(11697) <= (layer0_outputs(3838)) and (layer0_outputs(5130));
    outputs(11698) <= layer0_outputs(7194);
    outputs(11699) <= (layer0_outputs(9116)) and not (layer0_outputs(1588));
    outputs(11700) <= (layer0_outputs(10732)) and not (layer0_outputs(1283));
    outputs(11701) <= not(layer0_outputs(835)) or (layer0_outputs(9455));
    outputs(11702) <= (layer0_outputs(9315)) and not (layer0_outputs(11952));
    outputs(11703) <= layer0_outputs(3882);
    outputs(11704) <= not((layer0_outputs(11531)) xor (layer0_outputs(6958)));
    outputs(11705) <= layer0_outputs(3849);
    outputs(11706) <= not((layer0_outputs(669)) or (layer0_outputs(7877)));
    outputs(11707) <= layer0_outputs(3229);
    outputs(11708) <= not((layer0_outputs(3356)) xor (layer0_outputs(2778)));
    outputs(11709) <= not((layer0_outputs(3148)) xor (layer0_outputs(2009)));
    outputs(11710) <= not(layer0_outputs(3122));
    outputs(11711) <= (layer0_outputs(5962)) xor (layer0_outputs(12433));
    outputs(11712) <= layer0_outputs(6526);
    outputs(11713) <= not(layer0_outputs(8955));
    outputs(11714) <= not(layer0_outputs(8816));
    outputs(11715) <= not(layer0_outputs(2325)) or (layer0_outputs(11999));
    outputs(11716) <= not(layer0_outputs(10220));
    outputs(11717) <= not(layer0_outputs(6166));
    outputs(11718) <= (layer0_outputs(10529)) and (layer0_outputs(719));
    outputs(11719) <= (layer0_outputs(1900)) xor (layer0_outputs(383));
    outputs(11720) <= not((layer0_outputs(3538)) or (layer0_outputs(2082)));
    outputs(11721) <= layer0_outputs(5672);
    outputs(11722) <= (layer0_outputs(7954)) xor (layer0_outputs(852));
    outputs(11723) <= (layer0_outputs(7131)) and (layer0_outputs(8476));
    outputs(11724) <= (layer0_outputs(6070)) xor (layer0_outputs(60));
    outputs(11725) <= not((layer0_outputs(727)) xor (layer0_outputs(11128)));
    outputs(11726) <= (layer0_outputs(1803)) xor (layer0_outputs(5091));
    outputs(11727) <= not((layer0_outputs(7869)) xor (layer0_outputs(5972)));
    outputs(11728) <= (layer0_outputs(6553)) xor (layer0_outputs(10357));
    outputs(11729) <= not(layer0_outputs(424));
    outputs(11730) <= (layer0_outputs(1459)) xor (layer0_outputs(11594));
    outputs(11731) <= layer0_outputs(9623);
    outputs(11732) <= layer0_outputs(12276);
    outputs(11733) <= (layer0_outputs(9367)) and not (layer0_outputs(773));
    outputs(11734) <= not((layer0_outputs(3703)) xor (layer0_outputs(1474)));
    outputs(11735) <= (layer0_outputs(1576)) xor (layer0_outputs(2665));
    outputs(11736) <= not(layer0_outputs(3412));
    outputs(11737) <= not(layer0_outputs(3195));
    outputs(11738) <= (layer0_outputs(5882)) and not (layer0_outputs(8028));
    outputs(11739) <= (layer0_outputs(12125)) and not (layer0_outputs(4711));
    outputs(11740) <= not(layer0_outputs(2339));
    outputs(11741) <= not(layer0_outputs(1508)) or (layer0_outputs(4436));
    outputs(11742) <= not((layer0_outputs(11136)) and (layer0_outputs(9624)));
    outputs(11743) <= not((layer0_outputs(11338)) xor (layer0_outputs(5608)));
    outputs(11744) <= not(layer0_outputs(2455));
    outputs(11745) <= not(layer0_outputs(5678));
    outputs(11746) <= (layer0_outputs(3916)) xor (layer0_outputs(12716));
    outputs(11747) <= (layer0_outputs(5757)) or (layer0_outputs(10881));
    outputs(11748) <= layer0_outputs(10113);
    outputs(11749) <= (layer0_outputs(11790)) and (layer0_outputs(5122));
    outputs(11750) <= (layer0_outputs(11605)) xor (layer0_outputs(6767));
    outputs(11751) <= not(layer0_outputs(9611));
    outputs(11752) <= not((layer0_outputs(12084)) xor (layer0_outputs(5399)));
    outputs(11753) <= not(layer0_outputs(12658));
    outputs(11754) <= not(layer0_outputs(8539));
    outputs(11755) <= not((layer0_outputs(809)) xor (layer0_outputs(8410)));
    outputs(11756) <= (layer0_outputs(3246)) xor (layer0_outputs(7751));
    outputs(11757) <= layer0_outputs(11012);
    outputs(11758) <= not(layer0_outputs(1548));
    outputs(11759) <= (layer0_outputs(10139)) xor (layer0_outputs(8633));
    outputs(11760) <= not(layer0_outputs(7199)) or (layer0_outputs(4155));
    outputs(11761) <= not(layer0_outputs(6531)) or (layer0_outputs(4289));
    outputs(11762) <= (layer0_outputs(11585)) xor (layer0_outputs(11171));
    outputs(11763) <= (layer0_outputs(9767)) and not (layer0_outputs(895));
    outputs(11764) <= not((layer0_outputs(436)) or (layer0_outputs(6550)));
    outputs(11765) <= layer0_outputs(10230);
    outputs(11766) <= layer0_outputs(9939);
    outputs(11767) <= (layer0_outputs(1896)) and not (layer0_outputs(4701));
    outputs(11768) <= not(layer0_outputs(5769));
    outputs(11769) <= not(layer0_outputs(2566));
    outputs(11770) <= (layer0_outputs(3182)) xor (layer0_outputs(10359));
    outputs(11771) <= layer0_outputs(4489);
    outputs(11772) <= not((layer0_outputs(11500)) or (layer0_outputs(4568)));
    outputs(11773) <= not((layer0_outputs(5964)) xor (layer0_outputs(7509)));
    outputs(11774) <= layer0_outputs(6162);
    outputs(11775) <= not((layer0_outputs(8198)) xor (layer0_outputs(10830)));
    outputs(11776) <= (layer0_outputs(6107)) and not (layer0_outputs(12502));
    outputs(11777) <= (layer0_outputs(3098)) and not (layer0_outputs(2638));
    outputs(11778) <= (layer0_outputs(11350)) xor (layer0_outputs(8803));
    outputs(11779) <= (layer0_outputs(9426)) xor (layer0_outputs(12697));
    outputs(11780) <= not(layer0_outputs(6875)) or (layer0_outputs(2734));
    outputs(11781) <= not(layer0_outputs(500));
    outputs(11782) <= layer0_outputs(5377);
    outputs(11783) <= (layer0_outputs(10201)) xor (layer0_outputs(8752));
    outputs(11784) <= not(layer0_outputs(3786));
    outputs(11785) <= (layer0_outputs(9723)) and not (layer0_outputs(1648));
    outputs(11786) <= not((layer0_outputs(12634)) or (layer0_outputs(10720)));
    outputs(11787) <= not(layer0_outputs(12226));
    outputs(11788) <= (layer0_outputs(5131)) xor (layer0_outputs(11979));
    outputs(11789) <= layer0_outputs(5264);
    outputs(11790) <= layer0_outputs(9485);
    outputs(11791) <= not((layer0_outputs(9748)) xor (layer0_outputs(12008)));
    outputs(11792) <= not((layer0_outputs(10949)) xor (layer0_outputs(11759)));
    outputs(11793) <= not((layer0_outputs(9324)) xor (layer0_outputs(10456)));
    outputs(11794) <= not((layer0_outputs(11259)) xor (layer0_outputs(4345)));
    outputs(11795) <= not(layer0_outputs(8594));
    outputs(11796) <= not(layer0_outputs(7182));
    outputs(11797) <= layer0_outputs(6126);
    outputs(11798) <= not((layer0_outputs(489)) xor (layer0_outputs(1274)));
    outputs(11799) <= layer0_outputs(10852);
    outputs(11800) <= layer0_outputs(8471);
    outputs(11801) <= not((layer0_outputs(11182)) or (layer0_outputs(2921)));
    outputs(11802) <= (layer0_outputs(793)) xor (layer0_outputs(9449));
    outputs(11803) <= (layer0_outputs(1549)) and not (layer0_outputs(97));
    outputs(11804) <= not((layer0_outputs(12245)) xor (layer0_outputs(2806)));
    outputs(11805) <= (layer0_outputs(1422)) and not (layer0_outputs(3110));
    outputs(11806) <= not((layer0_outputs(6777)) and (layer0_outputs(9585)));
    outputs(11807) <= (layer0_outputs(3341)) or (layer0_outputs(12160));
    outputs(11808) <= layer0_outputs(6241);
    outputs(11809) <= layer0_outputs(3136);
    outputs(11810) <= (layer0_outputs(8041)) and (layer0_outputs(6976));
    outputs(11811) <= (layer0_outputs(6645)) xor (layer0_outputs(7843));
    outputs(11812) <= not(layer0_outputs(8727)) or (layer0_outputs(7328));
    outputs(11813) <= not(layer0_outputs(1458));
    outputs(11814) <= (layer0_outputs(611)) and not (layer0_outputs(4148));
    outputs(11815) <= not(layer0_outputs(8015));
    outputs(11816) <= not((layer0_outputs(10172)) or (layer0_outputs(5498)));
    outputs(11817) <= (layer0_outputs(3564)) xor (layer0_outputs(12669));
    outputs(11818) <= (layer0_outputs(12241)) xor (layer0_outputs(6727));
    outputs(11819) <= not((layer0_outputs(6093)) xor (layer0_outputs(6855)));
    outputs(11820) <= not((layer0_outputs(7681)) xor (layer0_outputs(2144)));
    outputs(11821) <= layer0_outputs(4943);
    outputs(11822) <= layer0_outputs(5956);
    outputs(11823) <= not((layer0_outputs(561)) xor (layer0_outputs(11223)));
    outputs(11824) <= not(layer0_outputs(8799));
    outputs(11825) <= layer0_outputs(3116);
    outputs(11826) <= (layer0_outputs(10202)) and (layer0_outputs(3081));
    outputs(11827) <= not((layer0_outputs(5615)) or (layer0_outputs(6229)));
    outputs(11828) <= not((layer0_outputs(6470)) xor (layer0_outputs(12751)));
    outputs(11829) <= not((layer0_outputs(11486)) xor (layer0_outputs(11748)));
    outputs(11830) <= not((layer0_outputs(9276)) xor (layer0_outputs(7703)));
    outputs(11831) <= not(layer0_outputs(1822));
    outputs(11832) <= layer0_outputs(7418);
    outputs(11833) <= (layer0_outputs(11839)) xor (layer0_outputs(5109));
    outputs(11834) <= not(layer0_outputs(4246)) or (layer0_outputs(4566));
    outputs(11835) <= layer0_outputs(9789);
    outputs(11836) <= not(layer0_outputs(7540));
    outputs(11837) <= not(layer0_outputs(3786));
    outputs(11838) <= not(layer0_outputs(7811)) or (layer0_outputs(1805));
    outputs(11839) <= layer0_outputs(3249);
    outputs(11840) <= (layer0_outputs(5714)) xor (layer0_outputs(8212));
    outputs(11841) <= not(layer0_outputs(12743));
    outputs(11842) <= layer0_outputs(12396);
    outputs(11843) <= layer0_outputs(9517);
    outputs(11844) <= (layer0_outputs(11531)) and not (layer0_outputs(9879));
    outputs(11845) <= layer0_outputs(870);
    outputs(11846) <= (layer0_outputs(4688)) and (layer0_outputs(11371));
    outputs(11847) <= layer0_outputs(10953);
    outputs(11848) <= (layer0_outputs(8609)) and (layer0_outputs(2926));
    outputs(11849) <= not((layer0_outputs(8073)) or (layer0_outputs(10443)));
    outputs(11850) <= not((layer0_outputs(9718)) xor (layer0_outputs(4690)));
    outputs(11851) <= (layer0_outputs(11354)) and not (layer0_outputs(11922));
    outputs(11852) <= not((layer0_outputs(1885)) xor (layer0_outputs(6527)));
    outputs(11853) <= layer0_outputs(84);
    outputs(11854) <= (layer0_outputs(2866)) and (layer0_outputs(1245));
    outputs(11855) <= not(layer0_outputs(5115)) or (layer0_outputs(5658));
    outputs(11856) <= layer0_outputs(951);
    outputs(11857) <= (layer0_outputs(7867)) xor (layer0_outputs(4139));
    outputs(11858) <= (layer0_outputs(11792)) and (layer0_outputs(11712));
    outputs(11859) <= (layer0_outputs(3571)) xor (layer0_outputs(6618));
    outputs(11860) <= (layer0_outputs(7127)) xor (layer0_outputs(969));
    outputs(11861) <= not((layer0_outputs(12379)) xor (layer0_outputs(1715)));
    outputs(11862) <= (layer0_outputs(2482)) xor (layer0_outputs(8523));
    outputs(11863) <= layer0_outputs(12673);
    outputs(11864) <= layer0_outputs(2766);
    outputs(11865) <= not(layer0_outputs(8102)) or (layer0_outputs(10947));
    outputs(11866) <= (layer0_outputs(9144)) and (layer0_outputs(2576));
    outputs(11867) <= (layer0_outputs(1556)) and not (layer0_outputs(12638));
    outputs(11868) <= layer0_outputs(1188);
    outputs(11869) <= not(layer0_outputs(8635)) or (layer0_outputs(3216));
    outputs(11870) <= layer0_outputs(9114);
    outputs(11871) <= layer0_outputs(9395);
    outputs(11872) <= not((layer0_outputs(11189)) or (layer0_outputs(5536)));
    outputs(11873) <= not(layer0_outputs(2183));
    outputs(11874) <= (layer0_outputs(4030)) and not (layer0_outputs(3502));
    outputs(11875) <= not(layer0_outputs(1200));
    outputs(11876) <= layer0_outputs(2916);
    outputs(11877) <= layer0_outputs(9647);
    outputs(11878) <= (layer0_outputs(8276)) xor (layer0_outputs(12325));
    outputs(11879) <= not((layer0_outputs(5058)) xor (layer0_outputs(3042)));
    outputs(11880) <= not((layer0_outputs(3045)) or (layer0_outputs(12170)));
    outputs(11881) <= layer0_outputs(993);
    outputs(11882) <= (layer0_outputs(12681)) or (layer0_outputs(6248));
    outputs(11883) <= not(layer0_outputs(12193));
    outputs(11884) <= (layer0_outputs(2617)) and not (layer0_outputs(6295));
    outputs(11885) <= not((layer0_outputs(592)) xor (layer0_outputs(10547)));
    outputs(11886) <= (layer0_outputs(7093)) xor (layer0_outputs(6233));
    outputs(11887) <= (layer0_outputs(12261)) xor (layer0_outputs(1218));
    outputs(11888) <= (layer0_outputs(10937)) and not (layer0_outputs(2376));
    outputs(11889) <= layer0_outputs(2501);
    outputs(11890) <= layer0_outputs(7888);
    outputs(11891) <= (layer0_outputs(591)) and not (layer0_outputs(2056));
    outputs(11892) <= (layer0_outputs(9214)) and (layer0_outputs(5594));
    outputs(11893) <= (layer0_outputs(4933)) and (layer0_outputs(11777));
    outputs(11894) <= not(layer0_outputs(9044));
    outputs(11895) <= not(layer0_outputs(11190));
    outputs(11896) <= not(layer0_outputs(8979));
    outputs(11897) <= (layer0_outputs(3892)) and not (layer0_outputs(10242));
    outputs(11898) <= not(layer0_outputs(10606)) or (layer0_outputs(10636));
    outputs(11899) <= (layer0_outputs(10722)) and not (layer0_outputs(9400));
    outputs(11900) <= layer0_outputs(8871);
    outputs(11901) <= layer0_outputs(6619);
    outputs(11902) <= not(layer0_outputs(6733));
    outputs(11903) <= not((layer0_outputs(4676)) or (layer0_outputs(10323)));
    outputs(11904) <= not(layer0_outputs(6427));
    outputs(11905) <= (layer0_outputs(5705)) and not (layer0_outputs(9226));
    outputs(11906) <= (layer0_outputs(10506)) and not (layer0_outputs(780));
    outputs(11907) <= not((layer0_outputs(2041)) and (layer0_outputs(4980)));
    outputs(11908) <= not(layer0_outputs(8269));
    outputs(11909) <= layer0_outputs(2157);
    outputs(11910) <= not(layer0_outputs(1010));
    outputs(11911) <= not((layer0_outputs(2982)) or (layer0_outputs(9742)));
    outputs(11912) <= layer0_outputs(4185);
    outputs(11913) <= layer0_outputs(11303);
    outputs(11914) <= layer0_outputs(6619);
    outputs(11915) <= (layer0_outputs(274)) and (layer0_outputs(2383));
    outputs(11916) <= (layer0_outputs(9951)) and (layer0_outputs(7924));
    outputs(11917) <= layer0_outputs(8872);
    outputs(11918) <= layer0_outputs(2970);
    outputs(11919) <= not(layer0_outputs(889));
    outputs(11920) <= not((layer0_outputs(3179)) or (layer0_outputs(10945)));
    outputs(11921) <= not(layer0_outputs(10259));
    outputs(11922) <= layer0_outputs(2448);
    outputs(11923) <= not((layer0_outputs(9710)) and (layer0_outputs(6205)));
    outputs(11924) <= (layer0_outputs(1210)) xor (layer0_outputs(4563));
    outputs(11925) <= not((layer0_outputs(4027)) xor (layer0_outputs(2163)));
    outputs(11926) <= layer0_outputs(4909);
    outputs(11927) <= not(layer0_outputs(11319));
    outputs(11928) <= layer0_outputs(6027);
    outputs(11929) <= layer0_outputs(7911);
    outputs(11930) <= (layer0_outputs(5174)) or (layer0_outputs(5715));
    outputs(11931) <= (layer0_outputs(5251)) and not (layer0_outputs(3887));
    outputs(11932) <= (layer0_outputs(4799)) and not (layer0_outputs(1501));
    outputs(11933) <= (layer0_outputs(10356)) and (layer0_outputs(3813));
    outputs(11934) <= (layer0_outputs(9659)) xor (layer0_outputs(7362));
    outputs(11935) <= not(layer0_outputs(5974));
    outputs(11936) <= layer0_outputs(9967);
    outputs(11937) <= not(layer0_outputs(31));
    outputs(11938) <= not((layer0_outputs(8726)) xor (layer0_outputs(12009)));
    outputs(11939) <= not(layer0_outputs(8649));
    outputs(11940) <= layer0_outputs(1185);
    outputs(11941) <= layer0_outputs(10386);
    outputs(11942) <= not((layer0_outputs(1007)) and (layer0_outputs(10174)));
    outputs(11943) <= (layer0_outputs(4284)) and (layer0_outputs(3625));
    outputs(11944) <= (layer0_outputs(3310)) and (layer0_outputs(12118));
    outputs(11945) <= (layer0_outputs(7544)) and (layer0_outputs(2700));
    outputs(11946) <= (layer0_outputs(9171)) and (layer0_outputs(5571));
    outputs(11947) <= layer0_outputs(9468);
    outputs(11948) <= not(layer0_outputs(12253));
    outputs(11949) <= layer0_outputs(7524);
    outputs(11950) <= not((layer0_outputs(1233)) xor (layer0_outputs(11431)));
    outputs(11951) <= layer0_outputs(1777);
    outputs(11952) <= (layer0_outputs(9240)) and (layer0_outputs(7916));
    outputs(11953) <= not((layer0_outputs(6035)) xor (layer0_outputs(10318)));
    outputs(11954) <= layer0_outputs(12224);
    outputs(11955) <= layer0_outputs(4893);
    outputs(11956) <= (layer0_outputs(9312)) xor (layer0_outputs(1676));
    outputs(11957) <= not(layer0_outputs(1727));
    outputs(11958) <= (layer0_outputs(3749)) xor (layer0_outputs(5664));
    outputs(11959) <= not((layer0_outputs(8026)) and (layer0_outputs(10217)));
    outputs(11960) <= not((layer0_outputs(2184)) or (layer0_outputs(10844)));
    outputs(11961) <= (layer0_outputs(845)) xor (layer0_outputs(191));
    outputs(11962) <= layer0_outputs(10006);
    outputs(11963) <= not(layer0_outputs(12201));
    outputs(11964) <= not(layer0_outputs(10904));
    outputs(11965) <= not(layer0_outputs(2377));
    outputs(11966) <= not((layer0_outputs(912)) xor (layer0_outputs(11422)));
    outputs(11967) <= not(layer0_outputs(199));
    outputs(11968) <= (layer0_outputs(11803)) and (layer0_outputs(7146));
    outputs(11969) <= (layer0_outputs(8448)) and not (layer0_outputs(12136));
    outputs(11970) <= (layer0_outputs(5628)) xor (layer0_outputs(2436));
    outputs(11971) <= not(layer0_outputs(1451));
    outputs(11972) <= not(layer0_outputs(5353));
    outputs(11973) <= (layer0_outputs(23)) or (layer0_outputs(12724));
    outputs(11974) <= layer0_outputs(12544);
    outputs(11975) <= layer0_outputs(822);
    outputs(11976) <= (layer0_outputs(6813)) xor (layer0_outputs(1662));
    outputs(11977) <= (layer0_outputs(1192)) xor (layer0_outputs(1481));
    outputs(11978) <= not((layer0_outputs(3730)) and (layer0_outputs(12394)));
    outputs(11979) <= (layer0_outputs(575)) and (layer0_outputs(7383));
    outputs(11980) <= layer0_outputs(11666);
    outputs(11981) <= layer0_outputs(2607);
    outputs(11982) <= (layer0_outputs(7711)) xor (layer0_outputs(1516));
    outputs(11983) <= (layer0_outputs(3763)) xor (layer0_outputs(8926));
    outputs(11984) <= (layer0_outputs(3585)) and not (layer0_outputs(5256));
    outputs(11985) <= layer0_outputs(7439);
    outputs(11986) <= not((layer0_outputs(2093)) xor (layer0_outputs(8475)));
    outputs(11987) <= (layer0_outputs(4347)) xor (layer0_outputs(1562));
    outputs(11988) <= not(layer0_outputs(3012));
    outputs(11989) <= not((layer0_outputs(7178)) xor (layer0_outputs(5183)));
    outputs(11990) <= layer0_outputs(149);
    outputs(11991) <= not(layer0_outputs(2755));
    outputs(11992) <= (layer0_outputs(8334)) xor (layer0_outputs(7448));
    outputs(11993) <= (layer0_outputs(8572)) xor (layer0_outputs(12172));
    outputs(11994) <= not(layer0_outputs(6478));
    outputs(11995) <= (layer0_outputs(12506)) xor (layer0_outputs(1776));
    outputs(11996) <= not((layer0_outputs(1780)) or (layer0_outputs(4883)));
    outputs(11997) <= layer0_outputs(1358);
    outputs(11998) <= not(layer0_outputs(7903));
    outputs(11999) <= not((layer0_outputs(9953)) xor (layer0_outputs(12173)));
    outputs(12000) <= not((layer0_outputs(11450)) xor (layer0_outputs(12275)));
    outputs(12001) <= layer0_outputs(7847);
    outputs(12002) <= (layer0_outputs(9963)) and not (layer0_outputs(11438));
    outputs(12003) <= not(layer0_outputs(9467));
    outputs(12004) <= layer0_outputs(5262);
    outputs(12005) <= not(layer0_outputs(393));
    outputs(12006) <= layer0_outputs(9871);
    outputs(12007) <= not((layer0_outputs(10734)) xor (layer0_outputs(6197)));
    outputs(12008) <= (layer0_outputs(7465)) or (layer0_outputs(1499));
    outputs(12009) <= not(layer0_outputs(1415));
    outputs(12010) <= not(layer0_outputs(4063)) or (layer0_outputs(4790));
    outputs(12011) <= (layer0_outputs(2977)) xor (layer0_outputs(11071));
    outputs(12012) <= not((layer0_outputs(7192)) xor (layer0_outputs(9035)));
    outputs(12013) <= (layer0_outputs(5887)) xor (layer0_outputs(1587));
    outputs(12014) <= not((layer0_outputs(322)) xor (layer0_outputs(1957)));
    outputs(12015) <= not(layer0_outputs(1316));
    outputs(12016) <= (layer0_outputs(887)) xor (layer0_outputs(9885));
    outputs(12017) <= layer0_outputs(11928);
    outputs(12018) <= (layer0_outputs(9550)) and (layer0_outputs(7482));
    outputs(12019) <= not(layer0_outputs(8185));
    outputs(12020) <= not((layer0_outputs(10716)) xor (layer0_outputs(12529)));
    outputs(12021) <= not((layer0_outputs(5329)) xor (layer0_outputs(7657)));
    outputs(12022) <= (layer0_outputs(2492)) xor (layer0_outputs(7498));
    outputs(12023) <= (layer0_outputs(8306)) and not (layer0_outputs(2031));
    outputs(12024) <= not(layer0_outputs(12691));
    outputs(12025) <= not(layer0_outputs(9940));
    outputs(12026) <= not(layer0_outputs(7122));
    outputs(12027) <= layer0_outputs(8909);
    outputs(12028) <= layer0_outputs(11587);
    outputs(12029) <= not((layer0_outputs(11123)) xor (layer0_outputs(8533)));
    outputs(12030) <= (layer0_outputs(10056)) xor (layer0_outputs(6118));
    outputs(12031) <= not((layer0_outputs(7561)) or (layer0_outputs(8768)));
    outputs(12032) <= layer0_outputs(402);
    outputs(12033) <= not(layer0_outputs(6625));
    outputs(12034) <= not(layer0_outputs(1045)) or (layer0_outputs(7713));
    outputs(12035) <= not((layer0_outputs(1814)) xor (layer0_outputs(2286)));
    outputs(12036) <= (layer0_outputs(6444)) xor (layer0_outputs(10315));
    outputs(12037) <= layer0_outputs(11461);
    outputs(12038) <= not(layer0_outputs(7742));
    outputs(12039) <= layer0_outputs(8320);
    outputs(12040) <= not((layer0_outputs(4712)) xor (layer0_outputs(12397)));
    outputs(12041) <= layer0_outputs(9572);
    outputs(12042) <= not(layer0_outputs(5504)) or (layer0_outputs(5123));
    outputs(12043) <= not((layer0_outputs(9494)) xor (layer0_outputs(3920)));
    outputs(12044) <= layer0_outputs(1833);
    outputs(12045) <= not((layer0_outputs(11413)) xor (layer0_outputs(1026)));
    outputs(12046) <= not((layer0_outputs(2627)) xor (layer0_outputs(1681)));
    outputs(12047) <= not(layer0_outputs(4177));
    outputs(12048) <= not((layer0_outputs(8889)) xor (layer0_outputs(6722)));
    outputs(12049) <= not(layer0_outputs(12530));
    outputs(12050) <= layer0_outputs(1105);
    outputs(12051) <= (layer0_outputs(8060)) xor (layer0_outputs(566));
    outputs(12052) <= layer0_outputs(6377);
    outputs(12053) <= not((layer0_outputs(8487)) xor (layer0_outputs(6706)));
    outputs(12054) <= not(layer0_outputs(11286));
    outputs(12055) <= (layer0_outputs(9725)) xor (layer0_outputs(10691));
    outputs(12056) <= not(layer0_outputs(5352)) or (layer0_outputs(1772));
    outputs(12057) <= not(layer0_outputs(12792));
    outputs(12058) <= not(layer0_outputs(683)) or (layer0_outputs(9900));
    outputs(12059) <= (layer0_outputs(4673)) xor (layer0_outputs(9264));
    outputs(12060) <= not((layer0_outputs(8104)) or (layer0_outputs(2692)));
    outputs(12061) <= not(layer0_outputs(4750));
    outputs(12062) <= layer0_outputs(6850);
    outputs(12063) <= layer0_outputs(1897);
    outputs(12064) <= layer0_outputs(9333);
    outputs(12065) <= not(layer0_outputs(7431)) or (layer0_outputs(3625));
    outputs(12066) <= not(layer0_outputs(11158));
    outputs(12067) <= not((layer0_outputs(10412)) or (layer0_outputs(9374)));
    outputs(12068) <= not((layer0_outputs(6192)) or (layer0_outputs(11257)));
    outputs(12069) <= not((layer0_outputs(1092)) or (layer0_outputs(4073)));
    outputs(12070) <= layer0_outputs(5286);
    outputs(12071) <= (layer0_outputs(874)) and not (layer0_outputs(290));
    outputs(12072) <= layer0_outputs(12659);
    outputs(12073) <= layer0_outputs(9587);
    outputs(12074) <= layer0_outputs(10300);
    outputs(12075) <= (layer0_outputs(11796)) and not (layer0_outputs(4178));
    outputs(12076) <= not(layer0_outputs(3893));
    outputs(12077) <= not(layer0_outputs(10573));
    outputs(12078) <= not((layer0_outputs(7495)) or (layer0_outputs(8991)));
    outputs(12079) <= not(layer0_outputs(10412));
    outputs(12080) <= not((layer0_outputs(1138)) or (layer0_outputs(11829)));
    outputs(12081) <= not(layer0_outputs(6681));
    outputs(12082) <= not((layer0_outputs(11550)) xor (layer0_outputs(1691)));
    outputs(12083) <= not(layer0_outputs(4735));
    outputs(12084) <= not((layer0_outputs(7137)) or (layer0_outputs(3027)));
    outputs(12085) <= (layer0_outputs(11927)) and not (layer0_outputs(12454));
    outputs(12086) <= (layer0_outputs(940)) and not (layer0_outputs(4003));
    outputs(12087) <= not(layer0_outputs(9825));
    outputs(12088) <= (layer0_outputs(6907)) xor (layer0_outputs(9453));
    outputs(12089) <= layer0_outputs(5701);
    outputs(12090) <= not(layer0_outputs(4402));
    outputs(12091) <= not((layer0_outputs(371)) xor (layer0_outputs(10888)));
    outputs(12092) <= layer0_outputs(11576);
    outputs(12093) <= not((layer0_outputs(1644)) xor (layer0_outputs(4064)));
    outputs(12094) <= (layer0_outputs(3032)) xor (layer0_outputs(11275));
    outputs(12095) <= not((layer0_outputs(7693)) xor (layer0_outputs(11911)));
    outputs(12096) <= not((layer0_outputs(1469)) xor (layer0_outputs(2531)));
    outputs(12097) <= not(layer0_outputs(10793));
    outputs(12098) <= not((layer0_outputs(1775)) xor (layer0_outputs(11785)));
    outputs(12099) <= (layer0_outputs(8661)) xor (layer0_outputs(5256));
    outputs(12100) <= not(layer0_outputs(1349)) or (layer0_outputs(4772));
    outputs(12101) <= layer0_outputs(7383);
    outputs(12102) <= not(layer0_outputs(10997));
    outputs(12103) <= not(layer0_outputs(12340));
    outputs(12104) <= (layer0_outputs(6123)) xor (layer0_outputs(12699));
    outputs(12105) <= not(layer0_outputs(10725));
    outputs(12106) <= layer0_outputs(11163);
    outputs(12107) <= layer0_outputs(4114);
    outputs(12108) <= (layer0_outputs(5408)) xor (layer0_outputs(6093));
    outputs(12109) <= (layer0_outputs(4476)) and not (layer0_outputs(1600));
    outputs(12110) <= not((layer0_outputs(5829)) xor (layer0_outputs(9167)));
    outputs(12111) <= layer0_outputs(9117);
    outputs(12112) <= (layer0_outputs(7056)) xor (layer0_outputs(6764));
    outputs(12113) <= not(layer0_outputs(5751));
    outputs(12114) <= (layer0_outputs(3762)) and (layer0_outputs(534));
    outputs(12115) <= not((layer0_outputs(7826)) xor (layer0_outputs(3139)));
    outputs(12116) <= (layer0_outputs(11029)) or (layer0_outputs(5625));
    outputs(12117) <= not(layer0_outputs(6244));
    outputs(12118) <= (layer0_outputs(8597)) xor (layer0_outputs(9724));
    outputs(12119) <= layer0_outputs(2034);
    outputs(12120) <= layer0_outputs(2299);
    outputs(12121) <= not(layer0_outputs(5542));
    outputs(12122) <= not((layer0_outputs(7033)) xor (layer0_outputs(10878)));
    outputs(12123) <= not(layer0_outputs(6004));
    outputs(12124) <= not((layer0_outputs(5842)) xor (layer0_outputs(7931)));
    outputs(12125) <= layer0_outputs(6893);
    outputs(12126) <= not(layer0_outputs(3469));
    outputs(12127) <= (layer0_outputs(2162)) and not (layer0_outputs(11234));
    outputs(12128) <= not((layer0_outputs(1702)) xor (layer0_outputs(10450)));
    outputs(12129) <= layer0_outputs(4065);
    outputs(12130) <= layer0_outputs(840);
    outputs(12131) <= (layer0_outputs(2848)) and not (layer0_outputs(9737));
    outputs(12132) <= not(layer0_outputs(11324)) or (layer0_outputs(12668));
    outputs(12133) <= not((layer0_outputs(4281)) xor (layer0_outputs(2919)));
    outputs(12134) <= (layer0_outputs(744)) and not (layer0_outputs(1503));
    outputs(12135) <= not(layer0_outputs(3665)) or (layer0_outputs(2032));
    outputs(12136) <= (layer0_outputs(10684)) and not (layer0_outputs(2601));
    outputs(12137) <= not((layer0_outputs(11995)) xor (layer0_outputs(8065)));
    outputs(12138) <= not((layer0_outputs(8758)) xor (layer0_outputs(12508)));
    outputs(12139) <= (layer0_outputs(2680)) and not (layer0_outputs(2631));
    outputs(12140) <= not((layer0_outputs(3450)) or (layer0_outputs(9981)));
    outputs(12141) <= layer0_outputs(9769);
    outputs(12142) <= not((layer0_outputs(5169)) or (layer0_outputs(11125)));
    outputs(12143) <= not(layer0_outputs(197));
    outputs(12144) <= (layer0_outputs(6914)) and (layer0_outputs(10163));
    outputs(12145) <= (layer0_outputs(4464)) xor (layer0_outputs(2652));
    outputs(12146) <= (layer0_outputs(10108)) and not (layer0_outputs(11155));
    outputs(12147) <= (layer0_outputs(1597)) xor (layer0_outputs(3879));
    outputs(12148) <= layer0_outputs(9451);
    outputs(12149) <= (layer0_outputs(11672)) and not (layer0_outputs(6435));
    outputs(12150) <= not(layer0_outputs(12259));
    outputs(12151) <= (layer0_outputs(12684)) xor (layer0_outputs(11798));
    outputs(12152) <= not((layer0_outputs(5725)) xor (layer0_outputs(1582)));
    outputs(12153) <= (layer0_outputs(6513)) xor (layer0_outputs(8356));
    outputs(12154) <= not((layer0_outputs(9881)) and (layer0_outputs(2459)));
    outputs(12155) <= not(layer0_outputs(9030));
    outputs(12156) <= not(layer0_outputs(5272)) or (layer0_outputs(4713));
    outputs(12157) <= (layer0_outputs(4202)) xor (layer0_outputs(494));
    outputs(12158) <= not((layer0_outputs(9619)) xor (layer0_outputs(4595)));
    outputs(12159) <= not(layer0_outputs(10015));
    outputs(12160) <= not((layer0_outputs(10650)) xor (layer0_outputs(4224)));
    outputs(12161) <= not(layer0_outputs(5110));
    outputs(12162) <= not(layer0_outputs(6411));
    outputs(12163) <= layer0_outputs(12212);
    outputs(12164) <= (layer0_outputs(4751)) or (layer0_outputs(2965));
    outputs(12165) <= (layer0_outputs(9425)) or (layer0_outputs(3935));
    outputs(12166) <= (layer0_outputs(4695)) and (layer0_outputs(11970));
    outputs(12167) <= not(layer0_outputs(9111));
    outputs(12168) <= not(layer0_outputs(12061));
    outputs(12169) <= layer0_outputs(1111);
    outputs(12170) <= layer0_outputs(10556);
    outputs(12171) <= not((layer0_outputs(11247)) or (layer0_outputs(3776)));
    outputs(12172) <= not(layer0_outputs(8820));
    outputs(12173) <= not(layer0_outputs(10210));
    outputs(12174) <= not((layer0_outputs(8646)) xor (layer0_outputs(4992)));
    outputs(12175) <= not(layer0_outputs(1118));
    outputs(12176) <= (layer0_outputs(8977)) xor (layer0_outputs(7502));
    outputs(12177) <= not((layer0_outputs(9589)) xor (layer0_outputs(7565)));
    outputs(12178) <= not(layer0_outputs(4179));
    outputs(12179) <= not((layer0_outputs(4260)) xor (layer0_outputs(6017)));
    outputs(12180) <= not(layer0_outputs(10698));
    outputs(12181) <= not(layer0_outputs(1570));
    outputs(12182) <= layer0_outputs(557);
    outputs(12183) <= layer0_outputs(2283);
    outputs(12184) <= (layer0_outputs(3118)) xor (layer0_outputs(9337));
    outputs(12185) <= (layer0_outputs(11543)) and not (layer0_outputs(3333));
    outputs(12186) <= not(layer0_outputs(2784));
    outputs(12187) <= not((layer0_outputs(9336)) xor (layer0_outputs(5819)));
    outputs(12188) <= not(layer0_outputs(8322));
    outputs(12189) <= layer0_outputs(10551);
    outputs(12190) <= not((layer0_outputs(1908)) or (layer0_outputs(2427)));
    outputs(12191) <= not(layer0_outputs(8993)) or (layer0_outputs(674));
    outputs(12192) <= not((layer0_outputs(11996)) xor (layer0_outputs(11166)));
    outputs(12193) <= layer0_outputs(12123);
    outputs(12194) <= layer0_outputs(2365);
    outputs(12195) <= not((layer0_outputs(737)) xor (layer0_outputs(5503)));
    outputs(12196) <= not((layer0_outputs(12606)) and (layer0_outputs(9488)));
    outputs(12197) <= (layer0_outputs(4835)) xor (layer0_outputs(4880));
    outputs(12198) <= layer0_outputs(10336);
    outputs(12199) <= not(layer0_outputs(4387));
    outputs(12200) <= not(layer0_outputs(11513));
    outputs(12201) <= (layer0_outputs(9399)) xor (layer0_outputs(8201));
    outputs(12202) <= not((layer0_outputs(9521)) xor (layer0_outputs(2939)));
    outputs(12203) <= (layer0_outputs(4798)) and not (layer0_outputs(473));
    outputs(12204) <= not((layer0_outputs(3102)) xor (layer0_outputs(6604)));
    outputs(12205) <= (layer0_outputs(174)) xor (layer0_outputs(3611));
    outputs(12206) <= layer0_outputs(1291);
    outputs(12207) <= (layer0_outputs(5279)) xor (layer0_outputs(6996));
    outputs(12208) <= not(layer0_outputs(7123)) or (layer0_outputs(10620));
    outputs(12209) <= not((layer0_outputs(11432)) xor (layer0_outputs(12643)));
    outputs(12210) <= layer0_outputs(5640);
    outputs(12211) <= not(layer0_outputs(12423));
    outputs(12212) <= not((layer0_outputs(10635)) or (layer0_outputs(457)));
    outputs(12213) <= not(layer0_outputs(5685));
    outputs(12214) <= (layer0_outputs(335)) xor (layer0_outputs(875));
    outputs(12215) <= not((layer0_outputs(2517)) or (layer0_outputs(8114)));
    outputs(12216) <= (layer0_outputs(7754)) xor (layer0_outputs(9865));
    outputs(12217) <= (layer0_outputs(11321)) xor (layer0_outputs(10334));
    outputs(12218) <= not(layer0_outputs(2290));
    outputs(12219) <= (layer0_outputs(7200)) and (layer0_outputs(5170));
    outputs(12220) <= not((layer0_outputs(10305)) or (layer0_outputs(6418)));
    outputs(12221) <= not(layer0_outputs(7884));
    outputs(12222) <= not((layer0_outputs(8884)) and (layer0_outputs(8200)));
    outputs(12223) <= not((layer0_outputs(9974)) xor (layer0_outputs(6477)));
    outputs(12224) <= (layer0_outputs(1250)) xor (layer0_outputs(8403));
    outputs(12225) <= not(layer0_outputs(11866));
    outputs(12226) <= (layer0_outputs(10810)) xor (layer0_outputs(4974));
    outputs(12227) <= (layer0_outputs(8321)) xor (layer0_outputs(2710));
    outputs(12228) <= (layer0_outputs(10915)) and not (layer0_outputs(2506));
    outputs(12229) <= (layer0_outputs(1854)) xor (layer0_outputs(221));
    outputs(12230) <= not((layer0_outputs(6448)) xor (layer0_outputs(10593)));
    outputs(12231) <= not((layer0_outputs(3429)) or (layer0_outputs(9639)));
    outputs(12232) <= layer0_outputs(4070);
    outputs(12233) <= not((layer0_outputs(3375)) xor (layer0_outputs(12793)));
    outputs(12234) <= not((layer0_outputs(6555)) and (layer0_outputs(9557)));
    outputs(12235) <= layer0_outputs(1163);
    outputs(12236) <= layer0_outputs(4550);
    outputs(12237) <= not(layer0_outputs(3557)) or (layer0_outputs(1829));
    outputs(12238) <= layer0_outputs(7666);
    outputs(12239) <= not(layer0_outputs(3904));
    outputs(12240) <= not((layer0_outputs(6713)) and (layer0_outputs(6149)));
    outputs(12241) <= layer0_outputs(2775);
    outputs(12242) <= not((layer0_outputs(10752)) xor (layer0_outputs(7339)));
    outputs(12243) <= not(layer0_outputs(3770));
    outputs(12244) <= not((layer0_outputs(10756)) xor (layer0_outputs(12071)));
    outputs(12245) <= (layer0_outputs(9023)) xor (layer0_outputs(3809));
    outputs(12246) <= not((layer0_outputs(10779)) xor (layer0_outputs(10211)));
    outputs(12247) <= (layer0_outputs(7965)) and (layer0_outputs(12384));
    outputs(12248) <= (layer0_outputs(6979)) and (layer0_outputs(4787));
    outputs(12249) <= (layer0_outputs(2550)) xor (layer0_outputs(7551));
    outputs(12250) <= (layer0_outputs(8880)) and not (layer0_outputs(7226));
    outputs(12251) <= (layer0_outputs(5955)) and not (layer0_outputs(2865));
    outputs(12252) <= not(layer0_outputs(8343));
    outputs(12253) <= not((layer0_outputs(3793)) xor (layer0_outputs(9886)));
    outputs(12254) <= not((layer0_outputs(9818)) xor (layer0_outputs(4906)));
    outputs(12255) <= not(layer0_outputs(8179));
    outputs(12256) <= not(layer0_outputs(10934));
    outputs(12257) <= (layer0_outputs(2442)) and (layer0_outputs(1718));
    outputs(12258) <= not(layer0_outputs(565));
    outputs(12259) <= not((layer0_outputs(7403)) xor (layer0_outputs(3481)));
    outputs(12260) <= (layer0_outputs(1574)) xor (layer0_outputs(12765));
    outputs(12261) <= (layer0_outputs(6033)) and not (layer0_outputs(1981));
    outputs(12262) <= not((layer0_outputs(6702)) xor (layer0_outputs(11246)));
    outputs(12263) <= (layer0_outputs(5191)) xor (layer0_outputs(9694));
    outputs(12264) <= not((layer0_outputs(10654)) xor (layer0_outputs(10358)));
    outputs(12265) <= not(layer0_outputs(12617));
    outputs(12266) <= (layer0_outputs(851)) and (layer0_outputs(8112));
    outputs(12267) <= layer0_outputs(6442);
    outputs(12268) <= (layer0_outputs(9490)) and not (layer0_outputs(2921));
    outputs(12269) <= layer0_outputs(6668);
    outputs(12270) <= (layer0_outputs(3244)) xor (layer0_outputs(10155));
    outputs(12271) <= (layer0_outputs(6856)) and not (layer0_outputs(8488));
    outputs(12272) <= not(layer0_outputs(2703));
    outputs(12273) <= layer0_outputs(1571);
    outputs(12274) <= (layer0_outputs(9489)) and not (layer0_outputs(10038));
    outputs(12275) <= not((layer0_outputs(6537)) xor (layer0_outputs(9233)));
    outputs(12276) <= layer0_outputs(11517);
    outputs(12277) <= not((layer0_outputs(3720)) xor (layer0_outputs(2506)));
    outputs(12278) <= not((layer0_outputs(8875)) xor (layer0_outputs(11956)));
    outputs(12279) <= (layer0_outputs(11556)) and not (layer0_outputs(5528));
    outputs(12280) <= (layer0_outputs(5929)) xor (layer0_outputs(12242));
    outputs(12281) <= layer0_outputs(11562);
    outputs(12282) <= (layer0_outputs(9473)) and (layer0_outputs(1749));
    outputs(12283) <= not((layer0_outputs(3928)) xor (layer0_outputs(3932)));
    outputs(12284) <= (layer0_outputs(11934)) xor (layer0_outputs(12213));
    outputs(12285) <= (layer0_outputs(8903)) xor (layer0_outputs(6225));
    outputs(12286) <= layer0_outputs(1927);
    outputs(12287) <= (layer0_outputs(7958)) xor (layer0_outputs(5752));
    outputs(12288) <= not((layer0_outputs(3251)) xor (layer0_outputs(12321)));
    outputs(12289) <= not(layer0_outputs(10166)) or (layer0_outputs(9874));
    outputs(12290) <= (layer0_outputs(4184)) xor (layer0_outputs(7020));
    outputs(12291) <= not((layer0_outputs(4250)) xor (layer0_outputs(12673)));
    outputs(12292) <= (layer0_outputs(2693)) and not (layer0_outputs(2246));
    outputs(12293) <= not(layer0_outputs(1342));
    outputs(12294) <= not(layer0_outputs(6845));
    outputs(12295) <= not((layer0_outputs(4935)) and (layer0_outputs(7891)));
    outputs(12296) <= layer0_outputs(4205);
    outputs(12297) <= not(layer0_outputs(10041));
    outputs(12298) <= layer0_outputs(11262);
    outputs(12299) <= not(layer0_outputs(3082));
    outputs(12300) <= (layer0_outputs(12365)) xor (layer0_outputs(1685));
    outputs(12301) <= layer0_outputs(9298);
    outputs(12302) <= (layer0_outputs(3114)) xor (layer0_outputs(10298));
    outputs(12303) <= (layer0_outputs(7590)) xor (layer0_outputs(409));
    outputs(12304) <= not(layer0_outputs(4371));
    outputs(12305) <= (layer0_outputs(7852)) and not (layer0_outputs(2851));
    outputs(12306) <= not(layer0_outputs(2041));
    outputs(12307) <= not(layer0_outputs(10872));
    outputs(12308) <= layer0_outputs(3542);
    outputs(12309) <= layer0_outputs(11109);
    outputs(12310) <= layer0_outputs(5211);
    outputs(12311) <= not(layer0_outputs(4690));
    outputs(12312) <= layer0_outputs(11561);
    outputs(12313) <= (layer0_outputs(2911)) and not (layer0_outputs(8622));
    outputs(12314) <= (layer0_outputs(12195)) and (layer0_outputs(5043));
    outputs(12315) <= not((layer0_outputs(253)) xor (layer0_outputs(5782)));
    outputs(12316) <= layer0_outputs(7560);
    outputs(12317) <= not(layer0_outputs(10180));
    outputs(12318) <= not(layer0_outputs(4129));
    outputs(12319) <= not((layer0_outputs(4693)) xor (layer0_outputs(3730)));
    outputs(12320) <= (layer0_outputs(4013)) and not (layer0_outputs(6236));
    outputs(12321) <= not((layer0_outputs(7469)) xor (layer0_outputs(2642)));
    outputs(12322) <= not((layer0_outputs(6603)) xor (layer0_outputs(6754)));
    outputs(12323) <= not((layer0_outputs(2582)) xor (layer0_outputs(1745)));
    outputs(12324) <= not((layer0_outputs(9649)) xor (layer0_outputs(10670)));
    outputs(12325) <= (layer0_outputs(12588)) and not (layer0_outputs(3199));
    outputs(12326) <= not(layer0_outputs(9343)) or (layer0_outputs(10617));
    outputs(12327) <= (layer0_outputs(6050)) xor (layer0_outputs(2523));
    outputs(12328) <= (layer0_outputs(12330)) xor (layer0_outputs(9457));
    outputs(12329) <= not(layer0_outputs(7914));
    outputs(12330) <= not((layer0_outputs(8499)) xor (layer0_outputs(11347)));
    outputs(12331) <= layer0_outputs(1078);
    outputs(12332) <= not(layer0_outputs(11376));
    outputs(12333) <= layer0_outputs(6848);
    outputs(12334) <= not(layer0_outputs(10418));
    outputs(12335) <= not((layer0_outputs(6449)) xor (layer0_outputs(4134)));
    outputs(12336) <= (layer0_outputs(12083)) xor (layer0_outputs(12427));
    outputs(12337) <= (layer0_outputs(10339)) and not (layer0_outputs(1616));
    outputs(12338) <= layer0_outputs(9247);
    outputs(12339) <= not(layer0_outputs(10297));
    outputs(12340) <= not(layer0_outputs(5146));
    outputs(12341) <= (layer0_outputs(1367)) xor (layer0_outputs(1997));
    outputs(12342) <= not((layer0_outputs(5467)) or (layer0_outputs(8953)));
    outputs(12343) <= not((layer0_outputs(6974)) and (layer0_outputs(4248)));
    outputs(12344) <= not((layer0_outputs(5393)) xor (layer0_outputs(7440)));
    outputs(12345) <= (layer0_outputs(6003)) xor (layer0_outputs(5362));
    outputs(12346) <= not((layer0_outputs(7270)) or (layer0_outputs(6353)));
    outputs(12347) <= not(layer0_outputs(12221)) or (layer0_outputs(5778));
    outputs(12348) <= not(layer0_outputs(3263));
    outputs(12349) <= layer0_outputs(10267);
    outputs(12350) <= (layer0_outputs(838)) xor (layer0_outputs(10840));
    outputs(12351) <= (layer0_outputs(12148)) and not (layer0_outputs(1040));
    outputs(12352) <= not(layer0_outputs(7649)) or (layer0_outputs(5001));
    outputs(12353) <= not(layer0_outputs(11964));
    outputs(12354) <= (layer0_outputs(10626)) xor (layer0_outputs(7115));
    outputs(12355) <= not((layer0_outputs(6699)) xor (layer0_outputs(2700)));
    outputs(12356) <= not((layer0_outputs(583)) or (layer0_outputs(2675)));
    outputs(12357) <= not((layer0_outputs(4814)) xor (layer0_outputs(2359)));
    outputs(12358) <= (layer0_outputs(8674)) xor (layer0_outputs(4533));
    outputs(12359) <= not(layer0_outputs(11600));
    outputs(12360) <= layer0_outputs(6278);
    outputs(12361) <= (layer0_outputs(288)) xor (layer0_outputs(8599));
    outputs(12362) <= layer0_outputs(605);
    outputs(12363) <= (layer0_outputs(8425)) and (layer0_outputs(3780));
    outputs(12364) <= not((layer0_outputs(3699)) xor (layer0_outputs(2871)));
    outputs(12365) <= (layer0_outputs(8238)) and not (layer0_outputs(3227));
    outputs(12366) <= not((layer0_outputs(7646)) xor (layer0_outputs(3517)));
    outputs(12367) <= not(layer0_outputs(2884)) or (layer0_outputs(3531));
    outputs(12368) <= (layer0_outputs(2528)) and not (layer0_outputs(9281));
    outputs(12369) <= (layer0_outputs(1361)) xor (layer0_outputs(1231));
    outputs(12370) <= layer0_outputs(4421);
    outputs(12371) <= not(layer0_outputs(8001));
    outputs(12372) <= (layer0_outputs(12769)) xor (layer0_outputs(329));
    outputs(12373) <= (layer0_outputs(11921)) xor (layer0_outputs(12222));
    outputs(12374) <= not(layer0_outputs(3669));
    outputs(12375) <= layer0_outputs(10964);
    outputs(12376) <= (layer0_outputs(8553)) xor (layer0_outputs(3922));
    outputs(12377) <= layer0_outputs(2276);
    outputs(12378) <= (layer0_outputs(11039)) or (layer0_outputs(7986));
    outputs(12379) <= not((layer0_outputs(9613)) or (layer0_outputs(11584)));
    outputs(12380) <= not(layer0_outputs(12722));
    outputs(12381) <= (layer0_outputs(11325)) and (layer0_outputs(1305));
    outputs(12382) <= not((layer0_outputs(5537)) or (layer0_outputs(7625)));
    outputs(12383) <= not((layer0_outputs(2100)) and (layer0_outputs(6411)));
    outputs(12384) <= (layer0_outputs(879)) xor (layer0_outputs(9123));
    outputs(12385) <= not(layer0_outputs(1845)) or (layer0_outputs(11049));
    outputs(12386) <= not((layer0_outputs(2941)) or (layer0_outputs(2367)));
    outputs(12387) <= (layer0_outputs(4204)) or (layer0_outputs(8848));
    outputs(12388) <= layer0_outputs(4238);
    outputs(12389) <= (layer0_outputs(10351)) xor (layer0_outputs(9758));
    outputs(12390) <= layer0_outputs(8007);
    outputs(12391) <= (layer0_outputs(10073)) xor (layer0_outputs(273));
    outputs(12392) <= layer0_outputs(9165);
    outputs(12393) <= not((layer0_outputs(12700)) or (layer0_outputs(12084)));
    outputs(12394) <= layer0_outputs(11230);
    outputs(12395) <= (layer0_outputs(8912)) xor (layer0_outputs(10359));
    outputs(12396) <= not((layer0_outputs(278)) xor (layer0_outputs(861)));
    outputs(12397) <= not(layer0_outputs(5307));
    outputs(12398) <= not(layer0_outputs(3757)) or (layer0_outputs(12452));
    outputs(12399) <= layer0_outputs(6617);
    outputs(12400) <= not(layer0_outputs(5078));
    outputs(12401) <= not(layer0_outputs(6142)) or (layer0_outputs(691));
    outputs(12402) <= not((layer0_outputs(772)) and (layer0_outputs(7094)));
    outputs(12403) <= layer0_outputs(7295);
    outputs(12404) <= (layer0_outputs(4954)) or (layer0_outputs(11616));
    outputs(12405) <= not(layer0_outputs(145));
    outputs(12406) <= not((layer0_outputs(6646)) xor (layer0_outputs(1865)));
    outputs(12407) <= layer0_outputs(4289);
    outputs(12408) <= (layer0_outputs(8461)) and not (layer0_outputs(10470));
    outputs(12409) <= not((layer0_outputs(6219)) xor (layer0_outputs(1466)));
    outputs(12410) <= not(layer0_outputs(3649));
    outputs(12411) <= layer0_outputs(5721);
    outputs(12412) <= (layer0_outputs(730)) and not (layer0_outputs(8114));
    outputs(12413) <= not((layer0_outputs(12104)) xor (layer0_outputs(12423)));
    outputs(12414) <= (layer0_outputs(8244)) and (layer0_outputs(11754));
    outputs(12415) <= (layer0_outputs(6380)) xor (layer0_outputs(8459));
    outputs(12416) <= not((layer0_outputs(8807)) xor (layer0_outputs(795)));
    outputs(12417) <= not(layer0_outputs(2310));
    outputs(12418) <= not((layer0_outputs(786)) and (layer0_outputs(1944)));
    outputs(12419) <= not((layer0_outputs(4663)) xor (layer0_outputs(6189)));
    outputs(12420) <= layer0_outputs(156);
    outputs(12421) <= layer0_outputs(7555);
    outputs(12422) <= layer0_outputs(10788);
    outputs(12423) <= (layer0_outputs(2862)) and not (layer0_outputs(2631));
    outputs(12424) <= not((layer0_outputs(12547)) xor (layer0_outputs(994)));
    outputs(12425) <= (layer0_outputs(3334)) and not (layer0_outputs(10212));
    outputs(12426) <= layer0_outputs(11769);
    outputs(12427) <= not(layer0_outputs(152));
    outputs(12428) <= layer0_outputs(7984);
    outputs(12429) <= (layer0_outputs(4426)) or (layer0_outputs(2076));
    outputs(12430) <= (layer0_outputs(1480)) xor (layer0_outputs(1679));
    outputs(12431) <= not(layer0_outputs(5652)) or (layer0_outputs(2016));
    outputs(12432) <= not((layer0_outputs(326)) or (layer0_outputs(6923)));
    outputs(12433) <= layer0_outputs(10790);
    outputs(12434) <= (layer0_outputs(3169)) or (layer0_outputs(2107));
    outputs(12435) <= (layer0_outputs(3066)) xor (layer0_outputs(1135));
    outputs(12436) <= not(layer0_outputs(5741)) or (layer0_outputs(11281));
    outputs(12437) <= layer0_outputs(5245);
    outputs(12438) <= not(layer0_outputs(776));
    outputs(12439) <= not(layer0_outputs(12109));
    outputs(12440) <= (layer0_outputs(5157)) and not (layer0_outputs(7710));
    outputs(12441) <= (layer0_outputs(6986)) and not (layer0_outputs(8885));
    outputs(12442) <= (layer0_outputs(146)) xor (layer0_outputs(5088));
    outputs(12443) <= not(layer0_outputs(12261));
    outputs(12444) <= layer0_outputs(3477);
    outputs(12445) <= (layer0_outputs(5511)) and (layer0_outputs(11898));
    outputs(12446) <= (layer0_outputs(12287)) xor (layer0_outputs(9342));
    outputs(12447) <= not((layer0_outputs(9026)) or (layer0_outputs(9780)));
    outputs(12448) <= (layer0_outputs(9107)) or (layer0_outputs(6014));
    outputs(12449) <= (layer0_outputs(8314)) xor (layer0_outputs(4783));
    outputs(12450) <= not(layer0_outputs(9325));
    outputs(12451) <= (layer0_outputs(12681)) and not (layer0_outputs(8277));
    outputs(12452) <= not(layer0_outputs(7878));
    outputs(12453) <= (layer0_outputs(6095)) or (layer0_outputs(3434));
    outputs(12454) <= (layer0_outputs(10651)) or (layer0_outputs(6382));
    outputs(12455) <= layer0_outputs(7484);
    outputs(12456) <= layer0_outputs(10285);
    outputs(12457) <= layer0_outputs(9530);
    outputs(12458) <= not((layer0_outputs(2653)) xor (layer0_outputs(8437)));
    outputs(12459) <= not((layer0_outputs(6434)) xor (layer0_outputs(1576)));
    outputs(12460) <= not((layer0_outputs(238)) xor (layer0_outputs(4585)));
    outputs(12461) <= layer0_outputs(9455);
    outputs(12462) <= not((layer0_outputs(7047)) xor (layer0_outputs(5653)));
    outputs(12463) <= (layer0_outputs(4005)) xor (layer0_outputs(2856));
    outputs(12464) <= layer0_outputs(1905);
    outputs(12465) <= not((layer0_outputs(7431)) and (layer0_outputs(8381)));
    outputs(12466) <= not(layer0_outputs(3298));
    outputs(12467) <= (layer0_outputs(8409)) and not (layer0_outputs(11509));
    outputs(12468) <= layer0_outputs(6243);
    outputs(12469) <= (layer0_outputs(4715)) or (layer0_outputs(8238));
    outputs(12470) <= layer0_outputs(5297);
    outputs(12471) <= not((layer0_outputs(5199)) or (layer0_outputs(1891)));
    outputs(12472) <= not(layer0_outputs(1593));
    outputs(12473) <= not((layer0_outputs(11497)) and (layer0_outputs(5451)));
    outputs(12474) <= not(layer0_outputs(3475));
    outputs(12475) <= not((layer0_outputs(9880)) xor (layer0_outputs(593)));
    outputs(12476) <= not((layer0_outputs(8799)) or (layer0_outputs(3674)));
    outputs(12477) <= not(layer0_outputs(10208));
    outputs(12478) <= (layer0_outputs(10165)) xor (layer0_outputs(7673));
    outputs(12479) <= (layer0_outputs(2333)) and not (layer0_outputs(5467));
    outputs(12480) <= not(layer0_outputs(9052));
    outputs(12481) <= layer0_outputs(2766);
    outputs(12482) <= (layer0_outputs(4875)) and not (layer0_outputs(4466));
    outputs(12483) <= not(layer0_outputs(848));
    outputs(12484) <= (layer0_outputs(9873)) xor (layer0_outputs(12393));
    outputs(12485) <= not(layer0_outputs(3783));
    outputs(12486) <= layer0_outputs(12272);
    outputs(12487) <= not(layer0_outputs(8506));
    outputs(12488) <= (layer0_outputs(12181)) and not (layer0_outputs(12440));
    outputs(12489) <= layer0_outputs(9634);
    outputs(12490) <= not((layer0_outputs(647)) xor (layer0_outputs(5940)));
    outputs(12491) <= layer0_outputs(933);
    outputs(12492) <= (layer0_outputs(10483)) xor (layer0_outputs(9920));
    outputs(12493) <= (layer0_outputs(7872)) xor (layer0_outputs(4666));
    outputs(12494) <= layer0_outputs(6779);
    outputs(12495) <= not((layer0_outputs(7942)) xor (layer0_outputs(3573)));
    outputs(12496) <= not(layer0_outputs(2932));
    outputs(12497) <= layer0_outputs(7154);
    outputs(12498) <= (layer0_outputs(11690)) and not (layer0_outputs(1933));
    outputs(12499) <= layer0_outputs(3490);
    outputs(12500) <= not((layer0_outputs(5466)) xor (layer0_outputs(6185)));
    outputs(12501) <= not((layer0_outputs(3804)) xor (layer0_outputs(360)));
    outputs(12502) <= (layer0_outputs(384)) xor (layer0_outputs(3850));
    outputs(12503) <= layer0_outputs(2542);
    outputs(12504) <= (layer0_outputs(10420)) and not (layer0_outputs(1092));
    outputs(12505) <= not((layer0_outputs(6276)) or (layer0_outputs(8843)));
    outputs(12506) <= not((layer0_outputs(10183)) xor (layer0_outputs(5471)));
    outputs(12507) <= (layer0_outputs(2672)) xor (layer0_outputs(5489));
    outputs(12508) <= layer0_outputs(6949);
    outputs(12509) <= (layer0_outputs(4720)) xor (layer0_outputs(8528));
    outputs(12510) <= (layer0_outputs(8088)) xor (layer0_outputs(8467));
    outputs(12511) <= not((layer0_outputs(6015)) xor (layer0_outputs(2059)));
    outputs(12512) <= not(layer0_outputs(567));
    outputs(12513) <= layer0_outputs(3096);
    outputs(12514) <= layer0_outputs(1935);
    outputs(12515) <= not((layer0_outputs(11020)) xor (layer0_outputs(12665)));
    outputs(12516) <= (layer0_outputs(6116)) xor (layer0_outputs(2263));
    outputs(12517) <= (layer0_outputs(1476)) and not (layer0_outputs(1260));
    outputs(12518) <= not(layer0_outputs(4472));
    outputs(12519) <= not(layer0_outputs(4572));
    outputs(12520) <= layer0_outputs(1273);
    outputs(12521) <= (layer0_outputs(375)) and (layer0_outputs(523));
    outputs(12522) <= not((layer0_outputs(7641)) xor (layer0_outputs(4702)));
    outputs(12523) <= (layer0_outputs(8787)) xor (layer0_outputs(2165));
    outputs(12524) <= layer0_outputs(10130);
    outputs(12525) <= layer0_outputs(11444);
    outputs(12526) <= (layer0_outputs(6131)) or (layer0_outputs(4140));
    outputs(12527) <= not(layer0_outputs(9807));
    outputs(12528) <= not((layer0_outputs(12143)) xor (layer0_outputs(9708)));
    outputs(12529) <= not((layer0_outputs(1718)) and (layer0_outputs(1540)));
    outputs(12530) <= not(layer0_outputs(5053));
    outputs(12531) <= (layer0_outputs(5367)) xor (layer0_outputs(10643));
    outputs(12532) <= not((layer0_outputs(9379)) or (layer0_outputs(3404)));
    outputs(12533) <= not(layer0_outputs(4589));
    outputs(12534) <= (layer0_outputs(4643)) or (layer0_outputs(7765));
    outputs(12535) <= layer0_outputs(2792);
    outputs(12536) <= not((layer0_outputs(9617)) xor (layer0_outputs(4132)));
    outputs(12537) <= (layer0_outputs(6734)) xor (layer0_outputs(8020));
    outputs(12538) <= not((layer0_outputs(1264)) xor (layer0_outputs(2597)));
    outputs(12539) <= layer0_outputs(8838);
    outputs(12540) <= not(layer0_outputs(3796));
    outputs(12541) <= not(layer0_outputs(8979));
    outputs(12542) <= layer0_outputs(5449);
    outputs(12543) <= layer0_outputs(9990);
    outputs(12544) <= layer0_outputs(2247);
    outputs(12545) <= not(layer0_outputs(6645));
    outputs(12546) <= not(layer0_outputs(7459));
    outputs(12547) <= layer0_outputs(6736);
    outputs(12548) <= not((layer0_outputs(10765)) xor (layer0_outputs(1304)));
    outputs(12549) <= (layer0_outputs(4958)) and (layer0_outputs(7081));
    outputs(12550) <= (layer0_outputs(10337)) xor (layer0_outputs(3252));
    outputs(12551) <= not(layer0_outputs(12606));
    outputs(12552) <= layer0_outputs(8684);
    outputs(12553) <= not(layer0_outputs(1438));
    outputs(12554) <= layer0_outputs(915);
    outputs(12555) <= (layer0_outputs(814)) and not (layer0_outputs(733));
    outputs(12556) <= layer0_outputs(2968);
    outputs(12557) <= not((layer0_outputs(10983)) or (layer0_outputs(4704)));
    outputs(12558) <= not(layer0_outputs(3339));
    outputs(12559) <= (layer0_outputs(9206)) and not (layer0_outputs(7536));
    outputs(12560) <= (layer0_outputs(7326)) and (layer0_outputs(334));
    outputs(12561) <= not(layer0_outputs(513));
    outputs(12562) <= not(layer0_outputs(5562));
    outputs(12563) <= layer0_outputs(2411);
    outputs(12564) <= not((layer0_outputs(2526)) xor (layer0_outputs(5045)));
    outputs(12565) <= (layer0_outputs(12356)) xor (layer0_outputs(9074));
    outputs(12566) <= (layer0_outputs(6074)) or (layer0_outputs(7355));
    outputs(12567) <= not(layer0_outputs(5661));
    outputs(12568) <= (layer0_outputs(8816)) xor (layer0_outputs(2751));
    outputs(12569) <= (layer0_outputs(4199)) xor (layer0_outputs(3200));
    outputs(12570) <= (layer0_outputs(12457)) and not (layer0_outputs(6395));
    outputs(12571) <= not(layer0_outputs(7417));
    outputs(12572) <= not((layer0_outputs(2322)) xor (layer0_outputs(7996)));
    outputs(12573) <= not(layer0_outputs(11503)) or (layer0_outputs(4653));
    outputs(12574) <= layer0_outputs(8421);
    outputs(12575) <= layer0_outputs(3146);
    outputs(12576) <= layer0_outputs(9655);
    outputs(12577) <= not((layer0_outputs(1225)) xor (layer0_outputs(3394)));
    outputs(12578) <= not((layer0_outputs(1788)) xor (layer0_outputs(1382)));
    outputs(12579) <= not((layer0_outputs(12090)) xor (layer0_outputs(4646)));
    outputs(12580) <= not((layer0_outputs(762)) or (layer0_outputs(2716)));
    outputs(12581) <= not(layer0_outputs(8615));
    outputs(12582) <= not(layer0_outputs(8009));
    outputs(12583) <= not((layer0_outputs(7805)) or (layer0_outputs(2024)));
    outputs(12584) <= not(layer0_outputs(6270));
    outputs(12585) <= (layer0_outputs(7467)) and not (layer0_outputs(1342));
    outputs(12586) <= (layer0_outputs(6747)) xor (layer0_outputs(4445));
    outputs(12587) <= (layer0_outputs(5029)) and not (layer0_outputs(9405));
    outputs(12588) <= layer0_outputs(952);
    outputs(12589) <= (layer0_outputs(6496)) xor (layer0_outputs(4493));
    outputs(12590) <= not((layer0_outputs(8993)) xor (layer0_outputs(2967)));
    outputs(12591) <= not(layer0_outputs(12730));
    outputs(12592) <= not(layer0_outputs(2036));
    outputs(12593) <= not(layer0_outputs(6143));
    outputs(12594) <= layer0_outputs(1365);
    outputs(12595) <= layer0_outputs(11075);
    outputs(12596) <= (layer0_outputs(6422)) and (layer0_outputs(3513));
    outputs(12597) <= layer0_outputs(1464);
    outputs(12598) <= not((layer0_outputs(6798)) xor (layer0_outputs(2421)));
    outputs(12599) <= not((layer0_outputs(9448)) xor (layer0_outputs(6253)));
    outputs(12600) <= not((layer0_outputs(9309)) or (layer0_outputs(1258)));
    outputs(12601) <= not((layer0_outputs(6855)) xor (layer0_outputs(11693)));
    outputs(12602) <= (layer0_outputs(4058)) xor (layer0_outputs(1122));
    outputs(12603) <= not(layer0_outputs(3861));
    outputs(12604) <= (layer0_outputs(6047)) and not (layer0_outputs(10236));
    outputs(12605) <= (layer0_outputs(12085)) and not (layer0_outputs(2012));
    outputs(12606) <= not(layer0_outputs(8451));
    outputs(12607) <= not(layer0_outputs(9065));
    outputs(12608) <= (layer0_outputs(5134)) and not (layer0_outputs(5047));
    outputs(12609) <= not((layer0_outputs(6136)) or (layer0_outputs(12359)));
    outputs(12610) <= not(layer0_outputs(12070)) or (layer0_outputs(3003));
    outputs(12611) <= not((layer0_outputs(3746)) and (layer0_outputs(2946)));
    outputs(12612) <= layer0_outputs(4930);
    outputs(12613) <= layer0_outputs(10724);
    outputs(12614) <= not(layer0_outputs(11947));
    outputs(12615) <= (layer0_outputs(9471)) and not (layer0_outputs(9228));
    outputs(12616) <= (layer0_outputs(2015)) and (layer0_outputs(2658));
    outputs(12617) <= not(layer0_outputs(1686));
    outputs(12618) <= not(layer0_outputs(2661));
    outputs(12619) <= layer0_outputs(3477);
    outputs(12620) <= layer0_outputs(9699);
    outputs(12621) <= (layer0_outputs(2323)) and not (layer0_outputs(6871));
    outputs(12622) <= not(layer0_outputs(11101)) or (layer0_outputs(10397));
    outputs(12623) <= (layer0_outputs(58)) and not (layer0_outputs(4867));
    outputs(12624) <= not(layer0_outputs(5694));
    outputs(12625) <= (layer0_outputs(2225)) and not (layer0_outputs(5517));
    outputs(12626) <= not(layer0_outputs(4542));
    outputs(12627) <= not(layer0_outputs(11153));
    outputs(12628) <= (layer0_outputs(3498)) and (layer0_outputs(3556));
    outputs(12629) <= (layer0_outputs(9872)) xor (layer0_outputs(12745));
    outputs(12630) <= layer0_outputs(10557);
    outputs(12631) <= not((layer0_outputs(6002)) xor (layer0_outputs(4524)));
    outputs(12632) <= not(layer0_outputs(8604));
    outputs(12633) <= not((layer0_outputs(1536)) and (layer0_outputs(5309)));
    outputs(12634) <= not((layer0_outputs(612)) and (layer0_outputs(7271)));
    outputs(12635) <= not((layer0_outputs(11546)) xor (layer0_outputs(12504)));
    outputs(12636) <= not(layer0_outputs(1873));
    outputs(12637) <= not(layer0_outputs(10118));
    outputs(12638) <= (layer0_outputs(6073)) xor (layer0_outputs(6056));
    outputs(12639) <= not((layer0_outputs(6457)) xor (layer0_outputs(10588)));
    outputs(12640) <= (layer0_outputs(983)) xor (layer0_outputs(11908));
    outputs(12641) <= layer0_outputs(6101);
    outputs(12642) <= (layer0_outputs(8063)) and not (layer0_outputs(10892));
    outputs(12643) <= layer0_outputs(5218);
    outputs(12644) <= (layer0_outputs(7766)) or (layer0_outputs(6888));
    outputs(12645) <= not((layer0_outputs(6946)) xor (layer0_outputs(12260)));
    outputs(12646) <= (layer0_outputs(5249)) xor (layer0_outputs(11273));
    outputs(12647) <= not(layer0_outputs(1881));
    outputs(12648) <= layer0_outputs(4433);
    outputs(12649) <= layer0_outputs(7883);
    outputs(12650) <= not(layer0_outputs(4970));
    outputs(12651) <= layer0_outputs(2135);
    outputs(12652) <= not(layer0_outputs(5853));
    outputs(12653) <= not(layer0_outputs(7923));
    outputs(12654) <= (layer0_outputs(10159)) and not (layer0_outputs(9175));
    outputs(12655) <= (layer0_outputs(3299)) xor (layer0_outputs(5629));
    outputs(12656) <= (layer0_outputs(4976)) and not (layer0_outputs(1752));
    outputs(12657) <= not((layer0_outputs(4424)) xor (layer0_outputs(11299)));
    outputs(12658) <= not((layer0_outputs(604)) xor (layer0_outputs(980)));
    outputs(12659) <= (layer0_outputs(8263)) xor (layer0_outputs(3560));
    outputs(12660) <= not((layer0_outputs(2424)) and (layer0_outputs(6548)));
    outputs(12661) <= (layer0_outputs(2138)) and (layer0_outputs(4463));
    outputs(12662) <= layer0_outputs(12549);
    outputs(12663) <= not(layer0_outputs(4879));
    outputs(12664) <= layer0_outputs(5072);
    outputs(12665) <= not((layer0_outputs(12763)) xor (layer0_outputs(11475)));
    outputs(12666) <= not(layer0_outputs(6902));
    outputs(12667) <= (layer0_outputs(1230)) and (layer0_outputs(556));
    outputs(12668) <= (layer0_outputs(12699)) or (layer0_outputs(11114));
    outputs(12669) <= not((layer0_outputs(10972)) xor (layer0_outputs(7056)));
    outputs(12670) <= not(layer0_outputs(35));
    outputs(12671) <= (layer0_outputs(4826)) and (layer0_outputs(11682));
    outputs(12672) <= not(layer0_outputs(7402));
    outputs(12673) <= (layer0_outputs(2196)) xor (layer0_outputs(12018));
    outputs(12674) <= (layer0_outputs(12410)) xor (layer0_outputs(5577));
    outputs(12675) <= (layer0_outputs(12060)) and not (layer0_outputs(11036));
    outputs(12676) <= (layer0_outputs(8062)) xor (layer0_outputs(9804));
    outputs(12677) <= not((layer0_outputs(10092)) or (layer0_outputs(8231)));
    outputs(12678) <= not((layer0_outputs(7282)) or (layer0_outputs(7255)));
    outputs(12679) <= (layer0_outputs(11615)) or (layer0_outputs(10617));
    outputs(12680) <= not(layer0_outputs(1838));
    outputs(12681) <= (layer0_outputs(6225)) or (layer0_outputs(7042));
    outputs(12682) <= (layer0_outputs(1053)) and not (layer0_outputs(9364));
    outputs(12683) <= (layer0_outputs(2085)) or (layer0_outputs(1238));
    outputs(12684) <= not(layer0_outputs(6531));
    outputs(12685) <= (layer0_outputs(4483)) or (layer0_outputs(4783));
    outputs(12686) <= (layer0_outputs(4987)) and (layer0_outputs(4857));
    outputs(12687) <= not(layer0_outputs(4970));
    outputs(12688) <= (layer0_outputs(10221)) xor (layer0_outputs(660));
    outputs(12689) <= (layer0_outputs(3403)) xor (layer0_outputs(2057));
    outputs(12690) <= not((layer0_outputs(7528)) xor (layer0_outputs(10859)));
    outputs(12691) <= not(layer0_outputs(7827)) or (layer0_outputs(10566));
    outputs(12692) <= layer0_outputs(11725);
    outputs(12693) <= not((layer0_outputs(12696)) xor (layer0_outputs(8160)));
    outputs(12694) <= layer0_outputs(10615);
    outputs(12695) <= (layer0_outputs(12232)) and not (layer0_outputs(2184));
    outputs(12696) <= (layer0_outputs(9555)) xor (layer0_outputs(6499));
    outputs(12697) <= (layer0_outputs(10540)) and not (layer0_outputs(12421));
    outputs(12698) <= (layer0_outputs(5860)) xor (layer0_outputs(12119));
    outputs(12699) <= not(layer0_outputs(9368)) or (layer0_outputs(2158));
    outputs(12700) <= not(layer0_outputs(4484));
    outputs(12701) <= (layer0_outputs(5747)) xor (layer0_outputs(4767));
    outputs(12702) <= not((layer0_outputs(12331)) or (layer0_outputs(368)));
    outputs(12703) <= (layer0_outputs(2822)) xor (layer0_outputs(1023));
    outputs(12704) <= not((layer0_outputs(6933)) or (layer0_outputs(3826)));
    outputs(12705) <= layer0_outputs(2496);
    outputs(12706) <= not((layer0_outputs(5119)) xor (layer0_outputs(3163)));
    outputs(12707) <= (layer0_outputs(3824)) xor (layer0_outputs(7241));
    outputs(12708) <= not((layer0_outputs(9230)) xor (layer0_outputs(1136)));
    outputs(12709) <= layer0_outputs(2003);
    outputs(12710) <= layer0_outputs(5366);
    outputs(12711) <= not(layer0_outputs(4457));
    outputs(12712) <= not(layer0_outputs(7262));
    outputs(12713) <= (layer0_outputs(10722)) or (layer0_outputs(5378));
    outputs(12714) <= not((layer0_outputs(10010)) or (layer0_outputs(12472)));
    outputs(12715) <= (layer0_outputs(1529)) and not (layer0_outputs(3672));
    outputs(12716) <= (layer0_outputs(9520)) and (layer0_outputs(10353));
    outputs(12717) <= not((layer0_outputs(3546)) or (layer0_outputs(9672)));
    outputs(12718) <= (layer0_outputs(11877)) and not (layer0_outputs(1126));
    outputs(12719) <= (layer0_outputs(4391)) xor (layer0_outputs(4453));
    outputs(12720) <= not((layer0_outputs(8526)) or (layer0_outputs(11139)));
    outputs(12721) <= (layer0_outputs(972)) xor (layer0_outputs(2725));
    outputs(12722) <= (layer0_outputs(535)) or (layer0_outputs(11025));
    outputs(12723) <= not(layer0_outputs(5775));
    outputs(12724) <= layer0_outputs(7483);
    outputs(12725) <= not(layer0_outputs(9286));
    outputs(12726) <= layer0_outputs(6057);
    outputs(12727) <= layer0_outputs(7398);
    outputs(12728) <= layer0_outputs(11294);
    outputs(12729) <= (layer0_outputs(9234)) xor (layer0_outputs(9725));
    outputs(12730) <= layer0_outputs(10759);
    outputs(12731) <= layer0_outputs(413);
    outputs(12732) <= not((layer0_outputs(8266)) or (layer0_outputs(3658)));
    outputs(12733) <= not(layer0_outputs(7105));
    outputs(12734) <= (layer0_outputs(7388)) and not (layer0_outputs(7848));
    outputs(12735) <= layer0_outputs(8983);
    outputs(12736) <= (layer0_outputs(4313)) xor (layer0_outputs(7488));
    outputs(12737) <= (layer0_outputs(3698)) and (layer0_outputs(5902));
    outputs(12738) <= (layer0_outputs(6796)) xor (layer0_outputs(7055));
    outputs(12739) <= (layer0_outputs(5979)) or (layer0_outputs(2763));
    outputs(12740) <= (layer0_outputs(12570)) and (layer0_outputs(3981));
    outputs(12741) <= layer0_outputs(957);
    outputs(12742) <= (layer0_outputs(5072)) and not (layer0_outputs(3040));
    outputs(12743) <= layer0_outputs(286);
    outputs(12744) <= not((layer0_outputs(1818)) xor (layer0_outputs(12567)));
    outputs(12745) <= layer0_outputs(740);
    outputs(12746) <= (layer0_outputs(9326)) and not (layer0_outputs(3265));
    outputs(12747) <= (layer0_outputs(8780)) xor (layer0_outputs(7731));
    outputs(12748) <= layer0_outputs(999);
    outputs(12749) <= not(layer0_outputs(2583));
    outputs(12750) <= (layer0_outputs(4176)) and not (layer0_outputs(5634));
    outputs(12751) <= not(layer0_outputs(12557));
    outputs(12752) <= not(layer0_outputs(10502));
    outputs(12753) <= (layer0_outputs(1321)) and not (layer0_outputs(4387));
    outputs(12754) <= not((layer0_outputs(1899)) or (layer0_outputs(12210)));
    outputs(12755) <= (layer0_outputs(63)) and (layer0_outputs(12347));
    outputs(12756) <= not((layer0_outputs(3717)) xor (layer0_outputs(9504)));
    outputs(12757) <= (layer0_outputs(12378)) and (layer0_outputs(3250));
    outputs(12758) <= (layer0_outputs(1490)) xor (layer0_outputs(10621));
    outputs(12759) <= not(layer0_outputs(6113));
    outputs(12760) <= layer0_outputs(7177);
    outputs(12761) <= (layer0_outputs(6657)) and not (layer0_outputs(505));
    outputs(12762) <= not((layer0_outputs(2481)) or (layer0_outputs(5728)));
    outputs(12763) <= not(layer0_outputs(5549));
    outputs(12764) <= not(layer0_outputs(5204));
    outputs(12765) <= not(layer0_outputs(4978));
    outputs(12766) <= not(layer0_outputs(10367));
    outputs(12767) <= not(layer0_outputs(3361));
    outputs(12768) <= not(layer0_outputs(548));
    outputs(12769) <= (layer0_outputs(634)) xor (layer0_outputs(11865));
    outputs(12770) <= not((layer0_outputs(4995)) xor (layer0_outputs(6693)));
    outputs(12771) <= not(layer0_outputs(6556));
    outputs(12772) <= (layer0_outputs(5806)) xor (layer0_outputs(8127));
    outputs(12773) <= not((layer0_outputs(6458)) and (layer0_outputs(4)));
    outputs(12774) <= layer0_outputs(10981);
    outputs(12775) <= (layer0_outputs(4130)) xor (layer0_outputs(9697));
    outputs(12776) <= layer0_outputs(10996);
    outputs(12777) <= not(layer0_outputs(10140));
    outputs(12778) <= (layer0_outputs(3302)) and not (layer0_outputs(2055));
    outputs(12779) <= not((layer0_outputs(9122)) or (layer0_outputs(616)));
    outputs(12780) <= not(layer0_outputs(9607));
    outputs(12781) <= layer0_outputs(4054);
    outputs(12782) <= not(layer0_outputs(8469));
    outputs(12783) <= not((layer0_outputs(9898)) xor (layer0_outputs(1001)));
    outputs(12784) <= not(layer0_outputs(12607));
    outputs(12785) <= (layer0_outputs(3018)) xor (layer0_outputs(9979));
    outputs(12786) <= not(layer0_outputs(11758)) or (layer0_outputs(5338));
    outputs(12787) <= layer0_outputs(6623);
    outputs(12788) <= layer0_outputs(6454);
    outputs(12789) <= not((layer0_outputs(5096)) xor (layer0_outputs(2430)));
    outputs(12790) <= not(layer0_outputs(9056));
    outputs(12791) <= not(layer0_outputs(2521));
    outputs(12792) <= not(layer0_outputs(10376));
    outputs(12793) <= not((layer0_outputs(7653)) xor (layer0_outputs(11741)));
    outputs(12794) <= not((layer0_outputs(10289)) or (layer0_outputs(8350)));
    outputs(12795) <= layer0_outputs(4537);
    outputs(12796) <= not(layer0_outputs(3261));
    outputs(12797) <= layer0_outputs(12795);
    outputs(12798) <= (layer0_outputs(6509)) xor (layer0_outputs(373));
    outputs(12799) <= layer0_outputs(5574);

end Behavioral;
