library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(7679 downto 0);

begin

    layer0_outputs(0) <= (inputs(48)) xor (inputs(140));
    layer0_outputs(1) <= not(inputs(92));
    layer0_outputs(2) <= (inputs(91)) or (inputs(249));
    layer0_outputs(3) <= inputs(42);
    layer0_outputs(4) <= (inputs(152)) and not (inputs(115));
    layer0_outputs(5) <= inputs(22);
    layer0_outputs(6) <= inputs(103);
    layer0_outputs(7) <= not(inputs(145));
    layer0_outputs(8) <= (inputs(137)) xor (inputs(17));
    layer0_outputs(9) <= not(inputs(75)) or (inputs(39));
    layer0_outputs(10) <= not((inputs(85)) xor (inputs(226)));
    layer0_outputs(11) <= not(inputs(89)) or (inputs(16));
    layer0_outputs(12) <= not(inputs(12)) or (inputs(238));
    layer0_outputs(13) <= inputs(24);
    layer0_outputs(14) <= '1';
    layer0_outputs(15) <= (inputs(23)) and not (inputs(160));
    layer0_outputs(16) <= inputs(19);
    layer0_outputs(17) <= not(inputs(179)) or (inputs(88));
    layer0_outputs(18) <= not(inputs(54));
    layer0_outputs(19) <= not(inputs(100));
    layer0_outputs(20) <= not(inputs(139));
    layer0_outputs(21) <= not((inputs(107)) xor (inputs(76)));
    layer0_outputs(22) <= (inputs(200)) xor (inputs(20));
    layer0_outputs(23) <= not((inputs(96)) or (inputs(202)));
    layer0_outputs(24) <= inputs(117);
    layer0_outputs(25) <= (inputs(223)) and not (inputs(126));
    layer0_outputs(26) <= not(inputs(168));
    layer0_outputs(27) <= not(inputs(202)) or (inputs(29));
    layer0_outputs(28) <= (inputs(76)) or (inputs(164));
    layer0_outputs(29) <= (inputs(55)) and not (inputs(100));
    layer0_outputs(30) <= not(inputs(182));
    layer0_outputs(31) <= inputs(31);
    layer0_outputs(32) <= not(inputs(70));
    layer0_outputs(33) <= not((inputs(167)) or (inputs(30)));
    layer0_outputs(34) <= (inputs(101)) or (inputs(107));
    layer0_outputs(35) <= (inputs(208)) and not (inputs(79));
    layer0_outputs(36) <= not((inputs(75)) or (inputs(52)));
    layer0_outputs(37) <= (inputs(220)) and not (inputs(53));
    layer0_outputs(38) <= (inputs(118)) xor (inputs(6));
    layer0_outputs(39) <= '0';
    layer0_outputs(40) <= inputs(130);
    layer0_outputs(41) <= inputs(43);
    layer0_outputs(42) <= inputs(124);
    layer0_outputs(43) <= not(inputs(93));
    layer0_outputs(44) <= (inputs(137)) and (inputs(183));
    layer0_outputs(45) <= (inputs(234)) or (inputs(166));
    layer0_outputs(46) <= not(inputs(70));
    layer0_outputs(47) <= not(inputs(219)) or (inputs(235));
    layer0_outputs(48) <= inputs(93);
    layer0_outputs(49) <= not((inputs(25)) or (inputs(110)));
    layer0_outputs(50) <= not(inputs(105));
    layer0_outputs(51) <= not(inputs(121)) or (inputs(19));
    layer0_outputs(52) <= (inputs(179)) xor (inputs(34));
    layer0_outputs(53) <= not(inputs(189));
    layer0_outputs(54) <= (inputs(108)) and not (inputs(132));
    layer0_outputs(55) <= (inputs(35)) and not (inputs(59));
    layer0_outputs(56) <= (inputs(243)) or (inputs(104));
    layer0_outputs(57) <= inputs(234);
    layer0_outputs(58) <= not((inputs(134)) or (inputs(14)));
    layer0_outputs(59) <= '0';
    layer0_outputs(60) <= not(inputs(203)) or (inputs(236));
    layer0_outputs(61) <= (inputs(62)) xor (inputs(68));
    layer0_outputs(62) <= inputs(149);
    layer0_outputs(63) <= (inputs(40)) or (inputs(135));
    layer0_outputs(64) <= inputs(42);
    layer0_outputs(65) <= (inputs(106)) or (inputs(128));
    layer0_outputs(66) <= not(inputs(114));
    layer0_outputs(67) <= (inputs(24)) and not (inputs(159));
    layer0_outputs(68) <= not((inputs(104)) or (inputs(144)));
    layer0_outputs(69) <= (inputs(147)) and not (inputs(252));
    layer0_outputs(70) <= (inputs(92)) xor (inputs(27));
    layer0_outputs(71) <= not(inputs(141));
    layer0_outputs(72) <= not(inputs(71)) or (inputs(110));
    layer0_outputs(73) <= not(inputs(21));
    layer0_outputs(74) <= '0';
    layer0_outputs(75) <= (inputs(243)) and not (inputs(11));
    layer0_outputs(76) <= (inputs(92)) xor (inputs(90));
    layer0_outputs(77) <= (inputs(248)) or (inputs(138));
    layer0_outputs(78) <= (inputs(74)) and (inputs(46));
    layer0_outputs(79) <= inputs(211);
    layer0_outputs(80) <= inputs(233);
    layer0_outputs(81) <= not(inputs(117)) or (inputs(193));
    layer0_outputs(82) <= not(inputs(42)) or (inputs(63));
    layer0_outputs(83) <= not((inputs(163)) or (inputs(178)));
    layer0_outputs(84) <= (inputs(204)) or (inputs(115));
    layer0_outputs(85) <= (inputs(141)) xor (inputs(230));
    layer0_outputs(86) <= (inputs(45)) and not (inputs(140));
    layer0_outputs(87) <= not(inputs(167)) or (inputs(231));
    layer0_outputs(88) <= not((inputs(182)) or (inputs(14)));
    layer0_outputs(89) <= (inputs(176)) xor (inputs(103));
    layer0_outputs(90) <= inputs(180);
    layer0_outputs(91) <= (inputs(108)) and not (inputs(241));
    layer0_outputs(92) <= not((inputs(128)) xor (inputs(225)));
    layer0_outputs(93) <= not(inputs(121)) or (inputs(162));
    layer0_outputs(94) <= not(inputs(117));
    layer0_outputs(95) <= inputs(119);
    layer0_outputs(96) <= '1';
    layer0_outputs(97) <= '0';
    layer0_outputs(98) <= (inputs(196)) and not (inputs(177));
    layer0_outputs(99) <= not((inputs(105)) xor (inputs(91)));
    layer0_outputs(100) <= (inputs(104)) or (inputs(235));
    layer0_outputs(101) <= not((inputs(132)) xor (inputs(18)));
    layer0_outputs(102) <= not(inputs(149)) or (inputs(236));
    layer0_outputs(103) <= inputs(116);
    layer0_outputs(104) <= (inputs(60)) xor (inputs(14));
    layer0_outputs(105) <= not(inputs(236)) or (inputs(36));
    layer0_outputs(106) <= not(inputs(90)) or (inputs(165));
    layer0_outputs(107) <= not(inputs(88));
    layer0_outputs(108) <= not((inputs(164)) xor (inputs(226)));
    layer0_outputs(109) <= (inputs(228)) or (inputs(69));
    layer0_outputs(110) <= (inputs(153)) or (inputs(250));
    layer0_outputs(111) <= '0';
    layer0_outputs(112) <= not(inputs(172));
    layer0_outputs(113) <= inputs(62);
    layer0_outputs(114) <= inputs(168);
    layer0_outputs(115) <= (inputs(146)) or (inputs(23));
    layer0_outputs(116) <= (inputs(92)) and not (inputs(207));
    layer0_outputs(117) <= (inputs(72)) and not (inputs(48));
    layer0_outputs(118) <= not(inputs(163));
    layer0_outputs(119) <= not(inputs(155));
    layer0_outputs(120) <= (inputs(85)) or (inputs(97));
    layer0_outputs(121) <= (inputs(36)) or (inputs(209));
    layer0_outputs(122) <= not(inputs(167)) or (inputs(62));
    layer0_outputs(123) <= (inputs(161)) and (inputs(89));
    layer0_outputs(124) <= not(inputs(37));
    layer0_outputs(125) <= (inputs(28)) or (inputs(174));
    layer0_outputs(126) <= not((inputs(81)) or (inputs(104)));
    layer0_outputs(127) <= not(inputs(122)) or (inputs(63));
    layer0_outputs(128) <= (inputs(14)) or (inputs(16));
    layer0_outputs(129) <= (inputs(150)) and not (inputs(210));
    layer0_outputs(130) <= not(inputs(87)) or (inputs(61));
    layer0_outputs(131) <= inputs(46);
    layer0_outputs(132) <= inputs(104);
    layer0_outputs(133) <= (inputs(45)) or (inputs(67));
    layer0_outputs(134) <= (inputs(101)) xor (inputs(202));
    layer0_outputs(135) <= not(inputs(125));
    layer0_outputs(136) <= (inputs(212)) and not (inputs(253));
    layer0_outputs(137) <= (inputs(55)) or (inputs(118));
    layer0_outputs(138) <= not((inputs(172)) xor (inputs(205)));
    layer0_outputs(139) <= not((inputs(58)) and (inputs(24)));
    layer0_outputs(140) <= inputs(246);
    layer0_outputs(141) <= not(inputs(16));
    layer0_outputs(142) <= (inputs(11)) or (inputs(183));
    layer0_outputs(143) <= not((inputs(153)) and (inputs(106)));
    layer0_outputs(144) <= not((inputs(203)) or (inputs(49)));
    layer0_outputs(145) <= not((inputs(39)) or (inputs(206)));
    layer0_outputs(146) <= not(inputs(186));
    layer0_outputs(147) <= not(inputs(88)) or (inputs(126));
    layer0_outputs(148) <= (inputs(104)) xor (inputs(155));
    layer0_outputs(149) <= inputs(211);
    layer0_outputs(150) <= (inputs(206)) xor (inputs(230));
    layer0_outputs(151) <= not((inputs(208)) and (inputs(34)));
    layer0_outputs(152) <= (inputs(55)) or (inputs(75));
    layer0_outputs(153) <= (inputs(180)) or (inputs(126));
    layer0_outputs(154) <= (inputs(136)) and not (inputs(68));
    layer0_outputs(155) <= not((inputs(24)) xor (inputs(40)));
    layer0_outputs(156) <= not(inputs(180)) or (inputs(65));
    layer0_outputs(157) <= not(inputs(136));
    layer0_outputs(158) <= not((inputs(242)) xor (inputs(10)));
    layer0_outputs(159) <= inputs(84);
    layer0_outputs(160) <= not(inputs(145)) or (inputs(178));
    layer0_outputs(161) <= not((inputs(242)) or (inputs(144)));
    layer0_outputs(162) <= not(inputs(56)) or (inputs(228));
    layer0_outputs(163) <= not((inputs(186)) xor (inputs(238)));
    layer0_outputs(164) <= not(inputs(248)) or (inputs(79));
    layer0_outputs(165) <= not(inputs(52)) or (inputs(7));
    layer0_outputs(166) <= (inputs(243)) and not (inputs(7));
    layer0_outputs(167) <= inputs(239);
    layer0_outputs(168) <= (inputs(148)) and not (inputs(99));
    layer0_outputs(169) <= (inputs(74)) or (inputs(2));
    layer0_outputs(170) <= not(inputs(243)) or (inputs(203));
    layer0_outputs(171) <= not((inputs(94)) or (inputs(56)));
    layer0_outputs(172) <= not(inputs(105)) or (inputs(132));
    layer0_outputs(173) <= (inputs(195)) and (inputs(222));
    layer0_outputs(174) <= not(inputs(252));
    layer0_outputs(175) <= not(inputs(59));
    layer0_outputs(176) <= not((inputs(161)) or (inputs(223)));
    layer0_outputs(177) <= not((inputs(183)) or (inputs(25)));
    layer0_outputs(178) <= not(inputs(185));
    layer0_outputs(179) <= (inputs(10)) xor (inputs(25));
    layer0_outputs(180) <= inputs(100);
    layer0_outputs(181) <= (inputs(219)) xor (inputs(17));
    layer0_outputs(182) <= not(inputs(85)) or (inputs(21));
    layer0_outputs(183) <= (inputs(26)) xor (inputs(134));
    layer0_outputs(184) <= (inputs(188)) xor (inputs(253));
    layer0_outputs(185) <= '1';
    layer0_outputs(186) <= not(inputs(151));
    layer0_outputs(187) <= not(inputs(136)) or (inputs(64));
    layer0_outputs(188) <= (inputs(49)) and not (inputs(232));
    layer0_outputs(189) <= (inputs(106)) xor (inputs(50));
    layer0_outputs(190) <= not((inputs(216)) xor (inputs(23)));
    layer0_outputs(191) <= (inputs(202)) and (inputs(37));
    layer0_outputs(192) <= not((inputs(175)) xor (inputs(57)));
    layer0_outputs(193) <= not(inputs(218));
    layer0_outputs(194) <= inputs(226);
    layer0_outputs(195) <= inputs(238);
    layer0_outputs(196) <= inputs(182);
    layer0_outputs(197) <= not(inputs(83));
    layer0_outputs(198) <= (inputs(122)) xor (inputs(251));
    layer0_outputs(199) <= (inputs(210)) and not (inputs(62));
    layer0_outputs(200) <= not(inputs(36));
    layer0_outputs(201) <= not(inputs(105)) or (inputs(52));
    layer0_outputs(202) <= (inputs(153)) or (inputs(14));
    layer0_outputs(203) <= not(inputs(164)) or (inputs(220));
    layer0_outputs(204) <= (inputs(188)) and not (inputs(253));
    layer0_outputs(205) <= (inputs(63)) and not (inputs(97));
    layer0_outputs(206) <= not((inputs(225)) or (inputs(85)));
    layer0_outputs(207) <= not(inputs(255));
    layer0_outputs(208) <= (inputs(35)) xor (inputs(69));
    layer0_outputs(209) <= '1';
    layer0_outputs(210) <= not((inputs(207)) and (inputs(250)));
    layer0_outputs(211) <= (inputs(98)) or (inputs(168));
    layer0_outputs(212) <= not((inputs(191)) or (inputs(21)));
    layer0_outputs(213) <= not(inputs(119)) or (inputs(245));
    layer0_outputs(214) <= not((inputs(33)) xor (inputs(41)));
    layer0_outputs(215) <= not((inputs(118)) xor (inputs(158)));
    layer0_outputs(216) <= (inputs(40)) xor (inputs(173));
    layer0_outputs(217) <= (inputs(6)) or (inputs(137));
    layer0_outputs(218) <= '1';
    layer0_outputs(219) <= inputs(197);
    layer0_outputs(220) <= (inputs(193)) and not (inputs(2));
    layer0_outputs(221) <= not(inputs(106));
    layer0_outputs(222) <= not((inputs(171)) xor (inputs(220)));
    layer0_outputs(223) <= inputs(42);
    layer0_outputs(224) <= not(inputs(119));
    layer0_outputs(225) <= inputs(178);
    layer0_outputs(226) <= not((inputs(21)) or (inputs(189)));
    layer0_outputs(227) <= not(inputs(57)) or (inputs(53));
    layer0_outputs(228) <= not(inputs(135));
    layer0_outputs(229) <= (inputs(134)) or (inputs(224));
    layer0_outputs(230) <= '1';
    layer0_outputs(231) <= not(inputs(131)) or (inputs(142));
    layer0_outputs(232) <= (inputs(136)) and not (inputs(159));
    layer0_outputs(233) <= inputs(212);
    layer0_outputs(234) <= not(inputs(10)) or (inputs(159));
    layer0_outputs(235) <= inputs(43);
    layer0_outputs(236) <= not(inputs(101));
    layer0_outputs(237) <= (inputs(11)) and not (inputs(31));
    layer0_outputs(238) <= inputs(220);
    layer0_outputs(239) <= (inputs(233)) or (inputs(254));
    layer0_outputs(240) <= not(inputs(124)) or (inputs(110));
    layer0_outputs(241) <= not((inputs(233)) or (inputs(171)));
    layer0_outputs(242) <= not(inputs(125));
    layer0_outputs(243) <= not(inputs(117)) or (inputs(42));
    layer0_outputs(244) <= not((inputs(48)) xor (inputs(123)));
    layer0_outputs(245) <= '1';
    layer0_outputs(246) <= inputs(94);
    layer0_outputs(247) <= not((inputs(212)) or (inputs(176)));
    layer0_outputs(248) <= inputs(132);
    layer0_outputs(249) <= not(inputs(60)) or (inputs(227));
    layer0_outputs(250) <= not(inputs(231));
    layer0_outputs(251) <= (inputs(4)) xor (inputs(142));
    layer0_outputs(252) <= not(inputs(9)) or (inputs(97));
    layer0_outputs(253) <= not(inputs(166));
    layer0_outputs(254) <= not(inputs(35)) or (inputs(29));
    layer0_outputs(255) <= (inputs(103)) or (inputs(24));
    layer0_outputs(256) <= not(inputs(160));
    layer0_outputs(257) <= not(inputs(79));
    layer0_outputs(258) <= (inputs(73)) and (inputs(39));
    layer0_outputs(259) <= '1';
    layer0_outputs(260) <= not(inputs(41));
    layer0_outputs(261) <= not((inputs(228)) xor (inputs(213)));
    layer0_outputs(262) <= not(inputs(62)) or (inputs(239));
    layer0_outputs(263) <= not(inputs(122));
    layer0_outputs(264) <= (inputs(25)) xor (inputs(204));
    layer0_outputs(265) <= not(inputs(173)) or (inputs(252));
    layer0_outputs(266) <= not(inputs(218));
    layer0_outputs(267) <= not((inputs(72)) and (inputs(69)));
    layer0_outputs(268) <= not((inputs(255)) or (inputs(159)));
    layer0_outputs(269) <= (inputs(204)) or (inputs(55));
    layer0_outputs(270) <= not(inputs(138)) or (inputs(61));
    layer0_outputs(271) <= not((inputs(204)) or (inputs(132)));
    layer0_outputs(272) <= (inputs(254)) and not (inputs(23));
    layer0_outputs(273) <= not(inputs(61)) or (inputs(225));
    layer0_outputs(274) <= (inputs(153)) or (inputs(176));
    layer0_outputs(275) <= '0';
    layer0_outputs(276) <= not(inputs(57)) or (inputs(68));
    layer0_outputs(277) <= (inputs(23)) or (inputs(119));
    layer0_outputs(278) <= (inputs(249)) xor (inputs(144));
    layer0_outputs(279) <= not((inputs(190)) xor (inputs(77)));
    layer0_outputs(280) <= (inputs(77)) xor (inputs(247));
    layer0_outputs(281) <= not(inputs(82)) or (inputs(239));
    layer0_outputs(282) <= (inputs(69)) and not (inputs(232));
    layer0_outputs(283) <= not(inputs(122)) or (inputs(207));
    layer0_outputs(284) <= not(inputs(101));
    layer0_outputs(285) <= inputs(136);
    layer0_outputs(286) <= (inputs(107)) xor (inputs(209));
    layer0_outputs(287) <= (inputs(230)) and not (inputs(93));
    layer0_outputs(288) <= (inputs(234)) xor (inputs(69));
    layer0_outputs(289) <= (inputs(91)) and not (inputs(180));
    layer0_outputs(290) <= not(inputs(152)) or (inputs(11));
    layer0_outputs(291) <= not((inputs(165)) or (inputs(117)));
    layer0_outputs(292) <= inputs(176);
    layer0_outputs(293) <= not(inputs(197)) or (inputs(100));
    layer0_outputs(294) <= not((inputs(67)) and (inputs(145)));
    layer0_outputs(295) <= not(inputs(194));
    layer0_outputs(296) <= not(inputs(213)) or (inputs(61));
    layer0_outputs(297) <= not((inputs(108)) or (inputs(233)));
    layer0_outputs(298) <= not((inputs(115)) xor (inputs(192)));
    layer0_outputs(299) <= (inputs(235)) and not (inputs(79));
    layer0_outputs(300) <= (inputs(125)) or (inputs(115));
    layer0_outputs(301) <= inputs(39);
    layer0_outputs(302) <= not((inputs(174)) or (inputs(211)));
    layer0_outputs(303) <= not(inputs(114)) or (inputs(7));
    layer0_outputs(304) <= (inputs(151)) or (inputs(67));
    layer0_outputs(305) <= (inputs(53)) or (inputs(63));
    layer0_outputs(306) <= not((inputs(79)) or (inputs(169)));
    layer0_outputs(307) <= not(inputs(116));
    layer0_outputs(308) <= (inputs(197)) and not (inputs(145));
    layer0_outputs(309) <= '0';
    layer0_outputs(310) <= (inputs(32)) xor (inputs(43));
    layer0_outputs(311) <= not(inputs(93));
    layer0_outputs(312) <= not((inputs(240)) xor (inputs(188)));
    layer0_outputs(313) <= not((inputs(48)) or (inputs(51)));
    layer0_outputs(314) <= (inputs(89)) or (inputs(234));
    layer0_outputs(315) <= not(inputs(132));
    layer0_outputs(316) <= not(inputs(93)) or (inputs(126));
    layer0_outputs(317) <= '0';
    layer0_outputs(318) <= (inputs(4)) and not (inputs(225));
    layer0_outputs(319) <= not((inputs(212)) or (inputs(179)));
    layer0_outputs(320) <= (inputs(82)) or (inputs(37));
    layer0_outputs(321) <= inputs(13);
    layer0_outputs(322) <= not((inputs(241)) and (inputs(32)));
    layer0_outputs(323) <= not(inputs(174));
    layer0_outputs(324) <= not(inputs(176));
    layer0_outputs(325) <= (inputs(120)) and not (inputs(143));
    layer0_outputs(326) <= not(inputs(165));
    layer0_outputs(327) <= not((inputs(43)) xor (inputs(181)));
    layer0_outputs(328) <= not(inputs(92)) or (inputs(45));
    layer0_outputs(329) <= not(inputs(88));
    layer0_outputs(330) <= not((inputs(215)) or (inputs(230)));
    layer0_outputs(331) <= (inputs(13)) or (inputs(159));
    layer0_outputs(332) <= not(inputs(165));
    layer0_outputs(333) <= not(inputs(202));
    layer0_outputs(334) <= not(inputs(232)) or (inputs(16));
    layer0_outputs(335) <= (inputs(66)) and not (inputs(112));
    layer0_outputs(336) <= (inputs(26)) and not (inputs(20));
    layer0_outputs(337) <= not(inputs(201)) or (inputs(220));
    layer0_outputs(338) <= not(inputs(91)) or (inputs(46));
    layer0_outputs(339) <= '0';
    layer0_outputs(340) <= inputs(119);
    layer0_outputs(341) <= not((inputs(64)) xor (inputs(122)));
    layer0_outputs(342) <= not((inputs(38)) and (inputs(111)));
    layer0_outputs(343) <= not((inputs(101)) xor (inputs(163)));
    layer0_outputs(344) <= not(inputs(56));
    layer0_outputs(345) <= inputs(135);
    layer0_outputs(346) <= not(inputs(200));
    layer0_outputs(347) <= not((inputs(84)) and (inputs(191)));
    layer0_outputs(348) <= not((inputs(76)) xor (inputs(105)));
    layer0_outputs(349) <= (inputs(163)) or (inputs(6));
    layer0_outputs(350) <= not((inputs(67)) or (inputs(162)));
    layer0_outputs(351) <= not(inputs(94)) or (inputs(175));
    layer0_outputs(352) <= not((inputs(207)) or (inputs(89)));
    layer0_outputs(353) <= not(inputs(73)) or (inputs(220));
    layer0_outputs(354) <= not((inputs(27)) xor (inputs(71)));
    layer0_outputs(355) <= (inputs(148)) or (inputs(207));
    layer0_outputs(356) <= (inputs(115)) or (inputs(246));
    layer0_outputs(357) <= (inputs(50)) xor (inputs(108));
    layer0_outputs(358) <= inputs(165);
    layer0_outputs(359) <= (inputs(237)) or (inputs(104));
    layer0_outputs(360) <= inputs(147);
    layer0_outputs(361) <= not(inputs(150));
    layer0_outputs(362) <= (inputs(7)) and not (inputs(21));
    layer0_outputs(363) <= not((inputs(248)) or (inputs(200)));
    layer0_outputs(364) <= not(inputs(190));
    layer0_outputs(365) <= not(inputs(167)) or (inputs(253));
    layer0_outputs(366) <= (inputs(85)) and not (inputs(177));
    layer0_outputs(367) <= (inputs(48)) and not (inputs(9));
    layer0_outputs(368) <= not(inputs(177)) or (inputs(236));
    layer0_outputs(369) <= (inputs(58)) or (inputs(66));
    layer0_outputs(370) <= not(inputs(104));
    layer0_outputs(371) <= not(inputs(10)) or (inputs(249));
    layer0_outputs(372) <= not((inputs(39)) xor (inputs(95)));
    layer0_outputs(373) <= not(inputs(255)) or (inputs(112));
    layer0_outputs(374) <= '1';
    layer0_outputs(375) <= not((inputs(183)) or (inputs(9)));
    layer0_outputs(376) <= not((inputs(152)) xor (inputs(141)));
    layer0_outputs(377) <= (inputs(231)) and not (inputs(13));
    layer0_outputs(378) <= inputs(197);
    layer0_outputs(379) <= not((inputs(112)) or (inputs(187)));
    layer0_outputs(380) <= (inputs(27)) xor (inputs(211));
    layer0_outputs(381) <= not((inputs(240)) and (inputs(126)));
    layer0_outputs(382) <= '1';
    layer0_outputs(383) <= (inputs(147)) xor (inputs(174));
    layer0_outputs(384) <= not(inputs(61)) or (inputs(242));
    layer0_outputs(385) <= (inputs(172)) or (inputs(107));
    layer0_outputs(386) <= '1';
    layer0_outputs(387) <= not((inputs(177)) xor (inputs(41)));
    layer0_outputs(388) <= (inputs(94)) or (inputs(55));
    layer0_outputs(389) <= not(inputs(45));
    layer0_outputs(390) <= inputs(99);
    layer0_outputs(391) <= not((inputs(18)) and (inputs(245)));
    layer0_outputs(392) <= (inputs(164)) and not (inputs(242));
    layer0_outputs(393) <= not(inputs(148));
    layer0_outputs(394) <= not((inputs(244)) or (inputs(44)));
    layer0_outputs(395) <= (inputs(153)) xor (inputs(191));
    layer0_outputs(396) <= not(inputs(2));
    layer0_outputs(397) <= inputs(183);
    layer0_outputs(398) <= (inputs(143)) xor (inputs(72));
    layer0_outputs(399) <= not((inputs(226)) or (inputs(50)));
    layer0_outputs(400) <= inputs(94);
    layer0_outputs(401) <= (inputs(240)) or (inputs(152));
    layer0_outputs(402) <= not((inputs(178)) or (inputs(240)));
    layer0_outputs(403) <= (inputs(34)) and (inputs(235));
    layer0_outputs(404) <= not(inputs(215)) or (inputs(94));
    layer0_outputs(405) <= not((inputs(82)) or (inputs(68)));
    layer0_outputs(406) <= not((inputs(67)) xor (inputs(25)));
    layer0_outputs(407) <= inputs(148);
    layer0_outputs(408) <= not((inputs(208)) xor (inputs(165)));
    layer0_outputs(409) <= (inputs(73)) or (inputs(178));
    layer0_outputs(410) <= inputs(180);
    layer0_outputs(411) <= (inputs(118)) xor (inputs(175));
    layer0_outputs(412) <= not((inputs(47)) or (inputs(126)));
    layer0_outputs(413) <= not((inputs(83)) or (inputs(170)));
    layer0_outputs(414) <= (inputs(234)) xor (inputs(100));
    layer0_outputs(415) <= inputs(143);
    layer0_outputs(416) <= (inputs(198)) or (inputs(6));
    layer0_outputs(417) <= (inputs(98)) and not (inputs(216));
    layer0_outputs(418) <= inputs(55);
    layer0_outputs(419) <= not((inputs(250)) or (inputs(177)));
    layer0_outputs(420) <= (inputs(2)) and not (inputs(50));
    layer0_outputs(421) <= (inputs(223)) xor (inputs(59));
    layer0_outputs(422) <= (inputs(152)) and (inputs(201));
    layer0_outputs(423) <= (inputs(190)) or (inputs(39));
    layer0_outputs(424) <= not((inputs(14)) xor (inputs(60)));
    layer0_outputs(425) <= (inputs(116)) or (inputs(153));
    layer0_outputs(426) <= not((inputs(63)) xor (inputs(147)));
    layer0_outputs(427) <= '1';
    layer0_outputs(428) <= inputs(166);
    layer0_outputs(429) <= not(inputs(171)) or (inputs(233));
    layer0_outputs(430) <= '1';
    layer0_outputs(431) <= not(inputs(29));
    layer0_outputs(432) <= not((inputs(186)) xor (inputs(79)));
    layer0_outputs(433) <= inputs(120);
    layer0_outputs(434) <= (inputs(8)) and not (inputs(178));
    layer0_outputs(435) <= '0';
    layer0_outputs(436) <= (inputs(241)) or (inputs(26));
    layer0_outputs(437) <= (inputs(97)) or (inputs(178));
    layer0_outputs(438) <= (inputs(235)) and not (inputs(220));
    layer0_outputs(439) <= inputs(181);
    layer0_outputs(440) <= not((inputs(248)) xor (inputs(182)));
    layer0_outputs(441) <= not(inputs(175)) or (inputs(245));
    layer0_outputs(442) <= (inputs(54)) or (inputs(60));
    layer0_outputs(443) <= (inputs(39)) and (inputs(109));
    layer0_outputs(444) <= not(inputs(106));
    layer0_outputs(445) <= (inputs(85)) or (inputs(111));
    layer0_outputs(446) <= not((inputs(152)) or (inputs(39)));
    layer0_outputs(447) <= '0';
    layer0_outputs(448) <= not(inputs(161)) or (inputs(98));
    layer0_outputs(449) <= (inputs(83)) and (inputs(165));
    layer0_outputs(450) <= not((inputs(121)) and (inputs(57)));
    layer0_outputs(451) <= (inputs(63)) or (inputs(124));
    layer0_outputs(452) <= not(inputs(156)) or (inputs(241));
    layer0_outputs(453) <= (inputs(211)) xor (inputs(114));
    layer0_outputs(454) <= (inputs(64)) and not (inputs(205));
    layer0_outputs(455) <= (inputs(88)) or (inputs(96));
    layer0_outputs(456) <= (inputs(219)) xor (inputs(255));
    layer0_outputs(457) <= inputs(39);
    layer0_outputs(458) <= not(inputs(166));
    layer0_outputs(459) <= '0';
    layer0_outputs(460) <= not((inputs(20)) or (inputs(169)));
    layer0_outputs(461) <= '1';
    layer0_outputs(462) <= (inputs(25)) and not (inputs(29));
    layer0_outputs(463) <= inputs(93);
    layer0_outputs(464) <= (inputs(75)) or (inputs(37));
    layer0_outputs(465) <= (inputs(193)) or (inputs(194));
    layer0_outputs(466) <= (inputs(177)) xor (inputs(112));
    layer0_outputs(467) <= (inputs(58)) xor (inputs(191));
    layer0_outputs(468) <= (inputs(36)) xor (inputs(98));
    layer0_outputs(469) <= inputs(92);
    layer0_outputs(470) <= inputs(236);
    layer0_outputs(471) <= not((inputs(156)) or (inputs(87)));
    layer0_outputs(472) <= not((inputs(184)) xor (inputs(251)));
    layer0_outputs(473) <= (inputs(96)) or (inputs(185));
    layer0_outputs(474) <= not(inputs(75));
    layer0_outputs(475) <= not(inputs(184)) or (inputs(174));
    layer0_outputs(476) <= not(inputs(232));
    layer0_outputs(477) <= not((inputs(55)) or (inputs(255)));
    layer0_outputs(478) <= inputs(161);
    layer0_outputs(479) <= not((inputs(14)) and (inputs(250)));
    layer0_outputs(480) <= not(inputs(132));
    layer0_outputs(481) <= inputs(119);
    layer0_outputs(482) <= '0';
    layer0_outputs(483) <= not(inputs(167));
    layer0_outputs(484) <= not((inputs(8)) or (inputs(213)));
    layer0_outputs(485) <= (inputs(206)) xor (inputs(57));
    layer0_outputs(486) <= not((inputs(6)) xor (inputs(218)));
    layer0_outputs(487) <= not(inputs(80));
    layer0_outputs(488) <= '0';
    layer0_outputs(489) <= not(inputs(86)) or (inputs(197));
    layer0_outputs(490) <= inputs(91);
    layer0_outputs(491) <= (inputs(137)) or (inputs(81));
    layer0_outputs(492) <= (inputs(218)) and not (inputs(126));
    layer0_outputs(493) <= (inputs(218)) xor (inputs(87));
    layer0_outputs(494) <= not(inputs(41));
    layer0_outputs(495) <= not((inputs(220)) and (inputs(5)));
    layer0_outputs(496) <= not(inputs(10));
    layer0_outputs(497) <= not((inputs(35)) or (inputs(54)));
    layer0_outputs(498) <= inputs(31);
    layer0_outputs(499) <= not(inputs(69));
    layer0_outputs(500) <= (inputs(163)) or (inputs(84));
    layer0_outputs(501) <= (inputs(115)) and not (inputs(48));
    layer0_outputs(502) <= '0';
    layer0_outputs(503) <= inputs(109);
    layer0_outputs(504) <= (inputs(53)) or (inputs(228));
    layer0_outputs(505) <= not(inputs(108)) or (inputs(248));
    layer0_outputs(506) <= inputs(101);
    layer0_outputs(507) <= (inputs(17)) xor (inputs(105));
    layer0_outputs(508) <= (inputs(246)) or (inputs(47));
    layer0_outputs(509) <= not(inputs(130));
    layer0_outputs(510) <= inputs(245);
    layer0_outputs(511) <= not(inputs(193));
    layer0_outputs(512) <= (inputs(76)) or (inputs(67));
    layer0_outputs(513) <= not((inputs(84)) or (inputs(126)));
    layer0_outputs(514) <= not((inputs(32)) and (inputs(1)));
    layer0_outputs(515) <= (inputs(132)) or (inputs(167));
    layer0_outputs(516) <= (inputs(133)) and not (inputs(68));
    layer0_outputs(517) <= inputs(179);
    layer0_outputs(518) <= not(inputs(44)) or (inputs(1));
    layer0_outputs(519) <= (inputs(55)) and not (inputs(126));
    layer0_outputs(520) <= not((inputs(182)) or (inputs(36)));
    layer0_outputs(521) <= not(inputs(133));
    layer0_outputs(522) <= (inputs(162)) and (inputs(127));
    layer0_outputs(523) <= not((inputs(63)) or (inputs(117)));
    layer0_outputs(524) <= not((inputs(250)) xor (inputs(133)));
    layer0_outputs(525) <= (inputs(77)) xor (inputs(75));
    layer0_outputs(526) <= (inputs(66)) or (inputs(43));
    layer0_outputs(527) <= inputs(38);
    layer0_outputs(528) <= not(inputs(154)) or (inputs(62));
    layer0_outputs(529) <= not(inputs(41)) or (inputs(205));
    layer0_outputs(530) <= (inputs(100)) and not (inputs(238));
    layer0_outputs(531) <= (inputs(230)) and not (inputs(13));
    layer0_outputs(532) <= (inputs(243)) or (inputs(141));
    layer0_outputs(533) <= (inputs(19)) and (inputs(98));
    layer0_outputs(534) <= (inputs(74)) and not (inputs(201));
    layer0_outputs(535) <= not((inputs(112)) or (inputs(30)));
    layer0_outputs(536) <= inputs(121);
    layer0_outputs(537) <= not(inputs(163));
    layer0_outputs(538) <= not(inputs(234)) or (inputs(172));
    layer0_outputs(539) <= (inputs(73)) and not (inputs(81));
    layer0_outputs(540) <= not(inputs(189));
    layer0_outputs(541) <= not(inputs(44));
    layer0_outputs(542) <= (inputs(167)) and not (inputs(242));
    layer0_outputs(543) <= inputs(137);
    layer0_outputs(544) <= '1';
    layer0_outputs(545) <= not(inputs(180)) or (inputs(21));
    layer0_outputs(546) <= not((inputs(42)) or (inputs(124)));
    layer0_outputs(547) <= inputs(188);
    layer0_outputs(548) <= (inputs(197)) and not (inputs(8));
    layer0_outputs(549) <= (inputs(251)) xor (inputs(12));
    layer0_outputs(550) <= '1';
    layer0_outputs(551) <= (inputs(137)) and not (inputs(217));
    layer0_outputs(552) <= (inputs(231)) xor (inputs(78));
    layer0_outputs(553) <= not(inputs(98)) or (inputs(35));
    layer0_outputs(554) <= inputs(197);
    layer0_outputs(555) <= not(inputs(200));
    layer0_outputs(556) <= not((inputs(191)) xor (inputs(90)));
    layer0_outputs(557) <= (inputs(231)) or (inputs(187));
    layer0_outputs(558) <= not(inputs(117)) or (inputs(67));
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= not((inputs(253)) and (inputs(227)));
    layer0_outputs(561) <= (inputs(179)) or (inputs(144));
    layer0_outputs(562) <= (inputs(10)) xor (inputs(23));
    layer0_outputs(563) <= (inputs(150)) and not (inputs(217));
    layer0_outputs(564) <= '1';
    layer0_outputs(565) <= inputs(116);
    layer0_outputs(566) <= not((inputs(247)) or (inputs(125)));
    layer0_outputs(567) <= (inputs(92)) and not (inputs(247));
    layer0_outputs(568) <= inputs(134);
    layer0_outputs(569) <= (inputs(67)) and not (inputs(168));
    layer0_outputs(570) <= (inputs(233)) xor (inputs(178));
    layer0_outputs(571) <= (inputs(38)) or (inputs(159));
    layer0_outputs(572) <= inputs(153);
    layer0_outputs(573) <= inputs(8);
    layer0_outputs(574) <= (inputs(9)) xor (inputs(243));
    layer0_outputs(575) <= (inputs(225)) xor (inputs(245));
    layer0_outputs(576) <= not(inputs(105));
    layer0_outputs(577) <= not(inputs(35));
    layer0_outputs(578) <= '1';
    layer0_outputs(579) <= (inputs(110)) or (inputs(205));
    layer0_outputs(580) <= inputs(182);
    layer0_outputs(581) <= inputs(247);
    layer0_outputs(582) <= inputs(197);
    layer0_outputs(583) <= not(inputs(120));
    layer0_outputs(584) <= not(inputs(64)) or (inputs(51));
    layer0_outputs(585) <= not(inputs(97));
    layer0_outputs(586) <= (inputs(171)) xor (inputs(57));
    layer0_outputs(587) <= not(inputs(140)) or (inputs(206));
    layer0_outputs(588) <= not(inputs(219));
    layer0_outputs(589) <= not(inputs(17));
    layer0_outputs(590) <= not((inputs(143)) and (inputs(236)));
    layer0_outputs(591) <= (inputs(100)) xor (inputs(5));
    layer0_outputs(592) <= (inputs(64)) and (inputs(97));
    layer0_outputs(593) <= not((inputs(93)) or (inputs(227)));
    layer0_outputs(594) <= not((inputs(117)) or (inputs(229)));
    layer0_outputs(595) <= inputs(5);
    layer0_outputs(596) <= not(inputs(150)) or (inputs(54));
    layer0_outputs(597) <= not((inputs(23)) and (inputs(8)));
    layer0_outputs(598) <= inputs(120);
    layer0_outputs(599) <= not(inputs(39));
    layer0_outputs(600) <= (inputs(201)) xor (inputs(137));
    layer0_outputs(601) <= (inputs(227)) or (inputs(106));
    layer0_outputs(602) <= not((inputs(145)) or (inputs(117)));
    layer0_outputs(603) <= inputs(103);
    layer0_outputs(604) <= (inputs(2)) or (inputs(156));
    layer0_outputs(605) <= inputs(121);
    layer0_outputs(606) <= not((inputs(60)) or (inputs(85)));
    layer0_outputs(607) <= (inputs(151)) and not (inputs(205));
    layer0_outputs(608) <= (inputs(230)) or (inputs(39));
    layer0_outputs(609) <= '1';
    layer0_outputs(610) <= (inputs(16)) xor (inputs(234));
    layer0_outputs(611) <= not(inputs(159)) or (inputs(217));
    layer0_outputs(612) <= '0';
    layer0_outputs(613) <= not((inputs(31)) and (inputs(140)));
    layer0_outputs(614) <= (inputs(145)) and not (inputs(62));
    layer0_outputs(615) <= (inputs(182)) and not (inputs(103));
    layer0_outputs(616) <= (inputs(186)) or (inputs(156));
    layer0_outputs(617) <= not(inputs(151));
    layer0_outputs(618) <= not((inputs(225)) xor (inputs(148)));
    layer0_outputs(619) <= (inputs(29)) or (inputs(213));
    layer0_outputs(620) <= not((inputs(51)) xor (inputs(175)));
    layer0_outputs(621) <= not(inputs(115)) or (inputs(190));
    layer0_outputs(622) <= (inputs(202)) or (inputs(53));
    layer0_outputs(623) <= (inputs(228)) and not (inputs(8));
    layer0_outputs(624) <= not((inputs(97)) and (inputs(126)));
    layer0_outputs(625) <= (inputs(75)) xor (inputs(123));
    layer0_outputs(626) <= (inputs(58)) xor (inputs(93));
    layer0_outputs(627) <= not(inputs(27)) or (inputs(60));
    layer0_outputs(628) <= not((inputs(101)) xor (inputs(175)));
    layer0_outputs(629) <= (inputs(172)) or (inputs(198));
    layer0_outputs(630) <= (inputs(198)) and not (inputs(99));
    layer0_outputs(631) <= '1';
    layer0_outputs(632) <= (inputs(208)) xor (inputs(61));
    layer0_outputs(633) <= (inputs(80)) xor (inputs(186));
    layer0_outputs(634) <= (inputs(193)) and not (inputs(205));
    layer0_outputs(635) <= (inputs(107)) and not (inputs(63));
    layer0_outputs(636) <= not((inputs(150)) or (inputs(64)));
    layer0_outputs(637) <= not((inputs(17)) or (inputs(145)));
    layer0_outputs(638) <= (inputs(121)) and not (inputs(164));
    layer0_outputs(639) <= not((inputs(17)) xor (inputs(210)));
    layer0_outputs(640) <= (inputs(196)) or (inputs(29));
    layer0_outputs(641) <= (inputs(184)) and not (inputs(130));
    layer0_outputs(642) <= not((inputs(139)) or (inputs(14)));
    layer0_outputs(643) <= (inputs(247)) or (inputs(240));
    layer0_outputs(644) <= (inputs(221)) and not (inputs(254));
    layer0_outputs(645) <= not(inputs(183)) or (inputs(10));
    layer0_outputs(646) <= not(inputs(137)) or (inputs(231));
    layer0_outputs(647) <= not((inputs(168)) or (inputs(20)));
    layer0_outputs(648) <= not((inputs(14)) and (inputs(73)));
    layer0_outputs(649) <= (inputs(37)) and not (inputs(53));
    layer0_outputs(650) <= not((inputs(56)) or (inputs(160)));
    layer0_outputs(651) <= (inputs(249)) or (inputs(176));
    layer0_outputs(652) <= not(inputs(149));
    layer0_outputs(653) <= not((inputs(156)) xor (inputs(65)));
    layer0_outputs(654) <= not(inputs(235)) or (inputs(35));
    layer0_outputs(655) <= '0';
    layer0_outputs(656) <= (inputs(151)) or (inputs(158));
    layer0_outputs(657) <= not(inputs(136));
    layer0_outputs(658) <= inputs(167);
    layer0_outputs(659) <= not((inputs(60)) or (inputs(139)));
    layer0_outputs(660) <= (inputs(241)) xor (inputs(118));
    layer0_outputs(661) <= not((inputs(148)) or (inputs(43)));
    layer0_outputs(662) <= not(inputs(231));
    layer0_outputs(663) <= not(inputs(94)) or (inputs(33));
    layer0_outputs(664) <= not(inputs(38));
    layer0_outputs(665) <= not(inputs(173)) or (inputs(146));
    layer0_outputs(666) <= (inputs(100)) or (inputs(206));
    layer0_outputs(667) <= not((inputs(229)) or (inputs(240)));
    layer0_outputs(668) <= (inputs(234)) or (inputs(124));
    layer0_outputs(669) <= not((inputs(22)) xor (inputs(146)));
    layer0_outputs(670) <= (inputs(108)) or (inputs(107));
    layer0_outputs(671) <= inputs(124);
    layer0_outputs(672) <= not((inputs(55)) xor (inputs(238)));
    layer0_outputs(673) <= not(inputs(67));
    layer0_outputs(674) <= (inputs(92)) and not (inputs(235));
    layer0_outputs(675) <= not(inputs(180));
    layer0_outputs(676) <= not((inputs(36)) or (inputs(45)));
    layer0_outputs(677) <= not(inputs(120));
    layer0_outputs(678) <= (inputs(77)) xor (inputs(202));
    layer0_outputs(679) <= not(inputs(216)) or (inputs(143));
    layer0_outputs(680) <= (inputs(254)) xor (inputs(200));
    layer0_outputs(681) <= not((inputs(98)) or (inputs(229)));
    layer0_outputs(682) <= '0';
    layer0_outputs(683) <= (inputs(236)) xor (inputs(66));
    layer0_outputs(684) <= '0';
    layer0_outputs(685) <= not((inputs(69)) or (inputs(213)));
    layer0_outputs(686) <= inputs(144);
    layer0_outputs(687) <= not(inputs(78));
    layer0_outputs(688) <= (inputs(54)) and not (inputs(131));
    layer0_outputs(689) <= not(inputs(128));
    layer0_outputs(690) <= inputs(140);
    layer0_outputs(691) <= not((inputs(23)) or (inputs(148)));
    layer0_outputs(692) <= not(inputs(233)) or (inputs(253));
    layer0_outputs(693) <= (inputs(61)) or (inputs(89));
    layer0_outputs(694) <= not(inputs(43)) or (inputs(162));
    layer0_outputs(695) <= (inputs(44)) and not (inputs(13));
    layer0_outputs(696) <= (inputs(44)) or (inputs(0));
    layer0_outputs(697) <= not((inputs(185)) or (inputs(156)));
    layer0_outputs(698) <= not(inputs(0)) or (inputs(24));
    layer0_outputs(699) <= inputs(32);
    layer0_outputs(700) <= not(inputs(215)) or (inputs(237));
    layer0_outputs(701) <= not(inputs(105));
    layer0_outputs(702) <= inputs(250);
    layer0_outputs(703) <= not(inputs(132));
    layer0_outputs(704) <= not(inputs(91)) or (inputs(219));
    layer0_outputs(705) <= (inputs(252)) or (inputs(166));
    layer0_outputs(706) <= inputs(184);
    layer0_outputs(707) <= not(inputs(97)) or (inputs(25));
    layer0_outputs(708) <= not((inputs(143)) or (inputs(53)));
    layer0_outputs(709) <= not(inputs(93)) or (inputs(1));
    layer0_outputs(710) <= not((inputs(161)) xor (inputs(157)));
    layer0_outputs(711) <= '0';
    layer0_outputs(712) <= inputs(12);
    layer0_outputs(713) <= not(inputs(144)) or (inputs(129));
    layer0_outputs(714) <= (inputs(153)) and not (inputs(163));
    layer0_outputs(715) <= not((inputs(181)) or (inputs(180)));
    layer0_outputs(716) <= (inputs(78)) or (inputs(18));
    layer0_outputs(717) <= (inputs(142)) and not (inputs(184));
    layer0_outputs(718) <= not((inputs(98)) or (inputs(24)));
    layer0_outputs(719) <= not(inputs(119)) or (inputs(32));
    layer0_outputs(720) <= not((inputs(205)) xor (inputs(230)));
    layer0_outputs(721) <= not((inputs(96)) xor (inputs(84)));
    layer0_outputs(722) <= not(inputs(99));
    layer0_outputs(723) <= '0';
    layer0_outputs(724) <= not((inputs(86)) or (inputs(78)));
    layer0_outputs(725) <= inputs(118);
    layer0_outputs(726) <= (inputs(88)) xor (inputs(42));
    layer0_outputs(727) <= not((inputs(0)) or (inputs(75)));
    layer0_outputs(728) <= (inputs(120)) or (inputs(5));
    layer0_outputs(729) <= (inputs(85)) and not (inputs(146));
    layer0_outputs(730) <= inputs(55);
    layer0_outputs(731) <= not((inputs(248)) xor (inputs(167)));
    layer0_outputs(732) <= not(inputs(218));
    layer0_outputs(733) <= not((inputs(17)) and (inputs(186)));
    layer0_outputs(734) <= (inputs(115)) and (inputs(243));
    layer0_outputs(735) <= not((inputs(123)) or (inputs(108)));
    layer0_outputs(736) <= (inputs(134)) and not (inputs(7));
    layer0_outputs(737) <= inputs(133);
    layer0_outputs(738) <= (inputs(0)) xor (inputs(198));
    layer0_outputs(739) <= '1';
    layer0_outputs(740) <= not(inputs(183));
    layer0_outputs(741) <= not(inputs(55));
    layer0_outputs(742) <= inputs(53);
    layer0_outputs(743) <= (inputs(179)) and not (inputs(179));
    layer0_outputs(744) <= not((inputs(20)) and (inputs(226)));
    layer0_outputs(745) <= not(inputs(228));
    layer0_outputs(746) <= not(inputs(149)) or (inputs(8));
    layer0_outputs(747) <= not(inputs(202)) or (inputs(80));
    layer0_outputs(748) <= (inputs(48)) or (inputs(104));
    layer0_outputs(749) <= (inputs(23)) and not (inputs(146));
    layer0_outputs(750) <= '1';
    layer0_outputs(751) <= not(inputs(54));
    layer0_outputs(752) <= not((inputs(11)) and (inputs(127)));
    layer0_outputs(753) <= inputs(89);
    layer0_outputs(754) <= (inputs(203)) xor (inputs(170));
    layer0_outputs(755) <= not((inputs(46)) xor (inputs(191)));
    layer0_outputs(756) <= not((inputs(141)) and (inputs(31)));
    layer0_outputs(757) <= not(inputs(110)) or (inputs(18));
    layer0_outputs(758) <= (inputs(157)) xor (inputs(41));
    layer0_outputs(759) <= not(inputs(87)) or (inputs(226));
    layer0_outputs(760) <= not(inputs(253)) or (inputs(27));
    layer0_outputs(761) <= (inputs(69)) and not (inputs(223));
    layer0_outputs(762) <= (inputs(57)) or (inputs(186));
    layer0_outputs(763) <= not((inputs(77)) or (inputs(14)));
    layer0_outputs(764) <= (inputs(35)) and (inputs(18));
    layer0_outputs(765) <= (inputs(19)) or (inputs(55));
    layer0_outputs(766) <= (inputs(161)) and not (inputs(209));
    layer0_outputs(767) <= not((inputs(1)) xor (inputs(151)));
    layer0_outputs(768) <= not(inputs(122)) or (inputs(18));
    layer0_outputs(769) <= not(inputs(131));
    layer0_outputs(770) <= inputs(14);
    layer0_outputs(771) <= (inputs(191)) or (inputs(99));
    layer0_outputs(772) <= not(inputs(242)) or (inputs(173));
    layer0_outputs(773) <= (inputs(232)) xor (inputs(203));
    layer0_outputs(774) <= (inputs(182)) xor (inputs(15));
    layer0_outputs(775) <= not(inputs(142)) or (inputs(152));
    layer0_outputs(776) <= inputs(160);
    layer0_outputs(777) <= not((inputs(53)) and (inputs(56)));
    layer0_outputs(778) <= inputs(196);
    layer0_outputs(779) <= not((inputs(7)) xor (inputs(240)));
    layer0_outputs(780) <= not(inputs(27));
    layer0_outputs(781) <= (inputs(111)) and (inputs(20));
    layer0_outputs(782) <= not((inputs(45)) xor (inputs(69)));
    layer0_outputs(783) <= (inputs(15)) or (inputs(162));
    layer0_outputs(784) <= (inputs(197)) and not (inputs(234));
    layer0_outputs(785) <= not((inputs(125)) or (inputs(194)));
    layer0_outputs(786) <= not(inputs(33)) or (inputs(127));
    layer0_outputs(787) <= not((inputs(231)) or (inputs(170)));
    layer0_outputs(788) <= not(inputs(225));
    layer0_outputs(789) <= (inputs(215)) and not (inputs(44));
    layer0_outputs(790) <= inputs(206);
    layer0_outputs(791) <= (inputs(228)) and (inputs(224));
    layer0_outputs(792) <= (inputs(231)) or (inputs(63));
    layer0_outputs(793) <= (inputs(246)) and not (inputs(185));
    layer0_outputs(794) <= not(inputs(139)) or (inputs(16));
    layer0_outputs(795) <= (inputs(18)) or (inputs(122));
    layer0_outputs(796) <= (inputs(231)) and not (inputs(219));
    layer0_outputs(797) <= (inputs(238)) and not (inputs(126));
    layer0_outputs(798) <= not((inputs(55)) and (inputs(152)));
    layer0_outputs(799) <= (inputs(174)) or (inputs(211));
    layer0_outputs(800) <= (inputs(214)) or (inputs(108));
    layer0_outputs(801) <= (inputs(202)) or (inputs(38));
    layer0_outputs(802) <= not(inputs(42));
    layer0_outputs(803) <= not((inputs(70)) or (inputs(194)));
    layer0_outputs(804) <= inputs(107);
    layer0_outputs(805) <= inputs(133);
    layer0_outputs(806) <= (inputs(103)) or (inputs(161));
    layer0_outputs(807) <= not(inputs(38));
    layer0_outputs(808) <= (inputs(140)) or (inputs(61));
    layer0_outputs(809) <= not(inputs(216)) or (inputs(109));
    layer0_outputs(810) <= inputs(73);
    layer0_outputs(811) <= (inputs(51)) and not (inputs(191));
    layer0_outputs(812) <= inputs(223);
    layer0_outputs(813) <= (inputs(101)) xor (inputs(9));
    layer0_outputs(814) <= not((inputs(119)) xor (inputs(204)));
    layer0_outputs(815) <= (inputs(158)) or (inputs(167));
    layer0_outputs(816) <= not((inputs(164)) or (inputs(207)));
    layer0_outputs(817) <= (inputs(253)) xor (inputs(38));
    layer0_outputs(818) <= not((inputs(248)) or (inputs(70)));
    layer0_outputs(819) <= (inputs(171)) xor (inputs(196));
    layer0_outputs(820) <= inputs(131);
    layer0_outputs(821) <= (inputs(178)) xor (inputs(251));
    layer0_outputs(822) <= not(inputs(131)) or (inputs(23));
    layer0_outputs(823) <= '0';
    layer0_outputs(824) <= inputs(65);
    layer0_outputs(825) <= not((inputs(39)) or (inputs(11)));
    layer0_outputs(826) <= (inputs(205)) or (inputs(233));
    layer0_outputs(827) <= (inputs(120)) and not (inputs(84));
    layer0_outputs(828) <= inputs(243);
    layer0_outputs(829) <= not((inputs(81)) and (inputs(119)));
    layer0_outputs(830) <= (inputs(3)) and not (inputs(146));
    layer0_outputs(831) <= (inputs(30)) xor (inputs(78));
    layer0_outputs(832) <= not((inputs(4)) xor (inputs(198)));
    layer0_outputs(833) <= not(inputs(115)) or (inputs(57));
    layer0_outputs(834) <= (inputs(31)) xor (inputs(177));
    layer0_outputs(835) <= (inputs(177)) and not (inputs(64));
    layer0_outputs(836) <= (inputs(202)) and not (inputs(28));
    layer0_outputs(837) <= (inputs(147)) and not (inputs(19));
    layer0_outputs(838) <= not((inputs(199)) or (inputs(241)));
    layer0_outputs(839) <= (inputs(173)) or (inputs(5));
    layer0_outputs(840) <= not((inputs(176)) or (inputs(209)));
    layer0_outputs(841) <= inputs(178);
    layer0_outputs(842) <= inputs(156);
    layer0_outputs(843) <= not(inputs(163));
    layer0_outputs(844) <= not((inputs(242)) and (inputs(251)));
    layer0_outputs(845) <= not((inputs(216)) or (inputs(246)));
    layer0_outputs(846) <= not(inputs(174)) or (inputs(117));
    layer0_outputs(847) <= not(inputs(43)) or (inputs(12));
    layer0_outputs(848) <= not((inputs(192)) or (inputs(18)));
    layer0_outputs(849) <= (inputs(190)) xor (inputs(90));
    layer0_outputs(850) <= inputs(92);
    layer0_outputs(851) <= not((inputs(9)) or (inputs(155)));
    layer0_outputs(852) <= not(inputs(240)) or (inputs(12));
    layer0_outputs(853) <= not(inputs(167));
    layer0_outputs(854) <= not(inputs(36)) or (inputs(19));
    layer0_outputs(855) <= (inputs(132)) and not (inputs(95));
    layer0_outputs(856) <= not(inputs(199)) or (inputs(156));
    layer0_outputs(857) <= (inputs(74)) or (inputs(246));
    layer0_outputs(858) <= (inputs(188)) xor (inputs(90));
    layer0_outputs(859) <= (inputs(182)) and not (inputs(114));
    layer0_outputs(860) <= (inputs(220)) or (inputs(193));
    layer0_outputs(861) <= not(inputs(246)) or (inputs(64));
    layer0_outputs(862) <= (inputs(7)) or (inputs(254));
    layer0_outputs(863) <= not((inputs(40)) xor (inputs(196)));
    layer0_outputs(864) <= not(inputs(169)) or (inputs(220));
    layer0_outputs(865) <= not(inputs(72));
    layer0_outputs(866) <= inputs(86);
    layer0_outputs(867) <= not(inputs(212)) or (inputs(82));
    layer0_outputs(868) <= not(inputs(114)) or (inputs(241));
    layer0_outputs(869) <= inputs(114);
    layer0_outputs(870) <= not(inputs(83));
    layer0_outputs(871) <= '1';
    layer0_outputs(872) <= (inputs(180)) or (inputs(210));
    layer0_outputs(873) <= not(inputs(28));
    layer0_outputs(874) <= not(inputs(215));
    layer0_outputs(875) <= (inputs(44)) xor (inputs(15));
    layer0_outputs(876) <= not((inputs(253)) or (inputs(166)));
    layer0_outputs(877) <= (inputs(55)) or (inputs(159));
    layer0_outputs(878) <= (inputs(250)) and (inputs(163));
    layer0_outputs(879) <= not(inputs(182));
    layer0_outputs(880) <= not(inputs(107));
    layer0_outputs(881) <= inputs(23);
    layer0_outputs(882) <= not(inputs(243));
    layer0_outputs(883) <= (inputs(77)) and not (inputs(40));
    layer0_outputs(884) <= not((inputs(114)) xor (inputs(67)));
    layer0_outputs(885) <= (inputs(50)) xor (inputs(41));
    layer0_outputs(886) <= (inputs(109)) or (inputs(25));
    layer0_outputs(887) <= inputs(124);
    layer0_outputs(888) <= not(inputs(253));
    layer0_outputs(889) <= (inputs(94)) xor (inputs(106));
    layer0_outputs(890) <= (inputs(175)) or (inputs(198));
    layer0_outputs(891) <= not(inputs(101));
    layer0_outputs(892) <= (inputs(228)) and not (inputs(174));
    layer0_outputs(893) <= (inputs(162)) and not (inputs(144));
    layer0_outputs(894) <= (inputs(41)) xor (inputs(187));
    layer0_outputs(895) <= not((inputs(185)) xor (inputs(235)));
    layer0_outputs(896) <= not(inputs(103));
    layer0_outputs(897) <= inputs(116);
    layer0_outputs(898) <= (inputs(237)) or (inputs(192));
    layer0_outputs(899) <= (inputs(90)) and (inputs(0));
    layer0_outputs(900) <= (inputs(148)) or (inputs(51));
    layer0_outputs(901) <= (inputs(153)) and not (inputs(179));
    layer0_outputs(902) <= not(inputs(86));
    layer0_outputs(903) <= not(inputs(61));
    layer0_outputs(904) <= not((inputs(129)) or (inputs(165)));
    layer0_outputs(905) <= not((inputs(242)) xor (inputs(38)));
    layer0_outputs(906) <= not((inputs(206)) xor (inputs(8)));
    layer0_outputs(907) <= not(inputs(93)) or (inputs(15));
    layer0_outputs(908) <= (inputs(210)) and not (inputs(9));
    layer0_outputs(909) <= (inputs(122)) or (inputs(255));
    layer0_outputs(910) <= not(inputs(4)) or (inputs(253));
    layer0_outputs(911) <= not(inputs(159));
    layer0_outputs(912) <= (inputs(71)) xor (inputs(91));
    layer0_outputs(913) <= not(inputs(18)) or (inputs(191));
    layer0_outputs(914) <= inputs(121);
    layer0_outputs(915) <= not(inputs(70));
    layer0_outputs(916) <= '0';
    layer0_outputs(917) <= not((inputs(214)) xor (inputs(215)));
    layer0_outputs(918) <= inputs(100);
    layer0_outputs(919) <= '1';
    layer0_outputs(920) <= (inputs(244)) or (inputs(195));
    layer0_outputs(921) <= (inputs(197)) and not (inputs(24));
    layer0_outputs(922) <= '0';
    layer0_outputs(923) <= not((inputs(225)) or (inputs(83)));
    layer0_outputs(924) <= not(inputs(169)) or (inputs(160));
    layer0_outputs(925) <= (inputs(45)) xor (inputs(95));
    layer0_outputs(926) <= (inputs(231)) or (inputs(246));
    layer0_outputs(927) <= not(inputs(64));
    layer0_outputs(928) <= not(inputs(139));
    layer0_outputs(929) <= (inputs(249)) or (inputs(144));
    layer0_outputs(930) <= not(inputs(185));
    layer0_outputs(931) <= (inputs(80)) and not (inputs(1));
    layer0_outputs(932) <= not(inputs(204)) or (inputs(109));
    layer0_outputs(933) <= not(inputs(124));
    layer0_outputs(934) <= not((inputs(24)) and (inputs(36)));
    layer0_outputs(935) <= (inputs(101)) xor (inputs(222));
    layer0_outputs(936) <= '1';
    layer0_outputs(937) <= not((inputs(151)) xor (inputs(246)));
    layer0_outputs(938) <= not((inputs(196)) or (inputs(9)));
    layer0_outputs(939) <= (inputs(238)) xor (inputs(7));
    layer0_outputs(940) <= (inputs(250)) xor (inputs(64));
    layer0_outputs(941) <= not(inputs(216));
    layer0_outputs(942) <= (inputs(153)) or (inputs(147));
    layer0_outputs(943) <= '1';
    layer0_outputs(944) <= not((inputs(64)) or (inputs(218)));
    layer0_outputs(945) <= (inputs(227)) or (inputs(74));
    layer0_outputs(946) <= not((inputs(45)) xor (inputs(159)));
    layer0_outputs(947) <= not((inputs(158)) xor (inputs(51)));
    layer0_outputs(948) <= (inputs(1)) xor (inputs(169));
    layer0_outputs(949) <= (inputs(122)) and not (inputs(214));
    layer0_outputs(950) <= (inputs(216)) and not (inputs(194));
    layer0_outputs(951) <= not((inputs(151)) xor (inputs(29)));
    layer0_outputs(952) <= (inputs(41)) or (inputs(6));
    layer0_outputs(953) <= not((inputs(65)) or (inputs(159)));
    layer0_outputs(954) <= not((inputs(168)) xor (inputs(207)));
    layer0_outputs(955) <= (inputs(184)) xor (inputs(129));
    layer0_outputs(956) <= not((inputs(142)) or (inputs(141)));
    layer0_outputs(957) <= (inputs(70)) and not (inputs(174));
    layer0_outputs(958) <= (inputs(105)) or (inputs(83));
    layer0_outputs(959) <= not(inputs(202));
    layer0_outputs(960) <= not(inputs(32));
    layer0_outputs(961) <= (inputs(197)) or (inputs(78));
    layer0_outputs(962) <= inputs(77);
    layer0_outputs(963) <= not(inputs(61));
    layer0_outputs(964) <= (inputs(202)) or (inputs(145));
    layer0_outputs(965) <= inputs(143);
    layer0_outputs(966) <= not(inputs(132)) or (inputs(48));
    layer0_outputs(967) <= (inputs(55)) or (inputs(195));
    layer0_outputs(968) <= not((inputs(27)) or (inputs(187)));
    layer0_outputs(969) <= inputs(65);
    layer0_outputs(970) <= not((inputs(89)) or (inputs(127)));
    layer0_outputs(971) <= not((inputs(56)) xor (inputs(78)));
    layer0_outputs(972) <= not((inputs(152)) or (inputs(44)));
    layer0_outputs(973) <= not(inputs(103));
    layer0_outputs(974) <= (inputs(214)) and not (inputs(159));
    layer0_outputs(975) <= (inputs(186)) and not (inputs(192));
    layer0_outputs(976) <= not((inputs(59)) or (inputs(248)));
    layer0_outputs(977) <= not(inputs(187));
    layer0_outputs(978) <= not(inputs(18));
    layer0_outputs(979) <= not(inputs(170)) or (inputs(86));
    layer0_outputs(980) <= (inputs(103)) and not (inputs(8));
    layer0_outputs(981) <= (inputs(207)) and not (inputs(33));
    layer0_outputs(982) <= (inputs(185)) and not (inputs(142));
    layer0_outputs(983) <= (inputs(202)) and not (inputs(114));
    layer0_outputs(984) <= not((inputs(26)) or (inputs(149)));
    layer0_outputs(985) <= not((inputs(247)) or (inputs(4)));
    layer0_outputs(986) <= inputs(122);
    layer0_outputs(987) <= (inputs(165)) or (inputs(82));
    layer0_outputs(988) <= '0';
    layer0_outputs(989) <= (inputs(65)) xor (inputs(180));
    layer0_outputs(990) <= (inputs(247)) xor (inputs(164));
    layer0_outputs(991) <= not((inputs(122)) or (inputs(230)));
    layer0_outputs(992) <= not((inputs(140)) or (inputs(15)));
    layer0_outputs(993) <= not(inputs(119));
    layer0_outputs(994) <= not(inputs(86)) or (inputs(139));
    layer0_outputs(995) <= (inputs(71)) and not (inputs(112));
    layer0_outputs(996) <= '0';
    layer0_outputs(997) <= (inputs(165)) or (inputs(175));
    layer0_outputs(998) <= (inputs(125)) or (inputs(187));
    layer0_outputs(999) <= (inputs(91)) xor (inputs(22));
    layer0_outputs(1000) <= (inputs(144)) and not (inputs(31));
    layer0_outputs(1001) <= inputs(47);
    layer0_outputs(1002) <= (inputs(71)) and not (inputs(68));
    layer0_outputs(1003) <= not(inputs(133));
    layer0_outputs(1004) <= not(inputs(32));
    layer0_outputs(1005) <= not(inputs(130));
    layer0_outputs(1006) <= not((inputs(250)) xor (inputs(44)));
    layer0_outputs(1007) <= '1';
    layer0_outputs(1008) <= not(inputs(121));
    layer0_outputs(1009) <= not((inputs(162)) xor (inputs(179)));
    layer0_outputs(1010) <= not(inputs(59)) or (inputs(225));
    layer0_outputs(1011) <= (inputs(158)) and not (inputs(0));
    layer0_outputs(1012) <= (inputs(210)) or (inputs(60));
    layer0_outputs(1013) <= (inputs(154)) or (inputs(27));
    layer0_outputs(1014) <= (inputs(116)) and not (inputs(232));
    layer0_outputs(1015) <= not((inputs(110)) or (inputs(44)));
    layer0_outputs(1016) <= '1';
    layer0_outputs(1017) <= (inputs(75)) and (inputs(18));
    layer0_outputs(1018) <= not((inputs(25)) xor (inputs(68)));
    layer0_outputs(1019) <= not((inputs(136)) or (inputs(109)));
    layer0_outputs(1020) <= inputs(106);
    layer0_outputs(1021) <= not(inputs(117)) or (inputs(205));
    layer0_outputs(1022) <= (inputs(56)) and not (inputs(123));
    layer0_outputs(1023) <= not(inputs(214));
    layer0_outputs(1024) <= not((inputs(118)) or (inputs(63)));
    layer0_outputs(1025) <= not(inputs(229));
    layer0_outputs(1026) <= not(inputs(171)) or (inputs(195));
    layer0_outputs(1027) <= not(inputs(166)) or (inputs(218));
    layer0_outputs(1028) <= not(inputs(27)) or (inputs(237));
    layer0_outputs(1029) <= not(inputs(172));
    layer0_outputs(1030) <= (inputs(115)) and (inputs(160));
    layer0_outputs(1031) <= (inputs(17)) and not (inputs(37));
    layer0_outputs(1032) <= not((inputs(59)) xor (inputs(183)));
    layer0_outputs(1033) <= inputs(164);
    layer0_outputs(1034) <= not(inputs(12)) or (inputs(29));
    layer0_outputs(1035) <= inputs(171);
    layer0_outputs(1036) <= '1';
    layer0_outputs(1037) <= not(inputs(101)) or (inputs(177));
    layer0_outputs(1038) <= not(inputs(17));
    layer0_outputs(1039) <= not((inputs(199)) or (inputs(140)));
    layer0_outputs(1040) <= not((inputs(70)) xor (inputs(105)));
    layer0_outputs(1041) <= (inputs(41)) or (inputs(61));
    layer0_outputs(1042) <= (inputs(61)) or (inputs(138));
    layer0_outputs(1043) <= not((inputs(222)) xor (inputs(39)));
    layer0_outputs(1044) <= not(inputs(40)) or (inputs(246));
    layer0_outputs(1045) <= not((inputs(66)) and (inputs(88)));
    layer0_outputs(1046) <= not(inputs(71));
    layer0_outputs(1047) <= inputs(166);
    layer0_outputs(1048) <= inputs(38);
    layer0_outputs(1049) <= (inputs(180)) or (inputs(7));
    layer0_outputs(1050) <= inputs(39);
    layer0_outputs(1051) <= not(inputs(209)) or (inputs(180));
    layer0_outputs(1052) <= inputs(121);
    layer0_outputs(1053) <= not(inputs(175)) or (inputs(175));
    layer0_outputs(1054) <= not((inputs(143)) or (inputs(48)));
    layer0_outputs(1055) <= (inputs(188)) and (inputs(22));
    layer0_outputs(1056) <= not(inputs(109)) or (inputs(244));
    layer0_outputs(1057) <= not((inputs(9)) or (inputs(33)));
    layer0_outputs(1058) <= not(inputs(41));
    layer0_outputs(1059) <= (inputs(35)) xor (inputs(179));
    layer0_outputs(1060) <= (inputs(245)) and (inputs(152));
    layer0_outputs(1061) <= '1';
    layer0_outputs(1062) <= inputs(101);
    layer0_outputs(1063) <= not(inputs(100));
    layer0_outputs(1064) <= not(inputs(118)) or (inputs(228));
    layer0_outputs(1065) <= not((inputs(222)) xor (inputs(134)));
    layer0_outputs(1066) <= (inputs(169)) and not (inputs(109));
    layer0_outputs(1067) <= (inputs(75)) xor (inputs(106));
    layer0_outputs(1068) <= not(inputs(22));
    layer0_outputs(1069) <= (inputs(196)) and not (inputs(115));
    layer0_outputs(1070) <= (inputs(3)) or (inputs(251));
    layer0_outputs(1071) <= inputs(33);
    layer0_outputs(1072) <= (inputs(215)) or (inputs(140));
    layer0_outputs(1073) <= (inputs(137)) and not (inputs(207));
    layer0_outputs(1074) <= (inputs(8)) and (inputs(30));
    layer0_outputs(1075) <= not(inputs(143)) or (inputs(155));
    layer0_outputs(1076) <= (inputs(123)) or (inputs(124));
    layer0_outputs(1077) <= not((inputs(23)) or (inputs(121)));
    layer0_outputs(1078) <= not(inputs(76));
    layer0_outputs(1079) <= not((inputs(104)) xor (inputs(73)));
    layer0_outputs(1080) <= not(inputs(119));
    layer0_outputs(1081) <= (inputs(113)) or (inputs(252));
    layer0_outputs(1082) <= (inputs(222)) and not (inputs(225));
    layer0_outputs(1083) <= not(inputs(193));
    layer0_outputs(1084) <= (inputs(74)) or (inputs(105));
    layer0_outputs(1085) <= '0';
    layer0_outputs(1086) <= (inputs(147)) xor (inputs(145));
    layer0_outputs(1087) <= not(inputs(182)) or (inputs(116));
    layer0_outputs(1088) <= not((inputs(37)) or (inputs(1)));
    layer0_outputs(1089) <= (inputs(235)) or (inputs(159));
    layer0_outputs(1090) <= inputs(123);
    layer0_outputs(1091) <= (inputs(216)) xor (inputs(192));
    layer0_outputs(1092) <= '1';
    layer0_outputs(1093) <= not((inputs(116)) or (inputs(101)));
    layer0_outputs(1094) <= (inputs(19)) xor (inputs(252));
    layer0_outputs(1095) <= not((inputs(125)) or (inputs(244)));
    layer0_outputs(1096) <= not((inputs(16)) xor (inputs(245)));
    layer0_outputs(1097) <= (inputs(108)) or (inputs(135));
    layer0_outputs(1098) <= not((inputs(89)) or (inputs(120)));
    layer0_outputs(1099) <= not(inputs(72));
    layer0_outputs(1100) <= not(inputs(42));
    layer0_outputs(1101) <= not(inputs(227));
    layer0_outputs(1102) <= not(inputs(201));
    layer0_outputs(1103) <= (inputs(233)) or (inputs(201));
    layer0_outputs(1104) <= not(inputs(250)) or (inputs(156));
    layer0_outputs(1105) <= inputs(155);
    layer0_outputs(1106) <= (inputs(166)) and not (inputs(142));
    layer0_outputs(1107) <= not((inputs(136)) or (inputs(194)));
    layer0_outputs(1108) <= (inputs(65)) xor (inputs(111));
    layer0_outputs(1109) <= not(inputs(130));
    layer0_outputs(1110) <= (inputs(82)) or (inputs(144));
    layer0_outputs(1111) <= not(inputs(201)) or (inputs(9));
    layer0_outputs(1112) <= inputs(86);
    layer0_outputs(1113) <= inputs(207);
    layer0_outputs(1114) <= inputs(208);
    layer0_outputs(1115) <= inputs(247);
    layer0_outputs(1116) <= not(inputs(135));
    layer0_outputs(1117) <= inputs(153);
    layer0_outputs(1118) <= not((inputs(86)) xor (inputs(129)));
    layer0_outputs(1119) <= (inputs(56)) and not (inputs(93));
    layer0_outputs(1120) <= not(inputs(46));
    layer0_outputs(1121) <= inputs(89);
    layer0_outputs(1122) <= (inputs(222)) or (inputs(28));
    layer0_outputs(1123) <= not((inputs(87)) or (inputs(16)));
    layer0_outputs(1124) <= not(inputs(192));
    layer0_outputs(1125) <= inputs(231);
    layer0_outputs(1126) <= not((inputs(65)) or (inputs(144)));
    layer0_outputs(1127) <= not((inputs(154)) xor (inputs(108)));
    layer0_outputs(1128) <= (inputs(149)) and not (inputs(45));
    layer0_outputs(1129) <= (inputs(27)) and not (inputs(97));
    layer0_outputs(1130) <= (inputs(53)) or (inputs(124));
    layer0_outputs(1131) <= inputs(90);
    layer0_outputs(1132) <= not((inputs(163)) and (inputs(163)));
    layer0_outputs(1133) <= not((inputs(53)) xor (inputs(21)));
    layer0_outputs(1134) <= (inputs(57)) or (inputs(109));
    layer0_outputs(1135) <= not(inputs(156)) or (inputs(223));
    layer0_outputs(1136) <= (inputs(20)) or (inputs(223));
    layer0_outputs(1137) <= not(inputs(75));
    layer0_outputs(1138) <= not(inputs(133)) or (inputs(159));
    layer0_outputs(1139) <= (inputs(115)) and not (inputs(77));
    layer0_outputs(1140) <= not((inputs(118)) xor (inputs(241)));
    layer0_outputs(1141) <= not(inputs(31)) or (inputs(22));
    layer0_outputs(1142) <= (inputs(185)) and not (inputs(81));
    layer0_outputs(1143) <= '0';
    layer0_outputs(1144) <= (inputs(27)) or (inputs(103));
    layer0_outputs(1145) <= (inputs(41)) and not (inputs(125));
    layer0_outputs(1146) <= not(inputs(204)) or (inputs(212));
    layer0_outputs(1147) <= (inputs(32)) xor (inputs(44));
    layer0_outputs(1148) <= not(inputs(173));
    layer0_outputs(1149) <= not(inputs(116));
    layer0_outputs(1150) <= not(inputs(175));
    layer0_outputs(1151) <= not(inputs(37));
    layer0_outputs(1152) <= (inputs(149)) or (inputs(28));
    layer0_outputs(1153) <= not((inputs(188)) or (inputs(254)));
    layer0_outputs(1154) <= (inputs(30)) or (inputs(192));
    layer0_outputs(1155) <= (inputs(223)) and (inputs(249));
    layer0_outputs(1156) <= inputs(13);
    layer0_outputs(1157) <= (inputs(54)) and not (inputs(205));
    layer0_outputs(1158) <= inputs(175);
    layer0_outputs(1159) <= (inputs(149)) and not (inputs(177));
    layer0_outputs(1160) <= not((inputs(72)) and (inputs(238)));
    layer0_outputs(1161) <= (inputs(184)) and not (inputs(113));
    layer0_outputs(1162) <= inputs(108);
    layer0_outputs(1163) <= not(inputs(25)) or (inputs(50));
    layer0_outputs(1164) <= (inputs(128)) xor (inputs(219));
    layer0_outputs(1165) <= not(inputs(244)) or (inputs(222));
    layer0_outputs(1166) <= not((inputs(117)) or (inputs(118)));
    layer0_outputs(1167) <= not((inputs(65)) xor (inputs(172)));
    layer0_outputs(1168) <= (inputs(125)) and not (inputs(8));
    layer0_outputs(1169) <= not((inputs(61)) xor (inputs(205)));
    layer0_outputs(1170) <= not((inputs(224)) and (inputs(225)));
    layer0_outputs(1171) <= not((inputs(10)) xor (inputs(84)));
    layer0_outputs(1172) <= inputs(152);
    layer0_outputs(1173) <= inputs(118);
    layer0_outputs(1174) <= (inputs(167)) or (inputs(98));
    layer0_outputs(1175) <= not((inputs(159)) xor (inputs(130)));
    layer0_outputs(1176) <= not((inputs(58)) or (inputs(3)));
    layer0_outputs(1177) <= '1';
    layer0_outputs(1178) <= not((inputs(25)) xor (inputs(8)));
    layer0_outputs(1179) <= not((inputs(108)) or (inputs(130)));
    layer0_outputs(1180) <= not((inputs(207)) and (inputs(63)));
    layer0_outputs(1181) <= not((inputs(94)) or (inputs(59)));
    layer0_outputs(1182) <= (inputs(101)) or (inputs(69));
    layer0_outputs(1183) <= (inputs(99)) and (inputs(82));
    layer0_outputs(1184) <= not(inputs(87)) or (inputs(126));
    layer0_outputs(1185) <= not((inputs(220)) or (inputs(151)));
    layer0_outputs(1186) <= not((inputs(76)) or (inputs(183)));
    layer0_outputs(1187) <= inputs(171);
    layer0_outputs(1188) <= (inputs(53)) or (inputs(62));
    layer0_outputs(1189) <= not(inputs(90));
    layer0_outputs(1190) <= (inputs(131)) or (inputs(117));
    layer0_outputs(1191) <= (inputs(103)) and not (inputs(35));
    layer0_outputs(1192) <= not((inputs(88)) or (inputs(57)));
    layer0_outputs(1193) <= (inputs(38)) and not (inputs(38));
    layer0_outputs(1194) <= not(inputs(216));
    layer0_outputs(1195) <= not((inputs(28)) xor (inputs(192)));
    layer0_outputs(1196) <= inputs(198);
    layer0_outputs(1197) <= (inputs(214)) and not (inputs(68));
    layer0_outputs(1198) <= not(inputs(60));
    layer0_outputs(1199) <= '1';
    layer0_outputs(1200) <= (inputs(117)) and not (inputs(83));
    layer0_outputs(1201) <= not(inputs(27)) or (inputs(242));
    layer0_outputs(1202) <= not((inputs(250)) xor (inputs(138)));
    layer0_outputs(1203) <= inputs(55);
    layer0_outputs(1204) <= (inputs(117)) xor (inputs(79));
    layer0_outputs(1205) <= inputs(82);
    layer0_outputs(1206) <= (inputs(14)) or (inputs(200));
    layer0_outputs(1207) <= (inputs(213)) and not (inputs(221));
    layer0_outputs(1208) <= not(inputs(179)) or (inputs(80));
    layer0_outputs(1209) <= inputs(102);
    layer0_outputs(1210) <= not(inputs(140)) or (inputs(190));
    layer0_outputs(1211) <= not((inputs(190)) xor (inputs(229)));
    layer0_outputs(1212) <= inputs(219);
    layer0_outputs(1213) <= (inputs(211)) and not (inputs(63));
    layer0_outputs(1214) <= not(inputs(31)) or (inputs(127));
    layer0_outputs(1215) <= inputs(68);
    layer0_outputs(1216) <= inputs(186);
    layer0_outputs(1217) <= not(inputs(199));
    layer0_outputs(1218) <= inputs(108);
    layer0_outputs(1219) <= not(inputs(150));
    layer0_outputs(1220) <= not(inputs(194)) or (inputs(49));
    layer0_outputs(1221) <= not(inputs(97)) or (inputs(32));
    layer0_outputs(1222) <= (inputs(81)) and (inputs(248));
    layer0_outputs(1223) <= not((inputs(42)) or (inputs(25)));
    layer0_outputs(1224) <= (inputs(119)) xor (inputs(14));
    layer0_outputs(1225) <= not(inputs(163)) or (inputs(99));
    layer0_outputs(1226) <= not((inputs(93)) xor (inputs(169)));
    layer0_outputs(1227) <= not((inputs(137)) xor (inputs(112)));
    layer0_outputs(1228) <= inputs(122);
    layer0_outputs(1229) <= not((inputs(87)) or (inputs(115)));
    layer0_outputs(1230) <= not(inputs(226));
    layer0_outputs(1231) <= not((inputs(75)) xor (inputs(37)));
    layer0_outputs(1232) <= '1';
    layer0_outputs(1233) <= not(inputs(73));
    layer0_outputs(1234) <= not(inputs(138)) or (inputs(77));
    layer0_outputs(1235) <= not(inputs(92));
    layer0_outputs(1236) <= not((inputs(223)) or (inputs(163)));
    layer0_outputs(1237) <= not(inputs(195)) or (inputs(141));
    layer0_outputs(1238) <= inputs(161);
    layer0_outputs(1239) <= (inputs(174)) or (inputs(29));
    layer0_outputs(1240) <= not((inputs(108)) xor (inputs(152)));
    layer0_outputs(1241) <= inputs(233);
    layer0_outputs(1242) <= inputs(110);
    layer0_outputs(1243) <= not((inputs(220)) or (inputs(37)));
    layer0_outputs(1244) <= not(inputs(242)) or (inputs(65));
    layer0_outputs(1245) <= not(inputs(240));
    layer0_outputs(1246) <= (inputs(210)) and not (inputs(198));
    layer0_outputs(1247) <= inputs(81);
    layer0_outputs(1248) <= (inputs(236)) and not (inputs(21));
    layer0_outputs(1249) <= (inputs(16)) xor (inputs(140));
    layer0_outputs(1250) <= (inputs(165)) xor (inputs(206));
    layer0_outputs(1251) <= not(inputs(147));
    layer0_outputs(1252) <= (inputs(39)) and not (inputs(31));
    layer0_outputs(1253) <= not(inputs(120));
    layer0_outputs(1254) <= (inputs(161)) xor (inputs(172));
    layer0_outputs(1255) <= not(inputs(21));
    layer0_outputs(1256) <= not((inputs(33)) or (inputs(69)));
    layer0_outputs(1257) <= inputs(248);
    layer0_outputs(1258) <= not(inputs(216));
    layer0_outputs(1259) <= not(inputs(151));
    layer0_outputs(1260) <= not((inputs(12)) xor (inputs(56)));
    layer0_outputs(1261) <= not(inputs(69)) or (inputs(251));
    layer0_outputs(1262) <= (inputs(1)) xor (inputs(224));
    layer0_outputs(1263) <= inputs(164);
    layer0_outputs(1264) <= inputs(200);
    layer0_outputs(1265) <= not(inputs(96)) or (inputs(239));
    layer0_outputs(1266) <= (inputs(136)) and not (inputs(172));
    layer0_outputs(1267) <= (inputs(80)) or (inputs(192));
    layer0_outputs(1268) <= (inputs(184)) or (inputs(36));
    layer0_outputs(1269) <= (inputs(3)) xor (inputs(42));
    layer0_outputs(1270) <= (inputs(178)) or (inputs(155));
    layer0_outputs(1271) <= not((inputs(91)) xor (inputs(89)));
    layer0_outputs(1272) <= not(inputs(168)) or (inputs(252));
    layer0_outputs(1273) <= not((inputs(114)) xor (inputs(200)));
    layer0_outputs(1274) <= not(inputs(147));
    layer0_outputs(1275) <= not((inputs(123)) xor (inputs(172)));
    layer0_outputs(1276) <= not((inputs(81)) xor (inputs(167)));
    layer0_outputs(1277) <= (inputs(62)) xor (inputs(105));
    layer0_outputs(1278) <= (inputs(248)) or (inputs(57));
    layer0_outputs(1279) <= (inputs(177)) and (inputs(143));
    layer0_outputs(1280) <= not((inputs(207)) xor (inputs(39)));
    layer0_outputs(1281) <= not((inputs(203)) xor (inputs(94)));
    layer0_outputs(1282) <= not((inputs(240)) xor (inputs(134)));
    layer0_outputs(1283) <= (inputs(50)) xor (inputs(5));
    layer0_outputs(1284) <= not(inputs(45)) or (inputs(19));
    layer0_outputs(1285) <= (inputs(40)) or (inputs(22));
    layer0_outputs(1286) <= not(inputs(167)) or (inputs(35));
    layer0_outputs(1287) <= not(inputs(4)) or (inputs(76));
    layer0_outputs(1288) <= (inputs(121)) or (inputs(205));
    layer0_outputs(1289) <= not(inputs(153)) or (inputs(11));
    layer0_outputs(1290) <= not(inputs(103));
    layer0_outputs(1291) <= not(inputs(36)) or (inputs(111));
    layer0_outputs(1292) <= not(inputs(29));
    layer0_outputs(1293) <= (inputs(87)) or (inputs(234));
    layer0_outputs(1294) <= not((inputs(96)) xor (inputs(251)));
    layer0_outputs(1295) <= not((inputs(178)) or (inputs(228)));
    layer0_outputs(1296) <= (inputs(163)) and (inputs(222));
    layer0_outputs(1297) <= inputs(141);
    layer0_outputs(1298) <= inputs(178);
    layer0_outputs(1299) <= (inputs(186)) xor (inputs(144));
    layer0_outputs(1300) <= (inputs(84)) or (inputs(94));
    layer0_outputs(1301) <= (inputs(105)) xor (inputs(154));
    layer0_outputs(1302) <= not((inputs(40)) or (inputs(31)));
    layer0_outputs(1303) <= not((inputs(60)) or (inputs(84)));
    layer0_outputs(1304) <= (inputs(222)) xor (inputs(103));
    layer0_outputs(1305) <= (inputs(116)) xor (inputs(245));
    layer0_outputs(1306) <= (inputs(142)) or (inputs(101));
    layer0_outputs(1307) <= not(inputs(101)) or (inputs(228));
    layer0_outputs(1308) <= inputs(226);
    layer0_outputs(1309) <= not((inputs(13)) xor (inputs(247)));
    layer0_outputs(1310) <= not(inputs(102));
    layer0_outputs(1311) <= not(inputs(83)) or (inputs(114));
    layer0_outputs(1312) <= not((inputs(25)) or (inputs(158)));
    layer0_outputs(1313) <= (inputs(117)) and not (inputs(209));
    layer0_outputs(1314) <= (inputs(215)) or (inputs(123));
    layer0_outputs(1315) <= not(inputs(239)) or (inputs(160));
    layer0_outputs(1316) <= '1';
    layer0_outputs(1317) <= not((inputs(244)) or (inputs(30)));
    layer0_outputs(1318) <= inputs(27);
    layer0_outputs(1319) <= not((inputs(108)) or (inputs(119)));
    layer0_outputs(1320) <= (inputs(63)) xor (inputs(108));
    layer0_outputs(1321) <= not((inputs(199)) xor (inputs(70)));
    layer0_outputs(1322) <= (inputs(51)) or (inputs(170));
    layer0_outputs(1323) <= not((inputs(75)) and (inputs(251)));
    layer0_outputs(1324) <= (inputs(171)) and not (inputs(209));
    layer0_outputs(1325) <= not(inputs(64)) or (inputs(58));
    layer0_outputs(1326) <= inputs(243);
    layer0_outputs(1327) <= not(inputs(192));
    layer0_outputs(1328) <= (inputs(130)) xor (inputs(132));
    layer0_outputs(1329) <= (inputs(79)) and (inputs(251));
    layer0_outputs(1330) <= not(inputs(92)) or (inputs(241));
    layer0_outputs(1331) <= not((inputs(175)) xor (inputs(125)));
    layer0_outputs(1332) <= (inputs(154)) xor (inputs(125));
    layer0_outputs(1333) <= not((inputs(165)) xor (inputs(222)));
    layer0_outputs(1334) <= not(inputs(175));
    layer0_outputs(1335) <= inputs(252);
    layer0_outputs(1336) <= inputs(138);
    layer0_outputs(1337) <= not(inputs(119)) or (inputs(127));
    layer0_outputs(1338) <= (inputs(62)) or (inputs(134));
    layer0_outputs(1339) <= (inputs(252)) and not (inputs(141));
    layer0_outputs(1340) <= not((inputs(240)) xor (inputs(213)));
    layer0_outputs(1341) <= not((inputs(252)) or (inputs(1)));
    layer0_outputs(1342) <= (inputs(214)) and not (inputs(112));
    layer0_outputs(1343) <= not(inputs(195)) or (inputs(250));
    layer0_outputs(1344) <= not(inputs(155)) or (inputs(68));
    layer0_outputs(1345) <= not(inputs(167)) or (inputs(193));
    layer0_outputs(1346) <= (inputs(107)) and not (inputs(97));
    layer0_outputs(1347) <= (inputs(112)) or (inputs(108));
    layer0_outputs(1348) <= '0';
    layer0_outputs(1349) <= not(inputs(71)) or (inputs(167));
    layer0_outputs(1350) <= '1';
    layer0_outputs(1351) <= (inputs(89)) and not (inputs(233));
    layer0_outputs(1352) <= not(inputs(147));
    layer0_outputs(1353) <= not((inputs(227)) and (inputs(46)));
    layer0_outputs(1354) <= inputs(57);
    layer0_outputs(1355) <= (inputs(123)) xor (inputs(244));
    layer0_outputs(1356) <= inputs(204);
    layer0_outputs(1357) <= not((inputs(145)) or (inputs(156)));
    layer0_outputs(1358) <= (inputs(142)) or (inputs(234));
    layer0_outputs(1359) <= not(inputs(246)) or (inputs(128));
    layer0_outputs(1360) <= (inputs(48)) or (inputs(245));
    layer0_outputs(1361) <= (inputs(246)) xor (inputs(232));
    layer0_outputs(1362) <= inputs(40);
    layer0_outputs(1363) <= not(inputs(134));
    layer0_outputs(1364) <= (inputs(52)) and not (inputs(48));
    layer0_outputs(1365) <= (inputs(56)) or (inputs(99));
    layer0_outputs(1366) <= not((inputs(164)) or (inputs(67)));
    layer0_outputs(1367) <= inputs(153);
    layer0_outputs(1368) <= not((inputs(135)) or (inputs(208)));
    layer0_outputs(1369) <= not((inputs(212)) xor (inputs(109)));
    layer0_outputs(1370) <= inputs(59);
    layer0_outputs(1371) <= inputs(64);
    layer0_outputs(1372) <= (inputs(171)) and not (inputs(45));
    layer0_outputs(1373) <= not((inputs(93)) xor (inputs(130)));
    layer0_outputs(1374) <= not((inputs(40)) or (inputs(108)));
    layer0_outputs(1375) <= inputs(93);
    layer0_outputs(1376) <= not((inputs(200)) and (inputs(137)));
    layer0_outputs(1377) <= (inputs(226)) or (inputs(230));
    layer0_outputs(1378) <= inputs(220);
    layer0_outputs(1379) <= inputs(86);
    layer0_outputs(1380) <= not((inputs(154)) xor (inputs(107)));
    layer0_outputs(1381) <= inputs(102);
    layer0_outputs(1382) <= not(inputs(249));
    layer0_outputs(1383) <= not(inputs(13)) or (inputs(0));
    layer0_outputs(1384) <= inputs(60);
    layer0_outputs(1385) <= (inputs(162)) or (inputs(170));
    layer0_outputs(1386) <= (inputs(185)) or (inputs(138));
    layer0_outputs(1387) <= not((inputs(74)) or (inputs(50)));
    layer0_outputs(1388) <= (inputs(133)) or (inputs(79));
    layer0_outputs(1389) <= not((inputs(179)) xor (inputs(50)));
    layer0_outputs(1390) <= not((inputs(80)) xor (inputs(61)));
    layer0_outputs(1391) <= (inputs(214)) and not (inputs(183));
    layer0_outputs(1392) <= not(inputs(12)) or (inputs(205));
    layer0_outputs(1393) <= inputs(102);
    layer0_outputs(1394) <= (inputs(235)) or (inputs(202));
    layer0_outputs(1395) <= not((inputs(163)) xor (inputs(98)));
    layer0_outputs(1396) <= inputs(122);
    layer0_outputs(1397) <= (inputs(98)) or (inputs(136));
    layer0_outputs(1398) <= not(inputs(136));
    layer0_outputs(1399) <= not((inputs(149)) xor (inputs(220)));
    layer0_outputs(1400) <= (inputs(188)) and not (inputs(2));
    layer0_outputs(1401) <= not(inputs(29)) or (inputs(221));
    layer0_outputs(1402) <= not((inputs(211)) and (inputs(244)));
    layer0_outputs(1403) <= (inputs(249)) xor (inputs(210));
    layer0_outputs(1404) <= not(inputs(239)) or (inputs(25));
    layer0_outputs(1405) <= not(inputs(234));
    layer0_outputs(1406) <= not(inputs(43)) or (inputs(66));
    layer0_outputs(1407) <= not(inputs(84)) or (inputs(3));
    layer0_outputs(1408) <= (inputs(156)) xor (inputs(189));
    layer0_outputs(1409) <= not((inputs(54)) xor (inputs(247)));
    layer0_outputs(1410) <= (inputs(133)) and not (inputs(52));
    layer0_outputs(1411) <= inputs(207);
    layer0_outputs(1412) <= (inputs(127)) and not (inputs(113));
    layer0_outputs(1413) <= inputs(36);
    layer0_outputs(1414) <= (inputs(119)) and not (inputs(167));
    layer0_outputs(1415) <= not((inputs(193)) xor (inputs(6)));
    layer0_outputs(1416) <= inputs(157);
    layer0_outputs(1417) <= inputs(165);
    layer0_outputs(1418) <= (inputs(20)) or (inputs(74));
    layer0_outputs(1419) <= not(inputs(188)) or (inputs(11));
    layer0_outputs(1420) <= not(inputs(103)) or (inputs(98));
    layer0_outputs(1421) <= not(inputs(150));
    layer0_outputs(1422) <= inputs(221);
    layer0_outputs(1423) <= not((inputs(221)) xor (inputs(135)));
    layer0_outputs(1424) <= (inputs(137)) xor (inputs(122));
    layer0_outputs(1425) <= inputs(195);
    layer0_outputs(1426) <= (inputs(126)) xor (inputs(247));
    layer0_outputs(1427) <= not(inputs(107));
    layer0_outputs(1428) <= not(inputs(217)) or (inputs(20));
    layer0_outputs(1429) <= (inputs(215)) and not (inputs(10));
    layer0_outputs(1430) <= inputs(88);
    layer0_outputs(1431) <= not(inputs(146)) or (inputs(236));
    layer0_outputs(1432) <= '1';
    layer0_outputs(1433) <= (inputs(74)) xor (inputs(139));
    layer0_outputs(1434) <= not(inputs(217));
    layer0_outputs(1435) <= inputs(168);
    layer0_outputs(1436) <= inputs(185);
    layer0_outputs(1437) <= (inputs(108)) and not (inputs(205));
    layer0_outputs(1438) <= not((inputs(67)) or (inputs(70)));
    layer0_outputs(1439) <= not(inputs(81)) or (inputs(46));
    layer0_outputs(1440) <= not(inputs(147));
    layer0_outputs(1441) <= (inputs(76)) and not (inputs(147));
    layer0_outputs(1442) <= (inputs(187)) or (inputs(195));
    layer0_outputs(1443) <= not((inputs(90)) or (inputs(162)));
    layer0_outputs(1444) <= inputs(234);
    layer0_outputs(1445) <= not(inputs(37)) or (inputs(244));
    layer0_outputs(1446) <= not(inputs(120)) or (inputs(158));
    layer0_outputs(1447) <= not((inputs(188)) or (inputs(213)));
    layer0_outputs(1448) <= (inputs(181)) and not (inputs(159));
    layer0_outputs(1449) <= (inputs(35)) or (inputs(55));
    layer0_outputs(1450) <= not((inputs(140)) xor (inputs(255)));
    layer0_outputs(1451) <= not((inputs(166)) xor (inputs(148)));
    layer0_outputs(1452) <= not((inputs(179)) or (inputs(158)));
    layer0_outputs(1453) <= inputs(132);
    layer0_outputs(1454) <= not(inputs(124)) or (inputs(129));
    layer0_outputs(1455) <= not((inputs(204)) xor (inputs(225)));
    layer0_outputs(1456) <= not(inputs(191)) or (inputs(253));
    layer0_outputs(1457) <= not(inputs(141));
    layer0_outputs(1458) <= (inputs(238)) and not (inputs(159));
    layer0_outputs(1459) <= not(inputs(151)) or (inputs(57));
    layer0_outputs(1460) <= not((inputs(160)) or (inputs(213)));
    layer0_outputs(1461) <= not(inputs(115));
    layer0_outputs(1462) <= (inputs(6)) or (inputs(28));
    layer0_outputs(1463) <= (inputs(52)) or (inputs(6));
    layer0_outputs(1464) <= not(inputs(57)) or (inputs(154));
    layer0_outputs(1465) <= not((inputs(154)) xor (inputs(1)));
    layer0_outputs(1466) <= (inputs(63)) and (inputs(234));
    layer0_outputs(1467) <= (inputs(138)) or (inputs(230));
    layer0_outputs(1468) <= inputs(136);
    layer0_outputs(1469) <= not((inputs(103)) xor (inputs(17)));
    layer0_outputs(1470) <= not(inputs(159)) or (inputs(5));
    layer0_outputs(1471) <= (inputs(249)) xor (inputs(238));
    layer0_outputs(1472) <= not(inputs(100));
    layer0_outputs(1473) <= (inputs(140)) and not (inputs(203));
    layer0_outputs(1474) <= (inputs(44)) and not (inputs(29));
    layer0_outputs(1475) <= (inputs(202)) or (inputs(174));
    layer0_outputs(1476) <= (inputs(199)) and not (inputs(126));
    layer0_outputs(1477) <= (inputs(82)) or (inputs(246));
    layer0_outputs(1478) <= inputs(152);
    layer0_outputs(1479) <= inputs(42);
    layer0_outputs(1480) <= (inputs(164)) and not (inputs(130));
    layer0_outputs(1481) <= not(inputs(229));
    layer0_outputs(1482) <= not(inputs(163));
    layer0_outputs(1483) <= inputs(73);
    layer0_outputs(1484) <= (inputs(105)) and not (inputs(96));
    layer0_outputs(1485) <= (inputs(207)) and (inputs(192));
    layer0_outputs(1486) <= inputs(199);
    layer0_outputs(1487) <= not((inputs(56)) or (inputs(193)));
    layer0_outputs(1488) <= '0';
    layer0_outputs(1489) <= (inputs(118)) and not (inputs(66));
    layer0_outputs(1490) <= (inputs(229)) and not (inputs(43));
    layer0_outputs(1491) <= inputs(90);
    layer0_outputs(1492) <= (inputs(168)) and not (inputs(179));
    layer0_outputs(1493) <= '0';
    layer0_outputs(1494) <= '0';
    layer0_outputs(1495) <= not((inputs(15)) xor (inputs(116)));
    layer0_outputs(1496) <= inputs(92);
    layer0_outputs(1497) <= not((inputs(78)) or (inputs(239)));
    layer0_outputs(1498) <= (inputs(236)) xor (inputs(122));
    layer0_outputs(1499) <= inputs(99);
    layer0_outputs(1500) <= not(inputs(215));
    layer0_outputs(1501) <= '0';
    layer0_outputs(1502) <= not((inputs(190)) and (inputs(32)));
    layer0_outputs(1503) <= inputs(249);
    layer0_outputs(1504) <= not(inputs(76));
    layer0_outputs(1505) <= (inputs(207)) and not (inputs(8));
    layer0_outputs(1506) <= not((inputs(10)) xor (inputs(36)));
    layer0_outputs(1507) <= not((inputs(226)) or (inputs(151)));
    layer0_outputs(1508) <= not((inputs(24)) and (inputs(79)));
    layer0_outputs(1509) <= not(inputs(44)) or (inputs(4));
    layer0_outputs(1510) <= '0';
    layer0_outputs(1511) <= inputs(97);
    layer0_outputs(1512) <= (inputs(2)) or (inputs(135));
    layer0_outputs(1513) <= (inputs(228)) and not (inputs(248));
    layer0_outputs(1514) <= '1';
    layer0_outputs(1515) <= not(inputs(104)) or (inputs(99));
    layer0_outputs(1516) <= not((inputs(166)) or (inputs(30)));
    layer0_outputs(1517) <= '0';
    layer0_outputs(1518) <= (inputs(80)) xor (inputs(250));
    layer0_outputs(1519) <= not(inputs(13)) or (inputs(45));
    layer0_outputs(1520) <= (inputs(73)) and not (inputs(113));
    layer0_outputs(1521) <= not(inputs(46)) or (inputs(185));
    layer0_outputs(1522) <= not(inputs(175));
    layer0_outputs(1523) <= (inputs(139)) xor (inputs(156));
    layer0_outputs(1524) <= not(inputs(192));
    layer0_outputs(1525) <= (inputs(201)) or (inputs(110));
    layer0_outputs(1526) <= not(inputs(222));
    layer0_outputs(1527) <= (inputs(218)) xor (inputs(24));
    layer0_outputs(1528) <= not((inputs(160)) and (inputs(29)));
    layer0_outputs(1529) <= (inputs(17)) and not (inputs(10));
    layer0_outputs(1530) <= not(inputs(237)) or (inputs(110));
    layer0_outputs(1531) <= (inputs(154)) and not (inputs(30));
    layer0_outputs(1532) <= not((inputs(46)) or (inputs(197)));
    layer0_outputs(1533) <= not((inputs(63)) xor (inputs(188)));
    layer0_outputs(1534) <= not(inputs(22));
    layer0_outputs(1535) <= (inputs(57)) or (inputs(79));
    layer0_outputs(1536) <= (inputs(94)) and not (inputs(211));
    layer0_outputs(1537) <= (inputs(113)) xor (inputs(137));
    layer0_outputs(1538) <= (inputs(232)) or (inputs(86));
    layer0_outputs(1539) <= (inputs(153)) xor (inputs(60));
    layer0_outputs(1540) <= '0';
    layer0_outputs(1541) <= not((inputs(90)) and (inputs(136)));
    layer0_outputs(1542) <= not((inputs(37)) or (inputs(227)));
    layer0_outputs(1543) <= not((inputs(113)) or (inputs(127)));
    layer0_outputs(1544) <= (inputs(131)) or (inputs(49));
    layer0_outputs(1545) <= (inputs(101)) and not (inputs(24));
    layer0_outputs(1546) <= (inputs(92)) xor (inputs(198));
    layer0_outputs(1547) <= '0';
    layer0_outputs(1548) <= inputs(124);
    layer0_outputs(1549) <= not((inputs(230)) xor (inputs(28)));
    layer0_outputs(1550) <= (inputs(182)) or (inputs(231));
    layer0_outputs(1551) <= not((inputs(247)) or (inputs(10)));
    layer0_outputs(1552) <= not((inputs(208)) xor (inputs(136)));
    layer0_outputs(1553) <= (inputs(190)) and (inputs(223));
    layer0_outputs(1554) <= (inputs(107)) or (inputs(146));
    layer0_outputs(1555) <= (inputs(192)) xor (inputs(90));
    layer0_outputs(1556) <= inputs(188);
    layer0_outputs(1557) <= (inputs(131)) or (inputs(124));
    layer0_outputs(1558) <= not((inputs(195)) or (inputs(146)));
    layer0_outputs(1559) <= (inputs(166)) or (inputs(101));
    layer0_outputs(1560) <= (inputs(217)) and not (inputs(155));
    layer0_outputs(1561) <= not(inputs(38)) or (inputs(83));
    layer0_outputs(1562) <= not((inputs(201)) or (inputs(182)));
    layer0_outputs(1563) <= not(inputs(136));
    layer0_outputs(1564) <= (inputs(205)) or (inputs(151));
    layer0_outputs(1565) <= (inputs(84)) and not (inputs(235));
    layer0_outputs(1566) <= inputs(42);
    layer0_outputs(1567) <= inputs(198);
    layer0_outputs(1568) <= (inputs(212)) and (inputs(28));
    layer0_outputs(1569) <= (inputs(186)) and not (inputs(117));
    layer0_outputs(1570) <= (inputs(84)) or (inputs(165));
    layer0_outputs(1571) <= not((inputs(203)) or (inputs(82)));
    layer0_outputs(1572) <= not(inputs(190));
    layer0_outputs(1573) <= not((inputs(252)) and (inputs(111)));
    layer0_outputs(1574) <= not(inputs(48)) or (inputs(98));
    layer0_outputs(1575) <= (inputs(2)) or (inputs(188));
    layer0_outputs(1576) <= (inputs(113)) and not (inputs(29));
    layer0_outputs(1577) <= (inputs(169)) and not (inputs(36));
    layer0_outputs(1578) <= inputs(233);
    layer0_outputs(1579) <= not(inputs(185));
    layer0_outputs(1580) <= not(inputs(202)) or (inputs(48));
    layer0_outputs(1581) <= not((inputs(57)) or (inputs(104)));
    layer0_outputs(1582) <= not(inputs(155));
    layer0_outputs(1583) <= not(inputs(9)) or (inputs(45));
    layer0_outputs(1584) <= '1';
    layer0_outputs(1585) <= not((inputs(86)) or (inputs(102)));
    layer0_outputs(1586) <= not((inputs(89)) xor (inputs(5)));
    layer0_outputs(1587) <= not(inputs(194)) or (inputs(66));
    layer0_outputs(1588) <= not((inputs(10)) or (inputs(142)));
    layer0_outputs(1589) <= (inputs(204)) xor (inputs(28));
    layer0_outputs(1590) <= (inputs(23)) and not (inputs(42));
    layer0_outputs(1591) <= (inputs(158)) or (inputs(105));
    layer0_outputs(1592) <= '0';
    layer0_outputs(1593) <= not((inputs(14)) xor (inputs(23)));
    layer0_outputs(1594) <= (inputs(140)) or (inputs(76));
    layer0_outputs(1595) <= inputs(57);
    layer0_outputs(1596) <= not((inputs(7)) xor (inputs(166)));
    layer0_outputs(1597) <= not(inputs(13));
    layer0_outputs(1598) <= not(inputs(200));
    layer0_outputs(1599) <= (inputs(171)) xor (inputs(247));
    layer0_outputs(1600) <= not((inputs(215)) xor (inputs(230)));
    layer0_outputs(1601) <= not((inputs(207)) xor (inputs(33)));
    layer0_outputs(1602) <= (inputs(148)) or (inputs(24));
    layer0_outputs(1603) <= not((inputs(107)) xor (inputs(254)));
    layer0_outputs(1604) <= (inputs(121)) and (inputs(195));
    layer0_outputs(1605) <= not((inputs(105)) xor (inputs(17)));
    layer0_outputs(1606) <= not((inputs(69)) xor (inputs(139)));
    layer0_outputs(1607) <= (inputs(219)) xor (inputs(12));
    layer0_outputs(1608) <= not(inputs(177)) or (inputs(241));
    layer0_outputs(1609) <= inputs(156);
    layer0_outputs(1610) <= (inputs(26)) and not (inputs(222));
    layer0_outputs(1611) <= (inputs(101)) and not (inputs(242));
    layer0_outputs(1612) <= not(inputs(184));
    layer0_outputs(1613) <= not(inputs(214));
    layer0_outputs(1614) <= not(inputs(15)) or (inputs(124));
    layer0_outputs(1615) <= not((inputs(78)) xor (inputs(237)));
    layer0_outputs(1616) <= not((inputs(1)) xor (inputs(213)));
    layer0_outputs(1617) <= inputs(128);
    layer0_outputs(1618) <= not((inputs(72)) or (inputs(135)));
    layer0_outputs(1619) <= not(inputs(82)) or (inputs(64));
    layer0_outputs(1620) <= not(inputs(132));
    layer0_outputs(1621) <= inputs(197);
    layer0_outputs(1622) <= not(inputs(152));
    layer0_outputs(1623) <= (inputs(136)) or (inputs(93));
    layer0_outputs(1624) <= not((inputs(103)) or (inputs(228)));
    layer0_outputs(1625) <= (inputs(220)) or (inputs(155));
    layer0_outputs(1626) <= not((inputs(56)) xor (inputs(205)));
    layer0_outputs(1627) <= not((inputs(23)) or (inputs(98)));
    layer0_outputs(1628) <= not(inputs(105)) or (inputs(5));
    layer0_outputs(1629) <= not((inputs(93)) or (inputs(141)));
    layer0_outputs(1630) <= (inputs(226)) xor (inputs(95));
    layer0_outputs(1631) <= not((inputs(98)) xor (inputs(96)));
    layer0_outputs(1632) <= not((inputs(114)) xor (inputs(148)));
    layer0_outputs(1633) <= not((inputs(90)) or (inputs(73)));
    layer0_outputs(1634) <= not(inputs(137));
    layer0_outputs(1635) <= (inputs(38)) or (inputs(171));
    layer0_outputs(1636) <= (inputs(67)) or (inputs(38));
    layer0_outputs(1637) <= not((inputs(216)) xor (inputs(114)));
    layer0_outputs(1638) <= not((inputs(239)) or (inputs(186)));
    layer0_outputs(1639) <= (inputs(25)) xor (inputs(161));
    layer0_outputs(1640) <= not((inputs(17)) xor (inputs(53)));
    layer0_outputs(1641) <= (inputs(120)) and not (inputs(35));
    layer0_outputs(1642) <= not((inputs(55)) or (inputs(185)));
    layer0_outputs(1643) <= not(inputs(181));
    layer0_outputs(1644) <= (inputs(164)) or (inputs(13));
    layer0_outputs(1645) <= (inputs(212)) or (inputs(145));
    layer0_outputs(1646) <= (inputs(235)) and (inputs(81));
    layer0_outputs(1647) <= not(inputs(49));
    layer0_outputs(1648) <= inputs(164);
    layer0_outputs(1649) <= not(inputs(208));
    layer0_outputs(1650) <= inputs(51);
    layer0_outputs(1651) <= (inputs(201)) and not (inputs(190));
    layer0_outputs(1652) <= (inputs(238)) and (inputs(66));
    layer0_outputs(1653) <= not((inputs(5)) or (inputs(146)));
    layer0_outputs(1654) <= not((inputs(123)) xor (inputs(255)));
    layer0_outputs(1655) <= (inputs(138)) or (inputs(4));
    layer0_outputs(1656) <= (inputs(133)) xor (inputs(3));
    layer0_outputs(1657) <= inputs(140);
    layer0_outputs(1658) <= (inputs(214)) xor (inputs(129));
    layer0_outputs(1659) <= (inputs(151)) and not (inputs(67));
    layer0_outputs(1660) <= not((inputs(66)) or (inputs(89)));
    layer0_outputs(1661) <= (inputs(203)) or (inputs(38));
    layer0_outputs(1662) <= (inputs(178)) or (inputs(49));
    layer0_outputs(1663) <= (inputs(67)) xor (inputs(102));
    layer0_outputs(1664) <= (inputs(22)) and not (inputs(251));
    layer0_outputs(1665) <= not((inputs(202)) xor (inputs(15)));
    layer0_outputs(1666) <= (inputs(26)) or (inputs(134));
    layer0_outputs(1667) <= inputs(174);
    layer0_outputs(1668) <= not(inputs(161)) or (inputs(65));
    layer0_outputs(1669) <= not(inputs(183)) or (inputs(237));
    layer0_outputs(1670) <= not(inputs(135)) or (inputs(113));
    layer0_outputs(1671) <= (inputs(52)) and not (inputs(227));
    layer0_outputs(1672) <= (inputs(38)) xor (inputs(159));
    layer0_outputs(1673) <= not((inputs(89)) or (inputs(195)));
    layer0_outputs(1674) <= not((inputs(30)) or (inputs(113)));
    layer0_outputs(1675) <= not((inputs(165)) or (inputs(225)));
    layer0_outputs(1676) <= inputs(75);
    layer0_outputs(1677) <= inputs(172);
    layer0_outputs(1678) <= not((inputs(209)) and (inputs(254)));
    layer0_outputs(1679) <= not(inputs(186));
    layer0_outputs(1680) <= not((inputs(60)) or (inputs(166)));
    layer0_outputs(1681) <= not((inputs(53)) xor (inputs(107)));
    layer0_outputs(1682) <= not(inputs(206)) or (inputs(48));
    layer0_outputs(1683) <= (inputs(135)) and not (inputs(40));
    layer0_outputs(1684) <= not((inputs(90)) or (inputs(250)));
    layer0_outputs(1685) <= not(inputs(88)) or (inputs(62));
    layer0_outputs(1686) <= inputs(29);
    layer0_outputs(1687) <= not(inputs(40)) or (inputs(65));
    layer0_outputs(1688) <= (inputs(164)) xor (inputs(120));
    layer0_outputs(1689) <= not((inputs(23)) or (inputs(183)));
    layer0_outputs(1690) <= (inputs(112)) xor (inputs(157));
    layer0_outputs(1691) <= (inputs(231)) or (inputs(86));
    layer0_outputs(1692) <= not(inputs(202));
    layer0_outputs(1693) <= not((inputs(121)) or (inputs(79)));
    layer0_outputs(1694) <= not(inputs(206)) or (inputs(73));
    layer0_outputs(1695) <= not(inputs(102));
    layer0_outputs(1696) <= not((inputs(76)) or (inputs(139)));
    layer0_outputs(1697) <= not((inputs(197)) or (inputs(69)));
    layer0_outputs(1698) <= not((inputs(144)) or (inputs(112)));
    layer0_outputs(1699) <= not((inputs(197)) and (inputs(252)));
    layer0_outputs(1700) <= (inputs(7)) or (inputs(249));
    layer0_outputs(1701) <= (inputs(232)) and not (inputs(211));
    layer0_outputs(1702) <= (inputs(50)) and (inputs(210));
    layer0_outputs(1703) <= not((inputs(219)) or (inputs(93)));
    layer0_outputs(1704) <= not(inputs(171)) or (inputs(34));
    layer0_outputs(1705) <= not(inputs(222));
    layer0_outputs(1706) <= (inputs(94)) or (inputs(215));
    layer0_outputs(1707) <= (inputs(190)) and not (inputs(242));
    layer0_outputs(1708) <= not(inputs(101)) or (inputs(82));
    layer0_outputs(1709) <= inputs(105);
    layer0_outputs(1710) <= not((inputs(150)) xor (inputs(45)));
    layer0_outputs(1711) <= (inputs(175)) xor (inputs(186));
    layer0_outputs(1712) <= inputs(120);
    layer0_outputs(1713) <= '1';
    layer0_outputs(1714) <= inputs(79);
    layer0_outputs(1715) <= (inputs(171)) xor (inputs(30));
    layer0_outputs(1716) <= not((inputs(217)) and (inputs(167)));
    layer0_outputs(1717) <= inputs(63);
    layer0_outputs(1718) <= (inputs(7)) and not (inputs(250));
    layer0_outputs(1719) <= not(inputs(2)) or (inputs(207));
    layer0_outputs(1720) <= '1';
    layer0_outputs(1721) <= not((inputs(193)) and (inputs(234)));
    layer0_outputs(1722) <= not(inputs(110)) or (inputs(241));
    layer0_outputs(1723) <= not(inputs(128));
    layer0_outputs(1724) <= inputs(109);
    layer0_outputs(1725) <= inputs(210);
    layer0_outputs(1726) <= not((inputs(159)) or (inputs(138)));
    layer0_outputs(1727) <= not((inputs(53)) or (inputs(184)));
    layer0_outputs(1728) <= not(inputs(103));
    layer0_outputs(1729) <= not((inputs(197)) or (inputs(76)));
    layer0_outputs(1730) <= not(inputs(85));
    layer0_outputs(1731) <= not(inputs(124)) or (inputs(109));
    layer0_outputs(1732) <= inputs(104);
    layer0_outputs(1733) <= (inputs(215)) or (inputs(77));
    layer0_outputs(1734) <= (inputs(234)) or (inputs(33));
    layer0_outputs(1735) <= not(inputs(135));
    layer0_outputs(1736) <= inputs(237);
    layer0_outputs(1737) <= not(inputs(122));
    layer0_outputs(1738) <= inputs(76);
    layer0_outputs(1739) <= (inputs(170)) or (inputs(30));
    layer0_outputs(1740) <= not(inputs(75)) or (inputs(94));
    layer0_outputs(1741) <= (inputs(171)) and not (inputs(61));
    layer0_outputs(1742) <= not((inputs(137)) or (inputs(232)));
    layer0_outputs(1743) <= (inputs(245)) and not (inputs(12));
    layer0_outputs(1744) <= inputs(150);
    layer0_outputs(1745) <= not((inputs(253)) and (inputs(158)));
    layer0_outputs(1746) <= (inputs(202)) or (inputs(252));
    layer0_outputs(1747) <= inputs(134);
    layer0_outputs(1748) <= not(inputs(131));
    layer0_outputs(1749) <= not((inputs(58)) xor (inputs(29)));
    layer0_outputs(1750) <= (inputs(28)) and not (inputs(226));
    layer0_outputs(1751) <= '1';
    layer0_outputs(1752) <= (inputs(105)) xor (inputs(145));
    layer0_outputs(1753) <= not((inputs(104)) or (inputs(196)));
    layer0_outputs(1754) <= (inputs(151)) and not (inputs(27));
    layer0_outputs(1755) <= (inputs(83)) xor (inputs(32));
    layer0_outputs(1756) <= inputs(92);
    layer0_outputs(1757) <= (inputs(41)) or (inputs(228));
    layer0_outputs(1758) <= (inputs(201)) and not (inputs(150));
    layer0_outputs(1759) <= '0';
    layer0_outputs(1760) <= (inputs(37)) xor (inputs(149));
    layer0_outputs(1761) <= not((inputs(212)) xor (inputs(3)));
    layer0_outputs(1762) <= not((inputs(211)) or (inputs(236)));
    layer0_outputs(1763) <= not(inputs(169)) or (inputs(216));
    layer0_outputs(1764) <= not(inputs(218));
    layer0_outputs(1765) <= not(inputs(167)) or (inputs(162));
    layer0_outputs(1766) <= not((inputs(120)) xor (inputs(9)));
    layer0_outputs(1767) <= (inputs(76)) and (inputs(173));
    layer0_outputs(1768) <= (inputs(106)) and not (inputs(246));
    layer0_outputs(1769) <= not(inputs(155)) or (inputs(18));
    layer0_outputs(1770) <= not((inputs(169)) xor (inputs(127)));
    layer0_outputs(1771) <= not(inputs(154));
    layer0_outputs(1772) <= not(inputs(90)) or (inputs(114));
    layer0_outputs(1773) <= not(inputs(75));
    layer0_outputs(1774) <= inputs(227);
    layer0_outputs(1775) <= not(inputs(87)) or (inputs(152));
    layer0_outputs(1776) <= inputs(56);
    layer0_outputs(1777) <= not(inputs(118));
    layer0_outputs(1778) <= not((inputs(223)) xor (inputs(197)));
    layer0_outputs(1779) <= (inputs(235)) xor (inputs(221));
    layer0_outputs(1780) <= not((inputs(169)) or (inputs(126)));
    layer0_outputs(1781) <= inputs(181);
    layer0_outputs(1782) <= not(inputs(231)) or (inputs(59));
    layer0_outputs(1783) <= not((inputs(1)) and (inputs(112)));
    layer0_outputs(1784) <= not((inputs(75)) xor (inputs(52)));
    layer0_outputs(1785) <= (inputs(218)) and not (inputs(212));
    layer0_outputs(1786) <= (inputs(74)) or (inputs(214));
    layer0_outputs(1787) <= (inputs(236)) xor (inputs(152));
    layer0_outputs(1788) <= (inputs(109)) xor (inputs(76));
    layer0_outputs(1789) <= not(inputs(72)) or (inputs(26));
    layer0_outputs(1790) <= not((inputs(103)) xor (inputs(79)));
    layer0_outputs(1791) <= inputs(59);
    layer0_outputs(1792) <= (inputs(198)) or (inputs(33));
    layer0_outputs(1793) <= (inputs(246)) xor (inputs(214));
    layer0_outputs(1794) <= not(inputs(236)) or (inputs(209));
    layer0_outputs(1795) <= not(inputs(118));
    layer0_outputs(1796) <= inputs(85);
    layer0_outputs(1797) <= (inputs(46)) and not (inputs(30));
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= not(inputs(187)) or (inputs(98));
    layer0_outputs(1800) <= not((inputs(35)) or (inputs(201)));
    layer0_outputs(1801) <= not((inputs(187)) or (inputs(206)));
    layer0_outputs(1802) <= not((inputs(181)) or (inputs(189)));
    layer0_outputs(1803) <= (inputs(168)) and not (inputs(217));
    layer0_outputs(1804) <= (inputs(132)) xor (inputs(241));
    layer0_outputs(1805) <= not(inputs(59)) or (inputs(234));
    layer0_outputs(1806) <= (inputs(38)) xor (inputs(252));
    layer0_outputs(1807) <= inputs(94);
    layer0_outputs(1808) <= (inputs(201)) and not (inputs(98));
    layer0_outputs(1809) <= not(inputs(55));
    layer0_outputs(1810) <= not(inputs(200)) or (inputs(24));
    layer0_outputs(1811) <= not((inputs(58)) or (inputs(180)));
    layer0_outputs(1812) <= not(inputs(177));
    layer0_outputs(1813) <= (inputs(194)) or (inputs(165));
    layer0_outputs(1814) <= (inputs(59)) or (inputs(149));
    layer0_outputs(1815) <= not(inputs(202));
    layer0_outputs(1816) <= '1';
    layer0_outputs(1817) <= not(inputs(78));
    layer0_outputs(1818) <= not(inputs(54));
    layer0_outputs(1819) <= inputs(93);
    layer0_outputs(1820) <= inputs(100);
    layer0_outputs(1821) <= not(inputs(134)) or (inputs(6));
    layer0_outputs(1822) <= not((inputs(204)) xor (inputs(86)));
    layer0_outputs(1823) <= (inputs(158)) xor (inputs(239));
    layer0_outputs(1824) <= (inputs(87)) and not (inputs(139));
    layer0_outputs(1825) <= not(inputs(121)) or (inputs(166));
    layer0_outputs(1826) <= not((inputs(203)) or (inputs(232)));
    layer0_outputs(1827) <= not(inputs(186));
    layer0_outputs(1828) <= not((inputs(46)) xor (inputs(197)));
    layer0_outputs(1829) <= not((inputs(63)) xor (inputs(125)));
    layer0_outputs(1830) <= not((inputs(212)) or (inputs(191)));
    layer0_outputs(1831) <= not(inputs(147));
    layer0_outputs(1832) <= (inputs(152)) or (inputs(10));
    layer0_outputs(1833) <= (inputs(160)) and (inputs(191));
    layer0_outputs(1834) <= '1';
    layer0_outputs(1835) <= not((inputs(236)) and (inputs(158)));
    layer0_outputs(1836) <= not((inputs(169)) or (inputs(91)));
    layer0_outputs(1837) <= not((inputs(241)) or (inputs(93)));
    layer0_outputs(1838) <= (inputs(221)) or (inputs(96));
    layer0_outputs(1839) <= (inputs(142)) xor (inputs(156));
    layer0_outputs(1840) <= (inputs(185)) or (inputs(73));
    layer0_outputs(1841) <= (inputs(129)) or (inputs(93));
    layer0_outputs(1842) <= not(inputs(123));
    layer0_outputs(1843) <= (inputs(173)) and (inputs(27));
    layer0_outputs(1844) <= not((inputs(67)) or (inputs(67)));
    layer0_outputs(1845) <= (inputs(199)) or (inputs(66));
    layer0_outputs(1846) <= (inputs(98)) and not (inputs(8));
    layer0_outputs(1847) <= (inputs(174)) and (inputs(237));
    layer0_outputs(1848) <= not((inputs(247)) or (inputs(170)));
    layer0_outputs(1849) <= (inputs(249)) xor (inputs(93));
    layer0_outputs(1850) <= not((inputs(56)) or (inputs(40)));
    layer0_outputs(1851) <= not(inputs(198)) or (inputs(97));
    layer0_outputs(1852) <= (inputs(150)) xor (inputs(157));
    layer0_outputs(1853) <= not(inputs(203)) or (inputs(237));
    layer0_outputs(1854) <= not(inputs(181)) or (inputs(45));
    layer0_outputs(1855) <= inputs(76);
    layer0_outputs(1856) <= not((inputs(105)) and (inputs(142)));
    layer0_outputs(1857) <= (inputs(54)) and not (inputs(227));
    layer0_outputs(1858) <= not((inputs(139)) xor (inputs(172)));
    layer0_outputs(1859) <= (inputs(21)) and not (inputs(72));
    layer0_outputs(1860) <= (inputs(96)) or (inputs(199));
    layer0_outputs(1861) <= (inputs(126)) or (inputs(115));
    layer0_outputs(1862) <= not(inputs(128)) or (inputs(8));
    layer0_outputs(1863) <= (inputs(17)) xor (inputs(137));
    layer0_outputs(1864) <= not((inputs(92)) xor (inputs(113)));
    layer0_outputs(1865) <= not((inputs(163)) and (inputs(254)));
    layer0_outputs(1866) <= (inputs(221)) xor (inputs(101));
    layer0_outputs(1867) <= inputs(118);
    layer0_outputs(1868) <= (inputs(115)) or (inputs(187));
    layer0_outputs(1869) <= not(inputs(206));
    layer0_outputs(1870) <= (inputs(212)) or (inputs(171));
    layer0_outputs(1871) <= not((inputs(239)) and (inputs(98)));
    layer0_outputs(1872) <= (inputs(75)) and not (inputs(82));
    layer0_outputs(1873) <= not(inputs(107));
    layer0_outputs(1874) <= (inputs(86)) or (inputs(244));
    layer0_outputs(1875) <= inputs(135);
    layer0_outputs(1876) <= (inputs(66)) xor (inputs(76));
    layer0_outputs(1877) <= not((inputs(110)) xor (inputs(124)));
    layer0_outputs(1878) <= (inputs(2)) and not (inputs(211));
    layer0_outputs(1879) <= inputs(106);
    layer0_outputs(1880) <= inputs(166);
    layer0_outputs(1881) <= not((inputs(99)) and (inputs(16)));
    layer0_outputs(1882) <= (inputs(117)) xor (inputs(114));
    layer0_outputs(1883) <= (inputs(164)) or (inputs(57));
    layer0_outputs(1884) <= (inputs(182)) and not (inputs(228));
    layer0_outputs(1885) <= (inputs(54)) xor (inputs(234));
    layer0_outputs(1886) <= (inputs(170)) xor (inputs(37));
    layer0_outputs(1887) <= (inputs(203)) or (inputs(4));
    layer0_outputs(1888) <= (inputs(237)) xor (inputs(58));
    layer0_outputs(1889) <= (inputs(7)) or (inputs(254));
    layer0_outputs(1890) <= inputs(165);
    layer0_outputs(1891) <= (inputs(230)) or (inputs(67));
    layer0_outputs(1892) <= (inputs(149)) and not (inputs(189));
    layer0_outputs(1893) <= (inputs(87)) or (inputs(4));
    layer0_outputs(1894) <= (inputs(213)) xor (inputs(191));
    layer0_outputs(1895) <= not(inputs(131)) or (inputs(245));
    layer0_outputs(1896) <= not((inputs(10)) xor (inputs(83)));
    layer0_outputs(1897) <= not((inputs(140)) or (inputs(25)));
    layer0_outputs(1898) <= '1';
    layer0_outputs(1899) <= not(inputs(208)) or (inputs(102));
    layer0_outputs(1900) <= not(inputs(166));
    layer0_outputs(1901) <= not((inputs(38)) xor (inputs(210)));
    layer0_outputs(1902) <= not((inputs(34)) or (inputs(212)));
    layer0_outputs(1903) <= (inputs(198)) and not (inputs(100));
    layer0_outputs(1904) <= '1';
    layer0_outputs(1905) <= (inputs(228)) xor (inputs(231));
    layer0_outputs(1906) <= not((inputs(176)) or (inputs(96)));
    layer0_outputs(1907) <= inputs(81);
    layer0_outputs(1908) <= (inputs(229)) xor (inputs(56));
    layer0_outputs(1909) <= (inputs(24)) and not (inputs(204));
    layer0_outputs(1910) <= (inputs(87)) and not (inputs(129));
    layer0_outputs(1911) <= not((inputs(212)) or (inputs(196)));
    layer0_outputs(1912) <= not(inputs(157)) or (inputs(250));
    layer0_outputs(1913) <= not((inputs(232)) or (inputs(131)));
    layer0_outputs(1914) <= inputs(90);
    layer0_outputs(1915) <= (inputs(26)) and not (inputs(130));
    layer0_outputs(1916) <= '0';
    layer0_outputs(1917) <= (inputs(93)) and not (inputs(131));
    layer0_outputs(1918) <= not(inputs(252)) or (inputs(186));
    layer0_outputs(1919) <= (inputs(71)) and not (inputs(49));
    layer0_outputs(1920) <= not(inputs(51)) or (inputs(29));
    layer0_outputs(1921) <= not((inputs(128)) xor (inputs(192)));
    layer0_outputs(1922) <= not(inputs(108));
    layer0_outputs(1923) <= not(inputs(181));
    layer0_outputs(1924) <= not((inputs(189)) or (inputs(206)));
    layer0_outputs(1925) <= (inputs(46)) and not (inputs(214));
    layer0_outputs(1926) <= '0';
    layer0_outputs(1927) <= not((inputs(11)) or (inputs(233)));
    layer0_outputs(1928) <= (inputs(29)) or (inputs(215));
    layer0_outputs(1929) <= (inputs(112)) xor (inputs(90));
    layer0_outputs(1930) <= not((inputs(16)) xor (inputs(141)));
    layer0_outputs(1931) <= inputs(85);
    layer0_outputs(1932) <= not((inputs(203)) and (inputs(127)));
    layer0_outputs(1933) <= not(inputs(109)) or (inputs(132));
    layer0_outputs(1934) <= not(inputs(116));
    layer0_outputs(1935) <= inputs(73);
    layer0_outputs(1936) <= (inputs(211)) or (inputs(22));
    layer0_outputs(1937) <= (inputs(40)) and not (inputs(7));
    layer0_outputs(1938) <= not(inputs(122));
    layer0_outputs(1939) <= (inputs(33)) or (inputs(105));
    layer0_outputs(1940) <= not((inputs(177)) xor (inputs(212)));
    layer0_outputs(1941) <= not((inputs(228)) or (inputs(119)));
    layer0_outputs(1942) <= not((inputs(17)) xor (inputs(140)));
    layer0_outputs(1943) <= (inputs(162)) or (inputs(180));
    layer0_outputs(1944) <= not((inputs(217)) or (inputs(62)));
    layer0_outputs(1945) <= (inputs(156)) xor (inputs(187));
    layer0_outputs(1946) <= (inputs(245)) and not (inputs(7));
    layer0_outputs(1947) <= (inputs(53)) and not (inputs(110));
    layer0_outputs(1948) <= inputs(135);
    layer0_outputs(1949) <= not((inputs(51)) or (inputs(161)));
    layer0_outputs(1950) <= not((inputs(62)) xor (inputs(145)));
    layer0_outputs(1951) <= not(inputs(150));
    layer0_outputs(1952) <= not(inputs(67)) or (inputs(239));
    layer0_outputs(1953) <= (inputs(226)) and not (inputs(237));
    layer0_outputs(1954) <= not(inputs(207));
    layer0_outputs(1955) <= not(inputs(168)) or (inputs(222));
    layer0_outputs(1956) <= not((inputs(211)) or (inputs(249)));
    layer0_outputs(1957) <= (inputs(72)) or (inputs(35));
    layer0_outputs(1958) <= (inputs(218)) and not (inputs(192));
    layer0_outputs(1959) <= (inputs(165)) and not (inputs(153));
    layer0_outputs(1960) <= not(inputs(91));
    layer0_outputs(1961) <= not(inputs(219)) or (inputs(30));
    layer0_outputs(1962) <= not((inputs(217)) or (inputs(130)));
    layer0_outputs(1963) <= '1';
    layer0_outputs(1964) <= (inputs(54)) or (inputs(60));
    layer0_outputs(1965) <= not((inputs(120)) or (inputs(186)));
    layer0_outputs(1966) <= inputs(57);
    layer0_outputs(1967) <= not((inputs(48)) or (inputs(234)));
    layer0_outputs(1968) <= (inputs(149)) and not (inputs(109));
    layer0_outputs(1969) <= not(inputs(247));
    layer0_outputs(1970) <= (inputs(35)) xor (inputs(120));
    layer0_outputs(1971) <= not((inputs(97)) xor (inputs(49)));
    layer0_outputs(1972) <= not(inputs(84));
    layer0_outputs(1973) <= not(inputs(102)) or (inputs(145));
    layer0_outputs(1974) <= not((inputs(174)) or (inputs(90)));
    layer0_outputs(1975) <= not((inputs(168)) or (inputs(42)));
    layer0_outputs(1976) <= inputs(107);
    layer0_outputs(1977) <= not(inputs(153)) or (inputs(103));
    layer0_outputs(1978) <= (inputs(104)) xor (inputs(208));
    layer0_outputs(1979) <= inputs(136);
    layer0_outputs(1980) <= not(inputs(184)) or (inputs(246));
    layer0_outputs(1981) <= not(inputs(146));
    layer0_outputs(1982) <= (inputs(242)) and not (inputs(238));
    layer0_outputs(1983) <= inputs(33);
    layer0_outputs(1984) <= not((inputs(253)) and (inputs(145)));
    layer0_outputs(1985) <= not(inputs(154));
    layer0_outputs(1986) <= not((inputs(193)) and (inputs(192)));
    layer0_outputs(1987) <= not(inputs(116)) or (inputs(180));
    layer0_outputs(1988) <= inputs(219);
    layer0_outputs(1989) <= (inputs(162)) xor (inputs(158));
    layer0_outputs(1990) <= (inputs(126)) xor (inputs(142));
    layer0_outputs(1991) <= (inputs(91)) and not (inputs(74));
    layer0_outputs(1992) <= (inputs(9)) or (inputs(186));
    layer0_outputs(1993) <= (inputs(224)) or (inputs(172));
    layer0_outputs(1994) <= not((inputs(183)) xor (inputs(224)));
    layer0_outputs(1995) <= not(inputs(40)) or (inputs(244));
    layer0_outputs(1996) <= '0';
    layer0_outputs(1997) <= inputs(133);
    layer0_outputs(1998) <= not((inputs(138)) xor (inputs(8)));
    layer0_outputs(1999) <= not(inputs(194)) or (inputs(225));
    layer0_outputs(2000) <= not(inputs(22));
    layer0_outputs(2001) <= (inputs(223)) or (inputs(186));
    layer0_outputs(2002) <= (inputs(135)) and not (inputs(156));
    layer0_outputs(2003) <= (inputs(183)) and not (inputs(91));
    layer0_outputs(2004) <= not(inputs(131)) or (inputs(10));
    layer0_outputs(2005) <= not(inputs(230)) or (inputs(204));
    layer0_outputs(2006) <= (inputs(20)) xor (inputs(101));
    layer0_outputs(2007) <= not((inputs(19)) xor (inputs(216)));
    layer0_outputs(2008) <= not((inputs(176)) and (inputs(19)));
    layer0_outputs(2009) <= not((inputs(22)) or (inputs(148)));
    layer0_outputs(2010) <= not(inputs(204)) or (inputs(29));
    layer0_outputs(2011) <= inputs(106);
    layer0_outputs(2012) <= not((inputs(164)) or (inputs(54)));
    layer0_outputs(2013) <= not((inputs(139)) and (inputs(93)));
    layer0_outputs(2014) <= (inputs(79)) and (inputs(127));
    layer0_outputs(2015) <= not((inputs(49)) xor (inputs(20)));
    layer0_outputs(2016) <= not((inputs(34)) or (inputs(200)));
    layer0_outputs(2017) <= (inputs(123)) xor (inputs(127));
    layer0_outputs(2018) <= not(inputs(37)) or (inputs(231));
    layer0_outputs(2019) <= '1';
    layer0_outputs(2020) <= not(inputs(89));
    layer0_outputs(2021) <= not(inputs(134)) or (inputs(115));
    layer0_outputs(2022) <= (inputs(128)) xor (inputs(133));
    layer0_outputs(2023) <= inputs(74);
    layer0_outputs(2024) <= not((inputs(8)) xor (inputs(203)));
    layer0_outputs(2025) <= inputs(181);
    layer0_outputs(2026) <= (inputs(98)) and not (inputs(18));
    layer0_outputs(2027) <= not((inputs(100)) or (inputs(45)));
    layer0_outputs(2028) <= not((inputs(132)) or (inputs(209)));
    layer0_outputs(2029) <= not(inputs(237));
    layer0_outputs(2030) <= (inputs(23)) or (inputs(84));
    layer0_outputs(2031) <= (inputs(169)) or (inputs(255));
    layer0_outputs(2032) <= (inputs(130)) xor (inputs(127));
    layer0_outputs(2033) <= inputs(56);
    layer0_outputs(2034) <= '0';
    layer0_outputs(2035) <= not((inputs(155)) xor (inputs(182)));
    layer0_outputs(2036) <= not((inputs(106)) or (inputs(131)));
    layer0_outputs(2037) <= not(inputs(40));
    layer0_outputs(2038) <= not(inputs(168)) or (inputs(130));
    layer0_outputs(2039) <= '0';
    layer0_outputs(2040) <= not((inputs(124)) and (inputs(23)));
    layer0_outputs(2041) <= not((inputs(38)) or (inputs(4)));
    layer0_outputs(2042) <= not(inputs(171)) or (inputs(71));
    layer0_outputs(2043) <= inputs(188);
    layer0_outputs(2044) <= (inputs(246)) and not (inputs(88));
    layer0_outputs(2045) <= not(inputs(29));
    layer0_outputs(2046) <= '1';
    layer0_outputs(2047) <= (inputs(251)) and (inputs(160));
    layer0_outputs(2048) <= (inputs(88)) or (inputs(37));
    layer0_outputs(2049) <= (inputs(198)) xor (inputs(40));
    layer0_outputs(2050) <= not((inputs(171)) or (inputs(207)));
    layer0_outputs(2051) <= not((inputs(160)) or (inputs(89)));
    layer0_outputs(2052) <= (inputs(139)) xor (inputs(96));
    layer0_outputs(2053) <= not((inputs(128)) or (inputs(248)));
    layer0_outputs(2054) <= not((inputs(255)) and (inputs(36)));
    layer0_outputs(2055) <= inputs(196);
    layer0_outputs(2056) <= inputs(125);
    layer0_outputs(2057) <= (inputs(255)) and (inputs(218));
    layer0_outputs(2058) <= inputs(148);
    layer0_outputs(2059) <= (inputs(3)) or (inputs(121));
    layer0_outputs(2060) <= (inputs(68)) or (inputs(68));
    layer0_outputs(2061) <= not((inputs(98)) or (inputs(152)));
    layer0_outputs(2062) <= inputs(177);
    layer0_outputs(2063) <= not((inputs(205)) xor (inputs(222)));
    layer0_outputs(2064) <= not(inputs(147));
    layer0_outputs(2065) <= (inputs(42)) xor (inputs(231));
    layer0_outputs(2066) <= not((inputs(39)) or (inputs(245)));
    layer0_outputs(2067) <= inputs(226);
    layer0_outputs(2068) <= (inputs(160)) or (inputs(209));
    layer0_outputs(2069) <= not(inputs(88)) or (inputs(221));
    layer0_outputs(2070) <= (inputs(105)) and not (inputs(240));
    layer0_outputs(2071) <= (inputs(75)) xor (inputs(254));
    layer0_outputs(2072) <= not((inputs(178)) and (inputs(64)));
    layer0_outputs(2073) <= inputs(102);
    layer0_outputs(2074) <= not(inputs(224)) or (inputs(218));
    layer0_outputs(2075) <= (inputs(66)) and not (inputs(22));
    layer0_outputs(2076) <= inputs(73);
    layer0_outputs(2077) <= (inputs(84)) or (inputs(102));
    layer0_outputs(2078) <= inputs(68);
    layer0_outputs(2079) <= (inputs(177)) and (inputs(146));
    layer0_outputs(2080) <= not((inputs(147)) or (inputs(62)));
    layer0_outputs(2081) <= not((inputs(94)) xor (inputs(125)));
    layer0_outputs(2082) <= not(inputs(51));
    layer0_outputs(2083) <= (inputs(116)) and not (inputs(244));
    layer0_outputs(2084) <= (inputs(189)) or (inputs(75));
    layer0_outputs(2085) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(2086) <= inputs(243);
    layer0_outputs(2087) <= (inputs(106)) and not (inputs(125));
    layer0_outputs(2088) <= (inputs(11)) and (inputs(242));
    layer0_outputs(2089) <= not((inputs(129)) xor (inputs(5)));
    layer0_outputs(2090) <= not(inputs(134)) or (inputs(239));
    layer0_outputs(2091) <= inputs(202);
    layer0_outputs(2092) <= (inputs(46)) or (inputs(165));
    layer0_outputs(2093) <= not(inputs(251)) or (inputs(107));
    layer0_outputs(2094) <= (inputs(50)) xor (inputs(118));
    layer0_outputs(2095) <= (inputs(96)) and (inputs(64));
    layer0_outputs(2096) <= not(inputs(193)) or (inputs(246));
    layer0_outputs(2097) <= inputs(153);
    layer0_outputs(2098) <= not((inputs(100)) or (inputs(6)));
    layer0_outputs(2099) <= (inputs(137)) or (inputs(169));
    layer0_outputs(2100) <= not(inputs(167));
    layer0_outputs(2101) <= (inputs(2)) and not (inputs(140));
    layer0_outputs(2102) <= not(inputs(77)) or (inputs(205));
    layer0_outputs(2103) <= not(inputs(102)) or (inputs(57));
    layer0_outputs(2104) <= not(inputs(141));
    layer0_outputs(2105) <= (inputs(186)) and not (inputs(18));
    layer0_outputs(2106) <= not((inputs(63)) xor (inputs(246)));
    layer0_outputs(2107) <= (inputs(223)) or (inputs(148));
    layer0_outputs(2108) <= not((inputs(29)) or (inputs(119)));
    layer0_outputs(2109) <= not(inputs(170));
    layer0_outputs(2110) <= not(inputs(77)) or (inputs(206));
    layer0_outputs(2111) <= not((inputs(127)) or (inputs(36)));
    layer0_outputs(2112) <= not((inputs(23)) or (inputs(82)));
    layer0_outputs(2113) <= (inputs(181)) xor (inputs(10));
    layer0_outputs(2114) <= not(inputs(3));
    layer0_outputs(2115) <= not((inputs(131)) and (inputs(221)));
    layer0_outputs(2116) <= not((inputs(178)) or (inputs(83)));
    layer0_outputs(2117) <= inputs(65);
    layer0_outputs(2118) <= inputs(183);
    layer0_outputs(2119) <= not(inputs(163));
    layer0_outputs(2120) <= inputs(214);
    layer0_outputs(2121) <= not((inputs(68)) xor (inputs(43)));
    layer0_outputs(2122) <= not(inputs(148));
    layer0_outputs(2123) <= (inputs(247)) or (inputs(176));
    layer0_outputs(2124) <= not(inputs(85)) or (inputs(33));
    layer0_outputs(2125) <= (inputs(94)) or (inputs(186));
    layer0_outputs(2126) <= not(inputs(80));
    layer0_outputs(2127) <= not((inputs(130)) or (inputs(168)));
    layer0_outputs(2128) <= not((inputs(34)) or (inputs(181)));
    layer0_outputs(2129) <= (inputs(174)) and (inputs(243));
    layer0_outputs(2130) <= inputs(156);
    layer0_outputs(2131) <= (inputs(114)) and not (inputs(255));
    layer0_outputs(2132) <= (inputs(203)) and not (inputs(70));
    layer0_outputs(2133) <= not((inputs(185)) or (inputs(27)));
    layer0_outputs(2134) <= not(inputs(100));
    layer0_outputs(2135) <= '0';
    layer0_outputs(2136) <= inputs(232);
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= (inputs(9)) or (inputs(109));
    layer0_outputs(2139) <= not(inputs(156));
    layer0_outputs(2140) <= not(inputs(136));
    layer0_outputs(2141) <= not((inputs(112)) and (inputs(176)));
    layer0_outputs(2142) <= (inputs(63)) and (inputs(49));
    layer0_outputs(2143) <= not((inputs(43)) xor (inputs(42)));
    layer0_outputs(2144) <= not(inputs(184));
    layer0_outputs(2145) <= (inputs(139)) xor (inputs(252));
    layer0_outputs(2146) <= not(inputs(33));
    layer0_outputs(2147) <= not((inputs(8)) or (inputs(224)));
    layer0_outputs(2148) <= not(inputs(102)) or (inputs(211));
    layer0_outputs(2149) <= not((inputs(51)) xor (inputs(140)));
    layer0_outputs(2150) <= '1';
    layer0_outputs(2151) <= (inputs(234)) xor (inputs(41));
    layer0_outputs(2152) <= not((inputs(19)) or (inputs(186)));
    layer0_outputs(2153) <= (inputs(99)) xor (inputs(188));
    layer0_outputs(2154) <= (inputs(146)) or (inputs(58));
    layer0_outputs(2155) <= inputs(14);
    layer0_outputs(2156) <= (inputs(118)) or (inputs(174));
    layer0_outputs(2157) <= not((inputs(123)) xor (inputs(119)));
    layer0_outputs(2158) <= (inputs(92)) and (inputs(221));
    layer0_outputs(2159) <= inputs(108);
    layer0_outputs(2160) <= not((inputs(153)) or (inputs(228)));
    layer0_outputs(2161) <= not((inputs(253)) xor (inputs(68)));
    layer0_outputs(2162) <= not((inputs(167)) or (inputs(64)));
    layer0_outputs(2163) <= not((inputs(151)) xor (inputs(221)));
    layer0_outputs(2164) <= (inputs(202)) or (inputs(127));
    layer0_outputs(2165) <= not((inputs(88)) or (inputs(49)));
    layer0_outputs(2166) <= (inputs(236)) and not (inputs(205));
    layer0_outputs(2167) <= not((inputs(164)) or (inputs(125)));
    layer0_outputs(2168) <= '0';
    layer0_outputs(2169) <= not(inputs(108));
    layer0_outputs(2170) <= not((inputs(4)) xor (inputs(156)));
    layer0_outputs(2171) <= (inputs(227)) or (inputs(220));
    layer0_outputs(2172) <= (inputs(215)) xor (inputs(19));
    layer0_outputs(2173) <= not((inputs(65)) or (inputs(139)));
    layer0_outputs(2174) <= not((inputs(237)) xor (inputs(119)));
    layer0_outputs(2175) <= (inputs(142)) xor (inputs(90));
    layer0_outputs(2176) <= (inputs(88)) and not (inputs(62));
    layer0_outputs(2177) <= (inputs(214)) and not (inputs(252));
    layer0_outputs(2178) <= not((inputs(200)) xor (inputs(212)));
    layer0_outputs(2179) <= inputs(226);
    layer0_outputs(2180) <= not(inputs(141));
    layer0_outputs(2181) <= (inputs(137)) xor (inputs(153));
    layer0_outputs(2182) <= inputs(90);
    layer0_outputs(2183) <= not(inputs(72));
    layer0_outputs(2184) <= '1';
    layer0_outputs(2185) <= not((inputs(119)) xor (inputs(80)));
    layer0_outputs(2186) <= (inputs(95)) and not (inputs(249));
    layer0_outputs(2187) <= not((inputs(239)) xor (inputs(112)));
    layer0_outputs(2188) <= inputs(16);
    layer0_outputs(2189) <= inputs(9);
    layer0_outputs(2190) <= inputs(88);
    layer0_outputs(2191) <= (inputs(239)) and not (inputs(62));
    layer0_outputs(2192) <= not(inputs(19)) or (inputs(191));
    layer0_outputs(2193) <= (inputs(130)) and not (inputs(241));
    layer0_outputs(2194) <= (inputs(215)) or (inputs(124));
    layer0_outputs(2195) <= not(inputs(29));
    layer0_outputs(2196) <= not(inputs(217));
    layer0_outputs(2197) <= not(inputs(165));
    layer0_outputs(2198) <= (inputs(85)) and not (inputs(127));
    layer0_outputs(2199) <= not((inputs(70)) or (inputs(231)));
    layer0_outputs(2200) <= (inputs(131)) or (inputs(245));
    layer0_outputs(2201) <= not((inputs(214)) or (inputs(215)));
    layer0_outputs(2202) <= inputs(31);
    layer0_outputs(2203) <= not((inputs(111)) or (inputs(86)));
    layer0_outputs(2204) <= (inputs(31)) and (inputs(9));
    layer0_outputs(2205) <= (inputs(172)) xor (inputs(188));
    layer0_outputs(2206) <= not((inputs(148)) xor (inputs(181)));
    layer0_outputs(2207) <= not(inputs(23)) or (inputs(189));
    layer0_outputs(2208) <= (inputs(181)) and not (inputs(243));
    layer0_outputs(2209) <= not((inputs(93)) xor (inputs(4)));
    layer0_outputs(2210) <= not(inputs(59)) or (inputs(192));
    layer0_outputs(2211) <= (inputs(47)) xor (inputs(86));
    layer0_outputs(2212) <= not((inputs(211)) xor (inputs(13)));
    layer0_outputs(2213) <= (inputs(249)) and not (inputs(19));
    layer0_outputs(2214) <= (inputs(125)) or (inputs(196));
    layer0_outputs(2215) <= (inputs(255)) and (inputs(253));
    layer0_outputs(2216) <= (inputs(242)) and not (inputs(177));
    layer0_outputs(2217) <= not(inputs(234)) or (inputs(221));
    layer0_outputs(2218) <= not((inputs(164)) xor (inputs(153)));
    layer0_outputs(2219) <= (inputs(113)) xor (inputs(138));
    layer0_outputs(2220) <= (inputs(86)) and not (inputs(158));
    layer0_outputs(2221) <= (inputs(193)) or (inputs(227));
    layer0_outputs(2222) <= '1';
    layer0_outputs(2223) <= (inputs(99)) and not (inputs(139));
    layer0_outputs(2224) <= inputs(85);
    layer0_outputs(2225) <= not(inputs(196));
    layer0_outputs(2226) <= not(inputs(179)) or (inputs(40));
    layer0_outputs(2227) <= inputs(71);
    layer0_outputs(2228) <= not(inputs(223)) or (inputs(129));
    layer0_outputs(2229) <= (inputs(220)) and (inputs(178));
    layer0_outputs(2230) <= not((inputs(87)) xor (inputs(129)));
    layer0_outputs(2231) <= not(inputs(98)) or (inputs(31));
    layer0_outputs(2232) <= not(inputs(72)) or (inputs(193));
    layer0_outputs(2233) <= not(inputs(117));
    layer0_outputs(2234) <= not((inputs(231)) or (inputs(123)));
    layer0_outputs(2235) <= not((inputs(44)) or (inputs(99)));
    layer0_outputs(2236) <= not((inputs(254)) or (inputs(97)));
    layer0_outputs(2237) <= (inputs(127)) xor (inputs(57));
    layer0_outputs(2238) <= not(inputs(138)) or (inputs(253));
    layer0_outputs(2239) <= (inputs(104)) xor (inputs(53));
    layer0_outputs(2240) <= not(inputs(119));
    layer0_outputs(2241) <= (inputs(170)) or (inputs(213));
    layer0_outputs(2242) <= not((inputs(11)) or (inputs(209)));
    layer0_outputs(2243) <= (inputs(123)) and not (inputs(39));
    layer0_outputs(2244) <= (inputs(76)) or (inputs(44));
    layer0_outputs(2245) <= (inputs(14)) or (inputs(139));
    layer0_outputs(2246) <= (inputs(114)) or (inputs(234));
    layer0_outputs(2247) <= not(inputs(151)) or (inputs(81));
    layer0_outputs(2248) <= (inputs(60)) and not (inputs(244));
    layer0_outputs(2249) <= (inputs(76)) and not (inputs(224));
    layer0_outputs(2250) <= (inputs(201)) and not (inputs(13));
    layer0_outputs(2251) <= inputs(230);
    layer0_outputs(2252) <= (inputs(195)) or (inputs(203));
    layer0_outputs(2253) <= not(inputs(164));
    layer0_outputs(2254) <= not((inputs(151)) xor (inputs(221)));
    layer0_outputs(2255) <= (inputs(58)) xor (inputs(224));
    layer0_outputs(2256) <= '1';
    layer0_outputs(2257) <= (inputs(126)) xor (inputs(35));
    layer0_outputs(2258) <= not((inputs(124)) or (inputs(190)));
    layer0_outputs(2259) <= not((inputs(5)) xor (inputs(219)));
    layer0_outputs(2260) <= not(inputs(56));
    layer0_outputs(2261) <= (inputs(21)) or (inputs(171));
    layer0_outputs(2262) <= not(inputs(115));
    layer0_outputs(2263) <= not((inputs(24)) or (inputs(181)));
    layer0_outputs(2264) <= not(inputs(114));
    layer0_outputs(2265) <= not(inputs(138)) or (inputs(109));
    layer0_outputs(2266) <= inputs(10);
    layer0_outputs(2267) <= (inputs(130)) or (inputs(9));
    layer0_outputs(2268) <= inputs(160);
    layer0_outputs(2269) <= (inputs(253)) or (inputs(234));
    layer0_outputs(2270) <= inputs(88);
    layer0_outputs(2271) <= (inputs(220)) and not (inputs(19));
    layer0_outputs(2272) <= not(inputs(71));
    layer0_outputs(2273) <= (inputs(197)) xor (inputs(236));
    layer0_outputs(2274) <= inputs(99);
    layer0_outputs(2275) <= not((inputs(174)) or (inputs(181)));
    layer0_outputs(2276) <= not((inputs(160)) or (inputs(183)));
    layer0_outputs(2277) <= not(inputs(160)) or (inputs(27));
    layer0_outputs(2278) <= not(inputs(28)) or (inputs(178));
    layer0_outputs(2279) <= not((inputs(65)) and (inputs(143)));
    layer0_outputs(2280) <= inputs(82);
    layer0_outputs(2281) <= '0';
    layer0_outputs(2282) <= (inputs(176)) and (inputs(219));
    layer0_outputs(2283) <= inputs(118);
    layer0_outputs(2284) <= (inputs(22)) and not (inputs(209));
    layer0_outputs(2285) <= (inputs(199)) or (inputs(145));
    layer0_outputs(2286) <= not((inputs(54)) or (inputs(202)));
    layer0_outputs(2287) <= not(inputs(36));
    layer0_outputs(2288) <= (inputs(205)) xor (inputs(119));
    layer0_outputs(2289) <= not(inputs(6));
    layer0_outputs(2290) <= not(inputs(69));
    layer0_outputs(2291) <= (inputs(111)) and (inputs(7));
    layer0_outputs(2292) <= (inputs(195)) and not (inputs(237));
    layer0_outputs(2293) <= not(inputs(40));
    layer0_outputs(2294) <= inputs(170);
    layer0_outputs(2295) <= not((inputs(127)) or (inputs(32)));
    layer0_outputs(2296) <= not((inputs(157)) or (inputs(40)));
    layer0_outputs(2297) <= not(inputs(106));
    layer0_outputs(2298) <= (inputs(217)) and not (inputs(160));
    layer0_outputs(2299) <= not(inputs(42));
    layer0_outputs(2300) <= (inputs(85)) or (inputs(7));
    layer0_outputs(2301) <= (inputs(247)) or (inputs(204));
    layer0_outputs(2302) <= inputs(150);
    layer0_outputs(2303) <= not((inputs(190)) or (inputs(121)));
    layer0_outputs(2304) <= not(inputs(147));
    layer0_outputs(2305) <= not((inputs(6)) xor (inputs(162)));
    layer0_outputs(2306) <= (inputs(0)) and not (inputs(31));
    layer0_outputs(2307) <= not(inputs(150)) or (inputs(48));
    layer0_outputs(2308) <= inputs(186);
    layer0_outputs(2309) <= (inputs(137)) and not (inputs(222));
    layer0_outputs(2310) <= (inputs(173)) xor (inputs(194));
    layer0_outputs(2311) <= (inputs(148)) and (inputs(63));
    layer0_outputs(2312) <= (inputs(138)) xor (inputs(12));
    layer0_outputs(2313) <= inputs(214);
    layer0_outputs(2314) <= not(inputs(233)) or (inputs(13));
    layer0_outputs(2315) <= not(inputs(155)) or (inputs(208));
    layer0_outputs(2316) <= (inputs(54)) or (inputs(21));
    layer0_outputs(2317) <= not(inputs(167)) or (inputs(229));
    layer0_outputs(2318) <= not(inputs(212)) or (inputs(28));
    layer0_outputs(2319) <= not(inputs(191)) or (inputs(34));
    layer0_outputs(2320) <= not(inputs(68));
    layer0_outputs(2321) <= not(inputs(70));
    layer0_outputs(2322) <= not(inputs(149)) or (inputs(18));
    layer0_outputs(2323) <= not(inputs(185));
    layer0_outputs(2324) <= not(inputs(71)) or (inputs(30));
    layer0_outputs(2325) <= not((inputs(252)) and (inputs(112)));
    layer0_outputs(2326) <= not((inputs(4)) xor (inputs(48)));
    layer0_outputs(2327) <= (inputs(124)) and not (inputs(67));
    layer0_outputs(2328) <= (inputs(157)) xor (inputs(173));
    layer0_outputs(2329) <= not((inputs(39)) or (inputs(248)));
    layer0_outputs(2330) <= (inputs(25)) or (inputs(81));
    layer0_outputs(2331) <= (inputs(39)) and not (inputs(5));
    layer0_outputs(2332) <= not((inputs(244)) and (inputs(75)));
    layer0_outputs(2333) <= not(inputs(85)) or (inputs(177));
    layer0_outputs(2334) <= not(inputs(105)) or (inputs(225));
    layer0_outputs(2335) <= '1';
    layer0_outputs(2336) <= (inputs(86)) and (inputs(86));
    layer0_outputs(2337) <= not((inputs(199)) xor (inputs(128)));
    layer0_outputs(2338) <= not(inputs(57));
    layer0_outputs(2339) <= not((inputs(12)) or (inputs(135)));
    layer0_outputs(2340) <= not((inputs(67)) or (inputs(41)));
    layer0_outputs(2341) <= not((inputs(47)) xor (inputs(60)));
    layer0_outputs(2342) <= (inputs(230)) and not (inputs(187));
    layer0_outputs(2343) <= (inputs(5)) and not (inputs(19));
    layer0_outputs(2344) <= not((inputs(69)) or (inputs(22)));
    layer0_outputs(2345) <= not(inputs(85));
    layer0_outputs(2346) <= (inputs(103)) and not (inputs(242));
    layer0_outputs(2347) <= (inputs(79)) and not (inputs(82));
    layer0_outputs(2348) <= inputs(184);
    layer0_outputs(2349) <= inputs(101);
    layer0_outputs(2350) <= '0';
    layer0_outputs(2351) <= not((inputs(33)) xor (inputs(92)));
    layer0_outputs(2352) <= not((inputs(233)) xor (inputs(166)));
    layer0_outputs(2353) <= (inputs(87)) or (inputs(137));
    layer0_outputs(2354) <= not(inputs(102)) or (inputs(178));
    layer0_outputs(2355) <= not(inputs(123)) or (inputs(35));
    layer0_outputs(2356) <= not((inputs(113)) or (inputs(79)));
    layer0_outputs(2357) <= inputs(104);
    layer0_outputs(2358) <= not((inputs(118)) or (inputs(79)));
    layer0_outputs(2359) <= not(inputs(180));
    layer0_outputs(2360) <= not(inputs(96)) or (inputs(246));
    layer0_outputs(2361) <= inputs(165);
    layer0_outputs(2362) <= (inputs(129)) and not (inputs(125));
    layer0_outputs(2363) <= not((inputs(81)) xor (inputs(194)));
    layer0_outputs(2364) <= (inputs(146)) and (inputs(24));
    layer0_outputs(2365) <= (inputs(220)) or (inputs(193));
    layer0_outputs(2366) <= inputs(171);
    layer0_outputs(2367) <= inputs(218);
    layer0_outputs(2368) <= (inputs(209)) and not (inputs(125));
    layer0_outputs(2369) <= (inputs(242)) or (inputs(169));
    layer0_outputs(2370) <= (inputs(185)) and not (inputs(8));
    layer0_outputs(2371) <= (inputs(97)) and not (inputs(9));
    layer0_outputs(2372) <= not((inputs(34)) and (inputs(11)));
    layer0_outputs(2373) <= (inputs(26)) and not (inputs(114));
    layer0_outputs(2374) <= not(inputs(74));
    layer0_outputs(2375) <= not((inputs(151)) xor (inputs(255)));
    layer0_outputs(2376) <= not((inputs(118)) or (inputs(126)));
    layer0_outputs(2377) <= (inputs(22)) xor (inputs(101));
    layer0_outputs(2378) <= not(inputs(105)) or (inputs(103));
    layer0_outputs(2379) <= not(inputs(111));
    layer0_outputs(2380) <= not(inputs(63)) or (inputs(2));
    layer0_outputs(2381) <= not((inputs(34)) xor (inputs(151)));
    layer0_outputs(2382) <= not((inputs(110)) and (inputs(81)));
    layer0_outputs(2383) <= not(inputs(136)) or (inputs(173));
    layer0_outputs(2384) <= (inputs(190)) xor (inputs(124));
    layer0_outputs(2385) <= not(inputs(164)) or (inputs(220));
    layer0_outputs(2386) <= (inputs(102)) or (inputs(166));
    layer0_outputs(2387) <= (inputs(32)) xor (inputs(150));
    layer0_outputs(2388) <= (inputs(104)) or (inputs(230));
    layer0_outputs(2389) <= (inputs(162)) or (inputs(45));
    layer0_outputs(2390) <= (inputs(90)) or (inputs(228));
    layer0_outputs(2391) <= not(inputs(164)) or (inputs(254));
    layer0_outputs(2392) <= not((inputs(229)) or (inputs(230)));
    layer0_outputs(2393) <= not((inputs(71)) or (inputs(241)));
    layer0_outputs(2394) <= inputs(120);
    layer0_outputs(2395) <= '1';
    layer0_outputs(2396) <= not(inputs(185)) or (inputs(168));
    layer0_outputs(2397) <= not(inputs(232)) or (inputs(46));
    layer0_outputs(2398) <= not((inputs(221)) or (inputs(202)));
    layer0_outputs(2399) <= (inputs(50)) or (inputs(221));
    layer0_outputs(2400) <= inputs(131);
    layer0_outputs(2401) <= (inputs(177)) and not (inputs(51));
    layer0_outputs(2402) <= inputs(215);
    layer0_outputs(2403) <= inputs(88);
    layer0_outputs(2404) <= '0';
    layer0_outputs(2405) <= (inputs(99)) and not (inputs(62));
    layer0_outputs(2406) <= '0';
    layer0_outputs(2407) <= not(inputs(164)) or (inputs(30));
    layer0_outputs(2408) <= (inputs(236)) or (inputs(96));
    layer0_outputs(2409) <= inputs(123);
    layer0_outputs(2410) <= (inputs(187)) and not (inputs(238));
    layer0_outputs(2411) <= not((inputs(150)) or (inputs(40)));
    layer0_outputs(2412) <= not((inputs(108)) or (inputs(250)));
    layer0_outputs(2413) <= (inputs(233)) or (inputs(15));
    layer0_outputs(2414) <= inputs(184);
    layer0_outputs(2415) <= not(inputs(236));
    layer0_outputs(2416) <= not(inputs(88));
    layer0_outputs(2417) <= not((inputs(186)) xor (inputs(224)));
    layer0_outputs(2418) <= not(inputs(229));
    layer0_outputs(2419) <= inputs(4);
    layer0_outputs(2420) <= (inputs(189)) or (inputs(38));
    layer0_outputs(2421) <= inputs(232);
    layer0_outputs(2422) <= (inputs(0)) or (inputs(116));
    layer0_outputs(2423) <= (inputs(198)) and not (inputs(9));
    layer0_outputs(2424) <= not((inputs(253)) and (inputs(110)));
    layer0_outputs(2425) <= (inputs(23)) xor (inputs(105));
    layer0_outputs(2426) <= not(inputs(157));
    layer0_outputs(2427) <= not((inputs(188)) or (inputs(254)));
    layer0_outputs(2428) <= (inputs(24)) and not (inputs(238));
    layer0_outputs(2429) <= (inputs(40)) or (inputs(151));
    layer0_outputs(2430) <= not(inputs(89)) or (inputs(5));
    layer0_outputs(2431) <= not(inputs(126));
    layer0_outputs(2432) <= (inputs(223)) and not (inputs(51));
    layer0_outputs(2433) <= not((inputs(16)) xor (inputs(167)));
    layer0_outputs(2434) <= not(inputs(229));
    layer0_outputs(2435) <= (inputs(247)) and not (inputs(61));
    layer0_outputs(2436) <= not((inputs(51)) xor (inputs(185)));
    layer0_outputs(2437) <= not((inputs(203)) or (inputs(76)));
    layer0_outputs(2438) <= (inputs(219)) xor (inputs(187));
    layer0_outputs(2439) <= not(inputs(0)) or (inputs(142));
    layer0_outputs(2440) <= not((inputs(86)) or (inputs(41)));
    layer0_outputs(2441) <= (inputs(194)) xor (inputs(6));
    layer0_outputs(2442) <= (inputs(62)) or (inputs(106));
    layer0_outputs(2443) <= not(inputs(120));
    layer0_outputs(2444) <= (inputs(157)) and not (inputs(130));
    layer0_outputs(2445) <= not(inputs(16));
    layer0_outputs(2446) <= not(inputs(106));
    layer0_outputs(2447) <= inputs(196);
    layer0_outputs(2448) <= not((inputs(37)) xor (inputs(3)));
    layer0_outputs(2449) <= not(inputs(23));
    layer0_outputs(2450) <= not((inputs(120)) or (inputs(162)));
    layer0_outputs(2451) <= not((inputs(146)) or (inputs(52)));
    layer0_outputs(2452) <= not((inputs(134)) xor (inputs(50)));
    layer0_outputs(2453) <= (inputs(69)) or (inputs(78));
    layer0_outputs(2454) <= inputs(85);
    layer0_outputs(2455) <= not(inputs(86));
    layer0_outputs(2456) <= inputs(212);
    layer0_outputs(2457) <= (inputs(204)) or (inputs(135));
    layer0_outputs(2458) <= (inputs(93)) and not (inputs(93));
    layer0_outputs(2459) <= not(inputs(56)) or (inputs(94));
    layer0_outputs(2460) <= not(inputs(30));
    layer0_outputs(2461) <= inputs(247);
    layer0_outputs(2462) <= not(inputs(215)) or (inputs(225));
    layer0_outputs(2463) <= not((inputs(157)) xor (inputs(133)));
    layer0_outputs(2464) <= not(inputs(40)) or (inputs(244));
    layer0_outputs(2465) <= not((inputs(192)) or (inputs(230)));
    layer0_outputs(2466) <= (inputs(91)) and not (inputs(131));
    layer0_outputs(2467) <= not(inputs(140)) or (inputs(5));
    layer0_outputs(2468) <= '0';
    layer0_outputs(2469) <= (inputs(128)) xor (inputs(19));
    layer0_outputs(2470) <= not((inputs(146)) xor (inputs(60)));
    layer0_outputs(2471) <= not(inputs(214));
    layer0_outputs(2472) <= not((inputs(189)) xor (inputs(231)));
    layer0_outputs(2473) <= not((inputs(157)) or (inputs(194)));
    layer0_outputs(2474) <= not((inputs(164)) xor (inputs(175)));
    layer0_outputs(2475) <= not(inputs(151)) or (inputs(51));
    layer0_outputs(2476) <= (inputs(219)) and (inputs(225));
    layer0_outputs(2477) <= (inputs(49)) and (inputs(16));
    layer0_outputs(2478) <= inputs(115);
    layer0_outputs(2479) <= (inputs(139)) xor (inputs(31));
    layer0_outputs(2480) <= (inputs(127)) xor (inputs(64));
    layer0_outputs(2481) <= (inputs(90)) and not (inputs(28));
    layer0_outputs(2482) <= '0';
    layer0_outputs(2483) <= inputs(23);
    layer0_outputs(2484) <= (inputs(137)) and not (inputs(56));
    layer0_outputs(2485) <= (inputs(120)) or (inputs(53));
    layer0_outputs(2486) <= not((inputs(113)) xor (inputs(85)));
    layer0_outputs(2487) <= inputs(115);
    layer0_outputs(2488) <= (inputs(120)) and not (inputs(29));
    layer0_outputs(2489) <= not((inputs(109)) xor (inputs(15)));
    layer0_outputs(2490) <= inputs(89);
    layer0_outputs(2491) <= inputs(139);
    layer0_outputs(2492) <= (inputs(53)) or (inputs(83));
    layer0_outputs(2493) <= not(inputs(39)) or (inputs(27));
    layer0_outputs(2494) <= not((inputs(196)) xor (inputs(82)));
    layer0_outputs(2495) <= not((inputs(235)) or (inputs(150)));
    layer0_outputs(2496) <= (inputs(240)) and not (inputs(192));
    layer0_outputs(2497) <= inputs(41);
    layer0_outputs(2498) <= (inputs(57)) and not (inputs(93));
    layer0_outputs(2499) <= (inputs(13)) xor (inputs(199));
    layer0_outputs(2500) <= (inputs(85)) or (inputs(13));
    layer0_outputs(2501) <= (inputs(87)) and not (inputs(71));
    layer0_outputs(2502) <= (inputs(21)) or (inputs(33));
    layer0_outputs(2503) <= not((inputs(239)) or (inputs(93)));
    layer0_outputs(2504) <= not(inputs(193)) or (inputs(70));
    layer0_outputs(2505) <= (inputs(73)) and not (inputs(47));
    layer0_outputs(2506) <= (inputs(26)) and (inputs(161));
    layer0_outputs(2507) <= not(inputs(74)) or (inputs(132));
    layer0_outputs(2508) <= (inputs(106)) and not (inputs(143));
    layer0_outputs(2509) <= inputs(19);
    layer0_outputs(2510) <= (inputs(128)) and not (inputs(0));
    layer0_outputs(2511) <= not((inputs(237)) and (inputs(236)));
    layer0_outputs(2512) <= inputs(54);
    layer0_outputs(2513) <= (inputs(95)) or (inputs(201));
    layer0_outputs(2514) <= (inputs(24)) xor (inputs(252));
    layer0_outputs(2515) <= not((inputs(47)) or (inputs(20)));
    layer0_outputs(2516) <= not((inputs(55)) xor (inputs(64)));
    layer0_outputs(2517) <= (inputs(238)) xor (inputs(132));
    layer0_outputs(2518) <= '1';
    layer0_outputs(2519) <= (inputs(133)) or (inputs(159));
    layer0_outputs(2520) <= (inputs(175)) xor (inputs(47));
    layer0_outputs(2521) <= not((inputs(109)) or (inputs(67)));
    layer0_outputs(2522) <= not((inputs(189)) xor (inputs(242)));
    layer0_outputs(2523) <= inputs(230);
    layer0_outputs(2524) <= (inputs(233)) xor (inputs(39));
    layer0_outputs(2525) <= not(inputs(220)) or (inputs(110));
    layer0_outputs(2526) <= (inputs(137)) xor (inputs(237));
    layer0_outputs(2527) <= not(inputs(244)) or (inputs(115));
    layer0_outputs(2528) <= (inputs(209)) or (inputs(154));
    layer0_outputs(2529) <= (inputs(220)) or (inputs(153));
    layer0_outputs(2530) <= not(inputs(120));
    layer0_outputs(2531) <= not(inputs(141)) or (inputs(248));
    layer0_outputs(2532) <= inputs(49);
    layer0_outputs(2533) <= (inputs(103)) and not (inputs(10));
    layer0_outputs(2534) <= '0';
    layer0_outputs(2535) <= not((inputs(132)) xor (inputs(251)));
    layer0_outputs(2536) <= not((inputs(139)) or (inputs(186)));
    layer0_outputs(2537) <= not(inputs(41));
    layer0_outputs(2538) <= not((inputs(231)) or (inputs(134)));
    layer0_outputs(2539) <= (inputs(231)) and not (inputs(253));
    layer0_outputs(2540) <= (inputs(20)) or (inputs(71));
    layer0_outputs(2541) <= (inputs(179)) or (inputs(209));
    layer0_outputs(2542) <= not((inputs(163)) or (inputs(203)));
    layer0_outputs(2543) <= (inputs(252)) and not (inputs(52));
    layer0_outputs(2544) <= not(inputs(131)) or (inputs(190));
    layer0_outputs(2545) <= (inputs(73)) or (inputs(232));
    layer0_outputs(2546) <= not(inputs(104)) or (inputs(81));
    layer0_outputs(2547) <= inputs(228);
    layer0_outputs(2548) <= not(inputs(54)) or (inputs(26));
    layer0_outputs(2549) <= not(inputs(73));
    layer0_outputs(2550) <= inputs(135);
    layer0_outputs(2551) <= not(inputs(107));
    layer0_outputs(2552) <= (inputs(55)) xor (inputs(0));
    layer0_outputs(2553) <= not(inputs(59));
    layer0_outputs(2554) <= (inputs(199)) xor (inputs(16));
    layer0_outputs(2555) <= (inputs(236)) and not (inputs(21));
    layer0_outputs(2556) <= inputs(173);
    layer0_outputs(2557) <= inputs(187);
    layer0_outputs(2558) <= (inputs(61)) and not (inputs(12));
    layer0_outputs(2559) <= (inputs(127)) and (inputs(240));
    layer0_outputs(2560) <= (inputs(102)) or (inputs(232));
    layer0_outputs(2561) <= not((inputs(175)) xor (inputs(88)));
    layer0_outputs(2562) <= (inputs(232)) and not (inputs(17));
    layer0_outputs(2563) <= not((inputs(85)) xor (inputs(252)));
    layer0_outputs(2564) <= not(inputs(157)) or (inputs(66));
    layer0_outputs(2565) <= not(inputs(125));
    layer0_outputs(2566) <= (inputs(39)) xor (inputs(44));
    layer0_outputs(2567) <= (inputs(189)) and not (inputs(238));
    layer0_outputs(2568) <= not(inputs(123)) or (inputs(178));
    layer0_outputs(2569) <= (inputs(216)) or (inputs(199));
    layer0_outputs(2570) <= not((inputs(66)) or (inputs(33)));
    layer0_outputs(2571) <= not(inputs(185)) or (inputs(207));
    layer0_outputs(2572) <= not((inputs(93)) or (inputs(229)));
    layer0_outputs(2573) <= (inputs(186)) and not (inputs(47));
    layer0_outputs(2574) <= not(inputs(180));
    layer0_outputs(2575) <= inputs(235);
    layer0_outputs(2576) <= inputs(62);
    layer0_outputs(2577) <= not((inputs(223)) and (inputs(184)));
    layer0_outputs(2578) <= not(inputs(106)) or (inputs(42));
    layer0_outputs(2579) <= not(inputs(55));
    layer0_outputs(2580) <= not(inputs(125));
    layer0_outputs(2581) <= not(inputs(93));
    layer0_outputs(2582) <= (inputs(78)) and not (inputs(194));
    layer0_outputs(2583) <= (inputs(214)) and not (inputs(111));
    layer0_outputs(2584) <= not((inputs(141)) or (inputs(169)));
    layer0_outputs(2585) <= not(inputs(106));
    layer0_outputs(2586) <= inputs(215);
    layer0_outputs(2587) <= '0';
    layer0_outputs(2588) <= not(inputs(133)) or (inputs(32));
    layer0_outputs(2589) <= not((inputs(23)) xor (inputs(147)));
    layer0_outputs(2590) <= not((inputs(191)) xor (inputs(93)));
    layer0_outputs(2591) <= '0';
    layer0_outputs(2592) <= not(inputs(41));
    layer0_outputs(2593) <= (inputs(168)) and not (inputs(172));
    layer0_outputs(2594) <= not((inputs(207)) and (inputs(219)));
    layer0_outputs(2595) <= (inputs(76)) and not (inputs(188));
    layer0_outputs(2596) <= not(inputs(151)) or (inputs(232));
    layer0_outputs(2597) <= '0';
    layer0_outputs(2598) <= not(inputs(180));
    layer0_outputs(2599) <= (inputs(152)) and not (inputs(62));
    layer0_outputs(2600) <= not(inputs(107)) or (inputs(26));
    layer0_outputs(2601) <= '0';
    layer0_outputs(2602) <= (inputs(103)) and not (inputs(231));
    layer0_outputs(2603) <= (inputs(86)) or (inputs(142));
    layer0_outputs(2604) <= not((inputs(230)) xor (inputs(136)));
    layer0_outputs(2605) <= not(inputs(21));
    layer0_outputs(2606) <= (inputs(62)) or (inputs(132));
    layer0_outputs(2607) <= not(inputs(109)) or (inputs(78));
    layer0_outputs(2608) <= (inputs(127)) or (inputs(219));
    layer0_outputs(2609) <= '1';
    layer0_outputs(2610) <= not(inputs(83));
    layer0_outputs(2611) <= (inputs(252)) or (inputs(142));
    layer0_outputs(2612) <= (inputs(166)) xor (inputs(224));
    layer0_outputs(2613) <= not((inputs(155)) xor (inputs(29)));
    layer0_outputs(2614) <= (inputs(181)) or (inputs(129));
    layer0_outputs(2615) <= not((inputs(20)) xor (inputs(105)));
    layer0_outputs(2616) <= not((inputs(207)) xor (inputs(110)));
    layer0_outputs(2617) <= (inputs(162)) or (inputs(115));
    layer0_outputs(2618) <= not((inputs(2)) xor (inputs(201)));
    layer0_outputs(2619) <= not(inputs(212)) or (inputs(4));
    layer0_outputs(2620) <= (inputs(73)) and not (inputs(200));
    layer0_outputs(2621) <= (inputs(175)) or (inputs(32));
    layer0_outputs(2622) <= not((inputs(22)) or (inputs(104)));
    layer0_outputs(2623) <= '0';
    layer0_outputs(2624) <= not((inputs(121)) xor (inputs(65)));
    layer0_outputs(2625) <= (inputs(80)) and (inputs(54));
    layer0_outputs(2626) <= '0';
    layer0_outputs(2627) <= not(inputs(179)) or (inputs(96));
    layer0_outputs(2628) <= inputs(75);
    layer0_outputs(2629) <= (inputs(225)) xor (inputs(24));
    layer0_outputs(2630) <= (inputs(38)) and not (inputs(96));
    layer0_outputs(2631) <= (inputs(209)) and not (inputs(66));
    layer0_outputs(2632) <= (inputs(149)) and not (inputs(2));
    layer0_outputs(2633) <= not((inputs(54)) or (inputs(28)));
    layer0_outputs(2634) <= (inputs(195)) xor (inputs(126));
    layer0_outputs(2635) <= not((inputs(50)) and (inputs(93)));
    layer0_outputs(2636) <= not(inputs(214)) or (inputs(133));
    layer0_outputs(2637) <= (inputs(44)) or (inputs(2));
    layer0_outputs(2638) <= not((inputs(189)) xor (inputs(157)));
    layer0_outputs(2639) <= not(inputs(99)) or (inputs(237));
    layer0_outputs(2640) <= not(inputs(133)) or (inputs(177));
    layer0_outputs(2641) <= (inputs(223)) xor (inputs(184));
    layer0_outputs(2642) <= not((inputs(161)) xor (inputs(161)));
    layer0_outputs(2643) <= (inputs(96)) or (inputs(8));
    layer0_outputs(2644) <= (inputs(252)) xor (inputs(201));
    layer0_outputs(2645) <= (inputs(173)) and (inputs(161));
    layer0_outputs(2646) <= not((inputs(77)) xor (inputs(54)));
    layer0_outputs(2647) <= not(inputs(87));
    layer0_outputs(2648) <= not((inputs(111)) or (inputs(4)));
    layer0_outputs(2649) <= (inputs(84)) or (inputs(78));
    layer0_outputs(2650) <= not(inputs(197));
    layer0_outputs(2651) <= not((inputs(167)) or (inputs(253)));
    layer0_outputs(2652) <= (inputs(76)) xor (inputs(202));
    layer0_outputs(2653) <= not(inputs(131)) or (inputs(60));
    layer0_outputs(2654) <= (inputs(115)) and not (inputs(22));
    layer0_outputs(2655) <= not((inputs(56)) or (inputs(219)));
    layer0_outputs(2656) <= '1';
    layer0_outputs(2657) <= (inputs(186)) and not (inputs(143));
    layer0_outputs(2658) <= not((inputs(172)) and (inputs(160)));
    layer0_outputs(2659) <= inputs(193);
    layer0_outputs(2660) <= (inputs(138)) and not (inputs(104));
    layer0_outputs(2661) <= not((inputs(83)) and (inputs(160)));
    layer0_outputs(2662) <= not(inputs(83));
    layer0_outputs(2663) <= (inputs(123)) and not (inputs(50));
    layer0_outputs(2664) <= not(inputs(61));
    layer0_outputs(2665) <= not((inputs(255)) or (inputs(50)));
    layer0_outputs(2666) <= not(inputs(220));
    layer0_outputs(2667) <= not(inputs(135)) or (inputs(45));
    layer0_outputs(2668) <= inputs(2);
    layer0_outputs(2669) <= not(inputs(182)) or (inputs(223));
    layer0_outputs(2670) <= (inputs(123)) and not (inputs(110));
    layer0_outputs(2671) <= not((inputs(203)) or (inputs(58)));
    layer0_outputs(2672) <= (inputs(61)) xor (inputs(175));
    layer0_outputs(2673) <= not((inputs(134)) xor (inputs(36)));
    layer0_outputs(2674) <= not((inputs(229)) xor (inputs(31)));
    layer0_outputs(2675) <= not((inputs(147)) or (inputs(229)));
    layer0_outputs(2676) <= not(inputs(225)) or (inputs(14));
    layer0_outputs(2677) <= (inputs(221)) or (inputs(183));
    layer0_outputs(2678) <= not((inputs(51)) xor (inputs(178)));
    layer0_outputs(2679) <= not((inputs(137)) or (inputs(27)));
    layer0_outputs(2680) <= inputs(21);
    layer0_outputs(2681) <= (inputs(175)) or (inputs(24));
    layer0_outputs(2682) <= '1';
    layer0_outputs(2683) <= not(inputs(126));
    layer0_outputs(2684) <= not((inputs(28)) xor (inputs(146)));
    layer0_outputs(2685) <= (inputs(252)) xor (inputs(166));
    layer0_outputs(2686) <= not(inputs(97)) or (inputs(254));
    layer0_outputs(2687) <= not(inputs(138)) or (inputs(9));
    layer0_outputs(2688) <= inputs(125);
    layer0_outputs(2689) <= inputs(121);
    layer0_outputs(2690) <= not(inputs(76)) or (inputs(112));
    layer0_outputs(2691) <= (inputs(186)) xor (inputs(225));
    layer0_outputs(2692) <= (inputs(94)) or (inputs(164));
    layer0_outputs(2693) <= (inputs(108)) and not (inputs(77));
    layer0_outputs(2694) <= '0';
    layer0_outputs(2695) <= inputs(150);
    layer0_outputs(2696) <= (inputs(198)) or (inputs(151));
    layer0_outputs(2697) <= not(inputs(120)) or (inputs(82));
    layer0_outputs(2698) <= inputs(93);
    layer0_outputs(2699) <= not((inputs(110)) xor (inputs(220)));
    layer0_outputs(2700) <= not((inputs(163)) xor (inputs(251)));
    layer0_outputs(2701) <= not(inputs(188)) or (inputs(169));
    layer0_outputs(2702) <= not((inputs(189)) or (inputs(7)));
    layer0_outputs(2703) <= (inputs(18)) xor (inputs(187));
    layer0_outputs(2704) <= not(inputs(25));
    layer0_outputs(2705) <= inputs(165);
    layer0_outputs(2706) <= '1';
    layer0_outputs(2707) <= not(inputs(173));
    layer0_outputs(2708) <= (inputs(124)) or (inputs(107));
    layer0_outputs(2709) <= not((inputs(102)) xor (inputs(235)));
    layer0_outputs(2710) <= not(inputs(137));
    layer0_outputs(2711) <= not(inputs(59)) or (inputs(190));
    layer0_outputs(2712) <= not(inputs(166));
    layer0_outputs(2713) <= (inputs(100)) xor (inputs(47));
    layer0_outputs(2714) <= not(inputs(130));
    layer0_outputs(2715) <= (inputs(58)) and not (inputs(251));
    layer0_outputs(2716) <= (inputs(35)) or (inputs(140));
    layer0_outputs(2717) <= (inputs(252)) xor (inputs(124));
    layer0_outputs(2718) <= inputs(133);
    layer0_outputs(2719) <= (inputs(159)) xor (inputs(214));
    layer0_outputs(2720) <= (inputs(106)) xor (inputs(125));
    layer0_outputs(2721) <= not(inputs(71)) or (inputs(44));
    layer0_outputs(2722) <= (inputs(28)) or (inputs(141));
    layer0_outputs(2723) <= (inputs(179)) xor (inputs(21));
    layer0_outputs(2724) <= not(inputs(167));
    layer0_outputs(2725) <= not(inputs(170)) or (inputs(197));
    layer0_outputs(2726) <= not((inputs(107)) xor (inputs(95)));
    layer0_outputs(2727) <= (inputs(112)) xor (inputs(74));
    layer0_outputs(2728) <= (inputs(250)) or (inputs(169));
    layer0_outputs(2729) <= not(inputs(28)) or (inputs(130));
    layer0_outputs(2730) <= inputs(57);
    layer0_outputs(2731) <= '0';
    layer0_outputs(2732) <= '0';
    layer0_outputs(2733) <= not(inputs(177));
    layer0_outputs(2734) <= not(inputs(58)) or (inputs(224));
    layer0_outputs(2735) <= not(inputs(33));
    layer0_outputs(2736) <= not(inputs(197)) or (inputs(132));
    layer0_outputs(2737) <= (inputs(134)) and not (inputs(33));
    layer0_outputs(2738) <= not((inputs(125)) or (inputs(103)));
    layer0_outputs(2739) <= (inputs(33)) or (inputs(136));
    layer0_outputs(2740) <= (inputs(199)) xor (inputs(48));
    layer0_outputs(2741) <= (inputs(100)) or (inputs(186));
    layer0_outputs(2742) <= inputs(194);
    layer0_outputs(2743) <= not((inputs(228)) xor (inputs(23)));
    layer0_outputs(2744) <= inputs(184);
    layer0_outputs(2745) <= (inputs(30)) xor (inputs(187));
    layer0_outputs(2746) <= not((inputs(100)) and (inputs(216)));
    layer0_outputs(2747) <= (inputs(196)) xor (inputs(8));
    layer0_outputs(2748) <= not((inputs(29)) or (inputs(183)));
    layer0_outputs(2749) <= not(inputs(58));
    layer0_outputs(2750) <= (inputs(39)) and (inputs(61));
    layer0_outputs(2751) <= (inputs(118)) and not (inputs(217));
    layer0_outputs(2752) <= not(inputs(231)) or (inputs(3));
    layer0_outputs(2753) <= not((inputs(149)) xor (inputs(173)));
    layer0_outputs(2754) <= (inputs(54)) and not (inputs(146));
    layer0_outputs(2755) <= not((inputs(216)) and (inputs(205)));
    layer0_outputs(2756) <= not((inputs(32)) xor (inputs(56)));
    layer0_outputs(2757) <= not(inputs(195)) or (inputs(17));
    layer0_outputs(2758) <= not((inputs(229)) xor (inputs(118)));
    layer0_outputs(2759) <= not(inputs(21));
    layer0_outputs(2760) <= (inputs(232)) xor (inputs(228));
    layer0_outputs(2761) <= inputs(185);
    layer0_outputs(2762) <= not(inputs(17)) or (inputs(227));
    layer0_outputs(2763) <= not(inputs(159));
    layer0_outputs(2764) <= not(inputs(74));
    layer0_outputs(2765) <= (inputs(203)) and not (inputs(226));
    layer0_outputs(2766) <= not((inputs(164)) or (inputs(178)));
    layer0_outputs(2767) <= not(inputs(65));
    layer0_outputs(2768) <= not(inputs(252));
    layer0_outputs(2769) <= not(inputs(43));
    layer0_outputs(2770) <= '0';
    layer0_outputs(2771) <= not(inputs(232));
    layer0_outputs(2772) <= not(inputs(42)) or (inputs(255));
    layer0_outputs(2773) <= (inputs(76)) xor (inputs(30));
    layer0_outputs(2774) <= not(inputs(28)) or (inputs(143));
    layer0_outputs(2775) <= (inputs(24)) xor (inputs(145));
    layer0_outputs(2776) <= not((inputs(213)) or (inputs(76)));
    layer0_outputs(2777) <= not((inputs(80)) and (inputs(96)));
    layer0_outputs(2778) <= (inputs(133)) or (inputs(7));
    layer0_outputs(2779) <= not((inputs(5)) or (inputs(86)));
    layer0_outputs(2780) <= not((inputs(162)) or (inputs(198)));
    layer0_outputs(2781) <= (inputs(11)) and (inputs(144));
    layer0_outputs(2782) <= (inputs(172)) or (inputs(177));
    layer0_outputs(2783) <= inputs(106);
    layer0_outputs(2784) <= inputs(10);
    layer0_outputs(2785) <= (inputs(76)) or (inputs(158));
    layer0_outputs(2786) <= not(inputs(212));
    layer0_outputs(2787) <= not((inputs(104)) or (inputs(35)));
    layer0_outputs(2788) <= '1';
    layer0_outputs(2789) <= not(inputs(198));
    layer0_outputs(2790) <= (inputs(250)) and not (inputs(147));
    layer0_outputs(2791) <= not((inputs(205)) xor (inputs(117)));
    layer0_outputs(2792) <= (inputs(92)) and not (inputs(183));
    layer0_outputs(2793) <= not((inputs(149)) or (inputs(170)));
    layer0_outputs(2794) <= (inputs(4)) and not (inputs(13));
    layer0_outputs(2795) <= not((inputs(26)) or (inputs(163)));
    layer0_outputs(2796) <= (inputs(230)) and not (inputs(6));
    layer0_outputs(2797) <= not(inputs(31)) or (inputs(39));
    layer0_outputs(2798) <= not((inputs(233)) or (inputs(47)));
    layer0_outputs(2799) <= not(inputs(101)) or (inputs(18));
    layer0_outputs(2800) <= (inputs(76)) or (inputs(211));
    layer0_outputs(2801) <= (inputs(189)) xor (inputs(242));
    layer0_outputs(2802) <= (inputs(43)) xor (inputs(176));
    layer0_outputs(2803) <= inputs(216);
    layer0_outputs(2804) <= not((inputs(130)) and (inputs(238)));
    layer0_outputs(2805) <= inputs(148);
    layer0_outputs(2806) <= not(inputs(160));
    layer0_outputs(2807) <= not(inputs(88)) or (inputs(63));
    layer0_outputs(2808) <= not(inputs(240)) or (inputs(53));
    layer0_outputs(2809) <= inputs(9);
    layer0_outputs(2810) <= (inputs(42)) xor (inputs(23));
    layer0_outputs(2811) <= not((inputs(84)) or (inputs(143)));
    layer0_outputs(2812) <= inputs(137);
    layer0_outputs(2813) <= not(inputs(158)) or (inputs(239));
    layer0_outputs(2814) <= '0';
    layer0_outputs(2815) <= not((inputs(56)) and (inputs(211)));
    layer0_outputs(2816) <= (inputs(171)) and not (inputs(44));
    layer0_outputs(2817) <= (inputs(47)) or (inputs(169));
    layer0_outputs(2818) <= (inputs(191)) or (inputs(92));
    layer0_outputs(2819) <= (inputs(53)) or (inputs(174));
    layer0_outputs(2820) <= inputs(58);
    layer0_outputs(2821) <= not((inputs(190)) or (inputs(207)));
    layer0_outputs(2822) <= not((inputs(74)) or (inputs(221)));
    layer0_outputs(2823) <= not(inputs(171));
    layer0_outputs(2824) <= inputs(89);
    layer0_outputs(2825) <= not((inputs(186)) or (inputs(82)));
    layer0_outputs(2826) <= not(inputs(157));
    layer0_outputs(2827) <= (inputs(173)) and not (inputs(113));
    layer0_outputs(2828) <= not((inputs(49)) xor (inputs(70)));
    layer0_outputs(2829) <= (inputs(119)) and not (inputs(115));
    layer0_outputs(2830) <= (inputs(179)) and not (inputs(99));
    layer0_outputs(2831) <= not(inputs(187)) or (inputs(131));
    layer0_outputs(2832) <= inputs(71);
    layer0_outputs(2833) <= not((inputs(160)) or (inputs(73)));
    layer0_outputs(2834) <= (inputs(225)) or (inputs(123));
    layer0_outputs(2835) <= not(inputs(145)) or (inputs(252));
    layer0_outputs(2836) <= (inputs(196)) or (inputs(215));
    layer0_outputs(2837) <= not(inputs(168));
    layer0_outputs(2838) <= not((inputs(64)) xor (inputs(156)));
    layer0_outputs(2839) <= inputs(169);
    layer0_outputs(2840) <= not(inputs(60)) or (inputs(27));
    layer0_outputs(2841) <= not(inputs(241));
    layer0_outputs(2842) <= (inputs(133)) or (inputs(114));
    layer0_outputs(2843) <= not((inputs(188)) xor (inputs(212)));
    layer0_outputs(2844) <= inputs(115);
    layer0_outputs(2845) <= (inputs(82)) and not (inputs(28));
    layer0_outputs(2846) <= not(inputs(186)) or (inputs(146));
    layer0_outputs(2847) <= not((inputs(217)) xor (inputs(176)));
    layer0_outputs(2848) <= not((inputs(67)) or (inputs(37)));
    layer0_outputs(2849) <= not((inputs(238)) xor (inputs(199)));
    layer0_outputs(2850) <= (inputs(208)) xor (inputs(111));
    layer0_outputs(2851) <= (inputs(189)) or (inputs(60));
    layer0_outputs(2852) <= inputs(140);
    layer0_outputs(2853) <= not(inputs(217));
    layer0_outputs(2854) <= '0';
    layer0_outputs(2855) <= not((inputs(134)) xor (inputs(143)));
    layer0_outputs(2856) <= not((inputs(17)) and (inputs(20)));
    layer0_outputs(2857) <= not(inputs(0)) or (inputs(190));
    layer0_outputs(2858) <= not(inputs(71)) or (inputs(104));
    layer0_outputs(2859) <= not((inputs(206)) or (inputs(238)));
    layer0_outputs(2860) <= inputs(195);
    layer0_outputs(2861) <= not(inputs(42));
    layer0_outputs(2862) <= not(inputs(106));
    layer0_outputs(2863) <= (inputs(236)) xor (inputs(106));
    layer0_outputs(2864) <= not(inputs(165)) or (inputs(180));
    layer0_outputs(2865) <= inputs(121);
    layer0_outputs(2866) <= inputs(131);
    layer0_outputs(2867) <= (inputs(80)) and not (inputs(35));
    layer0_outputs(2868) <= not(inputs(198)) or (inputs(130));
    layer0_outputs(2869) <= not((inputs(185)) or (inputs(158)));
    layer0_outputs(2870) <= (inputs(33)) and not (inputs(128));
    layer0_outputs(2871) <= (inputs(132)) or (inputs(1));
    layer0_outputs(2872) <= inputs(61);
    layer0_outputs(2873) <= not((inputs(131)) or (inputs(124)));
    layer0_outputs(2874) <= (inputs(132)) or (inputs(207));
    layer0_outputs(2875) <= not((inputs(210)) xor (inputs(38)));
    layer0_outputs(2876) <= not(inputs(8));
    layer0_outputs(2877) <= not((inputs(187)) xor (inputs(210)));
    layer0_outputs(2878) <= not((inputs(22)) and (inputs(111)));
    layer0_outputs(2879) <= (inputs(27)) or (inputs(183));
    layer0_outputs(2880) <= not((inputs(112)) xor (inputs(138)));
    layer0_outputs(2881) <= inputs(19);
    layer0_outputs(2882) <= (inputs(191)) or (inputs(118));
    layer0_outputs(2883) <= not(inputs(153)) or (inputs(1));
    layer0_outputs(2884) <= not(inputs(73)) or (inputs(43));
    layer0_outputs(2885) <= inputs(136);
    layer0_outputs(2886) <= not((inputs(158)) xor (inputs(250)));
    layer0_outputs(2887) <= (inputs(180)) xor (inputs(237));
    layer0_outputs(2888) <= '1';
    layer0_outputs(2889) <= not(inputs(231)) or (inputs(26));
    layer0_outputs(2890) <= inputs(101);
    layer0_outputs(2891) <= (inputs(43)) xor (inputs(158));
    layer0_outputs(2892) <= (inputs(168)) or (inputs(37));
    layer0_outputs(2893) <= inputs(108);
    layer0_outputs(2894) <= inputs(168);
    layer0_outputs(2895) <= not((inputs(185)) xor (inputs(110)));
    layer0_outputs(2896) <= (inputs(87)) or (inputs(108));
    layer0_outputs(2897) <= inputs(19);
    layer0_outputs(2898) <= inputs(102);
    layer0_outputs(2899) <= (inputs(166)) xor (inputs(113));
    layer0_outputs(2900) <= not(inputs(133)) or (inputs(22));
    layer0_outputs(2901) <= (inputs(11)) and not (inputs(26));
    layer0_outputs(2902) <= (inputs(95)) or (inputs(241));
    layer0_outputs(2903) <= not((inputs(229)) or (inputs(140)));
    layer0_outputs(2904) <= '1';
    layer0_outputs(2905) <= not(inputs(25)) or (inputs(194));
    layer0_outputs(2906) <= not((inputs(192)) xor (inputs(135)));
    layer0_outputs(2907) <= not((inputs(65)) and (inputs(184)));
    layer0_outputs(2908) <= '0';
    layer0_outputs(2909) <= not((inputs(72)) xor (inputs(154)));
    layer0_outputs(2910) <= not(inputs(44));
    layer0_outputs(2911) <= (inputs(138)) or (inputs(232));
    layer0_outputs(2912) <= not((inputs(168)) xor (inputs(88)));
    layer0_outputs(2913) <= not((inputs(16)) or (inputs(244)));
    layer0_outputs(2914) <= (inputs(66)) xor (inputs(230));
    layer0_outputs(2915) <= (inputs(218)) or (inputs(133));
    layer0_outputs(2916) <= inputs(140);
    layer0_outputs(2917) <= (inputs(86)) or (inputs(0));
    layer0_outputs(2918) <= not(inputs(148));
    layer0_outputs(2919) <= (inputs(117)) and not (inputs(180));
    layer0_outputs(2920) <= not((inputs(190)) or (inputs(125)));
    layer0_outputs(2921) <= not((inputs(221)) or (inputs(81)));
    layer0_outputs(2922) <= (inputs(0)) or (inputs(21));
    layer0_outputs(2923) <= not(inputs(100));
    layer0_outputs(2924) <= not((inputs(252)) or (inputs(238)));
    layer0_outputs(2925) <= (inputs(21)) xor (inputs(216));
    layer0_outputs(2926) <= (inputs(103)) and not (inputs(254));
    layer0_outputs(2927) <= not(inputs(48)) or (inputs(8));
    layer0_outputs(2928) <= inputs(106);
    layer0_outputs(2929) <= not(inputs(151));
    layer0_outputs(2930) <= (inputs(235)) xor (inputs(207));
    layer0_outputs(2931) <= not(inputs(217));
    layer0_outputs(2932) <= '1';
    layer0_outputs(2933) <= not(inputs(104)) or (inputs(145));
    layer0_outputs(2934) <= '1';
    layer0_outputs(2935) <= (inputs(232)) and not (inputs(109));
    layer0_outputs(2936) <= not((inputs(182)) xor (inputs(10)));
    layer0_outputs(2937) <= (inputs(218)) or (inputs(255));
    layer0_outputs(2938) <= inputs(117);
    layer0_outputs(2939) <= not((inputs(92)) xor (inputs(123)));
    layer0_outputs(2940) <= not(inputs(228));
    layer0_outputs(2941) <= not((inputs(142)) or (inputs(183)));
    layer0_outputs(2942) <= '0';
    layer0_outputs(2943) <= not((inputs(203)) xor (inputs(115)));
    layer0_outputs(2944) <= (inputs(154)) and not (inputs(174));
    layer0_outputs(2945) <= (inputs(43)) xor (inputs(94));
    layer0_outputs(2946) <= not(inputs(85)) or (inputs(52));
    layer0_outputs(2947) <= '1';
    layer0_outputs(2948) <= (inputs(223)) and not (inputs(176));
    layer0_outputs(2949) <= not(inputs(197)) or (inputs(29));
    layer0_outputs(2950) <= (inputs(85)) and not (inputs(124));
    layer0_outputs(2951) <= not(inputs(74)) or (inputs(38));
    layer0_outputs(2952) <= not((inputs(167)) xor (inputs(10)));
    layer0_outputs(2953) <= (inputs(163)) xor (inputs(116));
    layer0_outputs(2954) <= '1';
    layer0_outputs(2955) <= (inputs(140)) and not (inputs(130));
    layer0_outputs(2956) <= (inputs(42)) and not (inputs(253));
    layer0_outputs(2957) <= not((inputs(47)) and (inputs(251)));
    layer0_outputs(2958) <= (inputs(183)) and not (inputs(194));
    layer0_outputs(2959) <= inputs(200);
    layer0_outputs(2960) <= (inputs(169)) and not (inputs(10));
    layer0_outputs(2961) <= not(inputs(114)) or (inputs(220));
    layer0_outputs(2962) <= (inputs(0)) and not (inputs(37));
    layer0_outputs(2963) <= (inputs(87)) and not (inputs(216));
    layer0_outputs(2964) <= (inputs(52)) and not (inputs(242));
    layer0_outputs(2965) <= inputs(89);
    layer0_outputs(2966) <= not((inputs(157)) xor (inputs(159)));
    layer0_outputs(2967) <= not(inputs(111)) or (inputs(14));
    layer0_outputs(2968) <= (inputs(113)) and not (inputs(250));
    layer0_outputs(2969) <= (inputs(161)) and not (inputs(205));
    layer0_outputs(2970) <= not((inputs(74)) or (inputs(92)));
    layer0_outputs(2971) <= (inputs(59)) and not (inputs(38));
    layer0_outputs(2972) <= not(inputs(128)) or (inputs(33));
    layer0_outputs(2973) <= not(inputs(59));
    layer0_outputs(2974) <= (inputs(1)) and not (inputs(195));
    layer0_outputs(2975) <= not((inputs(41)) or (inputs(172)));
    layer0_outputs(2976) <= not((inputs(172)) or (inputs(40)));
    layer0_outputs(2977) <= not(inputs(100));
    layer0_outputs(2978) <= not(inputs(100));
    layer0_outputs(2979) <= (inputs(58)) and not (inputs(44));
    layer0_outputs(2980) <= not(inputs(216)) or (inputs(17));
    layer0_outputs(2981) <= not((inputs(60)) and (inputs(63)));
    layer0_outputs(2982) <= (inputs(9)) or (inputs(225));
    layer0_outputs(2983) <= not((inputs(31)) or (inputs(248)));
    layer0_outputs(2984) <= (inputs(96)) xor (inputs(146));
    layer0_outputs(2985) <= not(inputs(71));
    layer0_outputs(2986) <= not(inputs(73));
    layer0_outputs(2987) <= (inputs(80)) xor (inputs(169));
    layer0_outputs(2988) <= inputs(58);
    layer0_outputs(2989) <= (inputs(146)) or (inputs(48));
    layer0_outputs(2990) <= '0';
    layer0_outputs(2991) <= (inputs(30)) xor (inputs(104));
    layer0_outputs(2992) <= not(inputs(184)) or (inputs(251));
    layer0_outputs(2993) <= (inputs(20)) or (inputs(37));
    layer0_outputs(2994) <= (inputs(156)) xor (inputs(211));
    layer0_outputs(2995) <= not(inputs(57));
    layer0_outputs(2996) <= inputs(126);
    layer0_outputs(2997) <= not(inputs(232)) or (inputs(158));
    layer0_outputs(2998) <= (inputs(79)) xor (inputs(133));
    layer0_outputs(2999) <= not(inputs(223));
    layer0_outputs(3000) <= (inputs(73)) xor (inputs(190));
    layer0_outputs(3001) <= not((inputs(26)) xor (inputs(75)));
    layer0_outputs(3002) <= '1';
    layer0_outputs(3003) <= inputs(133);
    layer0_outputs(3004) <= (inputs(121)) and not (inputs(102));
    layer0_outputs(3005) <= not(inputs(107)) or (inputs(210));
    layer0_outputs(3006) <= inputs(42);
    layer0_outputs(3007) <= not((inputs(113)) xor (inputs(86)));
    layer0_outputs(3008) <= inputs(199);
    layer0_outputs(3009) <= (inputs(46)) xor (inputs(199));
    layer0_outputs(3010) <= (inputs(233)) or (inputs(89));
    layer0_outputs(3011) <= not(inputs(241)) or (inputs(95));
    layer0_outputs(3012) <= inputs(71);
    layer0_outputs(3013) <= '0';
    layer0_outputs(3014) <= not(inputs(188)) or (inputs(94));
    layer0_outputs(3015) <= not(inputs(176));
    layer0_outputs(3016) <= (inputs(9)) and not (inputs(244));
    layer0_outputs(3017) <= not(inputs(85)) or (inputs(25));
    layer0_outputs(3018) <= (inputs(103)) or (inputs(97));
    layer0_outputs(3019) <= (inputs(145)) xor (inputs(138));
    layer0_outputs(3020) <= (inputs(77)) and not (inputs(161));
    layer0_outputs(3021) <= (inputs(23)) and not (inputs(1));
    layer0_outputs(3022) <= not(inputs(205)) or (inputs(18));
    layer0_outputs(3023) <= not(inputs(115)) or (inputs(14));
    layer0_outputs(3024) <= (inputs(217)) or (inputs(58));
    layer0_outputs(3025) <= not(inputs(249)) or (inputs(209));
    layer0_outputs(3026) <= not((inputs(95)) and (inputs(74)));
    layer0_outputs(3027) <= (inputs(55)) and not (inputs(62));
    layer0_outputs(3028) <= '0';
    layer0_outputs(3029) <= not(inputs(168)) or (inputs(246));
    layer0_outputs(3030) <= (inputs(167)) or (inputs(93));
    layer0_outputs(3031) <= not((inputs(178)) xor (inputs(63)));
    layer0_outputs(3032) <= not((inputs(235)) or (inputs(99)));
    layer0_outputs(3033) <= not(inputs(72));
    layer0_outputs(3034) <= '1';
    layer0_outputs(3035) <= inputs(195);
    layer0_outputs(3036) <= not(inputs(117));
    layer0_outputs(3037) <= not((inputs(131)) or (inputs(232)));
    layer0_outputs(3038) <= not((inputs(69)) or (inputs(39)));
    layer0_outputs(3039) <= (inputs(28)) or (inputs(180));
    layer0_outputs(3040) <= not(inputs(165));
    layer0_outputs(3041) <= not(inputs(175));
    layer0_outputs(3042) <= not(inputs(148)) or (inputs(38));
    layer0_outputs(3043) <= (inputs(164)) or (inputs(106));
    layer0_outputs(3044) <= not(inputs(42));
    layer0_outputs(3045) <= '0';
    layer0_outputs(3046) <= inputs(154);
    layer0_outputs(3047) <= '0';
    layer0_outputs(3048) <= inputs(66);
    layer0_outputs(3049) <= not(inputs(214));
    layer0_outputs(3050) <= not((inputs(188)) or (inputs(106)));
    layer0_outputs(3051) <= not(inputs(144)) or (inputs(253));
    layer0_outputs(3052) <= (inputs(145)) and (inputs(208));
    layer0_outputs(3053) <= not((inputs(232)) xor (inputs(233)));
    layer0_outputs(3054) <= (inputs(172)) and not (inputs(209));
    layer0_outputs(3055) <= inputs(183);
    layer0_outputs(3056) <= (inputs(226)) xor (inputs(131));
    layer0_outputs(3057) <= not((inputs(76)) or (inputs(171)));
    layer0_outputs(3058) <= (inputs(46)) and not (inputs(218));
    layer0_outputs(3059) <= not(inputs(223)) or (inputs(46));
    layer0_outputs(3060) <= not((inputs(30)) and (inputs(15)));
    layer0_outputs(3061) <= inputs(101);
    layer0_outputs(3062) <= not(inputs(75));
    layer0_outputs(3063) <= not(inputs(152)) or (inputs(162));
    layer0_outputs(3064) <= not((inputs(95)) xor (inputs(11)));
    layer0_outputs(3065) <= (inputs(211)) xor (inputs(47));
    layer0_outputs(3066) <= not((inputs(247)) or (inputs(150)));
    layer0_outputs(3067) <= inputs(172);
    layer0_outputs(3068) <= not((inputs(231)) xor (inputs(71)));
    layer0_outputs(3069) <= not(inputs(59)) or (inputs(22));
    layer0_outputs(3070) <= (inputs(3)) or (inputs(178));
    layer0_outputs(3071) <= not((inputs(218)) and (inputs(208)));
    layer0_outputs(3072) <= (inputs(12)) xor (inputs(254));
    layer0_outputs(3073) <= (inputs(141)) or (inputs(60));
    layer0_outputs(3074) <= inputs(134);
    layer0_outputs(3075) <= not(inputs(54));
    layer0_outputs(3076) <= inputs(122);
    layer0_outputs(3077) <= not((inputs(226)) or (inputs(38)));
    layer0_outputs(3078) <= not(inputs(189));
    layer0_outputs(3079) <= (inputs(222)) or (inputs(223));
    layer0_outputs(3080) <= (inputs(145)) and not (inputs(49));
    layer0_outputs(3081) <= not((inputs(56)) xor (inputs(40)));
    layer0_outputs(3082) <= (inputs(9)) and not (inputs(147));
    layer0_outputs(3083) <= inputs(99);
    layer0_outputs(3084) <= not((inputs(16)) or (inputs(154)));
    layer0_outputs(3085) <= (inputs(144)) or (inputs(222));
    layer0_outputs(3086) <= not(inputs(147)) or (inputs(81));
    layer0_outputs(3087) <= (inputs(201)) and not (inputs(193));
    layer0_outputs(3088) <= (inputs(226)) and not (inputs(13));
    layer0_outputs(3089) <= not((inputs(11)) or (inputs(154)));
    layer0_outputs(3090) <= not(inputs(180)) or (inputs(10));
    layer0_outputs(3091) <= inputs(87);
    layer0_outputs(3092) <= (inputs(92)) or (inputs(84));
    layer0_outputs(3093) <= inputs(215);
    layer0_outputs(3094) <= '0';
    layer0_outputs(3095) <= inputs(178);
    layer0_outputs(3096) <= '0';
    layer0_outputs(3097) <= not(inputs(132));
    layer0_outputs(3098) <= not((inputs(208)) or (inputs(45)));
    layer0_outputs(3099) <= '0';
    layer0_outputs(3100) <= inputs(132);
    layer0_outputs(3101) <= not(inputs(6)) or (inputs(115));
    layer0_outputs(3102) <= not(inputs(147));
    layer0_outputs(3103) <= (inputs(49)) xor (inputs(58));
    layer0_outputs(3104) <= inputs(77);
    layer0_outputs(3105) <= not(inputs(143));
    layer0_outputs(3106) <= inputs(86);
    layer0_outputs(3107) <= (inputs(175)) xor (inputs(75));
    layer0_outputs(3108) <= (inputs(187)) or (inputs(96));
    layer0_outputs(3109) <= not((inputs(64)) xor (inputs(88)));
    layer0_outputs(3110) <= not(inputs(145)) or (inputs(239));
    layer0_outputs(3111) <= not(inputs(80));
    layer0_outputs(3112) <= (inputs(108)) and not (inputs(254));
    layer0_outputs(3113) <= not((inputs(36)) or (inputs(155)));
    layer0_outputs(3114) <= not(inputs(86));
    layer0_outputs(3115) <= (inputs(57)) and not (inputs(178));
    layer0_outputs(3116) <= not(inputs(149));
    layer0_outputs(3117) <= (inputs(3)) or (inputs(163));
    layer0_outputs(3118) <= not(inputs(95));
    layer0_outputs(3119) <= not(inputs(102));
    layer0_outputs(3120) <= (inputs(100)) and not (inputs(116));
    layer0_outputs(3121) <= (inputs(233)) and not (inputs(226));
    layer0_outputs(3122) <= (inputs(118)) or (inputs(149));
    layer0_outputs(3123) <= not((inputs(232)) or (inputs(68)));
    layer0_outputs(3124) <= (inputs(112)) xor (inputs(88));
    layer0_outputs(3125) <= (inputs(96)) xor (inputs(206));
    layer0_outputs(3126) <= '0';
    layer0_outputs(3127) <= not(inputs(74)) or (inputs(129));
    layer0_outputs(3128) <= inputs(150);
    layer0_outputs(3129) <= (inputs(137)) and not (inputs(38));
    layer0_outputs(3130) <= inputs(76);
    layer0_outputs(3131) <= not(inputs(165)) or (inputs(2));
    layer0_outputs(3132) <= not((inputs(197)) or (inputs(46)));
    layer0_outputs(3133) <= not((inputs(75)) and (inputs(121)));
    layer0_outputs(3134) <= inputs(62);
    layer0_outputs(3135) <= not(inputs(53)) or (inputs(99));
    layer0_outputs(3136) <= (inputs(251)) and (inputs(12));
    layer0_outputs(3137) <= not(inputs(130)) or (inputs(14));
    layer0_outputs(3138) <= '0';
    layer0_outputs(3139) <= not((inputs(0)) and (inputs(251)));
    layer0_outputs(3140) <= not(inputs(118)) or (inputs(130));
    layer0_outputs(3141) <= not(inputs(217));
    layer0_outputs(3142) <= (inputs(57)) and not (inputs(44));
    layer0_outputs(3143) <= (inputs(55)) and not (inputs(190));
    layer0_outputs(3144) <= inputs(148);
    layer0_outputs(3145) <= inputs(210);
    layer0_outputs(3146) <= (inputs(245)) xor (inputs(158));
    layer0_outputs(3147) <= not(inputs(55));
    layer0_outputs(3148) <= (inputs(93)) xor (inputs(61));
    layer0_outputs(3149) <= (inputs(220)) xor (inputs(47));
    layer0_outputs(3150) <= (inputs(225)) xor (inputs(59));
    layer0_outputs(3151) <= not(inputs(166));
    layer0_outputs(3152) <= not(inputs(179));
    layer0_outputs(3153) <= inputs(200);
    layer0_outputs(3154) <= not((inputs(81)) or (inputs(234)));
    layer0_outputs(3155) <= not(inputs(13)) or (inputs(240));
    layer0_outputs(3156) <= not(inputs(154));
    layer0_outputs(3157) <= (inputs(238)) xor (inputs(106));
    layer0_outputs(3158) <= not(inputs(92));
    layer0_outputs(3159) <= not(inputs(53)) or (inputs(5));
    layer0_outputs(3160) <= not((inputs(158)) xor (inputs(242)));
    layer0_outputs(3161) <= (inputs(213)) or (inputs(187));
    layer0_outputs(3162) <= not(inputs(6));
    layer0_outputs(3163) <= (inputs(23)) xor (inputs(44));
    layer0_outputs(3164) <= (inputs(84)) and not (inputs(126));
    layer0_outputs(3165) <= (inputs(105)) and not (inputs(236));
    layer0_outputs(3166) <= (inputs(24)) or (inputs(69));
    layer0_outputs(3167) <= (inputs(179)) and not (inputs(36));
    layer0_outputs(3168) <= (inputs(21)) or (inputs(143));
    layer0_outputs(3169) <= not(inputs(106)) or (inputs(235));
    layer0_outputs(3170) <= (inputs(41)) or (inputs(229));
    layer0_outputs(3171) <= not((inputs(104)) xor (inputs(76)));
    layer0_outputs(3172) <= not((inputs(87)) or (inputs(252)));
    layer0_outputs(3173) <= not((inputs(19)) xor (inputs(207)));
    layer0_outputs(3174) <= not((inputs(3)) and (inputs(223)));
    layer0_outputs(3175) <= (inputs(229)) and not (inputs(170));
    layer0_outputs(3176) <= (inputs(204)) or (inputs(248));
    layer0_outputs(3177) <= (inputs(26)) or (inputs(152));
    layer0_outputs(3178) <= '0';
    layer0_outputs(3179) <= (inputs(198)) xor (inputs(5));
    layer0_outputs(3180) <= (inputs(81)) or (inputs(140));
    layer0_outputs(3181) <= not(inputs(250));
    layer0_outputs(3182) <= not((inputs(204)) or (inputs(89)));
    layer0_outputs(3183) <= not(inputs(4)) or (inputs(218));
    layer0_outputs(3184) <= '0';
    layer0_outputs(3185) <= (inputs(107)) or (inputs(217));
    layer0_outputs(3186) <= (inputs(160)) or (inputs(5));
    layer0_outputs(3187) <= not((inputs(24)) or (inputs(62)));
    layer0_outputs(3188) <= not((inputs(200)) and (inputs(111)));
    layer0_outputs(3189) <= not(inputs(182)) or (inputs(231));
    layer0_outputs(3190) <= not((inputs(172)) xor (inputs(42)));
    layer0_outputs(3191) <= not((inputs(141)) or (inputs(62)));
    layer0_outputs(3192) <= not(inputs(171));
    layer0_outputs(3193) <= inputs(120);
    layer0_outputs(3194) <= (inputs(170)) and not (inputs(240));
    layer0_outputs(3195) <= inputs(159);
    layer0_outputs(3196) <= (inputs(43)) or (inputs(190));
    layer0_outputs(3197) <= not(inputs(228));
    layer0_outputs(3198) <= '0';
    layer0_outputs(3199) <= not(inputs(99)) or (inputs(187));
    layer0_outputs(3200) <= not(inputs(85));
    layer0_outputs(3201) <= (inputs(127)) and (inputs(65));
    layer0_outputs(3202) <= (inputs(64)) xor (inputs(201));
    layer0_outputs(3203) <= (inputs(136)) or (inputs(5));
    layer0_outputs(3204) <= inputs(52);
    layer0_outputs(3205) <= not(inputs(241)) or (inputs(211));
    layer0_outputs(3206) <= not((inputs(190)) and (inputs(206)));
    layer0_outputs(3207) <= (inputs(196)) xor (inputs(201));
    layer0_outputs(3208) <= not(inputs(128));
    layer0_outputs(3209) <= (inputs(119)) or (inputs(205));
    layer0_outputs(3210) <= (inputs(235)) or (inputs(124));
    layer0_outputs(3211) <= (inputs(102)) or (inputs(238));
    layer0_outputs(3212) <= not((inputs(155)) or (inputs(186)));
    layer0_outputs(3213) <= (inputs(26)) and not (inputs(80));
    layer0_outputs(3214) <= (inputs(12)) xor (inputs(59));
    layer0_outputs(3215) <= not(inputs(10)) or (inputs(144));
    layer0_outputs(3216) <= not((inputs(123)) or (inputs(2)));
    layer0_outputs(3217) <= inputs(38);
    layer0_outputs(3218) <= not(inputs(251)) or (inputs(249));
    layer0_outputs(3219) <= (inputs(158)) xor (inputs(113));
    layer0_outputs(3220) <= (inputs(83)) or (inputs(171));
    layer0_outputs(3221) <= not(inputs(23)) or (inputs(48));
    layer0_outputs(3222) <= not(inputs(185)) or (inputs(236));
    layer0_outputs(3223) <= not(inputs(181)) or (inputs(95));
    layer0_outputs(3224) <= (inputs(141)) or (inputs(210));
    layer0_outputs(3225) <= (inputs(185)) xor (inputs(236));
    layer0_outputs(3226) <= (inputs(161)) or (inputs(118));
    layer0_outputs(3227) <= (inputs(197)) or (inputs(221));
    layer0_outputs(3228) <= inputs(47);
    layer0_outputs(3229) <= not(inputs(44));
    layer0_outputs(3230) <= (inputs(172)) or (inputs(46));
    layer0_outputs(3231) <= (inputs(109)) xor (inputs(209));
    layer0_outputs(3232) <= inputs(117);
    layer0_outputs(3233) <= inputs(89);
    layer0_outputs(3234) <= not(inputs(2));
    layer0_outputs(3235) <= (inputs(74)) xor (inputs(96));
    layer0_outputs(3236) <= not(inputs(73)) or (inputs(4));
    layer0_outputs(3237) <= not(inputs(201)) or (inputs(9));
    layer0_outputs(3238) <= not(inputs(198)) or (inputs(192));
    layer0_outputs(3239) <= not((inputs(100)) xor (inputs(209)));
    layer0_outputs(3240) <= (inputs(108)) xor (inputs(79));
    layer0_outputs(3241) <= '0';
    layer0_outputs(3242) <= (inputs(155)) and not (inputs(113));
    layer0_outputs(3243) <= not((inputs(201)) xor (inputs(248)));
    layer0_outputs(3244) <= (inputs(158)) xor (inputs(107));
    layer0_outputs(3245) <= not((inputs(42)) xor (inputs(55)));
    layer0_outputs(3246) <= (inputs(29)) or (inputs(132));
    layer0_outputs(3247) <= (inputs(124)) or (inputs(245));
    layer0_outputs(3248) <= not((inputs(172)) or (inputs(21)));
    layer0_outputs(3249) <= (inputs(112)) xor (inputs(107));
    layer0_outputs(3250) <= (inputs(137)) or (inputs(92));
    layer0_outputs(3251) <= inputs(135);
    layer0_outputs(3252) <= not((inputs(55)) xor (inputs(63)));
    layer0_outputs(3253) <= (inputs(35)) xor (inputs(34));
    layer0_outputs(3254) <= (inputs(17)) and not (inputs(103));
    layer0_outputs(3255) <= not(inputs(102)) or (inputs(168));
    layer0_outputs(3256) <= (inputs(105)) and not (inputs(78));
    layer0_outputs(3257) <= not((inputs(123)) or (inputs(209)));
    layer0_outputs(3258) <= not((inputs(135)) or (inputs(57)));
    layer0_outputs(3259) <= (inputs(13)) and not (inputs(231));
    layer0_outputs(3260) <= not((inputs(242)) and (inputs(235)));
    layer0_outputs(3261) <= (inputs(123)) xor (inputs(105));
    layer0_outputs(3262) <= (inputs(40)) or (inputs(41));
    layer0_outputs(3263) <= not(inputs(51)) or (inputs(79));
    layer0_outputs(3264) <= not(inputs(11));
    layer0_outputs(3265) <= (inputs(47)) or (inputs(245));
    layer0_outputs(3266) <= (inputs(231)) and not (inputs(244));
    layer0_outputs(3267) <= not(inputs(150));
    layer0_outputs(3268) <= (inputs(213)) and not (inputs(42));
    layer0_outputs(3269) <= inputs(45);
    layer0_outputs(3270) <= not((inputs(83)) or (inputs(71)));
    layer0_outputs(3271) <= not((inputs(6)) and (inputs(245)));
    layer0_outputs(3272) <= (inputs(6)) and not (inputs(82));
    layer0_outputs(3273) <= (inputs(121)) or (inputs(68));
    layer0_outputs(3274) <= not((inputs(52)) xor (inputs(19)));
    layer0_outputs(3275) <= (inputs(58)) or (inputs(155));
    layer0_outputs(3276) <= not(inputs(110));
    layer0_outputs(3277) <= (inputs(127)) and (inputs(222));
    layer0_outputs(3278) <= (inputs(186)) and not (inputs(150));
    layer0_outputs(3279) <= not((inputs(196)) and (inputs(236)));
    layer0_outputs(3280) <= not((inputs(72)) or (inputs(244)));
    layer0_outputs(3281) <= (inputs(182)) and not (inputs(47));
    layer0_outputs(3282) <= not((inputs(167)) or (inputs(191)));
    layer0_outputs(3283) <= (inputs(190)) and not (inputs(1));
    layer0_outputs(3284) <= not(inputs(176));
    layer0_outputs(3285) <= '1';
    layer0_outputs(3286) <= not((inputs(52)) xor (inputs(210)));
    layer0_outputs(3287) <= (inputs(34)) or (inputs(85));
    layer0_outputs(3288) <= not(inputs(225)) or (inputs(46));
    layer0_outputs(3289) <= inputs(149);
    layer0_outputs(3290) <= not((inputs(49)) or (inputs(60)));
    layer0_outputs(3291) <= (inputs(201)) or (inputs(129));
    layer0_outputs(3292) <= not((inputs(70)) or (inputs(106)));
    layer0_outputs(3293) <= (inputs(198)) and not (inputs(34));
    layer0_outputs(3294) <= not((inputs(199)) or (inputs(94)));
    layer0_outputs(3295) <= not(inputs(148));
    layer0_outputs(3296) <= not(inputs(148)) or (inputs(113));
    layer0_outputs(3297) <= not(inputs(59)) or (inputs(17));
    layer0_outputs(3298) <= not(inputs(173));
    layer0_outputs(3299) <= (inputs(85)) or (inputs(102));
    layer0_outputs(3300) <= (inputs(211)) or (inputs(125));
    layer0_outputs(3301) <= (inputs(161)) xor (inputs(179));
    layer0_outputs(3302) <= not(inputs(89)) or (inputs(5));
    layer0_outputs(3303) <= inputs(165);
    layer0_outputs(3304) <= not(inputs(249));
    layer0_outputs(3305) <= (inputs(174)) or (inputs(55));
    layer0_outputs(3306) <= (inputs(117)) and (inputs(242));
    layer0_outputs(3307) <= '0';
    layer0_outputs(3308) <= not(inputs(154)) or (inputs(70));
    layer0_outputs(3309) <= inputs(46);
    layer0_outputs(3310) <= not(inputs(3)) or (inputs(94));
    layer0_outputs(3311) <= (inputs(193)) xor (inputs(29));
    layer0_outputs(3312) <= (inputs(56)) and not (inputs(44));
    layer0_outputs(3313) <= '1';
    layer0_outputs(3314) <= not((inputs(244)) and (inputs(224)));
    layer0_outputs(3315) <= inputs(182);
    layer0_outputs(3316) <= inputs(120);
    layer0_outputs(3317) <= not(inputs(106)) or (inputs(62));
    layer0_outputs(3318) <= inputs(149);
    layer0_outputs(3319) <= not((inputs(3)) xor (inputs(155)));
    layer0_outputs(3320) <= not((inputs(172)) or (inputs(54)));
    layer0_outputs(3321) <= not((inputs(251)) or (inputs(80)));
    layer0_outputs(3322) <= not(inputs(96));
    layer0_outputs(3323) <= inputs(52);
    layer0_outputs(3324) <= not(inputs(121));
    layer0_outputs(3325) <= inputs(170);
    layer0_outputs(3326) <= not((inputs(237)) or (inputs(121)));
    layer0_outputs(3327) <= not(inputs(89));
    layer0_outputs(3328) <= not((inputs(119)) or (inputs(94)));
    layer0_outputs(3329) <= not(inputs(159)) or (inputs(227));
    layer0_outputs(3330) <= not((inputs(184)) or (inputs(174)));
    layer0_outputs(3331) <= not(inputs(181));
    layer0_outputs(3332) <= (inputs(213)) or (inputs(239));
    layer0_outputs(3333) <= not(inputs(136));
    layer0_outputs(3334) <= not(inputs(13)) or (inputs(223));
    layer0_outputs(3335) <= (inputs(34)) or (inputs(237));
    layer0_outputs(3336) <= (inputs(199)) and not (inputs(237));
    layer0_outputs(3337) <= (inputs(184)) and not (inputs(1));
    layer0_outputs(3338) <= (inputs(160)) xor (inputs(180));
    layer0_outputs(3339) <= not(inputs(31)) or (inputs(255));
    layer0_outputs(3340) <= (inputs(72)) and not (inputs(222));
    layer0_outputs(3341) <= (inputs(84)) and not (inputs(179));
    layer0_outputs(3342) <= (inputs(49)) and not (inputs(208));
    layer0_outputs(3343) <= (inputs(208)) or (inputs(81));
    layer0_outputs(3344) <= (inputs(91)) and not (inputs(84));
    layer0_outputs(3345) <= not(inputs(189));
    layer0_outputs(3346) <= inputs(133);
    layer0_outputs(3347) <= (inputs(2)) xor (inputs(111));
    layer0_outputs(3348) <= (inputs(180)) and not (inputs(224));
    layer0_outputs(3349) <= not(inputs(114));
    layer0_outputs(3350) <= not((inputs(216)) or (inputs(10)));
    layer0_outputs(3351) <= inputs(86);
    layer0_outputs(3352) <= not((inputs(35)) or (inputs(188)));
    layer0_outputs(3353) <= (inputs(234)) and not (inputs(216));
    layer0_outputs(3354) <= (inputs(45)) or (inputs(96));
    layer0_outputs(3355) <= not((inputs(138)) or (inputs(50)));
    layer0_outputs(3356) <= (inputs(234)) and not (inputs(5));
    layer0_outputs(3357) <= not((inputs(81)) and (inputs(14)));
    layer0_outputs(3358) <= not(inputs(77));
    layer0_outputs(3359) <= not((inputs(43)) xor (inputs(51)));
    layer0_outputs(3360) <= not(inputs(224));
    layer0_outputs(3361) <= not((inputs(95)) and (inputs(31)));
    layer0_outputs(3362) <= not(inputs(101)) or (inputs(49));
    layer0_outputs(3363) <= '1';
    layer0_outputs(3364) <= not((inputs(5)) and (inputs(22)));
    layer0_outputs(3365) <= not((inputs(222)) or (inputs(188)));
    layer0_outputs(3366) <= not(inputs(152));
    layer0_outputs(3367) <= inputs(90);
    layer0_outputs(3368) <= inputs(126);
    layer0_outputs(3369) <= '0';
    layer0_outputs(3370) <= (inputs(2)) and not (inputs(38));
    layer0_outputs(3371) <= (inputs(192)) xor (inputs(69));
    layer0_outputs(3372) <= not((inputs(169)) or (inputs(136)));
    layer0_outputs(3373) <= (inputs(67)) xor (inputs(199));
    layer0_outputs(3374) <= (inputs(6)) and not (inputs(232));
    layer0_outputs(3375) <= not((inputs(26)) xor (inputs(241)));
    layer0_outputs(3376) <= (inputs(123)) or (inputs(15));
    layer0_outputs(3377) <= not((inputs(103)) or (inputs(250)));
    layer0_outputs(3378) <= not((inputs(133)) or (inputs(99)));
    layer0_outputs(3379) <= '0';
    layer0_outputs(3380) <= not(inputs(140));
    layer0_outputs(3381) <= not((inputs(180)) or (inputs(1)));
    layer0_outputs(3382) <= inputs(207);
    layer0_outputs(3383) <= inputs(227);
    layer0_outputs(3384) <= (inputs(191)) xor (inputs(56));
    layer0_outputs(3385) <= not(inputs(7));
    layer0_outputs(3386) <= (inputs(38)) or (inputs(141));
    layer0_outputs(3387) <= not((inputs(242)) xor (inputs(129)));
    layer0_outputs(3388) <= not(inputs(196));
    layer0_outputs(3389) <= not(inputs(200)) or (inputs(90));
    layer0_outputs(3390) <= (inputs(222)) xor (inputs(69));
    layer0_outputs(3391) <= (inputs(179)) and not (inputs(81));
    layer0_outputs(3392) <= inputs(149);
    layer0_outputs(3393) <= not(inputs(124));
    layer0_outputs(3394) <= not(inputs(247));
    layer0_outputs(3395) <= (inputs(206)) xor (inputs(185));
    layer0_outputs(3396) <= inputs(137);
    layer0_outputs(3397) <= (inputs(94)) or (inputs(227));
    layer0_outputs(3398) <= not(inputs(104));
    layer0_outputs(3399) <= not(inputs(58)) or (inputs(135));
    layer0_outputs(3400) <= (inputs(191)) and not (inputs(193));
    layer0_outputs(3401) <= not(inputs(120));
    layer0_outputs(3402) <= (inputs(58)) xor (inputs(219));
    layer0_outputs(3403) <= not(inputs(229)) or (inputs(193));
    layer0_outputs(3404) <= (inputs(19)) or (inputs(243));
    layer0_outputs(3405) <= not((inputs(255)) xor (inputs(173)));
    layer0_outputs(3406) <= not((inputs(126)) and (inputs(98)));
    layer0_outputs(3407) <= (inputs(243)) or (inputs(126));
    layer0_outputs(3408) <= inputs(41);
    layer0_outputs(3409) <= (inputs(53)) xor (inputs(18));
    layer0_outputs(3410) <= not(inputs(76));
    layer0_outputs(3411) <= not((inputs(80)) xor (inputs(194)));
    layer0_outputs(3412) <= not((inputs(91)) xor (inputs(126)));
    layer0_outputs(3413) <= '0';
    layer0_outputs(3414) <= (inputs(153)) and not (inputs(174));
    layer0_outputs(3415) <= not(inputs(101));
    layer0_outputs(3416) <= (inputs(255)) and not (inputs(47));
    layer0_outputs(3417) <= not((inputs(230)) xor (inputs(132)));
    layer0_outputs(3418) <= '0';
    layer0_outputs(3419) <= not(inputs(151));
    layer0_outputs(3420) <= not((inputs(86)) or (inputs(94)));
    layer0_outputs(3421) <= inputs(133);
    layer0_outputs(3422) <= not(inputs(181));
    layer0_outputs(3423) <= inputs(225);
    layer0_outputs(3424) <= not(inputs(108)) or (inputs(111));
    layer0_outputs(3425) <= not((inputs(74)) or (inputs(37)));
    layer0_outputs(3426) <= inputs(223);
    layer0_outputs(3427) <= (inputs(211)) xor (inputs(51));
    layer0_outputs(3428) <= not((inputs(250)) and (inputs(215)));
    layer0_outputs(3429) <= (inputs(109)) or (inputs(198));
    layer0_outputs(3430) <= '0';
    layer0_outputs(3431) <= (inputs(29)) or (inputs(242));
    layer0_outputs(3432) <= (inputs(174)) and not (inputs(95));
    layer0_outputs(3433) <= not(inputs(27)) or (inputs(224));
    layer0_outputs(3434) <= (inputs(68)) or (inputs(65));
    layer0_outputs(3435) <= not((inputs(250)) or (inputs(113)));
    layer0_outputs(3436) <= not((inputs(247)) xor (inputs(211)));
    layer0_outputs(3437) <= (inputs(36)) or (inputs(239));
    layer0_outputs(3438) <= not((inputs(54)) or (inputs(182)));
    layer0_outputs(3439) <= (inputs(165)) and not (inputs(162));
    layer0_outputs(3440) <= (inputs(180)) and not (inputs(105));
    layer0_outputs(3441) <= not((inputs(83)) xor (inputs(17)));
    layer0_outputs(3442) <= not(inputs(200)) or (inputs(14));
    layer0_outputs(3443) <= inputs(125);
    layer0_outputs(3444) <= (inputs(217)) and not (inputs(226));
    layer0_outputs(3445) <= (inputs(109)) or (inputs(140));
    layer0_outputs(3446) <= (inputs(208)) or (inputs(153));
    layer0_outputs(3447) <= (inputs(200)) and not (inputs(209));
    layer0_outputs(3448) <= inputs(202);
    layer0_outputs(3449) <= not(inputs(131));
    layer0_outputs(3450) <= (inputs(150)) or (inputs(84));
    layer0_outputs(3451) <= (inputs(5)) xor (inputs(163));
    layer0_outputs(3452) <= inputs(171);
    layer0_outputs(3453) <= inputs(40);
    layer0_outputs(3454) <= not((inputs(96)) xor (inputs(57)));
    layer0_outputs(3455) <= not(inputs(164)) or (inputs(231));
    layer0_outputs(3456) <= not((inputs(204)) xor (inputs(232)));
    layer0_outputs(3457) <= '0';
    layer0_outputs(3458) <= not((inputs(0)) and (inputs(17)));
    layer0_outputs(3459) <= not(inputs(230));
    layer0_outputs(3460) <= not((inputs(128)) or (inputs(167)));
    layer0_outputs(3461) <= not(inputs(85)) or (inputs(64));
    layer0_outputs(3462) <= not(inputs(120)) or (inputs(141));
    layer0_outputs(3463) <= inputs(138);
    layer0_outputs(3464) <= inputs(168);
    layer0_outputs(3465) <= inputs(181);
    layer0_outputs(3466) <= (inputs(206)) or (inputs(48));
    layer0_outputs(3467) <= not((inputs(94)) and (inputs(239)));
    layer0_outputs(3468) <= (inputs(162)) xor (inputs(81));
    layer0_outputs(3469) <= not(inputs(85));
    layer0_outputs(3470) <= not((inputs(35)) xor (inputs(89)));
    layer0_outputs(3471) <= (inputs(184)) xor (inputs(76));
    layer0_outputs(3472) <= not((inputs(182)) xor (inputs(106)));
    layer0_outputs(3473) <= (inputs(228)) xor (inputs(102));
    layer0_outputs(3474) <= not((inputs(9)) and (inputs(109)));
    layer0_outputs(3475) <= not((inputs(38)) or (inputs(212)));
    layer0_outputs(3476) <= not(inputs(157)) or (inputs(178));
    layer0_outputs(3477) <= not(inputs(56));
    layer0_outputs(3478) <= '0';
    layer0_outputs(3479) <= not(inputs(195));
    layer0_outputs(3480) <= (inputs(54)) and (inputs(56));
    layer0_outputs(3481) <= inputs(87);
    layer0_outputs(3482) <= (inputs(50)) and (inputs(65));
    layer0_outputs(3483) <= not((inputs(202)) or (inputs(93)));
    layer0_outputs(3484) <= not((inputs(98)) xor (inputs(30)));
    layer0_outputs(3485) <= not((inputs(7)) or (inputs(253)));
    layer0_outputs(3486) <= not((inputs(82)) xor (inputs(104)));
    layer0_outputs(3487) <= not((inputs(134)) or (inputs(149)));
    layer0_outputs(3488) <= inputs(32);
    layer0_outputs(3489) <= not((inputs(96)) xor (inputs(161)));
    layer0_outputs(3490) <= not((inputs(23)) or (inputs(98)));
    layer0_outputs(3491) <= (inputs(190)) and not (inputs(207));
    layer0_outputs(3492) <= (inputs(40)) and not (inputs(242));
    layer0_outputs(3493) <= inputs(200);
    layer0_outputs(3494) <= not((inputs(6)) xor (inputs(26)));
    layer0_outputs(3495) <= not(inputs(166));
    layer0_outputs(3496) <= inputs(39);
    layer0_outputs(3497) <= not((inputs(74)) or (inputs(6)));
    layer0_outputs(3498) <= not((inputs(3)) xor (inputs(171)));
    layer0_outputs(3499) <= not(inputs(8));
    layer0_outputs(3500) <= (inputs(111)) and (inputs(16));
    layer0_outputs(3501) <= not(inputs(200)) or (inputs(38));
    layer0_outputs(3502) <= not((inputs(217)) or (inputs(105)));
    layer0_outputs(3503) <= not(inputs(126));
    layer0_outputs(3504) <= inputs(52);
    layer0_outputs(3505) <= not(inputs(168));
    layer0_outputs(3506) <= (inputs(245)) and (inputs(48));
    layer0_outputs(3507) <= inputs(63);
    layer0_outputs(3508) <= '1';
    layer0_outputs(3509) <= (inputs(22)) or (inputs(200));
    layer0_outputs(3510) <= not(inputs(87)) or (inputs(62));
    layer0_outputs(3511) <= not(inputs(170)) or (inputs(207));
    layer0_outputs(3512) <= (inputs(121)) or (inputs(79));
    layer0_outputs(3513) <= not((inputs(135)) xor (inputs(36)));
    layer0_outputs(3514) <= (inputs(231)) or (inputs(69));
    layer0_outputs(3515) <= not(inputs(116));
    layer0_outputs(3516) <= (inputs(170)) and not (inputs(210));
    layer0_outputs(3517) <= inputs(124);
    layer0_outputs(3518) <= not(inputs(254)) or (inputs(236));
    layer0_outputs(3519) <= inputs(216);
    layer0_outputs(3520) <= inputs(156);
    layer0_outputs(3521) <= (inputs(18)) xor (inputs(181));
    layer0_outputs(3522) <= not((inputs(119)) xor (inputs(31)));
    layer0_outputs(3523) <= (inputs(132)) and not (inputs(21));
    layer0_outputs(3524) <= not(inputs(145)) or (inputs(236));
    layer0_outputs(3525) <= not(inputs(105)) or (inputs(83));
    layer0_outputs(3526) <= (inputs(139)) or (inputs(245));
    layer0_outputs(3527) <= not(inputs(203)) or (inputs(16));
    layer0_outputs(3528) <= (inputs(192)) and not (inputs(201));
    layer0_outputs(3529) <= not((inputs(176)) xor (inputs(147)));
    layer0_outputs(3530) <= inputs(199);
    layer0_outputs(3531) <= (inputs(120)) and not (inputs(84));
    layer0_outputs(3532) <= not((inputs(156)) or (inputs(7)));
    layer0_outputs(3533) <= (inputs(24)) xor (inputs(254));
    layer0_outputs(3534) <= not(inputs(150));
    layer0_outputs(3535) <= inputs(151);
    layer0_outputs(3536) <= inputs(165);
    layer0_outputs(3537) <= (inputs(58)) or (inputs(115));
    layer0_outputs(3538) <= inputs(144);
    layer0_outputs(3539) <= not((inputs(193)) and (inputs(15)));
    layer0_outputs(3540) <= not(inputs(165));
    layer0_outputs(3541) <= not((inputs(106)) xor (inputs(224)));
    layer0_outputs(3542) <= '0';
    layer0_outputs(3543) <= inputs(26);
    layer0_outputs(3544) <= (inputs(0)) and (inputs(250));
    layer0_outputs(3545) <= (inputs(176)) or (inputs(166));
    layer0_outputs(3546) <= inputs(81);
    layer0_outputs(3547) <= not((inputs(233)) and (inputs(109)));
    layer0_outputs(3548) <= (inputs(71)) or (inputs(229));
    layer0_outputs(3549) <= inputs(40);
    layer0_outputs(3550) <= (inputs(72)) and not (inputs(82));
    layer0_outputs(3551) <= not(inputs(161));
    layer0_outputs(3552) <= not((inputs(84)) xor (inputs(20)));
    layer0_outputs(3553) <= not(inputs(194)) or (inputs(143));
    layer0_outputs(3554) <= (inputs(113)) xor (inputs(246));
    layer0_outputs(3555) <= (inputs(121)) and not (inputs(167));
    layer0_outputs(3556) <= (inputs(83)) xor (inputs(64));
    layer0_outputs(3557) <= not(inputs(41)) or (inputs(46));
    layer0_outputs(3558) <= not(inputs(241)) or (inputs(147));
    layer0_outputs(3559) <= not(inputs(9)) or (inputs(136));
    layer0_outputs(3560) <= not(inputs(37)) or (inputs(237));
    layer0_outputs(3561) <= not((inputs(224)) xor (inputs(161)));
    layer0_outputs(3562) <= not(inputs(120));
    layer0_outputs(3563) <= not(inputs(191)) or (inputs(161));
    layer0_outputs(3564) <= not((inputs(149)) xor (inputs(182)));
    layer0_outputs(3565) <= not((inputs(71)) or (inputs(231)));
    layer0_outputs(3566) <= not(inputs(171)) or (inputs(234));
    layer0_outputs(3567) <= not((inputs(244)) xor (inputs(80)));
    layer0_outputs(3568) <= not(inputs(152));
    layer0_outputs(3569) <= not(inputs(49));
    layer0_outputs(3570) <= not((inputs(122)) or (inputs(221)));
    layer0_outputs(3571) <= (inputs(125)) and not (inputs(129));
    layer0_outputs(3572) <= '0';
    layer0_outputs(3573) <= not(inputs(243)) or (inputs(32));
    layer0_outputs(3574) <= not((inputs(109)) or (inputs(109)));
    layer0_outputs(3575) <= (inputs(125)) xor (inputs(157));
    layer0_outputs(3576) <= not((inputs(122)) xor (inputs(59)));
    layer0_outputs(3577) <= (inputs(14)) xor (inputs(72));
    layer0_outputs(3578) <= inputs(165);
    layer0_outputs(3579) <= (inputs(74)) or (inputs(146));
    layer0_outputs(3580) <= not((inputs(148)) or (inputs(117)));
    layer0_outputs(3581) <= (inputs(25)) and not (inputs(157));
    layer0_outputs(3582) <= (inputs(54)) and not (inputs(124));
    layer0_outputs(3583) <= not((inputs(113)) or (inputs(164)));
    layer0_outputs(3584) <= (inputs(27)) and (inputs(245));
    layer0_outputs(3585) <= (inputs(186)) xor (inputs(2));
    layer0_outputs(3586) <= not((inputs(183)) or (inputs(27)));
    layer0_outputs(3587) <= (inputs(192)) xor (inputs(1));
    layer0_outputs(3588) <= (inputs(71)) xor (inputs(246));
    layer0_outputs(3589) <= not((inputs(160)) xor (inputs(68)));
    layer0_outputs(3590) <= inputs(96);
    layer0_outputs(3591) <= not(inputs(97));
    layer0_outputs(3592) <= (inputs(88)) and not (inputs(210));
    layer0_outputs(3593) <= (inputs(2)) or (inputs(77));
    layer0_outputs(3594) <= inputs(187);
    layer0_outputs(3595) <= not(inputs(105));
    layer0_outputs(3596) <= not(inputs(91)) or (inputs(175));
    layer0_outputs(3597) <= not((inputs(182)) xor (inputs(227)));
    layer0_outputs(3598) <= not(inputs(57));
    layer0_outputs(3599) <= (inputs(223)) xor (inputs(78));
    layer0_outputs(3600) <= not(inputs(60)) or (inputs(65));
    layer0_outputs(3601) <= (inputs(125)) or (inputs(130));
    layer0_outputs(3602) <= inputs(107);
    layer0_outputs(3603) <= (inputs(30)) and not (inputs(147));
    layer0_outputs(3604) <= (inputs(30)) or (inputs(126));
    layer0_outputs(3605) <= not((inputs(99)) xor (inputs(208)));
    layer0_outputs(3606) <= inputs(223);
    layer0_outputs(3607) <= (inputs(41)) and not (inputs(47));
    layer0_outputs(3608) <= (inputs(204)) and not (inputs(21));
    layer0_outputs(3609) <= not((inputs(184)) or (inputs(189)));
    layer0_outputs(3610) <= not((inputs(103)) or (inputs(29)));
    layer0_outputs(3611) <= not((inputs(114)) xor (inputs(211)));
    layer0_outputs(3612) <= not(inputs(170)) or (inputs(66));
    layer0_outputs(3613) <= (inputs(155)) xor (inputs(233));
    layer0_outputs(3614) <= inputs(53);
    layer0_outputs(3615) <= not((inputs(218)) or (inputs(91)));
    layer0_outputs(3616) <= not(inputs(26));
    layer0_outputs(3617) <= not((inputs(241)) or (inputs(75)));
    layer0_outputs(3618) <= not(inputs(132)) or (inputs(224));
    layer0_outputs(3619) <= not((inputs(139)) or (inputs(62)));
    layer0_outputs(3620) <= (inputs(1)) or (inputs(116));
    layer0_outputs(3621) <= not((inputs(200)) or (inputs(231)));
    layer0_outputs(3622) <= (inputs(41)) xor (inputs(13));
    layer0_outputs(3623) <= (inputs(183)) and not (inputs(89));
    layer0_outputs(3624) <= inputs(11);
    layer0_outputs(3625) <= not((inputs(196)) xor (inputs(92)));
    layer0_outputs(3626) <= (inputs(218)) and not (inputs(22));
    layer0_outputs(3627) <= not((inputs(119)) xor (inputs(26)));
    layer0_outputs(3628) <= not(inputs(137)) or (inputs(93));
    layer0_outputs(3629) <= not((inputs(175)) and (inputs(243)));
    layer0_outputs(3630) <= not(inputs(93));
    layer0_outputs(3631) <= (inputs(198)) xor (inputs(166));
    layer0_outputs(3632) <= (inputs(138)) and not (inputs(187));
    layer0_outputs(3633) <= '1';
    layer0_outputs(3634) <= (inputs(128)) xor (inputs(167));
    layer0_outputs(3635) <= '1';
    layer0_outputs(3636) <= not((inputs(21)) xor (inputs(253)));
    layer0_outputs(3637) <= (inputs(28)) or (inputs(79));
    layer0_outputs(3638) <= not(inputs(33));
    layer0_outputs(3639) <= not((inputs(41)) or (inputs(248)));
    layer0_outputs(3640) <= not(inputs(44)) or (inputs(6));
    layer0_outputs(3641) <= not(inputs(183));
    layer0_outputs(3642) <= not(inputs(59)) or (inputs(60));
    layer0_outputs(3643) <= not(inputs(91));
    layer0_outputs(3644) <= (inputs(162)) xor (inputs(68));
    layer0_outputs(3645) <= not(inputs(31)) or (inputs(126));
    layer0_outputs(3646) <= (inputs(242)) and not (inputs(189));
    layer0_outputs(3647) <= (inputs(109)) and not (inputs(145));
    layer0_outputs(3648) <= (inputs(199)) and not (inputs(238));
    layer0_outputs(3649) <= (inputs(250)) and not (inputs(81));
    layer0_outputs(3650) <= (inputs(26)) xor (inputs(2));
    layer0_outputs(3651) <= not((inputs(24)) and (inputs(247)));
    layer0_outputs(3652) <= not((inputs(1)) or (inputs(62)));
    layer0_outputs(3653) <= not((inputs(140)) xor (inputs(138)));
    layer0_outputs(3654) <= not(inputs(253)) or (inputs(18));
    layer0_outputs(3655) <= (inputs(39)) and not (inputs(6));
    layer0_outputs(3656) <= not(inputs(17)) or (inputs(195));
    layer0_outputs(3657) <= not((inputs(110)) or (inputs(38)));
    layer0_outputs(3658) <= not(inputs(149));
    layer0_outputs(3659) <= not((inputs(186)) xor (inputs(138)));
    layer0_outputs(3660) <= not(inputs(187));
    layer0_outputs(3661) <= inputs(94);
    layer0_outputs(3662) <= inputs(117);
    layer0_outputs(3663) <= inputs(184);
    layer0_outputs(3664) <= not(inputs(216));
    layer0_outputs(3665) <= not(inputs(15));
    layer0_outputs(3666) <= not((inputs(8)) and (inputs(193)));
    layer0_outputs(3667) <= not(inputs(160));
    layer0_outputs(3668) <= (inputs(37)) and not (inputs(4));
    layer0_outputs(3669) <= not((inputs(55)) or (inputs(110)));
    layer0_outputs(3670) <= inputs(39);
    layer0_outputs(3671) <= not(inputs(234));
    layer0_outputs(3672) <= (inputs(26)) xor (inputs(124));
    layer0_outputs(3673) <= '0';
    layer0_outputs(3674) <= '0';
    layer0_outputs(3675) <= not(inputs(124)) or (inputs(169));
    layer0_outputs(3676) <= not((inputs(164)) or (inputs(141)));
    layer0_outputs(3677) <= (inputs(139)) and not (inputs(0));
    layer0_outputs(3678) <= inputs(106);
    layer0_outputs(3679) <= not(inputs(69)) or (inputs(227));
    layer0_outputs(3680) <= (inputs(75)) xor (inputs(77));
    layer0_outputs(3681) <= (inputs(124)) and not (inputs(62));
    layer0_outputs(3682) <= not((inputs(63)) and (inputs(177)));
    layer0_outputs(3683) <= inputs(129);
    layer0_outputs(3684) <= (inputs(211)) or (inputs(177));
    layer0_outputs(3685) <= (inputs(21)) and not (inputs(176));
    layer0_outputs(3686) <= not(inputs(72)) or (inputs(97));
    layer0_outputs(3687) <= not(inputs(17)) or (inputs(1));
    layer0_outputs(3688) <= (inputs(180)) and not (inputs(25));
    layer0_outputs(3689) <= (inputs(127)) or (inputs(45));
    layer0_outputs(3690) <= not((inputs(71)) or (inputs(248)));
    layer0_outputs(3691) <= (inputs(155)) and not (inputs(82));
    layer0_outputs(3692) <= not(inputs(218));
    layer0_outputs(3693) <= not((inputs(170)) or (inputs(116)));
    layer0_outputs(3694) <= (inputs(186)) and not (inputs(247));
    layer0_outputs(3695) <= (inputs(183)) and not (inputs(2));
    layer0_outputs(3696) <= not(inputs(40)) or (inputs(206));
    layer0_outputs(3697) <= not(inputs(1));
    layer0_outputs(3698) <= (inputs(14)) and not (inputs(238));
    layer0_outputs(3699) <= not((inputs(246)) and (inputs(179)));
    layer0_outputs(3700) <= '0';
    layer0_outputs(3701) <= not((inputs(71)) xor (inputs(168)));
    layer0_outputs(3702) <= '1';
    layer0_outputs(3703) <= (inputs(213)) and not (inputs(27));
    layer0_outputs(3704) <= (inputs(88)) xor (inputs(79));
    layer0_outputs(3705) <= not(inputs(196));
    layer0_outputs(3706) <= inputs(176);
    layer0_outputs(3707) <= not(inputs(162)) or (inputs(13));
    layer0_outputs(3708) <= (inputs(33)) and (inputs(34));
    layer0_outputs(3709) <= (inputs(170)) xor (inputs(31));
    layer0_outputs(3710) <= not(inputs(169));
    layer0_outputs(3711) <= not((inputs(250)) or (inputs(207)));
    layer0_outputs(3712) <= not(inputs(157)) or (inputs(25));
    layer0_outputs(3713) <= (inputs(182)) and not (inputs(48));
    layer0_outputs(3714) <= not(inputs(170));
    layer0_outputs(3715) <= '1';
    layer0_outputs(3716) <= not(inputs(213)) or (inputs(229));
    layer0_outputs(3717) <= (inputs(104)) xor (inputs(57));
    layer0_outputs(3718) <= not((inputs(180)) or (inputs(109)));
    layer0_outputs(3719) <= not(inputs(170)) or (inputs(99));
    layer0_outputs(3720) <= not(inputs(117));
    layer0_outputs(3721) <= (inputs(241)) or (inputs(212));
    layer0_outputs(3722) <= not(inputs(78));
    layer0_outputs(3723) <= (inputs(237)) xor (inputs(84));
    layer0_outputs(3724) <= inputs(192);
    layer0_outputs(3725) <= inputs(143);
    layer0_outputs(3726) <= (inputs(26)) and (inputs(230));
    layer0_outputs(3727) <= not(inputs(150));
    layer0_outputs(3728) <= not(inputs(179)) or (inputs(47));
    layer0_outputs(3729) <= not((inputs(81)) or (inputs(78)));
    layer0_outputs(3730) <= not(inputs(66));
    layer0_outputs(3731) <= (inputs(120)) and not (inputs(173));
    layer0_outputs(3732) <= not((inputs(254)) or (inputs(142)));
    layer0_outputs(3733) <= not((inputs(187)) or (inputs(186)));
    layer0_outputs(3734) <= not(inputs(57)) or (inputs(25));
    layer0_outputs(3735) <= not(inputs(20)) or (inputs(113));
    layer0_outputs(3736) <= inputs(237);
    layer0_outputs(3737) <= not(inputs(179));
    layer0_outputs(3738) <= not((inputs(141)) or (inputs(90)));
    layer0_outputs(3739) <= (inputs(211)) and not (inputs(130));
    layer0_outputs(3740) <= (inputs(172)) xor (inputs(26));
    layer0_outputs(3741) <= not((inputs(33)) or (inputs(231)));
    layer0_outputs(3742) <= not((inputs(188)) and (inputs(157)));
    layer0_outputs(3743) <= not((inputs(7)) xor (inputs(188)));
    layer0_outputs(3744) <= (inputs(194)) and not (inputs(115));
    layer0_outputs(3745) <= inputs(71);
    layer0_outputs(3746) <= (inputs(224)) and not (inputs(226));
    layer0_outputs(3747) <= not(inputs(114)) or (inputs(4));
    layer0_outputs(3748) <= inputs(40);
    layer0_outputs(3749) <= not(inputs(153));
    layer0_outputs(3750) <= not(inputs(228));
    layer0_outputs(3751) <= inputs(167);
    layer0_outputs(3752) <= not((inputs(160)) xor (inputs(15)));
    layer0_outputs(3753) <= not(inputs(74)) or (inputs(46));
    layer0_outputs(3754) <= not(inputs(234)) or (inputs(75));
    layer0_outputs(3755) <= (inputs(161)) and not (inputs(193));
    layer0_outputs(3756) <= '0';
    layer0_outputs(3757) <= not(inputs(206));
    layer0_outputs(3758) <= not((inputs(114)) xor (inputs(230)));
    layer0_outputs(3759) <= inputs(165);
    layer0_outputs(3760) <= inputs(156);
    layer0_outputs(3761) <= not((inputs(144)) or (inputs(232)));
    layer0_outputs(3762) <= (inputs(59)) or (inputs(200));
    layer0_outputs(3763) <= not(inputs(202)) or (inputs(27));
    layer0_outputs(3764) <= not(inputs(53)) or (inputs(127));
    layer0_outputs(3765) <= (inputs(201)) xor (inputs(111));
    layer0_outputs(3766) <= (inputs(93)) xor (inputs(65));
    layer0_outputs(3767) <= inputs(124);
    layer0_outputs(3768) <= not(inputs(88));
    layer0_outputs(3769) <= not((inputs(75)) or (inputs(189)));
    layer0_outputs(3770) <= not(inputs(148));
    layer0_outputs(3771) <= inputs(79);
    layer0_outputs(3772) <= inputs(217);
    layer0_outputs(3773) <= not((inputs(216)) xor (inputs(253)));
    layer0_outputs(3774) <= (inputs(45)) xor (inputs(78));
    layer0_outputs(3775) <= not(inputs(194));
    layer0_outputs(3776) <= (inputs(18)) and not (inputs(13));
    layer0_outputs(3777) <= not((inputs(119)) or (inputs(244)));
    layer0_outputs(3778) <= (inputs(181)) xor (inputs(63));
    layer0_outputs(3779) <= not((inputs(20)) xor (inputs(43)));
    layer0_outputs(3780) <= not((inputs(114)) xor (inputs(64)));
    layer0_outputs(3781) <= (inputs(78)) or (inputs(78));
    layer0_outputs(3782) <= (inputs(3)) or (inputs(7));
    layer0_outputs(3783) <= not((inputs(252)) xor (inputs(122)));
    layer0_outputs(3784) <= not(inputs(89)) or (inputs(195));
    layer0_outputs(3785) <= not(inputs(55)) or (inputs(178));
    layer0_outputs(3786) <= inputs(109);
    layer0_outputs(3787) <= (inputs(140)) and (inputs(216));
    layer0_outputs(3788) <= (inputs(206)) and not (inputs(192));
    layer0_outputs(3789) <= not((inputs(111)) or (inputs(29)));
    layer0_outputs(3790) <= (inputs(162)) or (inputs(146));
    layer0_outputs(3791) <= not(inputs(73));
    layer0_outputs(3792) <= not((inputs(109)) or (inputs(213)));
    layer0_outputs(3793) <= (inputs(5)) xor (inputs(64));
    layer0_outputs(3794) <= not((inputs(99)) xor (inputs(160)));
    layer0_outputs(3795) <= not((inputs(139)) or (inputs(196)));
    layer0_outputs(3796) <= not(inputs(91)) or (inputs(205));
    layer0_outputs(3797) <= not((inputs(12)) xor (inputs(211)));
    layer0_outputs(3798) <= (inputs(152)) and not (inputs(226));
    layer0_outputs(3799) <= not(inputs(11)) or (inputs(174));
    layer0_outputs(3800) <= inputs(172);
    layer0_outputs(3801) <= (inputs(158)) or (inputs(164));
    layer0_outputs(3802) <= not((inputs(93)) xor (inputs(3)));
    layer0_outputs(3803) <= (inputs(125)) or (inputs(47));
    layer0_outputs(3804) <= '1';
    layer0_outputs(3805) <= inputs(148);
    layer0_outputs(3806) <= '0';
    layer0_outputs(3807) <= not(inputs(42)) or (inputs(47));
    layer0_outputs(3808) <= (inputs(152)) and not (inputs(176));
    layer0_outputs(3809) <= not((inputs(230)) xor (inputs(49)));
    layer0_outputs(3810) <= not((inputs(60)) or (inputs(6)));
    layer0_outputs(3811) <= not(inputs(151)) or (inputs(70));
    layer0_outputs(3812) <= not((inputs(212)) or (inputs(232)));
    layer0_outputs(3813) <= (inputs(180)) xor (inputs(28));
    layer0_outputs(3814) <= (inputs(14)) or (inputs(189));
    layer0_outputs(3815) <= (inputs(130)) xor (inputs(249));
    layer0_outputs(3816) <= not((inputs(78)) and (inputs(147)));
    layer0_outputs(3817) <= (inputs(229)) or (inputs(228));
    layer0_outputs(3818) <= not(inputs(243)) or (inputs(50));
    layer0_outputs(3819) <= not(inputs(138));
    layer0_outputs(3820) <= (inputs(22)) xor (inputs(130));
    layer0_outputs(3821) <= inputs(60);
    layer0_outputs(3822) <= (inputs(201)) and not (inputs(22));
    layer0_outputs(3823) <= (inputs(7)) or (inputs(55));
    layer0_outputs(3824) <= '0';
    layer0_outputs(3825) <= not(inputs(134));
    layer0_outputs(3826) <= not(inputs(47));
    layer0_outputs(3827) <= not(inputs(191)) or (inputs(127));
    layer0_outputs(3828) <= not((inputs(45)) xor (inputs(76)));
    layer0_outputs(3829) <= '0';
    layer0_outputs(3830) <= not((inputs(56)) xor (inputs(111)));
    layer0_outputs(3831) <= not((inputs(51)) and (inputs(143)));
    layer0_outputs(3832) <= (inputs(130)) or (inputs(39));
    layer0_outputs(3833) <= not(inputs(137));
    layer0_outputs(3834) <= not(inputs(116));
    layer0_outputs(3835) <= (inputs(59)) or (inputs(115));
    layer0_outputs(3836) <= not((inputs(240)) or (inputs(180)));
    layer0_outputs(3837) <= (inputs(102)) xor (inputs(84));
    layer0_outputs(3838) <= not(inputs(78)) or (inputs(96));
    layer0_outputs(3839) <= not((inputs(122)) or (inputs(229)));
    layer0_outputs(3840) <= not(inputs(167)) or (inputs(196));
    layer0_outputs(3841) <= not(inputs(13));
    layer0_outputs(3842) <= inputs(196);
    layer0_outputs(3843) <= (inputs(210)) or (inputs(194));
    layer0_outputs(3844) <= not((inputs(226)) xor (inputs(90)));
    layer0_outputs(3845) <= (inputs(181)) xor (inputs(220));
    layer0_outputs(3846) <= not(inputs(74));
    layer0_outputs(3847) <= not((inputs(47)) or (inputs(142)));
    layer0_outputs(3848) <= not(inputs(138)) or (inputs(62));
    layer0_outputs(3849) <= inputs(160);
    layer0_outputs(3850) <= not(inputs(32));
    layer0_outputs(3851) <= inputs(239);
    layer0_outputs(3852) <= inputs(187);
    layer0_outputs(3853) <= (inputs(240)) or (inputs(11));
    layer0_outputs(3854) <= (inputs(240)) or (inputs(161));
    layer0_outputs(3855) <= (inputs(171)) and not (inputs(204));
    layer0_outputs(3856) <= not(inputs(247));
    layer0_outputs(3857) <= not((inputs(118)) and (inputs(135)));
    layer0_outputs(3858) <= (inputs(12)) and not (inputs(156));
    layer0_outputs(3859) <= (inputs(225)) xor (inputs(92));
    layer0_outputs(3860) <= not(inputs(204)) or (inputs(119));
    layer0_outputs(3861) <= not(inputs(71));
    layer0_outputs(3862) <= (inputs(205)) or (inputs(71));
    layer0_outputs(3863) <= not((inputs(163)) or (inputs(53)));
    layer0_outputs(3864) <= not(inputs(137));
    layer0_outputs(3865) <= (inputs(70)) or (inputs(32));
    layer0_outputs(3866) <= (inputs(154)) xor (inputs(158));
    layer0_outputs(3867) <= not(inputs(64));
    layer0_outputs(3868) <= inputs(28);
    layer0_outputs(3869) <= not((inputs(161)) xor (inputs(140)));
    layer0_outputs(3870) <= not(inputs(133)) or (inputs(129));
    layer0_outputs(3871) <= inputs(247);
    layer0_outputs(3872) <= (inputs(140)) and not (inputs(97));
    layer0_outputs(3873) <= (inputs(244)) xor (inputs(202));
    layer0_outputs(3874) <= (inputs(251)) and not (inputs(110));
    layer0_outputs(3875) <= not(inputs(78)) or (inputs(192));
    layer0_outputs(3876) <= (inputs(157)) and not (inputs(177));
    layer0_outputs(3877) <= not((inputs(174)) xor (inputs(241)));
    layer0_outputs(3878) <= '1';
    layer0_outputs(3879) <= (inputs(53)) and not (inputs(17));
    layer0_outputs(3880) <= (inputs(6)) and not (inputs(62));
    layer0_outputs(3881) <= (inputs(145)) and (inputs(255));
    layer0_outputs(3882) <= not((inputs(32)) or (inputs(235)));
    layer0_outputs(3883) <= not((inputs(195)) and (inputs(106)));
    layer0_outputs(3884) <= (inputs(186)) or (inputs(109));
    layer0_outputs(3885) <= (inputs(240)) and not (inputs(95));
    layer0_outputs(3886) <= '0';
    layer0_outputs(3887) <= '0';
    layer0_outputs(3888) <= not(inputs(103)) or (inputs(18));
    layer0_outputs(3889) <= inputs(116);
    layer0_outputs(3890) <= not((inputs(164)) or (inputs(139)));
    layer0_outputs(3891) <= not((inputs(78)) or (inputs(92)));
    layer0_outputs(3892) <= not(inputs(136)) or (inputs(85));
    layer0_outputs(3893) <= not(inputs(172));
    layer0_outputs(3894) <= (inputs(47)) or (inputs(181));
    layer0_outputs(3895) <= not((inputs(55)) xor (inputs(33)));
    layer0_outputs(3896) <= inputs(175);
    layer0_outputs(3897) <= (inputs(149)) or (inputs(80));
    layer0_outputs(3898) <= not(inputs(122)) or (inputs(87));
    layer0_outputs(3899) <= not(inputs(225));
    layer0_outputs(3900) <= not((inputs(69)) xor (inputs(84)));
    layer0_outputs(3901) <= '1';
    layer0_outputs(3902) <= (inputs(52)) or (inputs(183));
    layer0_outputs(3903) <= not((inputs(2)) or (inputs(133)));
    layer0_outputs(3904) <= not(inputs(195));
    layer0_outputs(3905) <= (inputs(136)) and not (inputs(156));
    layer0_outputs(3906) <= inputs(87);
    layer0_outputs(3907) <= (inputs(103)) and not (inputs(39));
    layer0_outputs(3908) <= (inputs(189)) or (inputs(52));
    layer0_outputs(3909) <= (inputs(56)) xor (inputs(115));
    layer0_outputs(3910) <= (inputs(7)) xor (inputs(130));
    layer0_outputs(3911) <= inputs(132);
    layer0_outputs(3912) <= not(inputs(254));
    layer0_outputs(3913) <= not(inputs(132)) or (inputs(97));
    layer0_outputs(3914) <= not((inputs(216)) or (inputs(111)));
    layer0_outputs(3915) <= not(inputs(28)) or (inputs(66));
    layer0_outputs(3916) <= inputs(177);
    layer0_outputs(3917) <= (inputs(51)) and not (inputs(114));
    layer0_outputs(3918) <= not((inputs(181)) xor (inputs(224)));
    layer0_outputs(3919) <= not(inputs(86)) or (inputs(83));
    layer0_outputs(3920) <= not(inputs(121));
    layer0_outputs(3921) <= inputs(16);
    layer0_outputs(3922) <= inputs(133);
    layer0_outputs(3923) <= (inputs(185)) and not (inputs(98));
    layer0_outputs(3924) <= (inputs(107)) or (inputs(168));
    layer0_outputs(3925) <= (inputs(213)) xor (inputs(69));
    layer0_outputs(3926) <= not(inputs(208));
    layer0_outputs(3927) <= not((inputs(16)) or (inputs(138)));
    layer0_outputs(3928) <= not((inputs(141)) or (inputs(61)));
    layer0_outputs(3929) <= not(inputs(221));
    layer0_outputs(3930) <= (inputs(142)) or (inputs(164));
    layer0_outputs(3931) <= not((inputs(149)) or (inputs(67)));
    layer0_outputs(3932) <= not(inputs(56));
    layer0_outputs(3933) <= not(inputs(117)) or (inputs(177));
    layer0_outputs(3934) <= (inputs(5)) xor (inputs(198));
    layer0_outputs(3935) <= not((inputs(172)) xor (inputs(201)));
    layer0_outputs(3936) <= not((inputs(250)) or (inputs(60)));
    layer0_outputs(3937) <= (inputs(124)) or (inputs(97));
    layer0_outputs(3938) <= not(inputs(211)) or (inputs(26));
    layer0_outputs(3939) <= not((inputs(41)) or (inputs(32)));
    layer0_outputs(3940) <= not((inputs(104)) xor (inputs(252)));
    layer0_outputs(3941) <= not((inputs(103)) and (inputs(50)));
    layer0_outputs(3942) <= inputs(52);
    layer0_outputs(3943) <= (inputs(63)) or (inputs(43));
    layer0_outputs(3944) <= not(inputs(136));
    layer0_outputs(3945) <= (inputs(98)) or (inputs(80));
    layer0_outputs(3946) <= inputs(218);
    layer0_outputs(3947) <= not(inputs(176)) or (inputs(43));
    layer0_outputs(3948) <= not(inputs(150));
    layer0_outputs(3949) <= inputs(139);
    layer0_outputs(3950) <= not((inputs(240)) xor (inputs(194)));
    layer0_outputs(3951) <= inputs(131);
    layer0_outputs(3952) <= not((inputs(103)) or (inputs(84)));
    layer0_outputs(3953) <= (inputs(196)) xor (inputs(82));
    layer0_outputs(3954) <= not(inputs(67)) or (inputs(249));
    layer0_outputs(3955) <= not((inputs(212)) xor (inputs(36)));
    layer0_outputs(3956) <= inputs(235);
    layer0_outputs(3957) <= (inputs(113)) and not (inputs(178));
    layer0_outputs(3958) <= (inputs(188)) and not (inputs(254));
    layer0_outputs(3959) <= not((inputs(139)) xor (inputs(99)));
    layer0_outputs(3960) <= (inputs(83)) and (inputs(86));
    layer0_outputs(3961) <= (inputs(78)) or (inputs(101));
    layer0_outputs(3962) <= not(inputs(150)) or (inputs(19));
    layer0_outputs(3963) <= (inputs(106)) and not (inputs(161));
    layer0_outputs(3964) <= not(inputs(44));
    layer0_outputs(3965) <= inputs(178);
    layer0_outputs(3966) <= inputs(227);
    layer0_outputs(3967) <= inputs(212);
    layer0_outputs(3968) <= not(inputs(179));
    layer0_outputs(3969) <= (inputs(55)) or (inputs(254));
    layer0_outputs(3970) <= not((inputs(84)) xor (inputs(203)));
    layer0_outputs(3971) <= (inputs(230)) and not (inputs(157));
    layer0_outputs(3972) <= not((inputs(122)) or (inputs(145)));
    layer0_outputs(3973) <= (inputs(220)) or (inputs(202));
    layer0_outputs(3974) <= not((inputs(33)) or (inputs(188)));
    layer0_outputs(3975) <= not(inputs(178));
    layer0_outputs(3976) <= (inputs(121)) or (inputs(54));
    layer0_outputs(3977) <= (inputs(189)) or (inputs(116));
    layer0_outputs(3978) <= not((inputs(55)) or (inputs(12)));
    layer0_outputs(3979) <= inputs(132);
    layer0_outputs(3980) <= not(inputs(27));
    layer0_outputs(3981) <= not((inputs(111)) or (inputs(208)));
    layer0_outputs(3982) <= not(inputs(42)) or (inputs(224));
    layer0_outputs(3983) <= not((inputs(13)) or (inputs(176)));
    layer0_outputs(3984) <= (inputs(126)) or (inputs(163));
    layer0_outputs(3985) <= (inputs(3)) xor (inputs(119));
    layer0_outputs(3986) <= not(inputs(163));
    layer0_outputs(3987) <= (inputs(117)) or (inputs(131));
    layer0_outputs(3988) <= not(inputs(132));
    layer0_outputs(3989) <= (inputs(113)) or (inputs(111));
    layer0_outputs(3990) <= (inputs(213)) xor (inputs(39));
    layer0_outputs(3991) <= inputs(162);
    layer0_outputs(3992) <= (inputs(235)) and not (inputs(79));
    layer0_outputs(3993) <= (inputs(115)) and not (inputs(246));
    layer0_outputs(3994) <= (inputs(123)) xor (inputs(146));
    layer0_outputs(3995) <= (inputs(196)) and not (inputs(85));
    layer0_outputs(3996) <= (inputs(48)) and not (inputs(114));
    layer0_outputs(3997) <= (inputs(39)) xor (inputs(200));
    layer0_outputs(3998) <= not(inputs(216));
    layer0_outputs(3999) <= (inputs(26)) xor (inputs(4));
    layer0_outputs(4000) <= inputs(124);
    layer0_outputs(4001) <= inputs(203);
    layer0_outputs(4002) <= (inputs(215)) and not (inputs(108));
    layer0_outputs(4003) <= inputs(139);
    layer0_outputs(4004) <= '0';
    layer0_outputs(4005) <= not(inputs(203));
    layer0_outputs(4006) <= '1';
    layer0_outputs(4007) <= (inputs(139)) and not (inputs(205));
    layer0_outputs(4008) <= not((inputs(56)) or (inputs(146)));
    layer0_outputs(4009) <= not(inputs(194));
    layer0_outputs(4010) <= not((inputs(117)) or (inputs(62)));
    layer0_outputs(4011) <= not((inputs(88)) or (inputs(253)));
    layer0_outputs(4012) <= '1';
    layer0_outputs(4013) <= (inputs(182)) or (inputs(209));
    layer0_outputs(4014) <= not(inputs(165)) or (inputs(140));
    layer0_outputs(4015) <= not(inputs(89));
    layer0_outputs(4016) <= not(inputs(198)) or (inputs(9));
    layer0_outputs(4017) <= not(inputs(32)) or (inputs(99));
    layer0_outputs(4018) <= inputs(224);
    layer0_outputs(4019) <= not(inputs(182));
    layer0_outputs(4020) <= (inputs(178)) or (inputs(120));
    layer0_outputs(4021) <= (inputs(240)) or (inputs(162));
    layer0_outputs(4022) <= (inputs(146)) or (inputs(26));
    layer0_outputs(4023) <= inputs(131);
    layer0_outputs(4024) <= not((inputs(215)) or (inputs(200)));
    layer0_outputs(4025) <= (inputs(177)) or (inputs(9));
    layer0_outputs(4026) <= not((inputs(148)) or (inputs(207)));
    layer0_outputs(4027) <= (inputs(147)) and not (inputs(95));
    layer0_outputs(4028) <= (inputs(131)) or (inputs(251));
    layer0_outputs(4029) <= (inputs(73)) and not (inputs(223));
    layer0_outputs(4030) <= (inputs(135)) and not (inputs(234));
    layer0_outputs(4031) <= not(inputs(123));
    layer0_outputs(4032) <= not(inputs(67));
    layer0_outputs(4033) <= not(inputs(147)) or (inputs(221));
    layer0_outputs(4034) <= (inputs(72)) and not (inputs(127));
    layer0_outputs(4035) <= not(inputs(218));
    layer0_outputs(4036) <= (inputs(98)) xor (inputs(147));
    layer0_outputs(4037) <= not((inputs(95)) xor (inputs(229)));
    layer0_outputs(4038) <= not(inputs(54));
    layer0_outputs(4039) <= inputs(51);
    layer0_outputs(4040) <= not(inputs(151));
    layer0_outputs(4041) <= not(inputs(227)) or (inputs(110));
    layer0_outputs(4042) <= (inputs(173)) or (inputs(116));
    layer0_outputs(4043) <= (inputs(230)) xor (inputs(177));
    layer0_outputs(4044) <= inputs(133);
    layer0_outputs(4045) <= not((inputs(35)) or (inputs(97)));
    layer0_outputs(4046) <= not(inputs(246));
    layer0_outputs(4047) <= (inputs(10)) or (inputs(62));
    layer0_outputs(4048) <= (inputs(55)) or (inputs(10));
    layer0_outputs(4049) <= inputs(62);
    layer0_outputs(4050) <= (inputs(158)) and not (inputs(82));
    layer0_outputs(4051) <= not((inputs(170)) or (inputs(35)));
    layer0_outputs(4052) <= not((inputs(223)) or (inputs(129)));
    layer0_outputs(4053) <= (inputs(197)) and not (inputs(115));
    layer0_outputs(4054) <= (inputs(79)) and (inputs(174));
    layer0_outputs(4055) <= (inputs(241)) and not (inputs(222));
    layer0_outputs(4056) <= (inputs(180)) xor (inputs(73));
    layer0_outputs(4057) <= not((inputs(66)) xor (inputs(74)));
    layer0_outputs(4058) <= not(inputs(68));
    layer0_outputs(4059) <= inputs(134);
    layer0_outputs(4060) <= (inputs(116)) and not (inputs(143));
    layer0_outputs(4061) <= inputs(119);
    layer0_outputs(4062) <= (inputs(15)) or (inputs(218));
    layer0_outputs(4063) <= not(inputs(71));
    layer0_outputs(4064) <= (inputs(71)) and not (inputs(119));
    layer0_outputs(4065) <= not((inputs(130)) or (inputs(227)));
    layer0_outputs(4066) <= not((inputs(211)) or (inputs(80)));
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= not((inputs(137)) or (inputs(221)));
    layer0_outputs(4069) <= not((inputs(173)) xor (inputs(79)));
    layer0_outputs(4070) <= not((inputs(171)) xor (inputs(64)));
    layer0_outputs(4071) <= (inputs(172)) or (inputs(75));
    layer0_outputs(4072) <= not(inputs(163)) or (inputs(28));
    layer0_outputs(4073) <= not((inputs(35)) xor (inputs(154)));
    layer0_outputs(4074) <= not(inputs(90)) or (inputs(159));
    layer0_outputs(4075) <= (inputs(127)) and not (inputs(137));
    layer0_outputs(4076) <= (inputs(253)) and not (inputs(112));
    layer0_outputs(4077) <= (inputs(88)) or (inputs(230));
    layer0_outputs(4078) <= not((inputs(247)) or (inputs(34)));
    layer0_outputs(4079) <= not(inputs(2));
    layer0_outputs(4080) <= (inputs(36)) and not (inputs(189));
    layer0_outputs(4081) <= not((inputs(167)) or (inputs(219)));
    layer0_outputs(4082) <= not((inputs(203)) xor (inputs(179)));
    layer0_outputs(4083) <= not(inputs(62)) or (inputs(173));
    layer0_outputs(4084) <= not(inputs(224));
    layer0_outputs(4085) <= '1';
    layer0_outputs(4086) <= not((inputs(111)) and (inputs(13)));
    layer0_outputs(4087) <= not((inputs(150)) xor (inputs(36)));
    layer0_outputs(4088) <= (inputs(156)) and not (inputs(210));
    layer0_outputs(4089) <= (inputs(74)) and not (inputs(34));
    layer0_outputs(4090) <= (inputs(82)) or (inputs(25));
    layer0_outputs(4091) <= (inputs(185)) or (inputs(23));
    layer0_outputs(4092) <= '0';
    layer0_outputs(4093) <= (inputs(91)) and not (inputs(230));
    layer0_outputs(4094) <= (inputs(192)) and not (inputs(19));
    layer0_outputs(4095) <= not(inputs(121));
    layer0_outputs(4096) <= (inputs(118)) and not (inputs(3));
    layer0_outputs(4097) <= not(inputs(136));
    layer0_outputs(4098) <= (inputs(105)) and (inputs(213));
    layer0_outputs(4099) <= not(inputs(21));
    layer0_outputs(4100) <= not((inputs(189)) or (inputs(51)));
    layer0_outputs(4101) <= inputs(121);
    layer0_outputs(4102) <= not((inputs(37)) xor (inputs(81)));
    layer0_outputs(4103) <= inputs(187);
    layer0_outputs(4104) <= (inputs(16)) and not (inputs(63));
    layer0_outputs(4105) <= inputs(214);
    layer0_outputs(4106) <= inputs(113);
    layer0_outputs(4107) <= not((inputs(164)) or (inputs(137)));
    layer0_outputs(4108) <= not((inputs(30)) or (inputs(129)));
    layer0_outputs(4109) <= not(inputs(213)) or (inputs(77));
    layer0_outputs(4110) <= not(inputs(7)) or (inputs(97));
    layer0_outputs(4111) <= (inputs(173)) xor (inputs(50));
    layer0_outputs(4112) <= (inputs(219)) or (inputs(110));
    layer0_outputs(4113) <= (inputs(37)) xor (inputs(169));
    layer0_outputs(4114) <= not((inputs(194)) or (inputs(35)));
    layer0_outputs(4115) <= (inputs(30)) xor (inputs(166));
    layer0_outputs(4116) <= (inputs(220)) and not (inputs(217));
    layer0_outputs(4117) <= (inputs(58)) or (inputs(94));
    layer0_outputs(4118) <= '0';
    layer0_outputs(4119) <= not(inputs(87));
    layer0_outputs(4120) <= not((inputs(149)) xor (inputs(240)));
    layer0_outputs(4121) <= inputs(214);
    layer0_outputs(4122) <= not(inputs(151));
    layer0_outputs(4123) <= (inputs(179)) and not (inputs(134));
    layer0_outputs(4124) <= not((inputs(167)) or (inputs(10)));
    layer0_outputs(4125) <= not(inputs(233)) or (inputs(176));
    layer0_outputs(4126) <= '0';
    layer0_outputs(4127) <= (inputs(42)) or (inputs(197));
    layer0_outputs(4128) <= inputs(92);
    layer0_outputs(4129) <= (inputs(250)) or (inputs(238));
    layer0_outputs(4130) <= not(inputs(142));
    layer0_outputs(4131) <= inputs(249);
    layer0_outputs(4132) <= not(inputs(136)) or (inputs(26));
    layer0_outputs(4133) <= (inputs(126)) or (inputs(48));
    layer0_outputs(4134) <= not((inputs(35)) xor (inputs(224)));
    layer0_outputs(4135) <= not(inputs(228));
    layer0_outputs(4136) <= (inputs(198)) and (inputs(200));
    layer0_outputs(4137) <= (inputs(3)) and (inputs(233));
    layer0_outputs(4138) <= not(inputs(163)) or (inputs(225));
    layer0_outputs(4139) <= (inputs(8)) or (inputs(217));
    layer0_outputs(4140) <= (inputs(57)) or (inputs(29));
    layer0_outputs(4141) <= '0';
    layer0_outputs(4142) <= (inputs(162)) and (inputs(112));
    layer0_outputs(4143) <= '0';
    layer0_outputs(4144) <= (inputs(32)) xor (inputs(198));
    layer0_outputs(4145) <= (inputs(139)) xor (inputs(10));
    layer0_outputs(4146) <= not((inputs(22)) xor (inputs(49)));
    layer0_outputs(4147) <= not(inputs(132));
    layer0_outputs(4148) <= (inputs(191)) xor (inputs(84));
    layer0_outputs(4149) <= inputs(83);
    layer0_outputs(4150) <= not(inputs(231));
    layer0_outputs(4151) <= (inputs(202)) or (inputs(70));
    layer0_outputs(4152) <= (inputs(242)) and (inputs(74));
    layer0_outputs(4153) <= not(inputs(77)) or (inputs(7));
    layer0_outputs(4154) <= inputs(217);
    layer0_outputs(4155) <= (inputs(147)) and not (inputs(201));
    layer0_outputs(4156) <= (inputs(88)) and not (inputs(206));
    layer0_outputs(4157) <= not(inputs(110));
    layer0_outputs(4158) <= not(inputs(49));
    layer0_outputs(4159) <= (inputs(138)) xor (inputs(255));
    layer0_outputs(4160) <= not((inputs(138)) xor (inputs(46)));
    layer0_outputs(4161) <= not(inputs(140));
    layer0_outputs(4162) <= not((inputs(95)) xor (inputs(118)));
    layer0_outputs(4163) <= not((inputs(254)) and (inputs(104)));
    layer0_outputs(4164) <= not(inputs(133)) or (inputs(110));
    layer0_outputs(4165) <= inputs(234);
    layer0_outputs(4166) <= (inputs(181)) xor (inputs(118));
    layer0_outputs(4167) <= (inputs(139)) and not (inputs(189));
    layer0_outputs(4168) <= not(inputs(9));
    layer0_outputs(4169) <= (inputs(53)) or (inputs(194));
    layer0_outputs(4170) <= (inputs(134)) and not (inputs(246));
    layer0_outputs(4171) <= not((inputs(210)) xor (inputs(157)));
    layer0_outputs(4172) <= (inputs(78)) xor (inputs(255));
    layer0_outputs(4173) <= (inputs(28)) xor (inputs(32));
    layer0_outputs(4174) <= inputs(210);
    layer0_outputs(4175) <= (inputs(147)) and not (inputs(111));
    layer0_outputs(4176) <= (inputs(91)) and not (inputs(21));
    layer0_outputs(4177) <= not(inputs(53));
    layer0_outputs(4178) <= (inputs(187)) and not (inputs(228));
    layer0_outputs(4179) <= (inputs(90)) or (inputs(157));
    layer0_outputs(4180) <= not(inputs(99));
    layer0_outputs(4181) <= (inputs(213)) and not (inputs(126));
    layer0_outputs(4182) <= inputs(45);
    layer0_outputs(4183) <= (inputs(137)) or (inputs(230));
    layer0_outputs(4184) <= (inputs(200)) xor (inputs(80));
    layer0_outputs(4185) <= (inputs(31)) and not (inputs(20));
    layer0_outputs(4186) <= not((inputs(194)) or (inputs(191)));
    layer0_outputs(4187) <= inputs(86);
    layer0_outputs(4188) <= not((inputs(116)) or (inputs(192)));
    layer0_outputs(4189) <= not((inputs(132)) or (inputs(170)));
    layer0_outputs(4190) <= (inputs(38)) xor (inputs(69));
    layer0_outputs(4191) <= not((inputs(160)) xor (inputs(203)));
    layer0_outputs(4192) <= not((inputs(52)) or (inputs(6)));
    layer0_outputs(4193) <= not((inputs(224)) or (inputs(59)));
    layer0_outputs(4194) <= '1';
    layer0_outputs(4195) <= not((inputs(86)) or (inputs(224)));
    layer0_outputs(4196) <= (inputs(216)) and not (inputs(126));
    layer0_outputs(4197) <= not(inputs(80)) or (inputs(27));
    layer0_outputs(4198) <= (inputs(57)) and not (inputs(48));
    layer0_outputs(4199) <= inputs(94);
    layer0_outputs(4200) <= not((inputs(139)) or (inputs(154)));
    layer0_outputs(4201) <= not(inputs(7)) or (inputs(36));
    layer0_outputs(4202) <= (inputs(154)) xor (inputs(147));
    layer0_outputs(4203) <= (inputs(14)) and (inputs(3));
    layer0_outputs(4204) <= not(inputs(138)) or (inputs(43));
    layer0_outputs(4205) <= (inputs(17)) or (inputs(111));
    layer0_outputs(4206) <= not((inputs(127)) and (inputs(51)));
    layer0_outputs(4207) <= (inputs(86)) and not (inputs(52));
    layer0_outputs(4208) <= (inputs(154)) and (inputs(101));
    layer0_outputs(4209) <= (inputs(122)) and not (inputs(243));
    layer0_outputs(4210) <= not(inputs(71));
    layer0_outputs(4211) <= inputs(136);
    layer0_outputs(4212) <= inputs(184);
    layer0_outputs(4213) <= (inputs(106)) and not (inputs(72));
    layer0_outputs(4214) <= not((inputs(255)) or (inputs(230)));
    layer0_outputs(4215) <= not((inputs(173)) xor (inputs(215)));
    layer0_outputs(4216) <= not((inputs(231)) xor (inputs(4)));
    layer0_outputs(4217) <= (inputs(255)) or (inputs(191));
    layer0_outputs(4218) <= inputs(87);
    layer0_outputs(4219) <= inputs(82);
    layer0_outputs(4220) <= (inputs(120)) and not (inputs(141));
    layer0_outputs(4221) <= '0';
    layer0_outputs(4222) <= (inputs(253)) and not (inputs(178));
    layer0_outputs(4223) <= not(inputs(107)) or (inputs(115));
    layer0_outputs(4224) <= inputs(199);
    layer0_outputs(4225) <= (inputs(95)) xor (inputs(75));
    layer0_outputs(4226) <= '1';
    layer0_outputs(4227) <= not(inputs(123)) or (inputs(80));
    layer0_outputs(4228) <= not((inputs(237)) or (inputs(235)));
    layer0_outputs(4229) <= inputs(231);
    layer0_outputs(4230) <= not((inputs(18)) xor (inputs(234)));
    layer0_outputs(4231) <= not(inputs(61)) or (inputs(156));
    layer0_outputs(4232) <= (inputs(66)) xor (inputs(209));
    layer0_outputs(4233) <= (inputs(181)) and not (inputs(236));
    layer0_outputs(4234) <= not(inputs(30)) or (inputs(162));
    layer0_outputs(4235) <= not((inputs(217)) xor (inputs(241)));
    layer0_outputs(4236) <= not((inputs(221)) xor (inputs(47)));
    layer0_outputs(4237) <= (inputs(133)) xor (inputs(147));
    layer0_outputs(4238) <= (inputs(199)) xor (inputs(162));
    layer0_outputs(4239) <= not(inputs(170)) or (inputs(88));
    layer0_outputs(4240) <= not(inputs(134));
    layer0_outputs(4241) <= (inputs(31)) or (inputs(168));
    layer0_outputs(4242) <= (inputs(29)) and not (inputs(160));
    layer0_outputs(4243) <= not(inputs(252)) or (inputs(95));
    layer0_outputs(4244) <= not((inputs(16)) xor (inputs(151)));
    layer0_outputs(4245) <= not((inputs(118)) or (inputs(94)));
    layer0_outputs(4246) <= not(inputs(5));
    layer0_outputs(4247) <= (inputs(216)) and (inputs(213));
    layer0_outputs(4248) <= (inputs(81)) or (inputs(49));
    layer0_outputs(4249) <= not((inputs(38)) xor (inputs(128)));
    layer0_outputs(4250) <= '0';
    layer0_outputs(4251) <= (inputs(48)) xor (inputs(58));
    layer0_outputs(4252) <= not(inputs(101)) or (inputs(20));
    layer0_outputs(4253) <= inputs(150);
    layer0_outputs(4254) <= not((inputs(113)) or (inputs(203)));
    layer0_outputs(4255) <= not((inputs(25)) or (inputs(149)));
    layer0_outputs(4256) <= not(inputs(124)) or (inputs(160));
    layer0_outputs(4257) <= not(inputs(150));
    layer0_outputs(4258) <= (inputs(64)) xor (inputs(208));
    layer0_outputs(4259) <= not((inputs(70)) xor (inputs(134)));
    layer0_outputs(4260) <= '0';
    layer0_outputs(4261) <= (inputs(44)) or (inputs(82));
    layer0_outputs(4262) <= inputs(32);
    layer0_outputs(4263) <= inputs(110);
    layer0_outputs(4264) <= inputs(147);
    layer0_outputs(4265) <= (inputs(0)) and (inputs(93));
    layer0_outputs(4266) <= '0';
    layer0_outputs(4267) <= (inputs(96)) or (inputs(249));
    layer0_outputs(4268) <= not((inputs(112)) or (inputs(99)));
    layer0_outputs(4269) <= not((inputs(71)) or (inputs(190)));
    layer0_outputs(4270) <= not((inputs(56)) xor (inputs(46)));
    layer0_outputs(4271) <= inputs(208);
    layer0_outputs(4272) <= not((inputs(203)) or (inputs(177)));
    layer0_outputs(4273) <= not(inputs(157)) or (inputs(246));
    layer0_outputs(4274) <= not((inputs(36)) or (inputs(185)));
    layer0_outputs(4275) <= not(inputs(186)) or (inputs(13));
    layer0_outputs(4276) <= not((inputs(245)) or (inputs(233)));
    layer0_outputs(4277) <= (inputs(233)) and not (inputs(69));
    layer0_outputs(4278) <= not((inputs(94)) and (inputs(142)));
    layer0_outputs(4279) <= '1';
    layer0_outputs(4280) <= not(inputs(229)) or (inputs(61));
    layer0_outputs(4281) <= inputs(48);
    layer0_outputs(4282) <= (inputs(183)) or (inputs(233));
    layer0_outputs(4283) <= inputs(135);
    layer0_outputs(4284) <= inputs(99);
    layer0_outputs(4285) <= not((inputs(43)) xor (inputs(191)));
    layer0_outputs(4286) <= (inputs(205)) xor (inputs(164));
    layer0_outputs(4287) <= (inputs(68)) or (inputs(52));
    layer0_outputs(4288) <= not((inputs(78)) or (inputs(118)));
    layer0_outputs(4289) <= (inputs(252)) xor (inputs(42));
    layer0_outputs(4290) <= (inputs(113)) or (inputs(193));
    layer0_outputs(4291) <= not(inputs(193));
    layer0_outputs(4292) <= not((inputs(58)) xor (inputs(29)));
    layer0_outputs(4293) <= inputs(131);
    layer0_outputs(4294) <= inputs(102);
    layer0_outputs(4295) <= '0';
    layer0_outputs(4296) <= (inputs(183)) and not (inputs(193));
    layer0_outputs(4297) <= inputs(27);
    layer0_outputs(4298) <= not(inputs(252)) or (inputs(84));
    layer0_outputs(4299) <= not(inputs(59));
    layer0_outputs(4300) <= inputs(58);
    layer0_outputs(4301) <= (inputs(238)) or (inputs(157));
    layer0_outputs(4302) <= not(inputs(30));
    layer0_outputs(4303) <= not(inputs(219)) or (inputs(175));
    layer0_outputs(4304) <= not(inputs(72)) or (inputs(162));
    layer0_outputs(4305) <= (inputs(190)) or (inputs(69));
    layer0_outputs(4306) <= not(inputs(5));
    layer0_outputs(4307) <= inputs(215);
    layer0_outputs(4308) <= not(inputs(156));
    layer0_outputs(4309) <= not(inputs(29));
    layer0_outputs(4310) <= not(inputs(90));
    layer0_outputs(4311) <= (inputs(164)) and not (inputs(3));
    layer0_outputs(4312) <= not(inputs(217));
    layer0_outputs(4313) <= not((inputs(188)) and (inputs(13)));
    layer0_outputs(4314) <= (inputs(36)) xor (inputs(162));
    layer0_outputs(4315) <= not((inputs(249)) xor (inputs(241)));
    layer0_outputs(4316) <= (inputs(241)) xor (inputs(27));
    layer0_outputs(4317) <= inputs(136);
    layer0_outputs(4318) <= not((inputs(119)) or (inputs(204)));
    layer0_outputs(4319) <= not(inputs(135));
    layer0_outputs(4320) <= not((inputs(233)) or (inputs(193)));
    layer0_outputs(4321) <= not(inputs(152)) or (inputs(231));
    layer0_outputs(4322) <= not(inputs(206)) or (inputs(177));
    layer0_outputs(4323) <= not((inputs(24)) xor (inputs(227)));
    layer0_outputs(4324) <= (inputs(134)) and not (inputs(240));
    layer0_outputs(4325) <= (inputs(42)) and not (inputs(33));
    layer0_outputs(4326) <= (inputs(59)) and not (inputs(154));
    layer0_outputs(4327) <= not(inputs(64)) or (inputs(191));
    layer0_outputs(4328) <= not(inputs(181));
    layer0_outputs(4329) <= not(inputs(91)) or (inputs(210));
    layer0_outputs(4330) <= '1';
    layer0_outputs(4331) <= inputs(94);
    layer0_outputs(4332) <= inputs(121);
    layer0_outputs(4333) <= not(inputs(122)) or (inputs(7));
    layer0_outputs(4334) <= not((inputs(207)) or (inputs(70)));
    layer0_outputs(4335) <= (inputs(19)) or (inputs(68));
    layer0_outputs(4336) <= not(inputs(52));
    layer0_outputs(4337) <= (inputs(104)) and not (inputs(220));
    layer0_outputs(4338) <= not((inputs(67)) xor (inputs(94)));
    layer0_outputs(4339) <= (inputs(123)) or (inputs(93));
    layer0_outputs(4340) <= not(inputs(101)) or (inputs(226));
    layer0_outputs(4341) <= (inputs(85)) xor (inputs(151));
    layer0_outputs(4342) <= (inputs(148)) or (inputs(195));
    layer0_outputs(4343) <= inputs(59);
    layer0_outputs(4344) <= (inputs(159)) xor (inputs(165));
    layer0_outputs(4345) <= inputs(123);
    layer0_outputs(4346) <= not((inputs(200)) xor (inputs(214)));
    layer0_outputs(4347) <= (inputs(134)) xor (inputs(247));
    layer0_outputs(4348) <= '1';
    layer0_outputs(4349) <= inputs(60);
    layer0_outputs(4350) <= inputs(75);
    layer0_outputs(4351) <= inputs(214);
    layer0_outputs(4352) <= not((inputs(50)) xor (inputs(194)));
    layer0_outputs(4353) <= not((inputs(195)) or (inputs(134)));
    layer0_outputs(4354) <= inputs(217);
    layer0_outputs(4355) <= inputs(104);
    layer0_outputs(4356) <= not(inputs(180));
    layer0_outputs(4357) <= (inputs(85)) and not (inputs(174));
    layer0_outputs(4358) <= (inputs(108)) or (inputs(125));
    layer0_outputs(4359) <= not(inputs(89));
    layer0_outputs(4360) <= (inputs(149)) or (inputs(101));
    layer0_outputs(4361) <= not(inputs(79)) or (inputs(78));
    layer0_outputs(4362) <= not((inputs(252)) or (inputs(73)));
    layer0_outputs(4363) <= not(inputs(167));
    layer0_outputs(4364) <= (inputs(219)) and (inputs(222));
    layer0_outputs(4365) <= not(inputs(131));
    layer0_outputs(4366) <= inputs(146);
    layer0_outputs(4367) <= not(inputs(173)) or (inputs(0));
    layer0_outputs(4368) <= not((inputs(29)) or (inputs(36)));
    layer0_outputs(4369) <= (inputs(217)) or (inputs(78));
    layer0_outputs(4370) <= '1';
    layer0_outputs(4371) <= (inputs(90)) xor (inputs(47));
    layer0_outputs(4372) <= (inputs(0)) xor (inputs(184));
    layer0_outputs(4373) <= not(inputs(18));
    layer0_outputs(4374) <= not((inputs(54)) xor (inputs(9)));
    layer0_outputs(4375) <= inputs(156);
    layer0_outputs(4376) <= '1';
    layer0_outputs(4377) <= (inputs(247)) or (inputs(142));
    layer0_outputs(4378) <= not((inputs(190)) xor (inputs(242)));
    layer0_outputs(4379) <= not((inputs(80)) or (inputs(224)));
    layer0_outputs(4380) <= not((inputs(48)) and (inputs(65)));
    layer0_outputs(4381) <= not(inputs(92));
    layer0_outputs(4382) <= (inputs(136)) xor (inputs(70));
    layer0_outputs(4383) <= not(inputs(206));
    layer0_outputs(4384) <= inputs(56);
    layer0_outputs(4385) <= (inputs(43)) and (inputs(65));
    layer0_outputs(4386) <= not(inputs(131));
    layer0_outputs(4387) <= (inputs(131)) xor (inputs(15));
    layer0_outputs(4388) <= (inputs(40)) or (inputs(50));
    layer0_outputs(4389) <= (inputs(227)) and not (inputs(144));
    layer0_outputs(4390) <= (inputs(137)) or (inputs(224));
    layer0_outputs(4391) <= not(inputs(26));
    layer0_outputs(4392) <= (inputs(99)) and not (inputs(80));
    layer0_outputs(4393) <= not((inputs(10)) or (inputs(36)));
    layer0_outputs(4394) <= inputs(194);
    layer0_outputs(4395) <= (inputs(106)) xor (inputs(123));
    layer0_outputs(4396) <= (inputs(190)) or (inputs(234));
    layer0_outputs(4397) <= not(inputs(54)) or (inputs(87));
    layer0_outputs(4398) <= not(inputs(154));
    layer0_outputs(4399) <= not((inputs(213)) or (inputs(76)));
    layer0_outputs(4400) <= (inputs(91)) or (inputs(150));
    layer0_outputs(4401) <= (inputs(222)) or (inputs(41));
    layer0_outputs(4402) <= not((inputs(216)) or (inputs(91)));
    layer0_outputs(4403) <= '0';
    layer0_outputs(4404) <= not((inputs(170)) or (inputs(181)));
    layer0_outputs(4405) <= not(inputs(8));
    layer0_outputs(4406) <= (inputs(31)) xor (inputs(112));
    layer0_outputs(4407) <= not(inputs(6));
    layer0_outputs(4408) <= (inputs(71)) or (inputs(176));
    layer0_outputs(4409) <= not(inputs(230));
    layer0_outputs(4410) <= (inputs(58)) and (inputs(214));
    layer0_outputs(4411) <= (inputs(93)) and not (inputs(83));
    layer0_outputs(4412) <= inputs(62);
    layer0_outputs(4413) <= '1';
    layer0_outputs(4414) <= not(inputs(218)) or (inputs(167));
    layer0_outputs(4415) <= not(inputs(208));
    layer0_outputs(4416) <= not(inputs(214));
    layer0_outputs(4417) <= (inputs(188)) or (inputs(238));
    layer0_outputs(4418) <= '0';
    layer0_outputs(4419) <= (inputs(111)) and not (inputs(5));
    layer0_outputs(4420) <= (inputs(205)) or (inputs(84));
    layer0_outputs(4421) <= (inputs(36)) or (inputs(30));
    layer0_outputs(4422) <= inputs(235);
    layer0_outputs(4423) <= (inputs(117)) and not (inputs(41));
    layer0_outputs(4424) <= (inputs(126)) or (inputs(149));
    layer0_outputs(4425) <= not((inputs(73)) xor (inputs(67)));
    layer0_outputs(4426) <= not(inputs(217)) or (inputs(144));
    layer0_outputs(4427) <= not((inputs(192)) or (inputs(14)));
    layer0_outputs(4428) <= (inputs(154)) xor (inputs(124));
    layer0_outputs(4429) <= not((inputs(172)) xor (inputs(163)));
    layer0_outputs(4430) <= inputs(102);
    layer0_outputs(4431) <= '1';
    layer0_outputs(4432) <= not((inputs(219)) xor (inputs(196)));
    layer0_outputs(4433) <= inputs(71);
    layer0_outputs(4434) <= (inputs(171)) xor (inputs(12));
    layer0_outputs(4435) <= '0';
    layer0_outputs(4436) <= (inputs(238)) and not (inputs(177));
    layer0_outputs(4437) <= not(inputs(116)) or (inputs(221));
    layer0_outputs(4438) <= not((inputs(181)) or (inputs(176)));
    layer0_outputs(4439) <= (inputs(117)) and not (inputs(98));
    layer0_outputs(4440) <= (inputs(221)) and not (inputs(102));
    layer0_outputs(4441) <= not(inputs(70));
    layer0_outputs(4442) <= not((inputs(110)) xor (inputs(24)));
    layer0_outputs(4443) <= not(inputs(167));
    layer0_outputs(4444) <= '1';
    layer0_outputs(4445) <= not(inputs(150)) or (inputs(20));
    layer0_outputs(4446) <= (inputs(215)) and not (inputs(15));
    layer0_outputs(4447) <= not(inputs(48)) or (inputs(251));
    layer0_outputs(4448) <= (inputs(187)) or (inputs(40));
    layer0_outputs(4449) <= not((inputs(63)) xor (inputs(19)));
    layer0_outputs(4450) <= (inputs(41)) xor (inputs(34));
    layer0_outputs(4451) <= (inputs(11)) and not (inputs(1));
    layer0_outputs(4452) <= not(inputs(233));
    layer0_outputs(4453) <= (inputs(116)) and not (inputs(205));
    layer0_outputs(4454) <= not((inputs(239)) or (inputs(215)));
    layer0_outputs(4455) <= (inputs(110)) and not (inputs(192));
    layer0_outputs(4456) <= not((inputs(108)) and (inputs(164)));
    layer0_outputs(4457) <= '1';
    layer0_outputs(4458) <= (inputs(71)) or (inputs(224));
    layer0_outputs(4459) <= not(inputs(105));
    layer0_outputs(4460) <= (inputs(21)) xor (inputs(245));
    layer0_outputs(4461) <= not(inputs(201)) or (inputs(244));
    layer0_outputs(4462) <= (inputs(124)) or (inputs(199));
    layer0_outputs(4463) <= (inputs(68)) xor (inputs(222));
    layer0_outputs(4464) <= not(inputs(73)) or (inputs(32));
    layer0_outputs(4465) <= not(inputs(215)) or (inputs(128));
    layer0_outputs(4466) <= not((inputs(15)) or (inputs(74)));
    layer0_outputs(4467) <= (inputs(182)) and not (inputs(125));
    layer0_outputs(4468) <= not(inputs(75)) or (inputs(178));
    layer0_outputs(4469) <= not(inputs(216));
    layer0_outputs(4470) <= inputs(77);
    layer0_outputs(4471) <= not(inputs(27)) or (inputs(148));
    layer0_outputs(4472) <= not((inputs(180)) or (inputs(41)));
    layer0_outputs(4473) <= inputs(214);
    layer0_outputs(4474) <= (inputs(35)) xor (inputs(45));
    layer0_outputs(4475) <= not(inputs(123));
    layer0_outputs(4476) <= not((inputs(61)) or (inputs(114)));
    layer0_outputs(4477) <= not((inputs(125)) and (inputs(211)));
    layer0_outputs(4478) <= '0';
    layer0_outputs(4479) <= inputs(32);
    layer0_outputs(4480) <= inputs(96);
    layer0_outputs(4481) <= not(inputs(11)) or (inputs(63));
    layer0_outputs(4482) <= not((inputs(214)) xor (inputs(111)));
    layer0_outputs(4483) <= not((inputs(149)) or (inputs(219)));
    layer0_outputs(4484) <= not(inputs(59)) or (inputs(195));
    layer0_outputs(4485) <= (inputs(85)) and not (inputs(245));
    layer0_outputs(4486) <= not(inputs(27));
    layer0_outputs(4487) <= not((inputs(38)) and (inputs(120)));
    layer0_outputs(4488) <= inputs(73);
    layer0_outputs(4489) <= inputs(24);
    layer0_outputs(4490) <= not((inputs(97)) xor (inputs(180)));
    layer0_outputs(4491) <= (inputs(233)) or (inputs(161));
    layer0_outputs(4492) <= (inputs(171)) and not (inputs(6));
    layer0_outputs(4493) <= not((inputs(196)) or (inputs(118)));
    layer0_outputs(4494) <= (inputs(85)) or (inputs(242));
    layer0_outputs(4495) <= inputs(184);
    layer0_outputs(4496) <= not(inputs(182));
    layer0_outputs(4497) <= (inputs(179)) or (inputs(41));
    layer0_outputs(4498) <= (inputs(84)) or (inputs(127));
    layer0_outputs(4499) <= inputs(132);
    layer0_outputs(4500) <= (inputs(189)) and not (inputs(127));
    layer0_outputs(4501) <= inputs(114);
    layer0_outputs(4502) <= (inputs(9)) and not (inputs(161));
    layer0_outputs(4503) <= not(inputs(89));
    layer0_outputs(4504) <= not((inputs(22)) and (inputs(236)));
    layer0_outputs(4505) <= (inputs(204)) or (inputs(39));
    layer0_outputs(4506) <= inputs(51);
    layer0_outputs(4507) <= not((inputs(184)) or (inputs(179)));
    layer0_outputs(4508) <= (inputs(116)) and not (inputs(207));
    layer0_outputs(4509) <= inputs(125);
    layer0_outputs(4510) <= inputs(214);
    layer0_outputs(4511) <= not((inputs(100)) or (inputs(134)));
    layer0_outputs(4512) <= not(inputs(132));
    layer0_outputs(4513) <= (inputs(181)) and not (inputs(217));
    layer0_outputs(4514) <= (inputs(136)) and not (inputs(13));
    layer0_outputs(4515) <= (inputs(169)) xor (inputs(146));
    layer0_outputs(4516) <= (inputs(102)) xor (inputs(188));
    layer0_outputs(4517) <= inputs(59);
    layer0_outputs(4518) <= (inputs(216)) and not (inputs(243));
    layer0_outputs(4519) <= inputs(55);
    layer0_outputs(4520) <= not(inputs(61));
    layer0_outputs(4521) <= (inputs(201)) xor (inputs(161));
    layer0_outputs(4522) <= not(inputs(163));
    layer0_outputs(4523) <= not(inputs(171));
    layer0_outputs(4524) <= not(inputs(73)) or (inputs(124));
    layer0_outputs(4525) <= (inputs(55)) and not (inputs(83));
    layer0_outputs(4526) <= (inputs(172)) or (inputs(156));
    layer0_outputs(4527) <= (inputs(21)) xor (inputs(236));
    layer0_outputs(4528) <= not(inputs(5));
    layer0_outputs(4529) <= (inputs(218)) and not (inputs(225));
    layer0_outputs(4530) <= not((inputs(2)) xor (inputs(215)));
    layer0_outputs(4531) <= '1';
    layer0_outputs(4532) <= not(inputs(116)) or (inputs(9));
    layer0_outputs(4533) <= (inputs(235)) or (inputs(43));
    layer0_outputs(4534) <= not((inputs(192)) xor (inputs(218)));
    layer0_outputs(4535) <= not(inputs(112));
    layer0_outputs(4536) <= (inputs(202)) or (inputs(49));
    layer0_outputs(4537) <= inputs(238);
    layer0_outputs(4538) <= (inputs(104)) or (inputs(45));
    layer0_outputs(4539) <= not((inputs(15)) or (inputs(47)));
    layer0_outputs(4540) <= (inputs(55)) xor (inputs(136));
    layer0_outputs(4541) <= (inputs(143)) and (inputs(94));
    layer0_outputs(4542) <= not((inputs(188)) and (inputs(158)));
    layer0_outputs(4543) <= (inputs(119)) and not (inputs(250));
    layer0_outputs(4544) <= not(inputs(196)) or (inputs(190));
    layer0_outputs(4545) <= not((inputs(195)) or (inputs(37)));
    layer0_outputs(4546) <= not(inputs(185)) or (inputs(60));
    layer0_outputs(4547) <= inputs(152);
    layer0_outputs(4548) <= not(inputs(69));
    layer0_outputs(4549) <= not(inputs(112)) or (inputs(108));
    layer0_outputs(4550) <= (inputs(215)) or (inputs(14));
    layer0_outputs(4551) <= inputs(54);
    layer0_outputs(4552) <= '0';
    layer0_outputs(4553) <= not(inputs(39));
    layer0_outputs(4554) <= (inputs(189)) or (inputs(49));
    layer0_outputs(4555) <= (inputs(232)) and (inputs(29));
    layer0_outputs(4556) <= not((inputs(57)) or (inputs(78)));
    layer0_outputs(4557) <= not(inputs(153));
    layer0_outputs(4558) <= not(inputs(149)) or (inputs(175));
    layer0_outputs(4559) <= inputs(196);
    layer0_outputs(4560) <= '1';
    layer0_outputs(4561) <= not(inputs(219));
    layer0_outputs(4562) <= not((inputs(69)) xor (inputs(45)));
    layer0_outputs(4563) <= not((inputs(140)) or (inputs(65)));
    layer0_outputs(4564) <= not(inputs(61)) or (inputs(192));
    layer0_outputs(4565) <= not((inputs(210)) or (inputs(89)));
    layer0_outputs(4566) <= not((inputs(12)) xor (inputs(9)));
    layer0_outputs(4567) <= '0';
    layer0_outputs(4568) <= inputs(228);
    layer0_outputs(4569) <= (inputs(240)) and (inputs(143));
    layer0_outputs(4570) <= not(inputs(49));
    layer0_outputs(4571) <= not((inputs(132)) or (inputs(216)));
    layer0_outputs(4572) <= (inputs(208)) and not (inputs(15));
    layer0_outputs(4573) <= (inputs(199)) or (inputs(53));
    layer0_outputs(4574) <= (inputs(36)) and not (inputs(43));
    layer0_outputs(4575) <= (inputs(28)) xor (inputs(229));
    layer0_outputs(4576) <= (inputs(30)) xor (inputs(228));
    layer0_outputs(4577) <= not(inputs(118)) or (inputs(82));
    layer0_outputs(4578) <= inputs(182);
    layer0_outputs(4579) <= (inputs(187)) and not (inputs(148));
    layer0_outputs(4580) <= inputs(181);
    layer0_outputs(4581) <= not((inputs(234)) or (inputs(23)));
    layer0_outputs(4582) <= (inputs(78)) and (inputs(32));
    layer0_outputs(4583) <= not(inputs(66)) or (inputs(188));
    layer0_outputs(4584) <= not((inputs(101)) or (inputs(84)));
    layer0_outputs(4585) <= not(inputs(101)) or (inputs(174));
    layer0_outputs(4586) <= inputs(86);
    layer0_outputs(4587) <= (inputs(59)) or (inputs(242));
    layer0_outputs(4588) <= (inputs(77)) and not (inputs(35));
    layer0_outputs(4589) <= (inputs(129)) xor (inputs(222));
    layer0_outputs(4590) <= not((inputs(184)) or (inputs(213)));
    layer0_outputs(4591) <= (inputs(101)) or (inputs(174));
    layer0_outputs(4592) <= not((inputs(55)) or (inputs(195)));
    layer0_outputs(4593) <= not((inputs(54)) or (inputs(73)));
    layer0_outputs(4594) <= (inputs(210)) or (inputs(239));
    layer0_outputs(4595) <= not(inputs(214)) or (inputs(100));
    layer0_outputs(4596) <= not((inputs(68)) or (inputs(162)));
    layer0_outputs(4597) <= '1';
    layer0_outputs(4598) <= not((inputs(19)) xor (inputs(103)));
    layer0_outputs(4599) <= (inputs(59)) xor (inputs(240));
    layer0_outputs(4600) <= inputs(43);
    layer0_outputs(4601) <= not((inputs(18)) xor (inputs(27)));
    layer0_outputs(4602) <= not((inputs(150)) or (inputs(43)));
    layer0_outputs(4603) <= (inputs(39)) or (inputs(142));
    layer0_outputs(4604) <= inputs(3);
    layer0_outputs(4605) <= not(inputs(60));
    layer0_outputs(4606) <= (inputs(38)) and not (inputs(215));
    layer0_outputs(4607) <= inputs(1);
    layer0_outputs(4608) <= not((inputs(19)) xor (inputs(229)));
    layer0_outputs(4609) <= inputs(132);
    layer0_outputs(4610) <= not((inputs(42)) xor (inputs(206)));
    layer0_outputs(4611) <= inputs(141);
    layer0_outputs(4612) <= (inputs(150)) and (inputs(88));
    layer0_outputs(4613) <= (inputs(237)) and not (inputs(39));
    layer0_outputs(4614) <= (inputs(87)) and not (inputs(225));
    layer0_outputs(4615) <= inputs(148);
    layer0_outputs(4616) <= not((inputs(80)) or (inputs(136)));
    layer0_outputs(4617) <= not(inputs(222));
    layer0_outputs(4618) <= (inputs(116)) and not (inputs(222));
    layer0_outputs(4619) <= not((inputs(21)) or (inputs(90)));
    layer0_outputs(4620) <= not(inputs(57)) or (inputs(117));
    layer0_outputs(4621) <= not((inputs(37)) or (inputs(12)));
    layer0_outputs(4622) <= inputs(71);
    layer0_outputs(4623) <= not(inputs(133));
    layer0_outputs(4624) <= not(inputs(133));
    layer0_outputs(4625) <= inputs(216);
    layer0_outputs(4626) <= not(inputs(191));
    layer0_outputs(4627) <= not((inputs(136)) xor (inputs(148)));
    layer0_outputs(4628) <= (inputs(130)) and not (inputs(82));
    layer0_outputs(4629) <= '1';
    layer0_outputs(4630) <= (inputs(64)) and not (inputs(48));
    layer0_outputs(4631) <= (inputs(226)) and not (inputs(131));
    layer0_outputs(4632) <= (inputs(11)) or (inputs(158));
    layer0_outputs(4633) <= (inputs(106)) xor (inputs(97));
    layer0_outputs(4634) <= inputs(250);
    layer0_outputs(4635) <= not(inputs(167));
    layer0_outputs(4636) <= (inputs(187)) and (inputs(167));
    layer0_outputs(4637) <= (inputs(49)) and (inputs(1));
    layer0_outputs(4638) <= not((inputs(34)) xor (inputs(20)));
    layer0_outputs(4639) <= not(inputs(68));
    layer0_outputs(4640) <= not((inputs(98)) xor (inputs(252)));
    layer0_outputs(4641) <= not(inputs(142)) or (inputs(249));
    layer0_outputs(4642) <= not((inputs(28)) xor (inputs(221)));
    layer0_outputs(4643) <= not(inputs(152)) or (inputs(25));
    layer0_outputs(4644) <= (inputs(154)) and not (inputs(143));
    layer0_outputs(4645) <= not((inputs(70)) or (inputs(221)));
    layer0_outputs(4646) <= inputs(199);
    layer0_outputs(4647) <= inputs(78);
    layer0_outputs(4648) <= not(inputs(107)) or (inputs(237));
    layer0_outputs(4649) <= not(inputs(104)) or (inputs(0));
    layer0_outputs(4650) <= (inputs(102)) and not (inputs(235));
    layer0_outputs(4651) <= not(inputs(52));
    layer0_outputs(4652) <= not((inputs(209)) or (inputs(173)));
    layer0_outputs(4653) <= not(inputs(174)) or (inputs(181));
    layer0_outputs(4654) <= not(inputs(65)) or (inputs(235));
    layer0_outputs(4655) <= not(inputs(11));
    layer0_outputs(4656) <= (inputs(203)) xor (inputs(32));
    layer0_outputs(4657) <= not((inputs(144)) or (inputs(71)));
    layer0_outputs(4658) <= (inputs(178)) or (inputs(130));
    layer0_outputs(4659) <= not((inputs(61)) or (inputs(239)));
    layer0_outputs(4660) <= not(inputs(52)) or (inputs(79));
    layer0_outputs(4661) <= not((inputs(246)) or (inputs(94)));
    layer0_outputs(4662) <= not(inputs(140)) or (inputs(90));
    layer0_outputs(4663) <= (inputs(235)) or (inputs(141));
    layer0_outputs(4664) <= not(inputs(94));
    layer0_outputs(4665) <= (inputs(255)) and not (inputs(191));
    layer0_outputs(4666) <= not((inputs(27)) xor (inputs(50)));
    layer0_outputs(4667) <= not(inputs(120));
    layer0_outputs(4668) <= not(inputs(173));
    layer0_outputs(4669) <= (inputs(153)) and not (inputs(12));
    layer0_outputs(4670) <= not(inputs(17)) or (inputs(17));
    layer0_outputs(4671) <= inputs(166);
    layer0_outputs(4672) <= not((inputs(45)) or (inputs(112)));
    layer0_outputs(4673) <= not(inputs(31));
    layer0_outputs(4674) <= (inputs(71)) or (inputs(157));
    layer0_outputs(4675) <= '0';
    layer0_outputs(4676) <= not((inputs(189)) or (inputs(88)));
    layer0_outputs(4677) <= not(inputs(187));
    layer0_outputs(4678) <= (inputs(107)) and not (inputs(37));
    layer0_outputs(4679) <= not(inputs(31));
    layer0_outputs(4680) <= (inputs(70)) or (inputs(153));
    layer0_outputs(4681) <= not((inputs(216)) or (inputs(11)));
    layer0_outputs(4682) <= not((inputs(217)) or (inputs(151)));
    layer0_outputs(4683) <= (inputs(192)) and not (inputs(3));
    layer0_outputs(4684) <= (inputs(196)) and not (inputs(140));
    layer0_outputs(4685) <= (inputs(159)) xor (inputs(120));
    layer0_outputs(4686) <= '1';
    layer0_outputs(4687) <= inputs(182);
    layer0_outputs(4688) <= (inputs(86)) xor (inputs(33));
    layer0_outputs(4689) <= not(inputs(150));
    layer0_outputs(4690) <= (inputs(121)) and not (inputs(222));
    layer0_outputs(4691) <= (inputs(199)) or (inputs(100));
    layer0_outputs(4692) <= '1';
    layer0_outputs(4693) <= not((inputs(141)) and (inputs(42)));
    layer0_outputs(4694) <= not((inputs(35)) or (inputs(77)));
    layer0_outputs(4695) <= not(inputs(110)) or (inputs(239));
    layer0_outputs(4696) <= (inputs(197)) and not (inputs(36));
    layer0_outputs(4697) <= not((inputs(225)) xor (inputs(137)));
    layer0_outputs(4698) <= inputs(85);
    layer0_outputs(4699) <= not((inputs(255)) xor (inputs(187)));
    layer0_outputs(4700) <= (inputs(235)) and not (inputs(13));
    layer0_outputs(4701) <= (inputs(176)) and not (inputs(7));
    layer0_outputs(4702) <= (inputs(66)) and (inputs(221));
    layer0_outputs(4703) <= not((inputs(237)) xor (inputs(91)));
    layer0_outputs(4704) <= inputs(140);
    layer0_outputs(4705) <= not(inputs(157)) or (inputs(174));
    layer0_outputs(4706) <= not(inputs(152));
    layer0_outputs(4707) <= (inputs(94)) xor (inputs(218));
    layer0_outputs(4708) <= not(inputs(63)) or (inputs(112));
    layer0_outputs(4709) <= (inputs(243)) and not (inputs(254));
    layer0_outputs(4710) <= (inputs(81)) or (inputs(123));
    layer0_outputs(4711) <= (inputs(197)) or (inputs(77));
    layer0_outputs(4712) <= (inputs(246)) xor (inputs(27));
    layer0_outputs(4713) <= (inputs(95)) xor (inputs(111));
    layer0_outputs(4714) <= not((inputs(34)) xor (inputs(6)));
    layer0_outputs(4715) <= not((inputs(84)) or (inputs(85)));
    layer0_outputs(4716) <= inputs(136);
    layer0_outputs(4717) <= (inputs(53)) and not (inputs(94));
    layer0_outputs(4718) <= inputs(216);
    layer0_outputs(4719) <= not(inputs(155)) or (inputs(129));
    layer0_outputs(4720) <= not((inputs(127)) or (inputs(99)));
    layer0_outputs(4721) <= (inputs(221)) or (inputs(58));
    layer0_outputs(4722) <= not((inputs(172)) or (inputs(186)));
    layer0_outputs(4723) <= not(inputs(122)) or (inputs(20));
    layer0_outputs(4724) <= (inputs(147)) xor (inputs(10));
    layer0_outputs(4725) <= inputs(187);
    layer0_outputs(4726) <= not(inputs(216));
    layer0_outputs(4727) <= not(inputs(143)) or (inputs(82));
    layer0_outputs(4728) <= (inputs(69)) and not (inputs(96));
    layer0_outputs(4729) <= not(inputs(43));
    layer0_outputs(4730) <= (inputs(59)) and not (inputs(248));
    layer0_outputs(4731) <= not((inputs(5)) xor (inputs(213)));
    layer0_outputs(4732) <= inputs(25);
    layer0_outputs(4733) <= not(inputs(180));
    layer0_outputs(4734) <= inputs(165);
    layer0_outputs(4735) <= not((inputs(163)) or (inputs(57)));
    layer0_outputs(4736) <= (inputs(24)) or (inputs(81));
    layer0_outputs(4737) <= not((inputs(36)) and (inputs(218)));
    layer0_outputs(4738) <= inputs(235);
    layer0_outputs(4739) <= (inputs(156)) or (inputs(53));
    layer0_outputs(4740) <= not(inputs(135)) or (inputs(127));
    layer0_outputs(4741) <= (inputs(186)) and not (inputs(210));
    layer0_outputs(4742) <= not((inputs(49)) or (inputs(119)));
    layer0_outputs(4743) <= (inputs(244)) xor (inputs(76));
    layer0_outputs(4744) <= (inputs(72)) or (inputs(95));
    layer0_outputs(4745) <= (inputs(239)) and not (inputs(14));
    layer0_outputs(4746) <= inputs(55);
    layer0_outputs(4747) <= inputs(72);
    layer0_outputs(4748) <= (inputs(97)) xor (inputs(212));
    layer0_outputs(4749) <= not(inputs(241));
    layer0_outputs(4750) <= not((inputs(31)) or (inputs(217)));
    layer0_outputs(4751) <= not(inputs(0));
    layer0_outputs(4752) <= inputs(120);
    layer0_outputs(4753) <= not((inputs(166)) or (inputs(245)));
    layer0_outputs(4754) <= inputs(200);
    layer0_outputs(4755) <= not((inputs(17)) or (inputs(119)));
    layer0_outputs(4756) <= not((inputs(170)) and (inputs(9)));
    layer0_outputs(4757) <= inputs(5);
    layer0_outputs(4758) <= (inputs(41)) xor (inputs(185));
    layer0_outputs(4759) <= (inputs(241)) or (inputs(243));
    layer0_outputs(4760) <= not(inputs(77));
    layer0_outputs(4761) <= (inputs(168)) or (inputs(37));
    layer0_outputs(4762) <= (inputs(45)) or (inputs(236));
    layer0_outputs(4763) <= (inputs(66)) xor (inputs(11));
    layer0_outputs(4764) <= not((inputs(8)) or (inputs(100)));
    layer0_outputs(4765) <= not(inputs(255)) or (inputs(143));
    layer0_outputs(4766) <= not((inputs(112)) xor (inputs(238)));
    layer0_outputs(4767) <= (inputs(58)) and not (inputs(160));
    layer0_outputs(4768) <= not((inputs(241)) or (inputs(192)));
    layer0_outputs(4769) <= not(inputs(41)) or (inputs(124));
    layer0_outputs(4770) <= not(inputs(137));
    layer0_outputs(4771) <= inputs(125);
    layer0_outputs(4772) <= inputs(176);
    layer0_outputs(4773) <= (inputs(204)) or (inputs(203));
    layer0_outputs(4774) <= (inputs(7)) or (inputs(122));
    layer0_outputs(4775) <= (inputs(189)) or (inputs(167));
    layer0_outputs(4776) <= not(inputs(105));
    layer0_outputs(4777) <= inputs(231);
    layer0_outputs(4778) <= (inputs(242)) xor (inputs(158));
    layer0_outputs(4779) <= inputs(148);
    layer0_outputs(4780) <= inputs(199);
    layer0_outputs(4781) <= not(inputs(109));
    layer0_outputs(4782) <= not(inputs(50));
    layer0_outputs(4783) <= not(inputs(100)) or (inputs(51));
    layer0_outputs(4784) <= (inputs(111)) and (inputs(91));
    layer0_outputs(4785) <= (inputs(89)) or (inputs(234));
    layer0_outputs(4786) <= not((inputs(113)) xor (inputs(28)));
    layer0_outputs(4787) <= inputs(155);
    layer0_outputs(4788) <= inputs(139);
    layer0_outputs(4789) <= not(inputs(43)) or (inputs(65));
    layer0_outputs(4790) <= not((inputs(98)) or (inputs(217)));
    layer0_outputs(4791) <= (inputs(248)) xor (inputs(183));
    layer0_outputs(4792) <= '1';
    layer0_outputs(4793) <= '0';
    layer0_outputs(4794) <= not(inputs(209));
    layer0_outputs(4795) <= '0';
    layer0_outputs(4796) <= not(inputs(246));
    layer0_outputs(4797) <= not((inputs(210)) or (inputs(64)));
    layer0_outputs(4798) <= not((inputs(207)) or (inputs(97)));
    layer0_outputs(4799) <= not((inputs(1)) or (inputs(52)));
    layer0_outputs(4800) <= not(inputs(32)) or (inputs(44));
    layer0_outputs(4801) <= not((inputs(9)) xor (inputs(56)));
    layer0_outputs(4802) <= (inputs(2)) or (inputs(133));
    layer0_outputs(4803) <= not(inputs(168)) or (inputs(94));
    layer0_outputs(4804) <= (inputs(124)) and (inputs(26));
    layer0_outputs(4805) <= not((inputs(194)) or (inputs(203)));
    layer0_outputs(4806) <= (inputs(36)) and not (inputs(206));
    layer0_outputs(4807) <= (inputs(66)) and not (inputs(152));
    layer0_outputs(4808) <= (inputs(240)) or (inputs(118));
    layer0_outputs(4809) <= (inputs(81)) xor (inputs(151));
    layer0_outputs(4810) <= (inputs(182)) and (inputs(237));
    layer0_outputs(4811) <= not((inputs(120)) or (inputs(37)));
    layer0_outputs(4812) <= inputs(204);
    layer0_outputs(4813) <= not(inputs(44)) or (inputs(224));
    layer0_outputs(4814) <= inputs(43);
    layer0_outputs(4815) <= not(inputs(158));
    layer0_outputs(4816) <= (inputs(37)) xor (inputs(88));
    layer0_outputs(4817) <= not(inputs(211));
    layer0_outputs(4818) <= not(inputs(86)) or (inputs(126));
    layer0_outputs(4819) <= '1';
    layer0_outputs(4820) <= not(inputs(98));
    layer0_outputs(4821) <= (inputs(236)) or (inputs(131));
    layer0_outputs(4822) <= not((inputs(57)) or (inputs(12)));
    layer0_outputs(4823) <= (inputs(94)) or (inputs(180));
    layer0_outputs(4824) <= '0';
    layer0_outputs(4825) <= inputs(189);
    layer0_outputs(4826) <= inputs(78);
    layer0_outputs(4827) <= not((inputs(252)) or (inputs(166)));
    layer0_outputs(4828) <= not(inputs(182));
    layer0_outputs(4829) <= not((inputs(53)) or (inputs(199)));
    layer0_outputs(4830) <= not(inputs(116));
    layer0_outputs(4831) <= not((inputs(212)) and (inputs(201)));
    layer0_outputs(4832) <= not((inputs(203)) or (inputs(13)));
    layer0_outputs(4833) <= '0';
    layer0_outputs(4834) <= not((inputs(78)) xor (inputs(0)));
    layer0_outputs(4835) <= not((inputs(56)) or (inputs(13)));
    layer0_outputs(4836) <= (inputs(164)) xor (inputs(177));
    layer0_outputs(4837) <= (inputs(204)) or (inputs(157));
    layer0_outputs(4838) <= not(inputs(187));
    layer0_outputs(4839) <= inputs(39);
    layer0_outputs(4840) <= not((inputs(37)) or (inputs(158)));
    layer0_outputs(4841) <= '0';
    layer0_outputs(4842) <= not(inputs(117)) or (inputs(212));
    layer0_outputs(4843) <= (inputs(3)) and not (inputs(98));
    layer0_outputs(4844) <= not((inputs(153)) xor (inputs(1)));
    layer0_outputs(4845) <= not(inputs(143));
    layer0_outputs(4846) <= inputs(121);
    layer0_outputs(4847) <= (inputs(12)) or (inputs(252));
    layer0_outputs(4848) <= (inputs(171)) xor (inputs(115));
    layer0_outputs(4849) <= not(inputs(185));
    layer0_outputs(4850) <= not(inputs(144)) or (inputs(203));
    layer0_outputs(4851) <= '1';
    layer0_outputs(4852) <= (inputs(174)) and not (inputs(32));
    layer0_outputs(4853) <= not(inputs(73));
    layer0_outputs(4854) <= (inputs(12)) and not (inputs(62));
    layer0_outputs(4855) <= not(inputs(189));
    layer0_outputs(4856) <= (inputs(126)) xor (inputs(22));
    layer0_outputs(4857) <= (inputs(85)) or (inputs(98));
    layer0_outputs(4858) <= not(inputs(149));
    layer0_outputs(4859) <= not((inputs(204)) or (inputs(252)));
    layer0_outputs(4860) <= not(inputs(89));
    layer0_outputs(4861) <= inputs(140);
    layer0_outputs(4862) <= (inputs(131)) xor (inputs(166));
    layer0_outputs(4863) <= (inputs(47)) or (inputs(240));
    layer0_outputs(4864) <= inputs(233);
    layer0_outputs(4865) <= inputs(154);
    layer0_outputs(4866) <= (inputs(242)) xor (inputs(205));
    layer0_outputs(4867) <= not((inputs(213)) xor (inputs(18)));
    layer0_outputs(4868) <= (inputs(229)) xor (inputs(236));
    layer0_outputs(4869) <= inputs(92);
    layer0_outputs(4870) <= not((inputs(149)) xor (inputs(112)));
    layer0_outputs(4871) <= inputs(151);
    layer0_outputs(4872) <= (inputs(107)) xor (inputs(222));
    layer0_outputs(4873) <= '0';
    layer0_outputs(4874) <= (inputs(224)) and not (inputs(220));
    layer0_outputs(4875) <= not((inputs(210)) xor (inputs(82)));
    layer0_outputs(4876) <= not(inputs(31)) or (inputs(64));
    layer0_outputs(4877) <= not(inputs(230)) or (inputs(192));
    layer0_outputs(4878) <= not(inputs(222));
    layer0_outputs(4879) <= not((inputs(229)) or (inputs(228)));
    layer0_outputs(4880) <= (inputs(205)) or (inputs(13));
    layer0_outputs(4881) <= '1';
    layer0_outputs(4882) <= not((inputs(245)) xor (inputs(175)));
    layer0_outputs(4883) <= not((inputs(5)) and (inputs(128)));
    layer0_outputs(4884) <= not(inputs(214));
    layer0_outputs(4885) <= '0';
    layer0_outputs(4886) <= (inputs(245)) and (inputs(8));
    layer0_outputs(4887) <= not((inputs(99)) or (inputs(85)));
    layer0_outputs(4888) <= not(inputs(42));
    layer0_outputs(4889) <= (inputs(28)) or (inputs(166));
    layer0_outputs(4890) <= not(inputs(135)) or (inputs(132));
    layer0_outputs(4891) <= (inputs(226)) or (inputs(203));
    layer0_outputs(4892) <= not((inputs(189)) xor (inputs(181)));
    layer0_outputs(4893) <= not(inputs(102));
    layer0_outputs(4894) <= (inputs(145)) or (inputs(9));
    layer0_outputs(4895) <= (inputs(29)) and not (inputs(112));
    layer0_outputs(4896) <= inputs(109);
    layer0_outputs(4897) <= (inputs(153)) or (inputs(119));
    layer0_outputs(4898) <= inputs(163);
    layer0_outputs(4899) <= inputs(194);
    layer0_outputs(4900) <= not(inputs(86));
    layer0_outputs(4901) <= not(inputs(4));
    layer0_outputs(4902) <= (inputs(57)) and not (inputs(12));
    layer0_outputs(4903) <= (inputs(59)) or (inputs(162));
    layer0_outputs(4904) <= not(inputs(122));
    layer0_outputs(4905) <= (inputs(214)) and not (inputs(139));
    layer0_outputs(4906) <= (inputs(196)) and (inputs(43));
    layer0_outputs(4907) <= (inputs(30)) or (inputs(183));
    layer0_outputs(4908) <= not((inputs(15)) or (inputs(71)));
    layer0_outputs(4909) <= (inputs(78)) and not (inputs(124));
    layer0_outputs(4910) <= '0';
    layer0_outputs(4911) <= (inputs(166)) and not (inputs(114));
    layer0_outputs(4912) <= (inputs(185)) and not (inputs(6));
    layer0_outputs(4913) <= (inputs(204)) and not (inputs(96));
    layer0_outputs(4914) <= (inputs(133)) and not (inputs(212));
    layer0_outputs(4915) <= (inputs(195)) xor (inputs(8));
    layer0_outputs(4916) <= '1';
    layer0_outputs(4917) <= not(inputs(62)) or (inputs(66));
    layer0_outputs(4918) <= (inputs(83)) or (inputs(195));
    layer0_outputs(4919) <= inputs(0);
    layer0_outputs(4920) <= inputs(194);
    layer0_outputs(4921) <= not(inputs(118)) or (inputs(191));
    layer0_outputs(4922) <= not(inputs(137));
    layer0_outputs(4923) <= not(inputs(10));
    layer0_outputs(4924) <= (inputs(128)) xor (inputs(37));
    layer0_outputs(4925) <= (inputs(42)) or (inputs(160));
    layer0_outputs(4926) <= not(inputs(146)) or (inputs(114));
    layer0_outputs(4927) <= (inputs(229)) xor (inputs(18));
    layer0_outputs(4928) <= not((inputs(173)) or (inputs(51)));
    layer0_outputs(4929) <= '1';
    layer0_outputs(4930) <= (inputs(54)) or (inputs(69));
    layer0_outputs(4931) <= not(inputs(170)) or (inputs(226));
    layer0_outputs(4932) <= not((inputs(1)) or (inputs(102)));
    layer0_outputs(4933) <= (inputs(189)) or (inputs(66));
    layer0_outputs(4934) <= (inputs(173)) xor (inputs(76));
    layer0_outputs(4935) <= (inputs(3)) or (inputs(217));
    layer0_outputs(4936) <= not(inputs(161));
    layer0_outputs(4937) <= not((inputs(224)) xor (inputs(241)));
    layer0_outputs(4938) <= (inputs(191)) and not (inputs(68));
    layer0_outputs(4939) <= (inputs(234)) xor (inputs(25));
    layer0_outputs(4940) <= not((inputs(122)) or (inputs(165)));
    layer0_outputs(4941) <= (inputs(230)) xor (inputs(51));
    layer0_outputs(4942) <= inputs(169);
    layer0_outputs(4943) <= inputs(91);
    layer0_outputs(4944) <= inputs(188);
    layer0_outputs(4945) <= not((inputs(236)) or (inputs(141)));
    layer0_outputs(4946) <= (inputs(113)) or (inputs(73));
    layer0_outputs(4947) <= not((inputs(72)) xor (inputs(60)));
    layer0_outputs(4948) <= inputs(196);
    layer0_outputs(4949) <= inputs(142);
    layer0_outputs(4950) <= not(inputs(117)) or (inputs(244));
    layer0_outputs(4951) <= not((inputs(136)) xor (inputs(162)));
    layer0_outputs(4952) <= inputs(183);
    layer0_outputs(4953) <= not((inputs(90)) or (inputs(250)));
    layer0_outputs(4954) <= not((inputs(78)) xor (inputs(233)));
    layer0_outputs(4955) <= (inputs(56)) xor (inputs(80));
    layer0_outputs(4956) <= (inputs(6)) xor (inputs(34));
    layer0_outputs(4957) <= (inputs(199)) and not (inputs(66));
    layer0_outputs(4958) <= (inputs(233)) and not (inputs(249));
    layer0_outputs(4959) <= inputs(179);
    layer0_outputs(4960) <= not(inputs(90));
    layer0_outputs(4961) <= not(inputs(210));
    layer0_outputs(4962) <= (inputs(52)) or (inputs(184));
    layer0_outputs(4963) <= not((inputs(132)) xor (inputs(77)));
    layer0_outputs(4964) <= inputs(53);
    layer0_outputs(4965) <= not((inputs(55)) xor (inputs(153)));
    layer0_outputs(4966) <= not((inputs(59)) xor (inputs(242)));
    layer0_outputs(4967) <= '1';
    layer0_outputs(4968) <= not((inputs(217)) xor (inputs(37)));
    layer0_outputs(4969) <= not((inputs(20)) or (inputs(209)));
    layer0_outputs(4970) <= not((inputs(109)) or (inputs(30)));
    layer0_outputs(4971) <= not((inputs(25)) xor (inputs(170)));
    layer0_outputs(4972) <= not(inputs(219));
    layer0_outputs(4973) <= inputs(88);
    layer0_outputs(4974) <= (inputs(108)) or (inputs(57));
    layer0_outputs(4975) <= (inputs(204)) or (inputs(234));
    layer0_outputs(4976) <= (inputs(73)) or (inputs(239));
    layer0_outputs(4977) <= not(inputs(131));
    layer0_outputs(4978) <= not(inputs(84)) or (inputs(188));
    layer0_outputs(4979) <= '1';
    layer0_outputs(4980) <= inputs(151);
    layer0_outputs(4981) <= not((inputs(247)) or (inputs(30)));
    layer0_outputs(4982) <= (inputs(3)) or (inputs(63));
    layer0_outputs(4983) <= (inputs(240)) or (inputs(234));
    layer0_outputs(4984) <= (inputs(213)) and not (inputs(34));
    layer0_outputs(4985) <= (inputs(196)) and not (inputs(67));
    layer0_outputs(4986) <= (inputs(62)) xor (inputs(128));
    layer0_outputs(4987) <= not((inputs(16)) xor (inputs(234)));
    layer0_outputs(4988) <= not(inputs(173)) or (inputs(127));
    layer0_outputs(4989) <= not((inputs(224)) or (inputs(152)));
    layer0_outputs(4990) <= not(inputs(146));
    layer0_outputs(4991) <= not((inputs(49)) xor (inputs(120)));
    layer0_outputs(4992) <= (inputs(253)) and not (inputs(103));
    layer0_outputs(4993) <= (inputs(218)) and (inputs(142));
    layer0_outputs(4994) <= not((inputs(229)) or (inputs(84)));
    layer0_outputs(4995) <= not((inputs(8)) or (inputs(18)));
    layer0_outputs(4996) <= not(inputs(37)) or (inputs(159));
    layer0_outputs(4997) <= not(inputs(1));
    layer0_outputs(4998) <= (inputs(148)) and not (inputs(46));
    layer0_outputs(4999) <= not(inputs(34)) or (inputs(20));
    layer0_outputs(5000) <= (inputs(179)) xor (inputs(229));
    layer0_outputs(5001) <= (inputs(205)) or (inputs(130));
    layer0_outputs(5002) <= (inputs(102)) xor (inputs(239));
    layer0_outputs(5003) <= inputs(150);
    layer0_outputs(5004) <= not((inputs(167)) xor (inputs(0)));
    layer0_outputs(5005) <= not(inputs(147));
    layer0_outputs(5006) <= (inputs(130)) and not (inputs(82));
    layer0_outputs(5007) <= not(inputs(27));
    layer0_outputs(5008) <= '1';
    layer0_outputs(5009) <= (inputs(116)) or (inputs(128));
    layer0_outputs(5010) <= not(inputs(239)) or (inputs(250));
    layer0_outputs(5011) <= not((inputs(229)) xor (inputs(204)));
    layer0_outputs(5012) <= (inputs(63)) and not (inputs(100));
    layer0_outputs(5013) <= not((inputs(243)) or (inputs(112)));
    layer0_outputs(5014) <= inputs(117);
    layer0_outputs(5015) <= not(inputs(134));
    layer0_outputs(5016) <= not((inputs(199)) xor (inputs(230)));
    layer0_outputs(5017) <= not(inputs(153)) or (inputs(236));
    layer0_outputs(5018) <= inputs(201);
    layer0_outputs(5019) <= not((inputs(60)) xor (inputs(95)));
    layer0_outputs(5020) <= (inputs(130)) or (inputs(19));
    layer0_outputs(5021) <= (inputs(197)) and not (inputs(42));
    layer0_outputs(5022) <= (inputs(92)) xor (inputs(202));
    layer0_outputs(5023) <= (inputs(104)) xor (inputs(110));
    layer0_outputs(5024) <= not((inputs(80)) xor (inputs(126)));
    layer0_outputs(5025) <= (inputs(249)) and not (inputs(172));
    layer0_outputs(5026) <= (inputs(199)) xor (inputs(255));
    layer0_outputs(5027) <= not((inputs(53)) or (inputs(191)));
    layer0_outputs(5028) <= inputs(3);
    layer0_outputs(5029) <= not(inputs(40));
    layer0_outputs(5030) <= (inputs(254)) or (inputs(67));
    layer0_outputs(5031) <= (inputs(58)) or (inputs(195));
    layer0_outputs(5032) <= (inputs(190)) or (inputs(16));
    layer0_outputs(5033) <= '1';
    layer0_outputs(5034) <= not((inputs(14)) or (inputs(163)));
    layer0_outputs(5035) <= not(inputs(140));
    layer0_outputs(5036) <= (inputs(177)) or (inputs(222));
    layer0_outputs(5037) <= (inputs(149)) or (inputs(209));
    layer0_outputs(5038) <= (inputs(68)) or (inputs(44));
    layer0_outputs(5039) <= (inputs(94)) and not (inputs(159));
    layer0_outputs(5040) <= not((inputs(67)) or (inputs(226)));
    layer0_outputs(5041) <= not((inputs(154)) or (inputs(154)));
    layer0_outputs(5042) <= (inputs(152)) or (inputs(238));
    layer0_outputs(5043) <= (inputs(50)) or (inputs(39));
    layer0_outputs(5044) <= not((inputs(129)) and (inputs(127)));
    layer0_outputs(5045) <= (inputs(242)) and (inputs(68));
    layer0_outputs(5046) <= (inputs(97)) or (inputs(224));
    layer0_outputs(5047) <= not(inputs(41));
    layer0_outputs(5048) <= inputs(182);
    layer0_outputs(5049) <= not((inputs(123)) or (inputs(150)));
    layer0_outputs(5050) <= inputs(1);
    layer0_outputs(5051) <= '1';
    layer0_outputs(5052) <= not(inputs(93));
    layer0_outputs(5053) <= not((inputs(130)) and (inputs(227)));
    layer0_outputs(5054) <= inputs(108);
    layer0_outputs(5055) <= (inputs(111)) or (inputs(152));
    layer0_outputs(5056) <= (inputs(95)) or (inputs(153));
    layer0_outputs(5057) <= not((inputs(86)) xor (inputs(46)));
    layer0_outputs(5058) <= (inputs(121)) or (inputs(108));
    layer0_outputs(5059) <= (inputs(55)) xor (inputs(249));
    layer0_outputs(5060) <= not(inputs(181)) or (inputs(82));
    layer0_outputs(5061) <= not((inputs(226)) xor (inputs(28)));
    layer0_outputs(5062) <= (inputs(113)) xor (inputs(78));
    layer0_outputs(5063) <= inputs(88);
    layer0_outputs(5064) <= not(inputs(123)) or (inputs(217));
    layer0_outputs(5065) <= not((inputs(55)) or (inputs(179)));
    layer0_outputs(5066) <= (inputs(111)) and not (inputs(225));
    layer0_outputs(5067) <= not(inputs(118));
    layer0_outputs(5068) <= (inputs(136)) xor (inputs(4));
    layer0_outputs(5069) <= not(inputs(59)) or (inputs(177));
    layer0_outputs(5070) <= not((inputs(104)) or (inputs(186)));
    layer0_outputs(5071) <= not(inputs(17)) or (inputs(178));
    layer0_outputs(5072) <= (inputs(52)) or (inputs(198));
    layer0_outputs(5073) <= (inputs(76)) xor (inputs(217));
    layer0_outputs(5074) <= not((inputs(48)) xor (inputs(68)));
    layer0_outputs(5075) <= '0';
    layer0_outputs(5076) <= not(inputs(179));
    layer0_outputs(5077) <= inputs(3);
    layer0_outputs(5078) <= not((inputs(125)) or (inputs(160)));
    layer0_outputs(5079) <= inputs(212);
    layer0_outputs(5080) <= inputs(106);
    layer0_outputs(5081) <= not(inputs(146)) or (inputs(33));
    layer0_outputs(5082) <= (inputs(211)) or (inputs(66));
    layer0_outputs(5083) <= (inputs(235)) and not (inputs(34));
    layer0_outputs(5084) <= (inputs(204)) xor (inputs(145));
    layer0_outputs(5085) <= '1';
    layer0_outputs(5086) <= '0';
    layer0_outputs(5087) <= (inputs(117)) and not (inputs(107));
    layer0_outputs(5088) <= not(inputs(46)) or (inputs(2));
    layer0_outputs(5089) <= inputs(87);
    layer0_outputs(5090) <= not(inputs(196)) or (inputs(112));
    layer0_outputs(5091) <= (inputs(89)) xor (inputs(31));
    layer0_outputs(5092) <= (inputs(76)) xor (inputs(244));
    layer0_outputs(5093) <= not(inputs(229)) or (inputs(110));
    layer0_outputs(5094) <= not((inputs(123)) or (inputs(196)));
    layer0_outputs(5095) <= not(inputs(211)) or (inputs(176));
    layer0_outputs(5096) <= inputs(145);
    layer0_outputs(5097) <= not((inputs(153)) or (inputs(36)));
    layer0_outputs(5098) <= '1';
    layer0_outputs(5099) <= '0';
    layer0_outputs(5100) <= inputs(185);
    layer0_outputs(5101) <= not((inputs(46)) xor (inputs(50)));
    layer0_outputs(5102) <= not(inputs(158)) or (inputs(14));
    layer0_outputs(5103) <= (inputs(202)) xor (inputs(93));
    layer0_outputs(5104) <= not(inputs(56));
    layer0_outputs(5105) <= '0';
    layer0_outputs(5106) <= not((inputs(228)) or (inputs(94)));
    layer0_outputs(5107) <= (inputs(189)) or (inputs(101));
    layer0_outputs(5108) <= not((inputs(40)) or (inputs(166)));
    layer0_outputs(5109) <= (inputs(144)) xor (inputs(56));
    layer0_outputs(5110) <= not(inputs(185)) or (inputs(85));
    layer0_outputs(5111) <= inputs(70);
    layer0_outputs(5112) <= inputs(43);
    layer0_outputs(5113) <= not(inputs(190)) or (inputs(240));
    layer0_outputs(5114) <= (inputs(209)) and not (inputs(19));
    layer0_outputs(5115) <= inputs(169);
    layer0_outputs(5116) <= not(inputs(139));
    layer0_outputs(5117) <= (inputs(235)) xor (inputs(27));
    layer0_outputs(5118) <= (inputs(77)) or (inputs(229));
    layer0_outputs(5119) <= not((inputs(135)) or (inputs(144)));
    layer0_outputs(5120) <= '1';
    layer0_outputs(5121) <= not(inputs(197)) or (inputs(228));
    layer0_outputs(5122) <= (inputs(138)) and not (inputs(159));
    layer0_outputs(5123) <= (inputs(212)) xor (inputs(248));
    layer0_outputs(5124) <= not(inputs(100)) or (inputs(32));
    layer0_outputs(5125) <= (inputs(252)) or (inputs(1));
    layer0_outputs(5126) <= inputs(83);
    layer0_outputs(5127) <= inputs(89);
    layer0_outputs(5128) <= not(inputs(179));
    layer0_outputs(5129) <= inputs(2);
    layer0_outputs(5130) <= inputs(145);
    layer0_outputs(5131) <= (inputs(50)) and not (inputs(30));
    layer0_outputs(5132) <= (inputs(213)) xor (inputs(9));
    layer0_outputs(5133) <= not((inputs(32)) or (inputs(53)));
    layer0_outputs(5134) <= inputs(52);
    layer0_outputs(5135) <= inputs(61);
    layer0_outputs(5136) <= not(inputs(249));
    layer0_outputs(5137) <= not(inputs(180));
    layer0_outputs(5138) <= not(inputs(193)) or (inputs(123));
    layer0_outputs(5139) <= not((inputs(242)) xor (inputs(34)));
    layer0_outputs(5140) <= '1';
    layer0_outputs(5141) <= (inputs(85)) or (inputs(236));
    layer0_outputs(5142) <= not(inputs(234));
    layer0_outputs(5143) <= (inputs(232)) or (inputs(101));
    layer0_outputs(5144) <= not(inputs(2)) or (inputs(235));
    layer0_outputs(5145) <= not(inputs(48));
    layer0_outputs(5146) <= not((inputs(41)) or (inputs(198)));
    layer0_outputs(5147) <= not(inputs(225));
    layer0_outputs(5148) <= not(inputs(136));
    layer0_outputs(5149) <= (inputs(3)) or (inputs(168));
    layer0_outputs(5150) <= not((inputs(62)) or (inputs(161)));
    layer0_outputs(5151) <= (inputs(194)) or (inputs(203));
    layer0_outputs(5152) <= not(inputs(84));
    layer0_outputs(5153) <= (inputs(13)) and (inputs(12));
    layer0_outputs(5154) <= not((inputs(76)) xor (inputs(17)));
    layer0_outputs(5155) <= (inputs(139)) or (inputs(123));
    layer0_outputs(5156) <= not(inputs(72));
    layer0_outputs(5157) <= not(inputs(40));
    layer0_outputs(5158) <= not((inputs(219)) xor (inputs(126)));
    layer0_outputs(5159) <= (inputs(89)) and not (inputs(12));
    layer0_outputs(5160) <= (inputs(146)) or (inputs(47));
    layer0_outputs(5161) <= (inputs(64)) xor (inputs(229));
    layer0_outputs(5162) <= not(inputs(251)) or (inputs(62));
    layer0_outputs(5163) <= inputs(123);
    layer0_outputs(5164) <= inputs(106);
    layer0_outputs(5165) <= not(inputs(100));
    layer0_outputs(5166) <= not(inputs(154));
    layer0_outputs(5167) <= not((inputs(57)) or (inputs(134)));
    layer0_outputs(5168) <= (inputs(141)) or (inputs(81));
    layer0_outputs(5169) <= (inputs(41)) xor (inputs(254));
    layer0_outputs(5170) <= (inputs(228)) and not (inputs(221));
    layer0_outputs(5171) <= not(inputs(15)) or (inputs(49));
    layer0_outputs(5172) <= (inputs(83)) or (inputs(144));
    layer0_outputs(5173) <= inputs(99);
    layer0_outputs(5174) <= not(inputs(140));
    layer0_outputs(5175) <= not((inputs(62)) xor (inputs(18)));
    layer0_outputs(5176) <= '0';
    layer0_outputs(5177) <= not(inputs(197));
    layer0_outputs(5178) <= not((inputs(33)) xor (inputs(118)));
    layer0_outputs(5179) <= (inputs(65)) and not (inputs(240));
    layer0_outputs(5180) <= not(inputs(123)) or (inputs(225));
    layer0_outputs(5181) <= inputs(214);
    layer0_outputs(5182) <= inputs(215);
    layer0_outputs(5183) <= not(inputs(37)) or (inputs(17));
    layer0_outputs(5184) <= (inputs(173)) or (inputs(246));
    layer0_outputs(5185) <= (inputs(154)) and not (inputs(109));
    layer0_outputs(5186) <= not((inputs(242)) xor (inputs(12)));
    layer0_outputs(5187) <= (inputs(244)) xor (inputs(51));
    layer0_outputs(5188) <= not((inputs(219)) or (inputs(0)));
    layer0_outputs(5189) <= not(inputs(90)) or (inputs(36));
    layer0_outputs(5190) <= not((inputs(109)) or (inputs(164)));
    layer0_outputs(5191) <= (inputs(72)) xor (inputs(60));
    layer0_outputs(5192) <= (inputs(206)) xor (inputs(240));
    layer0_outputs(5193) <= not((inputs(211)) or (inputs(182)));
    layer0_outputs(5194) <= not(inputs(33)) or (inputs(226));
    layer0_outputs(5195) <= inputs(114);
    layer0_outputs(5196) <= '1';
    layer0_outputs(5197) <= (inputs(28)) and not (inputs(206));
    layer0_outputs(5198) <= inputs(101);
    layer0_outputs(5199) <= not((inputs(8)) and (inputs(220)));
    layer0_outputs(5200) <= (inputs(105)) and not (inputs(109));
    layer0_outputs(5201) <= not((inputs(205)) and (inputs(80)));
    layer0_outputs(5202) <= inputs(75);
    layer0_outputs(5203) <= not((inputs(204)) or (inputs(216)));
    layer0_outputs(5204) <= inputs(150);
    layer0_outputs(5205) <= not(inputs(196)) or (inputs(63));
    layer0_outputs(5206) <= not((inputs(214)) or (inputs(68)));
    layer0_outputs(5207) <= (inputs(231)) xor (inputs(22));
    layer0_outputs(5208) <= not(inputs(156)) or (inputs(230));
    layer0_outputs(5209) <= not((inputs(78)) or (inputs(165)));
    layer0_outputs(5210) <= not((inputs(24)) xor (inputs(228)));
    layer0_outputs(5211) <= not((inputs(153)) or (inputs(211)));
    layer0_outputs(5212) <= inputs(34);
    layer0_outputs(5213) <= (inputs(192)) and not (inputs(3));
    layer0_outputs(5214) <= not(inputs(3));
    layer0_outputs(5215) <= (inputs(102)) xor (inputs(72));
    layer0_outputs(5216) <= (inputs(169)) xor (inputs(137));
    layer0_outputs(5217) <= inputs(100);
    layer0_outputs(5218) <= '0';
    layer0_outputs(5219) <= (inputs(89)) or (inputs(0));
    layer0_outputs(5220) <= (inputs(2)) or (inputs(176));
    layer0_outputs(5221) <= inputs(19);
    layer0_outputs(5222) <= not((inputs(232)) xor (inputs(29)));
    layer0_outputs(5223) <= '0';
    layer0_outputs(5224) <= (inputs(175)) and (inputs(128));
    layer0_outputs(5225) <= '0';
    layer0_outputs(5226) <= (inputs(30)) and (inputs(175));
    layer0_outputs(5227) <= not(inputs(33));
    layer0_outputs(5228) <= (inputs(248)) and not (inputs(186));
    layer0_outputs(5229) <= not(inputs(171)) or (inputs(9));
    layer0_outputs(5230) <= (inputs(239)) and not (inputs(15));
    layer0_outputs(5231) <= not((inputs(1)) or (inputs(92)));
    layer0_outputs(5232) <= not((inputs(95)) xor (inputs(183)));
    layer0_outputs(5233) <= inputs(118);
    layer0_outputs(5234) <= not((inputs(213)) or (inputs(122)));
    layer0_outputs(5235) <= (inputs(223)) xor (inputs(186));
    layer0_outputs(5236) <= (inputs(67)) and not (inputs(245));
    layer0_outputs(5237) <= not((inputs(60)) xor (inputs(218)));
    layer0_outputs(5238) <= (inputs(120)) xor (inputs(247));
    layer0_outputs(5239) <= not(inputs(155));
    layer0_outputs(5240) <= inputs(135);
    layer0_outputs(5241) <= (inputs(113)) xor (inputs(181));
    layer0_outputs(5242) <= not(inputs(59)) or (inputs(194));
    layer0_outputs(5243) <= (inputs(236)) and not (inputs(191));
    layer0_outputs(5244) <= not(inputs(39)) or (inputs(208));
    layer0_outputs(5245) <= (inputs(101)) xor (inputs(48));
    layer0_outputs(5246) <= (inputs(123)) xor (inputs(195));
    layer0_outputs(5247) <= not((inputs(112)) and (inputs(218)));
    layer0_outputs(5248) <= not(inputs(92)) or (inputs(51));
    layer0_outputs(5249) <= not(inputs(73)) or (inputs(68));
    layer0_outputs(5250) <= inputs(80);
    layer0_outputs(5251) <= (inputs(204)) or (inputs(64));
    layer0_outputs(5252) <= not((inputs(91)) xor (inputs(65)));
    layer0_outputs(5253) <= '0';
    layer0_outputs(5254) <= not(inputs(255)) or (inputs(96));
    layer0_outputs(5255) <= (inputs(214)) and not (inputs(55));
    layer0_outputs(5256) <= not((inputs(65)) or (inputs(168)));
    layer0_outputs(5257) <= (inputs(7)) or (inputs(102));
    layer0_outputs(5258) <= (inputs(12)) and not (inputs(45));
    layer0_outputs(5259) <= (inputs(173)) and not (inputs(41));
    layer0_outputs(5260) <= (inputs(91)) and not (inputs(29));
    layer0_outputs(5261) <= (inputs(121)) or (inputs(52));
    layer0_outputs(5262) <= '0';
    layer0_outputs(5263) <= inputs(44);
    layer0_outputs(5264) <= (inputs(243)) or (inputs(92));
    layer0_outputs(5265) <= '1';
    layer0_outputs(5266) <= inputs(134);
    layer0_outputs(5267) <= (inputs(179)) and not (inputs(211));
    layer0_outputs(5268) <= (inputs(166)) or (inputs(116));
    layer0_outputs(5269) <= inputs(200);
    layer0_outputs(5270) <= not((inputs(107)) or (inputs(247)));
    layer0_outputs(5271) <= inputs(25);
    layer0_outputs(5272) <= not((inputs(229)) or (inputs(50)));
    layer0_outputs(5273) <= inputs(57);
    layer0_outputs(5274) <= (inputs(66)) xor (inputs(173));
    layer0_outputs(5275) <= not(inputs(37)) or (inputs(239));
    layer0_outputs(5276) <= '0';
    layer0_outputs(5277) <= (inputs(161)) and (inputs(174));
    layer0_outputs(5278) <= (inputs(80)) and not (inputs(66));
    layer0_outputs(5279) <= not((inputs(16)) xor (inputs(80)));
    layer0_outputs(5280) <= not((inputs(36)) or (inputs(69)));
    layer0_outputs(5281) <= not(inputs(16));
    layer0_outputs(5282) <= not(inputs(94)) or (inputs(31));
    layer0_outputs(5283) <= not(inputs(116));
    layer0_outputs(5284) <= inputs(39);
    layer0_outputs(5285) <= (inputs(229)) or (inputs(243));
    layer0_outputs(5286) <= (inputs(108)) or (inputs(90));
    layer0_outputs(5287) <= not(inputs(134));
    layer0_outputs(5288) <= not(inputs(87)) or (inputs(244));
    layer0_outputs(5289) <= not(inputs(230));
    layer0_outputs(5290) <= inputs(122);
    layer0_outputs(5291) <= (inputs(66)) and not (inputs(46));
    layer0_outputs(5292) <= not((inputs(135)) xor (inputs(200)));
    layer0_outputs(5293) <= not((inputs(174)) or (inputs(63)));
    layer0_outputs(5294) <= inputs(89);
    layer0_outputs(5295) <= (inputs(154)) and not (inputs(223));
    layer0_outputs(5296) <= (inputs(239)) or (inputs(77));
    layer0_outputs(5297) <= (inputs(67)) or (inputs(164));
    layer0_outputs(5298) <= (inputs(168)) and not (inputs(41));
    layer0_outputs(5299) <= not(inputs(12)) or (inputs(45));
    layer0_outputs(5300) <= (inputs(239)) xor (inputs(113));
    layer0_outputs(5301) <= (inputs(238)) xor (inputs(105));
    layer0_outputs(5302) <= (inputs(120)) and not (inputs(232));
    layer0_outputs(5303) <= not((inputs(169)) xor (inputs(38)));
    layer0_outputs(5304) <= not((inputs(129)) and (inputs(15)));
    layer0_outputs(5305) <= (inputs(166)) and not (inputs(146));
    layer0_outputs(5306) <= (inputs(203)) or (inputs(148));
    layer0_outputs(5307) <= (inputs(75)) xor (inputs(147));
    layer0_outputs(5308) <= (inputs(199)) xor (inputs(183));
    layer0_outputs(5309) <= inputs(242);
    layer0_outputs(5310) <= not((inputs(208)) xor (inputs(238)));
    layer0_outputs(5311) <= (inputs(102)) and not (inputs(28));
    layer0_outputs(5312) <= (inputs(151)) and not (inputs(237));
    layer0_outputs(5313) <= inputs(157);
    layer0_outputs(5314) <= (inputs(187)) and not (inputs(7));
    layer0_outputs(5315) <= not(inputs(202));
    layer0_outputs(5316) <= not((inputs(109)) or (inputs(215)));
    layer0_outputs(5317) <= not((inputs(154)) xor (inputs(84)));
    layer0_outputs(5318) <= not(inputs(19)) or (inputs(79));
    layer0_outputs(5319) <= not((inputs(9)) or (inputs(151)));
    layer0_outputs(5320) <= (inputs(100)) and not (inputs(160));
    layer0_outputs(5321) <= not(inputs(80)) or (inputs(157));
    layer0_outputs(5322) <= not((inputs(216)) or (inputs(38)));
    layer0_outputs(5323) <= not((inputs(181)) xor (inputs(195)));
    layer0_outputs(5324) <= not(inputs(75));
    layer0_outputs(5325) <= inputs(215);
    layer0_outputs(5326) <= not(inputs(2)) or (inputs(226));
    layer0_outputs(5327) <= not((inputs(154)) xor (inputs(188)));
    layer0_outputs(5328) <= (inputs(237)) and (inputs(100));
    layer0_outputs(5329) <= (inputs(193)) or (inputs(168));
    layer0_outputs(5330) <= (inputs(212)) and (inputs(136));
    layer0_outputs(5331) <= (inputs(20)) and not (inputs(209));
    layer0_outputs(5332) <= not(inputs(179)) or (inputs(255));
    layer0_outputs(5333) <= (inputs(92)) xor (inputs(37));
    layer0_outputs(5334) <= not(inputs(202));
    layer0_outputs(5335) <= inputs(103);
    layer0_outputs(5336) <= (inputs(110)) and not (inputs(22));
    layer0_outputs(5337) <= not(inputs(97)) or (inputs(5));
    layer0_outputs(5338) <= not(inputs(108));
    layer0_outputs(5339) <= inputs(139);
    layer0_outputs(5340) <= (inputs(86)) xor (inputs(224));
    layer0_outputs(5341) <= not(inputs(151)) or (inputs(141));
    layer0_outputs(5342) <= inputs(245);
    layer0_outputs(5343) <= (inputs(86)) xor (inputs(193));
    layer0_outputs(5344) <= inputs(148);
    layer0_outputs(5345) <= (inputs(192)) and (inputs(222));
    layer0_outputs(5346) <= (inputs(108)) and not (inputs(164));
    layer0_outputs(5347) <= not((inputs(71)) or (inputs(13)));
    layer0_outputs(5348) <= not(inputs(155));
    layer0_outputs(5349) <= not(inputs(41)) or (inputs(204));
    layer0_outputs(5350) <= not((inputs(146)) or (inputs(103)));
    layer0_outputs(5351) <= (inputs(99)) or (inputs(214));
    layer0_outputs(5352) <= (inputs(18)) and (inputs(48));
    layer0_outputs(5353) <= not(inputs(215)) or (inputs(45));
    layer0_outputs(5354) <= not(inputs(43));
    layer0_outputs(5355) <= not(inputs(156));
    layer0_outputs(5356) <= (inputs(146)) or (inputs(218));
    layer0_outputs(5357) <= not((inputs(158)) or (inputs(146)));
    layer0_outputs(5358) <= (inputs(238)) or (inputs(199));
    layer0_outputs(5359) <= not((inputs(178)) or (inputs(180)));
    layer0_outputs(5360) <= not(inputs(193));
    layer0_outputs(5361) <= (inputs(130)) xor (inputs(206));
    layer0_outputs(5362) <= not((inputs(26)) or (inputs(153)));
    layer0_outputs(5363) <= not((inputs(49)) and (inputs(22)));
    layer0_outputs(5364) <= (inputs(219)) and not (inputs(192));
    layer0_outputs(5365) <= not(inputs(59)) or (inputs(250));
    layer0_outputs(5366) <= (inputs(184)) xor (inputs(105));
    layer0_outputs(5367) <= (inputs(204)) or (inputs(65));
    layer0_outputs(5368) <= not(inputs(86));
    layer0_outputs(5369) <= not((inputs(129)) xor (inputs(227)));
    layer0_outputs(5370) <= (inputs(148)) and not (inputs(21));
    layer0_outputs(5371) <= not(inputs(233)) or (inputs(37));
    layer0_outputs(5372) <= (inputs(77)) or (inputs(188));
    layer0_outputs(5373) <= not((inputs(75)) or (inputs(89)));
    layer0_outputs(5374) <= (inputs(94)) or (inputs(103));
    layer0_outputs(5375) <= (inputs(46)) xor (inputs(130));
    layer0_outputs(5376) <= not(inputs(157)) or (inputs(239));
    layer0_outputs(5377) <= inputs(212);
    layer0_outputs(5378) <= not(inputs(168)) or (inputs(121));
    layer0_outputs(5379) <= (inputs(242)) or (inputs(35));
    layer0_outputs(5380) <= (inputs(231)) or (inputs(88));
    layer0_outputs(5381) <= not(inputs(40));
    layer0_outputs(5382) <= inputs(132);
    layer0_outputs(5383) <= (inputs(255)) or (inputs(66));
    layer0_outputs(5384) <= not((inputs(35)) or (inputs(62)));
    layer0_outputs(5385) <= not((inputs(225)) or (inputs(17)));
    layer0_outputs(5386) <= (inputs(233)) or (inputs(13));
    layer0_outputs(5387) <= (inputs(146)) or (inputs(155));
    layer0_outputs(5388) <= not(inputs(229)) or (inputs(67));
    layer0_outputs(5389) <= '1';
    layer0_outputs(5390) <= not(inputs(86));
    layer0_outputs(5391) <= not((inputs(57)) and (inputs(197)));
    layer0_outputs(5392) <= inputs(184);
    layer0_outputs(5393) <= not((inputs(108)) or (inputs(184)));
    layer0_outputs(5394) <= not((inputs(196)) or (inputs(206)));
    layer0_outputs(5395) <= (inputs(62)) or (inputs(18));
    layer0_outputs(5396) <= (inputs(245)) xor (inputs(181));
    layer0_outputs(5397) <= (inputs(184)) and not (inputs(48));
    layer0_outputs(5398) <= not(inputs(167)) or (inputs(241));
    layer0_outputs(5399) <= (inputs(158)) and not (inputs(29));
    layer0_outputs(5400) <= not((inputs(226)) xor (inputs(106)));
    layer0_outputs(5401) <= not((inputs(247)) xor (inputs(127)));
    layer0_outputs(5402) <= not(inputs(100)) or (inputs(212));
    layer0_outputs(5403) <= not((inputs(7)) or (inputs(131)));
    layer0_outputs(5404) <= not(inputs(209));
    layer0_outputs(5405) <= inputs(107);
    layer0_outputs(5406) <= not(inputs(59));
    layer0_outputs(5407) <= inputs(218);
    layer0_outputs(5408) <= '0';
    layer0_outputs(5409) <= not((inputs(183)) xor (inputs(53)));
    layer0_outputs(5410) <= not((inputs(201)) or (inputs(195)));
    layer0_outputs(5411) <= not(inputs(46));
    layer0_outputs(5412) <= not((inputs(145)) and (inputs(232)));
    layer0_outputs(5413) <= not((inputs(66)) or (inputs(24)));
    layer0_outputs(5414) <= inputs(118);
    layer0_outputs(5415) <= not(inputs(124));
    layer0_outputs(5416) <= not(inputs(151)) or (inputs(75));
    layer0_outputs(5417) <= (inputs(149)) or (inputs(87));
    layer0_outputs(5418) <= inputs(200);
    layer0_outputs(5419) <= not(inputs(124)) or (inputs(67));
    layer0_outputs(5420) <= (inputs(156)) xor (inputs(221));
    layer0_outputs(5421) <= (inputs(208)) and not (inputs(8));
    layer0_outputs(5422) <= not(inputs(167)) or (inputs(253));
    layer0_outputs(5423) <= (inputs(177)) and not (inputs(212));
    layer0_outputs(5424) <= inputs(123);
    layer0_outputs(5425) <= not(inputs(233));
    layer0_outputs(5426) <= (inputs(35)) and not (inputs(245));
    layer0_outputs(5427) <= not(inputs(190)) or (inputs(5));
    layer0_outputs(5428) <= not((inputs(99)) xor (inputs(87)));
    layer0_outputs(5429) <= not((inputs(12)) or (inputs(93)));
    layer0_outputs(5430) <= not((inputs(236)) or (inputs(206)));
    layer0_outputs(5431) <= not(inputs(59));
    layer0_outputs(5432) <= (inputs(138)) and not (inputs(15));
    layer0_outputs(5433) <= not((inputs(113)) or (inputs(139)));
    layer0_outputs(5434) <= (inputs(26)) and (inputs(3));
    layer0_outputs(5435) <= not(inputs(93));
    layer0_outputs(5436) <= not(inputs(84)) or (inputs(81));
    layer0_outputs(5437) <= not((inputs(213)) or (inputs(88)));
    layer0_outputs(5438) <= (inputs(27)) and not (inputs(130));
    layer0_outputs(5439) <= not(inputs(104));
    layer0_outputs(5440) <= (inputs(173)) or (inputs(70));
    layer0_outputs(5441) <= (inputs(119)) and not (inputs(233));
    layer0_outputs(5442) <= not((inputs(0)) xor (inputs(110)));
    layer0_outputs(5443) <= (inputs(133)) and not (inputs(47));
    layer0_outputs(5444) <= (inputs(49)) and not (inputs(1));
    layer0_outputs(5445) <= (inputs(44)) or (inputs(209));
    layer0_outputs(5446) <= not(inputs(134));
    layer0_outputs(5447) <= not((inputs(169)) or (inputs(65)));
    layer0_outputs(5448) <= (inputs(75)) xor (inputs(95));
    layer0_outputs(5449) <= not(inputs(166));
    layer0_outputs(5450) <= '0';
    layer0_outputs(5451) <= not(inputs(117));
    layer0_outputs(5452) <= inputs(56);
    layer0_outputs(5453) <= not(inputs(180)) or (inputs(143));
    layer0_outputs(5454) <= (inputs(11)) and not (inputs(67));
    layer0_outputs(5455) <= (inputs(122)) xor (inputs(125));
    layer0_outputs(5456) <= (inputs(13)) or (inputs(184));
    layer0_outputs(5457) <= (inputs(115)) and (inputs(143));
    layer0_outputs(5458) <= not(inputs(77));
    layer0_outputs(5459) <= inputs(112);
    layer0_outputs(5460) <= (inputs(190)) and not (inputs(250));
    layer0_outputs(5461) <= not((inputs(41)) xor (inputs(76)));
    layer0_outputs(5462) <= not((inputs(170)) or (inputs(7)));
    layer0_outputs(5463) <= (inputs(237)) xor (inputs(67));
    layer0_outputs(5464) <= (inputs(107)) and not (inputs(72));
    layer0_outputs(5465) <= not((inputs(61)) xor (inputs(50)));
    layer0_outputs(5466) <= '1';
    layer0_outputs(5467) <= (inputs(114)) or (inputs(51));
    layer0_outputs(5468) <= not(inputs(119));
    layer0_outputs(5469) <= (inputs(215)) and not (inputs(8));
    layer0_outputs(5470) <= not(inputs(202));
    layer0_outputs(5471) <= (inputs(52)) and not (inputs(52));
    layer0_outputs(5472) <= (inputs(125)) and not (inputs(152));
    layer0_outputs(5473) <= not((inputs(76)) or (inputs(28)));
    layer0_outputs(5474) <= (inputs(185)) or (inputs(141));
    layer0_outputs(5475) <= not((inputs(71)) xor (inputs(145)));
    layer0_outputs(5476) <= inputs(104);
    layer0_outputs(5477) <= not(inputs(55)) or (inputs(161));
    layer0_outputs(5478) <= (inputs(206)) xor (inputs(230));
    layer0_outputs(5479) <= not((inputs(194)) xor (inputs(233)));
    layer0_outputs(5480) <= (inputs(131)) or (inputs(46));
    layer0_outputs(5481) <= not((inputs(167)) or (inputs(208)));
    layer0_outputs(5482) <= (inputs(108)) or (inputs(169));
    layer0_outputs(5483) <= inputs(185);
    layer0_outputs(5484) <= not((inputs(79)) xor (inputs(152)));
    layer0_outputs(5485) <= not(inputs(107));
    layer0_outputs(5486) <= not(inputs(74)) or (inputs(242));
    layer0_outputs(5487) <= not(inputs(102)) or (inputs(227));
    layer0_outputs(5488) <= (inputs(41)) or (inputs(180));
    layer0_outputs(5489) <= not(inputs(187));
    layer0_outputs(5490) <= not(inputs(218)) or (inputs(128));
    layer0_outputs(5491) <= (inputs(254)) and not (inputs(249));
    layer0_outputs(5492) <= (inputs(164)) or (inputs(147));
    layer0_outputs(5493) <= (inputs(97)) or (inputs(13));
    layer0_outputs(5494) <= (inputs(58)) xor (inputs(47));
    layer0_outputs(5495) <= not(inputs(255));
    layer0_outputs(5496) <= (inputs(89)) and (inputs(223));
    layer0_outputs(5497) <= not(inputs(218)) or (inputs(254));
    layer0_outputs(5498) <= not(inputs(87));
    layer0_outputs(5499) <= not((inputs(185)) or (inputs(52)));
    layer0_outputs(5500) <= not((inputs(24)) or (inputs(20)));
    layer0_outputs(5501) <= (inputs(127)) xor (inputs(47));
    layer0_outputs(5502) <= not((inputs(114)) or (inputs(206)));
    layer0_outputs(5503) <= '1';
    layer0_outputs(5504) <= (inputs(72)) or (inputs(175));
    layer0_outputs(5505) <= (inputs(236)) or (inputs(35));
    layer0_outputs(5506) <= (inputs(135)) and not (inputs(85));
    layer0_outputs(5507) <= (inputs(185)) or (inputs(39));
    layer0_outputs(5508) <= (inputs(129)) xor (inputs(219));
    layer0_outputs(5509) <= '0';
    layer0_outputs(5510) <= (inputs(22)) or (inputs(53));
    layer0_outputs(5511) <= not((inputs(154)) or (inputs(185)));
    layer0_outputs(5512) <= (inputs(17)) xor (inputs(23));
    layer0_outputs(5513) <= (inputs(113)) and not (inputs(77));
    layer0_outputs(5514) <= not((inputs(161)) or (inputs(91)));
    layer0_outputs(5515) <= not((inputs(255)) or (inputs(220)));
    layer0_outputs(5516) <= not((inputs(107)) or (inputs(78)));
    layer0_outputs(5517) <= not(inputs(150)) or (inputs(100));
    layer0_outputs(5518) <= '1';
    layer0_outputs(5519) <= not(inputs(64)) or (inputs(243));
    layer0_outputs(5520) <= not(inputs(159));
    layer0_outputs(5521) <= (inputs(18)) and not (inputs(187));
    layer0_outputs(5522) <= (inputs(35)) or (inputs(151));
    layer0_outputs(5523) <= not(inputs(220));
    layer0_outputs(5524) <= (inputs(52)) or (inputs(147));
    layer0_outputs(5525) <= not(inputs(155)) or (inputs(180));
    layer0_outputs(5526) <= (inputs(61)) and not (inputs(247));
    layer0_outputs(5527) <= inputs(133);
    layer0_outputs(5528) <= inputs(218);
    layer0_outputs(5529) <= inputs(22);
    layer0_outputs(5530) <= (inputs(135)) and not (inputs(210));
    layer0_outputs(5531) <= '0';
    layer0_outputs(5532) <= (inputs(155)) or (inputs(80));
    layer0_outputs(5533) <= not(inputs(124)) or (inputs(122));
    layer0_outputs(5534) <= (inputs(196)) and not (inputs(50));
    layer0_outputs(5535) <= (inputs(176)) xor (inputs(82));
    layer0_outputs(5536) <= not((inputs(110)) or (inputs(212)));
    layer0_outputs(5537) <= (inputs(230)) xor (inputs(43));
    layer0_outputs(5538) <= not((inputs(86)) or (inputs(128)));
    layer0_outputs(5539) <= not((inputs(206)) xor (inputs(73)));
    layer0_outputs(5540) <= not(inputs(61));
    layer0_outputs(5541) <= (inputs(53)) xor (inputs(149));
    layer0_outputs(5542) <= (inputs(125)) and not (inputs(175));
    layer0_outputs(5543) <= not(inputs(199));
    layer0_outputs(5544) <= not((inputs(180)) or (inputs(2)));
    layer0_outputs(5545) <= (inputs(124)) and not (inputs(31));
    layer0_outputs(5546) <= inputs(102);
    layer0_outputs(5547) <= (inputs(9)) xor (inputs(43));
    layer0_outputs(5548) <= not((inputs(28)) xor (inputs(249)));
    layer0_outputs(5549) <= (inputs(146)) or (inputs(62));
    layer0_outputs(5550) <= (inputs(171)) and not (inputs(227));
    layer0_outputs(5551) <= (inputs(237)) and not (inputs(254));
    layer0_outputs(5552) <= not((inputs(54)) or (inputs(53)));
    layer0_outputs(5553) <= not(inputs(208));
    layer0_outputs(5554) <= not((inputs(181)) or (inputs(94)));
    layer0_outputs(5555) <= not(inputs(202)) or (inputs(169));
    layer0_outputs(5556) <= inputs(127);
    layer0_outputs(5557) <= not((inputs(184)) or (inputs(3)));
    layer0_outputs(5558) <= inputs(237);
    layer0_outputs(5559) <= inputs(174);
    layer0_outputs(5560) <= not((inputs(73)) or (inputs(190)));
    layer0_outputs(5561) <= (inputs(114)) or (inputs(46));
    layer0_outputs(5562) <= (inputs(62)) or (inputs(38));
    layer0_outputs(5563) <= (inputs(144)) xor (inputs(20));
    layer0_outputs(5564) <= not(inputs(49));
    layer0_outputs(5565) <= (inputs(220)) xor (inputs(214));
    layer0_outputs(5566) <= (inputs(163)) and not (inputs(81));
    layer0_outputs(5567) <= (inputs(158)) or (inputs(149));
    layer0_outputs(5568) <= (inputs(215)) or (inputs(81));
    layer0_outputs(5569) <= not(inputs(72));
    layer0_outputs(5570) <= not(inputs(133));
    layer0_outputs(5571) <= not(inputs(251)) or (inputs(97));
    layer0_outputs(5572) <= (inputs(116)) xor (inputs(138));
    layer0_outputs(5573) <= inputs(174);
    layer0_outputs(5574) <= not((inputs(47)) xor (inputs(125)));
    layer0_outputs(5575) <= not(inputs(68));
    layer0_outputs(5576) <= not((inputs(77)) and (inputs(77)));
    layer0_outputs(5577) <= inputs(192);
    layer0_outputs(5578) <= not(inputs(243)) or (inputs(5));
    layer0_outputs(5579) <= not((inputs(210)) and (inputs(9)));
    layer0_outputs(5580) <= inputs(101);
    layer0_outputs(5581) <= inputs(229);
    layer0_outputs(5582) <= (inputs(23)) and not (inputs(83));
    layer0_outputs(5583) <= (inputs(133)) or (inputs(28));
    layer0_outputs(5584) <= (inputs(158)) and (inputs(226));
    layer0_outputs(5585) <= (inputs(248)) or (inputs(189));
    layer0_outputs(5586) <= (inputs(159)) xor (inputs(213));
    layer0_outputs(5587) <= not(inputs(133));
    layer0_outputs(5588) <= (inputs(198)) and not (inputs(183));
    layer0_outputs(5589) <= (inputs(125)) and not (inputs(50));
    layer0_outputs(5590) <= not((inputs(100)) or (inputs(210)));
    layer0_outputs(5591) <= (inputs(230)) and not (inputs(111));
    layer0_outputs(5592) <= not((inputs(39)) and (inputs(180)));
    layer0_outputs(5593) <= (inputs(56)) and not (inputs(96));
    layer0_outputs(5594) <= (inputs(218)) and not (inputs(255));
    layer0_outputs(5595) <= inputs(205);
    layer0_outputs(5596) <= not((inputs(69)) or (inputs(208)));
    layer0_outputs(5597) <= (inputs(208)) or (inputs(16));
    layer0_outputs(5598) <= inputs(249);
    layer0_outputs(5599) <= not((inputs(22)) xor (inputs(89)));
    layer0_outputs(5600) <= (inputs(49)) or (inputs(150));
    layer0_outputs(5601) <= inputs(46);
    layer0_outputs(5602) <= inputs(106);
    layer0_outputs(5603) <= inputs(172);
    layer0_outputs(5604) <= inputs(198);
    layer0_outputs(5605) <= inputs(4);
    layer0_outputs(5606) <= not(inputs(136));
    layer0_outputs(5607) <= not((inputs(209)) xor (inputs(198)));
    layer0_outputs(5608) <= inputs(60);
    layer0_outputs(5609) <= not(inputs(134));
    layer0_outputs(5610) <= inputs(66);
    layer0_outputs(5611) <= (inputs(111)) or (inputs(154));
    layer0_outputs(5612) <= (inputs(177)) or (inputs(108));
    layer0_outputs(5613) <= inputs(184);
    layer0_outputs(5614) <= (inputs(171)) and not (inputs(99));
    layer0_outputs(5615) <= not((inputs(217)) or (inputs(160)));
    layer0_outputs(5616) <= (inputs(152)) or (inputs(150));
    layer0_outputs(5617) <= not(inputs(52)) or (inputs(99));
    layer0_outputs(5618) <= (inputs(53)) xor (inputs(10));
    layer0_outputs(5619) <= not(inputs(19));
    layer0_outputs(5620) <= not((inputs(247)) xor (inputs(118)));
    layer0_outputs(5621) <= (inputs(183)) xor (inputs(67));
    layer0_outputs(5622) <= not(inputs(2));
    layer0_outputs(5623) <= not(inputs(102));
    layer0_outputs(5624) <= not((inputs(114)) or (inputs(3)));
    layer0_outputs(5625) <= (inputs(228)) and not (inputs(96));
    layer0_outputs(5626) <= not(inputs(48));
    layer0_outputs(5627) <= not((inputs(150)) or (inputs(109)));
    layer0_outputs(5628) <= (inputs(12)) or (inputs(134));
    layer0_outputs(5629) <= inputs(39);
    layer0_outputs(5630) <= not(inputs(185));
    layer0_outputs(5631) <= not(inputs(38)) or (inputs(64));
    layer0_outputs(5632) <= not((inputs(198)) or (inputs(74)));
    layer0_outputs(5633) <= (inputs(97)) and not (inputs(145));
    layer0_outputs(5634) <= inputs(239);
    layer0_outputs(5635) <= not((inputs(171)) or (inputs(166)));
    layer0_outputs(5636) <= '0';
    layer0_outputs(5637) <= not(inputs(43));
    layer0_outputs(5638) <= (inputs(244)) xor (inputs(84));
    layer0_outputs(5639) <= (inputs(165)) xor (inputs(208));
    layer0_outputs(5640) <= not((inputs(172)) or (inputs(238)));
    layer0_outputs(5641) <= not(inputs(70));
    layer0_outputs(5642) <= not(inputs(150));
    layer0_outputs(5643) <= (inputs(225)) and not (inputs(3));
    layer0_outputs(5644) <= not(inputs(117)) or (inputs(114));
    layer0_outputs(5645) <= (inputs(145)) and (inputs(6));
    layer0_outputs(5646) <= not(inputs(245)) or (inputs(97));
    layer0_outputs(5647) <= not(inputs(107));
    layer0_outputs(5648) <= (inputs(147)) and not (inputs(158));
    layer0_outputs(5649) <= not(inputs(110)) or (inputs(47));
    layer0_outputs(5650) <= not(inputs(189)) or (inputs(127));
    layer0_outputs(5651) <= (inputs(103)) or (inputs(122));
    layer0_outputs(5652) <= not((inputs(8)) or (inputs(173)));
    layer0_outputs(5653) <= '1';
    layer0_outputs(5654) <= not((inputs(163)) or (inputs(169)));
    layer0_outputs(5655) <= inputs(136);
    layer0_outputs(5656) <= (inputs(99)) or (inputs(92));
    layer0_outputs(5657) <= not(inputs(218));
    layer0_outputs(5658) <= (inputs(228)) or (inputs(86));
    layer0_outputs(5659) <= not((inputs(98)) or (inputs(232)));
    layer0_outputs(5660) <= not((inputs(148)) xor (inputs(79)));
    layer0_outputs(5661) <= not((inputs(150)) xor (inputs(246)));
    layer0_outputs(5662) <= not((inputs(150)) or (inputs(201)));
    layer0_outputs(5663) <= not(inputs(102));
    layer0_outputs(5664) <= not((inputs(37)) or (inputs(142)));
    layer0_outputs(5665) <= (inputs(69)) or (inputs(115));
    layer0_outputs(5666) <= not((inputs(97)) or (inputs(36)));
    layer0_outputs(5667) <= not((inputs(62)) or (inputs(119)));
    layer0_outputs(5668) <= inputs(197);
    layer0_outputs(5669) <= not((inputs(161)) and (inputs(50)));
    layer0_outputs(5670) <= (inputs(227)) xor (inputs(50));
    layer0_outputs(5671) <= not((inputs(66)) xor (inputs(220)));
    layer0_outputs(5672) <= not(inputs(154));
    layer0_outputs(5673) <= (inputs(120)) xor (inputs(141));
    layer0_outputs(5674) <= (inputs(192)) or (inputs(210));
    layer0_outputs(5675) <= not((inputs(2)) xor (inputs(116)));
    layer0_outputs(5676) <= (inputs(65)) or (inputs(81));
    layer0_outputs(5677) <= inputs(141);
    layer0_outputs(5678) <= inputs(77);
    layer0_outputs(5679) <= inputs(106);
    layer0_outputs(5680) <= not(inputs(193)) or (inputs(178));
    layer0_outputs(5681) <= not((inputs(33)) xor (inputs(90)));
    layer0_outputs(5682) <= not(inputs(63));
    layer0_outputs(5683) <= (inputs(84)) and not (inputs(243));
    layer0_outputs(5684) <= inputs(145);
    layer0_outputs(5685) <= not((inputs(58)) xor (inputs(240)));
    layer0_outputs(5686) <= not(inputs(213)) or (inputs(80));
    layer0_outputs(5687) <= not(inputs(70));
    layer0_outputs(5688) <= '1';
    layer0_outputs(5689) <= not((inputs(234)) or (inputs(130)));
    layer0_outputs(5690) <= not(inputs(54));
    layer0_outputs(5691) <= inputs(174);
    layer0_outputs(5692) <= inputs(91);
    layer0_outputs(5693) <= (inputs(57)) and not (inputs(123));
    layer0_outputs(5694) <= '0';
    layer0_outputs(5695) <= '1';
    layer0_outputs(5696) <= (inputs(121)) and not (inputs(239));
    layer0_outputs(5697) <= not(inputs(91)) or (inputs(38));
    layer0_outputs(5698) <= not((inputs(170)) or (inputs(32)));
    layer0_outputs(5699) <= (inputs(7)) and (inputs(145));
    layer0_outputs(5700) <= not((inputs(122)) and (inputs(225)));
    layer0_outputs(5701) <= not((inputs(178)) or (inputs(251)));
    layer0_outputs(5702) <= (inputs(0)) and not (inputs(15));
    layer0_outputs(5703) <= (inputs(88)) and not (inputs(107));
    layer0_outputs(5704) <= (inputs(91)) and not (inputs(52));
    layer0_outputs(5705) <= inputs(86);
    layer0_outputs(5706) <= (inputs(190)) xor (inputs(217));
    layer0_outputs(5707) <= not((inputs(178)) or (inputs(66)));
    layer0_outputs(5708) <= not(inputs(132)) or (inputs(160));
    layer0_outputs(5709) <= (inputs(135)) xor (inputs(38));
    layer0_outputs(5710) <= '0';
    layer0_outputs(5711) <= not(inputs(107));
    layer0_outputs(5712) <= inputs(105);
    layer0_outputs(5713) <= (inputs(239)) xor (inputs(250));
    layer0_outputs(5714) <= (inputs(176)) and not (inputs(104));
    layer0_outputs(5715) <= (inputs(28)) xor (inputs(166));
    layer0_outputs(5716) <= not(inputs(56));
    layer0_outputs(5717) <= not((inputs(160)) or (inputs(186)));
    layer0_outputs(5718) <= (inputs(52)) and not (inputs(82));
    layer0_outputs(5719) <= inputs(139);
    layer0_outputs(5720) <= inputs(47);
    layer0_outputs(5721) <= not((inputs(139)) or (inputs(110)));
    layer0_outputs(5722) <= (inputs(135)) or (inputs(75));
    layer0_outputs(5723) <= not(inputs(69));
    layer0_outputs(5724) <= not((inputs(87)) or (inputs(43)));
    layer0_outputs(5725) <= '0';
    layer0_outputs(5726) <= not((inputs(87)) xor (inputs(205)));
    layer0_outputs(5727) <= (inputs(136)) and not (inputs(30));
    layer0_outputs(5728) <= not(inputs(230)) or (inputs(82));
    layer0_outputs(5729) <= not(inputs(123)) or (inputs(240));
    layer0_outputs(5730) <= not(inputs(89)) or (inputs(22));
    layer0_outputs(5731) <= not(inputs(167));
    layer0_outputs(5732) <= not(inputs(94));
    layer0_outputs(5733) <= not(inputs(195));
    layer0_outputs(5734) <= not(inputs(0)) or (inputs(76));
    layer0_outputs(5735) <= not(inputs(133)) or (inputs(79));
    layer0_outputs(5736) <= inputs(196);
    layer0_outputs(5737) <= not(inputs(117));
    layer0_outputs(5738) <= inputs(127);
    layer0_outputs(5739) <= not(inputs(68));
    layer0_outputs(5740) <= (inputs(126)) or (inputs(15));
    layer0_outputs(5741) <= (inputs(133)) and not (inputs(32));
    layer0_outputs(5742) <= inputs(85);
    layer0_outputs(5743) <= not(inputs(222));
    layer0_outputs(5744) <= (inputs(234)) or (inputs(183));
    layer0_outputs(5745) <= not((inputs(81)) and (inputs(18)));
    layer0_outputs(5746) <= not(inputs(211)) or (inputs(128));
    layer0_outputs(5747) <= not(inputs(117)) or (inputs(190));
    layer0_outputs(5748) <= '0';
    layer0_outputs(5749) <= (inputs(51)) or (inputs(72));
    layer0_outputs(5750) <= not((inputs(69)) xor (inputs(146)));
    layer0_outputs(5751) <= not(inputs(181));
    layer0_outputs(5752) <= not(inputs(183)) or (inputs(181));
    layer0_outputs(5753) <= not((inputs(30)) or (inputs(181)));
    layer0_outputs(5754) <= not(inputs(200));
    layer0_outputs(5755) <= (inputs(184)) and not (inputs(71));
    layer0_outputs(5756) <= inputs(31);
    layer0_outputs(5757) <= '1';
    layer0_outputs(5758) <= not(inputs(102));
    layer0_outputs(5759) <= not((inputs(2)) xor (inputs(127)));
    layer0_outputs(5760) <= '1';
    layer0_outputs(5761) <= not((inputs(66)) and (inputs(193)));
    layer0_outputs(5762) <= not(inputs(234));
    layer0_outputs(5763) <= not(inputs(191)) or (inputs(158));
    layer0_outputs(5764) <= not((inputs(186)) or (inputs(171)));
    layer0_outputs(5765) <= not(inputs(180));
    layer0_outputs(5766) <= inputs(135);
    layer0_outputs(5767) <= (inputs(122)) and not (inputs(196));
    layer0_outputs(5768) <= inputs(19);
    layer0_outputs(5769) <= not(inputs(119)) or (inputs(26));
    layer0_outputs(5770) <= not(inputs(112)) or (inputs(82));
    layer0_outputs(5771) <= (inputs(181)) or (inputs(63));
    layer0_outputs(5772) <= not((inputs(142)) and (inputs(98)));
    layer0_outputs(5773) <= not((inputs(137)) or (inputs(132)));
    layer0_outputs(5774) <= inputs(116);
    layer0_outputs(5775) <= not(inputs(117));
    layer0_outputs(5776) <= not(inputs(183));
    layer0_outputs(5777) <= (inputs(20)) and not (inputs(98));
    layer0_outputs(5778) <= '1';
    layer0_outputs(5779) <= not(inputs(102));
    layer0_outputs(5780) <= (inputs(209)) xor (inputs(162));
    layer0_outputs(5781) <= not(inputs(121)) or (inputs(23));
    layer0_outputs(5782) <= not(inputs(98));
    layer0_outputs(5783) <= (inputs(25)) and not (inputs(248));
    layer0_outputs(5784) <= (inputs(72)) and not (inputs(47));
    layer0_outputs(5785) <= not((inputs(211)) and (inputs(175)));
    layer0_outputs(5786) <= not((inputs(80)) and (inputs(127)));
    layer0_outputs(5787) <= not(inputs(56));
    layer0_outputs(5788) <= (inputs(166)) xor (inputs(30));
    layer0_outputs(5789) <= not((inputs(61)) and (inputs(64)));
    layer0_outputs(5790) <= (inputs(221)) xor (inputs(238));
    layer0_outputs(5791) <= not(inputs(167));
    layer0_outputs(5792) <= '1';
    layer0_outputs(5793) <= not(inputs(114)) or (inputs(219));
    layer0_outputs(5794) <= not((inputs(228)) xor (inputs(212)));
    layer0_outputs(5795) <= not((inputs(55)) xor (inputs(204)));
    layer0_outputs(5796) <= not(inputs(83));
    layer0_outputs(5797) <= not((inputs(113)) xor (inputs(178)));
    layer0_outputs(5798) <= not(inputs(115)) or (inputs(220));
    layer0_outputs(5799) <= (inputs(240)) or (inputs(35));
    layer0_outputs(5800) <= not((inputs(117)) or (inputs(236)));
    layer0_outputs(5801) <= not((inputs(15)) xor (inputs(4)));
    layer0_outputs(5802) <= not(inputs(124));
    layer0_outputs(5803) <= not((inputs(4)) xor (inputs(216)));
    layer0_outputs(5804) <= (inputs(138)) and not (inputs(188));
    layer0_outputs(5805) <= (inputs(150)) or (inputs(253));
    layer0_outputs(5806) <= inputs(233);
    layer0_outputs(5807) <= not(inputs(14));
    layer0_outputs(5808) <= not(inputs(75));
    layer0_outputs(5809) <= (inputs(118)) and not (inputs(111));
    layer0_outputs(5810) <= (inputs(86)) or (inputs(5));
    layer0_outputs(5811) <= '1';
    layer0_outputs(5812) <= inputs(200);
    layer0_outputs(5813) <= (inputs(133)) or (inputs(6));
    layer0_outputs(5814) <= not(inputs(255));
    layer0_outputs(5815) <= inputs(105);
    layer0_outputs(5816) <= (inputs(87)) and not (inputs(36));
    layer0_outputs(5817) <= inputs(149);
    layer0_outputs(5818) <= (inputs(34)) or (inputs(158));
    layer0_outputs(5819) <= not(inputs(2)) or (inputs(0));
    layer0_outputs(5820) <= inputs(184);
    layer0_outputs(5821) <= not((inputs(236)) and (inputs(7)));
    layer0_outputs(5822) <= not(inputs(112)) or (inputs(10));
    layer0_outputs(5823) <= inputs(111);
    layer0_outputs(5824) <= inputs(248);
    layer0_outputs(5825) <= (inputs(86)) or (inputs(137));
    layer0_outputs(5826) <= inputs(21);
    layer0_outputs(5827) <= (inputs(49)) or (inputs(172));
    layer0_outputs(5828) <= not(inputs(176)) or (inputs(145));
    layer0_outputs(5829) <= not((inputs(100)) xor (inputs(15)));
    layer0_outputs(5830) <= (inputs(118)) xor (inputs(14));
    layer0_outputs(5831) <= (inputs(27)) and not (inputs(19));
    layer0_outputs(5832) <= not(inputs(100)) or (inputs(189));
    layer0_outputs(5833) <= inputs(44);
    layer0_outputs(5834) <= (inputs(87)) and not (inputs(35));
    layer0_outputs(5835) <= (inputs(201)) or (inputs(177));
    layer0_outputs(5836) <= not((inputs(219)) xor (inputs(158)));
    layer0_outputs(5837) <= not((inputs(197)) xor (inputs(27)));
    layer0_outputs(5838) <= not(inputs(168)) or (inputs(214));
    layer0_outputs(5839) <= (inputs(241)) and (inputs(252));
    layer0_outputs(5840) <= not((inputs(184)) xor (inputs(64)));
    layer0_outputs(5841) <= inputs(23);
    layer0_outputs(5842) <= (inputs(254)) or (inputs(189));
    layer0_outputs(5843) <= inputs(148);
    layer0_outputs(5844) <= (inputs(231)) and not (inputs(145));
    layer0_outputs(5845) <= (inputs(217)) or (inputs(96));
    layer0_outputs(5846) <= inputs(139);
    layer0_outputs(5847) <= not((inputs(66)) xor (inputs(234)));
    layer0_outputs(5848) <= not((inputs(27)) or (inputs(60)));
    layer0_outputs(5849) <= not(inputs(138));
    layer0_outputs(5850) <= not(inputs(115));
    layer0_outputs(5851) <= (inputs(65)) and not (inputs(255));
    layer0_outputs(5852) <= not(inputs(205));
    layer0_outputs(5853) <= not((inputs(185)) or (inputs(27)));
    layer0_outputs(5854) <= not((inputs(45)) or (inputs(42)));
    layer0_outputs(5855) <= (inputs(155)) xor (inputs(56));
    layer0_outputs(5856) <= (inputs(199)) and not (inputs(52));
    layer0_outputs(5857) <= inputs(120);
    layer0_outputs(5858) <= not((inputs(160)) xor (inputs(153)));
    layer0_outputs(5859) <= not((inputs(46)) or (inputs(77)));
    layer0_outputs(5860) <= inputs(245);
    layer0_outputs(5861) <= not(inputs(242));
    layer0_outputs(5862) <= '1';
    layer0_outputs(5863) <= (inputs(85)) or (inputs(114));
    layer0_outputs(5864) <= (inputs(104)) and not (inputs(141));
    layer0_outputs(5865) <= (inputs(207)) xor (inputs(106));
    layer0_outputs(5866) <= (inputs(23)) xor (inputs(193));
    layer0_outputs(5867) <= (inputs(24)) and (inputs(243));
    layer0_outputs(5868) <= not((inputs(48)) xor (inputs(152)));
    layer0_outputs(5869) <= not((inputs(40)) or (inputs(164)));
    layer0_outputs(5870) <= not((inputs(25)) xor (inputs(203)));
    layer0_outputs(5871) <= not((inputs(39)) or (inputs(58)));
    layer0_outputs(5872) <= not((inputs(162)) or (inputs(191)));
    layer0_outputs(5873) <= (inputs(76)) and not (inputs(177));
    layer0_outputs(5874) <= (inputs(131)) xor (inputs(252));
    layer0_outputs(5875) <= not(inputs(27)) or (inputs(14));
    layer0_outputs(5876) <= (inputs(31)) xor (inputs(88));
    layer0_outputs(5877) <= not((inputs(25)) xor (inputs(110)));
    layer0_outputs(5878) <= (inputs(191)) and not (inputs(50));
    layer0_outputs(5879) <= inputs(44);
    layer0_outputs(5880) <= (inputs(162)) and not (inputs(250));
    layer0_outputs(5881) <= not(inputs(202)) or (inputs(8));
    layer0_outputs(5882) <= not(inputs(71)) or (inputs(114));
    layer0_outputs(5883) <= not(inputs(225));
    layer0_outputs(5884) <= (inputs(14)) or (inputs(71));
    layer0_outputs(5885) <= (inputs(0)) xor (inputs(194));
    layer0_outputs(5886) <= (inputs(152)) and not (inputs(212));
    layer0_outputs(5887) <= not((inputs(21)) xor (inputs(107)));
    layer0_outputs(5888) <= not(inputs(72)) or (inputs(163));
    layer0_outputs(5889) <= (inputs(0)) or (inputs(179));
    layer0_outputs(5890) <= not(inputs(215)) or (inputs(60));
    layer0_outputs(5891) <= inputs(105);
    layer0_outputs(5892) <= (inputs(30)) or (inputs(237));
    layer0_outputs(5893) <= (inputs(137)) or (inputs(234));
    layer0_outputs(5894) <= not(inputs(253)) or (inputs(114));
    layer0_outputs(5895) <= not(inputs(116));
    layer0_outputs(5896) <= (inputs(73)) and not (inputs(40));
    layer0_outputs(5897) <= inputs(67);
    layer0_outputs(5898) <= (inputs(33)) and not (inputs(183));
    layer0_outputs(5899) <= not(inputs(105)) or (inputs(103));
    layer0_outputs(5900) <= (inputs(59)) and not (inputs(219));
    layer0_outputs(5901) <= '0';
    layer0_outputs(5902) <= not(inputs(157)) or (inputs(127));
    layer0_outputs(5903) <= (inputs(75)) and not (inputs(240));
    layer0_outputs(5904) <= not(inputs(121));
    layer0_outputs(5905) <= (inputs(68)) or (inputs(51));
    layer0_outputs(5906) <= not(inputs(162)) or (inputs(250));
    layer0_outputs(5907) <= not((inputs(129)) xor (inputs(251)));
    layer0_outputs(5908) <= not((inputs(45)) xor (inputs(255)));
    layer0_outputs(5909) <= not((inputs(157)) xor (inputs(204)));
    layer0_outputs(5910) <= not((inputs(56)) or (inputs(162)));
    layer0_outputs(5911) <= (inputs(75)) or (inputs(163));
    layer0_outputs(5912) <= not((inputs(238)) xor (inputs(28)));
    layer0_outputs(5913) <= (inputs(230)) or (inputs(88));
    layer0_outputs(5914) <= not(inputs(94));
    layer0_outputs(5915) <= '1';
    layer0_outputs(5916) <= (inputs(66)) or (inputs(145));
    layer0_outputs(5917) <= (inputs(85)) xor (inputs(36));
    layer0_outputs(5918) <= (inputs(24)) and not (inputs(88));
    layer0_outputs(5919) <= (inputs(203)) xor (inputs(187));
    layer0_outputs(5920) <= not(inputs(77));
    layer0_outputs(5921) <= not((inputs(193)) or (inputs(95)));
    layer0_outputs(5922) <= not((inputs(91)) or (inputs(230)));
    layer0_outputs(5923) <= inputs(94);
    layer0_outputs(5924) <= (inputs(152)) xor (inputs(92));
    layer0_outputs(5925) <= not(inputs(54)) or (inputs(217));
    layer0_outputs(5926) <= (inputs(245)) xor (inputs(79));
    layer0_outputs(5927) <= not((inputs(88)) xor (inputs(222)));
    layer0_outputs(5928) <= (inputs(244)) and (inputs(101));
    layer0_outputs(5929) <= (inputs(213)) and not (inputs(208));
    layer0_outputs(5930) <= not(inputs(102));
    layer0_outputs(5931) <= (inputs(101)) and not (inputs(213));
    layer0_outputs(5932) <= (inputs(77)) xor (inputs(4));
    layer0_outputs(5933) <= (inputs(148)) xor (inputs(13));
    layer0_outputs(5934) <= (inputs(152)) and not (inputs(8));
    layer0_outputs(5935) <= (inputs(26)) and not (inputs(225));
    layer0_outputs(5936) <= inputs(223);
    layer0_outputs(5937) <= not(inputs(218)) or (inputs(109));
    layer0_outputs(5938) <= not(inputs(24));
    layer0_outputs(5939) <= not((inputs(48)) or (inputs(25)));
    layer0_outputs(5940) <= not((inputs(55)) or (inputs(205)));
    layer0_outputs(5941) <= not(inputs(109)) or (inputs(81));
    layer0_outputs(5942) <= (inputs(161)) and not (inputs(158));
    layer0_outputs(5943) <= not((inputs(28)) xor (inputs(118)));
    layer0_outputs(5944) <= not(inputs(41)) or (inputs(114));
    layer0_outputs(5945) <= (inputs(114)) xor (inputs(15));
    layer0_outputs(5946) <= not(inputs(84));
    layer0_outputs(5947) <= (inputs(95)) or (inputs(106));
    layer0_outputs(5948) <= inputs(197);
    layer0_outputs(5949) <= inputs(151);
    layer0_outputs(5950) <= not(inputs(69));
    layer0_outputs(5951) <= not(inputs(202));
    layer0_outputs(5952) <= (inputs(31)) and not (inputs(206));
    layer0_outputs(5953) <= not((inputs(81)) or (inputs(206)));
    layer0_outputs(5954) <= not((inputs(185)) xor (inputs(208)));
    layer0_outputs(5955) <= (inputs(172)) or (inputs(204));
    layer0_outputs(5956) <= not((inputs(199)) and (inputs(196)));
    layer0_outputs(5957) <= not((inputs(195)) xor (inputs(11)));
    layer0_outputs(5958) <= (inputs(120)) or (inputs(30));
    layer0_outputs(5959) <= (inputs(152)) and not (inputs(137));
    layer0_outputs(5960) <= not((inputs(188)) or (inputs(171)));
    layer0_outputs(5961) <= '0';
    layer0_outputs(5962) <= not((inputs(252)) xor (inputs(39)));
    layer0_outputs(5963) <= not(inputs(8)) or (inputs(129));
    layer0_outputs(5964) <= not(inputs(61)) or (inputs(143));
    layer0_outputs(5965) <= not(inputs(162)) or (inputs(237));
    layer0_outputs(5966) <= inputs(250);
    layer0_outputs(5967) <= inputs(72);
    layer0_outputs(5968) <= not((inputs(230)) or (inputs(218)));
    layer0_outputs(5969) <= (inputs(70)) and not (inputs(159));
    layer0_outputs(5970) <= not((inputs(201)) or (inputs(148)));
    layer0_outputs(5971) <= (inputs(156)) and (inputs(8));
    layer0_outputs(5972) <= inputs(212);
    layer0_outputs(5973) <= '1';
    layer0_outputs(5974) <= (inputs(21)) xor (inputs(203));
    layer0_outputs(5975) <= '0';
    layer0_outputs(5976) <= (inputs(129)) or (inputs(227));
    layer0_outputs(5977) <= not(inputs(134));
    layer0_outputs(5978) <= (inputs(97)) and not (inputs(4));
    layer0_outputs(5979) <= not(inputs(254));
    layer0_outputs(5980) <= not(inputs(73)) or (inputs(163));
    layer0_outputs(5981) <= (inputs(243)) xor (inputs(79));
    layer0_outputs(5982) <= (inputs(9)) xor (inputs(157));
    layer0_outputs(5983) <= not((inputs(40)) or (inputs(16)));
    layer0_outputs(5984) <= (inputs(88)) and not (inputs(78));
    layer0_outputs(5985) <= not(inputs(210)) or (inputs(64));
    layer0_outputs(5986) <= not(inputs(180));
    layer0_outputs(5987) <= not(inputs(201));
    layer0_outputs(5988) <= not(inputs(62)) or (inputs(37));
    layer0_outputs(5989) <= (inputs(101)) or (inputs(27));
    layer0_outputs(5990) <= not(inputs(185)) or (inputs(29));
    layer0_outputs(5991) <= (inputs(154)) and not (inputs(51));
    layer0_outputs(5992) <= not(inputs(88)) or (inputs(68));
    layer0_outputs(5993) <= (inputs(138)) and not (inputs(103));
    layer0_outputs(5994) <= not(inputs(22)) or (inputs(4));
    layer0_outputs(5995) <= inputs(124);
    layer0_outputs(5996) <= not((inputs(106)) xor (inputs(228)));
    layer0_outputs(5997) <= (inputs(95)) and (inputs(198));
    layer0_outputs(5998) <= '1';
    layer0_outputs(5999) <= not(inputs(211));
    layer0_outputs(6000) <= (inputs(192)) and not (inputs(4));
    layer0_outputs(6001) <= inputs(241);
    layer0_outputs(6002) <= not(inputs(136));
    layer0_outputs(6003) <= not(inputs(125)) or (inputs(7));
    layer0_outputs(6004) <= inputs(219);
    layer0_outputs(6005) <= (inputs(69)) or (inputs(161));
    layer0_outputs(6006) <= not((inputs(218)) or (inputs(197)));
    layer0_outputs(6007) <= not((inputs(5)) or (inputs(13)));
    layer0_outputs(6008) <= not((inputs(93)) xor (inputs(222)));
    layer0_outputs(6009) <= not(inputs(187));
    layer0_outputs(6010) <= '0';
    layer0_outputs(6011) <= (inputs(60)) and not (inputs(227));
    layer0_outputs(6012) <= (inputs(72)) xor (inputs(13));
    layer0_outputs(6013) <= (inputs(13)) or (inputs(178));
    layer0_outputs(6014) <= not(inputs(142)) or (inputs(30));
    layer0_outputs(6015) <= '0';
    layer0_outputs(6016) <= not((inputs(0)) xor (inputs(215)));
    layer0_outputs(6017) <= not((inputs(22)) and (inputs(68)));
    layer0_outputs(6018) <= not(inputs(103)) or (inputs(205));
    layer0_outputs(6019) <= (inputs(53)) xor (inputs(100));
    layer0_outputs(6020) <= (inputs(89)) and not (inputs(10));
    layer0_outputs(6021) <= not((inputs(109)) and (inputs(97)));
    layer0_outputs(6022) <= not(inputs(191)) or (inputs(12));
    layer0_outputs(6023) <= inputs(191);
    layer0_outputs(6024) <= (inputs(3)) or (inputs(214));
    layer0_outputs(6025) <= inputs(56);
    layer0_outputs(6026) <= (inputs(69)) xor (inputs(249));
    layer0_outputs(6027) <= not(inputs(192));
    layer0_outputs(6028) <= not(inputs(6));
    layer0_outputs(6029) <= not((inputs(93)) xor (inputs(196)));
    layer0_outputs(6030) <= not((inputs(229)) or (inputs(58)));
    layer0_outputs(6031) <= (inputs(70)) xor (inputs(96));
    layer0_outputs(6032) <= (inputs(69)) xor (inputs(199));
    layer0_outputs(6033) <= (inputs(14)) or (inputs(167));
    layer0_outputs(6034) <= not((inputs(255)) xor (inputs(210)));
    layer0_outputs(6035) <= (inputs(156)) and not (inputs(146));
    layer0_outputs(6036) <= not((inputs(180)) or (inputs(86)));
    layer0_outputs(6037) <= not(inputs(116)) or (inputs(141));
    layer0_outputs(6038) <= not((inputs(7)) or (inputs(188)));
    layer0_outputs(6039) <= (inputs(38)) and not (inputs(15));
    layer0_outputs(6040) <= not(inputs(42)) or (inputs(1));
    layer0_outputs(6041) <= inputs(57);
    layer0_outputs(6042) <= (inputs(168)) and not (inputs(251));
    layer0_outputs(6043) <= (inputs(242)) and (inputs(68));
    layer0_outputs(6044) <= not((inputs(50)) xor (inputs(243)));
    layer0_outputs(6045) <= not(inputs(181)) or (inputs(47));
    layer0_outputs(6046) <= not((inputs(164)) or (inputs(138)));
    layer0_outputs(6047) <= not((inputs(116)) or (inputs(130)));
    layer0_outputs(6048) <= not((inputs(193)) and (inputs(129)));
    layer0_outputs(6049) <= (inputs(191)) and not (inputs(63));
    layer0_outputs(6050) <= not((inputs(48)) xor (inputs(34)));
    layer0_outputs(6051) <= (inputs(173)) and (inputs(19));
    layer0_outputs(6052) <= not(inputs(133));
    layer0_outputs(6053) <= not((inputs(69)) or (inputs(162)));
    layer0_outputs(6054) <= not((inputs(205)) or (inputs(191)));
    layer0_outputs(6055) <= (inputs(80)) or (inputs(151));
    layer0_outputs(6056) <= (inputs(223)) xor (inputs(198));
    layer0_outputs(6057) <= not((inputs(205)) or (inputs(232)));
    layer0_outputs(6058) <= inputs(174);
    layer0_outputs(6059) <= not(inputs(181)) or (inputs(124));
    layer0_outputs(6060) <= not(inputs(221));
    layer0_outputs(6061) <= not((inputs(38)) xor (inputs(22)));
    layer0_outputs(6062) <= not(inputs(138)) or (inputs(109));
    layer0_outputs(6063) <= '1';
    layer0_outputs(6064) <= not((inputs(112)) xor (inputs(157)));
    layer0_outputs(6065) <= not(inputs(175)) or (inputs(3));
    layer0_outputs(6066) <= not((inputs(102)) or (inputs(224)));
    layer0_outputs(6067) <= not(inputs(175));
    layer0_outputs(6068) <= not(inputs(125));
    layer0_outputs(6069) <= not((inputs(230)) or (inputs(29)));
    layer0_outputs(6070) <= (inputs(245)) xor (inputs(50));
    layer0_outputs(6071) <= not(inputs(20)) or (inputs(203));
    layer0_outputs(6072) <= (inputs(217)) and not (inputs(244));
    layer0_outputs(6073) <= not(inputs(197));
    layer0_outputs(6074) <= not((inputs(58)) xor (inputs(2)));
    layer0_outputs(6075) <= not((inputs(176)) xor (inputs(66)));
    layer0_outputs(6076) <= not(inputs(120));
    layer0_outputs(6077) <= (inputs(45)) and (inputs(34));
    layer0_outputs(6078) <= not((inputs(43)) or (inputs(190)));
    layer0_outputs(6079) <= (inputs(211)) and not (inputs(65));
    layer0_outputs(6080) <= (inputs(133)) and not (inputs(59));
    layer0_outputs(6081) <= (inputs(100)) and not (inputs(223));
    layer0_outputs(6082) <= not(inputs(170));
    layer0_outputs(6083) <= not((inputs(172)) or (inputs(198)));
    layer0_outputs(6084) <= not((inputs(25)) or (inputs(156)));
    layer0_outputs(6085) <= inputs(112);
    layer0_outputs(6086) <= not((inputs(254)) or (inputs(241)));
    layer0_outputs(6087) <= not((inputs(199)) or (inputs(156)));
    layer0_outputs(6088) <= not((inputs(141)) xor (inputs(195)));
    layer0_outputs(6089) <= (inputs(177)) and (inputs(51));
    layer0_outputs(6090) <= not((inputs(15)) xor (inputs(101)));
    layer0_outputs(6091) <= (inputs(225)) and not (inputs(96));
    layer0_outputs(6092) <= not(inputs(143)) or (inputs(210));
    layer0_outputs(6093) <= '0';
    layer0_outputs(6094) <= (inputs(122)) and not (inputs(195));
    layer0_outputs(6095) <= '1';
    layer0_outputs(6096) <= not(inputs(215)) or (inputs(112));
    layer0_outputs(6097) <= (inputs(118)) and not (inputs(205));
    layer0_outputs(6098) <= not((inputs(174)) or (inputs(137)));
    layer0_outputs(6099) <= (inputs(199)) and not (inputs(45));
    layer0_outputs(6100) <= not(inputs(155));
    layer0_outputs(6101) <= inputs(82);
    layer0_outputs(6102) <= not((inputs(223)) xor (inputs(213)));
    layer0_outputs(6103) <= inputs(189);
    layer0_outputs(6104) <= not(inputs(195)) or (inputs(63));
    layer0_outputs(6105) <= not((inputs(64)) xor (inputs(50)));
    layer0_outputs(6106) <= (inputs(158)) and not (inputs(110));
    layer0_outputs(6107) <= (inputs(23)) or (inputs(229));
    layer0_outputs(6108) <= not((inputs(48)) or (inputs(119)));
    layer0_outputs(6109) <= not(inputs(69));
    layer0_outputs(6110) <= '0';
    layer0_outputs(6111) <= (inputs(52)) or (inputs(67));
    layer0_outputs(6112) <= (inputs(44)) or (inputs(2));
    layer0_outputs(6113) <= (inputs(54)) and not (inputs(153));
    layer0_outputs(6114) <= (inputs(16)) or (inputs(73));
    layer0_outputs(6115) <= '0';
    layer0_outputs(6116) <= not(inputs(87));
    layer0_outputs(6117) <= not(inputs(197)) or (inputs(45));
    layer0_outputs(6118) <= not(inputs(41)) or (inputs(69));
    layer0_outputs(6119) <= inputs(178);
    layer0_outputs(6120) <= (inputs(104)) and not (inputs(125));
    layer0_outputs(6121) <= inputs(244);
    layer0_outputs(6122) <= (inputs(19)) xor (inputs(142));
    layer0_outputs(6123) <= (inputs(192)) and not (inputs(211));
    layer0_outputs(6124) <= not((inputs(220)) or (inputs(135)));
    layer0_outputs(6125) <= not(inputs(134));
    layer0_outputs(6126) <= not((inputs(210)) and (inputs(47)));
    layer0_outputs(6127) <= not(inputs(26));
    layer0_outputs(6128) <= (inputs(90)) xor (inputs(13));
    layer0_outputs(6129) <= (inputs(28)) xor (inputs(182));
    layer0_outputs(6130) <= inputs(75);
    layer0_outputs(6131) <= not((inputs(69)) xor (inputs(203)));
    layer0_outputs(6132) <= not((inputs(150)) or (inputs(142)));
    layer0_outputs(6133) <= not(inputs(245)) or (inputs(255));
    layer0_outputs(6134) <= inputs(213);
    layer0_outputs(6135) <= not((inputs(126)) and (inputs(209)));
    layer0_outputs(6136) <= not((inputs(33)) xor (inputs(188)));
    layer0_outputs(6137) <= not((inputs(132)) or (inputs(31)));
    layer0_outputs(6138) <= not((inputs(28)) or (inputs(102)));
    layer0_outputs(6139) <= inputs(56);
    layer0_outputs(6140) <= (inputs(68)) and (inputs(45));
    layer0_outputs(6141) <= not((inputs(88)) or (inputs(18)));
    layer0_outputs(6142) <= not(inputs(74)) or (inputs(204));
    layer0_outputs(6143) <= not(inputs(207)) or (inputs(252));
    layer0_outputs(6144) <= (inputs(179)) and not (inputs(174));
    layer0_outputs(6145) <= (inputs(49)) and not (inputs(189));
    layer0_outputs(6146) <= (inputs(24)) or (inputs(35));
    layer0_outputs(6147) <= not(inputs(90));
    layer0_outputs(6148) <= inputs(133);
    layer0_outputs(6149) <= not(inputs(150)) or (inputs(157));
    layer0_outputs(6150) <= (inputs(161)) xor (inputs(231));
    layer0_outputs(6151) <= (inputs(89)) and not (inputs(79));
    layer0_outputs(6152) <= (inputs(166)) or (inputs(20));
    layer0_outputs(6153) <= not(inputs(165)) or (inputs(221));
    layer0_outputs(6154) <= not((inputs(146)) and (inputs(64)));
    layer0_outputs(6155) <= not((inputs(25)) xor (inputs(38)));
    layer0_outputs(6156) <= inputs(155);
    layer0_outputs(6157) <= not(inputs(2)) or (inputs(7));
    layer0_outputs(6158) <= (inputs(254)) and (inputs(43));
    layer0_outputs(6159) <= inputs(75);
    layer0_outputs(6160) <= not((inputs(116)) or (inputs(26)));
    layer0_outputs(6161) <= (inputs(251)) xor (inputs(117));
    layer0_outputs(6162) <= not(inputs(178)) or (inputs(83));
    layer0_outputs(6163) <= (inputs(105)) and not (inputs(251));
    layer0_outputs(6164) <= not((inputs(22)) xor (inputs(185)));
    layer0_outputs(6165) <= inputs(91);
    layer0_outputs(6166) <= not(inputs(98));
    layer0_outputs(6167) <= inputs(125);
    layer0_outputs(6168) <= not(inputs(137)) or (inputs(45));
    layer0_outputs(6169) <= not((inputs(129)) xor (inputs(203)));
    layer0_outputs(6170) <= not(inputs(94)) or (inputs(227));
    layer0_outputs(6171) <= (inputs(179)) and not (inputs(25));
    layer0_outputs(6172) <= inputs(170);
    layer0_outputs(6173) <= inputs(89);
    layer0_outputs(6174) <= (inputs(187)) or (inputs(110));
    layer0_outputs(6175) <= inputs(148);
    layer0_outputs(6176) <= (inputs(117)) xor (inputs(70));
    layer0_outputs(6177) <= (inputs(237)) xor (inputs(239));
    layer0_outputs(6178) <= not((inputs(86)) and (inputs(175)));
    layer0_outputs(6179) <= not(inputs(182));
    layer0_outputs(6180) <= not((inputs(9)) and (inputs(206)));
    layer0_outputs(6181) <= not(inputs(70)) or (inputs(117));
    layer0_outputs(6182) <= not((inputs(195)) or (inputs(76)));
    layer0_outputs(6183) <= inputs(122);
    layer0_outputs(6184) <= '1';
    layer0_outputs(6185) <= (inputs(111)) xor (inputs(83));
    layer0_outputs(6186) <= (inputs(18)) or (inputs(131));
    layer0_outputs(6187) <= (inputs(233)) and not (inputs(29));
    layer0_outputs(6188) <= not(inputs(132)) or (inputs(232));
    layer0_outputs(6189) <= (inputs(95)) xor (inputs(248));
    layer0_outputs(6190) <= (inputs(20)) and (inputs(81));
    layer0_outputs(6191) <= inputs(58);
    layer0_outputs(6192) <= '0';
    layer0_outputs(6193) <= inputs(180);
    layer0_outputs(6194) <= inputs(166);
    layer0_outputs(6195) <= (inputs(240)) xor (inputs(175));
    layer0_outputs(6196) <= not((inputs(157)) xor (inputs(225)));
    layer0_outputs(6197) <= (inputs(155)) or (inputs(49));
    layer0_outputs(6198) <= not((inputs(248)) or (inputs(240)));
    layer0_outputs(6199) <= (inputs(67)) and (inputs(251));
    layer0_outputs(6200) <= not(inputs(44)) or (inputs(246));
    layer0_outputs(6201) <= (inputs(53)) xor (inputs(174));
    layer0_outputs(6202) <= (inputs(41)) or (inputs(21));
    layer0_outputs(6203) <= (inputs(173)) xor (inputs(144));
    layer0_outputs(6204) <= (inputs(241)) and not (inputs(28));
    layer0_outputs(6205) <= (inputs(37)) or (inputs(60));
    layer0_outputs(6206) <= not(inputs(101)) or (inputs(83));
    layer0_outputs(6207) <= inputs(245);
    layer0_outputs(6208) <= (inputs(222)) xor (inputs(139));
    layer0_outputs(6209) <= not((inputs(120)) xor (inputs(48)));
    layer0_outputs(6210) <= (inputs(166)) xor (inputs(19));
    layer0_outputs(6211) <= (inputs(112)) and not (inputs(240));
    layer0_outputs(6212) <= (inputs(28)) and not (inputs(202));
    layer0_outputs(6213) <= inputs(37);
    layer0_outputs(6214) <= not(inputs(163));
    layer0_outputs(6215) <= (inputs(89)) or (inputs(172));
    layer0_outputs(6216) <= (inputs(96)) and not (inputs(113));
    layer0_outputs(6217) <= (inputs(155)) xor (inputs(146));
    layer0_outputs(6218) <= inputs(89);
    layer0_outputs(6219) <= not((inputs(55)) or (inputs(177)));
    layer0_outputs(6220) <= not(inputs(100));
    layer0_outputs(6221) <= '0';
    layer0_outputs(6222) <= '0';
    layer0_outputs(6223) <= not((inputs(230)) or (inputs(236)));
    layer0_outputs(6224) <= not(inputs(132)) or (inputs(27));
    layer0_outputs(6225) <= (inputs(110)) or (inputs(202));
    layer0_outputs(6226) <= (inputs(214)) and not (inputs(47));
    layer0_outputs(6227) <= not(inputs(135));
    layer0_outputs(6228) <= '1';
    layer0_outputs(6229) <= (inputs(109)) xor (inputs(138));
    layer0_outputs(6230) <= not(inputs(53)) or (inputs(9));
    layer0_outputs(6231) <= not((inputs(48)) or (inputs(217)));
    layer0_outputs(6232) <= (inputs(242)) and not (inputs(31));
    layer0_outputs(6233) <= inputs(66);
    layer0_outputs(6234) <= (inputs(57)) or (inputs(129));
    layer0_outputs(6235) <= not(inputs(141));
    layer0_outputs(6236) <= not((inputs(61)) or (inputs(10)));
    layer0_outputs(6237) <= not((inputs(190)) or (inputs(110)));
    layer0_outputs(6238) <= not(inputs(128)) or (inputs(198));
    layer0_outputs(6239) <= not((inputs(90)) xor (inputs(160)));
    layer0_outputs(6240) <= (inputs(108)) or (inputs(178));
    layer0_outputs(6241) <= (inputs(152)) and not (inputs(35));
    layer0_outputs(6242) <= not(inputs(86)) or (inputs(158));
    layer0_outputs(6243) <= not(inputs(102)) or (inputs(67));
    layer0_outputs(6244) <= inputs(65);
    layer0_outputs(6245) <= not(inputs(148)) or (inputs(63));
    layer0_outputs(6246) <= not(inputs(134)) or (inputs(28));
    layer0_outputs(6247) <= (inputs(209)) and not (inputs(253));
    layer0_outputs(6248) <= (inputs(196)) or (inputs(175));
    layer0_outputs(6249) <= (inputs(73)) or (inputs(178));
    layer0_outputs(6250) <= not(inputs(27));
    layer0_outputs(6251) <= not((inputs(211)) or (inputs(156)));
    layer0_outputs(6252) <= inputs(213);
    layer0_outputs(6253) <= (inputs(1)) or (inputs(168));
    layer0_outputs(6254) <= inputs(107);
    layer0_outputs(6255) <= '1';
    layer0_outputs(6256) <= not(inputs(95));
    layer0_outputs(6257) <= (inputs(86)) or (inputs(26));
    layer0_outputs(6258) <= (inputs(175)) xor (inputs(1));
    layer0_outputs(6259) <= (inputs(134)) and not (inputs(127));
    layer0_outputs(6260) <= not(inputs(173));
    layer0_outputs(6261) <= not(inputs(54));
    layer0_outputs(6262) <= not(inputs(247)) or (inputs(190));
    layer0_outputs(6263) <= not(inputs(106)) or (inputs(232));
    layer0_outputs(6264) <= (inputs(12)) and not (inputs(108));
    layer0_outputs(6265) <= inputs(41);
    layer0_outputs(6266) <= (inputs(4)) and not (inputs(229));
    layer0_outputs(6267) <= (inputs(52)) or (inputs(193));
    layer0_outputs(6268) <= '1';
    layer0_outputs(6269) <= not((inputs(201)) and (inputs(197)));
    layer0_outputs(6270) <= inputs(147);
    layer0_outputs(6271) <= not(inputs(1));
    layer0_outputs(6272) <= not(inputs(100));
    layer0_outputs(6273) <= not(inputs(214));
    layer0_outputs(6274) <= inputs(19);
    layer0_outputs(6275) <= not(inputs(79));
    layer0_outputs(6276) <= not(inputs(178)) or (inputs(15));
    layer0_outputs(6277) <= not((inputs(166)) or (inputs(218)));
    layer0_outputs(6278) <= not((inputs(162)) or (inputs(0)));
    layer0_outputs(6279) <= inputs(191);
    layer0_outputs(6280) <= not((inputs(54)) xor (inputs(204)));
    layer0_outputs(6281) <= (inputs(156)) xor (inputs(126));
    layer0_outputs(6282) <= (inputs(172)) and not (inputs(65));
    layer0_outputs(6283) <= (inputs(196)) and not (inputs(33));
    layer0_outputs(6284) <= '0';
    layer0_outputs(6285) <= (inputs(18)) and (inputs(81));
    layer0_outputs(6286) <= not((inputs(110)) or (inputs(153)));
    layer0_outputs(6287) <= (inputs(188)) xor (inputs(140));
    layer0_outputs(6288) <= (inputs(38)) or (inputs(225));
    layer0_outputs(6289) <= (inputs(126)) xor (inputs(189));
    layer0_outputs(6290) <= not((inputs(153)) or (inputs(68)));
    layer0_outputs(6291) <= inputs(232);
    layer0_outputs(6292) <= (inputs(148)) or (inputs(125));
    layer0_outputs(6293) <= not((inputs(119)) xor (inputs(222)));
    layer0_outputs(6294) <= (inputs(218)) and not (inputs(15));
    layer0_outputs(6295) <= not(inputs(243));
    layer0_outputs(6296) <= (inputs(237)) or (inputs(231));
    layer0_outputs(6297) <= (inputs(220)) or (inputs(31));
    layer0_outputs(6298) <= not(inputs(20));
    layer0_outputs(6299) <= not((inputs(148)) or (inputs(166)));
    layer0_outputs(6300) <= not(inputs(96));
    layer0_outputs(6301) <= not(inputs(171));
    layer0_outputs(6302) <= not(inputs(233));
    layer0_outputs(6303) <= '1';
    layer0_outputs(6304) <= (inputs(196)) and not (inputs(194));
    layer0_outputs(6305) <= not(inputs(181));
    layer0_outputs(6306) <= not(inputs(163)) or (inputs(151));
    layer0_outputs(6307) <= not((inputs(166)) or (inputs(35)));
    layer0_outputs(6308) <= not((inputs(81)) xor (inputs(172)));
    layer0_outputs(6309) <= inputs(107);
    layer0_outputs(6310) <= not((inputs(113)) or (inputs(255)));
    layer0_outputs(6311) <= inputs(149);
    layer0_outputs(6312) <= not(inputs(119));
    layer0_outputs(6313) <= not(inputs(181)) or (inputs(148));
    layer0_outputs(6314) <= (inputs(163)) or (inputs(107));
    layer0_outputs(6315) <= not((inputs(48)) xor (inputs(20)));
    layer0_outputs(6316) <= not(inputs(76)) or (inputs(39));
    layer0_outputs(6317) <= (inputs(183)) xor (inputs(104));
    layer0_outputs(6318) <= not((inputs(47)) xor (inputs(130)));
    layer0_outputs(6319) <= not((inputs(134)) xor (inputs(109)));
    layer0_outputs(6320) <= not((inputs(234)) xor (inputs(50)));
    layer0_outputs(6321) <= (inputs(70)) or (inputs(109));
    layer0_outputs(6322) <= (inputs(206)) or (inputs(190));
    layer0_outputs(6323) <= not((inputs(246)) and (inputs(238)));
    layer0_outputs(6324) <= inputs(4);
    layer0_outputs(6325) <= inputs(212);
    layer0_outputs(6326) <= not(inputs(21)) or (inputs(104));
    layer0_outputs(6327) <= not((inputs(245)) xor (inputs(62)));
    layer0_outputs(6328) <= inputs(197);
    layer0_outputs(6329) <= '1';
    layer0_outputs(6330) <= inputs(169);
    layer0_outputs(6331) <= not(inputs(121));
    layer0_outputs(6332) <= inputs(176);
    layer0_outputs(6333) <= (inputs(39)) or (inputs(206));
    layer0_outputs(6334) <= (inputs(83)) xor (inputs(231));
    layer0_outputs(6335) <= (inputs(34)) and not (inputs(1));
    layer0_outputs(6336) <= not(inputs(121)) or (inputs(28));
    layer0_outputs(6337) <= (inputs(61)) and not (inputs(174));
    layer0_outputs(6338) <= not((inputs(202)) xor (inputs(21)));
    layer0_outputs(6339) <= inputs(163);
    layer0_outputs(6340) <= (inputs(125)) or (inputs(90));
    layer0_outputs(6341) <= (inputs(245)) and (inputs(250));
    layer0_outputs(6342) <= not(inputs(11)) or (inputs(250));
    layer0_outputs(6343) <= not((inputs(198)) xor (inputs(53)));
    layer0_outputs(6344) <= not(inputs(48)) or (inputs(142));
    layer0_outputs(6345) <= not(inputs(196));
    layer0_outputs(6346) <= not(inputs(3)) or (inputs(211));
    layer0_outputs(6347) <= (inputs(204)) and not (inputs(246));
    layer0_outputs(6348) <= (inputs(147)) or (inputs(229));
    layer0_outputs(6349) <= not(inputs(134)) or (inputs(83));
    layer0_outputs(6350) <= not((inputs(130)) xor (inputs(51)));
    layer0_outputs(6351) <= inputs(169);
    layer0_outputs(6352) <= not(inputs(133)) or (inputs(195));
    layer0_outputs(6353) <= not((inputs(28)) or (inputs(44)));
    layer0_outputs(6354) <= (inputs(250)) and not (inputs(161));
    layer0_outputs(6355) <= inputs(82);
    layer0_outputs(6356) <= inputs(75);
    layer0_outputs(6357) <= not(inputs(118)) or (inputs(236));
    layer0_outputs(6358) <= not(inputs(227));
    layer0_outputs(6359) <= not((inputs(158)) or (inputs(74)));
    layer0_outputs(6360) <= not(inputs(141));
    layer0_outputs(6361) <= not(inputs(185));
    layer0_outputs(6362) <= not(inputs(120)) or (inputs(131));
    layer0_outputs(6363) <= not(inputs(134));
    layer0_outputs(6364) <= not((inputs(39)) or (inputs(25)));
    layer0_outputs(6365) <= not((inputs(158)) or (inputs(147)));
    layer0_outputs(6366) <= not((inputs(76)) or (inputs(100)));
    layer0_outputs(6367) <= not(inputs(58));
    layer0_outputs(6368) <= inputs(165);
    layer0_outputs(6369) <= not(inputs(200)) or (inputs(159));
    layer0_outputs(6370) <= (inputs(90)) and not (inputs(202));
    layer0_outputs(6371) <= not(inputs(131));
    layer0_outputs(6372) <= not((inputs(238)) and (inputs(2)));
    layer0_outputs(6373) <= (inputs(188)) or (inputs(149));
    layer0_outputs(6374) <= '0';
    layer0_outputs(6375) <= not(inputs(24));
    layer0_outputs(6376) <= inputs(176);
    layer0_outputs(6377) <= not((inputs(25)) and (inputs(129)));
    layer0_outputs(6378) <= inputs(119);
    layer0_outputs(6379) <= not(inputs(102));
    layer0_outputs(6380) <= (inputs(80)) and not (inputs(207));
    layer0_outputs(6381) <= (inputs(227)) and not (inputs(97));
    layer0_outputs(6382) <= '0';
    layer0_outputs(6383) <= (inputs(103)) xor (inputs(222));
    layer0_outputs(6384) <= (inputs(232)) and not (inputs(41));
    layer0_outputs(6385) <= (inputs(228)) xor (inputs(253));
    layer0_outputs(6386) <= not(inputs(72));
    layer0_outputs(6387) <= (inputs(21)) and not (inputs(45));
    layer0_outputs(6388) <= inputs(128);
    layer0_outputs(6389) <= (inputs(87)) and not (inputs(240));
    layer0_outputs(6390) <= inputs(165);
    layer0_outputs(6391) <= (inputs(87)) and not (inputs(174));
    layer0_outputs(6392) <= (inputs(104)) and (inputs(191));
    layer0_outputs(6393) <= not(inputs(147)) or (inputs(208));
    layer0_outputs(6394) <= inputs(226);
    layer0_outputs(6395) <= (inputs(138)) xor (inputs(250));
    layer0_outputs(6396) <= (inputs(123)) and not (inputs(221));
    layer0_outputs(6397) <= (inputs(53)) or (inputs(51));
    layer0_outputs(6398) <= not((inputs(2)) xor (inputs(44)));
    layer0_outputs(6399) <= (inputs(46)) xor (inputs(121));
    layer0_outputs(6400) <= (inputs(105)) or (inputs(33));
    layer0_outputs(6401) <= not(inputs(215));
    layer0_outputs(6402) <= (inputs(53)) and not (inputs(250));
    layer0_outputs(6403) <= (inputs(238)) and not (inputs(237));
    layer0_outputs(6404) <= not((inputs(36)) or (inputs(149)));
    layer0_outputs(6405) <= (inputs(95)) and not (inputs(169));
    layer0_outputs(6406) <= (inputs(219)) and not (inputs(145));
    layer0_outputs(6407) <= (inputs(37)) or (inputs(216));
    layer0_outputs(6408) <= not(inputs(152));
    layer0_outputs(6409) <= '0';
    layer0_outputs(6410) <= not((inputs(179)) or (inputs(54)));
    layer0_outputs(6411) <= not((inputs(255)) or (inputs(131)));
    layer0_outputs(6412) <= (inputs(216)) or (inputs(138));
    layer0_outputs(6413) <= '1';
    layer0_outputs(6414) <= inputs(205);
    layer0_outputs(6415) <= (inputs(71)) and not (inputs(31));
    layer0_outputs(6416) <= inputs(253);
    layer0_outputs(6417) <= not((inputs(85)) xor (inputs(153)));
    layer0_outputs(6418) <= '1';
    layer0_outputs(6419) <= (inputs(105)) and (inputs(195));
    layer0_outputs(6420) <= not((inputs(2)) xor (inputs(168)));
    layer0_outputs(6421) <= not((inputs(92)) or (inputs(87)));
    layer0_outputs(6422) <= not(inputs(124)) or (inputs(194));
    layer0_outputs(6423) <= inputs(25);
    layer0_outputs(6424) <= not((inputs(3)) or (inputs(200)));
    layer0_outputs(6425) <= (inputs(34)) or (inputs(227));
    layer0_outputs(6426) <= not(inputs(109));
    layer0_outputs(6427) <= not((inputs(53)) xor (inputs(223)));
    layer0_outputs(6428) <= not(inputs(88)) or (inputs(144));
    layer0_outputs(6429) <= (inputs(153)) and not (inputs(213));
    layer0_outputs(6430) <= not(inputs(255)) or (inputs(40));
    layer0_outputs(6431) <= not((inputs(82)) xor (inputs(14)));
    layer0_outputs(6432) <= (inputs(197)) xor (inputs(11));
    layer0_outputs(6433) <= inputs(201);
    layer0_outputs(6434) <= not((inputs(42)) xor (inputs(129)));
    layer0_outputs(6435) <= not((inputs(32)) xor (inputs(107)));
    layer0_outputs(6436) <= inputs(195);
    layer0_outputs(6437) <= (inputs(161)) or (inputs(195));
    layer0_outputs(6438) <= inputs(165);
    layer0_outputs(6439) <= (inputs(65)) xor (inputs(25));
    layer0_outputs(6440) <= (inputs(20)) and (inputs(176));
    layer0_outputs(6441) <= (inputs(224)) or (inputs(112));
    layer0_outputs(6442) <= not((inputs(117)) xor (inputs(37)));
    layer0_outputs(6443) <= (inputs(77)) or (inputs(205));
    layer0_outputs(6444) <= not(inputs(27)) or (inputs(218));
    layer0_outputs(6445) <= not(inputs(133)) or (inputs(50));
    layer0_outputs(6446) <= (inputs(88)) or (inputs(251));
    layer0_outputs(6447) <= (inputs(8)) xor (inputs(55));
    layer0_outputs(6448) <= (inputs(36)) and not (inputs(33));
    layer0_outputs(6449) <= inputs(179);
    layer0_outputs(6450) <= not(inputs(29));
    layer0_outputs(6451) <= not(inputs(231)) or (inputs(227));
    layer0_outputs(6452) <= not(inputs(194)) or (inputs(223));
    layer0_outputs(6453) <= not(inputs(216)) or (inputs(210));
    layer0_outputs(6454) <= (inputs(88)) and not (inputs(141));
    layer0_outputs(6455) <= not((inputs(80)) or (inputs(54)));
    layer0_outputs(6456) <= (inputs(203)) and (inputs(81));
    layer0_outputs(6457) <= inputs(41);
    layer0_outputs(6458) <= not(inputs(206));
    layer0_outputs(6459) <= inputs(39);
    layer0_outputs(6460) <= (inputs(191)) and (inputs(149));
    layer0_outputs(6461) <= (inputs(194)) or (inputs(184));
    layer0_outputs(6462) <= (inputs(40)) xor (inputs(176));
    layer0_outputs(6463) <= not(inputs(130));
    layer0_outputs(6464) <= not((inputs(67)) or (inputs(121)));
    layer0_outputs(6465) <= not(inputs(50)) or (inputs(89));
    layer0_outputs(6466) <= (inputs(168)) and not (inputs(173));
    layer0_outputs(6467) <= (inputs(245)) xor (inputs(144));
    layer0_outputs(6468) <= not((inputs(162)) or (inputs(165)));
    layer0_outputs(6469) <= not((inputs(104)) or (inputs(182)));
    layer0_outputs(6470) <= not(inputs(196));
    layer0_outputs(6471) <= (inputs(183)) and not (inputs(237));
    layer0_outputs(6472) <= (inputs(120)) and not (inputs(131));
    layer0_outputs(6473) <= not(inputs(96)) or (inputs(42));
    layer0_outputs(6474) <= (inputs(211)) or (inputs(248));
    layer0_outputs(6475) <= not(inputs(141)) or (inputs(211));
    layer0_outputs(6476) <= (inputs(142)) and (inputs(46));
    layer0_outputs(6477) <= not(inputs(203));
    layer0_outputs(6478) <= inputs(171);
    layer0_outputs(6479) <= (inputs(54)) and not (inputs(20));
    layer0_outputs(6480) <= not((inputs(20)) or (inputs(138)));
    layer0_outputs(6481) <= (inputs(29)) or (inputs(169));
    layer0_outputs(6482) <= (inputs(180)) or (inputs(103));
    layer0_outputs(6483) <= inputs(116);
    layer0_outputs(6484) <= not(inputs(105));
    layer0_outputs(6485) <= not((inputs(123)) or (inputs(148)));
    layer0_outputs(6486) <= not(inputs(79));
    layer0_outputs(6487) <= (inputs(216)) xor (inputs(142));
    layer0_outputs(6488) <= (inputs(239)) and not (inputs(1));
    layer0_outputs(6489) <= (inputs(194)) and (inputs(48));
    layer0_outputs(6490) <= inputs(40);
    layer0_outputs(6491) <= not((inputs(27)) or (inputs(204)));
    layer0_outputs(6492) <= inputs(250);
    layer0_outputs(6493) <= not(inputs(87));
    layer0_outputs(6494) <= not(inputs(10)) or (inputs(2));
    layer0_outputs(6495) <= not((inputs(57)) xor (inputs(17)));
    layer0_outputs(6496) <= not((inputs(43)) or (inputs(158)));
    layer0_outputs(6497) <= not(inputs(90)) or (inputs(142));
    layer0_outputs(6498) <= not((inputs(245)) xor (inputs(168)));
    layer0_outputs(6499) <= (inputs(115)) and not (inputs(79));
    layer0_outputs(6500) <= not((inputs(148)) or (inputs(253)));
    layer0_outputs(6501) <= (inputs(117)) or (inputs(23));
    layer0_outputs(6502) <= (inputs(246)) and not (inputs(186));
    layer0_outputs(6503) <= not(inputs(169)) or (inputs(223));
    layer0_outputs(6504) <= not(inputs(172)) or (inputs(237));
    layer0_outputs(6505) <= not(inputs(129));
    layer0_outputs(6506) <= not(inputs(204));
    layer0_outputs(6507) <= not((inputs(225)) or (inputs(172)));
    layer0_outputs(6508) <= (inputs(246)) or (inputs(173));
    layer0_outputs(6509) <= (inputs(39)) and (inputs(22));
    layer0_outputs(6510) <= not((inputs(43)) xor (inputs(188)));
    layer0_outputs(6511) <= (inputs(13)) or (inputs(77));
    layer0_outputs(6512) <= not(inputs(72));
    layer0_outputs(6513) <= inputs(119);
    layer0_outputs(6514) <= inputs(171);
    layer0_outputs(6515) <= inputs(179);
    layer0_outputs(6516) <= inputs(122);
    layer0_outputs(6517) <= inputs(54);
    layer0_outputs(6518) <= not((inputs(218)) xor (inputs(156)));
    layer0_outputs(6519) <= not((inputs(173)) xor (inputs(229)));
    layer0_outputs(6520) <= not(inputs(178)) or (inputs(42));
    layer0_outputs(6521) <= not(inputs(90)) or (inputs(45));
    layer0_outputs(6522) <= not(inputs(183)) or (inputs(217));
    layer0_outputs(6523) <= not(inputs(168)) or (inputs(102));
    layer0_outputs(6524) <= not(inputs(40)) or (inputs(8));
    layer0_outputs(6525) <= not((inputs(186)) xor (inputs(29)));
    layer0_outputs(6526) <= not(inputs(18)) or (inputs(66));
    layer0_outputs(6527) <= not(inputs(185)) or (inputs(3));
    layer0_outputs(6528) <= (inputs(60)) and not (inputs(158));
    layer0_outputs(6529) <= not((inputs(23)) and (inputs(249)));
    layer0_outputs(6530) <= inputs(118);
    layer0_outputs(6531) <= not(inputs(16));
    layer0_outputs(6532) <= (inputs(127)) or (inputs(104));
    layer0_outputs(6533) <= (inputs(227)) or (inputs(17));
    layer0_outputs(6534) <= not(inputs(136));
    layer0_outputs(6535) <= (inputs(156)) and not (inputs(34));
    layer0_outputs(6536) <= not(inputs(187));
    layer0_outputs(6537) <= (inputs(74)) and (inputs(181));
    layer0_outputs(6538) <= (inputs(82)) or (inputs(251));
    layer0_outputs(6539) <= (inputs(131)) and not (inputs(129));
    layer0_outputs(6540) <= (inputs(61)) xor (inputs(25));
    layer0_outputs(6541) <= not((inputs(142)) or (inputs(197)));
    layer0_outputs(6542) <= (inputs(108)) and not (inputs(143));
    layer0_outputs(6543) <= not(inputs(58)) or (inputs(211));
    layer0_outputs(6544) <= not(inputs(164)) or (inputs(34));
    layer0_outputs(6545) <= not((inputs(159)) xor (inputs(212)));
    layer0_outputs(6546) <= not((inputs(211)) xor (inputs(182)));
    layer0_outputs(6547) <= (inputs(168)) and not (inputs(178));
    layer0_outputs(6548) <= not((inputs(243)) or (inputs(205)));
    layer0_outputs(6549) <= not(inputs(87)) or (inputs(173));
    layer0_outputs(6550) <= not((inputs(168)) xor (inputs(188)));
    layer0_outputs(6551) <= not((inputs(105)) or (inputs(226)));
    layer0_outputs(6552) <= not((inputs(150)) or (inputs(236)));
    layer0_outputs(6553) <= (inputs(103)) xor (inputs(196));
    layer0_outputs(6554) <= (inputs(88)) or (inputs(159));
    layer0_outputs(6555) <= not(inputs(165)) or (inputs(226));
    layer0_outputs(6556) <= not(inputs(173));
    layer0_outputs(6557) <= inputs(39);
    layer0_outputs(6558) <= (inputs(176)) or (inputs(27));
    layer0_outputs(6559) <= not((inputs(107)) or (inputs(122)));
    layer0_outputs(6560) <= '1';
    layer0_outputs(6561) <= not((inputs(51)) or (inputs(173)));
    layer0_outputs(6562) <= not(inputs(130)) or (inputs(10));
    layer0_outputs(6563) <= not((inputs(99)) or (inputs(148)));
    layer0_outputs(6564) <= not(inputs(198));
    layer0_outputs(6565) <= not(inputs(48));
    layer0_outputs(6566) <= (inputs(140)) or (inputs(166));
    layer0_outputs(6567) <= (inputs(215)) or (inputs(189));
    layer0_outputs(6568) <= not(inputs(246));
    layer0_outputs(6569) <= (inputs(170)) or (inputs(103));
    layer0_outputs(6570) <= inputs(151);
    layer0_outputs(6571) <= not((inputs(26)) xor (inputs(153)));
    layer0_outputs(6572) <= not(inputs(222));
    layer0_outputs(6573) <= not((inputs(25)) xor (inputs(226)));
    layer0_outputs(6574) <= (inputs(205)) xor (inputs(76));
    layer0_outputs(6575) <= not((inputs(84)) xor (inputs(196)));
    layer0_outputs(6576) <= inputs(24);
    layer0_outputs(6577) <= (inputs(197)) and not (inputs(159));
    layer0_outputs(6578) <= not(inputs(225));
    layer0_outputs(6579) <= inputs(91);
    layer0_outputs(6580) <= not((inputs(159)) or (inputs(171)));
    layer0_outputs(6581) <= not(inputs(152));
    layer0_outputs(6582) <= (inputs(227)) xor (inputs(79));
    layer0_outputs(6583) <= inputs(219);
    layer0_outputs(6584) <= inputs(37);
    layer0_outputs(6585) <= not((inputs(143)) and (inputs(16)));
    layer0_outputs(6586) <= '0';
    layer0_outputs(6587) <= not(inputs(140)) or (inputs(232));
    layer0_outputs(6588) <= not(inputs(76));
    layer0_outputs(6589) <= not(inputs(182)) or (inputs(45));
    layer0_outputs(6590) <= (inputs(77)) xor (inputs(60));
    layer0_outputs(6591) <= (inputs(187)) or (inputs(61));
    layer0_outputs(6592) <= not((inputs(84)) xor (inputs(214)));
    layer0_outputs(6593) <= (inputs(238)) xor (inputs(201));
    layer0_outputs(6594) <= not(inputs(217));
    layer0_outputs(6595) <= (inputs(74)) or (inputs(130));
    layer0_outputs(6596) <= not(inputs(138)) or (inputs(220));
    layer0_outputs(6597) <= inputs(44);
    layer0_outputs(6598) <= (inputs(214)) or (inputs(32));
    layer0_outputs(6599) <= (inputs(107)) or (inputs(38));
    layer0_outputs(6600) <= inputs(91);
    layer0_outputs(6601) <= (inputs(189)) and (inputs(210));
    layer0_outputs(6602) <= not((inputs(37)) or (inputs(45)));
    layer0_outputs(6603) <= not((inputs(176)) xor (inputs(151)));
    layer0_outputs(6604) <= (inputs(202)) and not (inputs(32));
    layer0_outputs(6605) <= not(inputs(92));
    layer0_outputs(6606) <= not((inputs(50)) and (inputs(25)));
    layer0_outputs(6607) <= inputs(178);
    layer0_outputs(6608) <= (inputs(35)) and not (inputs(242));
    layer0_outputs(6609) <= '1';
    layer0_outputs(6610) <= not((inputs(92)) xor (inputs(210)));
    layer0_outputs(6611) <= not(inputs(100));
    layer0_outputs(6612) <= not(inputs(171)) or (inputs(15));
    layer0_outputs(6613) <= (inputs(198)) or (inputs(157));
    layer0_outputs(6614) <= not(inputs(70));
    layer0_outputs(6615) <= (inputs(58)) or (inputs(231));
    layer0_outputs(6616) <= (inputs(21)) and not (inputs(248));
    layer0_outputs(6617) <= (inputs(146)) xor (inputs(63));
    layer0_outputs(6618) <= not(inputs(74));
    layer0_outputs(6619) <= '1';
    layer0_outputs(6620) <= not((inputs(55)) or (inputs(165)));
    layer0_outputs(6621) <= (inputs(147)) and not (inputs(15));
    layer0_outputs(6622) <= (inputs(127)) xor (inputs(58));
    layer0_outputs(6623) <= '0';
    layer0_outputs(6624) <= (inputs(77)) and not (inputs(234));
    layer0_outputs(6625) <= inputs(169);
    layer0_outputs(6626) <= (inputs(254)) xor (inputs(163));
    layer0_outputs(6627) <= (inputs(121)) and not (inputs(25));
    layer0_outputs(6628) <= (inputs(165)) and not (inputs(195));
    layer0_outputs(6629) <= not((inputs(199)) or (inputs(230)));
    layer0_outputs(6630) <= inputs(138);
    layer0_outputs(6631) <= (inputs(53)) xor (inputs(127));
    layer0_outputs(6632) <= (inputs(15)) xor (inputs(233));
    layer0_outputs(6633) <= (inputs(154)) or (inputs(65));
    layer0_outputs(6634) <= inputs(26);
    layer0_outputs(6635) <= (inputs(9)) and (inputs(202));
    layer0_outputs(6636) <= not((inputs(121)) and (inputs(70)));
    layer0_outputs(6637) <= '1';
    layer0_outputs(6638) <= inputs(91);
    layer0_outputs(6639) <= not((inputs(115)) and (inputs(115)));
    layer0_outputs(6640) <= not(inputs(22));
    layer0_outputs(6641) <= not((inputs(35)) or (inputs(61)));
    layer0_outputs(6642) <= not((inputs(43)) and (inputs(137)));
    layer0_outputs(6643) <= '0';
    layer0_outputs(6644) <= (inputs(64)) and not (inputs(248));
    layer0_outputs(6645) <= inputs(73);
    layer0_outputs(6646) <= (inputs(80)) xor (inputs(83));
    layer0_outputs(6647) <= not(inputs(114));
    layer0_outputs(6648) <= inputs(39);
    layer0_outputs(6649) <= '0';
    layer0_outputs(6650) <= not(inputs(147));
    layer0_outputs(6651) <= not((inputs(153)) or (inputs(123)));
    layer0_outputs(6652) <= (inputs(235)) or (inputs(199));
    layer0_outputs(6653) <= inputs(100);
    layer0_outputs(6654) <= not(inputs(215)) or (inputs(244));
    layer0_outputs(6655) <= not(inputs(39)) or (inputs(112));
    layer0_outputs(6656) <= (inputs(235)) and (inputs(27));
    layer0_outputs(6657) <= inputs(119);
    layer0_outputs(6658) <= not(inputs(218)) or (inputs(41));
    layer0_outputs(6659) <= not(inputs(88)) or (inputs(121));
    layer0_outputs(6660) <= not(inputs(125)) or (inputs(16));
    layer0_outputs(6661) <= (inputs(25)) xor (inputs(153));
    layer0_outputs(6662) <= (inputs(135)) xor (inputs(145));
    layer0_outputs(6663) <= (inputs(134)) and not (inputs(248));
    layer0_outputs(6664) <= (inputs(98)) and not (inputs(48));
    layer0_outputs(6665) <= not((inputs(162)) or (inputs(38)));
    layer0_outputs(6666) <= (inputs(160)) and (inputs(53));
    layer0_outputs(6667) <= not((inputs(124)) or (inputs(117)));
    layer0_outputs(6668) <= inputs(118);
    layer0_outputs(6669) <= inputs(180);
    layer0_outputs(6670) <= not(inputs(144));
    layer0_outputs(6671) <= (inputs(129)) xor (inputs(43));
    layer0_outputs(6672) <= not((inputs(162)) xor (inputs(202)));
    layer0_outputs(6673) <= not(inputs(61));
    layer0_outputs(6674) <= (inputs(103)) or (inputs(100));
    layer0_outputs(6675) <= not((inputs(164)) or (inputs(244)));
    layer0_outputs(6676) <= not((inputs(220)) and (inputs(221)));
    layer0_outputs(6677) <= (inputs(110)) or (inputs(234));
    layer0_outputs(6678) <= not((inputs(190)) xor (inputs(220)));
    layer0_outputs(6679) <= not((inputs(183)) or (inputs(87)));
    layer0_outputs(6680) <= not(inputs(93));
    layer0_outputs(6681) <= not((inputs(98)) or (inputs(184)));
    layer0_outputs(6682) <= (inputs(183)) or (inputs(11));
    layer0_outputs(6683) <= (inputs(166)) or (inputs(182));
    layer0_outputs(6684) <= (inputs(112)) or (inputs(208));
    layer0_outputs(6685) <= not((inputs(162)) xor (inputs(160)));
    layer0_outputs(6686) <= not(inputs(182));
    layer0_outputs(6687) <= (inputs(137)) xor (inputs(156));
    layer0_outputs(6688) <= not((inputs(222)) xor (inputs(38)));
    layer0_outputs(6689) <= not(inputs(97)) or (inputs(216));
    layer0_outputs(6690) <= (inputs(166)) and not (inputs(89));
    layer0_outputs(6691) <= (inputs(84)) or (inputs(241));
    layer0_outputs(6692) <= not((inputs(96)) xor (inputs(85)));
    layer0_outputs(6693) <= (inputs(37)) and not (inputs(0));
    layer0_outputs(6694) <= not(inputs(190)) or (inputs(159));
    layer0_outputs(6695) <= not(inputs(43)) or (inputs(210));
    layer0_outputs(6696) <= (inputs(93)) and not (inputs(146));
    layer0_outputs(6697) <= '0';
    layer0_outputs(6698) <= inputs(56);
    layer0_outputs(6699) <= inputs(72);
    layer0_outputs(6700) <= not(inputs(158));
    layer0_outputs(6701) <= (inputs(14)) xor (inputs(34));
    layer0_outputs(6702) <= inputs(231);
    layer0_outputs(6703) <= (inputs(112)) xor (inputs(62));
    layer0_outputs(6704) <= not(inputs(248)) or (inputs(29));
    layer0_outputs(6705) <= inputs(10);
    layer0_outputs(6706) <= not(inputs(108));
    layer0_outputs(6707) <= (inputs(37)) and not (inputs(11));
    layer0_outputs(6708) <= not(inputs(138));
    layer0_outputs(6709) <= inputs(113);
    layer0_outputs(6710) <= inputs(168);
    layer0_outputs(6711) <= (inputs(134)) and (inputs(60));
    layer0_outputs(6712) <= (inputs(175)) xor (inputs(73));
    layer0_outputs(6713) <= (inputs(131)) or (inputs(43));
    layer0_outputs(6714) <= (inputs(135)) or (inputs(68));
    layer0_outputs(6715) <= (inputs(120)) and not (inputs(33));
    layer0_outputs(6716) <= not(inputs(98)) or (inputs(80));
    layer0_outputs(6717) <= (inputs(153)) or (inputs(114));
    layer0_outputs(6718) <= inputs(167);
    layer0_outputs(6719) <= not(inputs(241));
    layer0_outputs(6720) <= not((inputs(73)) or (inputs(112)));
    layer0_outputs(6721) <= '1';
    layer0_outputs(6722) <= '0';
    layer0_outputs(6723) <= (inputs(187)) or (inputs(53));
    layer0_outputs(6724) <= not((inputs(21)) or (inputs(166)));
    layer0_outputs(6725) <= not(inputs(182));
    layer0_outputs(6726) <= (inputs(25)) and not (inputs(155));
    layer0_outputs(6727) <= (inputs(132)) and not (inputs(211));
    layer0_outputs(6728) <= not(inputs(18)) or (inputs(53));
    layer0_outputs(6729) <= not((inputs(48)) xor (inputs(179)));
    layer0_outputs(6730) <= not(inputs(102));
    layer0_outputs(6731) <= (inputs(117)) and not (inputs(8));
    layer0_outputs(6732) <= not(inputs(91));
    layer0_outputs(6733) <= not(inputs(171)) or (inputs(96));
    layer0_outputs(6734) <= inputs(177);
    layer0_outputs(6735) <= not((inputs(178)) and (inputs(227)));
    layer0_outputs(6736) <= '1';
    layer0_outputs(6737) <= inputs(22);
    layer0_outputs(6738) <= not((inputs(228)) xor (inputs(24)));
    layer0_outputs(6739) <= inputs(214);
    layer0_outputs(6740) <= (inputs(91)) and not (inputs(41));
    layer0_outputs(6741) <= not(inputs(4)) or (inputs(161));
    layer0_outputs(6742) <= (inputs(119)) xor (inputs(235));
    layer0_outputs(6743) <= not(inputs(82));
    layer0_outputs(6744) <= (inputs(183)) or (inputs(171));
    layer0_outputs(6745) <= inputs(150);
    layer0_outputs(6746) <= not(inputs(212)) or (inputs(42));
    layer0_outputs(6747) <= not((inputs(8)) xor (inputs(80)));
    layer0_outputs(6748) <= not((inputs(204)) or (inputs(4)));
    layer0_outputs(6749) <= not(inputs(136));
    layer0_outputs(6750) <= not(inputs(68)) or (inputs(170));
    layer0_outputs(6751) <= not(inputs(215)) or (inputs(207));
    layer0_outputs(6752) <= (inputs(199)) or (inputs(216));
    layer0_outputs(6753) <= not((inputs(43)) xor (inputs(155)));
    layer0_outputs(6754) <= not(inputs(169)) or (inputs(75));
    layer0_outputs(6755) <= not(inputs(10));
    layer0_outputs(6756) <= inputs(152);
    layer0_outputs(6757) <= not((inputs(85)) or (inputs(21)));
    layer0_outputs(6758) <= not((inputs(108)) or (inputs(232)));
    layer0_outputs(6759) <= (inputs(156)) and not (inputs(253));
    layer0_outputs(6760) <= (inputs(108)) or (inputs(49));
    layer0_outputs(6761) <= not((inputs(68)) xor (inputs(187)));
    layer0_outputs(6762) <= (inputs(201)) and not (inputs(126));
    layer0_outputs(6763) <= not(inputs(225)) or (inputs(111));
    layer0_outputs(6764) <= not((inputs(45)) xor (inputs(78)));
    layer0_outputs(6765) <= not(inputs(229));
    layer0_outputs(6766) <= (inputs(165)) and not (inputs(243));
    layer0_outputs(6767) <= not(inputs(197)) or (inputs(169));
    layer0_outputs(6768) <= (inputs(23)) or (inputs(15));
    layer0_outputs(6769) <= inputs(231);
    layer0_outputs(6770) <= not(inputs(26)) or (inputs(182));
    layer0_outputs(6771) <= (inputs(59)) and not (inputs(244));
    layer0_outputs(6772) <= not((inputs(71)) and (inputs(49)));
    layer0_outputs(6773) <= (inputs(169)) and not (inputs(80));
    layer0_outputs(6774) <= inputs(151);
    layer0_outputs(6775) <= (inputs(136)) and not (inputs(249));
    layer0_outputs(6776) <= not(inputs(212));
    layer0_outputs(6777) <= not(inputs(104));
    layer0_outputs(6778) <= (inputs(205)) or (inputs(167));
    layer0_outputs(6779) <= not(inputs(118)) or (inputs(168));
    layer0_outputs(6780) <= (inputs(197)) or (inputs(190));
    layer0_outputs(6781) <= not((inputs(179)) or (inputs(246)));
    layer0_outputs(6782) <= (inputs(2)) or (inputs(29));
    layer0_outputs(6783) <= (inputs(72)) or (inputs(127));
    layer0_outputs(6784) <= (inputs(77)) or (inputs(204));
    layer0_outputs(6785) <= not(inputs(150)) or (inputs(243));
    layer0_outputs(6786) <= (inputs(102)) xor (inputs(210));
    layer0_outputs(6787) <= (inputs(220)) xor (inputs(233));
    layer0_outputs(6788) <= (inputs(156)) xor (inputs(207));
    layer0_outputs(6789) <= (inputs(123)) and not (inputs(236));
    layer0_outputs(6790) <= not((inputs(211)) or (inputs(104)));
    layer0_outputs(6791) <= not((inputs(49)) xor (inputs(93)));
    layer0_outputs(6792) <= inputs(168);
    layer0_outputs(6793) <= not(inputs(129)) or (inputs(143));
    layer0_outputs(6794) <= (inputs(217)) xor (inputs(95));
    layer0_outputs(6795) <= not((inputs(187)) or (inputs(197)));
    layer0_outputs(6796) <= inputs(218);
    layer0_outputs(6797) <= not((inputs(96)) xor (inputs(119)));
    layer0_outputs(6798) <= not((inputs(210)) xor (inputs(175)));
    layer0_outputs(6799) <= (inputs(44)) xor (inputs(52));
    layer0_outputs(6800) <= inputs(55);
    layer0_outputs(6801) <= (inputs(95)) xor (inputs(221));
    layer0_outputs(6802) <= (inputs(252)) or (inputs(164));
    layer0_outputs(6803) <= (inputs(227)) and not (inputs(46));
    layer0_outputs(6804) <= (inputs(90)) or (inputs(110));
    layer0_outputs(6805) <= (inputs(128)) and not (inputs(35));
    layer0_outputs(6806) <= not((inputs(250)) and (inputs(66)));
    layer0_outputs(6807) <= (inputs(131)) and not (inputs(162));
    layer0_outputs(6808) <= (inputs(25)) and not (inputs(6));
    layer0_outputs(6809) <= (inputs(184)) and not (inputs(217));
    layer0_outputs(6810) <= inputs(135);
    layer0_outputs(6811) <= inputs(17);
    layer0_outputs(6812) <= (inputs(79)) xor (inputs(141));
    layer0_outputs(6813) <= (inputs(228)) or (inputs(89));
    layer0_outputs(6814) <= not(inputs(79)) or (inputs(209));
    layer0_outputs(6815) <= not(inputs(68)) or (inputs(6));
    layer0_outputs(6816) <= not((inputs(69)) and (inputs(245)));
    layer0_outputs(6817) <= (inputs(128)) or (inputs(6));
    layer0_outputs(6818) <= inputs(156);
    layer0_outputs(6819) <= (inputs(226)) xor (inputs(165));
    layer0_outputs(6820) <= inputs(149);
    layer0_outputs(6821) <= (inputs(170)) or (inputs(156));
    layer0_outputs(6822) <= (inputs(120)) or (inputs(67));
    layer0_outputs(6823) <= (inputs(3)) xor (inputs(174));
    layer0_outputs(6824) <= not(inputs(69));
    layer0_outputs(6825) <= not((inputs(54)) xor (inputs(17)));
    layer0_outputs(6826) <= not(inputs(6));
    layer0_outputs(6827) <= inputs(216);
    layer0_outputs(6828) <= not((inputs(213)) or (inputs(95)));
    layer0_outputs(6829) <= not(inputs(56)) or (inputs(229));
    layer0_outputs(6830) <= (inputs(34)) and not (inputs(35));
    layer0_outputs(6831) <= not((inputs(233)) or (inputs(255)));
    layer0_outputs(6832) <= not((inputs(248)) and (inputs(87)));
    layer0_outputs(6833) <= not(inputs(167)) or (inputs(11));
    layer0_outputs(6834) <= inputs(170);
    layer0_outputs(6835) <= not((inputs(82)) and (inputs(18)));
    layer0_outputs(6836) <= (inputs(5)) or (inputs(61));
    layer0_outputs(6837) <= not(inputs(127));
    layer0_outputs(6838) <= (inputs(121)) or (inputs(131));
    layer0_outputs(6839) <= not((inputs(141)) xor (inputs(135)));
    layer0_outputs(6840) <= not(inputs(61));
    layer0_outputs(6841) <= (inputs(115)) and not (inputs(20));
    layer0_outputs(6842) <= not((inputs(219)) or (inputs(51)));
    layer0_outputs(6843) <= not(inputs(185));
    layer0_outputs(6844) <= (inputs(171)) or (inputs(158));
    layer0_outputs(6845) <= inputs(37);
    layer0_outputs(6846) <= (inputs(144)) or (inputs(216));
    layer0_outputs(6847) <= (inputs(224)) and (inputs(129));
    layer0_outputs(6848) <= (inputs(51)) xor (inputs(97));
    layer0_outputs(6849) <= (inputs(180)) and not (inputs(113));
    layer0_outputs(6850) <= (inputs(209)) xor (inputs(106));
    layer0_outputs(6851) <= not(inputs(148)) or (inputs(203));
    layer0_outputs(6852) <= not((inputs(250)) or (inputs(140)));
    layer0_outputs(6853) <= not(inputs(239)) or (inputs(0));
    layer0_outputs(6854) <= not((inputs(15)) xor (inputs(202)));
    layer0_outputs(6855) <= (inputs(30)) xor (inputs(79));
    layer0_outputs(6856) <= (inputs(49)) and not (inputs(16));
    layer0_outputs(6857) <= (inputs(137)) and not (inputs(201));
    layer0_outputs(6858) <= (inputs(164)) xor (inputs(135));
    layer0_outputs(6859) <= not(inputs(107)) or (inputs(141));
    layer0_outputs(6860) <= not((inputs(120)) xor (inputs(171)));
    layer0_outputs(6861) <= not((inputs(242)) xor (inputs(185)));
    layer0_outputs(6862) <= (inputs(83)) xor (inputs(2));
    layer0_outputs(6863) <= not((inputs(144)) or (inputs(84)));
    layer0_outputs(6864) <= (inputs(159)) and not (inputs(113));
    layer0_outputs(6865) <= not(inputs(86));
    layer0_outputs(6866) <= not(inputs(174)) or (inputs(111));
    layer0_outputs(6867) <= inputs(200);
    layer0_outputs(6868) <= inputs(109);
    layer0_outputs(6869) <= not((inputs(203)) or (inputs(86)));
    layer0_outputs(6870) <= inputs(149);
    layer0_outputs(6871) <= inputs(139);
    layer0_outputs(6872) <= not(inputs(104)) or (inputs(232));
    layer0_outputs(6873) <= (inputs(205)) xor (inputs(247));
    layer0_outputs(6874) <= not(inputs(180)) or (inputs(208));
    layer0_outputs(6875) <= not((inputs(194)) or (inputs(200)));
    layer0_outputs(6876) <= not((inputs(223)) or (inputs(31)));
    layer0_outputs(6877) <= not((inputs(40)) xor (inputs(223)));
    layer0_outputs(6878) <= not(inputs(36)) or (inputs(237));
    layer0_outputs(6879) <= inputs(70);
    layer0_outputs(6880) <= not(inputs(5));
    layer0_outputs(6881) <= not(inputs(30)) or (inputs(26));
    layer0_outputs(6882) <= (inputs(123)) and not (inputs(37));
    layer0_outputs(6883) <= not(inputs(165)) or (inputs(218));
    layer0_outputs(6884) <= not(inputs(231));
    layer0_outputs(6885) <= (inputs(147)) or (inputs(229));
    layer0_outputs(6886) <= inputs(157);
    layer0_outputs(6887) <= not(inputs(106));
    layer0_outputs(6888) <= (inputs(203)) and not (inputs(63));
    layer0_outputs(6889) <= (inputs(228)) xor (inputs(107));
    layer0_outputs(6890) <= inputs(190);
    layer0_outputs(6891) <= (inputs(147)) and not (inputs(30));
    layer0_outputs(6892) <= not(inputs(198));
    layer0_outputs(6893) <= '1';
    layer0_outputs(6894) <= not(inputs(230)) or (inputs(82));
    layer0_outputs(6895) <= not((inputs(145)) or (inputs(59)));
    layer0_outputs(6896) <= not(inputs(55));
    layer0_outputs(6897) <= not(inputs(154));
    layer0_outputs(6898) <= (inputs(200)) xor (inputs(247));
    layer0_outputs(6899) <= not((inputs(46)) xor (inputs(188)));
    layer0_outputs(6900) <= (inputs(213)) or (inputs(250));
    layer0_outputs(6901) <= not(inputs(89));
    layer0_outputs(6902) <= not(inputs(182));
    layer0_outputs(6903) <= (inputs(66)) or (inputs(113));
    layer0_outputs(6904) <= not(inputs(19));
    layer0_outputs(6905) <= not((inputs(165)) or (inputs(199)));
    layer0_outputs(6906) <= (inputs(86)) and not (inputs(107));
    layer0_outputs(6907) <= (inputs(114)) and (inputs(255));
    layer0_outputs(6908) <= not(inputs(167)) or (inputs(9));
    layer0_outputs(6909) <= (inputs(72)) and (inputs(122));
    layer0_outputs(6910) <= not(inputs(200)) or (inputs(83));
    layer0_outputs(6911) <= not((inputs(64)) and (inputs(188)));
    layer0_outputs(6912) <= (inputs(184)) and not (inputs(205));
    layer0_outputs(6913) <= (inputs(128)) or (inputs(128));
    layer0_outputs(6914) <= (inputs(177)) or (inputs(182));
    layer0_outputs(6915) <= (inputs(189)) and not (inputs(244));
    layer0_outputs(6916) <= not((inputs(148)) xor (inputs(48)));
    layer0_outputs(6917) <= not(inputs(84)) or (inputs(20));
    layer0_outputs(6918) <= not(inputs(46));
    layer0_outputs(6919) <= (inputs(114)) or (inputs(248));
    layer0_outputs(6920) <= not((inputs(193)) and (inputs(96)));
    layer0_outputs(6921) <= not((inputs(252)) or (inputs(181)));
    layer0_outputs(6922) <= not(inputs(46));
    layer0_outputs(6923) <= not((inputs(208)) or (inputs(114)));
    layer0_outputs(6924) <= (inputs(56)) or (inputs(154));
    layer0_outputs(6925) <= not(inputs(198));
    layer0_outputs(6926) <= (inputs(87)) and not (inputs(221));
    layer0_outputs(6927) <= not((inputs(92)) or (inputs(141)));
    layer0_outputs(6928) <= not(inputs(58));
    layer0_outputs(6929) <= (inputs(189)) xor (inputs(156));
    layer0_outputs(6930) <= not((inputs(43)) or (inputs(193)));
    layer0_outputs(6931) <= (inputs(176)) and not (inputs(7));
    layer0_outputs(6932) <= not(inputs(162)) or (inputs(97));
    layer0_outputs(6933) <= not((inputs(240)) xor (inputs(185)));
    layer0_outputs(6934) <= not((inputs(113)) and (inputs(117)));
    layer0_outputs(6935) <= (inputs(80)) or (inputs(230));
    layer0_outputs(6936) <= not(inputs(172)) or (inputs(130));
    layer0_outputs(6937) <= not((inputs(213)) xor (inputs(125)));
    layer0_outputs(6938) <= (inputs(247)) xor (inputs(43));
    layer0_outputs(6939) <= '1';
    layer0_outputs(6940) <= (inputs(60)) or (inputs(208));
    layer0_outputs(6941) <= not(inputs(70));
    layer0_outputs(6942) <= not((inputs(101)) or (inputs(190)));
    layer0_outputs(6943) <= not(inputs(27)) or (inputs(235));
    layer0_outputs(6944) <= (inputs(152)) and not (inputs(90));
    layer0_outputs(6945) <= not((inputs(206)) or (inputs(186)));
    layer0_outputs(6946) <= (inputs(213)) and not (inputs(91));
    layer0_outputs(6947) <= (inputs(186)) and not (inputs(252));
    layer0_outputs(6948) <= (inputs(73)) xor (inputs(28));
    layer0_outputs(6949) <= not((inputs(141)) xor (inputs(161)));
    layer0_outputs(6950) <= not(inputs(214));
    layer0_outputs(6951) <= (inputs(213)) and not (inputs(66));
    layer0_outputs(6952) <= not((inputs(183)) xor (inputs(193)));
    layer0_outputs(6953) <= (inputs(23)) or (inputs(68));
    layer0_outputs(6954) <= (inputs(189)) or (inputs(197));
    layer0_outputs(6955) <= not(inputs(137));
    layer0_outputs(6956) <= inputs(100);
    layer0_outputs(6957) <= '0';
    layer0_outputs(6958) <= not((inputs(230)) xor (inputs(34)));
    layer0_outputs(6959) <= (inputs(95)) or (inputs(199));
    layer0_outputs(6960) <= (inputs(3)) or (inputs(172));
    layer0_outputs(6961) <= not(inputs(47));
    layer0_outputs(6962) <= (inputs(129)) xor (inputs(211));
    layer0_outputs(6963) <= (inputs(173)) xor (inputs(2));
    layer0_outputs(6964) <= (inputs(209)) and not (inputs(254));
    layer0_outputs(6965) <= not(inputs(105));
    layer0_outputs(6966) <= not((inputs(110)) or (inputs(99)));
    layer0_outputs(6967) <= not(inputs(66));
    layer0_outputs(6968) <= not(inputs(228));
    layer0_outputs(6969) <= '0';
    layer0_outputs(6970) <= not(inputs(157)) or (inputs(248));
    layer0_outputs(6971) <= not(inputs(27));
    layer0_outputs(6972) <= (inputs(103)) and (inputs(121));
    layer0_outputs(6973) <= (inputs(224)) xor (inputs(8));
    layer0_outputs(6974) <= not((inputs(23)) and (inputs(112)));
    layer0_outputs(6975) <= not((inputs(103)) or (inputs(170)));
    layer0_outputs(6976) <= '1';
    layer0_outputs(6977) <= (inputs(115)) and (inputs(1));
    layer0_outputs(6978) <= not((inputs(254)) and (inputs(67)));
    layer0_outputs(6979) <= not(inputs(254)) or (inputs(5));
    layer0_outputs(6980) <= (inputs(243)) xor (inputs(99));
    layer0_outputs(6981) <= (inputs(217)) xor (inputs(145));
    layer0_outputs(6982) <= (inputs(132)) xor (inputs(68));
    layer0_outputs(6983) <= not(inputs(122));
    layer0_outputs(6984) <= not(inputs(140));
    layer0_outputs(6985) <= (inputs(209)) and not (inputs(143));
    layer0_outputs(6986) <= not((inputs(201)) xor (inputs(93)));
    layer0_outputs(6987) <= not(inputs(155)) or (inputs(115));
    layer0_outputs(6988) <= not((inputs(153)) or (inputs(83)));
    layer0_outputs(6989) <= (inputs(38)) or (inputs(129));
    layer0_outputs(6990) <= not(inputs(153)) or (inputs(18));
    layer0_outputs(6991) <= inputs(65);
    layer0_outputs(6992) <= (inputs(195)) and not (inputs(219));
    layer0_outputs(6993) <= not(inputs(120));
    layer0_outputs(6994) <= inputs(71);
    layer0_outputs(6995) <= (inputs(122)) and not (inputs(92));
    layer0_outputs(6996) <= (inputs(59)) and not (inputs(44));
    layer0_outputs(6997) <= inputs(52);
    layer0_outputs(6998) <= '1';
    layer0_outputs(6999) <= (inputs(56)) or (inputs(223));
    layer0_outputs(7000) <= inputs(127);
    layer0_outputs(7001) <= not((inputs(12)) or (inputs(43)));
    layer0_outputs(7002) <= not((inputs(74)) or (inputs(68)));
    layer0_outputs(7003) <= (inputs(127)) xor (inputs(206));
    layer0_outputs(7004) <= not(inputs(169)) or (inputs(77));
    layer0_outputs(7005) <= '0';
    layer0_outputs(7006) <= not(inputs(38)) or (inputs(34));
    layer0_outputs(7007) <= not(inputs(87)) or (inputs(244));
    layer0_outputs(7008) <= not((inputs(191)) or (inputs(40)));
    layer0_outputs(7009) <= not(inputs(4)) or (inputs(238));
    layer0_outputs(7010) <= not((inputs(240)) or (inputs(234)));
    layer0_outputs(7011) <= not(inputs(121));
    layer0_outputs(7012) <= (inputs(169)) or (inputs(138));
    layer0_outputs(7013) <= not((inputs(174)) and (inputs(159)));
    layer0_outputs(7014) <= not(inputs(184)) or (inputs(139));
    layer0_outputs(7015) <= not(inputs(119));
    layer0_outputs(7016) <= not(inputs(104));
    layer0_outputs(7017) <= not((inputs(182)) or (inputs(72)));
    layer0_outputs(7018) <= not((inputs(0)) xor (inputs(217)));
    layer0_outputs(7019) <= not((inputs(91)) xor (inputs(66)));
    layer0_outputs(7020) <= (inputs(131)) and not (inputs(58));
    layer0_outputs(7021) <= not((inputs(164)) xor (inputs(213)));
    layer0_outputs(7022) <= not(inputs(122));
    layer0_outputs(7023) <= (inputs(153)) and not (inputs(151));
    layer0_outputs(7024) <= (inputs(37)) and not (inputs(63));
    layer0_outputs(7025) <= not((inputs(247)) or (inputs(142)));
    layer0_outputs(7026) <= (inputs(24)) xor (inputs(193));
    layer0_outputs(7027) <= (inputs(121)) or (inputs(203));
    layer0_outputs(7028) <= (inputs(101)) and not (inputs(60));
    layer0_outputs(7029) <= not(inputs(183));
    layer0_outputs(7030) <= (inputs(206)) xor (inputs(99));
    layer0_outputs(7031) <= not((inputs(175)) or (inputs(134)));
    layer0_outputs(7032) <= (inputs(13)) and not (inputs(248));
    layer0_outputs(7033) <= '0';
    layer0_outputs(7034) <= (inputs(3)) and (inputs(144));
    layer0_outputs(7035) <= not((inputs(142)) xor (inputs(149)));
    layer0_outputs(7036) <= not((inputs(74)) or (inputs(187)));
    layer0_outputs(7037) <= (inputs(244)) xor (inputs(221));
    layer0_outputs(7038) <= (inputs(0)) and (inputs(223));
    layer0_outputs(7039) <= not(inputs(100));
    layer0_outputs(7040) <= (inputs(153)) xor (inputs(113));
    layer0_outputs(7041) <= not(inputs(201));
    layer0_outputs(7042) <= (inputs(49)) or (inputs(124));
    layer0_outputs(7043) <= not((inputs(205)) or (inputs(180)));
    layer0_outputs(7044) <= (inputs(59)) and not (inputs(114));
    layer0_outputs(7045) <= not(inputs(9));
    layer0_outputs(7046) <= inputs(96);
    layer0_outputs(7047) <= not((inputs(175)) and (inputs(112)));
    layer0_outputs(7048) <= not(inputs(105));
    layer0_outputs(7049) <= not(inputs(53)) or (inputs(11));
    layer0_outputs(7050) <= (inputs(114)) and not (inputs(248));
    layer0_outputs(7051) <= not((inputs(120)) or (inputs(234)));
    layer0_outputs(7052) <= not(inputs(16)) or (inputs(44));
    layer0_outputs(7053) <= not(inputs(75));
    layer0_outputs(7054) <= not(inputs(29));
    layer0_outputs(7055) <= (inputs(85)) xor (inputs(51));
    layer0_outputs(7056) <= not((inputs(47)) or (inputs(247)));
    layer0_outputs(7057) <= (inputs(119)) or (inputs(160));
    layer0_outputs(7058) <= not((inputs(20)) and (inputs(174)));
    layer0_outputs(7059) <= (inputs(135)) and not (inputs(237));
    layer0_outputs(7060) <= (inputs(57)) or (inputs(97));
    layer0_outputs(7061) <= (inputs(83)) or (inputs(11));
    layer0_outputs(7062) <= (inputs(60)) or (inputs(97));
    layer0_outputs(7063) <= '0';
    layer0_outputs(7064) <= not((inputs(34)) or (inputs(221)));
    layer0_outputs(7065) <= inputs(85);
    layer0_outputs(7066) <= (inputs(151)) or (inputs(95));
    layer0_outputs(7067) <= (inputs(152)) xor (inputs(237));
    layer0_outputs(7068) <= inputs(107);
    layer0_outputs(7069) <= not((inputs(106)) or (inputs(105)));
    layer0_outputs(7070) <= inputs(121);
    layer0_outputs(7071) <= '0';
    layer0_outputs(7072) <= inputs(138);
    layer0_outputs(7073) <= not(inputs(12));
    layer0_outputs(7074) <= (inputs(144)) xor (inputs(26));
    layer0_outputs(7075) <= (inputs(134)) and not (inputs(246));
    layer0_outputs(7076) <= not(inputs(220));
    layer0_outputs(7077) <= (inputs(118)) and not (inputs(139));
    layer0_outputs(7078) <= '1';
    layer0_outputs(7079) <= (inputs(163)) and not (inputs(23));
    layer0_outputs(7080) <= not((inputs(203)) or (inputs(220)));
    layer0_outputs(7081) <= not(inputs(61));
    layer0_outputs(7082) <= (inputs(40)) or (inputs(203));
    layer0_outputs(7083) <= (inputs(94)) and not (inputs(226));
    layer0_outputs(7084) <= (inputs(213)) and not (inputs(111));
    layer0_outputs(7085) <= '0';
    layer0_outputs(7086) <= not(inputs(165));
    layer0_outputs(7087) <= (inputs(108)) and not (inputs(145));
    layer0_outputs(7088) <= not(inputs(140)) or (inputs(129));
    layer0_outputs(7089) <= not((inputs(20)) or (inputs(200)));
    layer0_outputs(7090) <= not((inputs(77)) or (inputs(231)));
    layer0_outputs(7091) <= not((inputs(50)) xor (inputs(161)));
    layer0_outputs(7092) <= not(inputs(206));
    layer0_outputs(7093) <= inputs(133);
    layer0_outputs(7094) <= not((inputs(148)) or (inputs(56)));
    layer0_outputs(7095) <= (inputs(50)) xor (inputs(215));
    layer0_outputs(7096) <= (inputs(165)) and not (inputs(64));
    layer0_outputs(7097) <= (inputs(7)) and (inputs(62));
    layer0_outputs(7098) <= inputs(117);
    layer0_outputs(7099) <= not(inputs(41)) or (inputs(246));
    layer0_outputs(7100) <= (inputs(200)) or (inputs(243));
    layer0_outputs(7101) <= (inputs(101)) and not (inputs(208));
    layer0_outputs(7102) <= not(inputs(76)) or (inputs(243));
    layer0_outputs(7103) <= inputs(164);
    layer0_outputs(7104) <= (inputs(101)) and not (inputs(227));
    layer0_outputs(7105) <= not(inputs(203)) or (inputs(178));
    layer0_outputs(7106) <= not(inputs(132)) or (inputs(71));
    layer0_outputs(7107) <= '0';
    layer0_outputs(7108) <= inputs(133);
    layer0_outputs(7109) <= (inputs(104)) and not (inputs(230));
    layer0_outputs(7110) <= not(inputs(42)) or (inputs(47));
    layer0_outputs(7111) <= not((inputs(61)) xor (inputs(110)));
    layer0_outputs(7112) <= not(inputs(189)) or (inputs(239));
    layer0_outputs(7113) <= '1';
    layer0_outputs(7114) <= (inputs(15)) xor (inputs(57));
    layer0_outputs(7115) <= not((inputs(249)) and (inputs(119)));
    layer0_outputs(7116) <= not(inputs(97));
    layer0_outputs(7117) <= not(inputs(205));
    layer0_outputs(7118) <= not(inputs(107));
    layer0_outputs(7119) <= (inputs(192)) xor (inputs(86));
    layer0_outputs(7120) <= not(inputs(121)) or (inputs(225));
    layer0_outputs(7121) <= '0';
    layer0_outputs(7122) <= not((inputs(122)) xor (inputs(36)));
    layer0_outputs(7123) <= not((inputs(45)) or (inputs(105)));
    layer0_outputs(7124) <= not(inputs(104));
    layer0_outputs(7125) <= (inputs(121)) and not (inputs(78));
    layer0_outputs(7126) <= not((inputs(7)) or (inputs(181)));
    layer0_outputs(7127) <= (inputs(179)) xor (inputs(79));
    layer0_outputs(7128) <= not((inputs(248)) or (inputs(115)));
    layer0_outputs(7129) <= (inputs(50)) or (inputs(43));
    layer0_outputs(7130) <= (inputs(213)) and not (inputs(6));
    layer0_outputs(7131) <= (inputs(70)) or (inputs(83));
    layer0_outputs(7132) <= inputs(186);
    layer0_outputs(7133) <= (inputs(248)) and not (inputs(209));
    layer0_outputs(7134) <= inputs(57);
    layer0_outputs(7135) <= (inputs(172)) or (inputs(214));
    layer0_outputs(7136) <= not(inputs(191));
    layer0_outputs(7137) <= inputs(170);
    layer0_outputs(7138) <= '0';
    layer0_outputs(7139) <= not(inputs(46));
    layer0_outputs(7140) <= inputs(201);
    layer0_outputs(7141) <= (inputs(156)) xor (inputs(110));
    layer0_outputs(7142) <= not(inputs(133)) or (inputs(219));
    layer0_outputs(7143) <= not(inputs(117));
    layer0_outputs(7144) <= (inputs(87)) xor (inputs(99));
    layer0_outputs(7145) <= not((inputs(134)) or (inputs(44)));
    layer0_outputs(7146) <= not((inputs(194)) xor (inputs(17)));
    layer0_outputs(7147) <= (inputs(160)) and not (inputs(221));
    layer0_outputs(7148) <= (inputs(85)) xor (inputs(148));
    layer0_outputs(7149) <= (inputs(22)) and (inputs(8));
    layer0_outputs(7150) <= not(inputs(128)) or (inputs(208));
    layer0_outputs(7151) <= not((inputs(162)) or (inputs(233)));
    layer0_outputs(7152) <= inputs(134);
    layer0_outputs(7153) <= not((inputs(142)) xor (inputs(198)));
    layer0_outputs(7154) <= not((inputs(219)) or (inputs(251)));
    layer0_outputs(7155) <= not((inputs(170)) or (inputs(60)));
    layer0_outputs(7156) <= not(inputs(64));
    layer0_outputs(7157) <= (inputs(46)) or (inputs(120));
    layer0_outputs(7158) <= not(inputs(54));
    layer0_outputs(7159) <= not((inputs(31)) xor (inputs(100)));
    layer0_outputs(7160) <= (inputs(206)) and not (inputs(0));
    layer0_outputs(7161) <= not(inputs(119)) or (inputs(65));
    layer0_outputs(7162) <= inputs(118);
    layer0_outputs(7163) <= (inputs(241)) or (inputs(103));
    layer0_outputs(7164) <= (inputs(26)) xor (inputs(101));
    layer0_outputs(7165) <= not(inputs(88)) or (inputs(21));
    layer0_outputs(7166) <= (inputs(76)) and not (inputs(169));
    layer0_outputs(7167) <= not(inputs(194));
    layer0_outputs(7168) <= (inputs(127)) and (inputs(41));
    layer0_outputs(7169) <= inputs(136);
    layer0_outputs(7170) <= (inputs(124)) xor (inputs(209));
    layer0_outputs(7171) <= (inputs(63)) xor (inputs(78));
    layer0_outputs(7172) <= inputs(100);
    layer0_outputs(7173) <= not((inputs(249)) and (inputs(166)));
    layer0_outputs(7174) <= not(inputs(118));
    layer0_outputs(7175) <= (inputs(174)) and (inputs(221));
    layer0_outputs(7176) <= (inputs(210)) and not (inputs(114));
    layer0_outputs(7177) <= not(inputs(136));
    layer0_outputs(7178) <= (inputs(102)) xor (inputs(193));
    layer0_outputs(7179) <= (inputs(82)) xor (inputs(45));
    layer0_outputs(7180) <= not(inputs(155));
    layer0_outputs(7181) <= not((inputs(30)) and (inputs(79)));
    layer0_outputs(7182) <= (inputs(229)) or (inputs(155));
    layer0_outputs(7183) <= not((inputs(64)) xor (inputs(37)));
    layer0_outputs(7184) <= (inputs(162)) or (inputs(103));
    layer0_outputs(7185) <= not(inputs(178));
    layer0_outputs(7186) <= inputs(26);
    layer0_outputs(7187) <= (inputs(163)) and not (inputs(45));
    layer0_outputs(7188) <= not((inputs(146)) or (inputs(114)));
    layer0_outputs(7189) <= not((inputs(61)) xor (inputs(209)));
    layer0_outputs(7190) <= (inputs(44)) xor (inputs(131));
    layer0_outputs(7191) <= '1';
    layer0_outputs(7192) <= not((inputs(55)) or (inputs(248)));
    layer0_outputs(7193) <= not(inputs(27)) or (inputs(63));
    layer0_outputs(7194) <= not(inputs(180)) or (inputs(129));
    layer0_outputs(7195) <= '1';
    layer0_outputs(7196) <= (inputs(16)) and not (inputs(30));
    layer0_outputs(7197) <= not(inputs(251));
    layer0_outputs(7198) <= not((inputs(26)) or (inputs(226)));
    layer0_outputs(7199) <= not((inputs(215)) xor (inputs(255)));
    layer0_outputs(7200) <= not((inputs(125)) or (inputs(181)));
    layer0_outputs(7201) <= not((inputs(222)) or (inputs(45)));
    layer0_outputs(7202) <= not(inputs(108));
    layer0_outputs(7203) <= not(inputs(236)) or (inputs(11));
    layer0_outputs(7204) <= (inputs(29)) and not (inputs(114));
    layer0_outputs(7205) <= not((inputs(133)) xor (inputs(58)));
    layer0_outputs(7206) <= not(inputs(151));
    layer0_outputs(7207) <= '0';
    layer0_outputs(7208) <= inputs(111);
    layer0_outputs(7209) <= (inputs(10)) xor (inputs(89));
    layer0_outputs(7210) <= (inputs(177)) xor (inputs(16));
    layer0_outputs(7211) <= (inputs(141)) and not (inputs(239));
    layer0_outputs(7212) <= not((inputs(150)) xor (inputs(243)));
    layer0_outputs(7213) <= not(inputs(85)) or (inputs(168));
    layer0_outputs(7214) <= (inputs(212)) and (inputs(56));
    layer0_outputs(7215) <= '1';
    layer0_outputs(7216) <= (inputs(187)) xor (inputs(25));
    layer0_outputs(7217) <= not((inputs(42)) or (inputs(20)));
    layer0_outputs(7218) <= (inputs(91)) and not (inputs(22));
    layer0_outputs(7219) <= (inputs(242)) xor (inputs(165));
    layer0_outputs(7220) <= inputs(111);
    layer0_outputs(7221) <= not(inputs(241));
    layer0_outputs(7222) <= not(inputs(9));
    layer0_outputs(7223) <= (inputs(84)) or (inputs(244));
    layer0_outputs(7224) <= not(inputs(125)) or (inputs(226));
    layer0_outputs(7225) <= not(inputs(207)) or (inputs(56));
    layer0_outputs(7226) <= inputs(151);
    layer0_outputs(7227) <= not(inputs(54)) or (inputs(129));
    layer0_outputs(7228) <= (inputs(27)) or (inputs(152));
    layer0_outputs(7229) <= (inputs(85)) xor (inputs(24));
    layer0_outputs(7230) <= inputs(169);
    layer0_outputs(7231) <= not((inputs(201)) or (inputs(170)));
    layer0_outputs(7232) <= (inputs(70)) xor (inputs(187));
    layer0_outputs(7233) <= not((inputs(210)) or (inputs(87)));
    layer0_outputs(7234) <= not(inputs(190));
    layer0_outputs(7235) <= not(inputs(239));
    layer0_outputs(7236) <= '0';
    layer0_outputs(7237) <= not(inputs(73));
    layer0_outputs(7238) <= not(inputs(140)) or (inputs(17));
    layer0_outputs(7239) <= not(inputs(128)) or (inputs(112));
    layer0_outputs(7240) <= (inputs(91)) xor (inputs(82));
    layer0_outputs(7241) <= not((inputs(36)) xor (inputs(247)));
    layer0_outputs(7242) <= not(inputs(52));
    layer0_outputs(7243) <= not((inputs(248)) or (inputs(72)));
    layer0_outputs(7244) <= not(inputs(51));
    layer0_outputs(7245) <= not(inputs(104));
    layer0_outputs(7246) <= not(inputs(121)) or (inputs(223));
    layer0_outputs(7247) <= (inputs(173)) or (inputs(23));
    layer0_outputs(7248) <= inputs(155);
    layer0_outputs(7249) <= not(inputs(167)) or (inputs(240));
    layer0_outputs(7250) <= inputs(139);
    layer0_outputs(7251) <= not((inputs(63)) or (inputs(172)));
    layer0_outputs(7252) <= inputs(163);
    layer0_outputs(7253) <= not((inputs(160)) xor (inputs(130)));
    layer0_outputs(7254) <= inputs(201);
    layer0_outputs(7255) <= inputs(244);
    layer0_outputs(7256) <= (inputs(102)) or (inputs(133));
    layer0_outputs(7257) <= (inputs(57)) and not (inputs(17));
    layer0_outputs(7258) <= not(inputs(92)) or (inputs(165));
    layer0_outputs(7259) <= not(inputs(57));
    layer0_outputs(7260) <= not(inputs(70)) or (inputs(25));
    layer0_outputs(7261) <= not(inputs(100));
    layer0_outputs(7262) <= (inputs(55)) and not (inputs(44));
    layer0_outputs(7263) <= (inputs(29)) and not (inputs(34));
    layer0_outputs(7264) <= not((inputs(68)) or (inputs(58)));
    layer0_outputs(7265) <= '0';
    layer0_outputs(7266) <= not((inputs(242)) or (inputs(139)));
    layer0_outputs(7267) <= (inputs(61)) xor (inputs(118));
    layer0_outputs(7268) <= (inputs(155)) and not (inputs(78));
    layer0_outputs(7269) <= (inputs(170)) xor (inputs(162));
    layer0_outputs(7270) <= not((inputs(70)) xor (inputs(151)));
    layer0_outputs(7271) <= not((inputs(191)) or (inputs(70)));
    layer0_outputs(7272) <= (inputs(106)) and (inputs(20));
    layer0_outputs(7273) <= '1';
    layer0_outputs(7274) <= not(inputs(202));
    layer0_outputs(7275) <= not((inputs(30)) xor (inputs(14)));
    layer0_outputs(7276) <= not(inputs(31));
    layer0_outputs(7277) <= (inputs(155)) and (inputs(220));
    layer0_outputs(7278) <= not(inputs(59)) or (inputs(18));
    layer0_outputs(7279) <= not((inputs(161)) xor (inputs(12)));
    layer0_outputs(7280) <= not(inputs(64));
    layer0_outputs(7281) <= (inputs(215)) or (inputs(228));
    layer0_outputs(7282) <= inputs(196);
    layer0_outputs(7283) <= not((inputs(23)) xor (inputs(65)));
    layer0_outputs(7284) <= (inputs(148)) and not (inputs(235));
    layer0_outputs(7285) <= '0';
    layer0_outputs(7286) <= (inputs(138)) and not (inputs(70));
    layer0_outputs(7287) <= not(inputs(234)) or (inputs(32));
    layer0_outputs(7288) <= inputs(85);
    layer0_outputs(7289) <= (inputs(144)) xor (inputs(76));
    layer0_outputs(7290) <= (inputs(43)) xor (inputs(53));
    layer0_outputs(7291) <= inputs(10);
    layer0_outputs(7292) <= '1';
    layer0_outputs(7293) <= not((inputs(187)) xor (inputs(58)));
    layer0_outputs(7294) <= not((inputs(161)) xor (inputs(132)));
    layer0_outputs(7295) <= not(inputs(46));
    layer0_outputs(7296) <= '0';
    layer0_outputs(7297) <= (inputs(185)) and (inputs(138));
    layer0_outputs(7298) <= not((inputs(254)) xor (inputs(136)));
    layer0_outputs(7299) <= (inputs(51)) and not (inputs(129));
    layer0_outputs(7300) <= (inputs(238)) or (inputs(51));
    layer0_outputs(7301) <= not((inputs(240)) or (inputs(147)));
    layer0_outputs(7302) <= not(inputs(253));
    layer0_outputs(7303) <= not((inputs(108)) xor (inputs(249)));
    layer0_outputs(7304) <= (inputs(83)) and not (inputs(209));
    layer0_outputs(7305) <= inputs(166);
    layer0_outputs(7306) <= (inputs(210)) xor (inputs(17));
    layer0_outputs(7307) <= not((inputs(190)) xor (inputs(247)));
    layer0_outputs(7308) <= (inputs(88)) and not (inputs(120));
    layer0_outputs(7309) <= not(inputs(156)) or (inputs(207));
    layer0_outputs(7310) <= not(inputs(92));
    layer0_outputs(7311) <= not(inputs(206)) or (inputs(144));
    layer0_outputs(7312) <= (inputs(52)) or (inputs(204));
    layer0_outputs(7313) <= (inputs(146)) xor (inputs(90));
    layer0_outputs(7314) <= not(inputs(151));
    layer0_outputs(7315) <= (inputs(145)) and not (inputs(224));
    layer0_outputs(7316) <= not((inputs(50)) and (inputs(11)));
    layer0_outputs(7317) <= (inputs(141)) or (inputs(92));
    layer0_outputs(7318) <= not(inputs(119)) or (inputs(44));
    layer0_outputs(7319) <= '1';
    layer0_outputs(7320) <= (inputs(41)) and not (inputs(62));
    layer0_outputs(7321) <= not((inputs(149)) or (inputs(150)));
    layer0_outputs(7322) <= not(inputs(164));
    layer0_outputs(7323) <= (inputs(6)) xor (inputs(208));
    layer0_outputs(7324) <= '1';
    layer0_outputs(7325) <= not(inputs(199));
    layer0_outputs(7326) <= inputs(244);
    layer0_outputs(7327) <= (inputs(32)) or (inputs(139));
    layer0_outputs(7328) <= (inputs(106)) xor (inputs(225));
    layer0_outputs(7329) <= not(inputs(242));
    layer0_outputs(7330) <= not(inputs(134));
    layer0_outputs(7331) <= (inputs(136)) and not (inputs(177));
    layer0_outputs(7332) <= not(inputs(194));
    layer0_outputs(7333) <= (inputs(106)) or (inputs(227));
    layer0_outputs(7334) <= not(inputs(132)) or (inputs(229));
    layer0_outputs(7335) <= inputs(63);
    layer0_outputs(7336) <= (inputs(5)) and (inputs(62));
    layer0_outputs(7337) <= inputs(222);
    layer0_outputs(7338) <= not(inputs(165)) or (inputs(28));
    layer0_outputs(7339) <= not(inputs(107)) or (inputs(23));
    layer0_outputs(7340) <= (inputs(20)) or (inputs(44));
    layer0_outputs(7341) <= (inputs(222)) or (inputs(232));
    layer0_outputs(7342) <= inputs(189);
    layer0_outputs(7343) <= '1';
    layer0_outputs(7344) <= (inputs(170)) and not (inputs(123));
    layer0_outputs(7345) <= not(inputs(85)) or (inputs(140));
    layer0_outputs(7346) <= not(inputs(74)) or (inputs(232));
    layer0_outputs(7347) <= (inputs(204)) and not (inputs(124));
    layer0_outputs(7348) <= inputs(117);
    layer0_outputs(7349) <= (inputs(9)) and not (inputs(190));
    layer0_outputs(7350) <= not((inputs(149)) xor (inputs(79)));
    layer0_outputs(7351) <= not((inputs(107)) xor (inputs(83)));
    layer0_outputs(7352) <= not(inputs(164));
    layer0_outputs(7353) <= (inputs(245)) xor (inputs(198));
    layer0_outputs(7354) <= not(inputs(33));
    layer0_outputs(7355) <= (inputs(134)) and not (inputs(221));
    layer0_outputs(7356) <= not((inputs(215)) or (inputs(223)));
    layer0_outputs(7357) <= '0';
    layer0_outputs(7358) <= not((inputs(157)) xor (inputs(182)));
    layer0_outputs(7359) <= (inputs(4)) or (inputs(249));
    layer0_outputs(7360) <= not(inputs(120));
    layer0_outputs(7361) <= not(inputs(197));
    layer0_outputs(7362) <= not(inputs(181)) or (inputs(78));
    layer0_outputs(7363) <= (inputs(249)) or (inputs(153));
    layer0_outputs(7364) <= not(inputs(147)) or (inputs(255));
    layer0_outputs(7365) <= (inputs(160)) or (inputs(156));
    layer0_outputs(7366) <= (inputs(213)) and (inputs(164));
    layer0_outputs(7367) <= not(inputs(77)) or (inputs(116));
    layer0_outputs(7368) <= not(inputs(218));
    layer0_outputs(7369) <= not(inputs(139));
    layer0_outputs(7370) <= not(inputs(118));
    layer0_outputs(7371) <= not(inputs(234));
    layer0_outputs(7372) <= not(inputs(138));
    layer0_outputs(7373) <= not((inputs(154)) xor (inputs(155)));
    layer0_outputs(7374) <= not(inputs(83)) or (inputs(128));
    layer0_outputs(7375) <= (inputs(51)) or (inputs(197));
    layer0_outputs(7376) <= inputs(76);
    layer0_outputs(7377) <= (inputs(90)) and not (inputs(239));
    layer0_outputs(7378) <= (inputs(253)) xor (inputs(36));
    layer0_outputs(7379) <= inputs(195);
    layer0_outputs(7380) <= not((inputs(130)) xor (inputs(131)));
    layer0_outputs(7381) <= inputs(131);
    layer0_outputs(7382) <= not((inputs(77)) or (inputs(18)));
    layer0_outputs(7383) <= not(inputs(215)) or (inputs(146));
    layer0_outputs(7384) <= (inputs(247)) xor (inputs(167));
    layer0_outputs(7385) <= not((inputs(89)) or (inputs(106)));
    layer0_outputs(7386) <= not(inputs(146));
    layer0_outputs(7387) <= (inputs(148)) and not (inputs(217));
    layer0_outputs(7388) <= (inputs(67)) or (inputs(108));
    layer0_outputs(7389) <= (inputs(83)) and not (inputs(34));
    layer0_outputs(7390) <= not((inputs(157)) or (inputs(165)));
    layer0_outputs(7391) <= not(inputs(84)) or (inputs(79));
    layer0_outputs(7392) <= inputs(117);
    layer0_outputs(7393) <= '0';
    layer0_outputs(7394) <= (inputs(164)) or (inputs(169));
    layer0_outputs(7395) <= (inputs(86)) and not (inputs(196));
    layer0_outputs(7396) <= (inputs(203)) and not (inputs(147));
    layer0_outputs(7397) <= not((inputs(34)) xor (inputs(116)));
    layer0_outputs(7398) <= inputs(59);
    layer0_outputs(7399) <= inputs(115);
    layer0_outputs(7400) <= (inputs(50)) and (inputs(177));
    layer0_outputs(7401) <= inputs(93);
    layer0_outputs(7402) <= (inputs(87)) and not (inputs(165));
    layer0_outputs(7403) <= not((inputs(197)) xor (inputs(112)));
    layer0_outputs(7404) <= not((inputs(226)) or (inputs(90)));
    layer0_outputs(7405) <= (inputs(98)) and not (inputs(243));
    layer0_outputs(7406) <= not(inputs(182));
    layer0_outputs(7407) <= not(inputs(134)) or (inputs(206));
    layer0_outputs(7408) <= not((inputs(144)) xor (inputs(35)));
    layer0_outputs(7409) <= not((inputs(204)) or (inputs(56)));
    layer0_outputs(7410) <= (inputs(39)) or (inputs(173));
    layer0_outputs(7411) <= not((inputs(116)) or (inputs(228)));
    layer0_outputs(7412) <= (inputs(1)) and (inputs(92));
    layer0_outputs(7413) <= not(inputs(137)) or (inputs(50));
    layer0_outputs(7414) <= (inputs(135)) and not (inputs(56));
    layer0_outputs(7415) <= (inputs(184)) and not (inputs(227));
    layer0_outputs(7416) <= (inputs(73)) and not (inputs(109));
    layer0_outputs(7417) <= (inputs(54)) or (inputs(195));
    layer0_outputs(7418) <= not(inputs(228));
    layer0_outputs(7419) <= (inputs(157)) or (inputs(181));
    layer0_outputs(7420) <= not((inputs(139)) xor (inputs(54)));
    layer0_outputs(7421) <= inputs(149);
    layer0_outputs(7422) <= inputs(125);
    layer0_outputs(7423) <= inputs(20);
    layer0_outputs(7424) <= inputs(183);
    layer0_outputs(7425) <= (inputs(3)) xor (inputs(211));
    layer0_outputs(7426) <= (inputs(175)) and not (inputs(245));
    layer0_outputs(7427) <= '0';
    layer0_outputs(7428) <= not((inputs(31)) and (inputs(237)));
    layer0_outputs(7429) <= not(inputs(70)) or (inputs(190));
    layer0_outputs(7430) <= (inputs(191)) or (inputs(153));
    layer0_outputs(7431) <= (inputs(52)) and not (inputs(207));
    layer0_outputs(7432) <= inputs(112);
    layer0_outputs(7433) <= (inputs(97)) and (inputs(244));
    layer0_outputs(7434) <= (inputs(224)) and not (inputs(28));
    layer0_outputs(7435) <= not(inputs(252)) or (inputs(219));
    layer0_outputs(7436) <= not(inputs(150));
    layer0_outputs(7437) <= not((inputs(165)) xor (inputs(195)));
    layer0_outputs(7438) <= (inputs(146)) and not (inputs(81));
    layer0_outputs(7439) <= '0';
    layer0_outputs(7440) <= (inputs(91)) or (inputs(212));
    layer0_outputs(7441) <= not(inputs(125));
    layer0_outputs(7442) <= not(inputs(181));
    layer0_outputs(7443) <= (inputs(58)) or (inputs(188));
    layer0_outputs(7444) <= not((inputs(63)) xor (inputs(64)));
    layer0_outputs(7445) <= not(inputs(216));
    layer0_outputs(7446) <= not((inputs(97)) or (inputs(152)));
    layer0_outputs(7447) <= (inputs(134)) or (inputs(12));
    layer0_outputs(7448) <= not(inputs(147)) or (inputs(143));
    layer0_outputs(7449) <= (inputs(254)) and not (inputs(193));
    layer0_outputs(7450) <= not(inputs(57)) or (inputs(227));
    layer0_outputs(7451) <= (inputs(9)) and not (inputs(226));
    layer0_outputs(7452) <= not(inputs(224));
    layer0_outputs(7453) <= (inputs(169)) or (inputs(45));
    layer0_outputs(7454) <= not((inputs(144)) xor (inputs(3)));
    layer0_outputs(7455) <= not(inputs(135));
    layer0_outputs(7456) <= not(inputs(220)) or (inputs(144));
    layer0_outputs(7457) <= (inputs(77)) and not (inputs(107));
    layer0_outputs(7458) <= not(inputs(171));
    layer0_outputs(7459) <= not(inputs(170)) or (inputs(14));
    layer0_outputs(7460) <= not(inputs(69));
    layer0_outputs(7461) <= not((inputs(168)) xor (inputs(28)));
    layer0_outputs(7462) <= '1';
    layer0_outputs(7463) <= (inputs(149)) or (inputs(199));
    layer0_outputs(7464) <= not((inputs(171)) and (inputs(137)));
    layer0_outputs(7465) <= (inputs(115)) and not (inputs(245));
    layer0_outputs(7466) <= (inputs(150)) xor (inputs(111));
    layer0_outputs(7467) <= (inputs(239)) xor (inputs(115));
    layer0_outputs(7468) <= (inputs(185)) or (inputs(72));
    layer0_outputs(7469) <= (inputs(104)) and not (inputs(241));
    layer0_outputs(7470) <= not(inputs(178));
    layer0_outputs(7471) <= not((inputs(128)) xor (inputs(33)));
    layer0_outputs(7472) <= not((inputs(163)) or (inputs(186)));
    layer0_outputs(7473) <= inputs(40);
    layer0_outputs(7474) <= not(inputs(102));
    layer0_outputs(7475) <= (inputs(203)) or (inputs(190));
    layer0_outputs(7476) <= not((inputs(7)) or (inputs(103)));
    layer0_outputs(7477) <= (inputs(63)) xor (inputs(18));
    layer0_outputs(7478) <= not((inputs(93)) xor (inputs(251)));
    layer0_outputs(7479) <= not(inputs(116));
    layer0_outputs(7480) <= not(inputs(124));
    layer0_outputs(7481) <= '1';
    layer0_outputs(7482) <= not(inputs(84)) or (inputs(223));
    layer0_outputs(7483) <= (inputs(42)) or (inputs(97));
    layer0_outputs(7484) <= not(inputs(138)) or (inputs(249));
    layer0_outputs(7485) <= not(inputs(251));
    layer0_outputs(7486) <= not((inputs(249)) or (inputs(131)));
    layer0_outputs(7487) <= not((inputs(223)) or (inputs(56)));
    layer0_outputs(7488) <= (inputs(181)) xor (inputs(177));
    layer0_outputs(7489) <= not((inputs(27)) xor (inputs(79)));
    layer0_outputs(7490) <= not((inputs(116)) or (inputs(151)));
    layer0_outputs(7491) <= not((inputs(38)) or (inputs(252)));
    layer0_outputs(7492) <= not((inputs(65)) or (inputs(237)));
    layer0_outputs(7493) <= (inputs(172)) or (inputs(182));
    layer0_outputs(7494) <= (inputs(226)) and not (inputs(49));
    layer0_outputs(7495) <= (inputs(188)) and not (inputs(237));
    layer0_outputs(7496) <= inputs(109);
    layer0_outputs(7497) <= not(inputs(77));
    layer0_outputs(7498) <= not(inputs(0));
    layer0_outputs(7499) <= not(inputs(67)) or (inputs(95));
    layer0_outputs(7500) <= not(inputs(70));
    layer0_outputs(7501) <= (inputs(63)) xor (inputs(212));
    layer0_outputs(7502) <= not(inputs(166)) or (inputs(33));
    layer0_outputs(7503) <= not((inputs(199)) or (inputs(179)));
    layer0_outputs(7504) <= not((inputs(120)) or (inputs(128)));
    layer0_outputs(7505) <= not((inputs(128)) or (inputs(99)));
    layer0_outputs(7506) <= not(inputs(149));
    layer0_outputs(7507) <= (inputs(229)) or (inputs(155));
    layer0_outputs(7508) <= not((inputs(83)) or (inputs(36)));
    layer0_outputs(7509) <= not((inputs(60)) or (inputs(159)));
    layer0_outputs(7510) <= not(inputs(251)) or (inputs(95));
    layer0_outputs(7511) <= not((inputs(97)) xor (inputs(149)));
    layer0_outputs(7512) <= '1';
    layer0_outputs(7513) <= (inputs(58)) xor (inputs(8));
    layer0_outputs(7514) <= not(inputs(66));
    layer0_outputs(7515) <= (inputs(1)) and (inputs(172));
    layer0_outputs(7516) <= (inputs(198)) and not (inputs(115));
    layer0_outputs(7517) <= not(inputs(30));
    layer0_outputs(7518) <= (inputs(100)) and not (inputs(95));
    layer0_outputs(7519) <= not(inputs(160)) or (inputs(32));
    layer0_outputs(7520) <= (inputs(198)) xor (inputs(192));
    layer0_outputs(7521) <= not((inputs(127)) xor (inputs(241)));
    layer0_outputs(7522) <= not(inputs(1)) or (inputs(31));
    layer0_outputs(7523) <= not(inputs(113));
    layer0_outputs(7524) <= not(inputs(104));
    layer0_outputs(7525) <= not((inputs(159)) xor (inputs(59)));
    layer0_outputs(7526) <= not((inputs(212)) or (inputs(3)));
    layer0_outputs(7527) <= (inputs(132)) and not (inputs(232));
    layer0_outputs(7528) <= (inputs(154)) xor (inputs(137));
    layer0_outputs(7529) <= not((inputs(109)) or (inputs(198)));
    layer0_outputs(7530) <= '0';
    layer0_outputs(7531) <= not(inputs(176)) or (inputs(193));
    layer0_outputs(7532) <= not(inputs(108)) or (inputs(22));
    layer0_outputs(7533) <= not((inputs(54)) or (inputs(154)));
    layer0_outputs(7534) <= not((inputs(93)) or (inputs(5)));
    layer0_outputs(7535) <= (inputs(236)) xor (inputs(38));
    layer0_outputs(7536) <= (inputs(99)) xor (inputs(34));
    layer0_outputs(7537) <= inputs(151);
    layer0_outputs(7538) <= '1';
    layer0_outputs(7539) <= '0';
    layer0_outputs(7540) <= (inputs(140)) or (inputs(148));
    layer0_outputs(7541) <= not((inputs(153)) or (inputs(220)));
    layer0_outputs(7542) <= not((inputs(80)) xor (inputs(40)));
    layer0_outputs(7543) <= inputs(212);
    layer0_outputs(7544) <= (inputs(93)) and not (inputs(251));
    layer0_outputs(7545) <= (inputs(27)) or (inputs(18));
    layer0_outputs(7546) <= '1';
    layer0_outputs(7547) <= not(inputs(237)) or (inputs(71));
    layer0_outputs(7548) <= not((inputs(21)) or (inputs(123)));
    layer0_outputs(7549) <= not((inputs(187)) xor (inputs(67)));
    layer0_outputs(7550) <= (inputs(253)) and (inputs(130));
    layer0_outputs(7551) <= (inputs(112)) xor (inputs(135));
    layer0_outputs(7552) <= (inputs(54)) xor (inputs(84));
    layer0_outputs(7553) <= not((inputs(1)) xor (inputs(219)));
    layer0_outputs(7554) <= not((inputs(23)) xor (inputs(151)));
    layer0_outputs(7555) <= (inputs(80)) or (inputs(93));
    layer0_outputs(7556) <= (inputs(86)) or (inputs(87));
    layer0_outputs(7557) <= not((inputs(166)) and (inputs(135)));
    layer0_outputs(7558) <= '0';
    layer0_outputs(7559) <= not(inputs(149)) or (inputs(217));
    layer0_outputs(7560) <= not(inputs(1)) or (inputs(130));
    layer0_outputs(7561) <= (inputs(120)) and not (inputs(93));
    layer0_outputs(7562) <= (inputs(16)) and (inputs(153));
    layer0_outputs(7563) <= not(inputs(238)) or (inputs(1));
    layer0_outputs(7564) <= not(inputs(116));
    layer0_outputs(7565) <= not((inputs(164)) or (inputs(13)));
    layer0_outputs(7566) <= not((inputs(143)) or (inputs(176)));
    layer0_outputs(7567) <= inputs(148);
    layer0_outputs(7568) <= inputs(40);
    layer0_outputs(7569) <= not((inputs(222)) or (inputs(171)));
    layer0_outputs(7570) <= (inputs(244)) and (inputs(4));
    layer0_outputs(7571) <= inputs(141);
    layer0_outputs(7572) <= not((inputs(183)) or (inputs(126)));
    layer0_outputs(7573) <= (inputs(87)) xor (inputs(6));
    layer0_outputs(7574) <= not(inputs(74)) or (inputs(232));
    layer0_outputs(7575) <= not(inputs(72));
    layer0_outputs(7576) <= (inputs(57)) and not (inputs(49));
    layer0_outputs(7577) <= inputs(171);
    layer0_outputs(7578) <= not((inputs(215)) xor (inputs(10)));
    layer0_outputs(7579) <= not((inputs(143)) xor (inputs(98)));
    layer0_outputs(7580) <= not(inputs(152));
    layer0_outputs(7581) <= not((inputs(94)) xor (inputs(23)));
    layer0_outputs(7582) <= not((inputs(228)) or (inputs(122)));
    layer0_outputs(7583) <= (inputs(194)) or (inputs(55));
    layer0_outputs(7584) <= not(inputs(167));
    layer0_outputs(7585) <= not(inputs(200)) or (inputs(133));
    layer0_outputs(7586) <= (inputs(200)) or (inputs(52));
    layer0_outputs(7587) <= inputs(118);
    layer0_outputs(7588) <= (inputs(181)) and not (inputs(230));
    layer0_outputs(7589) <= inputs(170);
    layer0_outputs(7590) <= (inputs(91)) or (inputs(175));
    layer0_outputs(7591) <= inputs(62);
    layer0_outputs(7592) <= (inputs(187)) or (inputs(209));
    layer0_outputs(7593) <= (inputs(104)) or (inputs(249));
    layer0_outputs(7594) <= not(inputs(92));
    layer0_outputs(7595) <= inputs(244);
    layer0_outputs(7596) <= (inputs(50)) and not (inputs(208));
    layer0_outputs(7597) <= inputs(187);
    layer0_outputs(7598) <= not((inputs(46)) and (inputs(222)));
    layer0_outputs(7599) <= inputs(111);
    layer0_outputs(7600) <= not(inputs(124));
    layer0_outputs(7601) <= not(inputs(118));
    layer0_outputs(7602) <= (inputs(180)) or (inputs(140));
    layer0_outputs(7603) <= inputs(89);
    layer0_outputs(7604) <= (inputs(49)) xor (inputs(17));
    layer0_outputs(7605) <= not((inputs(91)) or (inputs(47)));
    layer0_outputs(7606) <= (inputs(104)) and not (inputs(113));
    layer0_outputs(7607) <= not(inputs(90));
    layer0_outputs(7608) <= not(inputs(215)) or (inputs(243));
    layer0_outputs(7609) <= not(inputs(168));
    layer0_outputs(7610) <= inputs(34);
    layer0_outputs(7611) <= (inputs(196)) or (inputs(241));
    layer0_outputs(7612) <= not((inputs(214)) or (inputs(163)));
    layer0_outputs(7613) <= (inputs(173)) xor (inputs(137));
    layer0_outputs(7614) <= not(inputs(171));
    layer0_outputs(7615) <= not(inputs(153)) or (inputs(230));
    layer0_outputs(7616) <= not((inputs(232)) or (inputs(227)));
    layer0_outputs(7617) <= not((inputs(68)) or (inputs(10)));
    layer0_outputs(7618) <= not(inputs(90));
    layer0_outputs(7619) <= not(inputs(179)) or (inputs(129));
    layer0_outputs(7620) <= not((inputs(60)) xor (inputs(43)));
    layer0_outputs(7621) <= (inputs(78)) and (inputs(163));
    layer0_outputs(7622) <= not(inputs(247));
    layer0_outputs(7623) <= (inputs(22)) and (inputs(147));
    layer0_outputs(7624) <= inputs(176);
    layer0_outputs(7625) <= not(inputs(185));
    layer0_outputs(7626) <= (inputs(131)) or (inputs(131));
    layer0_outputs(7627) <= not((inputs(238)) or (inputs(92)));
    layer0_outputs(7628) <= (inputs(99)) xor (inputs(159));
    layer0_outputs(7629) <= (inputs(52)) or (inputs(184));
    layer0_outputs(7630) <= (inputs(133)) and not (inputs(8));
    layer0_outputs(7631) <= (inputs(65)) xor (inputs(233));
    layer0_outputs(7632) <= not((inputs(215)) or (inputs(114)));
    layer0_outputs(7633) <= (inputs(237)) and (inputs(64));
    layer0_outputs(7634) <= not(inputs(186)) or (inputs(138));
    layer0_outputs(7635) <= not(inputs(149));
    layer0_outputs(7636) <= (inputs(253)) xor (inputs(189));
    layer0_outputs(7637) <= not((inputs(157)) xor (inputs(209)));
    layer0_outputs(7638) <= not(inputs(77));
    layer0_outputs(7639) <= (inputs(87)) and not (inputs(179));
    layer0_outputs(7640) <= not(inputs(98)) or (inputs(209));
    layer0_outputs(7641) <= not((inputs(19)) or (inputs(104)));
    layer0_outputs(7642) <= not(inputs(152)) or (inputs(68));
    layer0_outputs(7643) <= not((inputs(209)) xor (inputs(244)));
    layer0_outputs(7644) <= (inputs(150)) or (inputs(132));
    layer0_outputs(7645) <= not(inputs(71)) or (inputs(219));
    layer0_outputs(7646) <= not(inputs(148)) or (inputs(39));
    layer0_outputs(7647) <= not(inputs(114));
    layer0_outputs(7648) <= (inputs(207)) or (inputs(108));
    layer0_outputs(7649) <= inputs(171);
    layer0_outputs(7650) <= not((inputs(191)) xor (inputs(6)));
    layer0_outputs(7651) <= not((inputs(42)) xor (inputs(44)));
    layer0_outputs(7652) <= inputs(124);
    layer0_outputs(7653) <= not(inputs(221)) or (inputs(49));
    layer0_outputs(7654) <= inputs(175);
    layer0_outputs(7655) <= not(inputs(206));
    layer0_outputs(7656) <= (inputs(89)) or (inputs(246));
    layer0_outputs(7657) <= not(inputs(137)) or (inputs(26));
    layer0_outputs(7658) <= not(inputs(62)) or (inputs(247));
    layer0_outputs(7659) <= not((inputs(85)) xor (inputs(47)));
    layer0_outputs(7660) <= not(inputs(149)) or (inputs(54));
    layer0_outputs(7661) <= (inputs(99)) or (inputs(145));
    layer0_outputs(7662) <= inputs(149);
    layer0_outputs(7663) <= not(inputs(153)) or (inputs(26));
    layer0_outputs(7664) <= (inputs(222)) or (inputs(189));
    layer0_outputs(7665) <= (inputs(191)) and (inputs(0));
    layer0_outputs(7666) <= (inputs(151)) and not (inputs(165));
    layer0_outputs(7667) <= not((inputs(1)) or (inputs(219)));
    layer0_outputs(7668) <= not((inputs(152)) or (inputs(80)));
    layer0_outputs(7669) <= '1';
    layer0_outputs(7670) <= (inputs(182)) or (inputs(111));
    layer0_outputs(7671) <= not(inputs(42));
    layer0_outputs(7672) <= not((inputs(182)) xor (inputs(254)));
    layer0_outputs(7673) <= inputs(215);
    layer0_outputs(7674) <= not((inputs(34)) and (inputs(224)));
    layer0_outputs(7675) <= '1';
    layer0_outputs(7676) <= not((inputs(16)) xor (inputs(98)));
    layer0_outputs(7677) <= (inputs(3)) and (inputs(76));
    layer0_outputs(7678) <= (inputs(212)) and (inputs(10));
    layer0_outputs(7679) <= not(inputs(248)) or (inputs(161));
    outputs(0) <= layer0_outputs(2113);
    outputs(1) <= not(layer0_outputs(4283));
    outputs(2) <= (layer0_outputs(743)) or (layer0_outputs(4779));
    outputs(3) <= (layer0_outputs(6878)) and not (layer0_outputs(6299));
    outputs(4) <= not(layer0_outputs(5229));
    outputs(5) <= layer0_outputs(348);
    outputs(6) <= not((layer0_outputs(7071)) or (layer0_outputs(5607)));
    outputs(7) <= not(layer0_outputs(4259));
    outputs(8) <= (layer0_outputs(2880)) and not (layer0_outputs(5366));
    outputs(9) <= not(layer0_outputs(4482));
    outputs(10) <= not((layer0_outputs(442)) or (layer0_outputs(5353)));
    outputs(11) <= (layer0_outputs(679)) xor (layer0_outputs(7478));
    outputs(12) <= layer0_outputs(2979);
    outputs(13) <= layer0_outputs(6600);
    outputs(14) <= not(layer0_outputs(7532));
    outputs(15) <= (layer0_outputs(2706)) and not (layer0_outputs(3062));
    outputs(16) <= (layer0_outputs(5914)) and (layer0_outputs(7496));
    outputs(17) <= layer0_outputs(4123);
    outputs(18) <= layer0_outputs(6217);
    outputs(19) <= not(layer0_outputs(3846));
    outputs(20) <= layer0_outputs(1410);
    outputs(21) <= (layer0_outputs(512)) xor (layer0_outputs(665));
    outputs(22) <= (layer0_outputs(3244)) and (layer0_outputs(3349));
    outputs(23) <= not(layer0_outputs(618));
    outputs(24) <= '1';
    outputs(25) <= (layer0_outputs(876)) and (layer0_outputs(386));
    outputs(26) <= not((layer0_outputs(2291)) or (layer0_outputs(2985)));
    outputs(27) <= (layer0_outputs(7453)) xor (layer0_outputs(3823));
    outputs(28) <= (layer0_outputs(6370)) xor (layer0_outputs(5400));
    outputs(29) <= (layer0_outputs(7241)) and not (layer0_outputs(2399));
    outputs(30) <= not((layer0_outputs(5294)) xor (layer0_outputs(2279)));
    outputs(31) <= not(layer0_outputs(2739));
    outputs(32) <= layer0_outputs(7166);
    outputs(33) <= layer0_outputs(4808);
    outputs(34) <= not((layer0_outputs(3418)) xor (layer0_outputs(2387)));
    outputs(35) <= layer0_outputs(3647);
    outputs(36) <= (layer0_outputs(1860)) and (layer0_outputs(2755));
    outputs(37) <= not(layer0_outputs(1583)) or (layer0_outputs(3748));
    outputs(38) <= not((layer0_outputs(5957)) xor (layer0_outputs(1108)));
    outputs(39) <= not(layer0_outputs(5685));
    outputs(40) <= layer0_outputs(6577);
    outputs(41) <= not(layer0_outputs(3385)) or (layer0_outputs(2384));
    outputs(42) <= (layer0_outputs(3034)) xor (layer0_outputs(1095));
    outputs(43) <= layer0_outputs(4124);
    outputs(44) <= not(layer0_outputs(1897));
    outputs(45) <= not(layer0_outputs(6970));
    outputs(46) <= layer0_outputs(3631);
    outputs(47) <= layer0_outputs(4363);
    outputs(48) <= layer0_outputs(1091);
    outputs(49) <= not(layer0_outputs(1274));
    outputs(50) <= layer0_outputs(212);
    outputs(51) <= not(layer0_outputs(696));
    outputs(52) <= layer0_outputs(6867);
    outputs(53) <= not((layer0_outputs(691)) and (layer0_outputs(1530)));
    outputs(54) <= not(layer0_outputs(1778));
    outputs(55) <= not(layer0_outputs(3791));
    outputs(56) <= not((layer0_outputs(1077)) xor (layer0_outputs(1963)));
    outputs(57) <= not(layer0_outputs(6732)) or (layer0_outputs(6790));
    outputs(58) <= not((layer0_outputs(4317)) and (layer0_outputs(96)));
    outputs(59) <= not((layer0_outputs(2046)) xor (layer0_outputs(6060)));
    outputs(60) <= (layer0_outputs(3438)) xor (layer0_outputs(5440));
    outputs(61) <= not((layer0_outputs(3504)) and (layer0_outputs(6260)));
    outputs(62) <= not(layer0_outputs(7532));
    outputs(63) <= not((layer0_outputs(7672)) and (layer0_outputs(5415)));
    outputs(64) <= not(layer0_outputs(5432));
    outputs(65) <= not((layer0_outputs(3353)) and (layer0_outputs(3364)));
    outputs(66) <= not((layer0_outputs(5873)) xor (layer0_outputs(6619)));
    outputs(67) <= not((layer0_outputs(6320)) xor (layer0_outputs(7566)));
    outputs(68) <= not(layer0_outputs(4766)) or (layer0_outputs(1615));
    outputs(69) <= not(layer0_outputs(7341));
    outputs(70) <= (layer0_outputs(5978)) or (layer0_outputs(2409));
    outputs(71) <= layer0_outputs(4446);
    outputs(72) <= layer0_outputs(5968);
    outputs(73) <= layer0_outputs(1906);
    outputs(74) <= (layer0_outputs(3766)) or (layer0_outputs(1281));
    outputs(75) <= not((layer0_outputs(1048)) or (layer0_outputs(2129)));
    outputs(76) <= not((layer0_outputs(5601)) xor (layer0_outputs(7152)));
    outputs(77) <= layer0_outputs(5168);
    outputs(78) <= not(layer0_outputs(2226)) or (layer0_outputs(1090));
    outputs(79) <= layer0_outputs(3568);
    outputs(80) <= not((layer0_outputs(3751)) or (layer0_outputs(2078)));
    outputs(81) <= not((layer0_outputs(6224)) and (layer0_outputs(602)));
    outputs(82) <= not((layer0_outputs(1862)) and (layer0_outputs(6111)));
    outputs(83) <= layer0_outputs(2952);
    outputs(84) <= layer0_outputs(6286);
    outputs(85) <= not(layer0_outputs(5493)) or (layer0_outputs(3904));
    outputs(86) <= (layer0_outputs(7098)) and not (layer0_outputs(6123));
    outputs(87) <= (layer0_outputs(6712)) xor (layer0_outputs(3356));
    outputs(88) <= (layer0_outputs(7508)) and not (layer0_outputs(4773));
    outputs(89) <= not(layer0_outputs(6997));
    outputs(90) <= layer0_outputs(5289);
    outputs(91) <= not(layer0_outputs(7450)) or (layer0_outputs(6193));
    outputs(92) <= not((layer0_outputs(4312)) xor (layer0_outputs(906)));
    outputs(93) <= not(layer0_outputs(7600));
    outputs(94) <= layer0_outputs(1453);
    outputs(95) <= layer0_outputs(3333);
    outputs(96) <= not(layer0_outputs(1755));
    outputs(97) <= not((layer0_outputs(5486)) xor (layer0_outputs(3241)));
    outputs(98) <= (layer0_outputs(4572)) and (layer0_outputs(7073));
    outputs(99) <= '0';
    outputs(100) <= not(layer0_outputs(6718)) or (layer0_outputs(725));
    outputs(101) <= (layer0_outputs(1176)) xor (layer0_outputs(2286));
    outputs(102) <= not(layer0_outputs(3132));
    outputs(103) <= not(layer0_outputs(5916));
    outputs(104) <= not((layer0_outputs(4360)) xor (layer0_outputs(4664)));
    outputs(105) <= (layer0_outputs(3857)) and not (layer0_outputs(5261));
    outputs(106) <= (layer0_outputs(37)) xor (layer0_outputs(2108));
    outputs(107) <= not(layer0_outputs(2995)) or (layer0_outputs(4300));
    outputs(108) <= not(layer0_outputs(3380));
    outputs(109) <= '1';
    outputs(110) <= layer0_outputs(3717);
    outputs(111) <= (layer0_outputs(3271)) and not (layer0_outputs(2544));
    outputs(112) <= layer0_outputs(5588);
    outputs(113) <= not(layer0_outputs(304));
    outputs(114) <= (layer0_outputs(7018)) xor (layer0_outputs(2561));
    outputs(115) <= layer0_outputs(4989);
    outputs(116) <= not(layer0_outputs(4464)) or (layer0_outputs(4704));
    outputs(117) <= not((layer0_outputs(1361)) or (layer0_outputs(7179)));
    outputs(118) <= (layer0_outputs(6029)) or (layer0_outputs(5420));
    outputs(119) <= (layer0_outputs(3654)) and (layer0_outputs(3268));
    outputs(120) <= not((layer0_outputs(2137)) xor (layer0_outputs(2115)));
    outputs(121) <= layer0_outputs(944);
    outputs(122) <= (layer0_outputs(6977)) xor (layer0_outputs(4333));
    outputs(123) <= (layer0_outputs(25)) or (layer0_outputs(1014));
    outputs(124) <= not(layer0_outputs(4001));
    outputs(125) <= (layer0_outputs(6129)) xor (layer0_outputs(5277));
    outputs(126) <= layer0_outputs(4473);
    outputs(127) <= (layer0_outputs(774)) xor (layer0_outputs(3874));
    outputs(128) <= layer0_outputs(6455);
    outputs(129) <= not(layer0_outputs(5149));
    outputs(130) <= (layer0_outputs(4640)) and not (layer0_outputs(7000));
    outputs(131) <= not((layer0_outputs(4749)) and (layer0_outputs(4796)));
    outputs(132) <= (layer0_outputs(6480)) and not (layer0_outputs(277));
    outputs(133) <= not(layer0_outputs(3184)) or (layer0_outputs(3475));
    outputs(134) <= not(layer0_outputs(1435));
    outputs(135) <= not(layer0_outputs(1192));
    outputs(136) <= not((layer0_outputs(1243)) xor (layer0_outputs(1634)));
    outputs(137) <= (layer0_outputs(1203)) and (layer0_outputs(1312));
    outputs(138) <= not(layer0_outputs(6253));
    outputs(139) <= not(layer0_outputs(1539));
    outputs(140) <= not(layer0_outputs(7442));
    outputs(141) <= (layer0_outputs(1859)) xor (layer0_outputs(6098));
    outputs(142) <= (layer0_outputs(7249)) and not (layer0_outputs(353));
    outputs(143) <= (layer0_outputs(3488)) or (layer0_outputs(7006));
    outputs(144) <= layer0_outputs(4811);
    outputs(145) <= (layer0_outputs(6610)) xor (layer0_outputs(7404));
    outputs(146) <= layer0_outputs(3589);
    outputs(147) <= not(layer0_outputs(246));
    outputs(148) <= layer0_outputs(2076);
    outputs(149) <= not(layer0_outputs(7259));
    outputs(150) <= not(layer0_outputs(5539));
    outputs(151) <= layer0_outputs(4291);
    outputs(152) <= not((layer0_outputs(5324)) xor (layer0_outputs(1356)));
    outputs(153) <= not(layer0_outputs(2086)) or (layer0_outputs(3218));
    outputs(154) <= (layer0_outputs(6081)) and not (layer0_outputs(4437));
    outputs(155) <= not(layer0_outputs(121));
    outputs(156) <= not(layer0_outputs(5533));
    outputs(157) <= (layer0_outputs(3159)) xor (layer0_outputs(3138));
    outputs(158) <= not(layer0_outputs(480)) or (layer0_outputs(1568));
    outputs(159) <= not(layer0_outputs(3716));
    outputs(160) <= not(layer0_outputs(7303));
    outputs(161) <= layer0_outputs(485);
    outputs(162) <= (layer0_outputs(3729)) and (layer0_outputs(2687));
    outputs(163) <= layer0_outputs(1742);
    outputs(164) <= not(layer0_outputs(6039)) or (layer0_outputs(2083));
    outputs(165) <= not(layer0_outputs(1260));
    outputs(166) <= layer0_outputs(2190);
    outputs(167) <= not(layer0_outputs(7466));
    outputs(168) <= (layer0_outputs(411)) and not (layer0_outputs(6671));
    outputs(169) <= (layer0_outputs(1984)) and (layer0_outputs(3375));
    outputs(170) <= not(layer0_outputs(1078)) or (layer0_outputs(1158));
    outputs(171) <= not(layer0_outputs(3097));
    outputs(172) <= not((layer0_outputs(4564)) xor (layer0_outputs(676)));
    outputs(173) <= layer0_outputs(937);
    outputs(174) <= not(layer0_outputs(7142));
    outputs(175) <= (layer0_outputs(472)) xor (layer0_outputs(2482));
    outputs(176) <= not((layer0_outputs(2373)) or (layer0_outputs(6850)));
    outputs(177) <= layer0_outputs(5843);
    outputs(178) <= not(layer0_outputs(5076));
    outputs(179) <= not(layer0_outputs(6745));
    outputs(180) <= not(layer0_outputs(3086));
    outputs(181) <= layer0_outputs(624);
    outputs(182) <= (layer0_outputs(4238)) xor (layer0_outputs(6119));
    outputs(183) <= not(layer0_outputs(6570));
    outputs(184) <= not(layer0_outputs(4897));
    outputs(185) <= not((layer0_outputs(3533)) xor (layer0_outputs(4637)));
    outputs(186) <= not(layer0_outputs(3659));
    outputs(187) <= layer0_outputs(1278);
    outputs(188) <= (layer0_outputs(4925)) xor (layer0_outputs(2541));
    outputs(189) <= not(layer0_outputs(404));
    outputs(190) <= not(layer0_outputs(491));
    outputs(191) <= not((layer0_outputs(6943)) xor (layer0_outputs(3315)));
    outputs(192) <= (layer0_outputs(4949)) xor (layer0_outputs(4202));
    outputs(193) <= not(layer0_outputs(6877)) or (layer0_outputs(5889));
    outputs(194) <= layer0_outputs(857);
    outputs(195) <= layer0_outputs(7662);
    outputs(196) <= not((layer0_outputs(3838)) xor (layer0_outputs(2662)));
    outputs(197) <= not(layer0_outputs(3639)) or (layer0_outputs(2967));
    outputs(198) <= layer0_outputs(153);
    outputs(199) <= not(layer0_outputs(5729)) or (layer0_outputs(7130));
    outputs(200) <= not(layer0_outputs(7040));
    outputs(201) <= not(layer0_outputs(1387));
    outputs(202) <= (layer0_outputs(4499)) xor (layer0_outputs(5639));
    outputs(203) <= (layer0_outputs(3705)) xor (layer0_outputs(1851));
    outputs(204) <= layer0_outputs(1825);
    outputs(205) <= layer0_outputs(866);
    outputs(206) <= layer0_outputs(5351);
    outputs(207) <= layer0_outputs(3691);
    outputs(208) <= not(layer0_outputs(7551));
    outputs(209) <= (layer0_outputs(3155)) and not (layer0_outputs(4139));
    outputs(210) <= (layer0_outputs(5041)) xor (layer0_outputs(3415));
    outputs(211) <= not(layer0_outputs(1749));
    outputs(212) <= not((layer0_outputs(5178)) xor (layer0_outputs(6189)));
    outputs(213) <= not(layer0_outputs(3624)) or (layer0_outputs(1223));
    outputs(214) <= layer0_outputs(7123);
    outputs(215) <= not(layer0_outputs(4901)) or (layer0_outputs(7209));
    outputs(216) <= layer0_outputs(4462);
    outputs(217) <= layer0_outputs(2615);
    outputs(218) <= (layer0_outputs(692)) xor (layer0_outputs(2310));
    outputs(219) <= not(layer0_outputs(4183));
    outputs(220) <= not((layer0_outputs(1840)) xor (layer0_outputs(7268)));
    outputs(221) <= layer0_outputs(1067);
    outputs(222) <= layer0_outputs(7140);
    outputs(223) <= layer0_outputs(6868);
    outputs(224) <= (layer0_outputs(4830)) xor (layer0_outputs(1770));
    outputs(225) <= (layer0_outputs(7049)) xor (layer0_outputs(4577));
    outputs(226) <= layer0_outputs(4611);
    outputs(227) <= layer0_outputs(5692);
    outputs(228) <= (layer0_outputs(1881)) xor (layer0_outputs(2669));
    outputs(229) <= not(layer0_outputs(6587));
    outputs(230) <= not(layer0_outputs(2807));
    outputs(231) <= not(layer0_outputs(1527));
    outputs(232) <= not(layer0_outputs(2900));
    outputs(233) <= not(layer0_outputs(6494));
    outputs(234) <= not(layer0_outputs(7380));
    outputs(235) <= layer0_outputs(7611);
    outputs(236) <= not(layer0_outputs(1331));
    outputs(237) <= not(layer0_outputs(4892)) or (layer0_outputs(6281));
    outputs(238) <= not(layer0_outputs(6717));
    outputs(239) <= not((layer0_outputs(5192)) xor (layer0_outputs(6682)));
    outputs(240) <= (layer0_outputs(206)) and not (layer0_outputs(5547));
    outputs(241) <= layer0_outputs(3934);
    outputs(242) <= not(layer0_outputs(7301));
    outputs(243) <= not(layer0_outputs(2950));
    outputs(244) <= not((layer0_outputs(4939)) or (layer0_outputs(5090)));
    outputs(245) <= not((layer0_outputs(3949)) xor (layer0_outputs(5254)));
    outputs(246) <= not(layer0_outputs(6225));
    outputs(247) <= not(layer0_outputs(5751));
    outputs(248) <= (layer0_outputs(6506)) or (layer0_outputs(4129));
    outputs(249) <= not((layer0_outputs(589)) xor (layer0_outputs(3517)));
    outputs(250) <= layer0_outputs(1605);
    outputs(251) <= not((layer0_outputs(7446)) xor (layer0_outputs(4226)));
    outputs(252) <= (layer0_outputs(7330)) and (layer0_outputs(7079));
    outputs(253) <= not(layer0_outputs(4463));
    outputs(254) <= layer0_outputs(4427);
    outputs(255) <= not((layer0_outputs(7221)) and (layer0_outputs(2367)));
    outputs(256) <= layer0_outputs(993);
    outputs(257) <= layer0_outputs(1941);
    outputs(258) <= not(layer0_outputs(2613));
    outputs(259) <= (layer0_outputs(3671)) xor (layer0_outputs(5296));
    outputs(260) <= (layer0_outputs(6128)) or (layer0_outputs(804));
    outputs(261) <= (layer0_outputs(6921)) xor (layer0_outputs(6008));
    outputs(262) <= not(layer0_outputs(4971));
    outputs(263) <= not(layer0_outputs(5949));
    outputs(264) <= not((layer0_outputs(6401)) and (layer0_outputs(3567)));
    outputs(265) <= layer0_outputs(5484);
    outputs(266) <= not(layer0_outputs(7390));
    outputs(267) <= layer0_outputs(5667);
    outputs(268) <= layer0_outputs(3366);
    outputs(269) <= layer0_outputs(1375);
    outputs(270) <= not(layer0_outputs(735)) or (layer0_outputs(7252));
    outputs(271) <= layer0_outputs(2921);
    outputs(272) <= (layer0_outputs(997)) or (layer0_outputs(4375));
    outputs(273) <= not((layer0_outputs(1734)) xor (layer0_outputs(7074)));
    outputs(274) <= '0';
    outputs(275) <= not(layer0_outputs(1147)) or (layer0_outputs(5328));
    outputs(276) <= not(layer0_outputs(1877));
    outputs(277) <= not((layer0_outputs(2686)) xor (layer0_outputs(2063)));
    outputs(278) <= (layer0_outputs(5597)) xor (layer0_outputs(5691));
    outputs(279) <= not((layer0_outputs(3626)) or (layer0_outputs(2417)));
    outputs(280) <= (layer0_outputs(861)) and not (layer0_outputs(7024));
    outputs(281) <= (layer0_outputs(1088)) xor (layer0_outputs(2271));
    outputs(282) <= (layer0_outputs(5801)) and not (layer0_outputs(1671));
    outputs(283) <= layer0_outputs(2761);
    outputs(284) <= not((layer0_outputs(2079)) xor (layer0_outputs(4563)));
    outputs(285) <= (layer0_outputs(5272)) xor (layer0_outputs(1248));
    outputs(286) <= not(layer0_outputs(3016)) or (layer0_outputs(5936));
    outputs(287) <= (layer0_outputs(1456)) xor (layer0_outputs(7078));
    outputs(288) <= not((layer0_outputs(1146)) xor (layer0_outputs(7353)));
    outputs(289) <= layer0_outputs(2546);
    outputs(290) <= not(layer0_outputs(1042));
    outputs(291) <= not(layer0_outputs(7070)) or (layer0_outputs(6951));
    outputs(292) <= layer0_outputs(5235);
    outputs(293) <= (layer0_outputs(2942)) or (layer0_outputs(2017));
    outputs(294) <= layer0_outputs(1391);
    outputs(295) <= not((layer0_outputs(1136)) or (layer0_outputs(5312)));
    outputs(296) <= layer0_outputs(1959);
    outputs(297) <= (layer0_outputs(3107)) and not (layer0_outputs(6495));
    outputs(298) <= not((layer0_outputs(5986)) and (layer0_outputs(2981)));
    outputs(299) <= not(layer0_outputs(4538)) or (layer0_outputs(3249));
    outputs(300) <= not(layer0_outputs(2701));
    outputs(301) <= (layer0_outputs(4874)) xor (layer0_outputs(6993));
    outputs(302) <= not(layer0_outputs(4761));
    outputs(303) <= not(layer0_outputs(352));
    outputs(304) <= not((layer0_outputs(6178)) and (layer0_outputs(2897)));
    outputs(305) <= not((layer0_outputs(1666)) or (layer0_outputs(61)));
    outputs(306) <= (layer0_outputs(4603)) or (layer0_outputs(2916));
    outputs(307) <= layer0_outputs(2628);
    outputs(308) <= not(layer0_outputs(7674)) or (layer0_outputs(3666));
    outputs(309) <= (layer0_outputs(2649)) xor (layer0_outputs(7368));
    outputs(310) <= not(layer0_outputs(1217));
    outputs(311) <= not((layer0_outputs(5496)) xor (layer0_outputs(992)));
    outputs(312) <= not((layer0_outputs(7050)) xor (layer0_outputs(2003)));
    outputs(313) <= not((layer0_outputs(7455)) xor (layer0_outputs(3711)));
    outputs(314) <= not(layer0_outputs(5533));
    outputs(315) <= (layer0_outputs(3047)) or (layer0_outputs(3743));
    outputs(316) <= not(layer0_outputs(7437));
    outputs(317) <= not((layer0_outputs(676)) xor (layer0_outputs(4792)));
    outputs(318) <= not(layer0_outputs(5891));
    outputs(319) <= layer0_outputs(718);
    outputs(320) <= not((layer0_outputs(608)) or (layer0_outputs(7535)));
    outputs(321) <= not(layer0_outputs(1495)) or (layer0_outputs(3347));
    outputs(322) <= layer0_outputs(4293);
    outputs(323) <= not((layer0_outputs(5885)) and (layer0_outputs(4268)));
    outputs(324) <= not((layer0_outputs(135)) xor (layer0_outputs(1798)));
    outputs(325) <= layer0_outputs(1812);
    outputs(326) <= (layer0_outputs(7399)) or (layer0_outputs(592));
    outputs(327) <= (layer0_outputs(4060)) or (layer0_outputs(3646));
    outputs(328) <= layer0_outputs(1379);
    outputs(329) <= not((layer0_outputs(5271)) xor (layer0_outputs(1248)));
    outputs(330) <= not((layer0_outputs(5887)) or (layer0_outputs(3890)));
    outputs(331) <= layer0_outputs(4946);
    outputs(332) <= not((layer0_outputs(6507)) xor (layer0_outputs(1888)));
    outputs(333) <= layer0_outputs(5067);
    outputs(334) <= (layer0_outputs(3824)) xor (layer0_outputs(2639));
    outputs(335) <= not(layer0_outputs(3742)) or (layer0_outputs(4088));
    outputs(336) <= layer0_outputs(6988);
    outputs(337) <= (layer0_outputs(7238)) xor (layer0_outputs(6883));
    outputs(338) <= not((layer0_outputs(5354)) xor (layer0_outputs(7520)));
    outputs(339) <= (layer0_outputs(5580)) and not (layer0_outputs(235));
    outputs(340) <= not(layer0_outputs(1288));
    outputs(341) <= layer0_outputs(263);
    outputs(342) <= not((layer0_outputs(1960)) xor (layer0_outputs(2509)));
    outputs(343) <= not(layer0_outputs(3163));
    outputs(344) <= (layer0_outputs(6630)) xor (layer0_outputs(3783));
    outputs(345) <= not(layer0_outputs(77));
    outputs(346) <= (layer0_outputs(1329)) xor (layer0_outputs(7320));
    outputs(347) <= not(layer0_outputs(3205)) or (layer0_outputs(7271));
    outputs(348) <= (layer0_outputs(4081)) xor (layer0_outputs(2974));
    outputs(349) <= not(layer0_outputs(3455));
    outputs(350) <= layer0_outputs(503);
    outputs(351) <= not(layer0_outputs(1705));
    outputs(352) <= layer0_outputs(2025);
    outputs(353) <= not(layer0_outputs(1589));
    outputs(354) <= (layer0_outputs(3975)) xor (layer0_outputs(4736));
    outputs(355) <= layer0_outputs(6328);
    outputs(356) <= not(layer0_outputs(1215));
    outputs(357) <= (layer0_outputs(1753)) xor (layer0_outputs(2007));
    outputs(358) <= (layer0_outputs(5448)) and (layer0_outputs(3605));
    outputs(359) <= layer0_outputs(7269);
    outputs(360) <= layer0_outputs(5876);
    outputs(361) <= not(layer0_outputs(6728)) or (layer0_outputs(1035));
    outputs(362) <= '1';
    outputs(363) <= layer0_outputs(52);
    outputs(364) <= not(layer0_outputs(2928));
    outputs(365) <= not(layer0_outputs(1712));
    outputs(366) <= layer0_outputs(7556);
    outputs(367) <= (layer0_outputs(4565)) xor (layer0_outputs(4747));
    outputs(368) <= layer0_outputs(6282);
    outputs(369) <= not(layer0_outputs(298)) or (layer0_outputs(968));
    outputs(370) <= not(layer0_outputs(1591));
    outputs(371) <= layer0_outputs(789);
    outputs(372) <= layer0_outputs(758);
    outputs(373) <= layer0_outputs(4244);
    outputs(374) <= (layer0_outputs(2881)) xor (layer0_outputs(418));
    outputs(375) <= layer0_outputs(3994);
    outputs(376) <= (layer0_outputs(2718)) and not (layer0_outputs(5892));
    outputs(377) <= layer0_outputs(1545);
    outputs(378) <= layer0_outputs(5072);
    outputs(379) <= layer0_outputs(7240);
    outputs(380) <= not(layer0_outputs(5068));
    outputs(381) <= layer0_outputs(7421);
    outputs(382) <= not(layer0_outputs(359));
    outputs(383) <= layer0_outputs(3883);
    outputs(384) <= layer0_outputs(6099);
    outputs(385) <= not(layer0_outputs(7637));
    outputs(386) <= not((layer0_outputs(2289)) and (layer0_outputs(4172)));
    outputs(387) <= layer0_outputs(1417);
    outputs(388) <= not(layer0_outputs(4960));
    outputs(389) <= layer0_outputs(701);
    outputs(390) <= not(layer0_outputs(6313)) or (layer0_outputs(6211));
    outputs(391) <= not((layer0_outputs(5097)) xor (layer0_outputs(1950)));
    outputs(392) <= layer0_outputs(2929);
    outputs(393) <= layer0_outputs(370);
    outputs(394) <= (layer0_outputs(4666)) and not (layer0_outputs(2171));
    outputs(395) <= (layer0_outputs(2589)) xor (layer0_outputs(4327));
    outputs(396) <= not((layer0_outputs(3069)) and (layer0_outputs(4758)));
    outputs(397) <= (layer0_outputs(6321)) or (layer0_outputs(91));
    outputs(398) <= not(layer0_outputs(1912));
    outputs(399) <= layer0_outputs(6286);
    outputs(400) <= (layer0_outputs(4449)) and not (layer0_outputs(2689));
    outputs(401) <= (layer0_outputs(7525)) xor (layer0_outputs(4270));
    outputs(402) <= not(layer0_outputs(6495));
    outputs(403) <= not(layer0_outputs(2385));
    outputs(404) <= (layer0_outputs(2075)) xor (layer0_outputs(5791));
    outputs(405) <= layer0_outputs(3343);
    outputs(406) <= not((layer0_outputs(770)) xor (layer0_outputs(3623)));
    outputs(407) <= not((layer0_outputs(6677)) xor (layer0_outputs(3902)));
    outputs(408) <= layer0_outputs(6209);
    outputs(409) <= not(layer0_outputs(4438)) or (layer0_outputs(3760));
    outputs(410) <= (layer0_outputs(5459)) or (layer0_outputs(3859));
    outputs(411) <= (layer0_outputs(2787)) and not (layer0_outputs(6753));
    outputs(412) <= (layer0_outputs(1223)) or (layer0_outputs(278));
    outputs(413) <= not(layer0_outputs(3644));
    outputs(414) <= (layer0_outputs(7081)) and not (layer0_outputs(6194));
    outputs(415) <= layer0_outputs(1398);
    outputs(416) <= not((layer0_outputs(7494)) and (layer0_outputs(5444)));
    outputs(417) <= not(layer0_outputs(3512));
    outputs(418) <= layer0_outputs(4887);
    outputs(419) <= layer0_outputs(7360);
    outputs(420) <= not(layer0_outputs(1598));
    outputs(421) <= (layer0_outputs(4985)) and not (layer0_outputs(129));
    outputs(422) <= not(layer0_outputs(2453));
    outputs(423) <= not(layer0_outputs(1878)) or (layer0_outputs(7190));
    outputs(424) <= not(layer0_outputs(6735)) or (layer0_outputs(1928));
    outputs(425) <= not((layer0_outputs(7050)) xor (layer0_outputs(4456)));
    outputs(426) <= (layer0_outputs(1074)) xor (layer0_outputs(848));
    outputs(427) <= not((layer0_outputs(5033)) and (layer0_outputs(372)));
    outputs(428) <= not(layer0_outputs(4558));
    outputs(429) <= not((layer0_outputs(1630)) xor (layer0_outputs(605)));
    outputs(430) <= (layer0_outputs(5848)) xor (layer0_outputs(3706));
    outputs(431) <= layer0_outputs(3093);
    outputs(432) <= not((layer0_outputs(1298)) xor (layer0_outputs(99)));
    outputs(433) <= not(layer0_outputs(2858)) or (layer0_outputs(6130));
    outputs(434) <= (layer0_outputs(2112)) and not (layer0_outputs(632));
    outputs(435) <= not(layer0_outputs(5060));
    outputs(436) <= layer0_outputs(186);
    outputs(437) <= (layer0_outputs(1596)) or (layer0_outputs(3587));
    outputs(438) <= not(layer0_outputs(3675));
    outputs(439) <= not((layer0_outputs(2141)) xor (layer0_outputs(6434)));
    outputs(440) <= not(layer0_outputs(2391));
    outputs(441) <= not((layer0_outputs(7105)) xor (layer0_outputs(5335)));
    outputs(442) <= not(layer0_outputs(6399));
    outputs(443) <= not(layer0_outputs(5514));
    outputs(444) <= layer0_outputs(3289);
    outputs(445) <= layer0_outputs(4272);
    outputs(446) <= layer0_outputs(927);
    outputs(447) <= not(layer0_outputs(6369));
    outputs(448) <= not(layer0_outputs(1294)) or (layer0_outputs(4959));
    outputs(449) <= (layer0_outputs(239)) xor (layer0_outputs(7080));
    outputs(450) <= not((layer0_outputs(7149)) xor (layer0_outputs(3734)));
    outputs(451) <= (layer0_outputs(767)) and not (layer0_outputs(3004));
    outputs(452) <= not((layer0_outputs(843)) and (layer0_outputs(3642)));
    outputs(453) <= (layer0_outputs(4810)) xor (layer0_outputs(4896));
    outputs(454) <= not((layer0_outputs(4861)) xor (layer0_outputs(1341)));
    outputs(455) <= not(layer0_outputs(3846));
    outputs(456) <= not(layer0_outputs(3285));
    outputs(457) <= layer0_outputs(4311);
    outputs(458) <= not(layer0_outputs(1854)) or (layer0_outputs(6282));
    outputs(459) <= layer0_outputs(998);
    outputs(460) <= layer0_outputs(3419);
    outputs(461) <= (layer0_outputs(5973)) or (layer0_outputs(3652));
    outputs(462) <= not((layer0_outputs(6485)) xor (layer0_outputs(4023)));
    outputs(463) <= not(layer0_outputs(5329));
    outputs(464) <= not((layer0_outputs(7346)) or (layer0_outputs(6409)));
    outputs(465) <= not(layer0_outputs(5712));
    outputs(466) <= not(layer0_outputs(1135));
    outputs(467) <= layer0_outputs(5988);
    outputs(468) <= not(layer0_outputs(2426));
    outputs(469) <= not((layer0_outputs(1044)) and (layer0_outputs(2139)));
    outputs(470) <= (layer0_outputs(736)) xor (layer0_outputs(620));
    outputs(471) <= (layer0_outputs(2336)) and (layer0_outputs(3516));
    outputs(472) <= (layer0_outputs(3725)) or (layer0_outputs(5872));
    outputs(473) <= (layer0_outputs(7591)) xor (layer0_outputs(3456));
    outputs(474) <= not((layer0_outputs(2401)) xor (layer0_outputs(3815)));
    outputs(475) <= layer0_outputs(3465);
    outputs(476) <= not(layer0_outputs(1021));
    outputs(477) <= not(layer0_outputs(296));
    outputs(478) <= (layer0_outputs(6357)) xor (layer0_outputs(7445));
    outputs(479) <= (layer0_outputs(4123)) or (layer0_outputs(4836));
    outputs(480) <= not((layer0_outputs(2128)) or (layer0_outputs(7574)));
    outputs(481) <= not(layer0_outputs(7338));
    outputs(482) <= not(layer0_outputs(7334));
    outputs(483) <= (layer0_outputs(6339)) and not (layer0_outputs(3198));
    outputs(484) <= layer0_outputs(463);
    outputs(485) <= not(layer0_outputs(5154));
    outputs(486) <= not((layer0_outputs(6657)) and (layer0_outputs(6071)));
    outputs(487) <= (layer0_outputs(5946)) and not (layer0_outputs(3));
    outputs(488) <= not((layer0_outputs(285)) xor (layer0_outputs(4248)));
    outputs(489) <= not(layer0_outputs(3738));
    outputs(490) <= not((layer0_outputs(2003)) xor (layer0_outputs(5591)));
    outputs(491) <= (layer0_outputs(2998)) and (layer0_outputs(1159));
    outputs(492) <= layer0_outputs(6368);
    outputs(493) <= (layer0_outputs(4510)) or (layer0_outputs(6161));
    outputs(494) <= (layer0_outputs(5592)) and not (layer0_outputs(5970));
    outputs(495) <= (layer0_outputs(3472)) xor (layer0_outputs(1650));
    outputs(496) <= not(layer0_outputs(4595));
    outputs(497) <= layer0_outputs(7573);
    outputs(498) <= not(layer0_outputs(203));
    outputs(499) <= (layer0_outputs(1244)) xor (layer0_outputs(2581));
    outputs(500) <= layer0_outputs(778);
    outputs(501) <= not(layer0_outputs(5682)) or (layer0_outputs(4129));
    outputs(502) <= layer0_outputs(2530);
    outputs(503) <= not(layer0_outputs(6690));
    outputs(504) <= not(layer0_outputs(5338)) or (layer0_outputs(6539));
    outputs(505) <= layer0_outputs(6669);
    outputs(506) <= not(layer0_outputs(7350));
    outputs(507) <= (layer0_outputs(7406)) xor (layer0_outputs(2283));
    outputs(508) <= (layer0_outputs(4745)) xor (layer0_outputs(1412));
    outputs(509) <= not((layer0_outputs(2370)) xor (layer0_outputs(672)));
    outputs(510) <= not(layer0_outputs(6159)) or (layer0_outputs(6900));
    outputs(511) <= not(layer0_outputs(505));
    outputs(512) <= layer0_outputs(2667);
    outputs(513) <= layer0_outputs(3144);
    outputs(514) <= layer0_outputs(7206);
    outputs(515) <= (layer0_outputs(2264)) xor (layer0_outputs(5000));
    outputs(516) <= not((layer0_outputs(7547)) and (layer0_outputs(315)));
    outputs(517) <= layer0_outputs(5325);
    outputs(518) <= not(layer0_outputs(5110)) or (layer0_outputs(894));
    outputs(519) <= (layer0_outputs(3755)) xor (layer0_outputs(599));
    outputs(520) <= layer0_outputs(4667);
    outputs(521) <= not(layer0_outputs(1789));
    outputs(522) <= layer0_outputs(7250);
    outputs(523) <= layer0_outputs(5500);
    outputs(524) <= (layer0_outputs(5356)) xor (layer0_outputs(4069));
    outputs(525) <= not((layer0_outputs(2923)) xor (layer0_outputs(2663)));
    outputs(526) <= layer0_outputs(6099);
    outputs(527) <= layer0_outputs(3240);
    outputs(528) <= (layer0_outputs(1844)) and (layer0_outputs(5948));
    outputs(529) <= not(layer0_outputs(1216)) or (layer0_outputs(6830));
    outputs(530) <= (layer0_outputs(5624)) and not (layer0_outputs(13));
    outputs(531) <= not(layer0_outputs(1367));
    outputs(532) <= (layer0_outputs(2513)) and (layer0_outputs(6302));
    outputs(533) <= not((layer0_outputs(1873)) or (layer0_outputs(2953)));
    outputs(534) <= (layer0_outputs(6980)) or (layer0_outputs(5854));
    outputs(535) <= not((layer0_outputs(1747)) xor (layer0_outputs(2291)));
    outputs(536) <= not(layer0_outputs(688));
    outputs(537) <= layer0_outputs(990);
    outputs(538) <= layer0_outputs(4696);
    outputs(539) <= (layer0_outputs(2082)) and (layer0_outputs(1665));
    outputs(540) <= not((layer0_outputs(5107)) xor (layer0_outputs(3136)));
    outputs(541) <= layer0_outputs(3194);
    outputs(542) <= not(layer0_outputs(1708)) or (layer0_outputs(5797));
    outputs(543) <= (layer0_outputs(3613)) and not (layer0_outputs(346));
    outputs(544) <= not(layer0_outputs(6650));
    outputs(545) <= layer0_outputs(7187);
    outputs(546) <= layer0_outputs(3935);
    outputs(547) <= not(layer0_outputs(1331));
    outputs(548) <= not(layer0_outputs(4828));
    outputs(549) <= layer0_outputs(4691);
    outputs(550) <= layer0_outputs(7603);
    outputs(551) <= not(layer0_outputs(3914));
    outputs(552) <= (layer0_outputs(4947)) xor (layer0_outputs(4246));
    outputs(553) <= not((layer0_outputs(4221)) xor (layer0_outputs(822)));
    outputs(554) <= '1';
    outputs(555) <= not(layer0_outputs(4522));
    outputs(556) <= (layer0_outputs(6358)) xor (layer0_outputs(1718));
    outputs(557) <= not(layer0_outputs(3510));
    outputs(558) <= not(layer0_outputs(3877)) or (layer0_outputs(5810));
    outputs(559) <= not(layer0_outputs(1457)) or (layer0_outputs(6123));
    outputs(560) <= layer0_outputs(738);
    outputs(561) <= not(layer0_outputs(1685));
    outputs(562) <= not(layer0_outputs(2918));
    outputs(563) <= not(layer0_outputs(7415)) or (layer0_outputs(859));
    outputs(564) <= not(layer0_outputs(1397));
    outputs(565) <= layer0_outputs(1346);
    outputs(566) <= layer0_outputs(2056);
    outputs(567) <= layer0_outputs(4068);
    outputs(568) <= not((layer0_outputs(557)) or (layer0_outputs(6589)));
    outputs(569) <= (layer0_outputs(6490)) or (layer0_outputs(6372));
    outputs(570) <= not(layer0_outputs(6079)) or (layer0_outputs(1664));
    outputs(571) <= layer0_outputs(6613);
    outputs(572) <= not(layer0_outputs(6852));
    outputs(573) <= layer0_outputs(2495);
    outputs(574) <= layer0_outputs(4410);
    outputs(575) <= (layer0_outputs(2237)) and not (layer0_outputs(7605));
    outputs(576) <= (layer0_outputs(5564)) and not (layer0_outputs(4043));
    outputs(577) <= not(layer0_outputs(1556));
    outputs(578) <= not((layer0_outputs(5446)) xor (layer0_outputs(4042)));
    outputs(579) <= (layer0_outputs(4983)) xor (layer0_outputs(3625));
    outputs(580) <= not(layer0_outputs(5140)) or (layer0_outputs(3167));
    outputs(581) <= not(layer0_outputs(709)) or (layer0_outputs(7172));
    outputs(582) <= (layer0_outputs(183)) xor (layer0_outputs(2736));
    outputs(583) <= not((layer0_outputs(1907)) xor (layer0_outputs(2930)));
    outputs(584) <= not(layer0_outputs(1585));
    outputs(585) <= (layer0_outputs(496)) xor (layer0_outputs(7131));
    outputs(586) <= not(layer0_outputs(618));
    outputs(587) <= not(layer0_outputs(4340)) or (layer0_outputs(2824));
    outputs(588) <= layer0_outputs(414);
    outputs(589) <= not((layer0_outputs(1450)) and (layer0_outputs(2756)));
    outputs(590) <= (layer0_outputs(4526)) xor (layer0_outputs(29));
    outputs(591) <= not((layer0_outputs(1034)) xor (layer0_outputs(2604)));
    outputs(592) <= layer0_outputs(1328);
    outputs(593) <= layer0_outputs(5311);
    outputs(594) <= not(layer0_outputs(1210));
    outputs(595) <= layer0_outputs(1622);
    outputs(596) <= layer0_outputs(4650);
    outputs(597) <= not((layer0_outputs(3222)) or (layer0_outputs(6847)));
    outputs(598) <= (layer0_outputs(5774)) and not (layer0_outputs(7129));
    outputs(599) <= (layer0_outputs(6789)) and not (layer0_outputs(1988));
    outputs(600) <= not(layer0_outputs(5390));
    outputs(601) <= (layer0_outputs(7123)) or (layer0_outputs(6579));
    outputs(602) <= not((layer0_outputs(109)) xor (layer0_outputs(1624)));
    outputs(603) <= not((layer0_outputs(5062)) xor (layer0_outputs(4162)));
    outputs(604) <= not(layer0_outputs(3926)) or (layer0_outputs(1388));
    outputs(605) <= not(layer0_outputs(1519));
    outputs(606) <= not(layer0_outputs(328));
    outputs(607) <= (layer0_outputs(3981)) and not (layer0_outputs(130));
    outputs(608) <= not(layer0_outputs(1642));
    outputs(609) <= (layer0_outputs(5370)) or (layer0_outputs(3303));
    outputs(610) <= not(layer0_outputs(71));
    outputs(611) <= not((layer0_outputs(7650)) xor (layer0_outputs(5670)));
    outputs(612) <= layer0_outputs(6373);
    outputs(613) <= not(layer0_outputs(5555));
    outputs(614) <= (layer0_outputs(974)) or (layer0_outputs(6502));
    outputs(615) <= not(layer0_outputs(4468)) or (layer0_outputs(3154));
    outputs(616) <= (layer0_outputs(1315)) xor (layer0_outputs(1880));
    outputs(617) <= not(layer0_outputs(1441));
    outputs(618) <= layer0_outputs(2182);
    outputs(619) <= not(layer0_outputs(3718));
    outputs(620) <= not(layer0_outputs(1309)) or (layer0_outputs(3530));
    outputs(621) <= not(layer0_outputs(6308)) or (layer0_outputs(1843));
    outputs(622) <= not(layer0_outputs(792));
    outputs(623) <= not(layer0_outputs(5808));
    outputs(624) <= (layer0_outputs(1507)) and not (layer0_outputs(7593));
    outputs(625) <= not(layer0_outputs(3399));
    outputs(626) <= (layer0_outputs(2886)) and (layer0_outputs(7374));
    outputs(627) <= not((layer0_outputs(6153)) xor (layer0_outputs(5480)));
    outputs(628) <= (layer0_outputs(6594)) xor (layer0_outputs(3886));
    outputs(629) <= not(layer0_outputs(817));
    outputs(630) <= (layer0_outputs(5474)) and (layer0_outputs(6994));
    outputs(631) <= not(layer0_outputs(7041)) or (layer0_outputs(5755));
    outputs(632) <= layer0_outputs(6491);
    outputs(633) <= (layer0_outputs(2402)) and not (layer0_outputs(5625));
    outputs(634) <= layer0_outputs(4442);
    outputs(635) <= not(layer0_outputs(7480));
    outputs(636) <= not((layer0_outputs(2819)) or (layer0_outputs(5218)));
    outputs(637) <= layer0_outputs(7287);
    outputs(638) <= not(layer0_outputs(3196));
    outputs(639) <= (layer0_outputs(1394)) xor (layer0_outputs(6329));
    outputs(640) <= not((layer0_outputs(2640)) and (layer0_outputs(2471)));
    outputs(641) <= not((layer0_outputs(5536)) or (layer0_outputs(6826)));
    outputs(642) <= not(layer0_outputs(3817));
    outputs(643) <= (layer0_outputs(1169)) and not (layer0_outputs(4369));
    outputs(644) <= layer0_outputs(4803);
    outputs(645) <= (layer0_outputs(1109)) and not (layer0_outputs(1403));
    outputs(646) <= (layer0_outputs(4625)) xor (layer0_outputs(4480));
    outputs(647) <= not((layer0_outputs(6835)) and (layer0_outputs(107)));
    outputs(648) <= not(layer0_outputs(1729));
    outputs(649) <= not(layer0_outputs(7363));
    outputs(650) <= not(layer0_outputs(1117));
    outputs(651) <= not(layer0_outputs(1578));
    outputs(652) <= not((layer0_outputs(6154)) xor (layer0_outputs(1593)));
    outputs(653) <= (layer0_outputs(3506)) or (layer0_outputs(1884));
    outputs(654) <= not((layer0_outputs(4697)) xor (layer0_outputs(550)));
    outputs(655) <= not(layer0_outputs(880));
    outputs(656) <= (layer0_outputs(3207)) and (layer0_outputs(994));
    outputs(657) <= not((layer0_outputs(3702)) xor (layer0_outputs(6169)));
    outputs(658) <= layer0_outputs(290);
    outputs(659) <= layer0_outputs(4301);
    outputs(660) <= not(layer0_outputs(4543));
    outputs(661) <= not(layer0_outputs(527));
    outputs(662) <= not(layer0_outputs(6461));
    outputs(663) <= not((layer0_outputs(7025)) and (layer0_outputs(5717)));
    outputs(664) <= layer0_outputs(6996);
    outputs(665) <= not(layer0_outputs(5249));
    outputs(666) <= not((layer0_outputs(227)) or (layer0_outputs(276)));
    outputs(667) <= not(layer0_outputs(1140));
    outputs(668) <= layer0_outputs(7541);
    outputs(669) <= not(layer0_outputs(4544)) or (layer0_outputs(5032));
    outputs(670) <= not(layer0_outputs(3918));
    outputs(671) <= not(layer0_outputs(2951));
    outputs(672) <= not(layer0_outputs(710));
    outputs(673) <= layer0_outputs(2906);
    outputs(674) <= layer0_outputs(1786);
    outputs(675) <= (layer0_outputs(5142)) xor (layer0_outputs(5618));
    outputs(676) <= (layer0_outputs(1489)) xor (layer0_outputs(1306));
    outputs(677) <= layer0_outputs(6482);
    outputs(678) <= not(layer0_outputs(5201)) or (layer0_outputs(5321));
    outputs(679) <= not(layer0_outputs(3535));
    outputs(680) <= not(layer0_outputs(5290));
    outputs(681) <= layer0_outputs(7673);
    outputs(682) <= not(layer0_outputs(189)) or (layer0_outputs(1018));
    outputs(683) <= layer0_outputs(4706);
    outputs(684) <= layer0_outputs(1483);
    outputs(685) <= (layer0_outputs(5690)) xor (layer0_outputs(5537));
    outputs(686) <= (layer0_outputs(7298)) and not (layer0_outputs(13));
    outputs(687) <= layer0_outputs(1437);
    outputs(688) <= not((layer0_outputs(25)) and (layer0_outputs(4365)));
    outputs(689) <= not(layer0_outputs(4496)) or (layer0_outputs(5898));
    outputs(690) <= not((layer0_outputs(7003)) xor (layer0_outputs(2474)));
    outputs(691) <= not(layer0_outputs(4671));
    outputs(692) <= (layer0_outputs(4245)) xor (layer0_outputs(1577));
    outputs(693) <= not(layer0_outputs(5042));
    outputs(694) <= layer0_outputs(5211);
    outputs(695) <= not((layer0_outputs(391)) xor (layer0_outputs(6180)));
    outputs(696) <= not((layer0_outputs(5285)) and (layer0_outputs(2711)));
    outputs(697) <= not(layer0_outputs(867)) or (layer0_outputs(4028));
    outputs(698) <= layer0_outputs(921);
    outputs(699) <= layer0_outputs(1657);
    outputs(700) <= not((layer0_outputs(5035)) xor (layer0_outputs(4632)));
    outputs(701) <= (layer0_outputs(3046)) xor (layer0_outputs(856));
    outputs(702) <= (layer0_outputs(1153)) xor (layer0_outputs(4858));
    outputs(703) <= layer0_outputs(4358);
    outputs(704) <= layer0_outputs(4840);
    outputs(705) <= not(layer0_outputs(1440)) or (layer0_outputs(7527));
    outputs(706) <= not((layer0_outputs(3818)) and (layer0_outputs(6460)));
    outputs(707) <= (layer0_outputs(4034)) and not (layer0_outputs(1915));
    outputs(708) <= (layer0_outputs(5671)) and (layer0_outputs(2436));
    outputs(709) <= not(layer0_outputs(6453)) or (layer0_outputs(565));
    outputs(710) <= not(layer0_outputs(3836)) or (layer0_outputs(3306));
    outputs(711) <= layer0_outputs(2392);
    outputs(712) <= (layer0_outputs(2614)) xor (layer0_outputs(7261));
    outputs(713) <= not((layer0_outputs(351)) xor (layer0_outputs(1949)));
    outputs(714) <= layer0_outputs(2861);
    outputs(715) <= (layer0_outputs(6923)) and (layer0_outputs(2538));
    outputs(716) <= (layer0_outputs(969)) and not (layer0_outputs(380));
    outputs(717) <= layer0_outputs(1259);
    outputs(718) <= not(layer0_outputs(5543));
    outputs(719) <= not((layer0_outputs(2610)) xor (layer0_outputs(3640)));
    outputs(720) <= (layer0_outputs(4453)) and (layer0_outputs(5762));
    outputs(721) <= (layer0_outputs(1894)) xor (layer0_outputs(5867));
    outputs(722) <= (layer0_outputs(5757)) xor (layer0_outputs(7560));
    outputs(723) <= not(layer0_outputs(3489)) or (layer0_outputs(2159));
    outputs(724) <= (layer0_outputs(4682)) or (layer0_outputs(3372));
    outputs(725) <= layer0_outputs(2042);
    outputs(726) <= not(layer0_outputs(1939));
    outputs(727) <= layer0_outputs(7422);
    outputs(728) <= (layer0_outputs(4071)) xor (layer0_outputs(5885));
    outputs(729) <= layer0_outputs(7652);
    outputs(730) <= not((layer0_outputs(4674)) xor (layer0_outputs(5957)));
    outputs(731) <= not((layer0_outputs(4133)) xor (layer0_outputs(440)));
    outputs(732) <= layer0_outputs(7108);
    outputs(733) <= not(layer0_outputs(5429));
    outputs(734) <= not(layer0_outputs(6927));
    outputs(735) <= (layer0_outputs(3777)) and not (layer0_outputs(6052));
    outputs(736) <= not(layer0_outputs(1498));
    outputs(737) <= (layer0_outputs(3757)) and not (layer0_outputs(3653));
    outputs(738) <= not(layer0_outputs(7340));
    outputs(739) <= layer0_outputs(3460);
    outputs(740) <= not((layer0_outputs(4448)) xor (layer0_outputs(5965)));
    outputs(741) <= not(layer0_outputs(7634));
    outputs(742) <= not(layer0_outputs(621));
    outputs(743) <= not(layer0_outputs(1755));
    outputs(744) <= layer0_outputs(4003);
    outputs(745) <= (layer0_outputs(681)) xor (layer0_outputs(6714));
    outputs(746) <= not(layer0_outputs(6357)) or (layer0_outputs(3647));
    outputs(747) <= not(layer0_outputs(3251));
    outputs(748) <= layer0_outputs(6740);
    outputs(749) <= not((layer0_outputs(711)) xor (layer0_outputs(1810)));
    outputs(750) <= not(layer0_outputs(2966));
    outputs(751) <= not(layer0_outputs(6767));
    outputs(752) <= not(layer0_outputs(1674)) or (layer0_outputs(7034));
    outputs(753) <= layer0_outputs(7100);
    outputs(754) <= layer0_outputs(5256);
    outputs(755) <= layer0_outputs(3272);
    outputs(756) <= not(layer0_outputs(7311)) or (layer0_outputs(4237));
    outputs(757) <= layer0_outputs(7582);
    outputs(758) <= not(layer0_outputs(2068));
    outputs(759) <= not((layer0_outputs(4108)) and (layer0_outputs(7451)));
    outputs(760) <= (layer0_outputs(1350)) and not (layer0_outputs(7294));
    outputs(761) <= (layer0_outputs(4198)) or (layer0_outputs(1086));
    outputs(762) <= not(layer0_outputs(6564));
    outputs(763) <= (layer0_outputs(2210)) or (layer0_outputs(2142));
    outputs(764) <= layer0_outputs(2530);
    outputs(765) <= layer0_outputs(6579);
    outputs(766) <= (layer0_outputs(5515)) and not (layer0_outputs(7228));
    outputs(767) <= (layer0_outputs(5612)) and not (layer0_outputs(428));
    outputs(768) <= (layer0_outputs(2841)) and (layer0_outputs(118));
    outputs(769) <= not(layer0_outputs(4890));
    outputs(770) <= not(layer0_outputs(7613));
    outputs(771) <= (layer0_outputs(6380)) and not (layer0_outputs(5247));
    outputs(772) <= not(layer0_outputs(5264));
    outputs(773) <= (layer0_outputs(5049)) and not (layer0_outputs(7317));
    outputs(774) <= not((layer0_outputs(2692)) or (layer0_outputs(6449)));
    outputs(775) <= (layer0_outputs(6400)) xor (layer0_outputs(2776));
    outputs(776) <= (layer0_outputs(236)) and not (layer0_outputs(1592));
    outputs(777) <= (layer0_outputs(2102)) and not (layer0_outputs(2953));
    outputs(778) <= not(layer0_outputs(678));
    outputs(779) <= (layer0_outputs(1037)) xor (layer0_outputs(5192));
    outputs(780) <= not((layer0_outputs(2676)) or (layer0_outputs(4866)));
    outputs(781) <= (layer0_outputs(7158)) xor (layer0_outputs(6489));
    outputs(782) <= not((layer0_outputs(6703)) or (layer0_outputs(5422)));
    outputs(783) <= not((layer0_outputs(4218)) xor (layer0_outputs(7572)));
    outputs(784) <= (layer0_outputs(7234)) and not (layer0_outputs(2782));
    outputs(785) <= not(layer0_outputs(6516));
    outputs(786) <= layer0_outputs(3274);
    outputs(787) <= not(layer0_outputs(5482));
    outputs(788) <= (layer0_outputs(7350)) and not (layer0_outputs(6664));
    outputs(789) <= (layer0_outputs(6318)) and not (layer0_outputs(7119));
    outputs(790) <= (layer0_outputs(5574)) and not (layer0_outputs(385));
    outputs(791) <= layer0_outputs(1266);
    outputs(792) <= (layer0_outputs(6944)) and not (layer0_outputs(6919));
    outputs(793) <= layer0_outputs(2425);
    outputs(794) <= (layer0_outputs(7319)) and (layer0_outputs(6969));
    outputs(795) <= layer0_outputs(2463);
    outputs(796) <= (layer0_outputs(6639)) and not (layer0_outputs(1993));
    outputs(797) <= (layer0_outputs(6832)) xor (layer0_outputs(1396));
    outputs(798) <= not((layer0_outputs(1616)) xor (layer0_outputs(3704)));
    outputs(799) <= (layer0_outputs(7479)) and (layer0_outputs(5055));
    outputs(800) <= not(layer0_outputs(1644));
    outputs(801) <= not((layer0_outputs(5306)) or (layer0_outputs(6886)));
    outputs(802) <= layer0_outputs(2012);
    outputs(803) <= not(layer0_outputs(2308));
    outputs(804) <= (layer0_outputs(5640)) and not (layer0_outputs(3766));
    outputs(805) <= not((layer0_outputs(3363)) xor (layer0_outputs(1224)));
    outputs(806) <= not((layer0_outputs(3799)) or (layer0_outputs(5676)));
    outputs(807) <= (layer0_outputs(4819)) and not (layer0_outputs(6514));
    outputs(808) <= (layer0_outputs(3045)) or (layer0_outputs(6471));
    outputs(809) <= (layer0_outputs(3193)) or (layer0_outputs(4863));
    outputs(810) <= not(layer0_outputs(972));
    outputs(811) <= (layer0_outputs(7138)) and not (layer0_outputs(514));
    outputs(812) <= not((layer0_outputs(6613)) or (layer0_outputs(7577)));
    outputs(813) <= layer0_outputs(7561);
    outputs(814) <= (layer0_outputs(1649)) and (layer0_outputs(3378));
    outputs(815) <= not(layer0_outputs(6402));
    outputs(816) <= (layer0_outputs(72)) xor (layer0_outputs(5642));
    outputs(817) <= (layer0_outputs(3619)) and (layer0_outputs(3798));
    outputs(818) <= (layer0_outputs(669)) and not (layer0_outputs(1866));
    outputs(819) <= (layer0_outputs(1196)) xor (layer0_outputs(6762));
    outputs(820) <= (layer0_outputs(1457)) and not (layer0_outputs(2635));
    outputs(821) <= not((layer0_outputs(4793)) or (layer0_outputs(3302)));
    outputs(822) <= not(layer0_outputs(2661)) or (layer0_outputs(3538));
    outputs(823) <= not(layer0_outputs(2973));
    outputs(824) <= (layer0_outputs(20)) and not (layer0_outputs(4347));
    outputs(825) <= (layer0_outputs(6469)) xor (layer0_outputs(6741));
    outputs(826) <= (layer0_outputs(3385)) and not (layer0_outputs(517));
    outputs(827) <= not((layer0_outputs(6847)) xor (layer0_outputs(2741)));
    outputs(828) <= not(layer0_outputs(3525));
    outputs(829) <= layer0_outputs(1697);
    outputs(830) <= (layer0_outputs(2315)) and not (layer0_outputs(5606));
    outputs(831) <= not(layer0_outputs(4400));
    outputs(832) <= (layer0_outputs(3368)) and not (layer0_outputs(6303));
    outputs(833) <= not(layer0_outputs(2105));
    outputs(834) <= (layer0_outputs(6520)) and (layer0_outputs(2939));
    outputs(835) <= (layer0_outputs(511)) and not (layer0_outputs(3997));
    outputs(836) <= (layer0_outputs(7501)) xor (layer0_outputs(7460));
    outputs(837) <= (layer0_outputs(3890)) and not (layer0_outputs(736));
    outputs(838) <= not((layer0_outputs(1513)) or (layer0_outputs(1214)));
    outputs(839) <= (layer0_outputs(2108)) and not (layer0_outputs(666));
    outputs(840) <= layer0_outputs(3825);
    outputs(841) <= (layer0_outputs(533)) and not (layer0_outputs(7410));
    outputs(842) <= not((layer0_outputs(5889)) or (layer0_outputs(3523)));
    outputs(843) <= not(layer0_outputs(7463));
    outputs(844) <= not(layer0_outputs(3043)) or (layer0_outputs(2965));
    outputs(845) <= not(layer0_outputs(6097));
    outputs(846) <= layer0_outputs(2376);
    outputs(847) <= not(layer0_outputs(3325));
    outputs(848) <= (layer0_outputs(4723)) and not (layer0_outputs(48));
    outputs(849) <= not(layer0_outputs(6833));
    outputs(850) <= not(layer0_outputs(3002));
    outputs(851) <= not((layer0_outputs(2628)) xor (layer0_outputs(3943)));
    outputs(852) <= (layer0_outputs(2978)) and (layer0_outputs(5334));
    outputs(853) <= (layer0_outputs(2149)) and (layer0_outputs(1449));
    outputs(854) <= (layer0_outputs(6109)) and (layer0_outputs(3762));
    outputs(855) <= layer0_outputs(3965);
    outputs(856) <= (layer0_outputs(5715)) and not (layer0_outputs(908));
    outputs(857) <= (layer0_outputs(4344)) xor (layer0_outputs(3962));
    outputs(858) <= (layer0_outputs(2807)) xor (layer0_outputs(5138));
    outputs(859) <= (layer0_outputs(7031)) and (layer0_outputs(3636));
    outputs(860) <= (layer0_outputs(1174)) and (layer0_outputs(7655));
    outputs(861) <= (layer0_outputs(7414)) xor (layer0_outputs(3704));
    outputs(862) <= not((layer0_outputs(4428)) or (layer0_outputs(7328)));
    outputs(863) <= (layer0_outputs(7624)) and (layer0_outputs(1816));
    outputs(864) <= not(layer0_outputs(5651));
    outputs(865) <= (layer0_outputs(41)) and (layer0_outputs(2459));
    outputs(866) <= not(layer0_outputs(7576));
    outputs(867) <= not((layer0_outputs(6248)) xor (layer0_outputs(2661)));
    outputs(868) <= not(layer0_outputs(7124));
    outputs(869) <= not(layer0_outputs(4727));
    outputs(870) <= (layer0_outputs(2996)) and not (layer0_outputs(4268));
    outputs(871) <= (layer0_outputs(3856)) and not (layer0_outputs(230));
    outputs(872) <= (layer0_outputs(2599)) and not (layer0_outputs(463));
    outputs(873) <= not(layer0_outputs(3830));
    outputs(874) <= '0';
    outputs(875) <= (layer0_outputs(5674)) and not (layer0_outputs(5136));
    outputs(876) <= layer0_outputs(2169);
    outputs(877) <= layer0_outputs(4893);
    outputs(878) <= '0';
    outputs(879) <= not(layer0_outputs(5817));
    outputs(880) <= (layer0_outputs(5543)) and not (layer0_outputs(3987));
    outputs(881) <= (layer0_outputs(5413)) and (layer0_outputs(6814));
    outputs(882) <= not((layer0_outputs(396)) xor (layer0_outputs(1409)));
    outputs(883) <= not(layer0_outputs(5216));
    outputs(884) <= (layer0_outputs(1640)) and not (layer0_outputs(7126));
    outputs(885) <= (layer0_outputs(7370)) and not (layer0_outputs(2410));
    outputs(886) <= (layer0_outputs(1233)) and not (layer0_outputs(4821));
    outputs(887) <= not(layer0_outputs(6105));
    outputs(888) <= not(layer0_outputs(729));
    outputs(889) <= (layer0_outputs(2115)) and not (layer0_outputs(617));
    outputs(890) <= not((layer0_outputs(116)) or (layer0_outputs(5002)));
    outputs(891) <= (layer0_outputs(334)) and not (layer0_outputs(6696));
    outputs(892) <= not(layer0_outputs(416));
    outputs(893) <= (layer0_outputs(4082)) and not (layer0_outputs(4857));
    outputs(894) <= (layer0_outputs(2869)) and (layer0_outputs(3257));
    outputs(895) <= layer0_outputs(3679);
    outputs(896) <= layer0_outputs(291);
    outputs(897) <= (layer0_outputs(4693)) and (layer0_outputs(6361));
    outputs(898) <= not(layer0_outputs(7280));
    outputs(899) <= (layer0_outputs(6454)) xor (layer0_outputs(695));
    outputs(900) <= (layer0_outputs(3839)) and not (layer0_outputs(5550));
    outputs(901) <= (layer0_outputs(6333)) and not (layer0_outputs(346));
    outputs(902) <= not((layer0_outputs(7461)) or (layer0_outputs(2938)));
    outputs(903) <= (layer0_outputs(2021)) and not (layer0_outputs(3504));
    outputs(904) <= (layer0_outputs(5630)) and not (layer0_outputs(6197));
    outputs(905) <= not((layer0_outputs(5927)) or (layer0_outputs(7072)));
    outputs(906) <= (layer0_outputs(1057)) and (layer0_outputs(3057));
    outputs(907) <= (layer0_outputs(5999)) xor (layer0_outputs(5381));
    outputs(908) <= (layer0_outputs(4031)) and not (layer0_outputs(7395));
    outputs(909) <= '0';
    outputs(910) <= (layer0_outputs(4838)) and not (layer0_outputs(3112));
    outputs(911) <= (layer0_outputs(262)) and not (layer0_outputs(1997));
    outputs(912) <= (layer0_outputs(6629)) and not (layer0_outputs(5480));
    outputs(913) <= not((layer0_outputs(2172)) or (layer0_outputs(4221)));
    outputs(914) <= layer0_outputs(7094);
    outputs(915) <= (layer0_outputs(1230)) and not (layer0_outputs(347));
    outputs(916) <= (layer0_outputs(3870)) xor (layer0_outputs(3624));
    outputs(917) <= layer0_outputs(728);
    outputs(918) <= not(layer0_outputs(358));
    outputs(919) <= not(layer0_outputs(5742));
    outputs(920) <= layer0_outputs(4020);
    outputs(921) <= (layer0_outputs(3848)) and (layer0_outputs(4086));
    outputs(922) <= not((layer0_outputs(6149)) xor (layer0_outputs(6263)));
    outputs(923) <= (layer0_outputs(2452)) and not (layer0_outputs(5827));
    outputs(924) <= layer0_outputs(5460);
    outputs(925) <= not(layer0_outputs(2378));
    outputs(926) <= (layer0_outputs(5322)) and not (layer0_outputs(6334));
    outputs(927) <= not((layer0_outputs(2091)) or (layer0_outputs(4081)));
    outputs(928) <= (layer0_outputs(708)) and not (layer0_outputs(3056));
    outputs(929) <= not(layer0_outputs(6408));
    outputs(930) <= (layer0_outputs(1593)) and not (layer0_outputs(1788));
    outputs(931) <= not((layer0_outputs(5741)) or (layer0_outputs(6964)));
    outputs(932) <= (layer0_outputs(22)) and not (layer0_outputs(6796));
    outputs(933) <= '0';
    outputs(934) <= (layer0_outputs(756)) and (layer0_outputs(7039));
    outputs(935) <= not(layer0_outputs(1338));
    outputs(936) <= not(layer0_outputs(4688));
    outputs(937) <= not(layer0_outputs(2163));
    outputs(938) <= '0';
    outputs(939) <= layer0_outputs(984);
    outputs(940) <= not((layer0_outputs(3852)) or (layer0_outputs(1544)));
    outputs(941) <= (layer0_outputs(7675)) and (layer0_outputs(5573));
    outputs(942) <= layer0_outputs(1604);
    outputs(943) <= (layer0_outputs(4338)) and not (layer0_outputs(1255));
    outputs(944) <= (layer0_outputs(4397)) and (layer0_outputs(4220));
    outputs(945) <= (layer0_outputs(6620)) and (layer0_outputs(5748));
    outputs(946) <= not((layer0_outputs(6849)) or (layer0_outputs(5678)));
    outputs(947) <= not((layer0_outputs(1150)) or (layer0_outputs(2856)));
    outputs(948) <= (layer0_outputs(4054)) and not (layer0_outputs(1466));
    outputs(949) <= (layer0_outputs(19)) and not (layer0_outputs(1314));
    outputs(950) <= not(layer0_outputs(1459));
    outputs(951) <= not(layer0_outputs(1044));
    outputs(952) <= not(layer0_outputs(6630));
    outputs(953) <= (layer0_outputs(5057)) and (layer0_outputs(5649));
    outputs(954) <= (layer0_outputs(461)) and not (layer0_outputs(2652));
    outputs(955) <= (layer0_outputs(5672)) and (layer0_outputs(7151));
    outputs(956) <= not((layer0_outputs(2694)) xor (layer0_outputs(5767)));
    outputs(957) <= not(layer0_outputs(3108));
    outputs(958) <= (layer0_outputs(4950)) and not (layer0_outputs(5267));
    outputs(959) <= (layer0_outputs(6563)) and not (layer0_outputs(568));
    outputs(960) <= not(layer0_outputs(3892));
    outputs(961) <= not((layer0_outputs(1797)) or (layer0_outputs(5761)));
    outputs(962) <= not(layer0_outputs(1537));
    outputs(963) <= (layer0_outputs(4878)) and not (layer0_outputs(3074));
    outputs(964) <= not((layer0_outputs(2377)) or (layer0_outputs(2723)));
    outputs(965) <= not(layer0_outputs(2445));
    outputs(966) <= not((layer0_outputs(5320)) or (layer0_outputs(2863)));
    outputs(967) <= layer0_outputs(1641);
    outputs(968) <= (layer0_outputs(217)) xor (layer0_outputs(3883));
    outputs(969) <= not(layer0_outputs(5510));
    outputs(970) <= layer0_outputs(7059);
    outputs(971) <= not(layer0_outputs(6184)) or (layer0_outputs(7423));
    outputs(972) <= layer0_outputs(3355);
    outputs(973) <= (layer0_outputs(3831)) and not (layer0_outputs(1800));
    outputs(974) <= not((layer0_outputs(4578)) or (layer0_outputs(911)));
    outputs(975) <= (layer0_outputs(3467)) and not (layer0_outputs(2131));
    outputs(976) <= (layer0_outputs(2726)) and not (layer0_outputs(6760));
    outputs(977) <= (layer0_outputs(844)) and not (layer0_outputs(622));
    outputs(978) <= (layer0_outputs(6694)) and not (layer0_outputs(475));
    outputs(979) <= '0';
    outputs(980) <= not((layer0_outputs(1876)) xor (layer0_outputs(1480)));
    outputs(981) <= (layer0_outputs(3316)) and not (layer0_outputs(6737));
    outputs(982) <= (layer0_outputs(3031)) and (layer0_outputs(452));
    outputs(983) <= layer0_outputs(6010);
    outputs(984) <= (layer0_outputs(541)) xor (layer0_outputs(6275));
    outputs(985) <= (layer0_outputs(6432)) and not (layer0_outputs(5001));
    outputs(986) <= (layer0_outputs(1995)) xor (layer0_outputs(5242));
    outputs(987) <= (layer0_outputs(1829)) and not (layer0_outputs(5319));
    outputs(988) <= layer0_outputs(5486);
    outputs(989) <= (layer0_outputs(2950)) xor (layer0_outputs(6689));
    outputs(990) <= (layer0_outputs(1319)) and (layer0_outputs(7623));
    outputs(991) <= (layer0_outputs(3281)) and (layer0_outputs(5315));
    outputs(992) <= not(layer0_outputs(5622)) or (layer0_outputs(4849));
    outputs(993) <= not((layer0_outputs(1813)) or (layer0_outputs(4924)));
    outputs(994) <= not(layer0_outputs(4714));
    outputs(995) <= (layer0_outputs(2934)) and (layer0_outputs(735));
    outputs(996) <= (layer0_outputs(6813)) and not (layer0_outputs(6787));
    outputs(997) <= (layer0_outputs(6907)) and not (layer0_outputs(5598));
    outputs(998) <= not(layer0_outputs(2560));
    outputs(999) <= not(layer0_outputs(647));
    outputs(1000) <= (layer0_outputs(4562)) and not (layer0_outputs(2410));
    outputs(1001) <= layer0_outputs(6266);
    outputs(1002) <= not(layer0_outputs(7587));
    outputs(1003) <= layer0_outputs(3720);
    outputs(1004) <= not((layer0_outputs(482)) xor (layer0_outputs(5953)));
    outputs(1005) <= (layer0_outputs(279)) and not (layer0_outputs(4567));
    outputs(1006) <= not(layer0_outputs(6234));
    outputs(1007) <= layer0_outputs(3081);
    outputs(1008) <= (layer0_outputs(3612)) and not (layer0_outputs(1190));
    outputs(1009) <= (layer0_outputs(1026)) and not (layer0_outputs(3000));
    outputs(1010) <= not((layer0_outputs(2690)) xor (layer0_outputs(142)));
    outputs(1011) <= not(layer0_outputs(1467));
    outputs(1012) <= (layer0_outputs(1873)) and not (layer0_outputs(5314));
    outputs(1013) <= not(layer0_outputs(6820));
    outputs(1014) <= layer0_outputs(3931);
    outputs(1015) <= layer0_outputs(2239);
    outputs(1016) <= (layer0_outputs(7511)) and not (layer0_outputs(2301));
    outputs(1017) <= layer0_outputs(4970);
    outputs(1018) <= layer0_outputs(5348);
    outputs(1019) <= not((layer0_outputs(2396)) xor (layer0_outputs(3527)));
    outputs(1020) <= not(layer0_outputs(5443));
    outputs(1021) <= layer0_outputs(1826);
    outputs(1022) <= (layer0_outputs(6915)) and not (layer0_outputs(2231));
    outputs(1023) <= not(layer0_outputs(7556));
    outputs(1024) <= not((layer0_outputs(1885)) or (layer0_outputs(4360)));
    outputs(1025) <= not(layer0_outputs(5731));
    outputs(1026) <= not((layer0_outputs(3371)) xor (layer0_outputs(5114)));
    outputs(1027) <= (layer0_outputs(7084)) and not (layer0_outputs(7252));
    outputs(1028) <= (layer0_outputs(7373)) and not (layer0_outputs(1429));
    outputs(1029) <= not((layer0_outputs(351)) or (layer0_outputs(3557)));
    outputs(1030) <= (layer0_outputs(4589)) xor (layer0_outputs(460));
    outputs(1031) <= layer0_outputs(816);
    outputs(1032) <= layer0_outputs(2062);
    outputs(1033) <= not((layer0_outputs(3579)) or (layer0_outputs(3627)));
    outputs(1034) <= not((layer0_outputs(2587)) or (layer0_outputs(4929)));
    outputs(1035) <= '0';
    outputs(1036) <= (layer0_outputs(759)) and not (layer0_outputs(2492));
    outputs(1037) <= (layer0_outputs(1433)) xor (layer0_outputs(253));
    outputs(1038) <= (layer0_outputs(3415)) and not (layer0_outputs(2442));
    outputs(1039) <= not((layer0_outputs(4753)) and (layer0_outputs(1316)));
    outputs(1040) <= not(layer0_outputs(4431));
    outputs(1041) <= not(layer0_outputs(3390));
    outputs(1042) <= (layer0_outputs(5703)) and (layer0_outputs(3474));
    outputs(1043) <= (layer0_outputs(5554)) and not (layer0_outputs(28));
    outputs(1044) <= layer0_outputs(4355);
    outputs(1045) <= (layer0_outputs(4735)) and (layer0_outputs(4746));
    outputs(1046) <= not(layer0_outputs(2492));
    outputs(1047) <= not(layer0_outputs(3633));
    outputs(1048) <= '0';
    outputs(1049) <= (layer0_outputs(4328)) and (layer0_outputs(1774));
    outputs(1050) <= (layer0_outputs(581)) and not (layer0_outputs(6115));
    outputs(1051) <= (layer0_outputs(303)) and not (layer0_outputs(536));
    outputs(1052) <= layer0_outputs(6409);
    outputs(1053) <= not((layer0_outputs(1701)) or (layer0_outputs(2952)));
    outputs(1054) <= '0';
    outputs(1055) <= not((layer0_outputs(3509)) xor (layer0_outputs(5251)));
    outputs(1056) <= (layer0_outputs(5853)) and (layer0_outputs(2432));
    outputs(1057) <= (layer0_outputs(6196)) and not (layer0_outputs(6947));
    outputs(1058) <= layer0_outputs(5949);
    outputs(1059) <= '0';
    outputs(1060) <= not(layer0_outputs(989));
    outputs(1061) <= layer0_outputs(21);
    outputs(1062) <= layer0_outputs(6090);
    outputs(1063) <= not((layer0_outputs(7336)) xor (layer0_outputs(1537)));
    outputs(1064) <= not(layer0_outputs(3745));
    outputs(1065) <= layer0_outputs(1771);
    outputs(1066) <= not(layer0_outputs(3055));
    outputs(1067) <= not((layer0_outputs(1994)) xor (layer0_outputs(3501)));
    outputs(1068) <= not((layer0_outputs(6356)) xor (layer0_outputs(6355)));
    outputs(1069) <= not(layer0_outputs(5730)) or (layer0_outputs(5082));
    outputs(1070) <= not(layer0_outputs(3949));
    outputs(1071) <= (layer0_outputs(7599)) xor (layer0_outputs(6990));
    outputs(1072) <= layer0_outputs(3718);
    outputs(1073) <= not(layer0_outputs(5372));
    outputs(1074) <= layer0_outputs(6446);
    outputs(1075) <= (layer0_outputs(5548)) and not (layer0_outputs(3104));
    outputs(1076) <= (layer0_outputs(1399)) and not (layer0_outputs(1164));
    outputs(1077) <= (layer0_outputs(6587)) xor (layer0_outputs(6481));
    outputs(1078) <= (layer0_outputs(6404)) and (layer0_outputs(4334));
    outputs(1079) <= not((layer0_outputs(3852)) or (layer0_outputs(2871)));
    outputs(1080) <= not((layer0_outputs(3586)) xor (layer0_outputs(78)));
    outputs(1081) <= not(layer0_outputs(3865));
    outputs(1082) <= not((layer0_outputs(3439)) or (layer0_outputs(1076)));
    outputs(1083) <= layer0_outputs(7369);
    outputs(1084) <= not(layer0_outputs(414));
    outputs(1085) <= not((layer0_outputs(1069)) or (layer0_outputs(5119)));
    outputs(1086) <= (layer0_outputs(5212)) and (layer0_outputs(1243));
    outputs(1087) <= (layer0_outputs(5904)) and not (layer0_outputs(6888));
    outputs(1088) <= '0';
    outputs(1089) <= '0';
    outputs(1090) <= (layer0_outputs(5074)) and not (layer0_outputs(4113));
    outputs(1091) <= not(layer0_outputs(1080));
    outputs(1092) <= (layer0_outputs(3379)) and not (layer0_outputs(4768));
    outputs(1093) <= not(layer0_outputs(5482));
    outputs(1094) <= not((layer0_outputs(7361)) xor (layer0_outputs(6102)));
    outputs(1095) <= (layer0_outputs(2297)) and not (layer0_outputs(464));
    outputs(1096) <= layer0_outputs(5315);
    outputs(1097) <= (layer0_outputs(6051)) and (layer0_outputs(5212));
    outputs(1098) <= not(layer0_outputs(2074));
    outputs(1099) <= not((layer0_outputs(5489)) xor (layer0_outputs(2412)));
    outputs(1100) <= (layer0_outputs(3828)) and (layer0_outputs(1029));
    outputs(1101) <= (layer0_outputs(7122)) xor (layer0_outputs(6649));
    outputs(1102) <= (layer0_outputs(3531)) or (layer0_outputs(2166));
    outputs(1103) <= (layer0_outputs(4630)) and not (layer0_outputs(4114));
    outputs(1104) <= (layer0_outputs(6126)) and not (layer0_outputs(3547));
    outputs(1105) <= not((layer0_outputs(288)) or (layer0_outputs(804)));
    outputs(1106) <= layer0_outputs(7067);
    outputs(1107) <= not(layer0_outputs(6176));
    outputs(1108) <= layer0_outputs(6417);
    outputs(1109) <= (layer0_outputs(5675)) and (layer0_outputs(3596));
    outputs(1110) <= layer0_outputs(1681);
    outputs(1111) <= (layer0_outputs(6225)) xor (layer0_outputs(2702));
    outputs(1112) <= layer0_outputs(5857);
    outputs(1113) <= not(layer0_outputs(1062));
    outputs(1114) <= (layer0_outputs(2791)) and not (layer0_outputs(4706));
    outputs(1115) <= (layer0_outputs(1713)) and (layer0_outputs(7491));
    outputs(1116) <= (layer0_outputs(881)) and (layer0_outputs(7496));
    outputs(1117) <= layer0_outputs(7596);
    outputs(1118) <= (layer0_outputs(2933)) xor (layer0_outputs(7010));
    outputs(1119) <= layer0_outputs(108);
    outputs(1120) <= (layer0_outputs(4100)) and (layer0_outputs(2199));
    outputs(1121) <= not((layer0_outputs(3993)) or (layer0_outputs(5307)));
    outputs(1122) <= (layer0_outputs(3587)) and not (layer0_outputs(498));
    outputs(1123) <= layer0_outputs(1179);
    outputs(1124) <= not(layer0_outputs(5414));
    outputs(1125) <= not((layer0_outputs(2087)) or (layer0_outputs(1496)));
    outputs(1126) <= not((layer0_outputs(2529)) xor (layer0_outputs(1060)));
    outputs(1127) <= (layer0_outputs(4180)) and not (layer0_outputs(2369));
    outputs(1128) <= (layer0_outputs(6554)) and not (layer0_outputs(2026));
    outputs(1129) <= not((layer0_outputs(3795)) xor (layer0_outputs(6904)));
    outputs(1130) <= (layer0_outputs(7225)) and not (layer0_outputs(7504));
    outputs(1131) <= (layer0_outputs(4)) and not (layer0_outputs(633));
    outputs(1132) <= (layer0_outputs(467)) and not (layer0_outputs(4085));
    outputs(1133) <= (layer0_outputs(7375)) and not (layer0_outputs(4905));
    outputs(1134) <= (layer0_outputs(6782)) and not (layer0_outputs(2329));
    outputs(1135) <= not((layer0_outputs(1160)) or (layer0_outputs(3445)));
    outputs(1136) <= not(layer0_outputs(7092));
    outputs(1137) <= not((layer0_outputs(2703)) or (layer0_outputs(1793)));
    outputs(1138) <= (layer0_outputs(2977)) and not (layer0_outputs(6872));
    outputs(1139) <= not((layer0_outputs(3034)) and (layer0_outputs(5292)));
    outputs(1140) <= not((layer0_outputs(411)) or (layer0_outputs(1768)));
    outputs(1141) <= '0';
    outputs(1142) <= (layer0_outputs(5828)) and not (layer0_outputs(1355));
    outputs(1143) <= (layer0_outputs(486)) and not (layer0_outputs(2562));
    outputs(1144) <= (layer0_outputs(2437)) and not (layer0_outputs(7075));
    outputs(1145) <= (layer0_outputs(628)) and not (layer0_outputs(5974));
    outputs(1146) <= not((layer0_outputs(5509)) or (layer0_outputs(2150)));
    outputs(1147) <= layer0_outputs(434);
    outputs(1148) <= '0';
    outputs(1149) <= not(layer0_outputs(6240));
    outputs(1150) <= '0';
    outputs(1151) <= not((layer0_outputs(7305)) xor (layer0_outputs(6340)));
    outputs(1152) <= not((layer0_outputs(6481)) xor (layer0_outputs(5706)));
    outputs(1153) <= not(layer0_outputs(7052)) or (layer0_outputs(3420));
    outputs(1154) <= not((layer0_outputs(4387)) or (layer0_outputs(5847)));
    outputs(1155) <= not(layer0_outputs(3392));
    outputs(1156) <= not((layer0_outputs(408)) xor (layer0_outputs(7462)));
    outputs(1157) <= (layer0_outputs(4031)) and not (layer0_outputs(5507));
    outputs(1158) <= '0';
    outputs(1159) <= not(layer0_outputs(2606));
    outputs(1160) <= (layer0_outputs(7188)) and not (layer0_outputs(189));
    outputs(1161) <= (layer0_outputs(421)) and not (layer0_outputs(7540));
    outputs(1162) <= not(layer0_outputs(2604));
    outputs(1163) <= not(layer0_outputs(3106));
    outputs(1164) <= (layer0_outputs(1846)) and (layer0_outputs(4594));
    outputs(1165) <= (layer0_outputs(3674)) and not (layer0_outputs(812));
    outputs(1166) <= (layer0_outputs(1387)) and not (layer0_outputs(2023));
    outputs(1167) <= not(layer0_outputs(5398));
    outputs(1168) <= not((layer0_outputs(1765)) or (layer0_outputs(6355)));
    outputs(1169) <= not((layer0_outputs(5665)) or (layer0_outputs(7447)));
    outputs(1170) <= not(layer0_outputs(1187));
    outputs(1171) <= layer0_outputs(7022);
    outputs(1172) <= not((layer0_outputs(1559)) or (layer0_outputs(442)));
    outputs(1173) <= (layer0_outputs(6431)) and not (layer0_outputs(4782));
    outputs(1174) <= layer0_outputs(5959);
    outputs(1175) <= (layer0_outputs(5575)) and not (layer0_outputs(6631));
    outputs(1176) <= (layer0_outputs(3403)) and (layer0_outputs(6592));
    outputs(1177) <= layer0_outputs(3528);
    outputs(1178) <= (layer0_outputs(2080)) and not (layer0_outputs(2785));
    outputs(1179) <= not(layer0_outputs(329));
    outputs(1180) <= not((layer0_outputs(206)) xor (layer0_outputs(868)));
    outputs(1181) <= layer0_outputs(7169);
    outputs(1182) <= (layer0_outputs(947)) and (layer0_outputs(6519));
    outputs(1183) <= not(layer0_outputs(6574));
    outputs(1184) <= (layer0_outputs(23)) and not (layer0_outputs(3648));
    outputs(1185) <= (layer0_outputs(2456)) or (layer0_outputs(2311));
    outputs(1186) <= not(layer0_outputs(1286));
    outputs(1187) <= (layer0_outputs(3939)) and not (layer0_outputs(5678));
    outputs(1188) <= not(layer0_outputs(1013));
    outputs(1189) <= not((layer0_outputs(3715)) or (layer0_outputs(6104)));
    outputs(1190) <= (layer0_outputs(3990)) xor (layer0_outputs(3793));
    outputs(1191) <= (layer0_outputs(5870)) and not (layer0_outputs(6533));
    outputs(1192) <= layer0_outputs(5641);
    outputs(1193) <= layer0_outputs(2991);
    outputs(1194) <= not(layer0_outputs(5527));
    outputs(1195) <= '0';
    outputs(1196) <= not((layer0_outputs(4516)) or (layer0_outputs(2630)));
    outputs(1197) <= not(layer0_outputs(2537));
    outputs(1198) <= (layer0_outputs(1384)) xor (layer0_outputs(2270));
    outputs(1199) <= (layer0_outputs(4531)) and (layer0_outputs(6815));
    outputs(1200) <= layer0_outputs(3156);
    outputs(1201) <= (layer0_outputs(287)) xor (layer0_outputs(5303));
    outputs(1202) <= not(layer0_outputs(4236));
    outputs(1203) <= not((layer0_outputs(7630)) and (layer0_outputs(2570)));
    outputs(1204) <= (layer0_outputs(1848)) and not (layer0_outputs(4680));
    outputs(1205) <= not((layer0_outputs(5026)) xor (layer0_outputs(952)));
    outputs(1206) <= not(layer0_outputs(5995));
    outputs(1207) <= not(layer0_outputs(3878));
    outputs(1208) <= (layer0_outputs(4188)) and not (layer0_outputs(6624));
    outputs(1209) <= not(layer0_outputs(2277));
    outputs(1210) <= layer0_outputs(6379);
    outputs(1211) <= (layer0_outputs(5801)) and not (layer0_outputs(5805));
    outputs(1212) <= (layer0_outputs(661)) and not (layer0_outputs(2382));
    outputs(1213) <= layer0_outputs(4288);
    outputs(1214) <= layer0_outputs(2572);
    outputs(1215) <= not(layer0_outputs(5838));
    outputs(1216) <= layer0_outputs(2290);
    outputs(1217) <= (layer0_outputs(537)) and (layer0_outputs(726));
    outputs(1218) <= (layer0_outputs(303)) xor (layer0_outputs(6345));
    outputs(1219) <= (layer0_outputs(58)) and not (layer0_outputs(999));
    outputs(1220) <= (layer0_outputs(3197)) and (layer0_outputs(2584));
    outputs(1221) <= not(layer0_outputs(2453));
    outputs(1222) <= (layer0_outputs(3931)) and not (layer0_outputs(4622));
    outputs(1223) <= layer0_outputs(1606);
    outputs(1224) <= (layer0_outputs(7276)) and not (layer0_outputs(4693));
    outputs(1225) <= (layer0_outputs(3957)) xor (layer0_outputs(7231));
    outputs(1226) <= not(layer0_outputs(5319));
    outputs(1227) <= not(layer0_outputs(1874));
    outputs(1228) <= (layer0_outputs(1904)) xor (layer0_outputs(2339));
    outputs(1229) <= not(layer0_outputs(7394));
    outputs(1230) <= not(layer0_outputs(4109));
    outputs(1231) <= (layer0_outputs(1529)) and not (layer0_outputs(2896));
    outputs(1232) <= not(layer0_outputs(4644));
    outputs(1233) <= layer0_outputs(2160);
    outputs(1234) <= not((layer0_outputs(5981)) or (layer0_outputs(3273)));
    outputs(1235) <= (layer0_outputs(3405)) and not (layer0_outputs(3747));
    outputs(1236) <= (layer0_outputs(1742)) and not (layer0_outputs(7138));
    outputs(1237) <= (layer0_outputs(1758)) and not (layer0_outputs(5182));
    outputs(1238) <= layer0_outputs(4374);
    outputs(1239) <= not(layer0_outputs(1386));
    outputs(1240) <= not((layer0_outputs(6479)) xor (layer0_outputs(1087)));
    outputs(1241) <= (layer0_outputs(5284)) and not (layer0_outputs(2508));
    outputs(1242) <= (layer0_outputs(521)) and (layer0_outputs(3203));
    outputs(1243) <= not((layer0_outputs(4499)) or (layer0_outputs(796)));
    outputs(1244) <= (layer0_outputs(669)) and not (layer0_outputs(6565));
    outputs(1245) <= not(layer0_outputs(964));
    outputs(1246) <= not((layer0_outputs(7298)) or (layer0_outputs(5472)));
    outputs(1247) <= (layer0_outputs(7603)) and not (layer0_outputs(731));
    outputs(1248) <= (layer0_outputs(2064)) and (layer0_outputs(6831));
    outputs(1249) <= (layer0_outputs(3438)) xor (layer0_outputs(4592));
    outputs(1250) <= (layer0_outputs(621)) and not (layer0_outputs(6413));
    outputs(1251) <= (layer0_outputs(3477)) and (layer0_outputs(2521));
    outputs(1252) <= not((layer0_outputs(5599)) xor (layer0_outputs(4554)));
    outputs(1253) <= (layer0_outputs(7608)) xor (layer0_outputs(355));
    outputs(1254) <= not((layer0_outputs(358)) or (layer0_outputs(6439)));
    outputs(1255) <= not((layer0_outputs(5917)) or (layer0_outputs(6707)));
    outputs(1256) <= layer0_outputs(7551);
    outputs(1257) <= not(layer0_outputs(2210));
    outputs(1258) <= not((layer0_outputs(2816)) xor (layer0_outputs(6885)));
    outputs(1259) <= not(layer0_outputs(5810));
    outputs(1260) <= layer0_outputs(459);
    outputs(1261) <= not(layer0_outputs(6415));
    outputs(1262) <= (layer0_outputs(3731)) xor (layer0_outputs(683));
    outputs(1263) <= (layer0_outputs(4602)) xor (layer0_outputs(954));
    outputs(1264) <= (layer0_outputs(709)) and not (layer0_outputs(5251));
    outputs(1265) <= not(layer0_outputs(6609));
    outputs(1266) <= layer0_outputs(5713);
    outputs(1267) <= (layer0_outputs(5190)) and not (layer0_outputs(1707));
    outputs(1268) <= not(layer0_outputs(6040)) or (layer0_outputs(1926));
    outputs(1269) <= (layer0_outputs(5225)) and not (layer0_outputs(4028));
    outputs(1270) <= (layer0_outputs(7335)) xor (layer0_outputs(5476));
    outputs(1271) <= (layer0_outputs(3053)) xor (layer0_outputs(1496));
    outputs(1272) <= (layer0_outputs(3869)) and not (layer0_outputs(5105));
    outputs(1273) <= layer0_outputs(4063);
    outputs(1274) <= not((layer0_outputs(6920)) and (layer0_outputs(3862)));
    outputs(1275) <= (layer0_outputs(5386)) and not (layer0_outputs(1817));
    outputs(1276) <= (layer0_outputs(2602)) and not (layer0_outputs(5778));
    outputs(1277) <= (layer0_outputs(715)) xor (layer0_outputs(7290));
    outputs(1278) <= (layer0_outputs(5322)) and not (layer0_outputs(4017));
    outputs(1279) <= not((layer0_outputs(4156)) xor (layer0_outputs(2018)));
    outputs(1280) <= not(layer0_outputs(4573));
    outputs(1281) <= (layer0_outputs(6233)) and (layer0_outputs(7315));
    outputs(1282) <= not((layer0_outputs(5270)) xor (layer0_outputs(6061)));
    outputs(1283) <= (layer0_outputs(821)) and (layer0_outputs(3756));
    outputs(1284) <= layer0_outputs(4162);
    outputs(1285) <= (layer0_outputs(428)) xor (layer0_outputs(6004));
    outputs(1286) <= not(layer0_outputs(1324));
    outputs(1287) <= (layer0_outputs(4441)) xor (layer0_outputs(1436));
    outputs(1288) <= not((layer0_outputs(3265)) or (layer0_outputs(3480)));
    outputs(1289) <= (layer0_outputs(874)) xor (layer0_outputs(2327));
    outputs(1290) <= layer0_outputs(5673);
    outputs(1291) <= not((layer0_outputs(5204)) or (layer0_outputs(1240)));
    outputs(1292) <= (layer0_outputs(6561)) and not (layer0_outputs(6094));
    outputs(1293) <= not(layer0_outputs(126));
    outputs(1294) <= (layer0_outputs(6774)) and (layer0_outputs(6556));
    outputs(1295) <= (layer0_outputs(5711)) and not (layer0_outputs(5694));
    outputs(1296) <= (layer0_outputs(2204)) xor (layer0_outputs(6252));
    outputs(1297) <= layer0_outputs(4211);
    outputs(1298) <= '0';
    outputs(1299) <= (layer0_outputs(1432)) and (layer0_outputs(3990));
    outputs(1300) <= not(layer0_outputs(1520));
    outputs(1301) <= (layer0_outputs(971)) xor (layer0_outputs(879));
    outputs(1302) <= not((layer0_outputs(6505)) or (layer0_outputs(2972)));
    outputs(1303) <= (layer0_outputs(3270)) xor (layer0_outputs(5501));
    outputs(1304) <= (layer0_outputs(1406)) xor (layer0_outputs(5910));
    outputs(1305) <= (layer0_outputs(7304)) and (layer0_outputs(4948));
    outputs(1306) <= (layer0_outputs(4094)) xor (layer0_outputs(605));
    outputs(1307) <= '0';
    outputs(1308) <= not((layer0_outputs(3022)) xor (layer0_outputs(4952)));
    outputs(1309) <= (layer0_outputs(7019)) and not (layer0_outputs(2898));
    outputs(1310) <= not((layer0_outputs(7439)) or (layer0_outputs(4964)));
    outputs(1311) <= (layer0_outputs(4809)) and (layer0_outputs(2550));
    outputs(1312) <= not((layer0_outputs(5100)) and (layer0_outputs(1197)));
    outputs(1313) <= layer0_outputs(2376);
    outputs(1314) <= (layer0_outputs(6941)) xor (layer0_outputs(492));
    outputs(1315) <= not((layer0_outputs(6021)) or (layer0_outputs(3697)));
    outputs(1316) <= layer0_outputs(5453);
    outputs(1317) <= (layer0_outputs(3113)) and not (layer0_outputs(2708));
    outputs(1318) <= (layer0_outputs(7349)) and (layer0_outputs(4555));
    outputs(1319) <= (layer0_outputs(6824)) and not (layer0_outputs(4339));
    outputs(1320) <= not((layer0_outputs(1639)) or (layer0_outputs(1635)));
    outputs(1321) <= layer0_outputs(1351);
    outputs(1322) <= layer0_outputs(2849);
    outputs(1323) <= layer0_outputs(4903);
    outputs(1324) <= not(layer0_outputs(4346));
    outputs(1325) <= not((layer0_outputs(264)) xor (layer0_outputs(3555)));
    outputs(1326) <= not((layer0_outputs(6476)) or (layer0_outputs(4179)));
    outputs(1327) <= (layer0_outputs(3875)) and not (layer0_outputs(1618));
    outputs(1328) <= (layer0_outputs(5701)) and not (layer0_outputs(6060));
    outputs(1329) <= (layer0_outputs(4239)) and (layer0_outputs(2394));
    outputs(1330) <= not((layer0_outputs(7507)) or (layer0_outputs(824)));
    outputs(1331) <= (layer0_outputs(2041)) and not (layer0_outputs(1061));
    outputs(1332) <= not(layer0_outputs(917));
    outputs(1333) <= not((layer0_outputs(2675)) xor (layer0_outputs(3616)));
    outputs(1334) <= (layer0_outputs(3319)) and not (layer0_outputs(552));
    outputs(1335) <= (layer0_outputs(595)) and not (layer0_outputs(7029));
    outputs(1336) <= not((layer0_outputs(4837)) or (layer0_outputs(3884)));
    outputs(1337) <= not(layer0_outputs(3041));
    outputs(1338) <= layer0_outputs(6125);
    outputs(1339) <= (layer0_outputs(7036)) and not (layer0_outputs(447));
    outputs(1340) <= not((layer0_outputs(4869)) or (layer0_outputs(4196)));
    outputs(1341) <= layer0_outputs(5329);
    outputs(1342) <= (layer0_outputs(3899)) and not (layer0_outputs(2927));
    outputs(1343) <= not(layer0_outputs(4128));
    outputs(1344) <= not(layer0_outputs(4813));
    outputs(1345) <= layer0_outputs(6792);
    outputs(1346) <= layer0_outputs(4010);
    outputs(1347) <= (layer0_outputs(5186)) and not (layer0_outputs(3466));
    outputs(1348) <= not((layer0_outputs(1114)) xor (layer0_outputs(6626)));
    outputs(1349) <= not((layer0_outputs(6959)) xor (layer0_outputs(3425)));
    outputs(1350) <= not((layer0_outputs(2930)) or (layer0_outputs(601)));
    outputs(1351) <= not((layer0_outputs(1002)) or (layer0_outputs(249)));
    outputs(1352) <= layer0_outputs(6811);
    outputs(1353) <= (layer0_outputs(1226)) and (layer0_outputs(1029));
    outputs(1354) <= layer0_outputs(6797);
    outputs(1355) <= (layer0_outputs(3510)) and (layer0_outputs(2306));
    outputs(1356) <= (layer0_outputs(5498)) and not (layer0_outputs(606));
    outputs(1357) <= not((layer0_outputs(6889)) or (layer0_outputs(7473)));
    outputs(1358) <= not(layer0_outputs(1436));
    outputs(1359) <= (layer0_outputs(785)) and not (layer0_outputs(1188));
    outputs(1360) <= (layer0_outputs(384)) and not (layer0_outputs(5483));
    outputs(1361) <= not(layer0_outputs(3631));
    outputs(1362) <= not(layer0_outputs(5056));
    outputs(1363) <= '0';
    outputs(1364) <= (layer0_outputs(497)) and (layer0_outputs(6477));
    outputs(1365) <= not((layer0_outputs(2856)) or (layer0_outputs(7523)));
    outputs(1366) <= not((layer0_outputs(3788)) xor (layer0_outputs(936)));
    outputs(1367) <= (layer0_outputs(6330)) xor (layer0_outputs(3754));
    outputs(1368) <= layer0_outputs(7449);
    outputs(1369) <= not((layer0_outputs(6041)) xor (layer0_outputs(5084)));
    outputs(1370) <= (layer0_outputs(3123)) and (layer0_outputs(433));
    outputs(1371) <= not(layer0_outputs(6838));
    outputs(1372) <= not(layer0_outputs(2682));
    outputs(1373) <= not(layer0_outputs(2619));
    outputs(1374) <= (layer0_outputs(7440)) xor (layer0_outputs(4432));
    outputs(1375) <= not((layer0_outputs(1336)) or (layer0_outputs(1263)));
    outputs(1376) <= (layer0_outputs(1281)) and (layer0_outputs(6242));
    outputs(1377) <= not(layer0_outputs(6908)) or (layer0_outputs(1714));
    outputs(1378) <= not((layer0_outputs(3317)) xor (layer0_outputs(545)));
    outputs(1379) <= not(layer0_outputs(2381));
    outputs(1380) <= (layer0_outputs(2183)) and not (layer0_outputs(998));
    outputs(1381) <= '0';
    outputs(1382) <= layer0_outputs(6553);
    outputs(1383) <= (layer0_outputs(4735)) and (layer0_outputs(4608));
    outputs(1384) <= (layer0_outputs(7508)) and (layer0_outputs(4303));
    outputs(1385) <= not((layer0_outputs(1925)) xor (layer0_outputs(3595)));
    outputs(1386) <= (layer0_outputs(1976)) xor (layer0_outputs(1899));
    outputs(1387) <= '0';
    outputs(1388) <= (layer0_outputs(5497)) and not (layer0_outputs(6287));
    outputs(1389) <= not(layer0_outputs(1117));
    outputs(1390) <= not((layer0_outputs(1702)) or (layer0_outputs(3450)));
    outputs(1391) <= (layer0_outputs(5916)) and not (layer0_outputs(730));
    outputs(1392) <= not((layer0_outputs(1682)) or (layer0_outputs(868)));
    outputs(1393) <= (layer0_outputs(2469)) and (layer0_outputs(7568));
    outputs(1394) <= (layer0_outputs(7241)) and not (layer0_outputs(2198));
    outputs(1395) <= layer0_outputs(6571);
    outputs(1396) <= not(layer0_outputs(5341));
    outputs(1397) <= not(layer0_outputs(6397));
    outputs(1398) <= (layer0_outputs(4383)) and not (layer0_outputs(5478));
    outputs(1399) <= layer0_outputs(86);
    outputs(1400) <= (layer0_outputs(6708)) and (layer0_outputs(2793));
    outputs(1401) <= not(layer0_outputs(2383));
    outputs(1402) <= layer0_outputs(3113);
    outputs(1403) <= not((layer0_outputs(4568)) or (layer0_outputs(7661)));
    outputs(1404) <= not((layer0_outputs(3908)) or (layer0_outputs(4616)));
    outputs(1405) <= layer0_outputs(2700);
    outputs(1406) <= (layer0_outputs(677)) xor (layer0_outputs(4570));
    outputs(1407) <= (layer0_outputs(7367)) and (layer0_outputs(3529));
    outputs(1408) <= layer0_outputs(5034);
    outputs(1409) <= (layer0_outputs(7324)) and (layer0_outputs(2753));
    outputs(1410) <= not(layer0_outputs(3486));
    outputs(1411) <= (layer0_outputs(6453)) and not (layer0_outputs(6412));
    outputs(1412) <= (layer0_outputs(4954)) and (layer0_outputs(3449));
    outputs(1413) <= layer0_outputs(1564);
    outputs(1414) <= not((layer0_outputs(449)) xor (layer0_outputs(120)));
    outputs(1415) <= layer0_outputs(4274);
    outputs(1416) <= not(layer0_outputs(409));
    outputs(1417) <= (layer0_outputs(96)) and (layer0_outputs(4354));
    outputs(1418) <= not(layer0_outputs(6895));
    outputs(1419) <= not((layer0_outputs(3172)) xor (layer0_outputs(7549)));
    outputs(1420) <= not((layer0_outputs(6789)) or (layer0_outputs(5905)));
    outputs(1421) <= not((layer0_outputs(6517)) or (layer0_outputs(3803)));
    outputs(1422) <= (layer0_outputs(2242)) and not (layer0_outputs(5656));
    outputs(1423) <= not(layer0_outputs(4878));
    outputs(1424) <= not((layer0_outputs(625)) or (layer0_outputs(6186)));
    outputs(1425) <= layer0_outputs(6654);
    outputs(1426) <= (layer0_outputs(7611)) and (layer0_outputs(3667));
    outputs(1427) <= not(layer0_outputs(7620));
    outputs(1428) <= not((layer0_outputs(6279)) or (layer0_outputs(1805)));
    outputs(1429) <= (layer0_outputs(4932)) and not (layer0_outputs(5311));
    outputs(1430) <= (layer0_outputs(1199)) and not (layer0_outputs(70));
    outputs(1431) <= not((layer0_outputs(2515)) xor (layer0_outputs(7666)));
    outputs(1432) <= (layer0_outputs(2908)) and not (layer0_outputs(1871));
    outputs(1433) <= layer0_outputs(6087);
    outputs(1434) <= not((layer0_outputs(7136)) xor (layer0_outputs(747)));
    outputs(1435) <= not((layer0_outputs(4823)) xor (layer0_outputs(3448)));
    outputs(1436) <= not(layer0_outputs(3111));
    outputs(1437) <= (layer0_outputs(6494)) xor (layer0_outputs(7099));
    outputs(1438) <= (layer0_outputs(101)) and (layer0_outputs(4610));
    outputs(1439) <= not((layer0_outputs(7230)) xor (layer0_outputs(137)));
    outputs(1440) <= layer0_outputs(2238);
    outputs(1441) <= (layer0_outputs(2688)) xor (layer0_outputs(1888));
    outputs(1442) <= layer0_outputs(4030);
    outputs(1443) <= layer0_outputs(4844);
    outputs(1444) <= (layer0_outputs(6337)) and (layer0_outputs(3823));
    outputs(1445) <= not(layer0_outputs(6659)) or (layer0_outputs(7537));
    outputs(1446) <= (layer0_outputs(2588)) and not (layer0_outputs(3440));
    outputs(1447) <= (layer0_outputs(5736)) and not (layer0_outputs(1529));
    outputs(1448) <= (layer0_outputs(2119)) and (layer0_outputs(7154));
    outputs(1449) <= (layer0_outputs(4561)) xor (layer0_outputs(2389));
    outputs(1450) <= (layer0_outputs(2815)) and (layer0_outputs(6393));
    outputs(1451) <= layer0_outputs(148);
    outputs(1452) <= not(layer0_outputs(3640));
    outputs(1453) <= (layer0_outputs(5058)) xor (layer0_outputs(6458));
    outputs(1454) <= not(layer0_outputs(5612));
    outputs(1455) <= (layer0_outputs(145)) and not (layer0_outputs(4246));
    outputs(1456) <= (layer0_outputs(6491)) and (layer0_outputs(5570));
    outputs(1457) <= layer0_outputs(4325);
    outputs(1458) <= (layer0_outputs(1299)) xor (layer0_outputs(6235));
    outputs(1459) <= '0';
    outputs(1460) <= (layer0_outputs(664)) and not (layer0_outputs(613));
    outputs(1461) <= not(layer0_outputs(1845));
    outputs(1462) <= (layer0_outputs(2877)) and (layer0_outputs(6038));
    outputs(1463) <= not((layer0_outputs(4740)) or (layer0_outputs(4725)));
    outputs(1464) <= layer0_outputs(2404);
    outputs(1465) <= layer0_outputs(4816);
    outputs(1466) <= (layer0_outputs(4467)) and (layer0_outputs(6127));
    outputs(1467) <= (layer0_outputs(1708)) and not (layer0_outputs(4155));
    outputs(1468) <= (layer0_outputs(2262)) and (layer0_outputs(982));
    outputs(1469) <= (layer0_outputs(2637)) xor (layer0_outputs(6359));
    outputs(1470) <= (layer0_outputs(2350)) and not (layer0_outputs(680));
    outputs(1471) <= not((layer0_outputs(2487)) or (layer0_outputs(3668)));
    outputs(1472) <= (layer0_outputs(3412)) xor (layer0_outputs(125));
    outputs(1473) <= not((layer0_outputs(44)) or (layer0_outputs(1013)));
    outputs(1474) <= layer0_outputs(1582);
    outputs(1475) <= (layer0_outputs(1494)) xor (layer0_outputs(6046));
    outputs(1476) <= not((layer0_outputs(2099)) or (layer0_outputs(7335)));
    outputs(1477) <= (layer0_outputs(3604)) and not (layer0_outputs(6186));
    outputs(1478) <= not(layer0_outputs(2156));
    outputs(1479) <= not((layer0_outputs(883)) or (layer0_outputs(1570)));
    outputs(1480) <= not((layer0_outputs(7299)) or (layer0_outputs(4631)));
    outputs(1481) <= not((layer0_outputs(3814)) or (layer0_outputs(2058)));
    outputs(1482) <= layer0_outputs(2814);
    outputs(1483) <= (layer0_outputs(4552)) and not (layer0_outputs(4629));
    outputs(1484) <= not(layer0_outputs(5541));
    outputs(1485) <= not(layer0_outputs(2580));
    outputs(1486) <= not(layer0_outputs(2094));
    outputs(1487) <= not((layer0_outputs(3098)) or (layer0_outputs(6711)));
    outputs(1488) <= (layer0_outputs(5220)) and (layer0_outputs(3406));
    outputs(1489) <= not((layer0_outputs(243)) xor (layer0_outputs(5047)));
    outputs(1490) <= not((layer0_outputs(1130)) or (layer0_outputs(2703)));
    outputs(1491) <= (layer0_outputs(4520)) and (layer0_outputs(1172));
    outputs(1492) <= (layer0_outputs(3062)) and (layer0_outputs(5901));
    outputs(1493) <= layer0_outputs(4699);
    outputs(1494) <= layer0_outputs(1973);
    outputs(1495) <= (layer0_outputs(5206)) and (layer0_outputs(724));
    outputs(1496) <= layer0_outputs(4334);
    outputs(1497) <= layer0_outputs(3379);
    outputs(1498) <= layer0_outputs(711);
    outputs(1499) <= (layer0_outputs(5428)) and (layer0_outputs(7619));
    outputs(1500) <= not(layer0_outputs(2911));
    outputs(1501) <= (layer0_outputs(7233)) and not (layer0_outputs(1766));
    outputs(1502) <= (layer0_outputs(5526)) and (layer0_outputs(1317));
    outputs(1503) <= (layer0_outputs(653)) and (layer0_outputs(1853));
    outputs(1504) <= (layer0_outputs(7614)) and not (layer0_outputs(4998));
    outputs(1505) <= (layer0_outputs(522)) xor (layer0_outputs(582));
    outputs(1506) <= not((layer0_outputs(398)) or (layer0_outputs(5545)));
    outputs(1507) <= not(layer0_outputs(1475));
    outputs(1508) <= (layer0_outputs(5553)) and not (layer0_outputs(6005));
    outputs(1509) <= '0';
    outputs(1510) <= not((layer0_outputs(3287)) or (layer0_outputs(1361)));
    outputs(1511) <= (layer0_outputs(7656)) xor (layer0_outputs(6030));
    outputs(1512) <= layer0_outputs(1936);
    outputs(1513) <= not(layer0_outputs(3597));
    outputs(1514) <= not(layer0_outputs(1628));
    outputs(1515) <= layer0_outputs(5112);
    outputs(1516) <= (layer0_outputs(3986)) and (layer0_outputs(1864));
    outputs(1517) <= layer0_outputs(6887);
    outputs(1518) <= (layer0_outputs(6988)) and not (layer0_outputs(2697));
    outputs(1519) <= (layer0_outputs(7469)) and not (layer0_outputs(445));
    outputs(1520) <= (layer0_outputs(4138)) and (layer0_outputs(5023));
    outputs(1521) <= not(layer0_outputs(7115));
    outputs(1522) <= not(layer0_outputs(4244));
    outputs(1523) <= not((layer0_outputs(5880)) or (layer0_outputs(4206)));
    outputs(1524) <= not((layer0_outputs(3983)) or (layer0_outputs(4843)));
    outputs(1525) <= not((layer0_outputs(4168)) and (layer0_outputs(5279)));
    outputs(1526) <= (layer0_outputs(2406)) and not (layer0_outputs(6656));
    outputs(1527) <= not(layer0_outputs(2540));
    outputs(1528) <= (layer0_outputs(3099)) xor (layer0_outputs(6500));
    outputs(1529) <= (layer0_outputs(2599)) and (layer0_outputs(5188));
    outputs(1530) <= layer0_outputs(2962);
    outputs(1531) <= (layer0_outputs(4511)) and not (layer0_outputs(4043));
    outputs(1532) <= (layer0_outputs(4064)) xor (layer0_outputs(2535));
    outputs(1533) <= not((layer0_outputs(2728)) or (layer0_outputs(1805)));
    outputs(1534) <= (layer0_outputs(3212)) and not (layer0_outputs(289));
    outputs(1535) <= not(layer0_outputs(7012));
    outputs(1536) <= not(layer0_outputs(3152));
    outputs(1537) <= (layer0_outputs(1525)) xor (layer0_outputs(2657));
    outputs(1538) <= layer0_outputs(3030);
    outputs(1539) <= (layer0_outputs(2389)) xor (layer0_outputs(3833));
    outputs(1540) <= layer0_outputs(3261);
    outputs(1541) <= not((layer0_outputs(4347)) and (layer0_outputs(5856)));
    outputs(1542) <= not(layer0_outputs(7385));
    outputs(1543) <= (layer0_outputs(7329)) xor (layer0_outputs(5039));
    outputs(1544) <= not(layer0_outputs(479)) or (layer0_outputs(3614));
    outputs(1545) <= not((layer0_outputs(3572)) and (layer0_outputs(3736)));
    outputs(1546) <= not((layer0_outputs(361)) and (layer0_outputs(7584)));
    outputs(1547) <= layer0_outputs(3600);
    outputs(1548) <= not(layer0_outputs(3056));
    outputs(1549) <= (layer0_outputs(3695)) and not (layer0_outputs(7158));
    outputs(1550) <= (layer0_outputs(3358)) and not (layer0_outputs(6094));
    outputs(1551) <= layer0_outputs(3338);
    outputs(1552) <= layer0_outputs(2420);
    outputs(1553) <= layer0_outputs(2174);
    outputs(1554) <= not((layer0_outputs(2817)) xor (layer0_outputs(6346)));
    outputs(1555) <= not(layer0_outputs(60));
    outputs(1556) <= layer0_outputs(4773);
    outputs(1557) <= not(layer0_outputs(3714));
    outputs(1558) <= (layer0_outputs(1661)) xor (layer0_outputs(4178));
    outputs(1559) <= not((layer0_outputs(4475)) xor (layer0_outputs(2759)));
    outputs(1560) <= not(layer0_outputs(4523));
    outputs(1561) <= (layer0_outputs(2060)) or (layer0_outputs(4048));
    outputs(1562) <= not(layer0_outputs(6338));
    outputs(1563) <= (layer0_outputs(3342)) xor (layer0_outputs(5886));
    outputs(1564) <= not(layer0_outputs(5137));
    outputs(1565) <= layer0_outputs(2027);
    outputs(1566) <= not(layer0_outputs(4691));
    outputs(1567) <= not((layer0_outputs(4714)) xor (layer0_outputs(2092)));
    outputs(1568) <= not(layer0_outputs(7256));
    outputs(1569) <= not(layer0_outputs(733)) or (layer0_outputs(3622));
    outputs(1570) <= not(layer0_outputs(2595));
    outputs(1571) <= not(layer0_outputs(3405)) or (layer0_outputs(517));
    outputs(1572) <= layer0_outputs(5620);
    outputs(1573) <= layer0_outputs(305);
    outputs(1574) <= not((layer0_outputs(116)) xor (layer0_outputs(7186)));
    outputs(1575) <= layer0_outputs(5800);
    outputs(1576) <= layer0_outputs(2233);
    outputs(1577) <= layer0_outputs(3920);
    outputs(1578) <= layer0_outputs(778);
    outputs(1579) <= layer0_outputs(6373);
    outputs(1580) <= not(layer0_outputs(2403)) or (layer0_outputs(9));
    outputs(1581) <= (layer0_outputs(2111)) xor (layer0_outputs(3986));
    outputs(1582) <= not(layer0_outputs(4971));
    outputs(1583) <= layer0_outputs(616);
    outputs(1584) <= not(layer0_outputs(6970)) or (layer0_outputs(6152));
    outputs(1585) <= layer0_outputs(7203);
    outputs(1586) <= not(layer0_outputs(3473));
    outputs(1587) <= not(layer0_outputs(5723)) or (layer0_outputs(1250));
    outputs(1588) <= not(layer0_outputs(3050));
    outputs(1589) <= not((layer0_outputs(3590)) xor (layer0_outputs(1197)));
    outputs(1590) <= layer0_outputs(6976);
    outputs(1591) <= (layer0_outputs(1660)) xor (layer0_outputs(2414));
    outputs(1592) <= not((layer0_outputs(1431)) and (layer0_outputs(2516)));
    outputs(1593) <= not((layer0_outputs(1352)) and (layer0_outputs(3022)));
    outputs(1594) <= not((layer0_outputs(6678)) and (layer0_outputs(5951)));
    outputs(1595) <= not((layer0_outputs(1763)) and (layer0_outputs(1974)));
    outputs(1596) <= not(layer0_outputs(6452)) or (layer0_outputs(6604));
    outputs(1597) <= layer0_outputs(773);
    outputs(1598) <= (layer0_outputs(5267)) xor (layer0_outputs(6907));
    outputs(1599) <= not(layer0_outputs(5156));
    outputs(1600) <= (layer0_outputs(2414)) and not (layer0_outputs(5961));
    outputs(1601) <= not(layer0_outputs(820));
    outputs(1602) <= not((layer0_outputs(375)) and (layer0_outputs(3282)));
    outputs(1603) <= (layer0_outputs(6647)) xor (layer0_outputs(1905));
    outputs(1604) <= (layer0_outputs(2997)) and not (layer0_outputs(2066));
    outputs(1605) <= not(layer0_outputs(4412)) or (layer0_outputs(1155));
    outputs(1606) <= layer0_outputs(6414);
    outputs(1607) <= not((layer0_outputs(583)) xor (layer0_outputs(4560)));
    outputs(1608) <= layer0_outputs(6723);
    outputs(1609) <= not((layer0_outputs(7157)) and (layer0_outputs(5293)));
    outputs(1610) <= not(layer0_outputs(3662));
    outputs(1611) <= not((layer0_outputs(2704)) xor (layer0_outputs(987)));
    outputs(1612) <= not((layer0_outputs(1280)) and (layer0_outputs(1209)));
    outputs(1613) <= not((layer0_outputs(3763)) and (layer0_outputs(4765)));
    outputs(1614) <= not((layer0_outputs(5740)) xor (layer0_outputs(4507)));
    outputs(1615) <= not((layer0_outputs(4619)) xor (layer0_outputs(1425)));
    outputs(1616) <= not(layer0_outputs(1275));
    outputs(1617) <= layer0_outputs(900);
    outputs(1618) <= not(layer0_outputs(2813));
    outputs(1619) <= layer0_outputs(1481);
    outputs(1620) <= not(layer0_outputs(2300));
    outputs(1621) <= layer0_outputs(269);
    outputs(1622) <= (layer0_outputs(3516)) xor (layer0_outputs(3566));
    outputs(1623) <= not(layer0_outputs(7080));
    outputs(1624) <= not(layer0_outputs(4008));
    outputs(1625) <= not(layer0_outputs(5861)) or (layer0_outputs(6914));
    outputs(1626) <= not(layer0_outputs(5117));
    outputs(1627) <= not(layer0_outputs(7565)) or (layer0_outputs(2801));
    outputs(1628) <= (layer0_outputs(4730)) xor (layer0_outputs(4373));
    outputs(1629) <= layer0_outputs(1636);
    outputs(1630) <= not(layer0_outputs(5770)) or (layer0_outputs(4408));
    outputs(1631) <= not(layer0_outputs(720)) or (layer0_outputs(415));
    outputs(1632) <= not(layer0_outputs(1594));
    outputs(1633) <= layer0_outputs(774);
    outputs(1634) <= not(layer0_outputs(4855)) or (layer0_outputs(2444));
    outputs(1635) <= not(layer0_outputs(5950));
    outputs(1636) <= not((layer0_outputs(4782)) and (layer0_outputs(6519)));
    outputs(1637) <= not(layer0_outputs(5443));
    outputs(1638) <= layer0_outputs(1194);
    outputs(1639) <= '1';
    outputs(1640) <= not(layer0_outputs(7307)) or (layer0_outputs(2165));
    outputs(1641) <= not((layer0_outputs(7619)) xor (layer0_outputs(2213)));
    outputs(1642) <= not(layer0_outputs(3961));
    outputs(1643) <= not(layer0_outputs(7465));
    outputs(1644) <= layer0_outputs(5254);
    outputs(1645) <= layer0_outputs(554);
    outputs(1646) <= layer0_outputs(4476);
    outputs(1647) <= (layer0_outputs(6974)) xor (layer0_outputs(1610));
    outputs(1648) <= not((layer0_outputs(3051)) and (layer0_outputs(3215)));
    outputs(1649) <= not(layer0_outputs(6389));
    outputs(1650) <= not(layer0_outputs(6214));
    outputs(1651) <= layer0_outputs(5106);
    outputs(1652) <= not(layer0_outputs(3083));
    outputs(1653) <= not((layer0_outputs(5900)) and (layer0_outputs(3686)));
    outputs(1654) <= not((layer0_outputs(2159)) xor (layer0_outputs(4177)));
    outputs(1655) <= (layer0_outputs(5321)) and not (layer0_outputs(6740));
    outputs(1656) <= not(layer0_outputs(4367));
    outputs(1657) <= layer0_outputs(3301);
    outputs(1658) <= (layer0_outputs(1063)) or (layer0_outputs(5276));
    outputs(1659) <= not((layer0_outputs(5545)) xor (layer0_outputs(5601)));
    outputs(1660) <= layer0_outputs(2892);
    outputs(1661) <= (layer0_outputs(6645)) and not (layer0_outputs(3581));
    outputs(1662) <= layer0_outputs(308);
    outputs(1663) <= layer0_outputs(1947);
    outputs(1664) <= not(layer0_outputs(6132)) or (layer0_outputs(1540));
    outputs(1665) <= layer0_outputs(373);
    outputs(1666) <= not((layer0_outputs(4054)) xor (layer0_outputs(35)));
    outputs(1667) <= not(layer0_outputs(7077));
    outputs(1668) <= (layer0_outputs(437)) or (layer0_outputs(5237));
    outputs(1669) <= layer0_outputs(392);
    outputs(1670) <= not(layer0_outputs(15)) or (layer0_outputs(3016));
    outputs(1671) <= not(layer0_outputs(6892));
    outputs(1672) <= not(layer0_outputs(1562)) or (layer0_outputs(3904));
    outputs(1673) <= layer0_outputs(1964);
    outputs(1674) <= not((layer0_outputs(5280)) and (layer0_outputs(1144)));
    outputs(1675) <= (layer0_outputs(3499)) and not (layer0_outputs(4445));
    outputs(1676) <= layer0_outputs(1968);
    outputs(1677) <= (layer0_outputs(3461)) and not (layer0_outputs(5445));
    outputs(1678) <= not(layer0_outputs(7227));
    outputs(1679) <= not(layer0_outputs(6858));
    outputs(1680) <= not((layer0_outputs(131)) or (layer0_outputs(429)));
    outputs(1681) <= (layer0_outputs(2498)) xor (layer0_outputs(4953));
    outputs(1682) <= not(layer0_outputs(2041));
    outputs(1683) <= (layer0_outputs(5854)) xor (layer0_outputs(7014));
    outputs(1684) <= (layer0_outputs(64)) or (layer0_outputs(3424));
    outputs(1685) <= not((layer0_outputs(2312)) xor (layer0_outputs(5445)));
    outputs(1686) <= layer0_outputs(3037);
    outputs(1687) <= not(layer0_outputs(6951));
    outputs(1688) <= layer0_outputs(1837);
    outputs(1689) <= (layer0_outputs(2122)) xor (layer0_outputs(1005));
    outputs(1690) <= layer0_outputs(5274);
    outputs(1691) <= layer0_outputs(1945);
    outputs(1692) <= layer0_outputs(6047);
    outputs(1693) <= not(layer0_outputs(1208)) or (layer0_outputs(3004));
    outputs(1694) <= not((layer0_outputs(5045)) and (layer0_outputs(4926)));
    outputs(1695) <= layer0_outputs(5729);
    outputs(1696) <= layer0_outputs(4115);
    outputs(1697) <= layer0_outputs(871);
    outputs(1698) <= not(layer0_outputs(2332)) or (layer0_outputs(4075));
    outputs(1699) <= layer0_outputs(5037);
    outputs(1700) <= not((layer0_outputs(5980)) xor (layer0_outputs(3275)));
    outputs(1701) <= layer0_outputs(4656);
    outputs(1702) <= layer0_outputs(4289);
    outputs(1703) <= (layer0_outputs(5562)) or (layer0_outputs(7134));
    outputs(1704) <= not(layer0_outputs(4139));
    outputs(1705) <= (layer0_outputs(2429)) and not (layer0_outputs(1774));
    outputs(1706) <= not(layer0_outputs(4470));
    outputs(1707) <= (layer0_outputs(4158)) or (layer0_outputs(2990));
    outputs(1708) <= layer0_outputs(106);
    outputs(1709) <= not((layer0_outputs(507)) and (layer0_outputs(3321)));
    outputs(1710) <= not(layer0_outputs(3982)) or (layer0_outputs(5490));
    outputs(1711) <= not((layer0_outputs(1737)) xor (layer0_outputs(7053)));
    outputs(1712) <= layer0_outputs(7504);
    outputs(1713) <= not(layer0_outputs(327));
    outputs(1714) <= not(layer0_outputs(6523));
    outputs(1715) <= (layer0_outputs(1084)) and not (layer0_outputs(6290));
    outputs(1716) <= not((layer0_outputs(6080)) and (layer0_outputs(1132)));
    outputs(1717) <= (layer0_outputs(4308)) xor (layer0_outputs(267));
    outputs(1718) <= layer0_outputs(371);
    outputs(1719) <= (layer0_outputs(6298)) and (layer0_outputs(7524));
    outputs(1720) <= not((layer0_outputs(2866)) and (layer0_outputs(431)));
    outputs(1721) <= layer0_outputs(4245);
    outputs(1722) <= not(layer0_outputs(4337));
    outputs(1723) <= (layer0_outputs(3283)) or (layer0_outputs(21));
    outputs(1724) <= not((layer0_outputs(1080)) xor (layer0_outputs(4067)));
    outputs(1725) <= layer0_outputs(7552);
    outputs(1726) <= not((layer0_outputs(4357)) or (layer0_outputs(1283)));
    outputs(1727) <= (layer0_outputs(7323)) or (layer0_outputs(2039));
    outputs(1728) <= layer0_outputs(330);
    outputs(1729) <= layer0_outputs(5134);
    outputs(1730) <= not((layer0_outputs(2548)) or (layer0_outputs(4518)));
    outputs(1731) <= not(layer0_outputs(4965));
    outputs(1732) <= not(layer0_outputs(1276));
    outputs(1733) <= not(layer0_outputs(2116));
    outputs(1734) <= layer0_outputs(4241);
    outputs(1735) <= not(layer0_outputs(2035));
    outputs(1736) <= not((layer0_outputs(1588)) and (layer0_outputs(2469)));
    outputs(1737) <= not(layer0_outputs(979)) or (layer0_outputs(3459));
    outputs(1738) <= (layer0_outputs(1048)) or (layer0_outputs(5151));
    outputs(1739) <= not((layer0_outputs(4639)) and (layer0_outputs(4490)));
    outputs(1740) <= layer0_outputs(5775);
    outputs(1741) <= not(layer0_outputs(632));
    outputs(1742) <= not((layer0_outputs(7232)) xor (layer0_outputs(7598)));
    outputs(1743) <= layer0_outputs(1021);
    outputs(1744) <= layer0_outputs(7356);
    outputs(1745) <= layer0_outputs(2105);
    outputs(1746) <= layer0_outputs(4178);
    outputs(1747) <= not((layer0_outputs(2345)) xor (layer0_outputs(3270)));
    outputs(1748) <= layer0_outputs(5778);
    outputs(1749) <= (layer0_outputs(7652)) xor (layer0_outputs(1025));
    outputs(1750) <= (layer0_outputs(4048)) and (layer0_outputs(219));
    outputs(1751) <= layer0_outputs(5933);
    outputs(1752) <= layer0_outputs(839);
    outputs(1753) <= layer0_outputs(7373);
    outputs(1754) <= not(layer0_outputs(951));
    outputs(1755) <= (layer0_outputs(5494)) or (layer0_outputs(2455));
    outputs(1756) <= not(layer0_outputs(2393)) or (layer0_outputs(7111));
    outputs(1757) <= layer0_outputs(1349);
    outputs(1758) <= (layer0_outputs(5573)) or (layer0_outputs(6884));
    outputs(1759) <= not((layer0_outputs(6522)) xor (layer0_outputs(2054)));
    outputs(1760) <= (layer0_outputs(6589)) xor (layer0_outputs(2940));
    outputs(1761) <= layer0_outputs(1832);
    outputs(1762) <= not(layer0_outputs(3298));
    outputs(1763) <= not(layer0_outputs(4441));
    outputs(1764) <= not(layer0_outputs(5330));
    outputs(1765) <= layer0_outputs(5308);
    outputs(1766) <= (layer0_outputs(4401)) or (layer0_outputs(1426));
    outputs(1767) <= layer0_outputs(4687);
    outputs(1768) <= layer0_outputs(4252);
    outputs(1769) <= layer0_outputs(1937);
    outputs(1770) <= not(layer0_outputs(2122));
    outputs(1771) <= layer0_outputs(6253);
    outputs(1772) <= not(layer0_outputs(2049));
    outputs(1773) <= (layer0_outputs(3398)) and not (layer0_outputs(808));
    outputs(1774) <= (layer0_outputs(7303)) xor (layer0_outputs(2202));
    outputs(1775) <= not((layer0_outputs(900)) xor (layer0_outputs(27)));
    outputs(1776) <= layer0_outputs(2218);
    outputs(1777) <= (layer0_outputs(648)) or (layer0_outputs(218));
    outputs(1778) <= (layer0_outputs(2255)) and (layer0_outputs(5724));
    outputs(1779) <= not(layer0_outputs(4875)) or (layer0_outputs(4344));
    outputs(1780) <= layer0_outputs(5600);
    outputs(1781) <= not(layer0_outputs(3300));
    outputs(1782) <= not(layer0_outputs(5047));
    outputs(1783) <= (layer0_outputs(5895)) and not (layer0_outputs(7561));
    outputs(1784) <= not(layer0_outputs(6257));
    outputs(1785) <= not(layer0_outputs(6881)) or (layer0_outputs(4021));
    outputs(1786) <= not((layer0_outputs(6657)) and (layer0_outputs(6300)));
    outputs(1787) <= (layer0_outputs(4651)) xor (layer0_outputs(1952));
    outputs(1788) <= not((layer0_outputs(7372)) xor (layer0_outputs(338)));
    outputs(1789) <= not(layer0_outputs(6511));
    outputs(1790) <= not(layer0_outputs(5255));
    outputs(1791) <= not(layer0_outputs(6655));
    outputs(1792) <= layer0_outputs(6888);
    outputs(1793) <= layer0_outputs(4519);
    outputs(1794) <= layer0_outputs(3442);
    outputs(1795) <= (layer0_outputs(1766)) xor (layer0_outputs(3266));
    outputs(1796) <= layer0_outputs(6288);
    outputs(1797) <= not((layer0_outputs(1218)) xor (layer0_outputs(4710)));
    outputs(1798) <= not(layer0_outputs(1724));
    outputs(1799) <= not(layer0_outputs(1912)) or (layer0_outputs(4913));
    outputs(1800) <= (layer0_outputs(5587)) and not (layer0_outputs(5976));
    outputs(1801) <= not(layer0_outputs(6552));
    outputs(1802) <= not(layer0_outputs(7401));
    outputs(1803) <= not(layer0_outputs(6009));
    outputs(1804) <= (layer0_outputs(4062)) xor (layer0_outputs(6958));
    outputs(1805) <= not(layer0_outputs(2886));
    outputs(1806) <= not(layer0_outputs(2459));
    outputs(1807) <= (layer0_outputs(1120)) or (layer0_outputs(3733));
    outputs(1808) <= not((layer0_outputs(4641)) xor (layer0_outputs(3670)));
    outputs(1809) <= (layer0_outputs(2107)) or (layer0_outputs(2690));
    outputs(1810) <= not((layer0_outputs(1360)) or (layer0_outputs(5173)));
    outputs(1811) <= not((layer0_outputs(7595)) xor (layer0_outputs(7265)));
    outputs(1812) <= not(layer0_outputs(1802));
    outputs(1813) <= not(layer0_outputs(7409));
    outputs(1814) <= not((layer0_outputs(1151)) and (layer0_outputs(5869)));
    outputs(1815) <= not(layer0_outputs(7194));
    outputs(1816) <= not(layer0_outputs(741));
    outputs(1817) <= not(layer0_outputs(5528)) or (layer0_outputs(5446));
    outputs(1818) <= layer0_outputs(5241);
    outputs(1819) <= (layer0_outputs(4528)) or (layer0_outputs(4116));
    outputs(1820) <= (layer0_outputs(485)) and (layer0_outputs(3591));
    outputs(1821) <= not(layer0_outputs(253));
    outputs(1822) <= not(layer0_outputs(6054));
    outputs(1823) <= (layer0_outputs(6448)) or (layer0_outputs(1934));
    outputs(1824) <= not((layer0_outputs(6175)) xor (layer0_outputs(1531)));
    outputs(1825) <= layer0_outputs(7082);
    outputs(1826) <= not((layer0_outputs(4862)) xor (layer0_outputs(4201)));
    outputs(1827) <= layer0_outputs(5439);
    outputs(1828) <= not(layer0_outputs(6348)) or (layer0_outputs(600));
    outputs(1829) <= layer0_outputs(1340);
    outputs(1830) <= not(layer0_outputs(7673));
    outputs(1831) <= (layer0_outputs(4205)) xor (layer0_outputs(4536));
    outputs(1832) <= not(layer0_outputs(11)) or (layer0_outputs(93));
    outputs(1833) <= not((layer0_outputs(1105)) xor (layer0_outputs(4165)));
    outputs(1834) <= not(layer0_outputs(7511));
    outputs(1835) <= not(layer0_outputs(156));
    outputs(1836) <= not((layer0_outputs(4695)) xor (layer0_outputs(5659)));
    outputs(1837) <= not(layer0_outputs(6150)) or (layer0_outputs(2168));
    outputs(1838) <= not((layer0_outputs(2852)) or (layer0_outputs(7362)));
    outputs(1839) <= not((layer0_outputs(6634)) xor (layer0_outputs(3925)));
    outputs(1840) <= not(layer0_outputs(6383));
    outputs(1841) <= (layer0_outputs(2825)) xor (layer0_outputs(3084));
    outputs(1842) <= not((layer0_outputs(5098)) xor (layer0_outputs(5506)));
    outputs(1843) <= (layer0_outputs(3001)) xor (layer0_outputs(2813));
    outputs(1844) <= '1';
    outputs(1845) <= not(layer0_outputs(5876));
    outputs(1846) <= (layer0_outputs(4241)) and (layer0_outputs(3630));
    outputs(1847) <= not((layer0_outputs(2251)) xor (layer0_outputs(7020)));
    outputs(1848) <= not(layer0_outputs(905));
    outputs(1849) <= layer0_outputs(4915);
    outputs(1850) <= (layer0_outputs(98)) or (layer0_outputs(5057));
    outputs(1851) <= not((layer0_outputs(4643)) and (layer0_outputs(1004)));
    outputs(1852) <= not(layer0_outputs(6061));
    outputs(1853) <= (layer0_outputs(7433)) or (layer0_outputs(7091));
    outputs(1854) <= not((layer0_outputs(5227)) xor (layer0_outputs(4361)));
    outputs(1855) <= not(layer0_outputs(7144));
    outputs(1856) <= (layer0_outputs(1887)) xor (layer0_outputs(1114));
    outputs(1857) <= not(layer0_outputs(1710)) or (layer0_outputs(114));
    outputs(1858) <= not(layer0_outputs(3517));
    outputs(1859) <= (layer0_outputs(4321)) xor (layer0_outputs(3002));
    outputs(1860) <= not(layer0_outputs(1558));
    outputs(1861) <= not((layer0_outputs(4702)) xor (layer0_outputs(1950)));
    outputs(1862) <= not((layer0_outputs(1918)) and (layer0_outputs(1955)));
    outputs(1863) <= not(layer0_outputs(7116)) or (layer0_outputs(7347));
    outputs(1864) <= not((layer0_outputs(2523)) xor (layer0_outputs(6677)));
    outputs(1865) <= not(layer0_outputs(5073));
    outputs(1866) <= layer0_outputs(2102);
    outputs(1867) <= not(layer0_outputs(14)) or (layer0_outputs(6055));
    outputs(1868) <= (layer0_outputs(6195)) or (layer0_outputs(3427));
    outputs(1869) <= (layer0_outputs(2462)) and not (layer0_outputs(4479));
    outputs(1870) <= not((layer0_outputs(7633)) or (layer0_outputs(5591)));
    outputs(1871) <= layer0_outputs(7382);
    outputs(1872) <= not(layer0_outputs(4122));
    outputs(1873) <= not(layer0_outputs(7182));
    outputs(1874) <= layer0_outputs(2178);
    outputs(1875) <= not(layer0_outputs(516)) or (layer0_outputs(1948));
    outputs(1876) <= not(layer0_outputs(3299));
    outputs(1877) <= (layer0_outputs(7351)) xor (layer0_outputs(2616));
    outputs(1878) <= layer0_outputs(2153);
    outputs(1879) <= not((layer0_outputs(2206)) xor (layer0_outputs(7208)));
    outputs(1880) <= not(layer0_outputs(2831));
    outputs(1881) <= not((layer0_outputs(1245)) xor (layer0_outputs(5703)));
    outputs(1882) <= not((layer0_outputs(7606)) xor (layer0_outputs(7432)));
    outputs(1883) <= not((layer0_outputs(42)) or (layer0_outputs(2479)));
    outputs(1884) <= layer0_outputs(5919);
    outputs(1885) <= not((layer0_outputs(1660)) and (layer0_outputs(1088)));
    outputs(1886) <= not((layer0_outputs(5908)) xor (layer0_outputs(5392)));
    outputs(1887) <= not((layer0_outputs(5516)) and (layer0_outputs(3014)));
    outputs(1888) <= (layer0_outputs(1659)) and (layer0_outputs(1927));
    outputs(1889) <= not(layer0_outputs(3946)) or (layer0_outputs(2268));
    outputs(1890) <= (layer0_outputs(1198)) and (layer0_outputs(3049));
    outputs(1891) <= layer0_outputs(4750);
    outputs(1892) <= not((layer0_outputs(3273)) and (layer0_outputs(7170)));
    outputs(1893) <= not(layer0_outputs(4522)) or (layer0_outputs(4785));
    outputs(1894) <= layer0_outputs(282);
    outputs(1895) <= not((layer0_outputs(4524)) xor (layer0_outputs(5040)));
    outputs(1896) <= (layer0_outputs(684)) xor (layer0_outputs(2234));
    outputs(1897) <= not(layer0_outputs(3345));
    outputs(1898) <= not(layer0_outputs(5625));
    outputs(1899) <= not(layer0_outputs(603));
    outputs(1900) <= layer0_outputs(284);
    outputs(1901) <= not((layer0_outputs(3157)) xor (layer0_outputs(151)));
    outputs(1902) <= not(layer0_outputs(7163));
    outputs(1903) <= layer0_outputs(298);
    outputs(1904) <= layer0_outputs(6924);
    outputs(1905) <= not(layer0_outputs(4382));
    outputs(1906) <= not(layer0_outputs(697)) or (layer0_outputs(5614));
    outputs(1907) <= not((layer0_outputs(6110)) xor (layer0_outputs(1975)));
    outputs(1908) <= not((layer0_outputs(1528)) and (layer0_outputs(453)));
    outputs(1909) <= layer0_outputs(7161);
    outputs(1910) <= (layer0_outputs(6849)) and not (layer0_outputs(1622));
    outputs(1911) <= not(layer0_outputs(3282)) or (layer0_outputs(4826));
    outputs(1912) <= not(layer0_outputs(6483));
    outputs(1913) <= not(layer0_outputs(2400));
    outputs(1914) <= (layer0_outputs(1962)) and not (layer0_outputs(4270));
    outputs(1915) <= not((layer0_outputs(3078)) xor (layer0_outputs(1041)));
    outputs(1916) <= not((layer0_outputs(5679)) and (layer0_outputs(5095)));
    outputs(1917) <= not((layer0_outputs(4821)) or (layer0_outputs(6423)));
    outputs(1918) <= (layer0_outputs(2592)) xor (layer0_outputs(6310));
    outputs(1919) <= not(layer0_outputs(3066));
    outputs(1920) <= layer0_outputs(7528);
    outputs(1921) <= layer0_outputs(6056);
    outputs(1922) <= layer0_outputs(902);
    outputs(1923) <= not(layer0_outputs(5157));
    outputs(1924) <= not(layer0_outputs(3659));
    outputs(1925) <= not(layer0_outputs(6384));
    outputs(1926) <= '1';
    outputs(1927) <= layer0_outputs(6954);
    outputs(1928) <= (layer0_outputs(1992)) or (layer0_outputs(5187));
    outputs(1929) <= not(layer0_outputs(6544)) or (layer0_outputs(7320));
    outputs(1930) <= (layer0_outputs(6070)) xor (layer0_outputs(4627));
    outputs(1931) <= (layer0_outputs(394)) and (layer0_outputs(2092));
    outputs(1932) <= (layer0_outputs(282)) xor (layer0_outputs(6886));
    outputs(1933) <= layer0_outputs(4980);
    outputs(1934) <= (layer0_outputs(6235)) and (layer0_outputs(6592));
    outputs(1935) <= not(layer0_outputs(5635));
    outputs(1936) <= layer0_outputs(4554);
    outputs(1937) <= (layer0_outputs(7321)) xor (layer0_outputs(963));
    outputs(1938) <= layer0_outputs(2730);
    outputs(1939) <= layer0_outputs(7516);
    outputs(1940) <= (layer0_outputs(6771)) or (layer0_outputs(6837));
    outputs(1941) <= (layer0_outputs(3210)) xor (layer0_outputs(4879));
    outputs(1942) <= layer0_outputs(3618);
    outputs(1943) <= not(layer0_outputs(483));
    outputs(1944) <= layer0_outputs(2110);
    outputs(1945) <= (layer0_outputs(4921)) and not (layer0_outputs(1192));
    outputs(1946) <= not(layer0_outputs(792));
    outputs(1947) <= (layer0_outputs(3263)) xor (layer0_outputs(267));
    outputs(1948) <= not(layer0_outputs(2394));
    outputs(1949) <= not(layer0_outputs(5481));
    outputs(1950) <= (layer0_outputs(839)) or (layer0_outputs(3953));
    outputs(1951) <= not((layer0_outputs(5705)) and (layer0_outputs(2446)));
    outputs(1952) <= not(layer0_outputs(5005)) or (layer0_outputs(3959));
    outputs(1953) <= (layer0_outputs(5647)) xor (layer0_outputs(1383));
    outputs(1954) <= (layer0_outputs(2997)) xor (layer0_outputs(4018));
    outputs(1955) <= layer0_outputs(6683);
    outputs(1956) <= layer0_outputs(571);
    outputs(1957) <= not(layer0_outputs(2549));
    outputs(1958) <= not(layer0_outputs(1225)) or (layer0_outputs(3407));
    outputs(1959) <= not(layer0_outputs(1910));
    outputs(1960) <= not(layer0_outputs(5999)) or (layer0_outputs(3963));
    outputs(1961) <= layer0_outputs(1944);
    outputs(1962) <= layer0_outputs(4469);
    outputs(1963) <= not(layer0_outputs(6548)) or (layer0_outputs(1493));
    outputs(1964) <= not((layer0_outputs(3712)) xor (layer0_outputs(1872)));
    outputs(1965) <= not(layer0_outputs(3863)) or (layer0_outputs(1049));
    outputs(1966) <= (layer0_outputs(4428)) xor (layer0_outputs(1486));
    outputs(1967) <= (layer0_outputs(4681)) and not (layer0_outputs(7004));
    outputs(1968) <= not(layer0_outputs(664));
    outputs(1969) <= (layer0_outputs(5019)) and (layer0_outputs(7521));
    outputs(1970) <= not(layer0_outputs(4494)) or (layer0_outputs(4224));
    outputs(1971) <= layer0_outputs(7445);
    outputs(1972) <= not(layer0_outputs(6513));
    outputs(1973) <= not(layer0_outputs(5198));
    outputs(1974) <= not(layer0_outputs(3935));
    outputs(1975) <= (layer0_outputs(1309)) and not (layer0_outputs(7072));
    outputs(1976) <= not(layer0_outputs(6725));
    outputs(1977) <= layer0_outputs(4115);
    outputs(1978) <= not((layer0_outputs(4670)) or (layer0_outputs(6500)));
    outputs(1979) <= layer0_outputs(3204);
    outputs(1980) <= not((layer0_outputs(4155)) xor (layer0_outputs(5557)));
    outputs(1981) <= not((layer0_outputs(1798)) xor (layer0_outputs(5661)));
    outputs(1982) <= layer0_outputs(1480);
    outputs(1983) <= not(layer0_outputs(226));
    outputs(1984) <= (layer0_outputs(4886)) and not (layer0_outputs(3684));
    outputs(1985) <= not(layer0_outputs(5816));
    outputs(1986) <= not(layer0_outputs(1977));
    outputs(1987) <= not(layer0_outputs(3351));
    outputs(1988) <= (layer0_outputs(7145)) or (layer0_outputs(3752));
    outputs(1989) <= not(layer0_outputs(2749));
    outputs(1990) <= (layer0_outputs(4234)) and not (layer0_outputs(2388));
    outputs(1991) <= not(layer0_outputs(4073)) or (layer0_outputs(6265));
    outputs(1992) <= not(layer0_outputs(7182)) or (layer0_outputs(7304));
    outputs(1993) <= not(layer0_outputs(5690));
    outputs(1994) <= (layer0_outputs(7659)) xor (layer0_outputs(595));
    outputs(1995) <= not(layer0_outputs(3478));
    outputs(1996) <= not(layer0_outputs(6164)) or (layer0_outputs(920));
    outputs(1997) <= layer0_outputs(2960);
    outputs(1998) <= (layer0_outputs(4724)) xor (layer0_outputs(7413));
    outputs(1999) <= not((layer0_outputs(4660)) xor (layer0_outputs(2441)));
    outputs(2000) <= layer0_outputs(3834);
    outputs(2001) <= not((layer0_outputs(5464)) xor (layer0_outputs(2272)));
    outputs(2002) <= not(layer0_outputs(5469));
    outputs(2003) <= (layer0_outputs(5646)) and not (layer0_outputs(2327));
    outputs(2004) <= not(layer0_outputs(3038));
    outputs(2005) <= not(layer0_outputs(4322)) or (layer0_outputs(3440));
    outputs(2006) <= not(layer0_outputs(625));
    outputs(2007) <= (layer0_outputs(3276)) xor (layer0_outputs(207));
    outputs(2008) <= not(layer0_outputs(2713));
    outputs(2009) <= (layer0_outputs(7658)) and not (layer0_outputs(5330));
    outputs(2010) <= layer0_outputs(3480);
    outputs(2011) <= layer0_outputs(5663);
    outputs(2012) <= not((layer0_outputs(4498)) xor (layer0_outputs(5380)));
    outputs(2013) <= not(layer0_outputs(4926)) or (layer0_outputs(4513));
    outputs(2014) <= (layer0_outputs(712)) xor (layer0_outputs(115));
    outputs(2015) <= not(layer0_outputs(6760));
    outputs(2016) <= not((layer0_outputs(3095)) xor (layer0_outputs(1723)));
    outputs(2017) <= not(layer0_outputs(6555)) or (layer0_outputs(385));
    outputs(2018) <= (layer0_outputs(3362)) and not (layer0_outputs(3082));
    outputs(2019) <= layer0_outputs(640);
    outputs(2020) <= (layer0_outputs(6173)) and not (layer0_outputs(977));
    outputs(2021) <= layer0_outputs(6756);
    outputs(2022) <= (layer0_outputs(6643)) xor (layer0_outputs(3940));
    outputs(2023) <= not((layer0_outputs(1638)) or (layer0_outputs(6439)));
    outputs(2024) <= not(layer0_outputs(807)) or (layer0_outputs(2820));
    outputs(2025) <= (layer0_outputs(4214)) xor (layer0_outputs(4316));
    outputs(2026) <= layer0_outputs(3610);
    outputs(2027) <= (layer0_outputs(5036)) xor (layer0_outputs(6351));
    outputs(2028) <= not(layer0_outputs(3202)) or (layer0_outputs(3237));
    outputs(2029) <= not(layer0_outputs(2035));
    outputs(2030) <= not((layer0_outputs(3163)) xor (layer0_outputs(6291)));
    outputs(2031) <= layer0_outputs(7187);
    outputs(2032) <= not(layer0_outputs(5378)) or (layer0_outputs(4812));
    outputs(2033) <= (layer0_outputs(615)) or (layer0_outputs(194));
    outputs(2034) <= not(layer0_outputs(1763));
    outputs(2035) <= not(layer0_outputs(1388));
    outputs(2036) <= (layer0_outputs(4762)) xor (layer0_outputs(3850));
    outputs(2037) <= not(layer0_outputs(6668));
    outputs(2038) <= (layer0_outputs(5433)) and not (layer0_outputs(6824));
    outputs(2039) <= layer0_outputs(6188);
    outputs(2040) <= not((layer0_outputs(5220)) or (layer0_outputs(4868)));
    outputs(2041) <= not(layer0_outputs(300));
    outputs(2042) <= not(layer0_outputs(5233));
    outputs(2043) <= not((layer0_outputs(4040)) xor (layer0_outputs(4793)));
    outputs(2044) <= (layer0_outputs(6791)) and not (layer0_outputs(3889));
    outputs(2045) <= not(layer0_outputs(503));
    outputs(2046) <= layer0_outputs(4767);
    outputs(2047) <= not(layer0_outputs(302)) or (layer0_outputs(862));
    outputs(2048) <= not((layer0_outputs(6006)) and (layer0_outputs(2594)));
    outputs(2049) <= not(layer0_outputs(6391));
    outputs(2050) <= layer0_outputs(7266);
    outputs(2051) <= not(layer0_outputs(6665));
    outputs(2052) <= not(layer0_outputs(2802)) or (layer0_outputs(7293));
    outputs(2053) <= layer0_outputs(4889);
    outputs(2054) <= not((layer0_outputs(2859)) and (layer0_outputs(2038)));
    outputs(2055) <= layer0_outputs(7262);
    outputs(2056) <= not(layer0_outputs(5499));
    outputs(2057) <= not((layer0_outputs(7202)) xor (layer0_outputs(7627)));
    outputs(2058) <= not(layer0_outputs(197)) or (layer0_outputs(6844));
    outputs(2059) <= not((layer0_outputs(7178)) or (layer0_outputs(446)));
    outputs(2060) <= not(layer0_outputs(6761));
    outputs(2061) <= layer0_outputs(7564);
    outputs(2062) <= not((layer0_outputs(5720)) or (layer0_outputs(2974)));
    outputs(2063) <= not(layer0_outputs(6906));
    outputs(2064) <= layer0_outputs(6402);
    outputs(2065) <= not((layer0_outputs(4014)) and (layer0_outputs(3641)));
    outputs(2066) <= not(layer0_outputs(4754));
    outputs(2067) <= not(layer0_outputs(1643));
    outputs(2068) <= (layer0_outputs(1160)) and (layer0_outputs(2980));
    outputs(2069) <= not(layer0_outputs(7351)) or (layer0_outputs(2408));
    outputs(2070) <= layer0_outputs(94);
    outputs(2071) <= (layer0_outputs(946)) xor (layer0_outputs(4501));
    outputs(2072) <= (layer0_outputs(1342)) xor (layer0_outputs(6968));
    outputs(2073) <= not(layer0_outputs(7557)) or (layer0_outputs(548));
    outputs(2074) <= not((layer0_outputs(2284)) xor (layer0_outputs(959)));
    outputs(2075) <= (layer0_outputs(549)) or (layer0_outputs(1102));
    outputs(2076) <= not(layer0_outputs(5925)) or (layer0_outputs(4053));
    outputs(2077) <= (layer0_outputs(2890)) xor (layer0_outputs(6342));
    outputs(2078) <= not(layer0_outputs(359));
    outputs(2079) <= layer0_outputs(6626);
    outputs(2080) <= (layer0_outputs(1033)) and not (layer0_outputs(6785));
    outputs(2081) <= not(layer0_outputs(2586)) or (layer0_outputs(6631));
    outputs(2082) <= (layer0_outputs(690)) xor (layer0_outputs(6349));
    outputs(2083) <= not((layer0_outputs(5229)) xor (layer0_outputs(1442)));
    outputs(2084) <= not(layer0_outputs(4718));
    outputs(2085) <= not(layer0_outputs(7472));
    outputs(2086) <= not(layer0_outputs(1404)) or (layer0_outputs(4505));
    outputs(2087) <= (layer0_outputs(6256)) xor (layer0_outputs(5193));
    outputs(2088) <= (layer0_outputs(5912)) xor (layer0_outputs(6691));
    outputs(2089) <= not(layer0_outputs(5730)) or (layer0_outputs(3179));
    outputs(2090) <= not((layer0_outputs(4130)) and (layer0_outputs(1208)));
    outputs(2091) <= (layer0_outputs(362)) xor (layer0_outputs(4394));
    outputs(2092) <= not(layer0_outputs(813));
    outputs(2093) <= not(layer0_outputs(1679));
    outputs(2094) <= layer0_outputs(4598);
    outputs(2095) <= not((layer0_outputs(6261)) or (layer0_outputs(6686)));
    outputs(2096) <= layer0_outputs(1184);
    outputs(2097) <= not(layer0_outputs(1129));
    outputs(2098) <= (layer0_outputs(35)) and (layer0_outputs(181));
    outputs(2099) <= layer0_outputs(4384);
    outputs(2100) <= (layer0_outputs(2215)) or (layer0_outputs(2457));
    outputs(2101) <= not((layer0_outputs(7365)) xor (layer0_outputs(3268)));
    outputs(2102) <= layer0_outputs(1163);
    outputs(2103) <= (layer0_outputs(5696)) xor (layer0_outputs(5295));
    outputs(2104) <= not((layer0_outputs(3656)) xor (layer0_outputs(2174)));
    outputs(2105) <= layer0_outputs(2531);
    outputs(2106) <= layer0_outputs(2903);
    outputs(2107) <= (layer0_outputs(3575)) or (layer0_outputs(6698));
    outputs(2108) <= layer0_outputs(6283);
    outputs(2109) <= layer0_outputs(305);
    outputs(2110) <= not(layer0_outputs(6391));
    outputs(2111) <= layer0_outputs(6311);
    outputs(2112) <= (layer0_outputs(7124)) xor (layer0_outputs(4527));
    outputs(2113) <= (layer0_outputs(1376)) and (layer0_outputs(1128));
    outputs(2114) <= layer0_outputs(7638);
    outputs(2115) <= layer0_outputs(2465);
    outputs(2116) <= not(layer0_outputs(7364)) or (layer0_outputs(2331));
    outputs(2117) <= not((layer0_outputs(3406)) xor (layer0_outputs(4917)));
    outputs(2118) <= not((layer0_outputs(1815)) xor (layer0_outputs(5634)));
    outputs(2119) <= (layer0_outputs(759)) and (layer0_outputs(7258));
    outputs(2120) <= not(layer0_outputs(1749));
    outputs(2121) <= not(layer0_outputs(1103)) or (layer0_outputs(2804));
    outputs(2122) <= not((layer0_outputs(1975)) and (layer0_outputs(209)));
    outputs(2123) <= layer0_outputs(3800);
    outputs(2124) <= (layer0_outputs(1273)) xor (layer0_outputs(2061));
    outputs(2125) <= not((layer0_outputs(6428)) xor (layer0_outputs(722)));
    outputs(2126) <= not(layer0_outputs(3232));
    outputs(2127) <= not(layer0_outputs(6917)) or (layer0_outputs(7312));
    outputs(2128) <= not(layer0_outputs(1732));
    outputs(2129) <= (layer0_outputs(662)) and not (layer0_outputs(7617));
    outputs(2130) <= not((layer0_outputs(5475)) xor (layer0_outputs(5584)));
    outputs(2131) <= layer0_outputs(3496);
    outputs(2132) <= not(layer0_outputs(652));
    outputs(2133) <= not((layer0_outputs(7243)) or (layer0_outputs(4077)));
    outputs(2134) <= (layer0_outputs(919)) and not (layer0_outputs(2172));
    outputs(2135) <= (layer0_outputs(1301)) and not (layer0_outputs(7094));
    outputs(2136) <= not(layer0_outputs(1801));
    outputs(2137) <= not(layer0_outputs(6781)) or (layer0_outputs(4607));
    outputs(2138) <= (layer0_outputs(5506)) xor (layer0_outputs(3693));
    outputs(2139) <= not((layer0_outputs(4904)) xor (layer0_outputs(2525)));
    outputs(2140) <= (layer0_outputs(2597)) or (layer0_outputs(4253));
    outputs(2141) <= (layer0_outputs(623)) or (layer0_outputs(766));
    outputs(2142) <= not((layer0_outputs(1502)) and (layer0_outputs(2925)));
    outputs(2143) <= not((layer0_outputs(7467)) xor (layer0_outputs(2501)));
    outputs(2144) <= not((layer0_outputs(5295)) xor (layer0_outputs(6309)));
    outputs(2145) <= not(layer0_outputs(2898));
    outputs(2146) <= layer0_outputs(705);
    outputs(2147) <= (layer0_outputs(6375)) and not (layer0_outputs(2077));
    outputs(2148) <= not(layer0_outputs(6503));
    outputs(2149) <= not((layer0_outputs(2872)) or (layer0_outputs(179)));
    outputs(2150) <= (layer0_outputs(3869)) and not (layer0_outputs(5863));
    outputs(2151) <= not(layer0_outputs(4832)) or (layer0_outputs(7431));
    outputs(2152) <= (layer0_outputs(6705)) xor (layer0_outputs(29));
    outputs(2153) <= (layer0_outputs(658)) and not (layer0_outputs(7543));
    outputs(2154) <= not(layer0_outputs(4060));
    outputs(2155) <= not(layer0_outputs(2844));
    outputs(2156) <= not(layer0_outputs(5128));
    outputs(2157) <= layer0_outputs(6667);
    outputs(2158) <= layer0_outputs(6915);
    outputs(2159) <= not(layer0_outputs(5118));
    outputs(2160) <= not(layer0_outputs(248));
    outputs(2161) <= not(layer0_outputs(5864));
    outputs(2162) <= not(layer0_outputs(3421));
    outputs(2163) <= not(layer0_outputs(4107)) or (layer0_outputs(7517));
    outputs(2164) <= not(layer0_outputs(100));
    outputs(2165) <= layer0_outputs(378);
    outputs(2166) <= not((layer0_outputs(3562)) xor (layer0_outputs(6659)));
    outputs(2167) <= not((layer0_outputs(4801)) or (layer0_outputs(7609)));
    outputs(2168) <= not(layer0_outputs(932));
    outputs(2169) <= not((layer0_outputs(4847)) xor (layer0_outputs(4509)));
    outputs(2170) <= layer0_outputs(1056);
    outputs(2171) <= not(layer0_outputs(5750));
    outputs(2172) <= (layer0_outputs(4236)) xor (layer0_outputs(4184));
    outputs(2173) <= not((layer0_outputs(3989)) or (layer0_outputs(4000)));
    outputs(2174) <= not((layer0_outputs(7510)) xor (layer0_outputs(1461)));
    outputs(2175) <= not((layer0_outputs(5117)) xor (layer0_outputs(3885)));
    outputs(2176) <= not(layer0_outputs(155));
    outputs(2177) <= not(layer0_outputs(3719)) or (layer0_outputs(3713));
    outputs(2178) <= (layer0_outputs(1776)) and (layer0_outputs(5735));
    outputs(2179) <= layer0_outputs(3984);
    outputs(2180) <= not(layer0_outputs(5320));
    outputs(2181) <= layer0_outputs(5305);
    outputs(2182) <= not((layer0_outputs(6764)) xor (layer0_outputs(6160)));
    outputs(2183) <= not(layer0_outputs(6082)) or (layer0_outputs(7300));
    outputs(2184) <= not(layer0_outputs(5422));
    outputs(2185) <= not((layer0_outputs(438)) or (layer0_outputs(159)));
    outputs(2186) <= layer0_outputs(2097);
    outputs(2187) <= (layer0_outputs(4282)) or (layer0_outputs(3595));
    outputs(2188) <= (layer0_outputs(6459)) or (layer0_outputs(4612));
    outputs(2189) <= not(layer0_outputs(6675)) or (layer0_outputs(1567));
    outputs(2190) <= not(layer0_outputs(5764));
    outputs(2191) <= layer0_outputs(5721);
    outputs(2192) <= (layer0_outputs(1882)) xor (layer0_outputs(535));
    outputs(2193) <= not(layer0_outputs(1072));
    outputs(2194) <= (layer0_outputs(2142)) xor (layer0_outputs(4127));
    outputs(2195) <= not(layer0_outputs(3835));
    outputs(2196) <= not((layer0_outputs(6344)) xor (layer0_outputs(5210)));
    outputs(2197) <= not(layer0_outputs(2338));
    outputs(2198) <= (layer0_outputs(1238)) or (layer0_outputs(288));
    outputs(2199) <= (layer0_outputs(7394)) or (layer0_outputs(5556));
    outputs(2200) <= layer0_outputs(593);
    outputs(2201) <= not(layer0_outputs(6032));
    outputs(2202) <= layer0_outputs(1145);
    outputs(2203) <= not((layer0_outputs(2251)) xor (layer0_outputs(3543)));
    outputs(2204) <= not((layer0_outputs(4044)) and (layer0_outputs(6752)));
    outputs(2205) <= not(layer0_outputs(1772)) or (layer0_outputs(6111));
    outputs(2206) <= (layer0_outputs(5477)) xor (layer0_outputs(1627));
    outputs(2207) <= (layer0_outputs(4110)) and not (layer0_outputs(575));
    outputs(2208) <= not(layer0_outputs(6458)) or (layer0_outputs(2099));
    outputs(2209) <= (layer0_outputs(1956)) xor (layer0_outputs(1772));
    outputs(2210) <= not(layer0_outputs(6921));
    outputs(2211) <= not(layer0_outputs(1853));
    outputs(2212) <= not(layer0_outputs(7006));
    outputs(2213) <= layer0_outputs(7488);
    outputs(2214) <= layer0_outputs(966);
    outputs(2215) <= not(layer0_outputs(7099));
    outputs(2216) <= not(layer0_outputs(6365)) or (layer0_outputs(7132));
    outputs(2217) <= (layer0_outputs(1967)) and not (layer0_outputs(7109));
    outputs(2218) <= layer0_outputs(1621);
    outputs(2219) <= layer0_outputs(416);
    outputs(2220) <= not(layer0_outputs(6972));
    outputs(2221) <= not(layer0_outputs(89));
    outputs(2222) <= (layer0_outputs(3499)) xor (layer0_outputs(3373));
    outputs(2223) <= layer0_outputs(6016);
    outputs(2224) <= not(layer0_outputs(1658));
    outputs(2225) <= (layer0_outputs(3174)) and not (layer0_outputs(7467));
    outputs(2226) <= layer0_outputs(7534);
    outputs(2227) <= not(layer0_outputs(141)) or (layer0_outputs(4912));
    outputs(2228) <= (layer0_outputs(3314)) xor (layer0_outputs(6973));
    outputs(2229) <= not((layer0_outputs(380)) or (layer0_outputs(699)));
    outputs(2230) <= layer0_outputs(2098);
    outputs(2231) <= not((layer0_outputs(2154)) xor (layer0_outputs(4234)));
    outputs(2232) <= not(layer0_outputs(1981)) or (layer0_outputs(2483));
    outputs(2233) <= not(layer0_outputs(122));
    outputs(2234) <= layer0_outputs(7497);
    outputs(2235) <= not(layer0_outputs(5856));
    outputs(2236) <= not(layer0_outputs(5113)) or (layer0_outputs(5992));
    outputs(2237) <= (layer0_outputs(2335)) and not (layer0_outputs(6059));
    outputs(2238) <= layer0_outputs(4395);
    outputs(2239) <= (layer0_outputs(1025)) xor (layer0_outputs(6786));
    outputs(2240) <= layer0_outputs(345);
    outputs(2241) <= (layer0_outputs(3304)) and (layer0_outputs(3496));
    outputs(2242) <= layer0_outputs(7159);
    outputs(2243) <= (layer0_outputs(4311)) and (layer0_outputs(7363));
    outputs(2244) <= layer0_outputs(2709);
    outputs(2245) <= not(layer0_outputs(4947)) or (layer0_outputs(787));
    outputs(2246) <= not((layer0_outputs(2368)) xor (layer0_outputs(2650)));
    outputs(2247) <= not((layer0_outputs(5118)) xor (layer0_outputs(6807)));
    outputs(2248) <= layer0_outputs(2205);
    outputs(2249) <= not(layer0_outputs(5090));
    outputs(2250) <= (layer0_outputs(2774)) and (layer0_outputs(168));
    outputs(2251) <= not(layer0_outputs(3691));
    outputs(2252) <= layer0_outputs(1782);
    outputs(2253) <= not((layer0_outputs(73)) and (layer0_outputs(2254)));
    outputs(2254) <= layer0_outputs(3384);
    outputs(2255) <= (layer0_outputs(1370)) xor (layer0_outputs(1084));
    outputs(2256) <= not(layer0_outputs(2493));
    outputs(2257) <= not(layer0_outputs(1901));
    outputs(2258) <= not(layer0_outputs(1424));
    outputs(2259) <= layer0_outputs(1754);
    outputs(2260) <= layer0_outputs(5067);
    outputs(2261) <= (layer0_outputs(2134)) and not (layer0_outputs(2809));
    outputs(2262) <= layer0_outputs(6438);
    outputs(2263) <= not((layer0_outputs(7251)) or (layer0_outputs(5250)));
    outputs(2264) <= (layer0_outputs(419)) xor (layer0_outputs(1458));
    outputs(2265) <= not(layer0_outputs(6269));
    outputs(2266) <= (layer0_outputs(2433)) xor (layer0_outputs(1963));
    outputs(2267) <= (layer0_outputs(3284)) xor (layer0_outputs(734));
    outputs(2268) <= not(layer0_outputs(1219));
    outputs(2269) <= not(layer0_outputs(1186));
    outputs(2270) <= (layer0_outputs(4072)) xor (layer0_outputs(5275));
    outputs(2271) <= layer0_outputs(1047);
    outputs(2272) <= not(layer0_outputs(5292));
    outputs(2273) <= not(layer0_outputs(5167));
    outputs(2274) <= (layer0_outputs(3619)) and not (layer0_outputs(4864));
    outputs(2275) <= layer0_outputs(117);
    outputs(2276) <= layer0_outputs(7024);
    outputs(2277) <= layer0_outputs(1564);
    outputs(2278) <= not(layer0_outputs(4815)) or (layer0_outputs(5426));
    outputs(2279) <= layer0_outputs(4492);
    outputs(2280) <= not((layer0_outputs(6900)) and (layer0_outputs(3563)));
    outputs(2281) <= not(layer0_outputs(5058)) or (layer0_outputs(6844));
    outputs(2282) <= (layer0_outputs(633)) or (layer0_outputs(6449));
    outputs(2283) <= layer0_outputs(852);
    outputs(2284) <= not(layer0_outputs(3418));
    outputs(2285) <= layer0_outputs(1913);
    outputs(2286) <= (layer0_outputs(2853)) and not (layer0_outputs(4014));
    outputs(2287) <= not(layer0_outputs(5467)) or (layer0_outputs(2679));
    outputs(2288) <= not((layer0_outputs(4814)) xor (layer0_outputs(3397)));
    outputs(2289) <= layer0_outputs(6424);
    outputs(2290) <= (layer0_outputs(6515)) or (layer0_outputs(2185));
    outputs(2291) <= not((layer0_outputs(1105)) or (layer0_outputs(3189)));
    outputs(2292) <= not((layer0_outputs(528)) xor (layer0_outputs(7377)));
    outputs(2293) <= not(layer0_outputs(2352)) or (layer0_outputs(885));
    outputs(2294) <= not(layer0_outputs(7348));
    outputs(2295) <= layer0_outputs(6330);
    outputs(2296) <= (layer0_outputs(5595)) or (layer0_outputs(4314));
    outputs(2297) <= not(layer0_outputs(7095));
    outputs(2298) <= not(layer0_outputs(3147));
    outputs(2299) <= not(layer0_outputs(469));
    outputs(2300) <= not((layer0_outputs(740)) or (layer0_outputs(4351)));
    outputs(2301) <= layer0_outputs(2027);
    outputs(2302) <= not(layer0_outputs(4704));
    outputs(2303) <= layer0_outputs(679);
    outputs(2304) <= (layer0_outputs(2761)) or (layer0_outputs(6201));
    outputs(2305) <= (layer0_outputs(5944)) and not (layer0_outputs(5716));
    outputs(2306) <= not((layer0_outputs(4302)) and (layer0_outputs(1321)));
    outputs(2307) <= layer0_outputs(7287);
    outputs(2308) <= layer0_outputs(3505);
    outputs(2309) <= not(layer0_outputs(7002)) or (layer0_outputs(3434));
    outputs(2310) <= layer0_outputs(1621);
    outputs(2311) <= not(layer0_outputs(228));
    outputs(2312) <= not(layer0_outputs(4591));
    outputs(2313) <= not((layer0_outputs(6075)) and (layer0_outputs(6112)));
    outputs(2314) <= not(layer0_outputs(2416)) or (layer0_outputs(3427));
    outputs(2315) <= not(layer0_outputs(3812));
    outputs(2316) <= not(layer0_outputs(1159));
    outputs(2317) <= layer0_outputs(2316);
    outputs(2318) <= not(layer0_outputs(4102)) or (layer0_outputs(3576));
    outputs(2319) <= (layer0_outputs(6526)) and (layer0_outputs(5775));
    outputs(2320) <= not((layer0_outputs(1170)) and (layer0_outputs(1392)));
    outputs(2321) <= not(layer0_outputs(5567));
    outputs(2322) <= layer0_outputs(2481);
    outputs(2323) <= layer0_outputs(3448);
    outputs(2324) <= layer0_outputs(3842);
    outputs(2325) <= layer0_outputs(5642);
    outputs(2326) <= (layer0_outputs(7359)) xor (layer0_outputs(3060));
    outputs(2327) <= not((layer0_outputs(3020)) or (layer0_outputs(4284)));
    outputs(2328) <= not(layer0_outputs(851));
    outputs(2329) <= (layer0_outputs(4094)) or (layer0_outputs(427));
    outputs(2330) <= (layer0_outputs(2617)) xor (layer0_outputs(5243));
    outputs(2331) <= (layer0_outputs(6160)) and not (layer0_outputs(747));
    outputs(2332) <= not(layer0_outputs(6872));
    outputs(2333) <= not(layer0_outputs(6164));
    outputs(2334) <= not(layer0_outputs(4914));
    outputs(2335) <= (layer0_outputs(5689)) and not (layer0_outputs(4466));
    outputs(2336) <= (layer0_outputs(5792)) xor (layer0_outputs(4429));
    outputs(2337) <= not(layer0_outputs(4862));
    outputs(2338) <= not(layer0_outputs(825));
    outputs(2339) <= layer0_outputs(7267);
    outputs(2340) <= layer0_outputs(7084);
    outputs(2341) <= layer0_outputs(4091);
    outputs(2342) <= not((layer0_outputs(2571)) xor (layer0_outputs(3593)));
    outputs(2343) <= not(layer0_outputs(5417));
    outputs(2344) <= not(layer0_outputs(4669));
    outputs(2345) <= not((layer0_outputs(5636)) xor (layer0_outputs(3649)));
    outputs(2346) <= layer0_outputs(3396);
    outputs(2347) <= layer0_outputs(5314);
    outputs(2348) <= layer0_outputs(629);
    outputs(2349) <= not((layer0_outputs(4871)) xor (layer0_outputs(4983)));
    outputs(2350) <= not(layer0_outputs(4588));
    outputs(2351) <= (layer0_outputs(3290)) xor (layer0_outputs(6504));
    outputs(2352) <= layer0_outputs(5403);
    outputs(2353) <= layer0_outputs(1569);
    outputs(2354) <= not(layer0_outputs(4187));
    outputs(2355) <= not((layer0_outputs(6671)) or (layer0_outputs(3240)));
    outputs(2356) <= (layer0_outputs(3758)) xor (layer0_outputs(6072));
    outputs(2357) <= (layer0_outputs(5525)) xor (layer0_outputs(1603));
    outputs(2358) <= layer0_outputs(5004);
    outputs(2359) <= (layer0_outputs(4067)) and not (layer0_outputs(5795));
    outputs(2360) <= layer0_outputs(1508);
    outputs(2361) <= not(layer0_outputs(5816));
    outputs(2362) <= not(layer0_outputs(6083));
    outputs(2363) <= layer0_outputs(6408);
    outputs(2364) <= (layer0_outputs(6271)) and (layer0_outputs(6650));
    outputs(2365) <= (layer0_outputs(760)) and not (layer0_outputs(6280));
    outputs(2366) <= layer0_outputs(7479);
    outputs(2367) <= layer0_outputs(5675);
    outputs(2368) <= (layer0_outputs(5007)) and not (layer0_outputs(3937));
    outputs(2369) <= not((layer0_outputs(369)) xor (layer0_outputs(6968)));
    outputs(2370) <= (layer0_outputs(6309)) xor (layer0_outputs(1411));
    outputs(2371) <= (layer0_outputs(5283)) and (layer0_outputs(1629));
    outputs(2372) <= (layer0_outputs(627)) xor (layer0_outputs(2472));
    outputs(2373) <= (layer0_outputs(3638)) xor (layer0_outputs(1382));
    outputs(2374) <= (layer0_outputs(3495)) xor (layer0_outputs(5817));
    outputs(2375) <= not((layer0_outputs(3201)) or (layer0_outputs(6542)));
    outputs(2376) <= layer0_outputs(3086);
    outputs(2377) <= not(layer0_outputs(1769));
    outputs(2378) <= not(layer0_outputs(4430)) or (layer0_outputs(3965));
    outputs(2379) <= (layer0_outputs(299)) xor (layer0_outputs(6063));
    outputs(2380) <= not(layer0_outputs(4356)) or (layer0_outputs(6775));
    outputs(2381) <= not(layer0_outputs(1852));
    outputs(2382) <= not(layer0_outputs(845)) or (layer0_outputs(651));
    outputs(2383) <= layer0_outputs(4340);
    outputs(2384) <= not(layer0_outputs(6812));
    outputs(2385) <= layer0_outputs(3469);
    outputs(2386) <= layer0_outputs(5661);
    outputs(2387) <= not((layer0_outputs(2557)) xor (layer0_outputs(3617)));
    outputs(2388) <= not(layer0_outputs(484));
    outputs(2389) <= (layer0_outputs(806)) xor (layer0_outputs(5207));
    outputs(2390) <= layer0_outputs(5722);
    outputs(2391) <= not((layer0_outputs(4058)) and (layer0_outputs(3625)));
    outputs(2392) <= layer0_outputs(3520);
    outputs(2393) <= (layer0_outputs(7672)) and not (layer0_outputs(1866));
    outputs(2394) <= (layer0_outputs(7411)) xor (layer0_outputs(2681));
    outputs(2395) <= not((layer0_outputs(4877)) and (layer0_outputs(7616)));
    outputs(2396) <= not(layer0_outputs(4791));
    outputs(2397) <= layer0_outputs(2250);
    outputs(2398) <= layer0_outputs(3143);
    outputs(2399) <= not((layer0_outputs(1598)) xor (layer0_outputs(2803)));
    outputs(2400) <= layer0_outputs(6660);
    outputs(2401) <= layer0_outputs(332);
    outputs(2402) <= (layer0_outputs(1351)) and not (layer0_outputs(2608));
    outputs(2403) <= not((layer0_outputs(166)) xor (layer0_outputs(7098)));
    outputs(2404) <= not((layer0_outputs(3278)) xor (layer0_outputs(6565)));
    outputs(2405) <= not((layer0_outputs(388)) xor (layer0_outputs(3804)));
    outputs(2406) <= not((layer0_outputs(5349)) and (layer0_outputs(6091)));
    outputs(2407) <= not(layer0_outputs(4911));
    outputs(2408) <= not(layer0_outputs(5990));
    outputs(2409) <= not(layer0_outputs(973));
    outputs(2410) <= (layer0_outputs(4065)) xor (layer0_outputs(6986));
    outputs(2411) <= (layer0_outputs(4698)) xor (layer0_outputs(4525));
    outputs(2412) <= (layer0_outputs(562)) xor (layer0_outputs(3314));
    outputs(2413) <= (layer0_outputs(5429)) and not (layer0_outputs(5989));
    outputs(2414) <= layer0_outputs(858);
    outputs(2415) <= not((layer0_outputs(1296)) xor (layer0_outputs(2895)));
    outputs(2416) <= layer0_outputs(2162);
    outputs(2417) <= (layer0_outputs(4653)) xor (layer0_outputs(1045));
    outputs(2418) <= not((layer0_outputs(6398)) xor (layer0_outputs(6327)));
    outputs(2419) <= not(layer0_outputs(1673));
    outputs(2420) <= not((layer0_outputs(4867)) xor (layer0_outputs(3472)));
    outputs(2421) <= not(layer0_outputs(75));
    outputs(2422) <= (layer0_outputs(4349)) xor (layer0_outputs(1504));
    outputs(2423) <= (layer0_outputs(6463)) xor (layer0_outputs(6368));
    outputs(2424) <= not((layer0_outputs(3775)) xor (layer0_outputs(7175)));
    outputs(2425) <= (layer0_outputs(1420)) xor (layer0_outputs(3741));
    outputs(2426) <= (layer0_outputs(525)) xor (layer0_outputs(5012));
    outputs(2427) <= not(layer0_outputs(1343));
    outputs(2428) <= not((layer0_outputs(2954)) xor (layer0_outputs(2739)));
    outputs(2429) <= not((layer0_outputs(2849)) xor (layer0_outputs(7095)));
    outputs(2430) <= not((layer0_outputs(1055)) xor (layer0_outputs(7044)));
    outputs(2431) <= not(layer0_outputs(4686)) or (layer0_outputs(4039));
    outputs(2432) <= not((layer0_outputs(3789)) xor (layer0_outputs(5260)));
    outputs(2433) <= not((layer0_outputs(6088)) xor (layer0_outputs(504)));
    outputs(2434) <= not(layer0_outputs(4776));
    outputs(2435) <= layer0_outputs(1451);
    outputs(2436) <= not((layer0_outputs(6770)) xor (layer0_outputs(335)));
    outputs(2437) <= not((layer0_outputs(1837)) xor (layer0_outputs(4610)));
    outputs(2438) <= not(layer0_outputs(3091));
    outputs(2439) <= layer0_outputs(5660);
    outputs(2440) <= not(layer0_outputs(6656)) or (layer0_outputs(2245));
    outputs(2441) <= (layer0_outputs(2055)) and not (layer0_outputs(2384));
    outputs(2442) <= not(layer0_outputs(51));
    outputs(2443) <= layer0_outputs(4195);
    outputs(2444) <= not(layer0_outputs(3464)) or (layer0_outputs(2480));
    outputs(2445) <= not((layer0_outputs(4634)) and (layer0_outputs(2773)));
    outputs(2446) <= not(layer0_outputs(1849));
    outputs(2447) <= layer0_outputs(4511);
    outputs(2448) <= not(layer0_outputs(6781));
    outputs(2449) <= not((layer0_outputs(4027)) xor (layer0_outputs(2123)));
    outputs(2450) <= not(layer0_outputs(3479)) or (layer0_outputs(2136));
    outputs(2451) <= (layer0_outputs(3490)) xor (layer0_outputs(2613));
    outputs(2452) <= (layer0_outputs(4764)) and (layer0_outputs(5109));
    outputs(2453) <= (layer0_outputs(3524)) xor (layer0_outputs(7048));
    outputs(2454) <= layer0_outputs(5540);
    outputs(2455) <= layer0_outputs(1451);
    outputs(2456) <= not(layer0_outputs(5764));
    outputs(2457) <= not(layer0_outputs(576));
    outputs(2458) <= not(layer0_outputs(779));
    outputs(2459) <= not(layer0_outputs(666));
    outputs(2460) <= not((layer0_outputs(4182)) xor (layer0_outputs(5163)));
    outputs(2461) <= (layer0_outputs(5390)) and not (layer0_outputs(3061));
    outputs(2462) <= not((layer0_outputs(493)) or (layer0_outputs(2958)));
    outputs(2463) <= not((layer0_outputs(3977)) or (layer0_outputs(2095)));
    outputs(2464) <= not(layer0_outputs(4592));
    outputs(2465) <= '1';
    outputs(2466) <= not(layer0_outputs(3530)) or (layer0_outputs(1779));
    outputs(2467) <= layer0_outputs(5749);
    outputs(2468) <= layer0_outputs(3800);
    outputs(2469) <= not((layer0_outputs(3262)) xor (layer0_outputs(1665)));
    outputs(2470) <= layer0_outputs(186);
    outputs(2471) <= (layer0_outputs(1921)) and not (layer0_outputs(2722));
    outputs(2472) <= not(layer0_outputs(7348));
    outputs(2473) <= not(layer0_outputs(4323)) or (layer0_outputs(5082));
    outputs(2474) <= not(layer0_outputs(2030));
    outputs(2475) <= (layer0_outputs(6997)) or (layer0_outputs(4576));
    outputs(2476) <= (layer0_outputs(882)) and (layer0_outputs(4190));
    outputs(2477) <= layer0_outputs(1680);
    outputs(2478) <= (layer0_outputs(4539)) xor (layer0_outputs(4527));
    outputs(2479) <= (layer0_outputs(2709)) and (layer0_outputs(3985));
    outputs(2480) <= (layer0_outputs(4278)) xor (layer0_outputs(7188));
    outputs(2481) <= (layer0_outputs(982)) xor (layer0_outputs(1400));
    outputs(2482) <= layer0_outputs(6215);
    outputs(2483) <= (layer0_outputs(3383)) or (layer0_outputs(7645));
    outputs(2484) <= not((layer0_outputs(3064)) or (layer0_outputs(6661)));
    outputs(2485) <= layer0_outputs(5693);
    outputs(2486) <= layer0_outputs(1851);
    outputs(2487) <= not((layer0_outputs(7641)) xor (layer0_outputs(233)));
    outputs(2488) <= layer0_outputs(1875);
    outputs(2489) <= layer0_outputs(1254);
    outputs(2490) <= (layer0_outputs(6977)) xor (layer0_outputs(2259));
    outputs(2491) <= not(layer0_outputs(4341));
    outputs(2492) <= not((layer0_outputs(3219)) xor (layer0_outputs(3394)));
    outputs(2493) <= not(layer0_outputs(366));
    outputs(2494) <= not(layer0_outputs(4524));
    outputs(2495) <= not(layer0_outputs(1077));
    outputs(2496) <= not(layer0_outputs(6717));
    outputs(2497) <= not((layer0_outputs(1881)) and (layer0_outputs(2109)));
    outputs(2498) <= layer0_outputs(2936);
    outputs(2499) <= not((layer0_outputs(1200)) or (layer0_outputs(2882)));
    outputs(2500) <= layer0_outputs(2829);
    outputs(2501) <= not(layer0_outputs(3723));
    outputs(2502) <= not(layer0_outputs(2051));
    outputs(2503) <= (layer0_outputs(2547)) and (layer0_outputs(1034));
    outputs(2504) <= not((layer0_outputs(5596)) and (layer0_outputs(4534)));
    outputs(2505) <= not(layer0_outputs(3464));
    outputs(2506) <= (layer0_outputs(5858)) xor (layer0_outputs(4709));
    outputs(2507) <= not(layer0_outputs(2851));
    outputs(2508) <= not((layer0_outputs(1456)) xor (layer0_outputs(3539)));
    outputs(2509) <= not(layer0_outputs(5492));
    outputs(2510) <= not(layer0_outputs(4615));
    outputs(2511) <= (layer0_outputs(4827)) xor (layer0_outputs(2872));
    outputs(2512) <= not((layer0_outputs(5552)) and (layer0_outputs(1172)));
    outputs(2513) <= layer0_outputs(7130);
    outputs(2514) <= layer0_outputs(3709);
    outputs(2515) <= layer0_outputs(2583);
    outputs(2516) <= not((layer0_outputs(1521)) xor (layer0_outputs(5004)));
    outputs(2517) <= not((layer0_outputs(3746)) xor (layer0_outputs(4114)));
    outputs(2518) <= (layer0_outputs(7391)) xor (layer0_outputs(7447));
    outputs(2519) <= layer0_outputs(7014);
    outputs(2520) <= layer0_outputs(3855);
    outputs(2521) <= not(layer0_outputs(4722)) or (layer0_outputs(2694));
    outputs(2522) <= not(layer0_outputs(1995)) or (layer0_outputs(2839));
    outputs(2523) <= layer0_outputs(2195);
    outputs(2524) <= not(layer0_outputs(4825));
    outputs(2525) <= not(layer0_outputs(4618));
    outputs(2526) <= not(layer0_outputs(5924));
    outputs(2527) <= not((layer0_outputs(6492)) xor (layer0_outputs(6065)));
    outputs(2528) <= not((layer0_outputs(5982)) xor (layer0_outputs(3354)));
    outputs(2529) <= (layer0_outputs(6866)) and (layer0_outputs(1171));
    outputs(2530) <= not(layer0_outputs(3171));
    outputs(2531) <= (layer0_outputs(2932)) or (layer0_outputs(1016));
    outputs(2532) <= not((layer0_outputs(2564)) and (layer0_outputs(421)));
    outputs(2533) <= layer0_outputs(1535);
    outputs(2534) <= layer0_outputs(490);
    outputs(2535) <= not(layer0_outputs(7582));
    outputs(2536) <= (layer0_outputs(4176)) xor (layer0_outputs(7678));
    outputs(2537) <= not(layer0_outputs(583));
    outputs(2538) <= (layer0_outputs(4466)) xor (layer0_outputs(7076));
    outputs(2539) <= '1';
    outputs(2540) <= layer0_outputs(1516);
    outputs(2541) <= layer0_outputs(6120);
    outputs(2542) <= not(layer0_outputs(5344));
    outputs(2543) <= (layer0_outputs(2045)) and not (layer0_outputs(7000));
    outputs(2544) <= not(layer0_outputs(1659));
    outputs(2545) <= layer0_outputs(6966);
    outputs(2546) <= not(layer0_outputs(5546));
    outputs(2547) <= not(layer0_outputs(7015));
    outputs(2548) <= not(layer0_outputs(2778));
    outputs(2549) <= not((layer0_outputs(3719)) and (layer0_outputs(4194)));
    outputs(2550) <= not(layer0_outputs(5539));
    outputs(2551) <= layer0_outputs(3919);
    outputs(2552) <= layer0_outputs(3609);
    outputs(2553) <= not(layer0_outputs(4799));
    outputs(2554) <= not(layer0_outputs(406)) or (layer0_outputs(1206));
    outputs(2555) <= not((layer0_outputs(6244)) xor (layer0_outputs(252)));
    outputs(2556) <= not(layer0_outputs(6547));
    outputs(2557) <= (layer0_outputs(6070)) and not (layer0_outputs(6136));
    outputs(2558) <= (layer0_outputs(3017)) and (layer0_outputs(3041));
    outputs(2559) <= layer0_outputs(4635);
    outputs(2560) <= layer0_outputs(2977);
    outputs(2561) <= (layer0_outputs(75)) xor (layer0_outputs(645));
    outputs(2562) <= not((layer0_outputs(6151)) xor (layer0_outputs(1506)));
    outputs(2563) <= not((layer0_outputs(2859)) xor (layer0_outputs(5000)));
    outputs(2564) <= not((layer0_outputs(6233)) xor (layer0_outputs(3160)));
    outputs(2565) <= not((layer0_outputs(2666)) xor (layer0_outputs(933)));
    outputs(2566) <= not(layer0_outputs(658));
    outputs(2567) <= not(layer0_outputs(6336));
    outputs(2568) <= not(layer0_outputs(6551));
    outputs(2569) <= (layer0_outputs(784)) and not (layer0_outputs(2138));
    outputs(2570) <= (layer0_outputs(465)) or (layer0_outputs(5588));
    outputs(2571) <= (layer0_outputs(4231)) and (layer0_outputs(5451));
    outputs(2572) <= layer0_outputs(4602);
    outputs(2573) <= not(layer0_outputs(4357));
    outputs(2574) <= (layer0_outputs(4158)) and not (layer0_outputs(407));
    outputs(2575) <= (layer0_outputs(2241)) xor (layer0_outputs(3306));
    outputs(2576) <= layer0_outputs(2253);
    outputs(2577) <= not(layer0_outputs(7612));
    outputs(2578) <= not(layer0_outputs(211));
    outputs(2579) <= (layer0_outputs(4629)) and not (layer0_outputs(7172));
    outputs(2580) <= not(layer0_outputs(413));
    outputs(2581) <= not(layer0_outputs(7192));
    outputs(2582) <= layer0_outputs(3515);
    outputs(2583) <= (layer0_outputs(4183)) and not (layer0_outputs(3607));
    outputs(2584) <= not((layer0_outputs(1014)) xor (layer0_outputs(3195)));
    outputs(2585) <= not(layer0_outputs(5540)) or (layer0_outputs(4135));
    outputs(2586) <= not(layer0_outputs(865));
    outputs(2587) <= layer0_outputs(2914);
    outputs(2588) <= not(layer0_outputs(6683));
    outputs(2589) <= not(layer0_outputs(3893));
    outputs(2590) <= not((layer0_outputs(744)) xor (layer0_outputs(3410)));
    outputs(2591) <= not(layer0_outputs(6876)) or (layer0_outputs(6430));
    outputs(2592) <= not(layer0_outputs(2212));
    outputs(2593) <= layer0_outputs(26);
    outputs(2594) <= not(layer0_outputs(4742));
    outputs(2595) <= not((layer0_outputs(7218)) xor (layer0_outputs(2988)));
    outputs(2596) <= (layer0_outputs(3821)) xor (layer0_outputs(6563));
    outputs(2597) <= (layer0_outputs(5598)) or (layer0_outputs(7649));
    outputs(2598) <= '1';
    outputs(2599) <= not(layer0_outputs(44));
    outputs(2600) <= not(layer0_outputs(7242));
    outputs(2601) <= not(layer0_outputs(1047));
    outputs(2602) <= not(layer0_outputs(677));
    outputs(2603) <= not(layer0_outputs(4871));
    outputs(2604) <= not((layer0_outputs(383)) xor (layer0_outputs(2891)));
    outputs(2605) <= not((layer0_outputs(7566)) xor (layer0_outputs(5083)));
    outputs(2606) <= not(layer0_outputs(3764));
    outputs(2607) <= not(layer0_outputs(1313));
    outputs(2608) <= not((layer0_outputs(4853)) and (layer0_outputs(4134)));
    outputs(2609) <= not(layer0_outputs(4459));
    outputs(2610) <= not((layer0_outputs(20)) and (layer0_outputs(4298)));
    outputs(2611) <= layer0_outputs(5737);
    outputs(2612) <= layer0_outputs(6954);
    outputs(2613) <= (layer0_outputs(3917)) and (layer0_outputs(5955));
    outputs(2614) <= not(layer0_outputs(2996));
    outputs(2615) <= not(layer0_outputs(5259)) or (layer0_outputs(3064));
    outputs(2616) <= not(layer0_outputs(6566));
    outputs(2617) <= not(layer0_outputs(1337));
    outputs(2618) <= layer0_outputs(6822);
    outputs(2619) <= not((layer0_outputs(6059)) xor (layer0_outputs(7088)));
    outputs(2620) <= not((layer0_outputs(2284)) or (layer0_outputs(6292)));
    outputs(2621) <= (layer0_outputs(2254)) and (layer0_outputs(1972));
    outputs(2622) <= '1';
    outputs(2623) <= not(layer0_outputs(3728)) or (layer0_outputs(6405));
    outputs(2624) <= layer0_outputs(7468);
    outputs(2625) <= layer0_outputs(5498);
    outputs(2626) <= layer0_outputs(4026);
    outputs(2627) <= layer0_outputs(4685);
    outputs(2628) <= layer0_outputs(5538);
    outputs(2629) <= layer0_outputs(7017);
    outputs(2630) <= not(layer0_outputs(2347));
    outputs(2631) <= not(layer0_outputs(3502));
    outputs(2632) <= not((layer0_outputs(3281)) xor (layer0_outputs(6802)));
    outputs(2633) <= layer0_outputs(2486);
    outputs(2634) <= (layer0_outputs(1635)) xor (layer0_outputs(6436));
    outputs(2635) <= not((layer0_outputs(1842)) xor (layer0_outputs(7139)));
    outputs(2636) <= layer0_outputs(7070);
    outputs(2637) <= (layer0_outputs(87)) and not (layer0_outputs(3593));
    outputs(2638) <= '0';
    outputs(2639) <= (layer0_outputs(841)) or (layer0_outputs(1700));
    outputs(2640) <= (layer0_outputs(3140)) xor (layer0_outputs(3133));
    outputs(2641) <= not(layer0_outputs(155));
    outputs(2642) <= layer0_outputs(5261);
    outputs(2643) <= (layer0_outputs(3615)) xor (layer0_outputs(3216));
    outputs(2644) <= not(layer0_outputs(6576));
    outputs(2645) <= (layer0_outputs(1710)) xor (layer0_outputs(3342));
    outputs(2646) <= not(layer0_outputs(5956));
    outputs(2647) <= layer0_outputs(6086);
    outputs(2648) <= layer0_outputs(6598);
    outputs(2649) <= not(layer0_outputs(5234)) or (layer0_outputs(6960));
    outputs(2650) <= (layer0_outputs(1858)) and (layer0_outputs(6981));
    outputs(2651) <= layer0_outputs(1093);
    outputs(2652) <= layer0_outputs(7112);
    outputs(2653) <= (layer0_outputs(891)) and not (layer0_outputs(3621));
    outputs(2654) <= not((layer0_outputs(7429)) xor (layer0_outputs(4401)));
    outputs(2655) <= not((layer0_outputs(5714)) xor (layer0_outputs(1787)));
    outputs(2656) <= not(layer0_outputs(6596));
    outputs(2657) <= layer0_outputs(5766);
    outputs(2658) <= layer0_outputs(7216);
    outputs(2659) <= layer0_outputs(5663);
    outputs(2660) <= '1';
    outputs(2661) <= not((layer0_outputs(7409)) xor (layer0_outputs(3973)));
    outputs(2662) <= not(layer0_outputs(1393));
    outputs(2663) <= not((layer0_outputs(7408)) or (layer0_outputs(3334)));
    outputs(2664) <= layer0_outputs(2463);
    outputs(2665) <= (layer0_outputs(4320)) xor (layer0_outputs(6527));
    outputs(2666) <= not((layer0_outputs(884)) xor (layer0_outputs(7210)));
    outputs(2667) <= not(layer0_outputs(6046)) or (layer0_outputs(4705));
    outputs(2668) <= (layer0_outputs(3065)) or (layer0_outputs(4217));
    outputs(2669) <= (layer0_outputs(3574)) xor (layer0_outputs(1538));
    outputs(2670) <= (layer0_outputs(174)) and not (layer0_outputs(2556));
    outputs(2671) <= layer0_outputs(3340);
    outputs(2672) <= layer0_outputs(4061);
    outputs(2673) <= (layer0_outputs(2359)) xor (layer0_outputs(4467));
    outputs(2674) <= not((layer0_outputs(3297)) xor (layer0_outputs(5447)));
    outputs(2675) <= layer0_outputs(3256);
    outputs(2676) <= layer0_outputs(6220);
    outputs(2677) <= (layer0_outputs(494)) and not (layer0_outputs(317));
    outputs(2678) <= layer0_outputs(754);
    outputs(2679) <= not((layer0_outputs(2878)) xor (layer0_outputs(7268)));
    outputs(2680) <= layer0_outputs(557);
    outputs(2681) <= not((layer0_outputs(4108)) and (layer0_outputs(4944)));
    outputs(2682) <= layer0_outputs(6052);
    outputs(2683) <= not(layer0_outputs(5206));
    outputs(2684) <= layer0_outputs(5551);
    outputs(2685) <= not(layer0_outputs(698)) or (layer0_outputs(4071));
    outputs(2686) <= not((layer0_outputs(5677)) xor (layer0_outputs(2274)));
    outputs(2687) <= (layer0_outputs(5538)) and not (layer0_outputs(6950));
    outputs(2688) <= not(layer0_outputs(1189));
    outputs(2689) <= not(layer0_outputs(4204)) or (layer0_outputs(3093));
    outputs(2690) <= layer0_outputs(6513);
    outputs(2691) <= not(layer0_outputs(2337)) or (layer0_outputs(2503));
    outputs(2692) <= layer0_outputs(3942);
    outputs(2693) <= not(layer0_outputs(2633));
    outputs(2694) <= not((layer0_outputs(3500)) xor (layer0_outputs(5520)));
    outputs(2695) <= (layer0_outputs(2230)) and not (layer0_outputs(7575));
    outputs(2696) <= not(layer0_outputs(2842));
    outputs(2697) <= layer0_outputs(2653);
    outputs(2698) <= layer0_outputs(6173);
    outputs(2699) <= not((layer0_outputs(4212)) xor (layer0_outputs(1722)));
    outputs(2700) <= not(layer0_outputs(3471));
    outputs(2701) <= (layer0_outputs(2648)) xor (layer0_outputs(1487));
    outputs(2702) <= not((layer0_outputs(6221)) xor (layer0_outputs(322)));
    outputs(2703) <= not(layer0_outputs(1500));
    outputs(2704) <= (layer0_outputs(6324)) or (layer0_outputs(237));
    outputs(2705) <= not((layer0_outputs(7371)) xor (layer0_outputs(1066)));
    outputs(2706) <= layer0_outputs(5920);
    outputs(2707) <= not(layer0_outputs(3539)) or (layer0_outputs(6979));
    outputs(2708) <= (layer0_outputs(3260)) xor (layer0_outputs(7171));
    outputs(2709) <= (layer0_outputs(4259)) and (layer0_outputs(3102));
    outputs(2710) <= (layer0_outputs(1270)) xor (layer0_outputs(2243));
    outputs(2711) <= (layer0_outputs(6863)) or (layer0_outputs(7501));
    outputs(2712) <= layer0_outputs(2495);
    outputs(2713) <= (layer0_outputs(3032)) and not (layer0_outputs(7019));
    outputs(2714) <= layer0_outputs(2010);
    outputs(2715) <= not(layer0_outputs(2899));
    outputs(2716) <= not(layer0_outputs(1606)) or (layer0_outputs(6437));
    outputs(2717) <= not((layer0_outputs(5627)) xor (layer0_outputs(5796)));
    outputs(2718) <= (layer0_outputs(3377)) xor (layer0_outputs(7645));
    outputs(2719) <= (layer0_outputs(7204)) or (layer0_outputs(4644));
    outputs(2720) <= not(layer0_outputs(6223));
    outputs(2721) <= layer0_outputs(5393);
    outputs(2722) <= (layer0_outputs(5614)) xor (layer0_outputs(4814));
    outputs(2723) <= (layer0_outputs(861)) or (layer0_outputs(7193));
    outputs(2724) <= layer0_outputs(236);
    outputs(2725) <= not((layer0_outputs(417)) xor (layer0_outputs(3681)));
    outputs(2726) <= (layer0_outputs(5490)) xor (layer0_outputs(5360));
    outputs(2727) <= not(layer0_outputs(855));
    outputs(2728) <= not(layer0_outputs(4991));
    outputs(2729) <= not(layer0_outputs(4566)) or (layer0_outputs(6538));
    outputs(2730) <= (layer0_outputs(5418)) and not (layer0_outputs(404));
    outputs(2731) <= not(layer0_outputs(4430));
    outputs(2732) <= not(layer0_outputs(918));
    outputs(2733) <= not(layer0_outputs(1446));
    outputs(2734) <= (layer0_outputs(2053)) and not (layer0_outputs(1673));
    outputs(2735) <= not((layer0_outputs(3841)) xor (layer0_outputs(2326)));
    outputs(2736) <= not(layer0_outputs(5076)) or (layer0_outputs(5634));
    outputs(2737) <= not((layer0_outputs(5824)) xor (layer0_outputs(2236)));
    outputs(2738) <= not((layer0_outputs(4880)) xor (layer0_outputs(5583)));
    outputs(2739) <= (layer0_outputs(6321)) xor (layer0_outputs(1776));
    outputs(2740) <= not((layer0_outputs(3431)) and (layer0_outputs(5352)));
    outputs(2741) <= layer0_outputs(4151);
    outputs(2742) <= not((layer0_outputs(1982)) xor (layer0_outputs(7295)));
    outputs(2743) <= (layer0_outputs(280)) xor (layer0_outputs(3469));
    outputs(2744) <= not(layer0_outputs(1256));
    outputs(2745) <= not(layer0_outputs(5617));
    outputs(2746) <= not((layer0_outputs(3429)) xor (layer0_outputs(2668)));
    outputs(2747) <= not(layer0_outputs(5410));
    outputs(2748) <= not((layer0_outputs(2582)) and (layer0_outputs(2117)));
    outputs(2749) <= layer0_outputs(564);
    outputs(2750) <= not((layer0_outputs(7076)) xor (layer0_outputs(6999)));
    outputs(2751) <= not(layer0_outputs(7041));
    outputs(2752) <= (layer0_outputs(706)) xor (layer0_outputs(3294));
    outputs(2753) <= not((layer0_outputs(6324)) xor (layer0_outputs(6101)));
    outputs(2754) <= not(layer0_outputs(1067));
    outputs(2755) <= layer0_outputs(5165);
    outputs(2756) <= (layer0_outputs(5948)) and (layer0_outputs(1028));
    outputs(2757) <= not(layer0_outputs(7403)) or (layer0_outputs(6762));
    outputs(2758) <= not(layer0_outputs(4402));
    outputs(2759) <= layer0_outputs(1822);
    outputs(2760) <= not((layer0_outputs(210)) and (layer0_outputs(3682)));
    outputs(2761) <= (layer0_outputs(1939)) and not (layer0_outputs(6410));
    outputs(2762) <= not(layer0_outputs(1443));
    outputs(2763) <= not((layer0_outputs(7083)) or (layer0_outputs(7087)));
    outputs(2764) <= layer0_outputs(5072);
    outputs(2765) <= (layer0_outputs(1651)) or (layer0_outputs(7396));
    outputs(2766) <= not((layer0_outputs(6856)) xor (layer0_outputs(2838)));
    outputs(2767) <= not((layer0_outputs(6611)) xor (layer0_outputs(203)));
    outputs(2768) <= (layer0_outputs(6578)) and not (layer0_outputs(251));
    outputs(2769) <= layer0_outputs(7352);
    outputs(2770) <= not((layer0_outputs(5617)) and (layer0_outputs(7271)));
    outputs(2771) <= layer0_outputs(6821);
    outputs(2772) <= not(layer0_outputs(3411));
    outputs(2773) <= not((layer0_outputs(927)) and (layer0_outputs(3328)));
    outputs(2774) <= (layer0_outputs(6622)) or (layer0_outputs(4728));
    outputs(2775) <= (layer0_outputs(958)) xor (layer0_outputs(5901));
    outputs(2776) <= (layer0_outputs(4656)) xor (layer0_outputs(2207));
    outputs(2777) <= (layer0_outputs(1900)) and (layer0_outputs(4624));
    outputs(2778) <= (layer0_outputs(6454)) or (layer0_outputs(1081));
    outputs(2779) <= layer0_outputs(2333);
    outputs(2780) <= not(layer0_outputs(4296));
    outputs(2781) <= not(layer0_outputs(146));
    outputs(2782) <= not((layer0_outputs(3368)) or (layer0_outputs(5556)));
    outputs(2783) <= (layer0_outputs(6048)) xor (layer0_outputs(2350));
    outputs(2784) <= not((layer0_outputs(3896)) or (layer0_outputs(2645)));
    outputs(2785) <= not(layer0_outputs(6009));
    outputs(2786) <= layer0_outputs(6378);
    outputs(2787) <= not(layer0_outputs(4042));
    outputs(2788) <= layer0_outputs(5219);
    outputs(2789) <= not((layer0_outputs(6747)) xor (layer0_outputs(1322)));
    outputs(2790) <= not(layer0_outputs(7415));
    outputs(2791) <= not(layer0_outputs(1369));
    outputs(2792) <= '0';
    outputs(2793) <= (layer0_outputs(2235)) and not (layer0_outputs(6875));
    outputs(2794) <= not(layer0_outputs(3951));
    outputs(2795) <= layer0_outputs(7132);
    outputs(2796) <= (layer0_outputs(7316)) and not (layer0_outputs(3774));
    outputs(2797) <= not(layer0_outputs(45));
    outputs(2798) <= not(layer0_outputs(60));
    outputs(2799) <= not(layer0_outputs(5093)) or (layer0_outputs(292));
    outputs(2800) <= layer0_outputs(2285);
    outputs(2801) <= (layer0_outputs(6222)) or (layer0_outputs(1362));
    outputs(2802) <= layer0_outputs(4483);
    outputs(2803) <= layer0_outputs(7554);
    outputs(2804) <= layer0_outputs(3161);
    outputs(2805) <= layer0_outputs(6138);
    outputs(2806) <= not(layer0_outputs(656));
    outputs(2807) <= not((layer0_outputs(750)) xor (layer0_outputs(3554)));
    outputs(2808) <= layer0_outputs(2486);
    outputs(2809) <= layer0_outputs(483);
    outputs(2810) <= not(layer0_outputs(5990));
    outputs(2811) <= not(layer0_outputs(4104));
    outputs(2812) <= (layer0_outputs(7531)) and not (layer0_outputs(4051));
    outputs(2813) <= not((layer0_outputs(4671)) xor (layer0_outputs(2558)));
    outputs(2814) <= (layer0_outputs(4186)) xor (layer0_outputs(3690));
    outputs(2815) <= not(layer0_outputs(5425)) or (layer0_outputs(3735));
    outputs(2816) <= layer0_outputs(2596);
    outputs(2817) <= layer0_outputs(5124);
    outputs(2818) <= layer0_outputs(3729);
    outputs(2819) <= (layer0_outputs(6953)) or (layer0_outputs(5930));
    outputs(2820) <= layer0_outputs(2508);
    outputs(2821) <= not(layer0_outputs(5048));
    outputs(2822) <= not(layer0_outputs(4595));
    outputs(2823) <= not((layer0_outputs(1558)) and (layer0_outputs(4323)));
    outputs(2824) <= not(layer0_outputs(372)) or (layer0_outputs(2432));
    outputs(2825) <= (layer0_outputs(259)) xor (layer0_outputs(4009));
    outputs(2826) <= not((layer0_outputs(1839)) xor (layer0_outputs(4923)));
    outputs(2827) <= not((layer0_outputs(1594)) xor (layer0_outputs(4084)));
    outputs(2828) <= not(layer0_outputs(4414)) or (layer0_outputs(6821));
    outputs(2829) <= layer0_outputs(5623);
    outputs(2830) <= layer0_outputs(2124);
    outputs(2831) <= not(layer0_outputs(6665));
    outputs(2832) <= (layer0_outputs(4520)) and not (layer0_outputs(3177));
    outputs(2833) <= layer0_outputs(5301);
    outputs(2834) <= (layer0_outputs(6230)) xor (layer0_outputs(934));
    outputs(2835) <= (layer0_outputs(3967)) or (layer0_outputs(6249));
    outputs(2836) <= layer0_outputs(7507);
    outputs(2837) <= layer0_outputs(2127);
    outputs(2838) <= layer0_outputs(4252);
    outputs(2839) <= not(layer0_outputs(5596));
    outputs(2840) <= layer0_outputs(4390);
    outputs(2841) <= (layer0_outputs(3980)) xor (layer0_outputs(5849));
    outputs(2842) <= not(layer0_outputs(2603));
    outputs(2843) <= (layer0_outputs(1397)) and not (layer0_outputs(4118));
    outputs(2844) <= not((layer0_outputs(3290)) xor (layer0_outputs(467)));
    outputs(2845) <= not((layer0_outputs(2282)) xor (layer0_outputs(2875)));
    outputs(2846) <= layer0_outputs(1022);
    outputs(2847) <= (layer0_outputs(4646)) xor (layer0_outputs(832));
    outputs(2848) <= not((layer0_outputs(6845)) xor (layer0_outputs(6133)));
    outputs(2849) <= not((layer0_outputs(3443)) or (layer0_outputs(515)));
    outputs(2850) <= not(layer0_outputs(5268));
    outputs(2851) <= not((layer0_outputs(6843)) xor (layer0_outputs(2280)));
    outputs(2852) <= not((layer0_outputs(2677)) and (layer0_outputs(3158)));
    outputs(2853) <= not(layer0_outputs(2831));
    outputs(2854) <= (layer0_outputs(3161)) and not (layer0_outputs(883));
    outputs(2855) <= layer0_outputs(4584);
    outputs(2856) <= not(layer0_outputs(2409));
    outputs(2857) <= not((layer0_outputs(6623)) or (layer0_outputs(3627)));
    outputs(2858) <= '1';
    outputs(2859) <= not((layer0_outputs(2752)) xor (layer0_outputs(1855)));
    outputs(2860) <= layer0_outputs(7572);
    outputs(2861) <= not((layer0_outputs(2656)) or (layer0_outputs(3571)));
    outputs(2862) <= layer0_outputs(3721);
    outputs(2863) <= (layer0_outputs(1740)) xor (layer0_outputs(7181));
    outputs(2864) <= not(layer0_outputs(1640));
    outputs(2865) <= (layer0_outputs(2631)) xor (layer0_outputs(6078));
    outputs(2866) <= not(layer0_outputs(1869)) or (layer0_outputs(1298));
    outputs(2867) <= layer0_outputs(5984);
    outputs(2868) <= not(layer0_outputs(4095));
    outputs(2869) <= not(layer0_outputs(1830));
    outputs(2870) <= (layer0_outputs(6420)) and not (layer0_outputs(5777));
    outputs(2871) <= not(layer0_outputs(7610)) or (layer0_outputs(2922));
    outputs(2872) <= (layer0_outputs(1406)) and not (layer0_outputs(6751));
    outputs(2873) <= not(layer0_outputs(3999));
    outputs(2874) <= not(layer0_outputs(611)) or (layer0_outputs(7326));
    outputs(2875) <= not(layer0_outputs(6181));
    outputs(2876) <= not(layer0_outputs(3894));
    outputs(2877) <= not(layer0_outputs(3077)) or (layer0_outputs(523));
    outputs(2878) <= not((layer0_outputs(2200)) or (layer0_outputs(4677)));
    outputs(2879) <= not(layer0_outputs(2058));
    outputs(2880) <= layer0_outputs(2657);
    outputs(2881) <= layer0_outputs(3312);
    outputs(2882) <= layer0_outputs(2388);
    outputs(2883) <= (layer0_outputs(1440)) and not (layer0_outputs(5934));
    outputs(2884) <= layer0_outputs(7490);
    outputs(2885) <= (layer0_outputs(584)) xor (layer0_outputs(768));
    outputs(2886) <= layer0_outputs(5722);
    outputs(2887) <= layer0_outputs(2652);
    outputs(2888) <= layer0_outputs(7270);
    outputs(2889) <= not((layer0_outputs(2245)) and (layer0_outputs(1225)));
    outputs(2890) <= (layer0_outputs(5298)) xor (layer0_outputs(5822));
    outputs(2891) <= (layer0_outputs(5281)) and (layer0_outputs(7235));
    outputs(2892) <= not(layer0_outputs(2786));
    outputs(2893) <= not((layer0_outputs(853)) xor (layer0_outputs(5915)));
    outputs(2894) <= not(layer0_outputs(7562)) or (layer0_outputs(1471));
    outputs(2895) <= layer0_outputs(661);
    outputs(2896) <= layer0_outputs(7007);
    outputs(2897) <= not((layer0_outputs(4591)) xor (layer0_outputs(1510)));
    outputs(2898) <= not(layer0_outputs(2622));
    outputs(2899) <= not(layer0_outputs(809));
    outputs(2900) <= (layer0_outputs(635)) xor (layer0_outputs(2100));
    outputs(2901) <= not(layer0_outputs(4734));
    outputs(2902) <= '1';
    outputs(2903) <= (layer0_outputs(836)) or (layer0_outputs(3259));
    outputs(2904) <= not(layer0_outputs(4620));
    outputs(2905) <= not(layer0_outputs(11));
    outputs(2906) <= (layer0_outputs(5368)) and not (layer0_outputs(6297));
    outputs(2907) <= not(layer0_outputs(2546));
    outputs(2908) <= not(layer0_outputs(3315));
    outputs(2909) <= not(layer0_outputs(2823));
    outputs(2910) <= not(layer0_outputs(700)) or (layer0_outputs(6808));
    outputs(2911) <= layer0_outputs(6245);
    outputs(2912) <= not((layer0_outputs(3601)) xor (layer0_outputs(3507)));
    outputs(2913) <= not((layer0_outputs(7065)) or (layer0_outputs(5512)));
    outputs(2914) <= (layer0_outputs(4887)) and not (layer0_outputs(337));
    outputs(2915) <= not((layer0_outputs(2765)) xor (layer0_outputs(2144)));
    outputs(2916) <= (layer0_outputs(4312)) and (layer0_outputs(5659));
    outputs(2917) <= not(layer0_outputs(1033));
    outputs(2918) <= not((layer0_outputs(1784)) and (layer0_outputs(4820)));
    outputs(2919) <= not(layer0_outputs(6790));
    outputs(2920) <= not(layer0_outputs(333));
    outputs(2921) <= not(layer0_outputs(2917));
    outputs(2922) <= not((layer0_outputs(313)) and (layer0_outputs(5061)));
    outputs(2923) <= not(layer0_outputs(1083));
    outputs(2924) <= not((layer0_outputs(6203)) or (layer0_outputs(2731)));
    outputs(2925) <= (layer0_outputs(6436)) or (layer0_outputs(2221));
    outputs(2926) <= not((layer0_outputs(546)) xor (layer0_outputs(7106)));
    outputs(2927) <= not(layer0_outputs(1209));
    outputs(2928) <= not(layer0_outputs(6168));
    outputs(2929) <= layer0_outputs(3582);
    outputs(2930) <= (layer0_outputs(682)) or (layer0_outputs(7589));
    outputs(2931) <= (layer0_outputs(2135)) or (layer0_outputs(854));
    outputs(2932) <= not(layer0_outputs(5348)) or (layer0_outputs(1119));
    outputs(2933) <= (layer0_outputs(742)) or (layer0_outputs(3996));
    outputs(2934) <= layer0_outputs(286);
    outputs(2935) <= layer0_outputs(2569);
    outputs(2936) <= layer0_outputs(4120);
    outputs(2937) <= not(layer0_outputs(4409)) or (layer0_outputs(2346));
    outputs(2938) <= not((layer0_outputs(3031)) and (layer0_outputs(2889)));
    outputs(2939) <= not(layer0_outputs(6338));
    outputs(2940) <= layer0_outputs(5060);
    outputs(2941) <= not((layer0_outputs(5834)) or (layer0_outputs(3849)));
    outputs(2942) <= (layer0_outputs(7503)) xor (layer0_outputs(7012));
    outputs(2943) <= not(layer0_outputs(1824));
    outputs(2944) <= layer0_outputs(481);
    outputs(2945) <= layer0_outputs(6072);
    outputs(2946) <= not(layer0_outputs(3033));
    outputs(2947) <= (layer0_outputs(6318)) and not (layer0_outputs(6621));
    outputs(2948) <= not(layer0_outputs(5119));
    outputs(2949) <= not((layer0_outputs(3133)) or (layer0_outputs(5230)));
    outputs(2950) <= not(layer0_outputs(7164));
    outputs(2951) <= not(layer0_outputs(938));
    outputs(2952) <= not(layer0_outputs(2871));
    outputs(2953) <= layer0_outputs(3116);
    outputs(2954) <= not(layer0_outputs(4838));
    outputs(2955) <= layer0_outputs(3046);
    outputs(2956) <= not(layer0_outputs(2880));
    outputs(2957) <= not(layer0_outputs(6944));
    outputs(2958) <= not(layer0_outputs(1532));
    outputs(2959) <= layer0_outputs(3594);
    outputs(2960) <= layer0_outputs(7212);
    outputs(2961) <= (layer0_outputs(1455)) xor (layer0_outputs(4491));
    outputs(2962) <= (layer0_outputs(1015)) and not (layer0_outputs(306));
    outputs(2963) <= not(layer0_outputs(5391));
    outputs(2964) <= not((layer0_outputs(501)) or (layer0_outputs(6501)));
    outputs(2965) <= layer0_outputs(7334);
    outputs(2966) <= layer0_outputs(437);
    outputs(2967) <= not((layer0_outputs(1624)) xor (layer0_outputs(7274)));
    outputs(2968) <= not(layer0_outputs(3190));
    outputs(2969) <= not(layer0_outputs(5620)) or (layer0_outputs(1604));
    outputs(2970) <= not((layer0_outputs(5606)) and (layer0_outputs(5733)));
    outputs(2971) <= not(layer0_outputs(474)) or (layer0_outputs(994));
    outputs(2972) <= not((layer0_outputs(6389)) xor (layer0_outputs(6049)));
    outputs(2973) <= not((layer0_outputs(7305)) xor (layer0_outputs(6802)));
    outputs(2974) <= not(layer0_outputs(6117));
    outputs(2975) <= layer0_outputs(1429);
    outputs(2976) <= not((layer0_outputs(2267)) xor (layer0_outputs(3753)));
    outputs(2977) <= not(layer0_outputs(5439));
    outputs(2978) <= layer0_outputs(3765);
    outputs(2979) <= not(layer0_outputs(3425));
    outputs(2980) <= layer0_outputs(1032);
    outputs(2981) <= (layer0_outputs(2071)) xor (layer0_outputs(6644));
    outputs(2982) <= layer0_outputs(5984);
    outputs(2983) <= not(layer0_outputs(5205));
    outputs(2984) <= not(layer0_outputs(6241));
    outputs(2985) <= layer0_outputs(6581);
    outputs(2986) <= not(layer0_outputs(4032));
    outputs(2987) <= not((layer0_outputs(1111)) and (layer0_outputs(6063)));
    outputs(2988) <= not(layer0_outputs(2021)) or (layer0_outputs(2742));
    outputs(2989) <= layer0_outputs(5132);
    outputs(2990) <= (layer0_outputs(5815)) and not (layer0_outputs(565));
    outputs(2991) <= layer0_outputs(2992);
    outputs(2992) <= (layer0_outputs(2477)) xor (layer0_outputs(6532));
    outputs(2993) <= not((layer0_outputs(1057)) and (layer0_outputs(2051)));
    outputs(2994) <= not((layer0_outputs(3213)) xor (layer0_outputs(2554)));
    outputs(2995) <= not((layer0_outputs(5569)) or (layer0_outputs(6053)));
    outputs(2996) <= (layer0_outputs(7031)) xor (layer0_outputs(7322));
    outputs(2997) <= layer0_outputs(398);
    outputs(2998) <= not(layer0_outputs(6480));
    outputs(2999) <= (layer0_outputs(7474)) or (layer0_outputs(3168));
    outputs(3000) <= layer0_outputs(3842);
    outputs(3001) <= not(layer0_outputs(1453));
    outputs(3002) <= layer0_outputs(6171);
    outputs(3003) <= not(layer0_outputs(1204));
    outputs(3004) <= (layer0_outputs(2609)) and not (layer0_outputs(7236));
    outputs(3005) <= not(layer0_outputs(2349));
    outputs(3006) <= not((layer0_outputs(2118)) xor (layer0_outputs(157)));
    outputs(3007) <= layer0_outputs(3585);
    outputs(3008) <= not((layer0_outputs(4267)) xor (layer0_outputs(4422)));
    outputs(3009) <= (layer0_outputs(5326)) xor (layer0_outputs(2567));
    outputs(3010) <= not(layer0_outputs(6429));
    outputs(3011) <= not(layer0_outputs(7239)) or (layer0_outputs(7275));
    outputs(3012) <= not((layer0_outputs(2855)) xor (layer0_outputs(4724)));
    outputs(3013) <= (layer0_outputs(7078)) or (layer0_outputs(2999));
    outputs(3014) <= not((layer0_outputs(3000)) xor (layer0_outputs(7671)));
    outputs(3015) <= not((layer0_outputs(6364)) and (layer0_outputs(47)));
    outputs(3016) <= layer0_outputs(6090);
    outputs(3017) <= (layer0_outputs(7153)) xor (layer0_outputs(3357));
    outputs(3018) <= not((layer0_outputs(2120)) xor (layer0_outputs(1284)));
    outputs(3019) <= not(layer0_outputs(3511));
    outputs(3020) <= not((layer0_outputs(4654)) xor (layer0_outputs(3858)));
    outputs(3021) <= not((layer0_outputs(2223)) xor (layer0_outputs(6882)));
    outputs(3022) <= not(layer0_outputs(4627));
    outputs(3023) <= (layer0_outputs(7667)) and not (layer0_outputs(6825));
    outputs(3024) <= not((layer0_outputs(1645)) xor (layer0_outputs(7224)));
    outputs(3025) <= not((layer0_outputs(409)) xor (layer0_outputs(3642)));
    outputs(3026) <= not(layer0_outputs(555));
    outputs(3027) <= (layer0_outputs(4905)) xor (layer0_outputs(6482));
    outputs(3028) <= (layer0_outputs(663)) or (layer0_outputs(559));
    outputs(3029) <= layer0_outputs(2447);
    outputs(3030) <= not((layer0_outputs(3832)) xor (layer0_outputs(5374)));
    outputs(3031) <= not((layer0_outputs(6170)) xor (layer0_outputs(7306)));
    outputs(3032) <= (layer0_outputs(2086)) xor (layer0_outputs(7461));
    outputs(3033) <= not((layer0_outputs(7518)) xor (layer0_outputs(5841)));
    outputs(3034) <= layer0_outputs(3739);
    outputs(3035) <= (layer0_outputs(2783)) and not (layer0_outputs(5014));
    outputs(3036) <= not((layer0_outputs(6707)) xor (layer0_outputs(4134)));
    outputs(3037) <= layer0_outputs(7209);
    outputs(3038) <= not(layer0_outputs(3171)) or (layer0_outputs(1207));
    outputs(3039) <= layer0_outputs(4021);
    outputs(3040) <= (layer0_outputs(200)) xor (layer0_outputs(7573));
    outputs(3041) <= (layer0_outputs(2773)) and not (layer0_outputs(4956));
    outputs(3042) <= not(layer0_outputs(4109));
    outputs(3043) <= not(layer0_outputs(5781));
    outputs(3044) <= not((layer0_outputs(180)) or (layer0_outputs(2827)));
    outputs(3045) <= not(layer0_outputs(2386));
    outputs(3046) <= not((layer0_outputs(5627)) xor (layer0_outputs(960)));
    outputs(3047) <= not((layer0_outputs(4922)) and (layer0_outputs(2624)));
    outputs(3048) <= not((layer0_outputs(6948)) xor (layer0_outputs(2081)));
    outputs(3049) <= layer0_outputs(6025);
    outputs(3050) <= not(layer0_outputs(143)) or (layer0_outputs(6931));
    outputs(3051) <= not(layer0_outputs(3401));
    outputs(3052) <= (layer0_outputs(4119)) xor (layer0_outputs(2224));
    outputs(3053) <= not(layer0_outputs(1920)) or (layer0_outputs(6598));
    outputs(3054) <= layer0_outputs(137);
    outputs(3055) <= not(layer0_outputs(7318));
    outputs(3056) <= (layer0_outputs(3776)) xor (layer0_outputs(5921));
    outputs(3057) <= not((layer0_outputs(5993)) or (layer0_outputs(237)));
    outputs(3058) <= not(layer0_outputs(5217));
    outputs(3059) <= (layer0_outputs(1514)) and not (layer0_outputs(111));
    outputs(3060) <= layer0_outputs(721);
    outputs(3061) <= layer0_outputs(1863);
    outputs(3062) <= layer0_outputs(4525);
    outputs(3063) <= not((layer0_outputs(7670)) xor (layer0_outputs(3801)));
    outputs(3064) <= (layer0_outputs(6928)) xor (layer0_outputs(5448));
    outputs(3065) <= not(layer0_outputs(2383));
    outputs(3066) <= not(layer0_outputs(1489));
    outputs(3067) <= not((layer0_outputs(5123)) xor (layer0_outputs(1721)));
    outputs(3068) <= not(layer0_outputs(4770)) or (layer0_outputs(1238));
    outputs(3069) <= not(layer0_outputs(3968));
    outputs(3070) <= not((layer0_outputs(1018)) and (layer0_outputs(6238)));
    outputs(3071) <= not(layer0_outputs(390));
    outputs(3072) <= (layer0_outputs(1409)) and not (layer0_outputs(2543));
    outputs(3073) <= layer0_outputs(4565);
    outputs(3074) <= (layer0_outputs(3213)) xor (layer0_outputs(1961));
    outputs(3075) <= not(layer0_outputs(1620));
    outputs(3076) <= not((layer0_outputs(7365)) or (layer0_outputs(6077)));
    outputs(3077) <= (layer0_outputs(1126)) xor (layer0_outputs(7660));
    outputs(3078) <= layer0_outputs(7192);
    outputs(3079) <= not(layer0_outputs(5043));
    outputs(3080) <= (layer0_outputs(3130)) xor (layer0_outputs(7513));
    outputs(3081) <= (layer0_outputs(913)) xor (layer0_outputs(4687));
    outputs(3082) <= not((layer0_outputs(6107)) xor (layer0_outputs(6234)));
    outputs(3083) <= not((layer0_outputs(5359)) xor (layer0_outputs(4640)));
    outputs(3084) <= (layer0_outputs(7265)) xor (layer0_outputs(7126));
    outputs(3085) <= not(layer0_outputs(659));
    outputs(3086) <= not((layer0_outputs(1572)) xor (layer0_outputs(4302)));
    outputs(3087) <= not((layer0_outputs(5451)) or (layer0_outputs(2717)));
    outputs(3088) <= not((layer0_outputs(1410)) xor (layer0_outputs(2000)));
    outputs(3089) <= not(layer0_outputs(732));
    outputs(3090) <= not((layer0_outputs(2211)) xor (layer0_outputs(6456)));
    outputs(3091) <= (layer0_outputs(6778)) and not (layer0_outputs(5558));
    outputs(3092) <= layer0_outputs(3621);
    outputs(3093) <= not((layer0_outputs(2374)) xor (layer0_outputs(4102)));
    outputs(3094) <= layer0_outputs(4470);
    outputs(3095) <= not((layer0_outputs(755)) and (layer0_outputs(4212)));
    outputs(3096) <= not((layer0_outputs(4015)) xor (layer0_outputs(2616)));
    outputs(3097) <= not(layer0_outputs(3898));
    outputs(3098) <= layer0_outputs(3318);
    outputs(3099) <= not((layer0_outputs(1268)) xor (layer0_outputs(4265)));
    outputs(3100) <= (layer0_outputs(6116)) xor (layer0_outputs(5452));
    outputs(3101) <= layer0_outputs(6469);
    outputs(3102) <= layer0_outputs(2890);
    outputs(3103) <= (layer0_outputs(261)) and not (layer0_outputs(6759));
    outputs(3104) <= (layer0_outputs(1463)) xor (layer0_outputs(3851));
    outputs(3105) <= (layer0_outputs(4404)) and not (layer0_outputs(2140));
    outputs(3106) <= layer0_outputs(6163);
    outputs(3107) <= not(layer0_outputs(3937)) or (layer0_outputs(5264));
    outputs(3108) <= (layer0_outputs(6610)) xor (layer0_outputs(4739));
    outputs(3109) <= not(layer0_outputs(523));
    outputs(3110) <= not((layer0_outputs(6145)) xor (layer0_outputs(6374)));
    outputs(3111) <= (layer0_outputs(6310)) xor (layer0_outputs(5603));
    outputs(3112) <= (layer0_outputs(6573)) and not (layer0_outputs(1477));
    outputs(3113) <= (layer0_outputs(2357)) xor (layer0_outputs(3750));
    outputs(3114) <= not((layer0_outputs(7026)) xor (layer0_outputs(3008)));
    outputs(3115) <= (layer0_outputs(4436)) xor (layer0_outputs(2551));
    outputs(3116) <= layer0_outputs(104);
    outputs(3117) <= not((layer0_outputs(6764)) xor (layer0_outputs(3895)));
    outputs(3118) <= not((layer0_outputs(4614)) or (layer0_outputs(1347)));
    outputs(3119) <= layer0_outputs(2937);
    outputs(3120) <= (layer0_outputs(1633)) and (layer0_outputs(2243));
    outputs(3121) <= (layer0_outputs(3836)) and (layer0_outputs(1531));
    outputs(3122) <= not((layer0_outputs(4057)) xor (layer0_outputs(2106)));
    outputs(3123) <= layer0_outputs(494);
    outputs(3124) <= not(layer0_outputs(3570));
    outputs(3125) <= (layer0_outputs(5489)) and not (layer0_outputs(521));
    outputs(3126) <= '0';
    outputs(3127) <= layer0_outputs(1623);
    outputs(3128) <= not((layer0_outputs(3888)) xor (layer0_outputs(1381)));
    outputs(3129) <= layer0_outputs(5809);
    outputs(3130) <= layer0_outputs(1533);
    outputs(3131) <= not((layer0_outputs(4601)) xor (layer0_outputs(675)));
    outputs(3132) <= not(layer0_outputs(1134));
    outputs(3133) <= not(layer0_outputs(4481));
    outputs(3134) <= not(layer0_outputs(1654));
    outputs(3135) <= layer0_outputs(4423);
    outputs(3136) <= (layer0_outputs(3271)) and not (layer0_outputs(2630));
    outputs(3137) <= layer0_outputs(27);
    outputs(3138) <= not((layer0_outputs(6289)) xor (layer0_outputs(6632)));
    outputs(3139) <= not(layer0_outputs(2741));
    outputs(3140) <= (layer0_outputs(2660)) and not (layer0_outputs(7419));
    outputs(3141) <= not(layer0_outputs(7184));
    outputs(3142) <= (layer0_outputs(51)) xor (layer0_outputs(5147));
    outputs(3143) <= (layer0_outputs(3807)) and not (layer0_outputs(2356));
    outputs(3144) <= not(layer0_outputs(1037));
    outputs(3145) <= (layer0_outputs(824)) xor (layer0_outputs(6620));
    outputs(3146) <= layer0_outputs(4593);
    outputs(3147) <= (layer0_outputs(2256)) and not (layer0_outputs(3308));
    outputs(3148) <= not((layer0_outputs(127)) xor (layer0_outputs(6991)));
    outputs(3149) <= not((layer0_outputs(6120)) or (layer0_outputs(6819)));
    outputs(3150) <= (layer0_outputs(4510)) xor (layer0_outputs(5194));
    outputs(3151) <= not(layer0_outputs(5568));
    outputs(3152) <= not((layer0_outputs(5474)) xor (layer0_outputs(4385)));
    outputs(3153) <= layer0_outputs(1577);
    outputs(3154) <= (layer0_outputs(7238)) xor (layer0_outputs(2255));
    outputs(3155) <= not((layer0_outputs(5440)) or (layer0_outputs(6405)));
    outputs(3156) <= not(layer0_outputs(4132));
    outputs(3157) <= not(layer0_outputs(1205));
    outputs(3158) <= layer0_outputs(2598);
    outputs(3159) <= layer0_outputs(1663);
    outputs(3160) <= not((layer0_outputs(1634)) xor (layer0_outputs(6576)));
    outputs(3161) <= (layer0_outputs(6531)) and (layer0_outputs(3159));
    outputs(3162) <= not((layer0_outputs(3170)) or (layer0_outputs(4533)));
    outputs(3163) <= not(layer0_outputs(3042));
    outputs(3164) <= (layer0_outputs(2497)) xor (layer0_outputs(1171));
    outputs(3165) <= not((layer0_outputs(1509)) and (layer0_outputs(1953)));
    outputs(3166) <= not((layer0_outputs(5269)) or (layer0_outputs(277)));
    outputs(3167) <= not((layer0_outputs(1565)) xor (layer0_outputs(6506)));
    outputs(3168) <= layer0_outputs(7644);
    outputs(3169) <= not(layer0_outputs(4257));
    outputs(3170) <= layer0_outputs(2561);
    outputs(3171) <= not(layer0_outputs(341));
    outputs(3172) <= (layer0_outputs(2334)) xor (layer0_outputs(3339));
    outputs(3173) <= not((layer0_outputs(5262)) xor (layer0_outputs(4484)));
    outputs(3174) <= not(layer0_outputs(7615));
    outputs(3175) <= layer0_outputs(6679);
    outputs(3176) <= not((layer0_outputs(3233)) and (layer0_outputs(7195)));
    outputs(3177) <= (layer0_outputs(5427)) and (layer0_outputs(3861));
    outputs(3178) <= layer0_outputs(3381);
    outputs(3179) <= not((layer0_outputs(6586)) or (layer0_outputs(3658)));
    outputs(3180) <= not((layer0_outputs(2285)) xor (layer0_outputs(3637)));
    outputs(3181) <= (layer0_outputs(1003)) xor (layer0_outputs(829));
    outputs(3182) <= not(layer0_outputs(1103)) or (layer0_outputs(7071));
    outputs(3183) <= not((layer0_outputs(2091)) xor (layer0_outputs(3928)));
    outputs(3184) <= not((layer0_outputs(5385)) and (layer0_outputs(4794)));
    outputs(3185) <= layer0_outputs(3236);
    outputs(3186) <= not(layer0_outputs(7516));
    outputs(3187) <= (layer0_outputs(1969)) and not (layer0_outputs(6129));
    outputs(3188) <= not((layer0_outputs(7360)) and (layer0_outputs(4192)));
    outputs(3189) <= (layer0_outputs(1460)) and (layer0_outputs(7056));
    outputs(3190) <= not(layer0_outputs(1998));
    outputs(3191) <= not(layer0_outputs(2080));
    outputs(3192) <= layer0_outputs(5155);
    outputs(3193) <= (layer0_outputs(3767)) and not (layer0_outputs(95));
    outputs(3194) <= not(layer0_outputs(6263)) or (layer0_outputs(4763));
    outputs(3195) <= layer0_outputs(2526);
    outputs(3196) <= layer0_outputs(5003);
    outputs(3197) <= not(layer0_outputs(1696));
    outputs(3198) <= not((layer0_outputs(4497)) xor (layer0_outputs(6963)));
    outputs(3199) <= (layer0_outputs(356)) and (layer0_outputs(6714));
    outputs(3200) <= not((layer0_outputs(1124)) xor (layer0_outputs(1625)));
    outputs(3201) <= (layer0_outputs(6395)) xor (layer0_outputs(3374));
    outputs(3202) <= not(layer0_outputs(4791));
    outputs(3203) <= layer0_outputs(805);
    outputs(3204) <= not((layer0_outputs(2485)) or (layer0_outputs(2601)));
    outputs(3205) <= (layer0_outputs(6962)) xor (layer0_outputs(2321));
    outputs(3206) <= (layer0_outputs(2424)) and (layer0_outputs(5650));
    outputs(3207) <= layer0_outputs(5641);
    outputs(3208) <= not(layer0_outputs(2544)) or (layer0_outputs(181));
    outputs(3209) <= not(layer0_outputs(4398));
    outputs(3210) <= (layer0_outputs(448)) and (layer0_outputs(916));
    outputs(3211) <= not((layer0_outputs(1348)) xor (layer0_outputs(4836)));
    outputs(3212) <= not(layer0_outputs(4977));
    outputs(3213) <= not((layer0_outputs(1522)) xor (layer0_outputs(4658)));
    outputs(3214) <= layer0_outputs(2646);
    outputs(3215) <= not((layer0_outputs(1358)) or (layer0_outputs(2827)));
    outputs(3216) <= not((layer0_outputs(318)) xor (layer0_outputs(3106)));
    outputs(3217) <= not(layer0_outputs(5015));
    outputs(3218) <= (layer0_outputs(6580)) xor (layer0_outputs(4411));
    outputs(3219) <= not(layer0_outputs(6615));
    outputs(3220) <= not((layer0_outputs(3945)) or (layer0_outputs(2405)));
    outputs(3221) <= layer0_outputs(5853);
    outputs(3222) <= not((layer0_outputs(2900)) or (layer0_outputs(2158)));
    outputs(3223) <= not((layer0_outputs(6470)) xor (layer0_outputs(265)));
    outputs(3224) <= layer0_outputs(5323);
    outputs(3225) <= not((layer0_outputs(4938)) xor (layer0_outputs(3071)));
    outputs(3226) <= (layer0_outputs(5771)) xor (layer0_outputs(2662));
    outputs(3227) <= (layer0_outputs(7388)) xor (layer0_outputs(4318));
    outputs(3228) <= layer0_outputs(3463);
    outputs(3229) <= layer0_outputs(3350);
    outputs(3230) <= not((layer0_outputs(80)) or (layer0_outputs(5633)));
    outputs(3231) <= not((layer0_outputs(5969)) xor (layer0_outputs(5981)));
    outputs(3232) <= not((layer0_outputs(1927)) xor (layer0_outputs(1545)));
    outputs(3233) <= '0';
    outputs(3234) <= not(layer0_outputs(7294));
    outputs(3235) <= (layer0_outputs(6223)) and not (layer0_outputs(220));
    outputs(3236) <= layer0_outputs(1020);
    outputs(3237) <= layer0_outputs(5135);
    outputs(3238) <= (layer0_outputs(2340)) and not (layer0_outputs(3708));
    outputs(3239) <= (layer0_outputs(1308)) and not (layer0_outputs(2114));
    outputs(3240) <= not(layer0_outputs(4156));
    outputs(3241) <= not((layer0_outputs(2441)) or (layer0_outputs(4446)));
    outputs(3242) <= not(layer0_outputs(4200));
    outputs(3243) <= not(layer0_outputs(6464));
    outputs(3244) <= not(layer0_outputs(4120));
    outputs(3245) <= (layer0_outputs(1407)) xor (layer0_outputs(7218));
    outputs(3246) <= layer0_outputs(3584);
    outputs(3247) <= layer0_outputs(2669);
    outputs(3248) <= (layer0_outputs(1619)) xor (layer0_outputs(5839));
    outputs(3249) <= layer0_outputs(6175);
    outputs(3250) <= not(layer0_outputs(762));
    outputs(3251) <= layer0_outputs(5177);
    outputs(3252) <= not(layer0_outputs(4961)) or (layer0_outputs(3165));
    outputs(3253) <= not((layer0_outputs(5287)) and (layer0_outputs(4881)));
    outputs(3254) <= not((layer0_outputs(1206)) xor (layer0_outputs(4899)));
    outputs(3255) <= layer0_outputs(3473);
    outputs(3256) <= not(layer0_outputs(3894));
    outputs(3257) <= not(layer0_outputs(4477)) or (layer0_outputs(4633));
    outputs(3258) <= not(layer0_outputs(2048)) or (layer0_outputs(6190));
    outputs(3259) <= (layer0_outputs(525)) and (layer0_outputs(2240));
    outputs(3260) <= layer0_outputs(4669);
    outputs(3261) <= not(layer0_outputs(7419));
    outputs(3262) <= (layer0_outputs(6092)) and not (layer0_outputs(7523));
    outputs(3263) <= not((layer0_outputs(5587)) xor (layer0_outputs(6043)));
    outputs(3264) <= (layer0_outputs(3808)) and not (layer0_outputs(1959));
    outputs(3265) <= (layer0_outputs(4256)) and not (layer0_outputs(5589));
    outputs(3266) <= (layer0_outputs(5611)) and not (layer0_outputs(2935));
    outputs(3267) <= layer0_outputs(1302);
    outputs(3268) <= not(layer0_outputs(1632));
    outputs(3269) <= (layer0_outputs(4720)) xor (layer0_outputs(2624));
    outputs(3270) <= not((layer0_outputs(6508)) or (layer0_outputs(5308)));
    outputs(3271) <= not(layer0_outputs(3305));
    outputs(3272) <= not(layer0_outputs(4444)) or (layer0_outputs(779));
    outputs(3273) <= not(layer0_outputs(45));
    outputs(3274) <= (layer0_outputs(4472)) and not (layer0_outputs(6846));
    outputs(3275) <= layer0_outputs(1498);
    outputs(3276) <= (layer0_outputs(4802)) and not (layer0_outputs(2612));
    outputs(3277) <= (layer0_outputs(1689)) and (layer0_outputs(4145));
    outputs(3278) <= (layer0_outputs(3396)) and (layer0_outputs(3003));
    outputs(3279) <= not(layer0_outputs(6695));
    outputs(3280) <= layer0_outputs(3255);
    outputs(3281) <= not(layer0_outputs(1541));
    outputs(3282) <= not((layer0_outputs(692)) xor (layer0_outputs(4416)));
    outputs(3283) <= (layer0_outputs(4720)) and not (layer0_outputs(3814));
    outputs(3284) <= layer0_outputs(879);
    outputs(3285) <= (layer0_outputs(3737)) and not (layer0_outputs(4448));
    outputs(3286) <= layer0_outputs(949);
    outputs(3287) <= (layer0_outputs(5846)) or (layer0_outputs(1492));
    outputs(3288) <= (layer0_outputs(4755)) and not (layer0_outputs(1662));
    outputs(3289) <= not(layer0_outputs(4445));
    outputs(3290) <= not(layer0_outputs(2799));
    outputs(3291) <= layer0_outputs(6841);
    outputs(3292) <= layer0_outputs(7361);
    outputs(3293) <= not((layer0_outputs(3974)) xor (layer0_outputs(5222)));
    outputs(3294) <= not(layer0_outputs(1006)) or (layer0_outputs(3104));
    outputs(3295) <= not(layer0_outputs(5366));
    outputs(3296) <= (layer0_outputs(4685)) xor (layer0_outputs(3011));
    outputs(3297) <= (layer0_outputs(4191)) and not (layer0_outputs(6474));
    outputs(3298) <= not((layer0_outputs(799)) xor (layer0_outputs(1739)));
    outputs(3299) <= not(layer0_outputs(2214));
    outputs(3300) <= (layer0_outputs(1817)) and not (layer0_outputs(7436));
    outputs(3301) <= (layer0_outputs(803)) and not (layer0_outputs(746));
    outputs(3302) <= not(layer0_outputs(3867)) or (layer0_outputs(5767));
    outputs(3303) <= (layer0_outputs(2015)) xor (layer0_outputs(7595));
    outputs(3304) <= layer0_outputs(6429);
    outputs(3305) <= not(layer0_outputs(762));
    outputs(3306) <= (layer0_outputs(3982)) and not (layer0_outputs(5834));
    outputs(3307) <= not((layer0_outputs(5807)) and (layer0_outputs(4582)));
    outputs(3308) <= (layer0_outputs(7313)) xor (layer0_outputs(3781));
    outputs(3309) <= (layer0_outputs(5012)) or (layer0_outputs(3910));
    outputs(3310) <= not(layer0_outputs(5018));
    outputs(3311) <= layer0_outputs(543);
    outputs(3312) <= layer0_outputs(4690);
    outputs(3313) <= not(layer0_outputs(1985));
    outputs(3314) <= layer0_outputs(2549);
    outputs(3315) <= not(layer0_outputs(3023)) or (layer0_outputs(1263));
    outputs(3316) <= (layer0_outputs(3555)) or (layer0_outputs(1098));
    outputs(3317) <= (layer0_outputs(3632)) and (layer0_outputs(1999));
    outputs(3318) <= (layer0_outputs(4677)) xor (layer0_outputs(4982));
    outputs(3319) <= (layer0_outputs(1087)) and not (layer0_outputs(5181));
    outputs(3320) <= (layer0_outputs(7168)) xor (layer0_outputs(6073));
    outputs(3321) <= not((layer0_outputs(6864)) xor (layer0_outputs(951)));
    outputs(3322) <= not((layer0_outputs(5169)) or (layer0_outputs(5781)));
    outputs(3323) <= layer0_outputs(7066);
    outputs(3324) <= (layer0_outputs(6466)) and not (layer0_outputs(7443));
    outputs(3325) <= not(layer0_outputs(2634));
    outputs(3326) <= not(layer0_outputs(4902)) or (layer0_outputs(1591));
    outputs(3327) <= not(layer0_outputs(1293));
    outputs(3328) <= not(layer0_outputs(5097));
    outputs(3329) <= not(layer0_outputs(397));
    outputs(3330) <= (layer0_outputs(1137)) xor (layer0_outputs(5923));
    outputs(3331) <= (layer0_outputs(6881)) xor (layer0_outputs(165));
    outputs(3332) <= not((layer0_outputs(1282)) or (layer0_outputs(1569)));
    outputs(3333) <= (layer0_outputs(239)) xor (layer0_outputs(2960));
    outputs(3334) <= not(layer0_outputs(7410)) or (layer0_outputs(1756));
    outputs(3335) <= '1';
    outputs(3336) <= (layer0_outputs(1235)) xor (layer0_outputs(981));
    outputs(3337) <= not((layer0_outputs(4698)) or (layer0_outputs(636)));
    outputs(3338) <= not(layer0_outputs(4578));
    outputs(3339) <= layer0_outputs(6894);
    outputs(3340) <= not(layer0_outputs(1748));
    outputs(3341) <= not(layer0_outputs(7667));
    outputs(3342) <= layer0_outputs(5837);
    outputs(3343) <= layer0_outputs(612);
    outputs(3344) <= (layer0_outputs(4009)) and not (layer0_outputs(3572));
    outputs(3345) <= not(layer0_outputs(2760));
    outputs(3346) <= not((layer0_outputs(7536)) or (layer0_outputs(6766)));
    outputs(3347) <= not(layer0_outputs(99));
    outputs(3348) <= (layer0_outputs(6117)) and not (layer0_outputs(3145));
    outputs(3349) <= not((layer0_outputs(2084)) xor (layer0_outputs(6026)));
    outputs(3350) <= not((layer0_outputs(3021)) or (layer0_outputs(1819)));
    outputs(3351) <= layer0_outputs(4914);
    outputs(3352) <= not((layer0_outputs(5937)) xor (layer0_outputs(413)));
    outputs(3353) <= not(layer0_outputs(4780));
    outputs(3354) <= (layer0_outputs(2823)) and not (layer0_outputs(4962));
    outputs(3355) <= layer0_outputs(6795);
    outputs(3356) <= not((layer0_outputs(6705)) or (layer0_outputs(2043)));
    outputs(3357) <= not((layer0_outputs(3599)) xor (layer0_outputs(2524)));
    outputs(3358) <= (layer0_outputs(69)) and not (layer0_outputs(561));
    outputs(3359) <= layer0_outputs(3511);
    outputs(3360) <= layer0_outputs(3109);
    outputs(3361) <= (layer0_outputs(3131)) and not (layer0_outputs(2514));
    outputs(3362) <= (layer0_outputs(6828)) and not (layer0_outputs(5744));
    outputs(3363) <= (layer0_outputs(875)) xor (layer0_outputs(6798));
    outputs(3364) <= not((layer0_outputs(2958)) and (layer0_outputs(230)));
    outputs(3365) <= '0';
    outputs(3366) <= (layer0_outputs(1038)) xor (layer0_outputs(457));
    outputs(3367) <= layer0_outputs(1982);
    outputs(3368) <= not(layer0_outputs(6289));
    outputs(3369) <= not((layer0_outputs(6508)) xor (layer0_outputs(67)));
    outputs(3370) <= not(layer0_outputs(102));
    outputs(3371) <= layer0_outputs(5942);
    outputs(3372) <= not(layer0_outputs(7407));
    outputs(3373) <= not(layer0_outputs(6744));
    outputs(3374) <= (layer0_outputs(4628)) xor (layer0_outputs(3157));
    outputs(3375) <= (layer0_outputs(2816)) xor (layer0_outputs(6104));
    outputs(3376) <= not(layer0_outputs(2981)) or (layer0_outputs(6905));
    outputs(3377) <= layer0_outputs(7051);
    outputs(3378) <= layer0_outputs(274);
    outputs(3379) <= not(layer0_outputs(307));
    outputs(3380) <= not(layer0_outputs(221));
    outputs(3381) <= not(layer0_outputs(1546));
    outputs(3382) <= (layer0_outputs(6306)) and (layer0_outputs(7286));
    outputs(3383) <= not((layer0_outputs(6079)) xor (layer0_outputs(2506)));
    outputs(3384) <= (layer0_outputs(3377)) and not (layer0_outputs(1425));
    outputs(3385) <= layer0_outputs(3753);
    outputs(3386) <= (layer0_outputs(4717)) xor (layer0_outputs(815));
    outputs(3387) <= not(layer0_outputs(1414)) or (layer0_outputs(3528));
    outputs(3388) <= not((layer0_outputs(1244)) xor (layer0_outputs(7498)));
    outputs(3389) <= not((layer0_outputs(5449)) xor (layer0_outputs(1333)));
    outputs(3390) <= not(layer0_outputs(1821));
    outputs(3391) <= not(layer0_outputs(5109));
    outputs(3392) <= layer0_outputs(7101);
    outputs(3393) <= layer0_outputs(2772);
    outputs(3394) <= not((layer0_outputs(1987)) and (layer0_outputs(7642)));
    outputs(3395) <= not((layer0_outputs(2101)) xor (layer0_outputs(3554)));
    outputs(3396) <= (layer0_outputs(1257)) xor (layer0_outputs(2072));
    outputs(3397) <= layer0_outputs(1381);
    outputs(3398) <= (layer0_outputs(6945)) and not (layer0_outputs(6024));
    outputs(3399) <= (layer0_outputs(6853)) xor (layer0_outputs(266));
    outputs(3400) <= (layer0_outputs(1516)) and not (layer0_outputs(7488));
    outputs(3401) <= layer0_outputs(5056);
    outputs(3402) <= not((layer0_outputs(4763)) xor (layer0_outputs(4455)));
    outputs(3403) <= layer0_outputs(2919);
    outputs(3404) <= not((layer0_outputs(3390)) or (layer0_outputs(4000)));
    outputs(3405) <= (layer0_outputs(149)) xor (layer0_outputs(7481));
    outputs(3406) <= not(layer0_outputs(4951));
    outputs(3407) <= not(layer0_outputs(5609));
    outputs(3408) <= not(layer0_outputs(1978));
    outputs(3409) <= (layer0_outputs(4751)) xor (layer0_outputs(489));
    outputs(3410) <= layer0_outputs(1237);
    outputs(3411) <= layer0_outputs(714);
    outputs(3412) <= (layer0_outputs(893)) xor (layer0_outputs(3435));
    outputs(3413) <= not(layer0_outputs(4346));
    outputs(3414) <= (layer0_outputs(5419)) and (layer0_outputs(1847));
    outputs(3415) <= layer0_outputs(2944);
    outputs(3416) <= not(layer0_outputs(1741));
    outputs(3417) <= not(layer0_outputs(1310));
    outputs(3418) <= layer0_outputs(1790);
    outputs(3419) <= (layer0_outputs(5077)) xor (layer0_outputs(1941));
    outputs(3420) <= (layer0_outputs(5725)) xor (layer0_outputs(2494));
    outputs(3421) <= not((layer0_outputs(2326)) and (layer0_outputs(3749)));
    outputs(3422) <= not(layer0_outputs(2237));
    outputs(3423) <= layer0_outputs(1557);
    outputs(3424) <= (layer0_outputs(7203)) or (layer0_outputs(7654));
    outputs(3425) <= not(layer0_outputs(2103));
    outputs(3426) <= (layer0_outputs(2938)) and not (layer0_outputs(199));
    outputs(3427) <= layer0_outputs(2894);
    outputs(3428) <= (layer0_outputs(3639)) and not (layer0_outputs(7281));
    outputs(3429) <= layer0_outputs(2606);
    outputs(3430) <= (layer0_outputs(3745)) xor (layer0_outputs(5007));
    outputs(3431) <= not((layer0_outputs(7342)) or (layer0_outputs(4940)));
    outputs(3432) <= (layer0_outputs(2825)) xor (layer0_outputs(3916));
    outputs(3433) <= not(layer0_outputs(2959));
    outputs(3434) <= not(layer0_outputs(6955));
    outputs(3435) <= not(layer0_outputs(4977));
    outputs(3436) <= not(layer0_outputs(4870));
    outputs(3437) <= not((layer0_outputs(2897)) xor (layer0_outputs(263)));
    outputs(3438) <= not(layer0_outputs(7660));
    outputs(3439) <= not(layer0_outputs(608));
    outputs(3440) <= layer0_outputs(4722);
    outputs(3441) <= not(layer0_outputs(4164));
    outputs(3442) <= not((layer0_outputs(7262)) or (layer0_outputs(3293)));
    outputs(3443) <= not((layer0_outputs(7471)) xor (layer0_outputs(6801)));
    outputs(3444) <= not(layer0_outputs(3124));
    outputs(3445) <= not((layer0_outputs(5013)) xor (layer0_outputs(6027)));
    outputs(3446) <= not(layer0_outputs(3326));
    outputs(3447) <= not(layer0_outputs(1620));
    outputs(3448) <= (layer0_outputs(4682)) xor (layer0_outputs(3527));
    outputs(3449) <= (layer0_outputs(4352)) and not (layer0_outputs(1300));
    outputs(3450) <= layer0_outputs(7016);
    outputs(3451) <= not(layer0_outputs(1241));
    outputs(3452) <= not(layer0_outputs(5404)) or (layer0_outputs(832));
    outputs(3453) <= (layer0_outputs(7390)) and not (layer0_outputs(4948));
    outputs(3454) <= layer0_outputs(6219);
    outputs(3455) <= not(layer0_outputs(769));
    outputs(3456) <= not(layer0_outputs(2065));
    outputs(3457) <= layer0_outputs(1828);
    outputs(3458) <= layer0_outputs(7017);
    outputs(3459) <= layer0_outputs(4320);
    outputs(3460) <= not(layer0_outputs(5465)) or (layer0_outputs(3725));
    outputs(3461) <= not(layer0_outputs(2190));
    outputs(3462) <= (layer0_outputs(6305)) and (layer0_outputs(304));
    outputs(3463) <= not((layer0_outputs(5813)) xor (layer0_outputs(5053)));
    outputs(3464) <= (layer0_outputs(1968)) and (layer0_outputs(2528));
    outputs(3465) <= layer0_outputs(3963);
    outputs(3466) <= layer0_outputs(1775);
    outputs(3467) <= not((layer0_outputs(1295)) xor (layer0_outputs(5202)));
    outputs(3468) <= layer0_outputs(1882);
    outputs(3469) <= not(layer0_outputs(6914));
    outputs(3470) <= not((layer0_outputs(4746)) or (layer0_outputs(377)));
    outputs(3471) <= (layer0_outputs(6777)) and not (layer0_outputs(2965));
    outputs(3472) <= not((layer0_outputs(7550)) xor (layer0_outputs(3412)));
    outputs(3473) <= (layer0_outputs(1247)) xor (layer0_outputs(4970));
    outputs(3474) <= layer0_outputs(942);
    outputs(3475) <= (layer0_outputs(3761)) and not (layer0_outputs(216));
    outputs(3476) <= layer0_outputs(3025);
    outputs(3477) <= not(layer0_outputs(6780));
    outputs(3478) <= not(layer0_outputs(6188));
    outputs(3479) <= layer0_outputs(6259);
    outputs(3480) <= layer0_outputs(5594);
    outputs(3481) <= not(layer0_outputs(4973));
    outputs(3482) <= not(layer0_outputs(6532));
    outputs(3483) <= not((layer0_outputs(6956)) xor (layer0_outputs(1918)));
    outputs(3484) <= (layer0_outputs(55)) or (layer0_outputs(3470));
    outputs(3485) <= not(layer0_outputs(726));
    outputs(3486) <= (layer0_outputs(312)) and (layer0_outputs(2260));
    outputs(3487) <= not(layer0_outputs(1504));
    outputs(3488) <= (layer0_outputs(1578)) xor (layer0_outputs(7529));
    outputs(3489) <= layer0_outputs(5934);
    outputs(3490) <= not(layer0_outputs(1121));
    outputs(3491) <= not((layer0_outputs(6830)) or (layer0_outputs(6199)));
    outputs(3492) <= (layer0_outputs(6306)) and not (layer0_outputs(94));
    outputs(3493) <= not((layer0_outputs(7653)) xor (layer0_outputs(7248)));
    outputs(3494) <= layer0_outputs(3462);
    outputs(3495) <= (layer0_outputs(3955)) and not (layer0_outputs(2754));
    outputs(3496) <= not(layer0_outputs(1550));
    outputs(3497) <= (layer0_outputs(2356)) xor (layer0_outputs(2601));
    outputs(3498) <= (layer0_outputs(1527)) xor (layer0_outputs(5613));
    outputs(3499) <= not((layer0_outputs(4149)) xor (layer0_outputs(4824)));
    outputs(3500) <= not((layer0_outputs(7133)) xor (layer0_outputs(5471)));
    outputs(3501) <= (layer0_outputs(393)) xor (layer0_outputs(6573));
    outputs(3502) <= (layer0_outputs(5967)) xor (layer0_outputs(7225));
    outputs(3503) <= (layer0_outputs(3135)) and not (layer0_outputs(6371));
    outputs(3504) <= layer0_outputs(82);
    outputs(3505) <= (layer0_outputs(1416)) xor (layer0_outputs(4171));
    outputs(3506) <= (layer0_outputs(3552)) and not (layer0_outputs(7586));
    outputs(3507) <= layer0_outputs(3134);
    outputs(3508) <= not((layer0_outputs(3437)) xor (layer0_outputs(5884)));
    outputs(3509) <= not(layer0_outputs(5188)) or (layer0_outputs(3374));
    outputs(3510) <= layer0_outputs(5029);
    outputs(3511) <= not(layer0_outputs(7135));
    outputs(3512) <= (layer0_outputs(3532)) and not (layer0_outputs(255));
    outputs(3513) <= (layer0_outputs(6074)) and (layer0_outputs(6064));
    outputs(3514) <= not((layer0_outputs(1372)) xor (layer0_outputs(4090)));
    outputs(3515) <= layer0_outputs(354);
    outputs(3516) <= (layer0_outputs(2449)) and (layer0_outputs(838));
    outputs(3517) <= not(layer0_outputs(6271));
    outputs(3518) <= not(layer0_outputs(967));
    outputs(3519) <= (layer0_outputs(5828)) xor (layer0_outputs(473));
    outputs(3520) <= (layer0_outputs(5837)) and not (layer0_outputs(7389));
    outputs(3521) <= not((layer0_outputs(2698)) or (layer0_outputs(3466)));
    outputs(3522) <= layer0_outputs(2219);
    outputs(3523) <= not(layer0_outputs(629));
    outputs(3524) <= not((layer0_outputs(5189)) xor (layer0_outputs(6335)));
    outputs(3525) <= not(layer0_outputs(152));
    outputs(3526) <= (layer0_outputs(3665)) and not (layer0_outputs(2640));
    outputs(3527) <= not(layer0_outputs(5827));
    outputs(3528) <= not(layer0_outputs(1895));
    outputs(3529) <= not((layer0_outputs(6308)) xor (layer0_outputs(3809)));
    outputs(3530) <= not(layer0_outputs(3534));
    outputs(3531) <= not(layer0_outputs(5977));
    outputs(3532) <= layer0_outputs(2416);
    outputs(3533) <= layer0_outputs(6278);
    outputs(3534) <= not((layer0_outputs(2357)) or (layer0_outputs(2316)));
    outputs(3535) <= (layer0_outputs(976)) and not (layer0_outputs(6723));
    outputs(3536) <= (layer0_outputs(7575)) and not (layer0_outputs(4606));
    outputs(3537) <= (layer0_outputs(5038)) or (layer0_outputs(5628));
    outputs(3538) <= (layer0_outputs(7021)) xor (layer0_outputs(7179));
    outputs(3539) <= layer0_outputs(395);
    outputs(3540) <= (layer0_outputs(5183)) xor (layer0_outputs(3124));
    outputs(3541) <= (layer0_outputs(6395)) and not (layer0_outputs(4282));
    outputs(3542) <= (layer0_outputs(970)) and not (layer0_outputs(1908));
    outputs(3543) <= not(layer0_outputs(5629));
    outputs(3544) <= not((layer0_outputs(2517)) xor (layer0_outputs(2888)));
    outputs(3545) <= not((layer0_outputs(4149)) xor (layer0_outputs(5666)));
    outputs(3546) <= not((layer0_outputs(4073)) and (layer0_outputs(2090)));
    outputs(3547) <= (layer0_outputs(5546)) xor (layer0_outputs(3544));
    outputs(3548) <= not((layer0_outputs(2269)) xor (layer0_outputs(3332)));
    outputs(3549) <= not(layer0_outputs(5123));
    outputs(3550) <= not(layer0_outputs(6744));
    outputs(3551) <= (layer0_outputs(5491)) xor (layer0_outputs(6621));
    outputs(3552) <= not(layer0_outputs(7120));
    outputs(3553) <= (layer0_outputs(4254)) and (layer0_outputs(1811));
    outputs(3554) <= (layer0_outputs(344)) and not (layer0_outputs(6137));
    outputs(3555) <= not(layer0_outputs(1385));
    outputs(3556) <= layer0_outputs(5830);
    outputs(3557) <= not(layer0_outputs(5015));
    outputs(3558) <= layer0_outputs(1340);
    outputs(3559) <= (layer0_outputs(76)) and not (layer0_outputs(4748));
    outputs(3560) <= not(layer0_outputs(102));
    outputs(3561) <= layer0_outputs(4846);
    outputs(3562) <= (layer0_outputs(960)) xor (layer0_outputs(3960));
    outputs(3563) <= not(layer0_outputs(7402));
    outputs(3564) <= not((layer0_outputs(773)) or (layer0_outputs(4144)));
    outputs(3565) <= not(layer0_outputs(6978)) or (layer0_outputs(5676));
    outputs(3566) <= layer0_outputs(2203);
    outputs(3567) <= not(layer0_outputs(3027));
    outputs(3568) <= not(layer0_outputs(5929));
    outputs(3569) <= (layer0_outputs(1815)) xor (layer0_outputs(1102));
    outputs(3570) <= not((layer0_outputs(6778)) xor (layer0_outputs(6638)));
    outputs(3571) <= not((layer0_outputs(6462)) or (layer0_outputs(5930)));
    outputs(3572) <= layer0_outputs(395);
    outputs(3573) <= not(layer0_outputs(1166));
    outputs(3574) <= not(layer0_outputs(6868));
    outputs(3575) <= layer0_outputs(6956);
    outputs(3576) <= not((layer0_outputs(7646)) xor (layer0_outputs(3070)));
    outputs(3577) <= layer0_outputs(1073);
    outputs(3578) <= not(layer0_outputs(3521));
    outputs(3579) <= (layer0_outputs(897)) xor (layer0_outputs(655));
    outputs(3580) <= (layer0_outputs(2987)) and (layer0_outputs(1096));
    outputs(3581) <= layer0_outputs(5055);
    outputs(3582) <= not(layer0_outputs(1486));
    outputs(3583) <= not(layer0_outputs(3039));
    outputs(3584) <= (layer0_outputs(7434)) and not (layer0_outputs(5505));
    outputs(3585) <= not(layer0_outputs(7114)) or (layer0_outputs(655));
    outputs(3586) <= not((layer0_outputs(2552)) xor (layer0_outputs(1725)));
    outputs(3587) <= (layer0_outputs(3882)) and not (layer0_outputs(1737));
    outputs(3588) <= (layer0_outputs(5760)) xor (layer0_outputs(576));
    outputs(3589) <= (layer0_outputs(7309)) xor (layer0_outputs(1472));
    outputs(3590) <= (layer0_outputs(6905)) and not (layer0_outputs(6819));
    outputs(3591) <= not((layer0_outputs(7459)) xor (layer0_outputs(5657)));
    outputs(3592) <= (layer0_outputs(5078)) and not (layer0_outputs(6446));
    outputs(3593) <= layer0_outputs(407);
    outputs(3594) <= not((layer0_outputs(6020)) or (layer0_outputs(2480)));
    outputs(3595) <= (layer0_outputs(6525)) xor (layer0_outputs(1475));
    outputs(3596) <= (layer0_outputs(3584)) xor (layer0_outputs(2954));
    outputs(3597) <= layer0_outputs(7632);
    outputs(3598) <= '0';
    outputs(3599) <= layer0_outputs(183);
    outputs(3600) <= (layer0_outputs(4197)) and (layer0_outputs(2975));
    outputs(3601) <= layer0_outputs(6870);
    outputs(3602) <= layer0_outputs(5245);
    outputs(3603) <= (layer0_outputs(5266)) and not (layer0_outputs(5273));
    outputs(3604) <= (layer0_outputs(7093)) and not (layer0_outputs(6296));
    outputs(3605) <= layer0_outputs(4170);
    outputs(3606) <= (layer0_outputs(117)) xor (layer0_outputs(6418));
    outputs(3607) <= (layer0_outputs(1452)) xor (layer0_outputs(1891));
    outputs(3608) <= not(layer0_outputs(3536));
    outputs(3609) <= not(layer0_outputs(1399));
    outputs(3610) <= not(layer0_outputs(6114));
    outputs(3611) <= not(layer0_outputs(966));
    outputs(3612) <= not((layer0_outputs(4261)) xor (layer0_outputs(3160)));
    outputs(3613) <= not((layer0_outputs(5203)) xor (layer0_outputs(7534)));
    outputs(3614) <= not(layer0_outputs(2837));
    outputs(3615) <= not(layer0_outputs(765));
    outputs(3616) <= not(layer0_outputs(6935));
    outputs(3617) <= not(layer0_outputs(2585));
    outputs(3618) <= '1';
    outputs(3619) <= layer0_outputs(1319);
    outputs(3620) <= not(layer0_outputs(1442));
    outputs(3621) <= layer0_outputs(2052);
    outputs(3622) <= not(layer0_outputs(6965)) or (layer0_outputs(2057));
    outputs(3623) <= layer0_outputs(3243);
    outputs(3624) <= not(layer0_outputs(4386));
    outputs(3625) <= not((layer0_outputs(2853)) or (layer0_outputs(1576)));
    outputs(3626) <= not(layer0_outputs(7474));
    outputs(3627) <= not((layer0_outputs(7229)) xor (layer0_outputs(4555)));
    outputs(3628) <= (layer0_outputs(4900)) xor (layer0_outputs(4771));
    outputs(3629) <= (layer0_outputs(2556)) xor (layer0_outputs(6672));
    outputs(3630) <= not((layer0_outputs(4177)) xor (layer0_outputs(4419)));
    outputs(3631) <= not(layer0_outputs(6442));
    outputs(3632) <= (layer0_outputs(1827)) xor (layer0_outputs(5285));
    outputs(3633) <= (layer0_outputs(319)) and not (layer0_outputs(1538));
    outputs(3634) <= (layer0_outputs(702)) xor (layer0_outputs(2047));
    outputs(3635) <= not(layer0_outputs(3338));
    outputs(3636) <= not(layer0_outputs(5586));
    outputs(3637) <= (layer0_outputs(6614)) and not (layer0_outputs(1191));
    outputs(3638) <= layer0_outputs(5437);
    outputs(3639) <= (layer0_outputs(3773)) and (layer0_outputs(5536));
    outputs(3640) <= (layer0_outputs(5532)) and (layer0_outputs(3711));
    outputs(3641) <= layer0_outputs(185);
    outputs(3642) <= layer0_outputs(4657);
    outputs(3643) <= not((layer0_outputs(2093)) xor (layer0_outputs(195)));
    outputs(3644) <= layer0_outputs(2491);
    outputs(3645) <= (layer0_outputs(5698)) and not (layer0_outputs(5153));
    outputs(3646) <= not((layer0_outputs(4358)) or (layer0_outputs(1069)));
    outputs(3647) <= (layer0_outputs(5468)) and (layer0_outputs(476));
    outputs(3648) <= not((layer0_outputs(6447)) and (layer0_outputs(1095)));
    outputs(3649) <= not(layer0_outputs(2710));
    outputs(3650) <= not(layer0_outputs(588)) or (layer0_outputs(5046));
    outputs(3651) <= not(layer0_outputs(4534));
    outputs(3652) <= layer0_outputs(4553);
    outputs(3653) <= not((layer0_outputs(6663)) xor (layer0_outputs(3279)));
    outputs(3654) <= (layer0_outputs(1940)) and (layer0_outputs(4119));
    outputs(3655) <= not(layer0_outputs(6037));
    outputs(3656) <= not(layer0_outputs(7601));
    outputs(3657) <= (layer0_outputs(6558)) xor (layer0_outputs(2850));
    outputs(3658) <= (layer0_outputs(2440)) and not (layer0_outputs(7631));
    outputs(3659) <= layer0_outputs(1512);
    outputs(3660) <= (layer0_outputs(1971)) and (layer0_outputs(3728));
    outputs(3661) <= layer0_outputs(3454);
    outputs(3662) <= layer0_outputs(3331);
    outputs(3663) <= not((layer0_outputs(6275)) xor (layer0_outputs(2765)));
    outputs(3664) <= not((layer0_outputs(1345)) or (layer0_outputs(3386)));
    outputs(3665) <= (layer0_outputs(7512)) and (layer0_outputs(5785));
    outputs(3666) <= not(layer0_outputs(4858));
    outputs(3667) <= (layer0_outputs(2766)) and not (layer0_outputs(3513));
    outputs(3668) <= layer0_outputs(5193);
    outputs(3669) <= not(layer0_outputs(4842));
    outputs(3670) <= not(layer0_outputs(6916));
    outputs(3671) <= layer0_outputs(5106);
    outputs(3672) <= layer0_outputs(4213);
    outputs(3673) <= (layer0_outputs(2573)) xor (layer0_outputs(1862));
    outputs(3674) <= (layer0_outputs(440)) and not (layer0_outputs(4321));
    outputs(3675) <= '0';
    outputs(3676) <= (layer0_outputs(5840)) and not (layer0_outputs(2760));
    outputs(3677) <= layer0_outputs(863);
    outputs(3678) <= layer0_outputs(1581);
    outputs(3679) <= layer0_outputs(353);
    outputs(3680) <= not((layer0_outputs(7122)) or (layer0_outputs(3048)));
    outputs(3681) <= (layer0_outputs(849)) xor (layer0_outputs(3994));
    outputs(3682) <= layer0_outputs(3784);
    outputs(3683) <= layer0_outputs(4269);
    outputs(3684) <= layer0_outputs(5236);
    outputs(3685) <= not((layer0_outputs(826)) or (layer0_outputs(6139)));
    outputs(3686) <= (layer0_outputs(7313)) and not (layer0_outputs(7001));
    outputs(3687) <= not(layer0_outputs(983));
    outputs(3688) <= (layer0_outputs(4456)) and not (layer0_outputs(3703));
    outputs(3689) <= not(layer0_outputs(5593));
    outputs(3690) <= (layer0_outputs(1794)) and not (layer0_outputs(390));
    outputs(3691) <= not(layer0_outputs(6783));
    outputs(3692) <= layer0_outputs(2260);
    outputs(3693) <= (layer0_outputs(6859)) xor (layer0_outputs(738));
    outputs(3694) <= layer0_outputs(3331);
    outputs(3695) <= not((layer0_outputs(6578)) xor (layer0_outputs(1173)));
    outputs(3696) <= (layer0_outputs(7462)) xor (layer0_outputs(3548));
    outputs(3697) <= not(layer0_outputs(3198));
    outputs(3698) <= layer0_outputs(6337);
    outputs(3699) <= layer0_outputs(3128);
    outputs(3700) <= not((layer0_outputs(2801)) or (layer0_outputs(2301)));
    outputs(3701) <= layer0_outputs(6720);
    outputs(3702) <= not(layer0_outputs(4437));
    outputs(3703) <= not(layer0_outputs(7128));
    outputs(3704) <= (layer0_outputs(6545)) and not (layer0_outputs(4377));
    outputs(3705) <= not((layer0_outputs(4005)) xor (layer0_outputs(5407)));
    outputs(3706) <= (layer0_outputs(4394)) or (layer0_outputs(3020));
    outputs(3707) <= layer0_outputs(5394);
    outputs(3708) <= not(layer0_outputs(3229));
    outputs(3709) <= not(layer0_outputs(7022));
    outputs(3710) <= (layer0_outputs(6628)) xor (layer0_outputs(772));
    outputs(3711) <= not((layer0_outputs(3743)) xor (layer0_outputs(4276)));
    outputs(3712) <= (layer0_outputs(674)) xor (layer0_outputs(7159));
    outputs(3713) <= not(layer0_outputs(4020));
    outputs(3714) <= layer0_outputs(5087);
    outputs(3715) <= not(layer0_outputs(7120));
    outputs(3716) <= not(layer0_outputs(587));
    outputs(3717) <= not(layer0_outputs(4201)) or (layer0_outputs(1752));
    outputs(3718) <= not(layer0_outputs(6236));
    outputs(3719) <= not(layer0_outputs(4458)) or (layer0_outputs(6530));
    outputs(3720) <= not((layer0_outputs(2130)) xor (layer0_outputs(6509)));
    outputs(3721) <= layer0_outputs(6297);
    outputs(3722) <= (layer0_outputs(6360)) xor (layer0_outputs(6441));
    outputs(3723) <= not(layer0_outputs(7127));
    outputs(3724) <= layer0_outputs(5185);
    outputs(3725) <= not((layer0_outputs(7498)) and (layer0_outputs(7417)));
    outputs(3726) <= layer0_outputs(6161);
    outputs(3727) <= (layer0_outputs(1011)) xor (layer0_outputs(7183));
    outputs(3728) <= not(layer0_outputs(2261));
    outputs(3729) <= not(layer0_outputs(810));
    outputs(3730) <= not((layer0_outputs(1605)) or (layer0_outputs(7593)));
    outputs(3731) <= not(layer0_outputs(5178));
    outputs(3732) <= (layer0_outputs(4165)) xor (layer0_outputs(5104));
    outputs(3733) <= (layer0_outputs(904)) or (layer0_outputs(6335));
    outputs(3734) <= layer0_outputs(3932);
    outputs(3735) <= (layer0_outputs(4435)) xor (layer0_outputs(3738));
    outputs(3736) <= not(layer0_outputs(5411)) or (layer0_outputs(3228));
    outputs(3737) <= not(layer0_outputs(5005));
    outputs(3738) <= not((layer0_outputs(5141)) and (layer0_outputs(2339)));
    outputs(3739) <= not(layer0_outputs(7145));
    outputs(3740) <= not((layer0_outputs(1178)) xor (layer0_outputs(718)));
    outputs(3741) <= (layer0_outputs(6166)) and not (layer0_outputs(4896));
    outputs(3742) <= layer0_outputs(6499);
    outputs(3743) <= not((layer0_outputs(5377)) xor (layer0_outputs(3543)));
    outputs(3744) <= layer0_outputs(3708);
    outputs(3745) <= not((layer0_outputs(2562)) or (layer0_outputs(4010)));
    outputs(3746) <= (layer0_outputs(241)) and not (layer0_outputs(6352));
    outputs(3747) <= layer0_outputs(7666);
    outputs(3748) <= not(layer0_outputs(424));
    outputs(3749) <= layer0_outputs(5002);
    outputs(3750) <= (layer0_outputs(1059)) xor (layer0_outputs(6923));
    outputs(3751) <= layer0_outputs(2471);
    outputs(3752) <= (layer0_outputs(297)) and (layer0_outputs(1148));
    outputs(3753) <= not(layer0_outputs(1278));
    outputs(3754) <= (layer0_outputs(356)) and (layer0_outputs(5652));
    outputs(3755) <= not(layer0_outputs(4414));
    outputs(3756) <= not((layer0_outputs(7355)) xor (layer0_outputs(1146)));
    outputs(3757) <= (layer0_outputs(3164)) xor (layer0_outputs(2749));
    outputs(3758) <= (layer0_outputs(3245)) and not (layer0_outputs(3447));
    outputs(3759) <= layer0_outputs(5727);
    outputs(3760) <= not(layer0_outputs(1089));
    outputs(3761) <= (layer0_outputs(144)) xor (layer0_outputs(2715));
    outputs(3762) <= (layer0_outputs(4195)) and not (layer0_outputs(39));
    outputs(3763) <= layer0_outputs(3987);
    outputs(3764) <= not(layer0_outputs(2265));
    outputs(3765) <= not((layer0_outputs(6920)) or (layer0_outputs(4936)));
    outputs(3766) <= (layer0_outputs(5592)) and not (layer0_outputs(3063));
    outputs(3767) <= (layer0_outputs(5718)) and (layer0_outputs(1990));
    outputs(3768) <= (layer0_outputs(1235)) and not (layer0_outputs(6378));
    outputs(3769) <= (layer0_outputs(1823)) xor (layer0_outputs(1902));
    outputs(3770) <= not((layer0_outputs(3822)) xor (layer0_outputs(1840)));
    outputs(3771) <= not(layer0_outputs(5116));
    outputs(3772) <= not(layer0_outputs(1390));
    outputs(3773) <= (layer0_outputs(3952)) xor (layer0_outputs(1344));
    outputs(3774) <= (layer0_outputs(4541)) and (layer0_outputs(2902));
    outputs(3775) <= (layer0_outputs(2183)) xor (layer0_outputs(3829));
    outputs(3776) <= not((layer0_outputs(5919)) xor (layer0_outputs(4748)));
    outputs(3777) <= not((layer0_outputs(2649)) or (layer0_outputs(4363)));
    outputs(3778) <= '0';
    outputs(3779) <= (layer0_outputs(227)) xor (layer0_outputs(4335));
    outputs(3780) <= layer0_outputs(1052);
    outputs(3781) <= (layer0_outputs(6936)) and not (layer0_outputs(4131));
    outputs(3782) <= (layer0_outputs(5523)) xor (layer0_outputs(4872));
    outputs(3783) <= not(layer0_outputs(3029));
    outputs(3784) <= not((layer0_outputs(6637)) xor (layer0_outputs(2817)));
    outputs(3785) <= not((layer0_outputs(622)) xor (layer0_outputs(1371)));
    outputs(3786) <= not((layer0_outputs(4035)) and (layer0_outputs(6200)));
    outputs(3787) <= (layer0_outputs(1944)) xor (layer0_outputs(6505));
    outputs(3788) <= (layer0_outputs(5382)) and not (layer0_outputs(7336));
    outputs(3789) <= not(layer0_outputs(5708));
    outputs(3790) <= not(layer0_outputs(2586));
    outputs(3791) <= (layer0_outputs(4928)) and not (layer0_outputs(4891));
    outputs(3792) <= (layer0_outputs(337)) and not (layer0_outputs(2693));
    outputs(3793) <= layer0_outputs(2625);
    outputs(3794) <= (layer0_outputs(5393)) and not (layer0_outputs(3956));
    outputs(3795) <= not(layer0_outputs(580));
    outputs(3796) <= not((layer0_outputs(2417)) xor (layer0_outputs(4415)));
    outputs(3797) <= layer0_outputs(1099);
    outputs(3798) <= not((layer0_outputs(7670)) xor (layer0_outputs(5089)));
    outputs(3799) <= layer0_outputs(808);
    outputs(3800) <= layer0_outputs(2283);
    outputs(3801) <= (layer0_outputs(2905)) and not (layer0_outputs(5258));
    outputs(3802) <= layer0_outputs(1073);
    outputs(3803) <= not(layer0_outputs(2090)) or (layer0_outputs(2805));
    outputs(3804) <= (layer0_outputs(2946)) xor (layer0_outputs(191));
    outputs(3805) <= not(layer0_outputs(628));
    outputs(3806) <= not((layer0_outputs(668)) or (layer0_outputs(3607)));
    outputs(3807) <= not(layer0_outputs(7607));
    outputs(3808) <= (layer0_outputs(5502)) and not (layer0_outputs(732));
    outputs(3809) <= layer0_outputs(2789);
    outputs(3810) <= (layer0_outputs(2781)) and not (layer0_outputs(6736));
    outputs(3811) <= not((layer0_outputs(301)) or (layer0_outputs(5955)));
    outputs(3812) <= not(layer0_outputs(2925)) or (layer0_outputs(6396));
    outputs(3813) <= not(layer0_outputs(5017));
    outputs(3814) <= layer0_outputs(1370);
    outputs(3815) <= layer0_outputs(1237);
    outputs(3816) <= (layer0_outputs(2748)) and not (layer0_outputs(4868));
    outputs(3817) <= (layer0_outputs(5079)) xor (layer0_outputs(4517));
    outputs(3818) <= (layer0_outputs(4275)) and (layer0_outputs(6761));
    outputs(3819) <= not((layer0_outputs(5650)) xor (layer0_outputs(4154)));
    outputs(3820) <= layer0_outputs(1079);
    outputs(3821) <= not(layer0_outputs(3284));
    outputs(3822) <= not(layer0_outputs(3988));
    outputs(3823) <= (layer0_outputs(2506)) or (layer0_outputs(5931));
    outputs(3824) <= not(layer0_outputs(1130));
    outputs(3825) <= (layer0_outputs(2397)) and not (layer0_outputs(908));
    outputs(3826) <= not(layer0_outputs(6842));
    outputs(3827) <= (layer0_outputs(124)) and (layer0_outputs(2192));
    outputs(3828) <= (layer0_outputs(2065)) xor (layer0_outputs(7529));
    outputs(3829) <= not((layer0_outputs(6203)) or (layer0_outputs(3036)));
    outputs(3830) <= not((layer0_outputs(5406)) or (layer0_outputs(6247)));
    outputs(3831) <= (layer0_outputs(4232)) and not (layer0_outputs(3803));
    outputs(3832) <= layer0_outputs(1200);
    outputs(3833) <= not(layer0_outputs(2423));
    outputs(3834) <= layer0_outputs(2321);
    outputs(3835) <= (layer0_outputs(3757)) and (layer0_outputs(7437));
    outputs(3836) <= (layer0_outputs(3761)) and not (layer0_outputs(348));
    outputs(3837) <= (layer0_outputs(4062)) xor (layer0_outputs(6489));
    outputs(3838) <= layer0_outputs(2484);
    outputs(3839) <= (layer0_outputs(3391)) xor (layer0_outputs(6057));
    outputs(3840) <= not(layer0_outputs(4145));
    outputs(3841) <= (layer0_outputs(4642)) and not (layer0_outputs(3536));
    outputs(3842) <= not((layer0_outputs(7393)) xor (layer0_outputs(6401)));
    outputs(3843) <= not((layer0_outputs(1868)) xor (layer0_outputs(930)));
    outputs(3844) <= not(layer0_outputs(3255)) or (layer0_outputs(6528));
    outputs(3845) <= not(layer0_outputs(1631)) or (layer0_outputs(4112));
    outputs(3846) <= not((layer0_outputs(7127)) xor (layer0_outputs(2822)));
    outputs(3847) <= (layer0_outputs(6829)) xor (layer0_outputs(5265));
    outputs(3848) <= not(layer0_outputs(4851)) or (layer0_outputs(2724));
    outputs(3849) <= not((layer0_outputs(4175)) or (layer0_outputs(6029)));
    outputs(3850) <= layer0_outputs(5962);
    outputs(3851) <= layer0_outputs(6404);
    outputs(3852) <= (layer0_outputs(5129)) and not (layer0_outputs(454));
    outputs(3853) <= not((layer0_outputs(6562)) xor (layer0_outputs(5652)));
    outputs(3854) <= (layer0_outputs(802)) xor (layer0_outputs(4399));
    outputs(3855) <= layer0_outputs(2273);
    outputs(3856) <= not(layer0_outputs(1728));
    outputs(3857) <= not(layer0_outputs(5655));
    outputs(3858) <= not(layer0_outputs(3483));
    outputs(3859) <= not(layer0_outputs(7156)) or (layer0_outputs(7379));
    outputs(3860) <= not((layer0_outputs(5164)) and (layer0_outputs(6178)));
    outputs(3861) <= not((layer0_outputs(4047)) xor (layer0_outputs(6533)));
    outputs(3862) <= (layer0_outputs(6615)) xor (layer0_outputs(6720));
    outputs(3863) <= (layer0_outputs(5830)) and (layer0_outputs(4558));
    outputs(3864) <= (layer0_outputs(3042)) and (layer0_outputs(3529));
    outputs(3865) <= (layer0_outputs(3307)) xor (layer0_outputs(6719));
    outputs(3866) <= layer0_outputs(4516);
    outputs(3867) <= not(layer0_outputs(343));
    outputs(3868) <= not(layer0_outputs(5914)) or (layer0_outputs(4152));
    outputs(3869) <= (layer0_outputs(122)) and (layer0_outputs(2217));
    outputs(3870) <= layer0_outputs(2313);
    outputs(3871) <= (layer0_outputs(3868)) or (layer0_outputs(4945));
    outputs(3872) <= not(layer0_outputs(3748));
    outputs(3873) <= not((layer0_outputs(6451)) and (layer0_outputs(5894)));
    outputs(3874) <= not(layer0_outputs(2382)) or (layer0_outputs(4822));
    outputs(3875) <= layer0_outputs(1271);
    outputs(3876) <= layer0_outputs(7580);
    outputs(3877) <= not((layer0_outputs(4515)) xor (layer0_outputs(6110)));
    outputs(3878) <= layer0_outputs(7457);
    outputs(3879) <= not((layer0_outputs(1688)) or (layer0_outputs(357)));
    outputs(3880) <= not(layer0_outputs(4785));
    outputs(3881) <= not(layer0_outputs(3208)) or (layer0_outputs(1872));
    outputs(3882) <= layer0_outputs(7435);
    outputs(3883) <= (layer0_outputs(5034)) xor (layer0_outputs(2812));
    outputs(3884) <= not(layer0_outputs(6773)) or (layer0_outputs(5278));
    outputs(3885) <= not(layer0_outputs(79));
    outputs(3886) <= not((layer0_outputs(3569)) xor (layer0_outputs(340)));
    outputs(3887) <= (layer0_outputs(1727)) or (layer0_outputs(3791));
    outputs(3888) <= not(layer0_outputs(6922)) or (layer0_outputs(4433));
    outputs(3889) <= (layer0_outputs(4786)) xor (layer0_outputs(3841));
    outputs(3890) <= (layer0_outputs(5904)) xor (layer0_outputs(2038));
    outputs(3891) <= not(layer0_outputs(5122)) or (layer0_outputs(2307));
    outputs(3892) <= layer0_outputs(5441);
    outputs(3893) <= (layer0_outputs(3887)) or (layer0_outputs(3211));
    outputs(3894) <= not(layer0_outputs(1806));
    outputs(3895) <= not((layer0_outputs(3344)) xor (layer0_outputs(6895)));
    outputs(3896) <= not((layer0_outputs(6779)) or (layer0_outputs(5522)));
    outputs(3897) <= (layer0_outputs(961)) and (layer0_outputs(6521));
    outputs(3898) <= not(layer0_outputs(2789)) or (layer0_outputs(5940));
    outputs(3899) <= layer0_outputs(7104);
    outputs(3900) <= not(layer0_outputs(4663));
    outputs(3901) <= (layer0_outputs(5590)) xor (layer0_outputs(6871));
    outputs(3902) <= (layer0_outputs(5046)) xor (layer0_outputs(1304));
    outputs(3903) <= not(layer0_outputs(1754));
    outputs(3904) <= layer0_outputs(1240);
    outputs(3905) <= not((layer0_outputs(1279)) xor (layer0_outputs(573)));
    outputs(3906) <= not((layer0_outputs(64)) xor (layer0_outputs(6848)));
    outputs(3907) <= not(layer0_outputs(7081));
    outputs(3908) <= not((layer0_outputs(6050)) or (layer0_outputs(3468)));
    outputs(3909) <= not((layer0_outputs(7125)) or (layer0_outputs(1285)));
    outputs(3910) <= layer0_outputs(6784);
    outputs(3911) <= (layer0_outputs(3295)) and not (layer0_outputs(5025));
    outputs(3912) <= not(layer0_outputs(6535)) or (layer0_outputs(2771));
    outputs(3913) <= not((layer0_outputs(6363)) xor (layer0_outputs(59)));
    outputs(3914) <= not(layer0_outputs(2361));
    outputs(3915) <= layer0_outputs(6498);
    outputs(3916) <= not(layer0_outputs(2230)) or (layer0_outputs(5333));
    outputs(3917) <= not(layer0_outputs(32));
    outputs(3918) <= layer0_outputs(1448);
    outputs(3919) <= not(layer0_outputs(7318));
    outputs(3920) <= not(layer0_outputs(1290));
    outputs(3921) <= not((layer0_outputs(3286)) xor (layer0_outputs(1694)));
    outputs(3922) <= layer0_outputs(2073);
    outputs(3923) <= (layer0_outputs(4744)) xor (layer0_outputs(6545));
    outputs(3924) <= (layer0_outputs(3796)) and (layer0_outputs(1543));
    outputs(3925) <= (layer0_outputs(1196)) and not (layer0_outputs(7422));
    outputs(3926) <= not(layer0_outputs(901));
    outputs(3927) <= not((layer0_outputs(457)) or (layer0_outputs(6542)));
    outputs(3928) <= layer0_outputs(2501);
    outputs(3929) <= (layer0_outputs(5976)) xor (layer0_outputs(4851));
    outputs(3930) <= (layer0_outputs(3348)) and not (layer0_outputs(5756));
    outputs(3931) <= not(layer0_outputs(6036));
    outputs(3932) <= not(layer0_outputs(1555)) or (layer0_outputs(1965));
    outputs(3933) <= (layer0_outputs(3409)) xor (layer0_outputs(5802));
    outputs(3934) <= not(layer0_outputs(6124));
    outputs(3935) <= not((layer0_outputs(1744)) or (layer0_outputs(7405)));
    outputs(3936) <= layer0_outputs(5107);
    outputs(3937) <= not(layer0_outputs(7201)) or (layer0_outputs(3833));
    outputs(3938) <= (layer0_outputs(4990)) and not (layer0_outputs(5643));
    outputs(3939) <= layer0_outputs(5103);
    outputs(3940) <= (layer0_outputs(2565)) and not (layer0_outputs(134));
    outputs(3941) <= layer0_outputs(1027);
    outputs(3942) <= layer0_outputs(5233);
    outputs(3943) <= not(layer0_outputs(7213)) or (layer0_outputs(4647));
    outputs(3944) <= not((layer0_outputs(4810)) or (layer0_outputs(2810)));
    outputs(3945) <= not(layer0_outputs(3726));
    outputs(3946) <= not((layer0_outputs(40)) xor (layer0_outputs(5126)));
    outputs(3947) <= not(layer0_outputs(4574));
    outputs(3948) <= layer0_outputs(7162);
    outputs(3949) <= (layer0_outputs(1076)) xor (layer0_outputs(1445));
    outputs(3950) <= layer0_outputs(5395);
    outputs(3951) <= not((layer0_outputs(2218)) xor (layer0_outputs(5389)));
    outputs(3952) <= not(layer0_outputs(4213));
    outputs(3953) <= layer0_outputs(984);
    outputs(3954) <= (layer0_outputs(6935)) xor (layer0_outputs(4233));
    outputs(3955) <= not(layer0_outputs(3231));
    outputs(3956) <= not((layer0_outputs(3514)) xor (layer0_outputs(2438)));
    outputs(3957) <= layer0_outputs(3040);
    outputs(3958) <= (layer0_outputs(5340)) xor (layer0_outputs(451));
    outputs(3959) <= not(layer0_outputs(4980));
    outputs(3960) <= layer0_outputs(6758);
    outputs(3961) <= '0';
    outputs(3962) <= not((layer0_outputs(6687)) xor (layer0_outputs(6601)));
    outputs(3963) <= not(layer0_outputs(891));
    outputs(3964) <= layer0_outputs(7246);
    outputs(3965) <= layer0_outputs(6003);
    outputs(3966) <= not(layer0_outputs(5726));
    outputs(3967) <= not((layer0_outputs(2617)) xor (layer0_outputs(77)));
    outputs(3968) <= (layer0_outputs(2889)) xor (layer0_outputs(6444));
    outputs(3969) <= not((layer0_outputs(4176)) and (layer0_outputs(1921)));
    outputs(3970) <= layer0_outputs(6706);
    outputs(3971) <= not(layer0_outputs(7228));
    outputs(3972) <= (layer0_outputs(2842)) or (layer0_outputs(4147));
    outputs(3973) <= not((layer0_outputs(5363)) xor (layer0_outputs(4033)));
    outputs(3974) <= not((layer0_outputs(5313)) or (layer0_outputs(3408)));
    outputs(3975) <= not(layer0_outputs(7571));
    outputs(3976) <= not(layer0_outputs(5696)) or (layer0_outputs(5038));
    outputs(3977) <= (layer0_outputs(7622)) and not (layer0_outputs(1168));
    outputs(3978) <= not(layer0_outputs(1215));
    outputs(3979) <= (layer0_outputs(3333)) and (layer0_outputs(6525));
    outputs(3980) <= not((layer0_outputs(6666)) xor (layer0_outputs(470)));
    outputs(3981) <= layer0_outputs(3596);
    outputs(3982) <= not((layer0_outputs(6392)) xor (layer0_outputs(6243)));
    outputs(3983) <= layer0_outputs(5249);
    outputs(3984) <= not(layer0_outputs(2758));
    outputs(3985) <= (layer0_outputs(6002)) and not (layer0_outputs(3492));
    outputs(3986) <= not(layer0_outputs(3602));
    outputs(3987) <= not(layer0_outputs(4514));
    outputs(3988) <= not(layer0_outputs(2319)) or (layer0_outputs(6696));
    outputs(3989) <= layer0_outputs(6581);
    outputs(3990) <= not(layer0_outputs(1655));
    outputs(3991) <= layer0_outputs(1656);
    outputs(3992) <= (layer0_outputs(1317)) xor (layer0_outputs(5430));
    outputs(3993) <= not((layer0_outputs(6146)) or (layer0_outputs(4779)));
    outputs(3994) <= layer0_outputs(4369);
    outputs(3995) <= not(layer0_outputs(3660));
    outputs(3996) <= not(layer0_outputs(7068));
    outputs(3997) <= layer0_outputs(2125);
    outputs(3998) <= not(layer0_outputs(2148));
    outputs(3999) <= layer0_outputs(5608);
    outputs(4000) <= (layer0_outputs(6540)) or (layer0_outputs(6304));
    outputs(4001) <= (layer0_outputs(6261)) xor (layer0_outputs(7060));
    outputs(4002) <= layer0_outputs(3393);
    outputs(4003) <= layer0_outputs(6484);
    outputs(4004) <= not(layer0_outputs(3810));
    outputs(4005) <= not(layer0_outputs(4240));
    outputs(4006) <= (layer0_outputs(3215)) and not (layer0_outputs(5913));
    outputs(4007) <= not(layer0_outputs(1869)) or (layer0_outputs(6590));
    outputs(4008) <= not((layer0_outputs(4332)) or (layer0_outputs(6448)));
    outputs(4009) <= not(layer0_outputs(3015)) or (layer0_outputs(2248));
    outputs(4010) <= layer0_outputs(6946);
    outputs(4011) <= (layer0_outputs(498)) or (layer0_outputs(410));
    outputs(4012) <= (layer0_outputs(5548)) or (layer0_outputs(7545));
    outputs(4013) <= not(layer0_outputs(1554));
    outputs(4014) <= (layer0_outputs(2320)) xor (layer0_outputs(6713));
    outputs(4015) <= layer0_outputs(4802);
    outputs(4016) <= layer0_outputs(1374);
    outputs(4017) <= (layer0_outputs(1949)) xor (layer0_outputs(1269));
    outputs(4018) <= layer0_outputs(3251);
    outputs(4019) <= (layer0_outputs(4557)) and (layer0_outputs(2009));
    outputs(4020) <= not((layer0_outputs(4742)) or (layer0_outputs(4118)));
    outputs(4021) <= (layer0_outputs(7321)) and (layer0_outputs(4487));
    outputs(4022) <= (layer0_outputs(6546)) or (layer0_outputs(3359));
    outputs(4023) <= not(layer0_outputs(6437)) or (layer0_outputs(5535));
    outputs(4024) <= not((layer0_outputs(3924)) or (layer0_outputs(3930)));
    outputs(4025) <= not(layer0_outputs(7397));
    outputs(4026) <= (layer0_outputs(2220)) or (layer0_outputs(6940));
    outputs(4027) <= layer0_outputs(3150);
    outputs(4028) <= not(layer0_outputs(6730)) or (layer0_outputs(5508));
    outputs(4029) <= (layer0_outputs(3102)) and not (layer0_outputs(491));
    outputs(4030) <= layer0_outputs(3066);
    outputs(4031) <= not((layer0_outputs(1930)) xor (layer0_outputs(7146)));
    outputs(4032) <= (layer0_outputs(6785)) and not (layer0_outputs(2132));
    outputs(4033) <= (layer0_outputs(4024)) xor (layer0_outputs(3996));
    outputs(4034) <= (layer0_outputs(4051)) xor (layer0_outputs(5708));
    outputs(4035) <= (layer0_outputs(569)) or (layer0_outputs(2073));
    outputs(4036) <= not((layer0_outputs(5695)) and (layer0_outputs(845)));
    outputs(4037) <= (layer0_outputs(7202)) and not (layer0_outputs(3698));
    outputs(4038) <= (layer0_outputs(1366)) and (layer0_outputs(2804));
    outputs(4039) <= not((layer0_outputs(1090)) or (layer0_outputs(7226)));
    outputs(4040) <= (layer0_outputs(5485)) and not (layer0_outputs(2281));
    outputs(4041) <= layer0_outputs(87);
    outputs(4042) <= (layer0_outputs(4388)) xor (layer0_outputs(917));
    outputs(4043) <= (layer0_outputs(4106)) xor (layer0_outputs(5665));
    outputs(4044) <= not(layer0_outputs(607));
    outputs(4045) <= (layer0_outputs(1414)) and not (layer0_outputs(97));
    outputs(4046) <= not(layer0_outputs(5950));
    outputs(4047) <= layer0_outputs(6603);
    outputs(4048) <= not((layer0_outputs(6611)) and (layer0_outputs(6986)));
    outputs(4049) <= not((layer0_outputs(3243)) xor (layer0_outputs(2189)));
    outputs(4050) <= not((layer0_outputs(7297)) and (layer0_outputs(706)));
    outputs(4051) <= layer0_outputs(2887);
    outputs(4052) <= not(layer0_outputs(2379)) or (layer0_outputs(24));
    outputs(4053) <= not(layer0_outputs(2695));
    outputs(4054) <= (layer0_outputs(685)) xor (layer0_outputs(2194));
    outputs(4055) <= layer0_outputs(5232);
    outputs(4056) <= not(layer0_outputs(2775));
    outputs(4057) <= not(layer0_outputs(2928));
    outputs(4058) <= (layer0_outputs(6325)) or (layer0_outputs(1870));
    outputs(4059) <= not((layer0_outputs(5044)) and (layer0_outputs(3810)));
    outputs(4060) <= layer0_outputs(3087);
    outputs(4061) <= (layer0_outputs(5387)) and not (layer0_outputs(5327));
    outputs(4062) <= (layer0_outputs(5518)) xor (layer0_outputs(5126));
    outputs(4063) <= (layer0_outputs(644)) xor (layer0_outputs(6068));
    outputs(4064) <= not(layer0_outputs(7043));
    outputs(4065) <= not(layer0_outputs(3847)) or (layer0_outputs(3285));
    outputs(4066) <= not(layer0_outputs(6854));
    outputs(4067) <= layer0_outputs(5733);
    outputs(4068) <= not((layer0_outputs(7665)) xor (layer0_outputs(4512)));
    outputs(4069) <= not(layer0_outputs(6229));
    outputs(4070) <= (layer0_outputs(224)) xor (layer0_outputs(1178));
    outputs(4071) <= not(layer0_outputs(5242));
    outputs(4072) <= not(layer0_outputs(963));
    outputs(4073) <= layer0_outputs(6239);
    outputs(4074) <= not(layer0_outputs(586));
    outputs(4075) <= (layer0_outputs(931)) or (layer0_outputs(5534));
    outputs(4076) <= not(layer0_outputs(6185));
    outputs(4077) <= layer0_outputs(5087);
    outputs(4078) <= not((layer0_outputs(5411)) and (layer0_outputs(43)));
    outputs(4079) <= not((layer0_outputs(2465)) xor (layer0_outputs(2623)));
    outputs(4080) <= not(layer0_outputs(5175)) or (layer0_outputs(7597));
    outputs(4081) <= not(layer0_outputs(5964));
    outputs(4082) <= (layer0_outputs(2848)) and (layer0_outputs(5953));
    outputs(4083) <= not((layer0_outputs(6098)) xor (layer0_outputs(276)));
    outputs(4084) <= not(layer0_outputs(5347));
    outputs(4085) <= not((layer0_outputs(4491)) xor (layer0_outputs(7388)));
    outputs(4086) <= not(layer0_outputs(4919));
    outputs(4087) <= layer0_outputs(7520);
    outputs(4088) <= not((layer0_outputs(4345)) or (layer0_outputs(7620)));
    outputs(4089) <= not((layer0_outputs(3889)) xor (layer0_outputs(1236)));
    outputs(4090) <= not((layer0_outputs(1556)) xor (layer0_outputs(1284)));
    outputs(4091) <= (layer0_outputs(3019)) xor (layer0_outputs(3075));
    outputs(4092) <= not(layer0_outputs(243));
    outputs(4093) <= not((layer0_outputs(2426)) xor (layer0_outputs(6130)));
    outputs(4094) <= (layer0_outputs(2421)) xor (layer0_outputs(3717));
    outputs(4095) <= not((layer0_outputs(7230)) xor (layer0_outputs(2548)));
    outputs(4096) <= not(layer0_outputs(6108));
    outputs(4097) <= layer0_outputs(6674);
    outputs(4098) <= layer0_outputs(2154);
    outputs(4099) <= layer0_outputs(214);
    outputs(4100) <= not(layer0_outputs(5063));
    outputs(4101) <= (layer0_outputs(6140)) xor (layer0_outputs(4232));
    outputs(4102) <= not(layer0_outputs(5163));
    outputs(4103) <= not((layer0_outputs(2226)) and (layer0_outputs(7492)));
    outputs(4104) <= not(layer0_outputs(2708));
    outputs(4105) <= layer0_outputs(1251);
    outputs(4106) <= not(layer0_outputs(7090));
    outputs(4107) <= layer0_outputs(2536);
    outputs(4108) <= not((layer0_outputs(6803)) and (layer0_outputs(2515)));
    outputs(4109) <= not(layer0_outputs(3259));
    outputs(4110) <= (layer0_outputs(520)) xor (layer0_outputs(7036));
    outputs(4111) <= (layer0_outputs(266)) xor (layer0_outputs(6960));
    outputs(4112) <= layer0_outputs(7668);
    outputs(4113) <= not((layer0_outputs(1768)) and (layer0_outputs(7302)));
    outputs(4114) <= not(layer0_outputs(6607));
    outputs(4115) <= not(layer0_outputs(3294));
    outputs(4116) <= (layer0_outputs(1163)) and not (layer0_outputs(6221));
    outputs(4117) <= not(layer0_outputs(3693)) or (layer0_outputs(6004));
    outputs(4118) <= not(layer0_outputs(3508)) or (layer0_outputs(4352));
    outputs(4119) <= (layer0_outputs(5604)) and not (layer0_outputs(2017));
    outputs(4120) <= layer0_outputs(270);
    outputs(4121) <= layer0_outputs(3576);
    outputs(4122) <= not((layer0_outputs(6196)) xor (layer0_outputs(6473)));
    outputs(4123) <= layer0_outputs(2247);
    outputs(4124) <= not(layer0_outputs(5365));
    outputs(4125) <= not(layer0_outputs(7205));
    outputs(4126) <= layer0_outputs(6916);
    outputs(4127) <= layer0_outputs(1004);
    outputs(4128) <= not(layer0_outputs(727));
    outputs(4129) <= not(layer0_outputs(6227)) or (layer0_outputs(2557));
    outputs(4130) <= layer0_outputs(7414);
    outputs(4131) <= not((layer0_outputs(430)) xor (layer0_outputs(2941)));
    outputs(4132) <= (layer0_outputs(2423)) and not (layer0_outputs(6270));
    outputs(4133) <= not((layer0_outputs(1732)) xor (layer0_outputs(500)));
    outputs(4134) <= not((layer0_outputs(6385)) or (layer0_outputs(167)));
    outputs(4135) <= not(layer0_outputs(3367));
    outputs(4136) <= not((layer0_outputs(6012)) and (layer0_outputs(174)));
    outputs(4137) <= (layer0_outputs(6228)) xor (layer0_outputs(1795));
    outputs(4138) <= layer0_outputs(3892);
    outputs(4139) <= not((layer0_outputs(7286)) or (layer0_outputs(5799)));
    outputs(4140) <= (layer0_outputs(953)) and not (layer0_outputs(6599));
    outputs(4141) <= (layer0_outputs(7060)) xor (layer0_outputs(6917));
    outputs(4142) <= (layer0_outputs(653)) xor (layer0_outputs(2059));
    outputs(4143) <= (layer0_outputs(6150)) xor (layer0_outputs(4295));
    outputs(4144) <= not(layer0_outputs(4846));
    outputs(4145) <= not(layer0_outputs(4253));
    outputs(4146) <= not((layer0_outputs(2552)) or (layer0_outputs(6817)));
    outputs(4147) <= not((layer0_outputs(3498)) xor (layer0_outputs(5203)));
    outputs(4148) <= (layer0_outputs(3422)) xor (layer0_outputs(4617));
    outputs(4149) <= layer0_outputs(4909);
    outputs(4150) <= not((layer0_outputs(4835)) xor (layer0_outputs(4348)));
    outputs(4151) <= not((layer0_outputs(3909)) xor (layer0_outputs(6385)));
    outputs(4152) <= not((layer0_outputs(1365)) xor (layer0_outputs(3537)));
    outputs(4153) <= (layer0_outputs(2790)) xor (layer0_outputs(1405));
    outputs(4154) <= not(layer0_outputs(3857));
    outputs(4155) <= not(layer0_outputs(6748));
    outputs(4156) <= (layer0_outputs(2683)) xor (layer0_outputs(3019));
    outputs(4157) <= not(layer0_outputs(724));
    outputs(4158) <= layer0_outputs(5647);
    outputs(4159) <= (layer0_outputs(7369)) and not (layer0_outputs(4747));
    outputs(4160) <= layer0_outputs(5108);
    outputs(4161) <= not((layer0_outputs(1107)) xor (layer0_outputs(7606)));
    outputs(4162) <= not(layer0_outputs(5054));
    outputs(4163) <= not(layer0_outputs(5128));
    outputs(4164) <= (layer0_outputs(2651)) xor (layer0_outputs(1247));
    outputs(4165) <= not((layer0_outputs(3668)) or (layer0_outputs(3289)));
    outputs(4166) <= (layer0_outputs(7037)) or (layer0_outputs(1738));
    outputs(4167) <= not(layer0_outputs(1428)) or (layer0_outputs(1762));
    outputs(4168) <= (layer0_outputs(1846)) xor (layer0_outputs(4553));
    outputs(4169) <= not((layer0_outputs(4570)) xor (layer0_outputs(819)));
    outputs(4170) <= not((layer0_outputs(34)) xor (layer0_outputs(4307)));
    outputs(4171) <= not(layer0_outputs(4884)) or (layer0_outputs(1788));
    outputs(4172) <= layer0_outputs(4294);
    outputs(4173) <= not(layer0_outputs(1973));
    outputs(4174) <= not(layer0_outputs(1075)) or (layer0_outputs(6959));
    outputs(4175) <= not(layer0_outputs(6975));
    outputs(4176) <= layer0_outputs(2220);
    outputs(4177) <= layer0_outputs(1807);
    outputs(4178) <= not((layer0_outputs(5783)) xor (layer0_outputs(2295)));
    outputs(4179) <= layer0_outputs(7057);
    outputs(4180) <= (layer0_outputs(3280)) xor (layer0_outputs(6487));
    outputs(4181) <= (layer0_outputs(5574)) xor (layer0_outputs(3672));
    outputs(4182) <= layer0_outputs(2464);
    outputs(4183) <= not(layer0_outputs(3256));
    outputs(4184) <= layer0_outputs(4117);
    outputs(4185) <= not(layer0_outputs(7023));
    outputs(4186) <= (layer0_outputs(6904)) xor (layer0_outputs(892));
    outputs(4187) <= not((layer0_outputs(3436)) xor (layer0_outputs(710)));
    outputs(4188) <= not((layer0_outputs(4854)) or (layer0_outputs(2011)));
    outputs(4189) <= layer0_outputs(7502);
    outputs(4190) <= layer0_outputs(3726);
    outputs(4191) <= (layer0_outputs(5059)) xor (layer0_outputs(902));
    outputs(4192) <= (layer0_outputs(967)) xor (layer0_outputs(6899));
    outputs(4193) <= not(layer0_outputs(4381));
    outputs(4194) <= (layer0_outputs(2909)) and not (layer0_outputs(3767));
    outputs(4195) <= not((layer0_outputs(4104)) xor (layer0_outputs(3080)));
    outputs(4196) <= not((layer0_outputs(1418)) xor (layer0_outputs(5207)));
    outputs(4197) <= not((layer0_outputs(6471)) xor (layer0_outputs(1133)));
    outputs(4198) <= (layer0_outputs(4006)) and not (layer0_outputs(4964));
    outputs(4199) <= not(layer0_outputs(7333));
    outputs(4200) <= not((layer0_outputs(6605)) xor (layer0_outputs(4721)));
    outputs(4201) <= not((layer0_outputs(7170)) or (layer0_outputs(1408)));
    outputs(4202) <= layer0_outputs(3417);
    outputs(4203) <= layer0_outputs(6860);
    outputs(4204) <= not((layer0_outputs(2802)) or (layer0_outputs(7189)));
    outputs(4205) <= (layer0_outputs(4041)) or (layer0_outputs(3485));
    outputs(4206) <= not((layer0_outputs(4509)) or (layer0_outputs(2110)));
    outputs(4207) <= not(layer0_outputs(6208));
    outputs(4208) <= (layer0_outputs(38)) xor (layer0_outputs(4406));
    outputs(4209) <= (layer0_outputs(1865)) xor (layer0_outputs(537));
    outputs(4210) <= not(layer0_outputs(3388));
    outputs(4211) <= not(layer0_outputs(7105)) or (layer0_outputs(2838));
    outputs(4212) <= not(layer0_outputs(360));
    outputs(4213) <= not(layer0_outputs(1695));
    outputs(4214) <= (layer0_outputs(1628)) xor (layer0_outputs(7103));
    outputs(4215) <= (layer0_outputs(2642)) xor (layer0_outputs(3307));
    outputs(4216) <= (layer0_outputs(3101)) and not (layer0_outputs(5134));
    outputs(4217) <= not(layer0_outputs(2152));
    outputs(4218) <= not((layer0_outputs(5686)) and (layer0_outputs(6170)));
    outputs(4219) <= not(layer0_outputs(3411));
    outputs(4220) <= not(layer0_outputs(6183));
    outputs(4221) <= not(layer0_outputs(6894)) or (layer0_outputs(7401));
    outputs(4222) <= not(layer0_outputs(4717));
    outputs(4223) <= not(layer0_outputs(5960)) or (layer0_outputs(459));
    outputs(4224) <= (layer0_outputs(7059)) and not (layer0_outputs(6128));
    outputs(4225) <= (layer0_outputs(1561)) xor (layer0_outputs(542));
    outputs(4226) <= (layer0_outputs(297)) and not (layer0_outputs(6425));
    outputs(4227) <= not((layer0_outputs(4332)) and (layer0_outputs(5751)));
    outputs(4228) <= not((layer0_outputs(2885)) xor (layer0_outputs(4284)));
    outputs(4229) <= not((layer0_outputs(2847)) xor (layer0_outputs(6672)));
    outputs(4230) <= (layer0_outputs(4004)) or (layer0_outputs(4848));
    outputs(4231) <= not(layer0_outputs(216));
    outputs(4232) <= not(layer0_outputs(7205));
    outputs(4233) <= (layer0_outputs(6245)) and not (layer0_outputs(5524));
    outputs(4234) <= (layer0_outputs(4741)) xor (layer0_outputs(2687));
    outputs(4235) <= not(layer0_outputs(5695)) or (layer0_outputs(2422));
    outputs(4236) <= (layer0_outputs(538)) and not (layer0_outputs(6266));
    outputs(4237) <= (layer0_outputs(1058)) and not (layer0_outputs(2611));
    outputs(4238) <= not(layer0_outputs(286));
    outputs(4239) <= (layer0_outputs(3419)) and not (layer0_outputs(7155));
    outputs(4240) <= not(layer0_outputs(2685));
    outputs(4241) <= not(layer0_outputs(6067)) or (layer0_outputs(2919));
    outputs(4242) <= not((layer0_outputs(2040)) xor (layer0_outputs(1304)));
    outputs(4243) <= not(layer0_outputs(4994)) or (layer0_outputs(5911));
    outputs(4244) <= not((layer0_outputs(3340)) or (layer0_outputs(6807)));
    outputs(4245) <= not(layer0_outputs(5823));
    outputs(4246) <= layer0_outputs(3003);
    outputs(4247) <= (layer0_outputs(1343)) and not (layer0_outputs(7250));
    outputs(4248) <= (layer0_outputs(6218)) xor (layer0_outputs(2001));
    outputs(4249) <= not((layer0_outputs(687)) and (layer0_outputs(1138)));
    outputs(4250) <= (layer0_outputs(5438)) xor (layer0_outputs(1713));
    outputs(4251) <= (layer0_outputs(5326)) or (layer0_outputs(4041));
    outputs(4252) <= not(layer0_outputs(5679));
    outputs(4253) <= not((layer0_outputs(3567)) and (layer0_outputs(6924)));
    outputs(4254) <= not((layer0_outputs(5379)) xor (layer0_outputs(1722)));
    outputs(4255) <= layer0_outputs(4136);
    outputs(4256) <= (layer0_outputs(730)) xor (layer0_outputs(6047));
    outputs(4257) <= not(layer0_outputs(6317));
    outputs(4258) <= not((layer0_outputs(196)) xor (layer0_outputs(1724)));
    outputs(4259) <= not((layer0_outputs(4405)) and (layer0_outputs(4263)));
    outputs(4260) <= not((layer0_outputs(5240)) xor (layer0_outputs(3184)));
    outputs(4261) <= layer0_outputs(2164);
    outputs(4262) <= (layer0_outputs(5252)) xor (layer0_outputs(5952));
    outputs(4263) <= not((layer0_outputs(6283)) xor (layer0_outputs(7627)));
    outputs(4264) <= not(layer0_outputs(320));
    outputs(4265) <= not((layer0_outputs(3802)) xor (layer0_outputs(1566)));
    outputs(4266) <= not((layer0_outputs(1613)) and (layer0_outputs(43)));
    outputs(4267) <= not(layer0_outputs(2885));
    outputs(4268) <= (layer0_outputs(3344)) xor (layer0_outputs(7358));
    outputs(4269) <= layer0_outputs(7616);
    outputs(4270) <= (layer0_outputs(4037)) xor (layer0_outputs(7331));
    outputs(4271) <= (layer0_outputs(933)) and not (layer0_outputs(4710));
    outputs(4272) <= not((layer0_outputs(6067)) xor (layer0_outputs(366)));
    outputs(4273) <= (layer0_outputs(5648)) xor (layer0_outputs(567));
    outputs(4274) <= not((layer0_outputs(2830)) xor (layer0_outputs(1613)));
    outputs(4275) <= not(layer0_outputs(6249));
    outputs(4276) <= layer0_outputs(1454);
    outputs(4277) <= layer0_outputs(6144);
    outputs(4278) <= not(layer0_outputs(3515)) or (layer0_outputs(2621));
    outputs(4279) <= not(layer0_outputs(1557));
    outputs(4280) <= not(layer0_outputs(6211));
    outputs(4281) <= not(layer0_outputs(6648));
    outputs(4282) <= layer0_outputs(5021);
    outputs(4283) <= layer0_outputs(6426);
    outputs(4284) <= not(layer0_outputs(4372));
    outputs(4285) <= layer0_outputs(716);
    outputs(4286) <= (layer0_outputs(919)) xor (layer0_outputs(5497));
    outputs(4287) <= not(layer0_outputs(3100));
    outputs(4288) <= not(layer0_outputs(7509)) or (layer0_outputs(6113));
    outputs(4289) <= not(layer0_outputs(85));
    outputs(4290) <= not(layer0_outputs(5473));
    outputs(4291) <= layer0_outputs(2352);
    outputs(4292) <= not((layer0_outputs(4410)) xor (layer0_outputs(7382)));
    outputs(4293) <= layer0_outputs(5660);
    outputs(4294) <= not((layer0_outputs(3737)) xor (layer0_outputs(2487)));
    outputs(4295) <= (layer0_outputs(2903)) xor (layer0_outputs(4050));
    outputs(4296) <= (layer0_outputs(180)) or (layer0_outputs(5263));
    outputs(4297) <= not(layer0_outputs(3140));
    outputs(4298) <= layer0_outputs(2197);
    outputs(4299) <= not((layer0_outputs(6805)) xor (layer0_outputs(5278)));
    outputs(4300) <= layer0_outputs(2651);
    outputs(4301) <= layer0_outputs(7163);
    outputs(4302) <= (layer0_outputs(2539)) xor (layer0_outputs(3109));
    outputs(4303) <= not((layer0_outputs(4264)) or (layer0_outputs(4732)));
    outputs(4304) <= layer0_outputs(5868);
    outputs(4305) <= (layer0_outputs(5027)) or (layer0_outputs(3822));
    outputs(4306) <= not(layer0_outputs(5737)) or (layer0_outputs(561));
    outputs(4307) <= layer0_outputs(3226);
    outputs(4308) <= not((layer0_outputs(2319)) and (layer0_outputs(3358)));
    outputs(4309) <= (layer0_outputs(538)) and (layer0_outputs(5064));
    outputs(4310) <= layer0_outputs(4411);
    outputs(4311) <= not(layer0_outputs(4918));
    outputs(4312) <= layer0_outputs(579);
    outputs(4313) <= (layer0_outputs(2452)) xor (layer0_outputs(2933));
    outputs(4314) <= not((layer0_outputs(4242)) or (layer0_outputs(4279)));
    outputs(4315) <= (layer0_outputs(6637)) xor (layer0_outputs(1804));
    outputs(4316) <= (layer0_outputs(2513)) and (layer0_outputs(6393));
    outputs(4317) <= (layer0_outputs(725)) or (layer0_outputs(5638));
    outputs(4318) <= not(layer0_outputs(757)) or (layer0_outputs(2100));
    outputs(4319) <= not(layer0_outputs(1505));
    outputs(4320) <= (layer0_outputs(5565)) and not (layer0_outputs(1471));
    outputs(4321) <= layer0_outputs(1062);
    outputs(4322) <= not(layer0_outputs(811)) or (layer0_outputs(2754));
    outputs(4323) <= not((layer0_outputs(6232)) or (layer0_outputs(6376)));
    outputs(4324) <= not((layer0_outputs(6738)) and (layer0_outputs(7251)));
    outputs(4325) <= layer0_outputs(1955);
    outputs(4326) <= not(layer0_outputs(1467));
    outputs(4327) <= not(layer0_outputs(6541));
    outputs(4328) <= not(layer0_outputs(6516));
    outputs(4329) <= not(layer0_outputs(1046)) or (layer0_outputs(2403));
    outputs(4330) <= not(layer0_outputs(2563));
    outputs(4331) <= (layer0_outputs(5187)) xor (layer0_outputs(88));
    outputs(4332) <= not(layer0_outputs(1258));
    outputs(4333) <= (layer0_outputs(2947)) xor (layer0_outputs(2840));
    outputs(4334) <= not((layer0_outputs(210)) xor (layer0_outputs(5421)));
    outputs(4335) <= layer0_outputs(4224);
    outputs(4336) <= layer0_outputs(4247);
    outputs(4337) <= (layer0_outputs(5530)) xor (layer0_outputs(2865));
    outputs(4338) <= (layer0_outputs(3907)) xor (layer0_outputs(7604));
    outputs(4339) <= layer0_outputs(1889);
    outputs(4340) <= layer0_outputs(2036);
    outputs(4341) <= (layer0_outputs(2375)) and (layer0_outputs(406));
    outputs(4342) <= not(layer0_outputs(6756));
    outputs(4343) <= not((layer0_outputs(3665)) xor (layer0_outputs(6420)));
    outputs(4344) <= not(layer0_outputs(6625));
    outputs(4345) <= not((layer0_outputs(4013)) or (layer0_outputs(202)));
    outputs(4346) <= not(layer0_outputs(6030));
    outputs(4347) <= not((layer0_outputs(1441)) xor (layer0_outputs(3750)));
    outputs(4348) <= (layer0_outputs(2638)) and (layer0_outputs(3742));
    outputs(4349) <= layer0_outputs(6738);
    outputs(4350) <= (layer0_outputs(2445)) and not (layer0_outputs(65));
    outputs(4351) <= '1';
    outputs(4352) <= (layer0_outputs(5111)) and not (layer0_outputs(4335));
    outputs(4353) <= (layer0_outputs(7086)) and not (layer0_outputs(4175));
    outputs(4354) <= (layer0_outputs(6697)) or (layer0_outputs(6452));
    outputs(4355) <= not(layer0_outputs(6570)) or (layer0_outputs(1193));
    outputs(4356) <= (layer0_outputs(3574)) and not (layer0_outputs(571));
    outputs(4357) <= (layer0_outputs(6675)) and (layer0_outputs(4797));
    outputs(4358) <= (layer0_outputs(798)) xor (layer0_outputs(7030));
    outputs(4359) <= not(layer0_outputs(3664));
    outputs(4360) <= not(layer0_outputs(6973)) or (layer0_outputs(2360));
    outputs(4361) <= (layer0_outputs(4556)) xor (layer0_outputs(5248));
    outputs(4362) <= not(layer0_outputs(6840));
    outputs(4363) <= '1';
    outputs(4364) <= layer0_outputs(626);
    outputs(4365) <= (layer0_outputs(7282)) and (layer0_outputs(6118));
    outputs(4366) <= (layer0_outputs(4665)) or (layer0_outputs(452));
    outputs(4367) <= layer0_outputs(5484);
    outputs(4368) <= '1';
    outputs(4369) <= layer0_outputs(3620);
    outputs(4370) <= (layer0_outputs(2622)) or (layer0_outputs(4452));
    outputs(4371) <= layer0_outputs(5899);
    outputs(4372) <= not(layer0_outputs(6566));
    outputs(4373) <= (layer0_outputs(4066)) xor (layer0_outputs(5450));
    outputs(4374) <= not((layer0_outputs(4293)) or (layer0_outputs(5749)));
    outputs(4375) <= not((layer0_outputs(2034)) xor (layer0_outputs(1065)));
    outputs(4376) <= not(layer0_outputs(7368)) or (layer0_outputs(3391));
    outputs(4377) <= layer0_outputs(4803);
    outputs(4378) <= not((layer0_outputs(5769)) and (layer0_outputs(294)));
    outputs(4379) <= layer0_outputs(1272);
    outputs(4380) <= (layer0_outputs(7550)) xor (layer0_outputs(6887));
    outputs(4381) <= not(layer0_outputs(910)) or (layer0_outputs(3341));
    outputs(4382) <= (layer0_outputs(1775)) xor (layer0_outputs(3365));
    outputs(4383) <= (layer0_outputs(2018)) and not (layer0_outputs(3851));
    outputs(4384) <= not(layer0_outputs(6311));
    outputs(4385) <= not((layer0_outputs(4721)) xor (layer0_outputs(6182)));
    outputs(4386) <= not(layer0_outputs(6929)) or (layer0_outputs(7545));
    outputs(4387) <= not((layer0_outputs(381)) xor (layer0_outputs(1715)));
    outputs(4388) <= not((layer0_outputs(4673)) and (layer0_outputs(9)));
    outputs(4389) <= not(layer0_outputs(5052));
    outputs(4390) <= not(layer0_outputs(1423));
    outputs(4391) <= not(layer0_outputs(1648));
    outputs(4392) <= (layer0_outputs(5802)) and (layer0_outputs(4708));
    outputs(4393) <= not((layer0_outputs(73)) xor (layer0_outputs(6168)));
    outputs(4394) <= (layer0_outputs(6147)) xor (layer0_outputs(6792));
    outputs(4395) <= not(layer0_outputs(758));
    outputs(4396) <= not(layer0_outputs(3680));
    outputs(4397) <= (layer0_outputs(836)) or (layer0_outputs(5135));
    outputs(4398) <= (layer0_outputs(7547)) and not (layer0_outputs(4603));
    outputs(4399) <= layer0_outputs(5868);
    outputs(4400) <= not(layer0_outputs(3100));
    outputs(4401) <= (layer0_outputs(334)) and not (layer0_outputs(5379));
    outputs(4402) <= layer0_outputs(7212);
    outputs(4403) <= not(layer0_outputs(3720));
    outputs(4404) <= not((layer0_outputs(4167)) or (layer0_outputs(5512)));
    outputs(4405) <= not((layer0_outputs(5566)) xor (layer0_outputs(6087)));
    outputs(4406) <= layer0_outputs(6147);
    outputs(4407) <= not((layer0_outputs(6759)) xor (layer0_outputs(634)));
    outputs(4408) <= layer0_outputs(4870);
    outputs(4409) <= not(layer0_outputs(1186));
    outputs(4410) <= (layer0_outputs(5760)) and not (layer0_outputs(4755));
    outputs(4411) <= not((layer0_outputs(5535)) xor (layer0_outputs(6022)));
    outputs(4412) <= (layer0_outputs(2125)) and not (layer0_outputs(1861));
    outputs(4413) <= layer0_outputs(957);
    outputs(4414) <= not(layer0_outputs(5855));
    outputs(4415) <= (layer0_outputs(7430)) xor (layer0_outputs(164));
    outputs(4416) <= (layer0_outputs(3794)) xor (layer0_outputs(7349));
    outputs(4417) <= not(layer0_outputs(1020));
    outputs(4418) <= (layer0_outputs(1886)) xor (layer0_outputs(5970));
    outputs(4419) <= (layer0_outputs(4993)) xor (layer0_outputs(3451));
    outputs(4420) <= layer0_outputs(50);
    outputs(4421) <= layer0_outputs(6590);
    outputs(4422) <= (layer0_outputs(1808)) and not (layer0_outputs(3096));
    outputs(4423) <= layer0_outputs(7338);
    outputs(4424) <= not(layer0_outputs(4007));
    outputs(4425) <= layer0_outputs(5416);
    outputs(4426) <= not(layer0_outputs(6316));
    outputs(4427) <= not((layer0_outputs(1819)) xor (layer0_outputs(6073)));
    outputs(4428) <= not(layer0_outputs(6774));
    outputs(4429) <= not(layer0_outputs(5779));
    outputs(4430) <= layer0_outputs(2378);
    outputs(4431) <= not(layer0_outputs(4943));
    outputs(4432) <= (layer0_outputs(4474)) or (layer0_outputs(6686));
    outputs(4433) <= layer0_outputs(3867);
    outputs(4434) <= not(layer0_outputs(3701));
    outputs(4435) <= (layer0_outputs(3970)) and not (layer0_outputs(1909));
    outputs(4436) <= not(layer0_outputs(3976)) or (layer0_outputs(3774));
    outputs(4437) <= not(layer0_outputs(4577));
    outputs(4438) <= layer0_outputs(1887);
    outputs(4439) <= not(layer0_outputs(1813));
    outputs(4440) <= layer0_outputs(755);
    outputs(4441) <= not(layer0_outputs(4921));
    outputs(4442) <= (layer0_outputs(5332)) xor (layer0_outputs(1415));
    outputs(4443) <= not(layer0_outputs(2348));
    outputs(4444) <= not((layer0_outputs(4023)) xor (layer0_outputs(1110)));
    outputs(4445) <= '0';
    outputs(4446) <= not((layer0_outputs(6375)) xor (layer0_outputs(6131)));
    outputs(4447) <= not(layer0_outputs(2664)) or (layer0_outputs(4076));
    outputs(4448) <= layer0_outputs(6906);
    outputs(4449) <= (layer0_outputs(1733)) and not (layer0_outputs(6537));
    outputs(4450) <= not((layer0_outputs(4856)) or (layer0_outputs(2129)));
    outputs(4451) <= not(layer0_outputs(6122));
    outputs(4452) <= not(layer0_outputs(7021));
    outputs(4453) <= layer0_outputs(775);
    outputs(4454) <= not((layer0_outputs(6891)) or (layer0_outputs(2689)));
    outputs(4455) <= not(layer0_outputs(4998));
    outputs(4456) <= (layer0_outputs(585)) xor (layer0_outputs(7196));
    outputs(4457) <= not((layer0_outputs(1752)) and (layer0_outputs(316)));
    outputs(4458) <= (layer0_outputs(3296)) and not (layer0_outputs(1777));
    outputs(4459) <= not(layer0_outputs(2647));
    outputs(4460) <= layer0_outputs(5840);
    outputs(4461) <= (layer0_outputs(5160)) xor (layer0_outputs(5022));
    outputs(4462) <= not((layer0_outputs(4708)) xor (layer0_outputs(4684)));
    outputs(4463) <= (layer0_outputs(3417)) xor (layer0_outputs(2881));
    outputs(4464) <= layer0_outputs(7480);
    outputs(4465) <= not((layer0_outputs(5673)) and (layer0_outputs(3298)));
    outputs(4466) <= not(layer0_outputs(1362));
    outputs(4467) <= (layer0_outputs(1490)) xor (layer0_outputs(4146));
    outputs(4468) <= (layer0_outputs(4756)) and not (layer0_outputs(5541));
    outputs(4469) <= (layer0_outputs(5338)) and not (layer0_outputs(4966));
    outputs(4470) <= not(layer0_outputs(7412));
    outputs(4471) <= not(layer0_outputs(1307));
    outputs(4472) <= not(layer0_outputs(4188)) or (layer0_outputs(130));
    outputs(4473) <= (layer0_outputs(7470)) and not (layer0_outputs(3786));
    outputs(4474) <= not(layer0_outputs(2868));
    outputs(4475) <= (layer0_outputs(1001)) or (layer0_outputs(1543));
    outputs(4476) <= not((layer0_outputs(835)) xor (layer0_outputs(3244)));
    outputs(4477) <= (layer0_outputs(6362)) xor (layer0_outputs(1599));
    outputs(4478) <= (layer0_outputs(1421)) and not (layer0_outputs(3381));
    outputs(4479) <= layer0_outputs(5416);
    outputs(4480) <= layer0_outputs(2757);
    outputs(4481) <= (layer0_outputs(5759)) and not (layer0_outputs(5542));
    outputs(4482) <= not(layer0_outputs(1052));
    outputs(4483) <= not(layer0_outputs(4093));
    outputs(4484) <= not(layer0_outputs(5224)) or (layer0_outputs(749));
    outputs(4485) <= not((layer0_outputs(837)) or (layer0_outputs(4841)));
    outputs(4486) <= not((layer0_outputs(6999)) xor (layer0_outputs(604)));
    outputs(4487) <= not((layer0_outputs(5148)) xor (layer0_outputs(4666)));
    outputs(4488) <= not((layer0_outputs(5069)) and (layer0_outputs(4209)));
    outputs(4489) <= (layer0_outputs(4550)) and not (layer0_outputs(3549));
    outputs(4490) <= not(layer0_outputs(3795)) or (layer0_outputs(82));
    outputs(4491) <= not((layer0_outputs(4478)) or (layer0_outputs(2668)));
    outputs(4492) <= not((layer0_outputs(578)) xor (layer0_outputs(1518)));
    outputs(4493) <= (layer0_outputs(3654)) and not (layer0_outputs(3678));
    outputs(4494) <= (layer0_outputs(2706)) xor (layer0_outputs(7026));
    outputs(4495) <= not(layer0_outputs(3832));
    outputs(4496) <= not(layer0_outputs(2390));
    outputs(4497) <= not(layer0_outputs(19));
    outputs(4498) <= (layer0_outputs(12)) and not (layer0_outputs(6348));
    outputs(4499) <= not(layer0_outputs(6366)) or (layer0_outputs(2587));
    outputs(4500) <= (layer0_outputs(1213)) xor (layer0_outputs(6524));
    outputs(4501) <= (layer0_outputs(308)) and (layer0_outputs(3651));
    outputs(4502) <= not(layer0_outputs(5069)) or (layer0_outputs(1552));
    outputs(4503) <= layer0_outputs(2580);
    outputs(4504) <= '1';
    outputs(4505) <= (layer0_outputs(4798)) and not (layer0_outputs(7389));
    outputs(4506) <= layer0_outputs(3845);
    outputs(4507) <= (layer0_outputs(7678)) xor (layer0_outputs(1685));
    outputs(4508) <= (layer0_outputs(63)) and not (layer0_outputs(2302));
    outputs(4509) <= (layer0_outputs(7101)) or (layer0_outputs(1375));
    outputs(4510) <= not((layer0_outputs(6982)) or (layer0_outputs(3512)));
    outputs(4511) <= not((layer0_outputs(1625)) xor (layer0_outputs(4325)));
    outputs(4512) <= not(layer0_outputs(7329)) or (layer0_outputs(3821));
    outputs(4513) <= not(layer0_outputs(3149)) or (layer0_outputs(3482));
    outputs(4514) <= layer0_outputs(2249);
    outputs(4515) <= (layer0_outputs(7229)) xor (layer0_outputs(3320));
    outputs(4516) <= not((layer0_outputs(5580)) xor (layer0_outputs(5190)));
    outputs(4517) <= (layer0_outputs(2798)) xor (layer0_outputs(1523));
    outputs(4518) <= (layer0_outputs(4225)) xor (layer0_outputs(5079));
    outputs(4519) <= not((layer0_outputs(873)) xor (layer0_outputs(1430)));
    outputs(4520) <= layer0_outputs(866);
    outputs(4521) <= not((layer0_outputs(649)) or (layer0_outputs(3650)));
    outputs(4522) <= (layer0_outputs(1333)) and not (layer0_outputs(2717));
    outputs(4523) <= layer0_outputs(5849);
    outputs(4524) <= (layer0_outputs(945)) xor (layer0_outputs(1646));
    outputs(4525) <= not((layer0_outputs(6371)) xor (layer0_outputs(1100)));
    outputs(4526) <= layer0_outputs(2912);
    outputs(4527) <= not(layer0_outputs(2151)) or (layer0_outputs(2458));
    outputs(4528) <= layer0_outputs(229);
    outputs(4529) <= (layer0_outputs(2143)) and (layer0_outputs(3541));
    outputs(4530) <= layer0_outputs(1546);
    outputs(4531) <= not(layer0_outputs(1662));
    outputs(4532) <= (layer0_outputs(5213)) or (layer0_outputs(3653));
    outputs(4533) <= layer0_outputs(912);
    outputs(4534) <= not(layer0_outputs(3376));
    outputs(4535) <= not(layer0_outputs(563));
    outputs(4536) <= not(layer0_outputs(3208)) or (layer0_outputs(3148));
    outputs(4537) <= (layer0_outputs(2511)) xor (layer0_outputs(175));
    outputs(4538) <= not((layer0_outputs(7487)) xor (layer0_outputs(4142)));
    outputs(4539) <= (layer0_outputs(5078)) and not (layer0_outputs(838));
    outputs(4540) <= not(layer0_outputs(5753));
    outputs(4541) <= (layer0_outputs(2584)) xor (layer0_outputs(5170));
    outputs(4542) <= (layer0_outputs(5713)) or (layer0_outputs(6947));
    outputs(4543) <= not(layer0_outputs(5920));
    outputs(4544) <= not(layer0_outputs(887));
    outputs(4545) <= not(layer0_outputs(6692));
    outputs(4546) <= not(layer0_outputs(545));
    outputs(4547) <= not((layer0_outputs(4757)) or (layer0_outputs(4761)));
    outputs(4548) <= (layer0_outputs(5074)) and not (layer0_outputs(702));
    outputs(4549) <= not(layer0_outputs(2577)) or (layer0_outputs(1793));
    outputs(4550) <= layer0_outputs(6833);
    outputs(4551) <= not((layer0_outputs(1492)) or (layer0_outputs(3581)));
    outputs(4552) <= not((layer0_outputs(2279)) and (layer0_outputs(5455)));
    outputs(4553) <= (layer0_outputs(3692)) xor (layer0_outputs(423));
    outputs(4554) <= layer0_outputs(4596);
    outputs(4555) <= not(layer0_outputs(1268));
    outputs(4556) <= not(layer0_outputs(6410));
    outputs(4557) <= (layer0_outputs(3)) xor (layer0_outputs(3324));
    outputs(4558) <= (layer0_outputs(1503)) or (layer0_outputs(4880));
    outputs(4559) <= layer0_outputs(3074);
    outputs(4560) <= not((layer0_outputs(5756)) xor (layer0_outputs(1500)));
    outputs(4561) <= (layer0_outputs(6716)) xor (layer0_outputs(4929));
    outputs(4562) <= not((layer0_outputs(3969)) xor (layer0_outputs(4505)));
    outputs(4563) <= not((layer0_outputs(3583)) xor (layer0_outputs(852)));
    outputs(4564) <= not((layer0_outputs(5566)) xor (layer0_outputs(6472)));
    outputs(4565) <= layer0_outputs(6754);
    outputs(4566) <= not((layer0_outputs(4832)) and (layer0_outputs(7655)));
    outputs(4567) <= not(layer0_outputs(4760));
    outputs(4568) <= (layer0_outputs(3562)) xor (layer0_outputs(6814));
    outputs(4569) <= not(layer0_outputs(3936));
    outputs(4570) <= not((layer0_outputs(1420)) or (layer0_outputs(671)));
    outputs(4571) <= not((layer0_outputs(1667)) or (layer0_outputs(5054)));
    outputs(4572) <= not(layer0_outputs(6379));
    outputs(4573) <= not((layer0_outputs(2855)) and (layer0_outputs(3177)));
    outputs(4574) <= layer0_outputs(5773);
    outputs(4575) <= not(layer0_outputs(6636)) or (layer0_outputs(1371));
    outputs(4576) <= (layer0_outputs(5793)) and (layer0_outputs(5095));
    outputs(4577) <= layer0_outputs(1383);
    outputs(4578) <= not(layer0_outputs(5310)) or (layer0_outputs(2211));
    outputs(4579) <= not((layer0_outputs(3670)) or (layer0_outputs(2819)));
    outputs(4580) <= not((layer0_outputs(6842)) and (layer0_outputs(1392)));
    outputs(4581) <= not(layer0_outputs(3431)) or (layer0_outputs(5399));
    outputs(4582) <= (layer0_outputs(3223)) xor (layer0_outputs(2677));
    outputs(4583) <= not(layer0_outputs(5016));
    outputs(4584) <= (layer0_outputs(229)) or (layer0_outputs(4759));
    outputs(4585) <= layer0_outputs(7289);
    outputs(4586) <= layer0_outputs(5340);
    outputs(4587) <= not(layer0_outputs(2152));
    outputs(4588) <= (layer0_outputs(6729)) xor (layer0_outputs(4729));
    outputs(4589) <= not((layer0_outputs(3503)) xor (layer0_outputs(1292)));
    outputs(4590) <= layer0_outputs(3263);
    outputs(4591) <= layer0_outputs(4674);
    outputs(4592) <= layer0_outputs(6724);
    outputs(4593) <= layer0_outputs(506);
    outputs(4594) <= (layer0_outputs(4586)) and (layer0_outputs(6468));
    outputs(4595) <= (layer0_outputs(1476)) and not (layer0_outputs(6962));
    outputs(4596) <= not((layer0_outputs(258)) or (layer0_outputs(5555)));
    outputs(4597) <= not((layer0_outputs(1122)) xor (layer0_outputs(3677)));
    outputs(4598) <= not(layer0_outputs(1728));
    outputs(4599) <= layer0_outputs(5021);
    outputs(4600) <= (layer0_outputs(6559)) and not (layer0_outputs(7493));
    outputs(4601) <= layer0_outputs(458);
    outputs(4602) <= not(layer0_outputs(4318));
    outputs(4603) <= (layer0_outputs(4418)) or (layer0_outputs(4494));
    outputs(4604) <= not(layer0_outputs(594));
    outputs(4605) <= not((layer0_outputs(5358)) xor (layer0_outputs(371)));
    outputs(4606) <= not((layer0_outputs(345)) xor (layer0_outputs(3416)));
    outputs(4607) <= (layer0_outputs(930)) or (layer0_outputs(7263));
    outputs(4608) <= layer0_outputs(2641);
    outputs(4609) <= not(layer0_outputs(6339));
    outputs(4610) <= not((layer0_outputs(6757)) xor (layer0_outputs(3660)));
    outputs(4611) <= (layer0_outputs(4943)) xor (layer0_outputs(3345));
    outputs(4612) <= layer0_outputs(6859);
    outputs(4613) <= (layer0_outputs(1261)) xor (layer0_outputs(6467));
    outputs(4614) <= not((layer0_outputs(627)) and (layer0_outputs(5611)));
    outputs(4615) <= '1';
    outputs(4616) <= not(layer0_outputs(540));
    outputs(4617) <= not((layer0_outputs(4354)) xor (layer0_outputs(1110)));
    outputs(4618) <= not(layer0_outputs(1255)) or (layer0_outputs(5935));
    outputs(4619) <= layer0_outputs(4464);
    outputs(4620) <= not((layer0_outputs(6415)) xor (layer0_outputs(5926)));
    outputs(4621) <= (layer0_outputs(5195)) xor (layer0_outputs(1221));
    outputs(4622) <= not((layer0_outputs(3487)) and (layer0_outputs(4379)));
    outputs(4623) <= not(layer0_outputs(3245));
    outputs(4624) <= not(layer0_outputs(30));
    outputs(4625) <= not((layer0_outputs(896)) xor (layer0_outputs(2336)));
    outputs(4626) <= (layer0_outputs(2759)) xor (layer0_outputs(6279));
    outputs(4627) <= not((layer0_outputs(1958)) xor (layer0_outputs(3992)));
    outputs(4628) <= not((layer0_outputs(1217)) or (layer0_outputs(2322)));
    outputs(4629) <= not((layer0_outputs(7443)) and (layer0_outputs(3944)));
    outputs(4630) <= layer0_outputs(2049);
    outputs(4631) <= layer0_outputs(3664);
    outputs(4632) <= layer0_outputs(477);
    outputs(4633) <= layer0_outputs(3884);
    outputs(4634) <= not(layer0_outputs(6445));
    outputs(4635) <= layer0_outputs(172);
    outputs(4636) <= (layer0_outputs(2216)) or (layer0_outputs(3447));
    outputs(4637) <= (layer0_outputs(3950)) and not (layer0_outputs(638));
    outputs(4638) <= (layer0_outputs(2922)) or (layer0_outputs(1082));
    outputs(4639) <= layer0_outputs(5344);
    outputs(4640) <= (layer0_outputs(1822)) and (layer0_outputs(3561));
    outputs(4641) <= (layer0_outputs(4125)) and (layer0_outputs(2707));
    outputs(4642) <= not(layer0_outputs(849));
    outputs(4643) <= (layer0_outputs(6680)) and not (layer0_outputs(4343));
    outputs(4644) <= not((layer0_outputs(612)) or (layer0_outputs(4738)));
    outputs(4645) <= not(layer0_outputs(5902)) or (layer0_outputs(3895));
    outputs(4646) <= not(layer0_outputs(5776));
    outputs(4647) <= not((layer0_outputs(6549)) xor (layer0_outputs(2422)));
    outputs(4648) <= not(layer0_outputs(5609));
    outputs(4649) <= (layer0_outputs(4707)) xor (layer0_outputs(5316));
    outputs(4650) <= not(layer0_outputs(4078)) or (layer0_outputs(5719));
    outputs(4651) <= not(layer0_outputs(6138));
    outputs(4652) <= not(layer0_outputs(7177));
    outputs(4653) <= not(layer0_outputs(6356));
    outputs(4654) <= (layer0_outputs(4533)) or (layer0_outputs(3542));
    outputs(4655) <= (layer0_outputs(2096)) and not (layer0_outputs(6012));
    outputs(4656) <= not(layer0_outputs(4124));
    outputs(4657) <= not(layer0_outputs(4380)) or (layer0_outputs(1599));
    outputs(4658) <= layer0_outputs(1753);
    outputs(4659) <= (layer0_outputs(1079)) and (layer0_outputs(6835));
    outputs(4660) <= not(layer0_outputs(642));
    outputs(4661) <= not(layer0_outputs(4273)) or (layer0_outputs(6202));
    outputs(4662) <= layer0_outputs(1803);
    outputs(4663) <= not((layer0_outputs(4166)) xor (layer0_outputs(5747)));
    outputs(4664) <= layer0_outputs(7111);
    outputs(4665) <= layer0_outputs(4439);
    outputs(4666) <= not(layer0_outputs(219));
    outputs(4667) <= (layer0_outputs(4216)) and not (layer0_outputs(3960));
    outputs(4668) <= (layer0_outputs(2400)) xor (layer0_outputs(1308));
    outputs(4669) <= (layer0_outputs(3553)) and (layer0_outputs(3565));
    outputs(4670) <= layer0_outputs(5732);
    outputs(4671) <= not(layer0_outputs(2992));
    outputs(4672) <= (layer0_outputs(907)) and not (layer0_outputs(534));
    outputs(4673) <= layer0_outputs(5687);
    outputs(4674) <= (layer0_outputs(7204)) or (layer0_outputs(6535));
    outputs(4675) <= layer0_outputs(2888);
    outputs(4676) <= layer0_outputs(7190);
    outputs(4677) <= (layer0_outputs(1859)) or (layer0_outputs(62));
    outputs(4678) <= (layer0_outputs(1580)) and not (layer0_outputs(6413));
    outputs(4679) <= not(layer0_outputs(4999)) or (layer0_outputs(3437));
    outputs(4680) <= (layer0_outputs(3650)) xor (layer0_outputs(1136));
    outputs(4681) <= not(layer0_outputs(5586));
    outputs(4682) <= not(layer0_outputs(3873)) or (layer0_outputs(2083));
    outputs(4683) <= layer0_outputs(2619);
    outputs(4684) <= not(layer0_outputs(6364));
    outputs(4685) <= not((layer0_outputs(5806)) or (layer0_outputs(1509)));
    outputs(4686) <= not(layer0_outputs(3628));
    outputs(4687) <= layer0_outputs(3897);
    outputs(4688) <= not(layer0_outputs(4355));
    outputs(4689) <= not(layer0_outputs(2009));
    outputs(4690) <= not(layer0_outputs(2712));
    outputs(4691) <= not(layer0_outputs(2738));
    outputs(4692) <= not(layer0_outputs(2565)) or (layer0_outputs(2056));
    outputs(4693) <= layer0_outputs(1325);
    outputs(4694) <= layer0_outputs(2519);
    outputs(4695) <= layer0_outputs(5639);
    outputs(4696) <= not(layer0_outputs(7289)) or (layer0_outputs(5066));
    outputs(4697) <= (layer0_outputs(3461)) xor (layer0_outputs(4036));
    outputs(4698) <= (layer0_outputs(1627)) xor (layer0_outputs(6343));
    outputs(4699) <= (layer0_outputs(3363)) and not (layer0_outputs(6445));
    outputs(4700) <= not(layer0_outputs(2323));
    outputs(4701) <= not((layer0_outputs(3930)) xor (layer0_outputs(5517)));
    outputs(4702) <= layer0_outputs(4648);
    outputs(4703) <= not(layer0_outputs(241));
    outputs(4704) <= not(layer0_outputs(469));
    outputs(4705) <= (layer0_outputs(616)) xor (layer0_outputs(5493));
    outputs(4706) <= layer0_outputs(3049);
    outputs(4707) <= layer0_outputs(859);
    outputs(4708) <= not(layer0_outputs(5668));
    outputs(4709) <= not((layer0_outputs(3992)) or (layer0_outputs(7625)));
    outputs(4710) <= (layer0_outputs(886)) xor (layer0_outputs(7400));
    outputs(4711) <= (layer0_outputs(6210)) and not (layer0_outputs(2836));
    outputs(4712) <= layer0_outputs(2751);
    outputs(4713) <= layer0_outputs(2646);
    outputs(4714) <= (layer0_outputs(4439)) and not (layer0_outputs(7548));
    outputs(4715) <= (layer0_outputs(5996)) and (layer0_outputs(840));
    outputs(4716) <= layer0_outputs(3663);
    outputs(4717) <= layer0_outputs(154);
    outputs(4718) <= layer0_outputs(4844);
    outputs(4719) <= (layer0_outputs(2472)) and (layer0_outputs(6967));
    outputs(4720) <= layer0_outputs(15);
    outputs(4721) <= layer0_outputs(4450);
    outputs(4722) <= not(layer0_outputs(3967));
    outputs(4723) <= not(layer0_outputs(2006)) or (layer0_outputs(3649));
    outputs(4724) <= (layer0_outputs(352)) and (layer0_outputs(4457));
    outputs(4725) <= (layer0_outputs(7288)) xor (layer0_outputs(3481));
    outputs(4726) <= not((layer0_outputs(3872)) xor (layer0_outputs(6044)));
    outputs(4727) <= (layer0_outputs(4681)) or (layer0_outputs(1318));
    outputs(4728) <= layer0_outputs(3707);
    outputs(4729) <= layer0_outputs(4235);
    outputs(4730) <= (layer0_outputs(5874)) xor (layer0_outputs(5809));
    outputs(4731) <= not(layer0_outputs(2793));
    outputs(4732) <= (layer0_outputs(6828)) and not (layer0_outputs(5173));
    outputs(4733) <= not((layer0_outputs(6226)) xor (layer0_outputs(16)));
    outputs(4734) <= layer0_outputs(7151);
    outputs(4735) <= layer0_outputs(3127);
    outputs(4736) <= (layer0_outputs(5977)) xor (layer0_outputs(803));
    outputs(4737) <= not(layer0_outputs(7413));
    outputs(4738) <= layer0_outputs(2650);
    outputs(4739) <= not(layer0_outputs(1064));
    outputs(4740) <= not(layer0_outputs(3366));
    outputs(4741) <= layer0_outputs(4811);
    outputs(4742) <= not(layer0_outputs(5754));
    outputs(4743) <= not((layer0_outputs(178)) xor (layer0_outputs(2496)));
    outputs(4744) <= not(layer0_outputs(831)) or (layer0_outputs(1736));
    outputs(4745) <= (layer0_outputs(5516)) and not (layer0_outputs(5844));
    outputs(4746) <= not((layer0_outputs(3155)) xor (layer0_outputs(5579)));
    outputs(4747) <= layer0_outputs(1479);
    outputs(4748) <= not((layer0_outputs(6607)) xor (layer0_outputs(7475)));
    outputs(4749) <= not(layer0_outputs(5958));
    outputs(4750) <= not((layer0_outputs(5927)) xor (layer0_outputs(4688)));
    outputs(4751) <= not((layer0_outputs(5226)) or (layer0_outputs(1394)));
    outputs(4752) <= (layer0_outputs(5479)) and (layer0_outputs(5231));
    outputs(4753) <= layer0_outputs(6276);
    outputs(4754) <= not((layer0_outputs(4585)) or (layer0_outputs(2555)));
    outputs(4755) <= layer0_outputs(7264);
    outputs(4756) <= not(layer0_outputs(945));
    outputs(4757) <= not(layer0_outputs(7543));
    outputs(4758) <= not((layer0_outputs(3696)) and (layer0_outputs(2564)));
    outputs(4759) <= layer0_outputs(4805);
    outputs(4760) <= not(layer0_outputs(215));
    outputs(4761) <= (layer0_outputs(563)) and not (layer0_outputs(5091));
    outputs(4762) <= not(layer0_outputs(694));
    outputs(4763) <= layer0_outputs(2554);
    outputs(4764) <= not(layer0_outputs(3402));
    outputs(4765) <= (layer0_outputs(1979)) and not (layer0_outputs(783));
    outputs(4766) <= layer0_outputs(7676);
    outputs(4767) <= not(layer0_outputs(5147)) or (layer0_outputs(4879));
    outputs(4768) <= not(layer0_outputs(850));
    outputs(4769) <= not((layer0_outputs(4835)) xor (layer0_outputs(2420)));
    outputs(4770) <= layer0_outputs(3247);
    outputs(4771) <= layer0_outputs(4495);
    outputs(4772) <= not(layer0_outputs(4205));
    outputs(4773) <= not(layer0_outputs(3840));
    outputs(4774) <= not(layer0_outputs(7148));
    outputs(4775) <= layer0_outputs(7137);
    outputs(4776) <= not((layer0_outputs(7379)) or (layer0_outputs(5505)));
    outputs(4777) <= not((layer0_outputs(479)) and (layer0_outputs(3375)));
    outputs(4778) <= not((layer0_outputs(4488)) xor (layer0_outputs(1348)));
    outputs(4779) <= not((layer0_outputs(3597)) and (layer0_outputs(4560)));
    outputs(4780) <= not(layer0_outputs(3703));
    outputs(4781) <= not(layer0_outputs(6724));
    outputs(4782) <= not(layer0_outputs(4711));
    outputs(4783) <= layer0_outputs(7137);
    outputs(4784) <= layer0_outputs(3128);
    outputs(4785) <= not((layer0_outputs(2031)) xor (layer0_outputs(3311)));
    outputs(4786) <= (layer0_outputs(5940)) and (layer0_outputs(5991));
    outputs(4787) <= not(layer0_outputs(1554));
    outputs(4788) <= not((layer0_outputs(831)) xor (layer0_outputs(6019)));
    outputs(4789) <= not((layer0_outputs(138)) and (layer0_outputs(635)));
    outputs(4790) <= layer0_outputs(2302);
    outputs(4791) <= layer0_outputs(5918);
    outputs(4792) <= (layer0_outputs(2764)) and not (layer0_outputs(48));
    outputs(4793) <= not((layer0_outputs(3092)) or (layer0_outputs(2087)));
    outputs(4794) <= not((layer0_outputs(5705)) or (layer0_outputs(1917)));
    outputs(4795) <= (layer0_outputs(2363)) and not (layer0_outputs(100));
    outputs(4796) <= not(layer0_outputs(387));
    outputs(4797) <= '0';
    outputs(4798) <= not(layer0_outputs(4161));
    outputs(4799) <= not((layer0_outputs(6450)) xor (layer0_outputs(542)));
    outputs(4800) <= (layer0_outputs(6966)) and not (layer0_outputs(1135));
    outputs(4801) <= layer0_outputs(310);
    outputs(4802) <= (layer0_outputs(364)) or (layer0_outputs(2150));
    outputs(4803) <= not((layer0_outputs(6528)) or (layer0_outputs(6296)));
    outputs(4804) <= not((layer0_outputs(2153)) or (layer0_outputs(61)));
    outputs(4805) <= layer0_outputs(3122);
    outputs(4806) <= layer0_outputs(7278);
    outputs(4807) <= layer0_outputs(2757);
    outputs(4808) <= not(layer0_outputs(4546));
    outputs(4809) <= (layer0_outputs(5910)) and not (layer0_outputs(790));
    outputs(4810) <= layer0_outputs(3805);
    outputs(4811) <= layer0_outputs(5986);
    outputs(4812) <= not(layer0_outputs(2910));
    outputs(4813) <= not((layer0_outputs(1379)) or (layer0_outputs(2323)));
    outputs(4814) <= not(layer0_outputs(3984));
    outputs(4815) <= not(layer0_outputs(3559));
    outputs(4816) <= layer0_outputs(6194);
    outputs(4817) <= layer0_outputs(5353);
    outputs(4818) <= (layer0_outputs(5252)) and (layer0_outputs(3403));
    outputs(4819) <= not(layer0_outputs(5528));
    outputs(4820) <= (layer0_outputs(5282)) and not (layer0_outputs(5031));
    outputs(4821) <= (layer0_outputs(5716)) xor (layer0_outputs(4038));
    outputs(4822) <= not(layer0_outputs(3582));
    outputs(4823) <= layer0_outputs(4649);
    outputs(4824) <= layer0_outputs(350);
    outputs(4825) <= not((layer0_outputs(961)) or (layer0_outputs(5075)));
    outputs(4826) <= (layer0_outputs(7426)) xor (layer0_outputs(7643));
    outputs(4827) <= layer0_outputs(1760);
    outputs(4828) <= layer0_outputs(7002);
    outputs(4829) <= not((layer0_outputs(6037)) xor (layer0_outputs(2096)));
    outputs(4830) <= not(layer0_outputs(1376));
    outputs(4831) <= not(layer0_outputs(3131));
    outputs(4832) <= layer0_outputs(2670);
    outputs(4833) <= not(layer0_outputs(524));
    outputs(4834) <= not((layer0_outputs(5637)) and (layer0_outputs(2050)));
    outputs(4835) <= not((layer0_outputs(6397)) xor (layer0_outputs(6243)));
    outputs(4836) <= (layer0_outputs(2658)) xor (layer0_outputs(1511));
    outputs(4837) <= not((layer0_outputs(5030)) and (layer0_outputs(1307)));
    outputs(4838) <= not(layer0_outputs(2276));
    outputs(4839) <= (layer0_outputs(6664)) xor (layer0_outputs(5133));
    outputs(4840) <= not(layer0_outputs(5202));
    outputs(4841) <= not(layer0_outputs(6307));
    outputs(4842) <= not(layer0_outputs(1553));
    outputs(4843) <= not(layer0_outputs(256)) or (layer0_outputs(6893));
    outputs(4844) <= not(layer0_outputs(4841));
    outputs(4845) <= not(layer0_outputs(895));
    outputs(4846) <= not(layer0_outputs(7055)) or (layer0_outputs(5790));
    outputs(4847) <= not(layer0_outputs(6314));
    outputs(4848) <= not(layer0_outputs(5381));
    outputs(4849) <= (layer0_outputs(4006)) and not (layer0_outputs(6011));
    outputs(4850) <= (layer0_outputs(323)) and (layer0_outputs(5697));
    outputs(4851) <= not(layer0_outputs(7035));
    outputs(4852) <= not(layer0_outputs(1277));
    outputs(4853) <= (layer0_outputs(1647)) and not (layer0_outputs(2727));
    outputs(4854) <= not(layer0_outputs(5151));
    outputs(4855) <= not(layer0_outputs(2162));
    outputs(4856) <= layer0_outputs(1216);
    outputs(4857) <= not(layer0_outputs(6353));
    outputs(4858) <= layer0_outputs(4712);
    outputs(4859) <= (layer0_outputs(3991)) xor (layer0_outputs(4465));
    outputs(4860) <= (layer0_outputs(2986)) and not (layer0_outputs(3626));
    outputs(4861) <= not(layer0_outputs(3310));
    outputs(4862) <= not(layer0_outputs(6567));
    outputs(4863) <= layer0_outputs(5787);
    outputs(4864) <= layer0_outputs(235);
    outputs(4865) <= layer0_outputs(293);
    outputs(4866) <= layer0_outputs(975);
    outputs(4867) <= (layer0_outputs(1427)) and (layer0_outputs(4082));
    outputs(4868) <= not(layer0_outputs(7025)) or (layer0_outputs(7354));
    outputs(4869) <= (layer0_outputs(6302)) and not (layer0_outputs(5380));
    outputs(4870) <= (layer0_outputs(3452)) and not (layer0_outputs(1827));
    outputs(4871) <= layer0_outputs(2443);
    outputs(4872) <= layer0_outputs(884);
    outputs(4873) <= not((layer0_outputs(6569)) xor (layer0_outputs(3794)));
    outputs(4874) <= not(layer0_outputs(7633));
    outputs(4875) <= not(layer0_outputs(6695));
    outputs(4876) <= layer0_outputs(397);
    outputs(4877) <= not(layer0_outputs(1484));
    outputs(4878) <= not(layer0_outputs(2941));
    outputs(4879) <= not(layer0_outputs(4976));
    outputs(4880) <= (layer0_outputs(3286)) xor (layer0_outputs(4331));
    outputs(4881) <= not((layer0_outputs(3436)) xor (layer0_outputs(4088)));
    outputs(4882) <= not((layer0_outputs(6646)) xor (layer0_outputs(1951)));
    outputs(4883) <= (layer0_outputs(4214)) xor (layer0_outputs(7300));
    outputs(4884) <= (layer0_outputs(4675)) xor (layer0_outputs(2151));
    outputs(4885) <= not(layer0_outputs(7362)) or (layer0_outputs(4059));
    outputs(4886) <= not(layer0_outputs(5351));
    outputs(4887) <= not(layer0_outputs(7464));
    outputs(4888) <= not(layer0_outputs(6804));
    outputs(4889) <= layer0_outputs(2119);
    outputs(4890) <= not(layer0_outputs(2449));
    outputs(4891) <= not(layer0_outputs(4121));
    outputs(4892) <= not(layer0_outputs(2464));
    outputs(4893) <= layer0_outputs(255);
    outputs(4894) <= not(layer0_outputs(531)) or (layer0_outputs(5471));
    outputs(4895) <= (layer0_outputs(3545)) and not (layer0_outputs(4098));
    outputs(4896) <= not((layer0_outputs(5175)) xor (layer0_outputs(3327)));
    outputs(4897) <= not((layer0_outputs(6851)) xor (layer0_outputs(1445)));
    outputs(4898) <= not(layer0_outputs(169));
    outputs(4899) <= (layer0_outputs(922)) and not (layer0_outputs(5852));
    outputs(4900) <= (layer0_outputs(5578)) and not (layer0_outputs(5557));
    outputs(4901) <= (layer0_outputs(401)) xor (layer0_outputs(3316));
    outputs(4902) <= (layer0_outputs(1182)) xor (layer0_outputs(446));
    outputs(4903) <= layer0_outputs(6055);
    outputs(4904) <= (layer0_outputs(2507)) and (layer0_outputs(4957));
    outputs(4905) <= layer0_outputs(7594);
    outputs(4906) <= layer0_outputs(4267);
    outputs(4907) <= not((layer0_outputs(6617)) and (layer0_outputs(5626)));
    outputs(4908) <= layer0_outputs(5396);
    outputs(4909) <= (layer0_outputs(3615)) xor (layer0_outputs(5463));
    outputs(4910) <= (layer0_outputs(860)) xor (layer0_outputs(3551));
    outputs(4911) <= (layer0_outputs(3643)) and not (layer0_outputs(4827));
    outputs(4912) <= not(layer0_outputs(928));
    outputs(4913) <= not((layer0_outputs(110)) and (layer0_outputs(6127)));
    outputs(4914) <= not(layer0_outputs(1065)) or (layer0_outputs(671));
    outputs(4915) <= (layer0_outputs(2374)) and not (layer0_outputs(4496));
    outputs(4916) <= not((layer0_outputs(1341)) and (layer0_outputs(6293)));
    outputs(4917) <= (layer0_outputs(7260)) and not (layer0_outputs(7583));
    outputs(4918) <= (layer0_outputs(2691)) and (layer0_outputs(4011));
    outputs(4919) <= layer0_outputs(2497);
    outputs(4920) <= not(layer0_outputs(4935));
    outputs(4921) <= layer0_outputs(4731);
    outputs(4922) <= not(layer0_outputs(5035));
    outputs(4923) <= not((layer0_outputs(606)) xor (layer0_outputs(3797)));
    outputs(4924) <= not(layer0_outputs(1756));
    outputs(4925) <= layer0_outputs(6809);
    outputs(4926) <= (layer0_outputs(3337)) and (layer0_outputs(3137));
    outputs(4927) <= (layer0_outputs(4322)) and not (layer0_outputs(492));
    outputs(4928) <= not(layer0_outputs(5398));
    outputs(4929) <= not(layer0_outputs(6045));
    outputs(4930) <= layer0_outputs(4434);
    outputs(4931) <= layer0_outputs(7067);
    outputs(4932) <= (layer0_outputs(6212)) or (layer0_outputs(5946));
    outputs(4933) <= not((layer0_outputs(6100)) and (layer0_outputs(1502)));
    outputs(4934) <= layer0_outputs(5922);
    outputs(4935) <= layer0_outputs(6035);
    outputs(4936) <= layer0_outputs(1839);
    outputs(4937) <= (layer0_outputs(3180)) and not (layer0_outputs(3550));
    outputs(4938) <= not((layer0_outputs(3623)) xor (layer0_outputs(1899)));
    outputs(4939) <= layer0_outputs(6490);
    outputs(4940) <= layer0_outputs(422);
    outputs(4941) <= layer0_outputs(4454);
    outputs(4942) <= not(layer0_outputs(596));
    outputs(4943) <= not(layer0_outputs(3519));
    outputs(4944) <= (layer0_outputs(7090)) and not (layer0_outputs(4056));
    outputs(4945) <= layer0_outputs(5011);
    outputs(4946) <= (layer0_outputs(6512)) and not (layer0_outputs(5952));
    outputs(4947) <= not(layer0_outputs(325));
    outputs(4948) <= layer0_outputs(1271);
    outputs(4949) <= (layer0_outputs(3954)) and not (layer0_outputs(7079));
    outputs(4950) <= not(layer0_outputs(4559));
    outputs(4951) <= not((layer0_outputs(5183)) and (layer0_outputs(794)));
    outputs(4952) <= not(layer0_outputs(1841)) or (layer0_outputs(6808));
    outputs(4953) <= not(layer0_outputs(1380));
    outputs(4954) <= (layer0_outputs(2418)) xor (layer0_outputs(7425));
    outputs(4955) <= (layer0_outputs(6628)) and not (layer0_outputs(4208));
    outputs(4956) <= layer0_outputs(6898);
    outputs(4957) <= not(layer0_outputs(3260));
    outputs(4958) <= not((layer0_outputs(2864)) or (layer0_outputs(610)));
    outputs(4959) <= layer0_outputs(1787);
    outputs(4960) <= layer0_outputs(2956);
    outputs(4961) <= not((layer0_outputs(6319)) or (layer0_outputs(6769)));
    outputs(4962) <= layer0_outputs(696);
    outputs(4963) <= (layer0_outputs(5230)) or (layer0_outputs(5456));
    outputs(4964) <= not(layer0_outputs(6118));
    outputs(4965) <= not((layer0_outputs(1312)) and (layer0_outputs(5146)));
    outputs(4966) <= layer0_outputs(3182);
    outputs(4967) <= layer0_outputs(2585);
    outputs(4968) <= layer0_outputs(2542);
    outputs(4969) <= layer0_outputs(6521);
    outputs(4970) <= not(layer0_outputs(6873));
    outputs(4971) <= (layer0_outputs(182)) and not (layer0_outputs(4389));
    outputs(4972) <= (layer0_outputs(3339)) and not (layer0_outputs(2317));
    outputs(4973) <= layer0_outputs(3533);
    outputs(4974) <= not((layer0_outputs(5059)) and (layer0_outputs(4705)));
    outputs(4975) <= not((layer0_outputs(3246)) xor (layer0_outputs(5495)));
    outputs(4976) <= layer0_outputs(5728);
    outputs(4977) <= layer0_outputs(5937);
    outputs(4978) <= (layer0_outputs(1147)) and not (layer0_outputs(3409));
    outputs(4979) <= layer0_outputs(6152);
    outputs(4980) <= not((layer0_outputs(920)) xor (layer0_outputs(4196)));
    outputs(4981) <= not((layer0_outputs(56)) or (layer0_outputs(6612)));
    outputs(4982) <= not(layer0_outputs(6250));
    outputs(4983) <= layer0_outputs(5572);
    outputs(4984) <= not((layer0_outputs(6550)) xor (layer0_outputs(5907)));
    outputs(4985) <= (layer0_outputs(7642)) xor (layer0_outputs(4617));
    outputs(4986) <= (layer0_outputs(2430)) and not (layer0_outputs(3164));
    outputs(4987) <= not(layer0_outputs(6426)) or (layer0_outputs(1890));
    outputs(4988) <= (layer0_outputs(1933)) and (layer0_outputs(6182));
    outputs(4989) <= not(layer0_outputs(1709));
    outputs(4990) <= not((layer0_outputs(781)) xor (layer0_outputs(1038)));
    outputs(4991) <= not((layer0_outputs(5358)) xor (layer0_outputs(807)));
    outputs(4992) <= not(layer0_outputs(163));
    outputs(4993) <= not((layer0_outputs(3148)) or (layer0_outputs(7341)));
    outputs(4994) <= layer0_outputs(777);
    outputs(4995) <= not((layer0_outputs(6507)) or (layer0_outputs(3531)));
    outputs(4996) <= not(layer0_outputs(3442));
    outputs(4997) <= (layer0_outputs(3880)) xor (layer0_outputs(6540));
    outputs(4998) <= (layer0_outputs(83)) and not (layer0_outputs(1203));
    outputs(4999) <= layer0_outputs(2294);
    outputs(5000) <= not(layer0_outputs(7240));
    outputs(5001) <= (layer0_outputs(3007)) xor (layer0_outputs(1780));
    outputs(5002) <= (layer0_outputs(2005)) xor (layer0_outputs(5706));
    outputs(5003) <= not((layer0_outputs(3178)) and (layer0_outputs(1652)));
    outputs(5004) <= layer0_outputs(1428);
    outputs(5005) <= layer0_outputs(4703);
    outputs(5006) <= (layer0_outputs(1043)) xor (layer0_outputs(1439));
    outputs(5007) <= (layer0_outputs(719)) xor (layer0_outputs(5758));
    outputs(5008) <= not((layer0_outputs(2674)) xor (layer0_outputs(5081)));
    outputs(5009) <= not(layer0_outputs(5911));
    outputs(5010) <= not(layer0_outputs(6669));
    outputs(5011) <= layer0_outputs(6732);
    outputs(5012) <= (layer0_outputs(1850)) and (layer0_outputs(5915));
    outputs(5013) <= not(layer0_outputs(6984));
    outputs(5014) <= layer0_outputs(4096);
    outputs(5015) <= (layer0_outputs(4153)) and (layer0_outputs(1010));
    outputs(5016) <= not(layer0_outputs(7671));
    outputs(5017) <= (layer0_outputs(2082)) and not (layer0_outputs(1311));
    outputs(5018) <= not(layer0_outputs(3953));
    outputs(5019) <= not(layer0_outputs(3040));
    outputs(5020) <= not((layer0_outputs(3070)) or (layer0_outputs(6536)));
    outputs(5021) <= layer0_outputs(193);
    outputs(5022) <= (layer0_outputs(980)) xor (layer0_outputs(771));
    outputs(5023) <= layer0_outputs(5396);
    outputs(5024) <= layer0_outputs(5373);
    outputs(5025) <= not(layer0_outputs(2588));
    outputs(5026) <= not((layer0_outputs(7558)) or (layer0_outputs(6527)));
    outputs(5027) <= (layer0_outputs(4990)) and (layer0_outputs(3837));
    outputs(5028) <= layer0_outputs(4074);
    outputs(5029) <= not(layer0_outputs(1795));
    outputs(5030) <= (layer0_outputs(1447)) xor (layer0_outputs(1193));
    outputs(5031) <= not((layer0_outputs(4642)) or (layer0_outputs(184)));
    outputs(5032) <= layer0_outputs(4462);
    outputs(5033) <= not((layer0_outputs(6646)) or (layer0_outputs(6734)));
    outputs(5034) <= not(layer0_outputs(1799));
    outputs(5035) <= not(layer0_outputs(6475)) or (layer0_outputs(7421));
    outputs(5036) <= layer0_outputs(1773);
    outputs(5037) <= (layer0_outputs(3090)) and not (layer0_outputs(1377));
    outputs(5038) <= layer0_outputs(6006);
    outputs(5039) <= not(layer0_outputs(4449)) or (layer0_outputs(1211));
    outputs(5040) <= (layer0_outputs(7553)) and not (layer0_outputs(3120));
    outputs(5041) <= not(layer0_outputs(2167));
    outputs(5042) <= (layer0_outputs(829)) xor (layer0_outputs(1733));
    outputs(5043) <= not(layer0_outputs(707)) or (layer0_outputs(4530));
    outputs(5044) <= layer0_outputs(1330);
    outputs(5045) <= not(layer0_outputs(4918)) or (layer0_outputs(4377));
    outputs(5046) <= not(layer0_outputs(2725));
    outputs(5047) <= not(layer0_outputs(3227));
    outputs(5048) <= not(layer0_outputs(2991));
    outputs(5049) <= not((layer0_outputs(6583)) or (layer0_outputs(1989)));
    outputs(5050) <= not((layer0_outputs(877)) or (layer0_outputs(644)));
    outputs(5051) <= layer0_outputs(6231);
    outputs(5052) <= (layer0_outputs(4025)) and not (layer0_outputs(159));
    outputs(5053) <= layer0_outputs(3760);
    outputs(5054) <= not(layer0_outputs(387));
    outputs(5055) <= (layer0_outputs(4193)) xor (layer0_outputs(2076));
    outputs(5056) <= (layer0_outputs(3388)) and not (layer0_outputs(1876));
    outputs(5057) <= (layer0_outputs(4650)) or (layer0_outputs(915));
    outputs(5058) <= not(layer0_outputs(4277));
    outputs(5059) <= layer0_outputs(532);
    outputs(5060) <= layer0_outputs(4402);
    outputs(5061) <= (layer0_outputs(1536)) xor (layer0_outputs(5406));
    outputs(5062) <= not(layer0_outputs(7143));
    outputs(5063) <= layer0_outputs(1417);
    outputs(5064) <= not(layer0_outputs(4934));
    outputs(5065) <= (layer0_outputs(3797)) and (layer0_outputs(1352));
    outputs(5066) <= (layer0_outputs(6692)) and not (layer0_outputs(5594));
    outputs(5067) <= not(layer0_outputs(2536));
    outputs(5068) <= not(layer0_outputs(3519));
    outputs(5069) <= (layer0_outputs(5470)) and not (layer0_outputs(4975));
    outputs(5070) <= layer0_outputs(6462);
    outputs(5071) <= layer0_outputs(3006);
    outputs(5072) <= (layer0_outputs(7033)) and not (layer0_outputs(7037));
    outputs(5073) <= layer0_outputs(310);
    outputs(5074) <= not(layer0_outputs(6640));
    outputs(5075) <= not(layer0_outputs(5717));
    outputs(5076) <= (layer0_outputs(2349)) xor (layer0_outputs(1595));
    outputs(5077) <= not(layer0_outputs(4351));
    outputs(5078) <= layer0_outputs(1305);
    outputs(5079) <= not(layer0_outputs(5821)) or (layer0_outputs(7453));
    outputs(5080) <= (layer0_outputs(7424)) xor (layer0_outputs(1903));
    outputs(5081) <= layer0_outputs(143);
    outputs(5082) <= not(layer0_outputs(2084));
    outputs(5083) <= not(layer0_outputs(3119));
    outputs(5084) <= layer0_outputs(232);
    outputs(5085) <= layer0_outputs(593);
    outputs(5086) <= layer0_outputs(172);
    outputs(5087) <= (layer0_outputs(7428)) xor (layer0_outputs(4815));
    outputs(5088) <= not(layer0_outputs(904));
    outputs(5089) <= not(layer0_outputs(5521)) or (layer0_outputs(6464));
    outputs(5090) <= not((layer0_outputs(1679)) xor (layer0_outputs(4579)));
    outputs(5091) <= not(layer0_outputs(864));
    outputs(5092) <= not(layer0_outputs(5891)) or (layer0_outputs(842));
    outputs(5093) <= (layer0_outputs(5389)) and (layer0_outputs(6231));
    outputs(5094) <= not(layer0_outputs(456));
    outputs(5095) <= not(layer0_outputs(3779));
    outputs(5096) <= (layer0_outputs(7559)) xor (layer0_outputs(4298));
    outputs(5097) <= not(layer0_outputs(6503));
    outputs(5098) <= (layer0_outputs(897)) and not (layer0_outputs(2202));
    outputs(5099) <= not((layer0_outputs(972)) xor (layer0_outputs(5691)));
    outputs(5100) <= (layer0_outputs(2227)) xor (layer0_outputs(95));
    outputs(5101) <= not((layer0_outputs(6985)) or (layer0_outputs(4872)));
    outputs(5102) <= layer0_outputs(3694);
    outputs(5103) <= (layer0_outputs(1154)) xor (layer0_outputs(5833));
    outputs(5104) <= not(layer0_outputs(7223));
    outputs(5105) <= layer0_outputs(4860);
    outputs(5106) <= not(layer0_outputs(5377)) or (layer0_outputs(4933));
    outputs(5107) <= layer0_outputs(4569);
    outputs(5108) <= layer0_outputs(5305);
    outputs(5109) <= not(layer0_outputs(783)) or (layer0_outputs(6963));
    outputs(5110) <= (layer0_outputs(1579)) xor (layer0_outputs(3078));
    outputs(5111) <= not(layer0_outputs(1227));
    outputs(5112) <= not(layer0_outputs(6784));
    outputs(5113) <= not(layer0_outputs(2299)) or (layer0_outputs(2670));
    outputs(5114) <= (layer0_outputs(279)) and not (layer0_outputs(5838));
    outputs(5115) <= layer0_outputs(6259);
    outputs(5116) <= (layer0_outputs(5310)) xor (layer0_outputs(1246));
    outputs(5117) <= layer0_outputs(7466);
    outputs(5118) <= (layer0_outputs(2666)) and not (layer0_outputs(5253));
    outputs(5119) <= not(layer0_outputs(6892));
    outputs(5120) <= layer0_outputs(5560);
    outputs(5121) <= (layer0_outputs(1977)) and not (layer0_outputs(3772));
    outputs(5122) <= layer0_outputs(4776);
    outputs(5123) <= not(layer0_outputs(3560)) or (layer0_outputs(7323));
    outputs(5124) <= not(layer0_outputs(5602));
    outputs(5125) <= not(layer0_outputs(956));
    outputs(5126) <= (layer0_outputs(4426)) and not (layer0_outputs(6643));
    outputs(5127) <= not(layer0_outputs(3579));
    outputs(5128) <= not((layer0_outputs(6972)) xor (layer0_outputs(2342)));
    outputs(5129) <= not(layer0_outputs(281));
    outputs(5130) <= layer0_outputs(5026);
    outputs(5131) <= (layer0_outputs(6865)) and (layer0_outputs(6320));
    outputs(5132) <= not((layer0_outputs(2780)) xor (layer0_outputs(4007)));
    outputs(5133) <= not((layer0_outputs(113)) or (layer0_outputs(2747)));
    outputs(5134) <= (layer0_outputs(4150)) and not (layer0_outputs(5487));
    outputs(5135) <= (layer0_outputs(5514)) and not (layer0_outputs(2442));
    outputs(5136) <= (layer0_outputs(1434)) and (layer0_outputs(6751));
    outputs(5137) <= not(layer0_outputs(92)) or (layer0_outputs(887));
    outputs(5138) <= not(layer0_outputs(7045)) or (layer0_outputs(2330));
    outputs(5139) <= (layer0_outputs(6272)) xor (layer0_outputs(4305));
    outputs(5140) <= not(layer0_outputs(4866));
    outputs(5141) <= not(layer0_outputs(3537));
    outputs(5142) <= not((layer0_outputs(3991)) xor (layer0_outputs(6734)));
    outputs(5143) <= layer0_outputs(2776);
    outputs(5144) <= (layer0_outputs(478)) xor (layer0_outputs(4645));
    outputs(5145) <= layer0_outputs(3526);
    outputs(5146) <= not(layer0_outputs(2917));
    outputs(5147) <= not((layer0_outputs(3254)) or (layer0_outputs(3165)));
    outputs(5148) <= (layer0_outputs(7061)) xor (layer0_outputs(5384));
    outputs(5149) <= not(layer0_outputs(3192));
    outputs(5150) <= not(layer0_outputs(7376));
    outputs(5151) <= layer0_outputs(6870);
    outputs(5152) <= (layer0_outputs(247)) and not (layer0_outputs(6349));
    outputs(5153) <= (layer0_outputs(5621)) and (layer0_outputs(4362));
    outputs(5154) <= not((layer0_outputs(2729)) xor (layer0_outputs(1305)));
    outputs(5155) <= layer0_outputs(965);
    outputs(5156) <= (layer0_outputs(647)) xor (layer0_outputs(1618));
    outputs(5157) <= not((layer0_outputs(2870)) xor (layer0_outputs(3592)));
    outputs(5158) <= not((layer0_outputs(4957)) xor (layer0_outputs(1920)));
    outputs(5159) <= not(layer0_outputs(225));
    outputs(5160) <= layer0_outputs(3876);
    outputs(5161) <= layer0_outputs(7075);
    outputs(5162) <= not((layer0_outputs(90)) xor (layer0_outputs(5508)));
    outputs(5163) <= (layer0_outputs(4079)) and not (layer0_outputs(2800));
    outputs(5164) <= not((layer0_outputs(6938)) xor (layer0_outputs(3657)));
    outputs(5165) <= not(layer0_outputs(691)) or (layer0_outputs(5438));
    outputs(5166) <= not(layer0_outputs(7257)) or (layer0_outputs(2522));
    outputs(5167) <= (layer0_outputs(6008)) and not (layer0_outputs(574));
    outputs(5168) <= not(layer0_outputs(3915)) or (layer0_outputs(7641));
    outputs(5169) <= layer0_outputs(5211);
    outputs(5170) <= not((layer0_outputs(995)) xor (layer0_outputs(1725)));
    outputs(5171) <= (layer0_outputs(89)) and not (layer0_outputs(1643));
    outputs(5172) <= not((layer0_outputs(4689)) and (layer0_outputs(4635)));
    outputs(5173) <= not(layer0_outputs(2490)) or (layer0_outputs(4260));
    outputs(5174) <= (layer0_outputs(932)) and not (layer0_outputs(814));
    outputs(5175) <= layer0_outputs(5347);
    outputs(5176) <= layer0_outputs(319);
    outputs(5177) <= not((layer0_outputs(7206)) or (layer0_outputs(863)));
    outputs(5178) <= (layer0_outputs(2256)) and not (layer0_outputs(926));
    outputs(5179) <= not(layer0_outputs(529));
    outputs(5180) <= not((layer0_outputs(3267)) and (layer0_outputs(7600)));
    outputs(5181) <= not((layer0_outputs(3008)) xor (layer0_outputs(2493)));
    outputs(5182) <= not((layer0_outputs(7247)) xor (layer0_outputs(719)));
    outputs(5183) <= (layer0_outputs(6588)) and not (layer0_outputs(7506));
    outputs(5184) <= not(layer0_outputs(3586));
    outputs(5185) <= (layer0_outputs(3652)) and not (layer0_outputs(6794));
    outputs(5186) <= not(layer0_outputs(2037));
    outputs(5187) <= not((layer0_outputs(7533)) or (layer0_outputs(5983)));
    outputs(5188) <= not(layer0_outputs(5260));
    outputs(5189) <= (layer0_outputs(5862)) and not (layer0_outputs(2365));
    outputs(5190) <= not((layer0_outputs(5602)) or (layer0_outputs(1072)));
    outputs(5191) <= (layer0_outputs(1354)) xor (layer0_outputs(3656));
    outputs(5192) <= (layer0_outputs(4180)) or (layer0_outputs(817));
    outputs(5193) <= not((layer0_outputs(7427)) or (layer0_outputs(4001)));
    outputs(5194) <= layer0_outputs(4503);
    outputs(5195) <= layer0_outputs(1711);
    outputs(5196) <= (layer0_outputs(7524)) and not (layer0_outputs(5375));
    outputs(5197) <= not(layer0_outputs(3959));
    outputs(5198) <= (layer0_outputs(3915)) xor (layer0_outputs(1201));
    outputs(5199) <= (layer0_outputs(2045)) xor (layer0_outputs(5127));
    outputs(5200) <= (layer0_outputs(7226)) and not (layer0_outputs(1377));
    outputs(5201) <= (layer0_outputs(2993)) xor (layer0_outputs(6553));
    outputs(5202) <= not((layer0_outputs(5028)) xor (layer0_outputs(566)));
    outputs(5203) <= not(layer0_outputs(49));
    outputs(5204) <= (layer0_outputs(1867)) and not (layer0_outputs(4774));
    outputs(5205) <= not((layer0_outputs(5318)) and (layer0_outputs(892)));
    outputs(5206) <= (layer0_outputs(1828)) and (layer0_outputs(5988));
    outputs(5207) <= not(layer0_outputs(3476)) or (layer0_outputs(6476));
    outputs(5208) <= (layer0_outputs(2519)) and not (layer0_outputs(4842));
    outputs(5209) <= layer0_outputs(2309);
    outputs(5210) <= not(layer0_outputs(177));
    outputs(5211) <= not((layer0_outputs(4826)) or (layer0_outputs(5585)));
    outputs(5212) <= not(layer0_outputs(3238)) or (layer0_outputs(6684));
    outputs(5213) <= not((layer0_outputs(2456)) or (layer0_outputs(6783)));
    outputs(5214) <= layer0_outputs(737);
    outputs(5215) <= layer0_outputs(2533);
    outputs(5216) <= not((layer0_outputs(7093)) xor (layer0_outputs(7598)));
    outputs(5217) <= layer0_outputs(3716);
    outputs(5218) <= not(layer0_outputs(4546));
    outputs(5219) <= (layer0_outputs(3730)) and not (layer0_outputs(4849));
    outputs(5220) <= (layer0_outputs(173)) xor (layer0_outputs(7284));
    outputs(5221) <= not(layer0_outputs(3222));
    outputs(5222) <= not(layer0_outputs(1360));
    outputs(5223) <= (layer0_outputs(941)) and not (layer0_outputs(5521));
    outputs(5224) <= not((layer0_outputs(5213)) xor (layer0_outputs(789)));
    outputs(5225) <= (layer0_outputs(7249)) xor (layer0_outputs(4086));
    outputs(5226) <= not(layer0_outputs(1914));
    outputs(5227) <= not(layer0_outputs(7217)) or (layer0_outputs(3590));
    outputs(5228) <= not(layer0_outputs(4189));
    outputs(5229) <= not(layer0_outputs(979));
    outputs(5230) <= (layer0_outputs(6939)) xor (layer0_outputs(7029));
    outputs(5231) <= not((layer0_outputs(4930)) xor (layer0_outputs(2593)));
    outputs(5232) <= layer0_outputs(881);
    outputs(5233) <= layer0_outputs(3741);
    outputs(5234) <= (layer0_outputs(3076)) and (layer0_outputs(1580));
    outputs(5235) <= (layer0_outputs(4407)) xor (layer0_outputs(7442));
    outputs(5236) <= not(layer0_outputs(1026));
    outputs(5237) <= layer0_outputs(5576);
    outputs(5238) <= not(layer0_outputs(475));
    outputs(5239) <= not(layer0_outputs(566)) or (layer0_outputs(2870));
    outputs(5240) <= (layer0_outputs(1152)) and not (layer0_outputs(1838));
    outputs(5241) <= not((layer0_outputs(2380)) xor (layer0_outputs(1633)));
    outputs(5242) <= layer0_outputs(6374);
    outputs(5243) <= not(layer0_outputs(1897));
    outputs(5244) <= layer0_outputs(4174);
    outputs(5245) <= layer0_outputs(3054);
    outputs(5246) <= (layer0_outputs(1050)) xor (layer0_outputs(594));
    outputs(5247) <= not(layer0_outputs(4473));
    outputs(5248) <= not(layer0_outputs(3301));
    outputs(5249) <= (layer0_outputs(818)) and not (layer0_outputs(5780));
    outputs(5250) <= not((layer0_outputs(2095)) xor (layer0_outputs(5973)));
    outputs(5251) <= layer0_outputs(6912);
    outputs(5252) <= layer0_outputs(4809);
    outputs(5253) <= not(layer0_outputs(5644)) or (layer0_outputs(6167));
    outputs(5254) <= not(layer0_outputs(6082));
    outputs(5255) <= layer0_outputs(201);
    outputs(5256) <= (layer0_outputs(3055)) and not (layer0_outputs(2189));
    outputs(5257) <= (layer0_outputs(3453)) and not (layer0_outputs(6284));
    outputs(5258) <= not(layer0_outputs(2545));
    outputs(5259) <= (layer0_outputs(3690)) and (layer0_outputs(207));
    outputs(5260) <= not(layer0_outputs(5631)) or (layer0_outputs(2397));
    outputs(5261) <= (layer0_outputs(3974)) xor (layer0_outputs(1790));
    outputs(5262) <= (layer0_outputs(4679)) or (layer0_outputs(1493));
    outputs(5263) <= (layer0_outputs(6143)) xor (layer0_outputs(4852));
    outputs(5264) <= not(layer0_outputs(7416));
    outputs(5265) <= not(layer0_outputs(4984));
    outputs(5266) <= (layer0_outputs(1407)) xor (layer0_outputs(6322));
    outputs(5267) <= (layer0_outputs(5331)) or (layer0_outputs(301));
    outputs(5268) <= (layer0_outputs(4454)) and not (layer0_outputs(1791));
    outputs(5269) <= not((layer0_outputs(1804)) xor (layer0_outputs(2553)));
    outputs(5270) <= (layer0_outputs(1335)) and not (layer0_outputs(5897));
    outputs(5271) <= not(layer0_outputs(2402));
    outputs(5272) <= not((layer0_outputs(2769)) xor (layer0_outputs(4551)));
    outputs(5273) <= layer0_outputs(7588);
    outputs(5274) <= (layer0_outputs(7509)) and (layer0_outputs(6767));
    outputs(5275) <= layer0_outputs(6965);
    outputs(5276) <= not((layer0_outputs(5709)) xor (layer0_outputs(5649)));
    outputs(5277) <= layer0_outputs(806);
    outputs(5278) <= layer0_outputs(997);
    outputs(5279) <= layer0_outputs(1455);
    outputs(5280) <= layer0_outputs(2705);
    outputs(5281) <= layer0_outputs(975);
    outputs(5282) <= (layer0_outputs(3878)) and not (layer0_outputs(6554));
    outputs(5283) <= not((layer0_outputs(4579)) and (layer0_outputs(4626)));
    outputs(5284) <= not((layer0_outputs(374)) and (layer0_outputs(6091)));
    outputs(5285) <= (layer0_outputs(4786)) xor (layer0_outputs(1698));
    outputs(5286) <= not((layer0_outputs(5581)) xor (layer0_outputs(6113)));
    outputs(5287) <= not((layer0_outputs(1676)) or (layer0_outputs(4563)));
    outputs(5288) <= not(layer0_outputs(6933));
    outputs(5289) <= not(layer0_outputs(6299));
    outputs(5290) <= (layer0_outputs(4757)) and not (layer0_outputs(5171));
    outputs(5291) <= not(layer0_outputs(4391)) or (layer0_outputs(4091));
    outputs(5292) <= not(layer0_outputs(6725));
    outputs(5293) <= layer0_outputs(4889);
    outputs(5294) <= layer0_outputs(2103);
    outputs(5295) <= not(layer0_outputs(5159));
    outputs(5296) <= not(layer0_outputs(3840));
    outputs(5297) <= not((layer0_outputs(2173)) xor (layer0_outputs(3919)));
    outputs(5298) <= layer0_outputs(6122);
    outputs(5299) <= (layer0_outputs(7274)) xor (layer0_outputs(3522));
    outputs(5300) <= not((layer0_outputs(2846)) and (layer0_outputs(6564)));
    outputs(5301) <= (layer0_outputs(2818)) xor (layer0_outputs(3900));
    outputs(5302) <= layer0_outputs(4942);
    outputs(5303) <= layer0_outputs(1729);
    outputs(5304) <= not((layer0_outputs(5864)) or (layer0_outputs(1879)));
    outputs(5305) <= (layer0_outputs(5689)) and not (layer0_outputs(2863));
    outputs(5306) <= layer0_outputs(1478);
    outputs(5307) <= not((layer0_outputs(4485)) xor (layer0_outputs(5164)));
    outputs(5308) <= layer0_outputs(3830);
    outputs(5309) <= not(layer0_outputs(5181));
    outputs(5310) <= not(layer0_outputs(2372)) or (layer0_outputs(7423));
    outputs(5311) <= layer0_outputs(7536);
    outputs(5312) <= layer0_outputs(7644);
    outputs(5313) <= (layer0_outputs(4561)) and (layer0_outputs(7392));
    outputs(5314) <= not(layer0_outputs(3446));
    outputs(5315) <= (layer0_outputs(4532)) xor (layer0_outputs(2322));
    outputs(5316) <= not(layer0_outputs(1638));
    outputs(5317) <= layer0_outputs(1214);
    outputs(5318) <= (layer0_outputs(3970)) xor (layer0_outputs(7027));
    outputs(5319) <= layer0_outputs(7186);
    outputs(5320) <= layer0_outputs(5843);
    outputs(5321) <= not((layer0_outputs(3248)) or (layer0_outputs(5367)));
    outputs(5322) <= (layer0_outputs(4326)) xor (layer0_outputs(1194));
    outputs(5323) <= layer0_outputs(5532);
    outputs(5324) <= not(layer0_outputs(4164));
    outputs(5325) <= (layer0_outputs(2517)) xor (layer0_outputs(915));
    outputs(5326) <= not(layer0_outputs(1658));
    outputs(5327) <= (layer0_outputs(2490)) xor (layer0_outputs(368));
    outputs(5328) <= not(layer0_outputs(7396));
    outputs(5329) <= (layer0_outputs(5228)) xor (layer0_outputs(4447));
    outputs(5330) <= not(layer0_outputs(332));
    outputs(5331) <= not((layer0_outputs(7370)) or (layer0_outputs(2753)));
    outputs(5332) <= not((layer0_outputs(1719)) and (layer0_outputs(412)));
    outputs(5333) <= (layer0_outputs(2688)) and not (layer0_outputs(6940));
    outputs(5334) <= not(layer0_outputs(6422));
    outputs(5335) <= layer0_outputs(5681);
    outputs(5336) <= (layer0_outputs(4504)) xor (layer0_outputs(985));
    outputs(5337) <= (layer0_outputs(6980)) xor (layer0_outputs(1148));
    outputs(5338) <= layer0_outputs(5825);
    outputs(5339) <= not(layer0_outputs(4668)) or (layer0_outputs(843));
    outputs(5340) <= not(layer0_outputs(974));
    outputs(5341) <= not((layer0_outputs(6645)) or (layer0_outputs(3233)));
    outputs(5342) <= not(layer0_outputs(4695)) or (layer0_outputs(6728));
    outputs(5343) <= not(layer0_outputs(2964));
    outputs(5344) <= (layer0_outputs(5888)) and not (layer0_outputs(2016));
    outputs(5345) <= not((layer0_outputs(6066)) or (layer0_outputs(208)));
    outputs(5346) <= not(layer0_outputs(30));
    outputs(5347) <= (layer0_outputs(2618)) xor (layer0_outputs(6198));
    outputs(5348) <= (layer0_outputs(2985)) and not (layer0_outputs(519));
    outputs(5349) <= (layer0_outputs(4535)) and not (layer0_outputs(5101));
    outputs(5350) <= not(layer0_outputs(7542)) or (layer0_outputs(684));
    outputs(5351) <= (layer0_outputs(1783)) and (layer0_outputs(3050));
    outputs(5352) <= not((layer0_outputs(1501)) xor (layer0_outputs(2070)));
    outputs(5353) <= layer0_outputs(7526);
    outputs(5354) <= not(layer0_outputs(2411));
    outputs(5355) <= not(layer0_outputs(7040));
    outputs(5356) <= (layer0_outputs(1902)) and not (layer0_outputs(4190));
    outputs(5357) <= (layer0_outputs(5359)) and (layer0_outputs(5782));
    outputs(5358) <= (layer0_outputs(715)) xor (layer0_outputs(4008));
    outputs(5359) <= not(layer0_outputs(4225));
    outputs(5360) <= not(layer0_outputs(4891));
    outputs(5361) <= (layer0_outputs(2145)) xor (layer0_outputs(5928));
    outputs(5362) <= layer0_outputs(4170);
    outputs(5363) <= (layer0_outputs(3399)) and (layer0_outputs(1711));
    outputs(5364) <= not((layer0_outputs(3636)) and (layer0_outputs(3362)));
    outputs(5365) <= not((layer0_outputs(2732)) or (layer0_outputs(4833)));
    outputs(5366) <= layer0_outputs(2450);
    outputs(5367) <= not((layer0_outputs(7189)) xor (layer0_outputs(6594)));
    outputs(5368) <= layer0_outputs(7424);
    outputs(5369) <= layer0_outputs(5335);
    outputs(5370) <= not(layer0_outputs(645));
    outputs(5371) <= (layer0_outputs(3009)) and not (layer0_outputs(1917));
    outputs(5372) <= (layer0_outputs(5337)) and not (layer0_outputs(5085));
    outputs(5373) <= not(layer0_outputs(5549));
    outputs(5374) <= (layer0_outputs(641)) and not (layer0_outputs(5884));
    outputs(5375) <= layer0_outputs(1548);
    outputs(5376) <= (layer0_outputs(3487)) or (layer0_outputs(1129));
    outputs(5377) <= not((layer0_outputs(5096)) xor (layer0_outputs(495)));
    outputs(5378) <= (layer0_outputs(6605)) xor (layer0_outputs(4144));
    outputs(5379) <= (layer0_outputs(600)) and not (layer0_outputs(5603));
    outputs(5380) <= not(layer0_outputs(444));
    outputs(5381) <= (layer0_outputs(4966)) and (layer0_outputs(4859));
    outputs(5382) <= (layer0_outputs(6363)) xor (layer0_outputs(3217));
    outputs(5383) <= not(layer0_outputs(1234));
    outputs(5384) <= (layer0_outputs(6262)) xor (layer0_outputs(36));
    outputs(5385) <= not((layer0_outputs(1068)) xor (layer0_outputs(4774)));
    outputs(5386) <= not(layer0_outputs(827));
    outputs(5387) <= (layer0_outputs(49)) and (layer0_outputs(213));
    outputs(5388) <= layer0_outputs(3249);
    outputs(5389) <= not(layer0_outputs(4600));
    outputs(5390) <= not((layer0_outputs(3746)) xor (layer0_outputs(3571)));
    outputs(5391) <= (layer0_outputs(7457)) xor (layer0_outputs(4876));
    outputs(5392) <= (layer0_outputs(2918)) and (layer0_outputs(1550));
    outputs(5393) <= (layer0_outputs(2828)) xor (layer0_outputs(1431));
    outputs(5394) <= (layer0_outputs(6040)) and not (layer0_outputs(7473));
    outputs(5395) <= layer0_outputs(3811);
    outputs(5396) <= (layer0_outputs(5196)) and not (layer0_outputs(2945));
    outputs(5397) <= (layer0_outputs(2673)) and not (layer0_outputs(2632));
    outputs(5398) <= not((layer0_outputs(4572)) or (layer0_outputs(7664)));
    outputs(5399) <= (layer0_outputs(1676)) and not (layer0_outputs(5618));
    outputs(5400) <= not(layer0_outputs(10)) or (layer0_outputs(3383));
    outputs(5401) <= not(layer0_outputs(6021));
    outputs(5402) <= (layer0_outputs(4319)) and (layer0_outputs(2358));
    outputs(5403) <= not(layer0_outputs(6148));
    outputs(5404) <= layer0_outputs(3834);
    outputs(5405) <= (layer0_outputs(432)) and not (layer0_outputs(4902));
    outputs(5406) <= not(layer0_outputs(4310));
    outputs(5407) <= not((layer0_outputs(1986)) xor (layer0_outputs(3264)));
    outputs(5408) <= (layer0_outputs(4805)) and not (layer0_outputs(1142));
    outputs(5409) <= not(layer0_outputs(4227));
    outputs(5410) <= not(layer0_outputs(1684));
    outputs(5411) <= layer0_outputs(2006);
    outputs(5412) <= (layer0_outputs(7332)) and not (layer0_outputs(1470));
    outputs(5413) <= layer0_outputs(847);
    outputs(5414) <= (layer0_outputs(3828)) xor (layer0_outputs(4417));
    outputs(5415) <= not(layer0_outputs(4903));
    outputs(5416) <= (layer0_outputs(2375)) and not (layer0_outputs(2595));
    outputs(5417) <= (layer0_outputs(3277)) and (layer0_outputs(244));
    outputs(5418) <= (layer0_outputs(2193)) and not (layer0_outputs(1770));
    outputs(5419) <= layer0_outputs(1563);
    outputs(5420) <= not((layer0_outputs(6101)) xor (layer0_outputs(6937)));
    outputs(5421) <= not(layer0_outputs(1008));
    outputs(5422) <= (layer0_outputs(3188)) and (layer0_outputs(7450));
    outputs(5423) <= not((layer0_outputs(2069)) or (layer0_outputs(3759)));
    outputs(5424) <= '0';
    outputs(5425) <= layer0_outputs(3588);
    outputs(5426) <= not(layer0_outputs(5653)) or (layer0_outputs(158));
    outputs(5427) <= not((layer0_outputs(589)) xor (layer0_outputs(4273)));
    outputs(5428) <= not(layer0_outputs(4994));
    outputs(5429) <= not((layer0_outputs(4204)) or (layer0_outputs(223)));
    outputs(5430) <= (layer0_outputs(1584)) and not (layer0_outputs(7618));
    outputs(5431) <= not((layer0_outputs(614)) xor (layer0_outputs(582)));
    outputs(5432) <= layer0_outputs(6910);
    outputs(5433) <= (layer0_outputs(2774)) xor (layer0_outputs(5371));
    outputs(5434) <= not((layer0_outputs(707)) xor (layer0_outputs(6857)));
    outputs(5435) <= not((layer0_outputs(4540)) or (layer0_outputs(2331)));
    outputs(5436) <= layer0_outputs(7051);
    outputs(5437) <= not(layer0_outputs(4342));
    outputs(5438) <= layer0_outputs(4292);
    outputs(5439) <= not(layer0_outputs(3740));
    outputs(5440) <= (layer0_outputs(5309)) or (layer0_outputs(3012));
    outputs(5441) <= layer0_outputs(7569);
    outputs(5442) <= not(layer0_outputs(659));
    outputs(5443) <= not(layer0_outputs(7134));
    outputs(5444) <= (layer0_outputs(3768)) xor (layer0_outputs(3651));
    outputs(5445) <= not(layer0_outputs(4597));
    outputs(5446) <= not(layer0_outputs(4987));
    outputs(5447) <= not(layer0_outputs(2730));
    outputs(5448) <= (layer0_outputs(4624)) xor (layer0_outputs(4262));
    outputs(5449) <= layer0_outputs(5685);
    outputs(5450) <= (layer0_outputs(2229)) xor (layer0_outputs(2004));
    outputs(5451) <= (layer0_outputs(480)) and (layer0_outputs(7288));
    outputs(5452) <= layer0_outputs(3939);
    outputs(5453) <= layer0_outputs(7133);
    outputs(5454) <= layer0_outputs(2620);
    outputs(5455) <= not(layer0_outputs(4103));
    outputs(5456) <= not((layer0_outputs(5162)) xor (layer0_outputs(1267)));
    outputs(5457) <= not(layer0_outputs(5888));
    outputs(5458) <= not(layer0_outputs(4300));
    outputs(5459) <= (layer0_outputs(938)) and not (layer0_outputs(3382));
    outputs(5460) <= (layer0_outputs(5447)) and not (layer0_outputs(3277));
    outputs(5461) <= not(layer0_outputs(6800));
    outputs(5462) <= not(layer0_outputs(6771));
    outputs(5463) <= layer0_outputs(2655);
    outputs(5464) <= layer0_outputs(914);
    outputs(5465) <= (layer0_outputs(7200)) and not (layer0_outputs(1736));
    outputs(5466) <= not((layer0_outputs(4557)) xor (layer0_outputs(1630)));
    outputs(5467) <= not((layer0_outputs(2989)) or (layer0_outputs(2308)));
    outputs(5468) <= not((layer0_outputs(4161)) xor (layer0_outputs(3235)));
    outputs(5469) <= not(layer0_outputs(5750));
    outputs(5470) <= (layer0_outputs(2598)) and not (layer0_outputs(2970));
    outputs(5471) <= (layer0_outputs(6546)) and not (layer0_outputs(349));
    outputs(5472) <= (layer0_outputs(5692)) and (layer0_outputs(6003));
    outputs(5473) <= layer0_outputs(2633);
    outputs(5474) <= (layer0_outputs(6945)) and (layer0_outputs(4931));
    outputs(5475) <= (layer0_outputs(7546)) and (layer0_outputs(1293));
    outputs(5476) <= layer0_outputs(4869);
    outputs(5477) <= (layer0_outputs(6825)) and (layer0_outputs(3071));
    outputs(5478) <= not(layer0_outputs(6148));
    outputs(5479) <= layer0_outputs(3580);
    outputs(5480) <= layer0_outputs(6710);
    outputs(5481) <= layer0_outputs(3957);
    outputs(5482) <= (layer0_outputs(6470)) and not (layer0_outputs(5189));
    outputs(5483) <= not(layer0_outputs(2498));
    outputs(5484) <= not(layer0_outputs(4573));
    outputs(5485) <= (layer0_outputs(1675)) and not (layer0_outputs(6103));
    outputs(5486) <= (layer0_outputs(4339)) and (layer0_outputs(7449));
    outputs(5487) <= not((layer0_outputs(3879)) or (layer0_outputs(3346)));
    outputs(5488) <= (layer0_outputs(6518)) and not (layer0_outputs(2865));
    outputs(5489) <= layer0_outputs(5960);
    outputs(5490) <= not((layer0_outputs(6041)) or (layer0_outputs(1468)));
    outputs(5491) <= not((layer0_outputs(7527)) or (layer0_outputs(184)));
    outputs(5492) <= layer0_outputs(5063);
    outputs(5493) <= not((layer0_outputs(6053)) and (layer0_outputs(1287)));
    outputs(5494) <= layer0_outputs(156);
    outputs(5495) <= not((layer0_outputs(5433)) and (layer0_outputs(5590)));
    outputs(5496) <= (layer0_outputs(6667)) and not (layer0_outputs(5001));
    outputs(5497) <= '0';
    outputs(5498) <= (layer0_outputs(4736)) xor (layer0_outputs(6838));
    outputs(5499) <= not((layer0_outputs(1294)) xor (layer0_outputs(2962)));
    outputs(5500) <= (layer0_outputs(320)) or (layer0_outputs(2846));
    outputs(5501) <= (layer0_outputs(6208)) xor (layer0_outputs(3204));
    outputs(5502) <= (layer0_outputs(1249)) xor (layer0_outputs(4040));
    outputs(5503) <= '0';
    outputs(5504) <= not(layer0_outputs(127));
    outputs(5505) <= layer0_outputs(1809);
    outputs(5506) <= (layer0_outputs(1437)) and (layer0_outputs(1137));
    outputs(5507) <= not(layer0_outputs(4342));
    outputs(5508) <= not((layer0_outputs(2371)) xor (layer0_outputs(1438)));
    outputs(5509) <= layer0_outputs(1321);
    outputs(5510) <= (layer0_outputs(5929)) and not (layer0_outputs(4222));
    outputs(5511) <= layer0_outputs(2593);
    outputs(5512) <= layer0_outputs(2766);
    outputs(5513) <= not(layer0_outputs(5562));
    outputs(5514) <= (layer0_outputs(700)) and (layer0_outputs(5553));
    outputs(5515) <= not((layer0_outputs(5239)) and (layer0_outputs(6323)));
    outputs(5516) <= not(layer0_outputs(2695));
    outputs(5517) <= (layer0_outputs(7217)) and not (layer0_outputs(4160));
    outputs(5518) <= not((layer0_outputs(5158)) xor (layer0_outputs(3414)));
    outputs(5519) <= layer0_outputs(6254);
    outputs(5520) <= (layer0_outputs(3948)) and (layer0_outputs(4208));
    outputs(5521) <= (layer0_outputs(6096)) and not (layer0_outputs(1619));
    outputs(5522) <= not((layer0_outputs(68)) xor (layer0_outputs(3084)));
    outputs(5523) <= not(layer0_outputs(7636));
    outputs(5524) <= not((layer0_outputs(6867)) xor (layer0_outputs(6856)));
    outputs(5525) <= (layer0_outputs(3248)) and not (layer0_outputs(4580));
    outputs(5526) <= not(layer0_outputs(4384));
    outputs(5527) <= (layer0_outputs(2920)) xor (layer0_outputs(5050));
    outputs(5528) <= not(layer0_outputs(2457));
    outputs(5529) <= (layer0_outputs(6136)) and not (layer0_outputs(4752));
    outputs(5530) <= not((layer0_outputs(1857)) or (layer0_outputs(6742)));
    outputs(5531) <= (layer0_outputs(3492)) xor (layer0_outputs(5848));
    outputs(5532) <= layer0_outputs(2078);
    outputs(5533) <= not((layer0_outputs(2369)) xor (layer0_outputs(7141)));
    outputs(5534) <= not((layer0_outputs(6438)) or (layer0_outputs(1422)));
    outputs(5535) <= (layer0_outputs(3488)) and (layer0_outputs(7489));
    outputs(5536) <= layer0_outputs(112);
    outputs(5537) <= layer0_outputs(2713);
    outputs(5538) <= layer0_outputs(4493);
    outputs(5539) <= (layer0_outputs(5947)) and not (layer0_outputs(7082));
    outputs(5540) <= (layer0_outputs(2858)) xor (layer0_outputs(1800));
    outputs(5541) <= not(layer0_outputs(7344));
    outputs(5542) <= not(layer0_outputs(7169));
    outputs(5543) <= not((layer0_outputs(6941)) or (layer0_outputs(3979)));
    outputs(5544) <= layer0_outputs(4019);
    outputs(5545) <= layer0_outputs(2834);
    outputs(5546) <= (layer0_outputs(4927)) and not (layer0_outputs(4039));
    outputs(5547) <= not((layer0_outputs(2860)) xor (layer0_outputs(3172)));
    outputs(5548) <= layer0_outputs(6555);
    outputs(5549) <= not(layer0_outputs(1884));
    outputs(5550) <= layer0_outputs(3566);
    outputs(5551) <= not(layer0_outputs(6987)) or (layer0_outputs(4367));
    outputs(5552) <= (layer0_outputs(5431)) xor (layer0_outputs(1356));
    outputs(5553) <= not(layer0_outputs(7096));
    outputs(5554) <= not((layer0_outputs(246)) or (layer0_outputs(3226)));
    outputs(5555) <= (layer0_outputs(1863)) and not (layer0_outputs(7245));
    outputs(5556) <= not((layer0_outputs(2634)) or (layer0_outputs(4203)));
    outputs(5557) <= not(layer0_outputs(5741));
    outputs(5558) <= layer0_outputs(1024);
    outputs(5559) <= layer0_outputs(5635);
    outputs(5560) <= not(layer0_outputs(3227));
    outputs(5561) <= (layer0_outputs(4789)) and not (layer0_outputs(6913));
    outputs(5562) <= (layer0_outputs(2589)) and (layer0_outputs(6300));
    outputs(5563) <= '0';
    outputs(5564) <= not(layer0_outputs(325));
    outputs(5565) <= not(layer0_outputs(5297));
    outputs(5566) <= (layer0_outputs(3351)) and not (layer0_outputs(2696));
    outputs(5567) <= not(layer0_outputs(3922));
    outputs(5568) <= not((layer0_outputs(2718)) xor (layer0_outputs(465)));
    outputs(5569) <= (layer0_outputs(630)) xor (layer0_outputs(4210));
    outputs(5570) <= not((layer0_outputs(5971)) xor (layer0_outputs(4046)));
    outputs(5571) <= (layer0_outputs(506)) or (layer0_outputs(1511));
    outputs(5572) <= not((layer0_outputs(484)) xor (layer0_outputs(2298)));
    outputs(5573) <= (layer0_outputs(983)) xor (layer0_outputs(3139));
    outputs(5574) <= not(layer0_outputs(3424));
    outputs(5575) <= (layer0_outputs(1306)) and (layer0_outputs(245));
    outputs(5576) <= layer0_outputs(2391);
    outputs(5577) <= not(layer0_outputs(3934));
    outputs(5578) <= not(layer0_outputs(4324));
    outputs(5579) <= not((layer0_outputs(7638)) xor (layer0_outputs(5052)));
    outputs(5580) <= (layer0_outputs(6050)) xor (layer0_outputs(3901));
    outputs(5581) <= not((layer0_outputs(4935)) xor (layer0_outputs(2806)));
    outputs(5582) <= (layer0_outputs(2398)) and (layer0_outputs(2359));
    outputs(5583) <= layer0_outputs(1181);
    outputs(5584) <= (layer0_outputs(5734)) xor (layer0_outputs(2276));
    outputs(5585) <= layer0_outputs(1874);
    outputs(5586) <= (layer0_outputs(2914)) xor (layer0_outputs(2026));
    outputs(5587) <= (layer0_outputs(260)) and not (layer0_outputs(4424));
    outputs(5588) <= (layer0_outputs(3183)) and (layer0_outputs(331));
    outputs(5589) <= layer0_outputs(6617);
    outputs(5590) <= not(layer0_outputs(248));
    outputs(5591) <= layer0_outputs(4472);
    outputs(5592) <= not(layer0_outputs(329));
    outputs(5593) <= not(layer0_outputs(6174));
    outputs(5594) <= not((layer0_outputs(1668)) xor (layer0_outputs(5262)));
    outputs(5595) <= (layer0_outputs(4271)) or (layer0_outputs(3264));
    outputs(5596) <= not((layer0_outputs(158)) xor (layer0_outputs(4567)));
    outputs(5597) <= not(layer0_outputs(5739));
    outputs(5598) <= layer0_outputs(1734);
    outputs(5599) <= not((layer0_outputs(1592)) xor (layer0_outputs(5936)));
    outputs(5600) <= layer0_outputs(3081);
    outputs(5601) <= (layer0_outputs(1980)) and not (layer0_outputs(5180));
    outputs(5602) <= (layer0_outputs(1900)) and not (layer0_outputs(4953));
    outputs(5603) <= (layer0_outputs(4141)) or (layer0_outputs(3556));
    outputs(5604) <= (layer0_outputs(5765)) and (layer0_outputs(5194));
    outputs(5605) <= (layer0_outputs(4215)) xor (layer0_outputs(6942));
    outputs(5606) <= not((layer0_outputs(4013)) or (layer0_outputs(4974)));
    outputs(5607) <= not((layer0_outputs(2514)) xor (layer0_outputs(7116)));
    outputs(5608) <= not((layer0_outputs(98)) or (layer0_outputs(2244)));
    outputs(5609) <= not(layer0_outputs(4730));
    outputs(5610) <= layer0_outputs(2257);
    outputs(5611) <= not((layer0_outputs(5293)) xor (layer0_outputs(5913)));
    outputs(5612) <= (layer0_outputs(2719)) and (layer0_outputs(7279));
    outputs(5613) <= not((layer0_outputs(4598)) xor (layer0_outputs(7039)));
    outputs(5614) <= (layer0_outputs(533)) xor (layer0_outputs(5632));
    outputs(5615) <= layer0_outputs(3612);
    outputs(5616) <= (layer0_outputs(7441)) xor (layer0_outputs(1595));
    outputs(5617) <= layer0_outputs(192);
    outputs(5618) <= layer0_outputs(4963);
    outputs(5619) <= layer0_outputs(529);
    outputs(5620) <= (layer0_outputs(1452)) and not (layer0_outputs(1474));
    outputs(5621) <= not((layer0_outputs(5300)) xor (layer0_outputs(3809)));
    outputs(5622) <= (layer0_outputs(2969)) and not (layer0_outputs(4004));
    outputs(5623) <= layer0_outputs(4070);
    outputs(5624) <= layer0_outputs(211);
    outputs(5625) <= (layer0_outputs(2435)) or (layer0_outputs(5464));
    outputs(5626) <= layer0_outputs(2);
    outputs(5627) <= (layer0_outputs(192)) and (layer0_outputs(1251));
    outputs(5628) <= not(layer0_outputs(1603));
    outputs(5629) <= layer0_outputs(497);
    outputs(5630) <= layer0_outputs(5662);
    outputs(5631) <= layer0_outputs(3192);
    outputs(5632) <= not(layer0_outputs(444));
    outputs(5633) <= not((layer0_outputs(2180)) xor (layer0_outputs(636)));
    outputs(5634) <= not((layer0_outputs(4366)) or (layer0_outputs(5768)));
    outputs(5635) <= layer0_outputs(1091);
    outputs(5636) <= layer0_outputs(4024);
    outputs(5637) <= not(layer0_outputs(1943));
    outputs(5638) <= layer0_outputs(5209);
    outputs(5639) <= layer0_outputs(3010);
    outputs(5640) <= not(layer0_outputs(4543));
    outputs(5641) <= layer0_outputs(5172);
    outputs(5642) <= not(layer0_outputs(5655));
    outputs(5643) <= layer0_outputs(6384);
    outputs(5644) <= not(layer0_outputs(7404));
    outputs(5645) <= not((layer0_outputs(7237)) xor (layer0_outputs(6498)));
    outputs(5646) <= (layer0_outputs(5062)) xor (layer0_outputs(5985));
    outputs(5647) <= (layer0_outputs(3087)) xor (layer0_outputs(1469));
    outputs(5648) <= not((layer0_outputs(4440)) or (layer0_outputs(6775)));
    outputs(5649) <= not(layer0_outputs(6750));
    outputs(5650) <= (layer0_outputs(4371)) and (layer0_outputs(907));
    outputs(5651) <= layer0_outputs(3658);
    outputs(5652) <= (layer0_outputs(2309)) and (layer0_outputs(4231));
    outputs(5653) <= not((layer0_outputs(6652)) or (layer0_outputs(3253)));
    outputs(5654) <= not(layer0_outputs(1656));
    outputs(5655) <= (layer0_outputs(2140)) and (layer0_outputs(5658));
    outputs(5656) <= not(layer0_outputs(1189));
    outputs(5657) <= (layer0_outputs(4683)) xor (layer0_outputs(4240));
    outputs(5658) <= not((layer0_outputs(6119)) xor (layer0_outputs(6390)));
    outputs(5659) <= not(layer0_outputs(3923));
    outputs(5660) <= not((layer0_outputs(4978)) and (layer0_outputs(7418)));
    outputs(5661) <= not((layer0_outputs(6549)) and (layer0_outputs(7471)));
    outputs(5662) <= (layer0_outputs(3913)) and not (layer0_outputs(4959));
    outputs(5663) <= layer0_outputs(1487);
    outputs(5664) <= layer0_outputs(2175);
    outputs(5665) <= not(layer0_outputs(2541));
    outputs(5666) <= (layer0_outputs(7110)) and not (layer0_outputs(66));
    outputs(5667) <= not(layer0_outputs(3142));
    outputs(5668) <= not((layer0_outputs(3880)) xor (layer0_outputs(7069)));
    outputs(5669) <= layer0_outputs(3962);
    outputs(5670) <= (layer0_outputs(7374)) xor (layer0_outputs(46));
    outputs(5671) <= not(layer0_outputs(818));
    outputs(5672) <= layer0_outputs(1929);
    outputs(5673) <= (layer0_outputs(4365)) and not (layer0_outputs(2451));
    outputs(5674) <= (layer0_outputs(80)) or (layer0_outputs(5638));
    outputs(5675) <= (layer0_outputs(2258)) and (layer0_outputs(311));
    outputs(5676) <= layer0_outputs(4859);
    outputs(5677) <= not((layer0_outputs(4452)) xor (layer0_outputs(6933)));
    outputs(5678) <= (layer0_outputs(3514)) and not (layer0_outputs(1575));
    outputs(5679) <= layer0_outputs(4740);
    outputs(5680) <= layer0_outputs(2516);
    outputs(5681) <= layer0_outputs(5683);
    outputs(5682) <= not(layer0_outputs(182));
    outputs(5683) <= layer0_outputs(5209);
    outputs(5684) <= layer0_outputs(7161);
    outputs(5685) <= layer0_outputs(2680);
    outputs(5686) <= layer0_outputs(5258);
    outputs(5687) <= not(layer0_outputs(1175)) or (layer0_outputs(1131));
    outputs(5688) <= not(layer0_outputs(1998));
    outputs(5689) <= not(layer0_outputs(3183)) or (layer0_outputs(7023));
    outputs(5690) <= not((layer0_outputs(1449)) xor (layer0_outputs(3150)));
    outputs(5691) <= (layer0_outputs(5287)) and not (layer0_outputs(5818));
    outputs(5692) <= not(layer0_outputs(5041));
    outputs(5693) <= (layer0_outputs(4804)) xor (layer0_outputs(3522));
    outputs(5694) <= not((layer0_outputs(6624)) or (layer0_outputs(3594)));
    outputs(5695) <= (layer0_outputs(2701)) or (layer0_outputs(2458));
    outputs(5696) <= layer0_outputs(4822);
    outputs(5697) <= not(layer0_outputs(394)) or (layer0_outputs(6949));
    outputs(5698) <= (layer0_outputs(7395)) and (layer0_outputs(5747));
    outputs(5699) <= layer0_outputs(6176);
    outputs(5700) <= '0';
    outputs(5701) <= not((layer0_outputs(3605)) xor (layer0_outputs(7131)));
    outputs(5702) <= not((layer0_outputs(125)) xor (layer0_outputs(6484)));
    outputs(5703) <= (layer0_outputs(2907)) xor (layer0_outputs(3459));
    outputs(5704) <= (layer0_outputs(1589)) xor (layer0_outputs(2574));
    outputs(5705) <= layer0_outputs(4828);
    outputs(5706) <= layer0_outputs(2411);
    outputs(5707) <= (layer0_outputs(5654)) and not (layer0_outputs(7091));
    outputs(5708) <= (layer0_outputs(1322)) xor (layer0_outputs(2436));
    outputs(5709) <= (layer0_outputs(3423)) and not (layer0_outputs(820));
    outputs(5710) <= not(layer0_outputs(4820));
    outputs(5711) <= not((layer0_outputs(609)) or (layer0_outputs(4566)));
    outputs(5712) <= not((layer0_outputs(5469)) xor (layer0_outputs(7463)));
    outputs(5713) <= (layer0_outputs(4239)) and not (layer0_outputs(3209));
    outputs(5714) <= not(layer0_outputs(5306));
    outputs(5715) <= (layer0_outputs(2197)) and not (layer0_outputs(499));
    outputs(5716) <= (layer0_outputs(1482)) and (layer0_outputs(5442));
    outputs(5717) <= not(layer0_outputs(3293));
    outputs(5718) <= not(layer0_outputs(430)) or (layer0_outputs(1477));
    outputs(5719) <= not(layer0_outputs(2737));
    outputs(5720) <= (layer0_outputs(6625)) and not (layer0_outputs(7010));
    outputs(5721) <= not(layer0_outputs(2710));
    outputs(5722) <= (layer0_outputs(4444)) and (layer0_outputs(7581));
    outputs(5723) <= not((layer0_outputs(7597)) or (layer0_outputs(7290)));
    outputs(5724) <= layer0_outputs(6417);
    outputs(5725) <= (layer0_outputs(6325)) or (layer0_outputs(5091));
    outputs(5726) <= not((layer0_outputs(5666)) xor (layer0_outputs(631)));
    outputs(5727) <= not((layer0_outputs(6260)) xor (layer0_outputs(1573)));
    outputs(5728) <= layer0_outputs(1935);
    outputs(5729) <= layer0_outputs(3341);
    outputs(5730) <= (layer0_outputs(3802)) and not (layer0_outputs(3395));
    outputs(5731) <= not((layer0_outputs(1195)) xor (layer0_outputs(272)));
    outputs(5732) <= layer0_outputs(4857);
    outputs(5733) <= (layer0_outputs(1767)) xor (layer0_outputs(2198));
    outputs(5734) <= (layer0_outputs(1692)) and (layer0_outputs(3129));
    outputs(5735) <= not((layer0_outputs(3231)) or (layer0_outputs(2512)));
    outputs(5736) <= layer0_outputs(3477);
    outputs(5737) <= (layer0_outputs(1499)) or (layer0_outputs(6702));
    outputs(5738) <= not((layer0_outputs(2680)) and (layer0_outputs(6075)));
    outputs(5739) <= (layer0_outputs(5552)) and (layer0_outputs(458));
    outputs(5740) <= (layer0_outputs(2246)) and not (layer0_outputs(280));
    outputs(5741) <= (layer0_outputs(5704)) and not (layer0_outputs(5720));
    outputs(5742) <= not((layer0_outputs(6103)) xor (layer0_outputs(383)));
    outputs(5743) <= layer0_outputs(3696);
    outputs(5744) <= (layer0_outputs(7055)) and (layer0_outputs(1259));
    outputs(5745) <= '0';
    outputs(5746) <= not(layer0_outputs(2566));
    outputs(5747) <= (layer0_outputs(2531)) and not (layer0_outputs(855));
    outputs(5748) <= not(layer0_outputs(7256));
    outputs(5749) <= not((layer0_outputs(2940)) and (layer0_outputs(4818)));
    outputs(5750) <= (layer0_outputs(6952)) xor (layer0_outputs(619));
    outputs(5751) <= (layer0_outputs(4148)) and not (layer0_outputs(2165));
    outputs(5752) <= layer0_outputs(5581);
    outputs(5753) <= not((layer0_outputs(5437)) or (layer0_outputs(2747)));
    outputs(5754) <= (layer0_outputs(1315)) and not (layer0_outputs(5256));
    outputs(5755) <= (layer0_outputs(5449)) and not (layer0_outputs(4126));
    outputs(5756) <= not(layer0_outputs(1586));
    outputs(5757) <= (layer0_outputs(7008)) xor (layer0_outputs(3781));
    outputs(5758) <= (layer0_outputs(6912)) and not (layer0_outputs(5024));
    outputs(5759) <= layer0_outputs(4438);
    outputs(5760) <= (layer0_outputs(1919)) xor (layer0_outputs(5699));
    outputs(5761) <= layer0_outputs(1166);
    outputs(5762) <= (layer0_outputs(2381)) and not (layer0_outputs(6946));
    outputs(5763) <= layer0_outputs(2010);
    outputs(5764) <= not((layer0_outputs(7269)) xor (layer0_outputs(6908)));
    outputs(5765) <= (layer0_outputs(2837)) xor (layer0_outputs(6670));
    outputs(5766) <= (layer0_outputs(5519)) and not (layer0_outputs(4812));
    outputs(5767) <= layer0_outputs(1596);
    outputs(5768) <= (layer0_outputs(4664)) and not (layer0_outputs(3569));
    outputs(5769) <= not(layer0_outputs(7579));
    outputs(5770) <= (layer0_outputs(4733)) and not (layer0_outputs(4920));
    outputs(5771) <= not(layer0_outputs(2020));
    outputs(5772) <= not((layer0_outputs(903)) xor (layer0_outputs(271)));
    outputs(5773) <= layer0_outputs(5662);
    outputs(5774) <= not(layer0_outputs(3392));
    outputs(5775) <= not((layer0_outputs(5907)) xor (layer0_outputs(460)));
    outputs(5776) <= layer0_outputs(4353);
    outputs(5777) <= layer0_outputs(750);
    outputs(5778) <= (layer0_outputs(3733)) and (layer0_outputs(7635));
    outputs(5779) <= layer0_outputs(314);
    outputs(5780) <= layer0_outputs(751);
    outputs(5781) <= (layer0_outputs(5822)) xor (layer0_outputs(69));
    outputs(5782) <= not((layer0_outputs(4734)) or (layer0_outputs(4286)));
    outputs(5783) <= layer0_outputs(6688);
    outputs(5784) <= layer0_outputs(2579);
    outputs(5785) <= layer0_outputs(6688);
    outputs(5786) <= (layer0_outputs(6305)) xor (layer0_outputs(3082));
    outputs(5787) <= layer0_outputs(1923);
    outputs(5788) <= (layer0_outputs(323)) and (layer0_outputs(4303));
    outputs(5789) <= layer0_outputs(3083);
    outputs(5790) <= (layer0_outputs(4991)) xor (layer0_outputs(3224));
    outputs(5791) <= (layer0_outputs(2712)) and not (layer0_outputs(464));
    outputs(5792) <= not(layer0_outputs(2600));
    outputs(5793) <= not((layer0_outputs(1933)) xor (layer0_outputs(6280)));
    outputs(5794) <= not((layer0_outputs(4479)) xor (layer0_outputs(3985)));
    outputs(5795) <= layer0_outputs(2269);
    outputs(5796) <= layer0_outputs(668);
    outputs(5797) <= not(layer0_outputs(4925));
    outputs(5798) <= not(layer0_outputs(7045));
    outputs(5799) <= layer0_outputs(1125);
    outputs(5800) <= (layer0_outputs(4831)) and not (layer0_outputs(568));
    outputs(5801) <= not(layer0_outputs(3768));
    outputs(5802) <= layer0_outputs(5754);
    outputs(5803) <= (layer0_outputs(5299)) and (layer0_outputs(274));
    outputs(5804) <= layer0_outputs(3564);
    outputs(5805) <= not(layer0_outputs(6708));
    outputs(5806) <= not((layer0_outputs(6273)) or (layer0_outputs(964)));
    outputs(5807) <= layer0_outputs(109);
    outputs(5808) <= not((layer0_outputs(3973)) xor (layer0_outputs(940)));
    outputs(5809) <= not(layer0_outputs(154));
    outputs(5810) <= (layer0_outputs(123)) or (layer0_outputs(7231));
    outputs(5811) <= (layer0_outputs(4095)) xor (layer0_outputs(5896));
    outputs(5812) <= not(layer0_outputs(1059));
    outputs(5813) <= not(layer0_outputs(4427)) or (layer0_outputs(6661));
    outputs(5814) <= (layer0_outputs(1320)) xor (layer0_outputs(4181));
    outputs(5815) <= not((layer0_outputs(106)) xor (layer0_outputs(3099)));
    outputs(5816) <= not(layer0_outputs(6166)) or (layer0_outputs(2716));
    outputs(5817) <= not(layer0_outputs(1979));
    outputs(5818) <= not(layer0_outputs(2001));
    outputs(5819) <= not(layer0_outputs(6431));
    outputs(5820) <= '0';
    outputs(5821) <= (layer0_outputs(5804)) xor (layer0_outputs(6392));
    outputs(5822) <= not(layer0_outputs(7398));
    outputs(5823) <= not(layer0_outputs(33));
    outputs(5824) <= not(layer0_outputs(7485)) or (layer0_outputs(1396));
    outputs(5825) <= (layer0_outputs(3787)) and not (layer0_outputs(4749));
    outputs(5826) <= not(layer0_outputs(1841));
    outputs(5827) <= (layer0_outputs(5237)) and not (layer0_outputs(6651));
    outputs(5828) <= not(layer0_outputs(1956)) or (layer0_outputs(2537));
    outputs(5829) <= (layer0_outputs(4413)) and not (layer0_outputs(2737));
    outputs(5830) <= (layer0_outputs(3763)) and (layer0_outputs(3705));
    outputs(5831) <= layer0_outputs(187);
    outputs(5832) <= not(layer0_outputs(7537));
    outputs(5833) <= (layer0_outputs(315)) and (layer0_outputs(957));
    outputs(5834) <= not(layer0_outputs(422));
    outputs(5835) <= (layer0_outputs(455)) and not (layer0_outputs(4141));
    outputs(5836) <= (layer0_outputs(429)) and not (layer0_outputs(3369));
    outputs(5837) <= not(layer0_outputs(991)) or (layer0_outputs(7068));
    outputs(5838) <= (layer0_outputs(6903)) xor (layer0_outputs(1320));
    outputs(5839) <= layer0_outputs(3988);
    outputs(5840) <= layer0_outputs(1821);
    outputs(5841) <= layer0_outputs(2270);
    outputs(5842) <= not(layer0_outputs(5755));
    outputs(5843) <= (layer0_outputs(4760)) and not (layer0_outputs(4600));
    outputs(5844) <= (layer0_outputs(7013)) and (layer0_outputs(1843));
    outputs(5845) <= layer0_outputs(6827);
    outputs(5846) <= not(layer0_outputs(3938));
    outputs(5847) <= (layer0_outputs(2029)) and not (layer0_outputs(6820));
    outputs(5848) <= not(layer0_outputs(1134));
    outputs(5849) <= (layer0_outputs(7472)) xor (layer0_outputs(2732));
    outputs(5850) <= layer0_outputs(1691);
    outputs(5851) <= (layer0_outputs(7064)) and not (layer0_outputs(3778));
    outputs(5852) <= not(layer0_outputs(405));
    outputs(5853) <= (layer0_outputs(3252)) and not (layer0_outputs(5616));
    outputs(5854) <= layer0_outputs(3678);
    outputs(5855) <= not(layer0_outputs(2430));
    outputs(5856) <= not(layer0_outputs(1234));
    outputs(5857) <= layer0_outputs(3826);
    outputs(5858) <= (layer0_outputs(4852)) and not (layer0_outputs(5998));
    outputs(5859) <= (layer0_outputs(6181)) xor (layer0_outputs(934));
    outputs(5860) <= not(layer0_outputs(1896));
    outputs(5861) <= layer0_outputs(5621);
    outputs(5862) <= (layer0_outputs(4443)) and not (layer0_outputs(5798));
    outputs(5863) <= layer0_outputs(6928);
    outputs(5864) <= (layer0_outputs(5143)) xor (layer0_outputs(2401));
    outputs(5865) <= (layer0_outputs(2700)) xor (layer0_outputs(1808));
    outputs(5866) <= (layer0_outputs(6818)) and (layer0_outputs(1232));
    outputs(5867) <= not((layer0_outputs(5093)) and (layer0_outputs(3435)));
    outputs(5868) <= not((layer0_outputs(4995)) and (layer0_outputs(7640)));
    outputs(5869) <= (layer0_outputs(5944)) and not (layer0_outputs(1814));
    outputs(5870) <= not(layer0_outputs(2429));
    outputs(5871) <= not(layer0_outputs(6569)) or (layer0_outputs(4435));
    outputs(5872) <= not(layer0_outputs(3067));
    outputs(5873) <= not(layer0_outputs(7663));
    outputs(5874) <= (layer0_outputs(2109)) and not (layer0_outputs(5032));
    outputs(5875) <= not((layer0_outputs(5526)) or (layer0_outputs(5488)));
    outputs(5876) <= layer0_outputs(2523);
    outputs(5877) <= layer0_outputs(3328);
    outputs(5878) <= layer0_outputs(971);
    outputs(5879) <= not((layer0_outputs(6501)) xor (layer0_outputs(6726)));
    outputs(5880) <= (layer0_outputs(2936)) and not (layer0_outputs(4015));
    outputs(5881) <= not(layer0_outputs(6704));
    outputs(5882) <= layer0_outputs(1125);
    outputs(5883) <= (layer0_outputs(2671)) and not (layer0_outputs(5922));
    outputs(5884) <= (layer0_outputs(2611)) or (layer0_outputs(2796));
    outputs(5885) <= (layer0_outputs(5384)) xor (layer0_outputs(1602));
    outputs(5886) <= not(layer0_outputs(6557));
    outputs(5887) <= layer0_outputs(3189);
    outputs(5888) <= layer0_outputs(1182);
    outputs(5889) <= layer0_outputs(570);
    outputs(5890) <= layer0_outputs(6399);
    outputs(5891) <= layer0_outputs(2929);
    outputs(5892) <= layer0_outputs(1107);
    outputs(5893) <= layer0_outputs(198);
    outputs(5894) <= layer0_outputs(4888);
    outputs(5895) <= layer0_outputs(4207);
    outputs(5896) <= (layer0_outputs(7497)) and (layer0_outputs(3458));
    outputs(5897) <= layer0_outputs(958);
    outputs(5898) <= layer0_outputs(6218);
    outputs(5899) <= (layer0_outputs(4969)) xor (layer0_outputs(2698));
    outputs(5900) <= layer0_outputs(909);
    outputs(5901) <= not(layer0_outputs(5044)) or (layer0_outputs(6396));
    outputs(5902) <= not((layer0_outputs(488)) or (layer0_outputs(2372)));
    outputs(5903) <= not((layer0_outputs(2799)) or (layer0_outputs(1330)));
    outputs(5904) <= (layer0_outputs(5244)) xor (layer0_outputs(6511));
    outputs(5905) <= (layer0_outputs(5513)) and (layer0_outputs(3912));
    outputs(5906) <= not((layer0_outputs(841)) or (layer0_outputs(1693)));
    outputs(5907) <= (layer0_outputs(7224)) and not (layer0_outputs(7544));
    outputs(5908) <= not((layer0_outputs(5361)) xor (layer0_outputs(5774)));
    outputs(5909) <= layer0_outputs(289);
    outputs(5910) <= not(layer0_outputs(2033));
    outputs(5911) <= layer0_outputs(7625);
    outputs(5912) <= (layer0_outputs(4193)) and (layer0_outputs(1675));
    outputs(5913) <= not((layer0_outputs(1472)) xor (layer0_outputs(2787)));
    outputs(5914) <= (layer0_outputs(2213)) or (layer0_outputs(2176));
    outputs(5915) <= not(layer0_outputs(3784));
    outputs(5916) <= not(layer0_outputs(5368));
    outputs(5917) <= (layer0_outputs(939)) or (layer0_outputs(4219));
    outputs(5918) <= (layer0_outputs(2857)) and not (layer0_outputs(1890));
    outputs(5919) <= layer0_outputs(3175);
    outputs(5920) <= layer0_outputs(5473);
    outputs(5921) <= layer0_outputs(5161);
    outputs(5922) <= layer0_outputs(602);
    outputs(5923) <= not(layer0_outputs(662));
    outputs(5924) <= (layer0_outputs(2522)) and not (layer0_outputs(6131));
    outputs(5925) <= not((layer0_outputs(1810)) xor (layer0_outputs(4571)));
    outputs(5926) <= not((layer0_outputs(6248)) or (layer0_outputs(3858)));
    outputs(5927) <= not((layer0_outputs(4258)) xor (layer0_outputs(790)));
    outputs(5928) <= (layer0_outputs(7454)) xor (layer0_outputs(2419));
    outputs(5929) <= not(layer0_outputs(1127));
    outputs(5930) <= layer0_outputs(802);
    outputs(5931) <= layer0_outputs(2893);
    outputs(5932) <= not(layer0_outputs(283));
    outputs(5933) <= (layer0_outputs(5244)) and not (layer0_outputs(1229));
    outputs(5934) <= not(layer0_outputs(6786));
    outputs(5935) <= not((layer0_outputs(2982)) xor (layer0_outputs(3186)));
    outputs(5936) <= not((layer0_outputs(969)) xor (layer0_outputs(5763)));
    outputs(5937) <= layer0_outputs(6442);
    outputs(5938) <= layer0_outputs(432);
    outputs(5939) <= (layer0_outputs(7053)) xor (layer0_outputs(5033));
    outputs(5940) <= (layer0_outputs(2273)) xor (layer0_outputs(5578));
    outputs(5941) <= not(layer0_outputs(285));
    outputs(5942) <= not((layer0_outputs(651)) xor (layer0_outputs(6092)));
    outputs(5943) <= not(layer0_outputs(2507));
    outputs(5944) <= not(layer0_outputs(1187));
    outputs(5945) <= layer0_outputs(3672);
    outputs(5946) <= not((layer0_outputs(4759)) or (layer0_outputs(3144)));
    outputs(5947) <= (layer0_outputs(7035)) and not (layer0_outputs(7535));
    outputs(5948) <= not((layer0_outputs(2217)) and (layer0_outputs(3123)));
    outputs(5949) <= layer0_outputs(5670);
    outputs(5950) <= layer0_outputs(4077);
    outputs(5951) <= not(layer0_outputs(3798));
    outputs(5952) <= not((layer0_outputs(2252)) or (layer0_outputs(10)));
    outputs(5953) <= (layer0_outputs(2427)) and not (layer0_outputs(5702));
    outputs(5954) <= not((layer0_outputs(5395)) or (layer0_outputs(3089)));
    outputs(5955) <= not((layer0_outputs(1162)) xor (layer0_outputs(6383)));
    outputs(5956) <= not((layer0_outputs(6772)) and (layer0_outputs(4415)));
    outputs(5957) <= not(layer0_outputs(3778));
    outputs(5958) <= layer0_outputs(3918);
    outputs(5959) <= (layer0_outputs(6994)) xor (layer0_outputs(32));
    outputs(5960) <= layer0_outputs(4623);
    outputs(5961) <= not((layer0_outputs(90)) xor (layer0_outputs(2310)));
    outputs(5962) <= (layer0_outputs(7198)) and not (layer0_outputs(2568));
    outputs(5963) <= not((layer0_outputs(2510)) xor (layer0_outputs(6347)));
    outputs(5964) <= not(layer0_outputs(476)) or (layer0_outputs(551));
    outputs(5965) <= layer0_outputs(558);
    outputs(5966) <= layer0_outputs(6926);
    outputs(5967) <= (layer0_outputs(3692)) and (layer0_outputs(6301));
    outputs(5968) <= not(layer0_outputs(2915));
    outputs(5969) <= layer0_outputs(5405);
    outputs(5970) <= not((layer0_outputs(2252)) or (layer0_outputs(3916)));
    outputs(5971) <= (layer0_outputs(1981)) xor (layer0_outputs(247));
    outputs(5972) <= layer0_outputs(3913);
    outputs(5973) <= (layer0_outputs(2742)) xor (layer0_outputs(2783));
    outputs(5974) <= (layer0_outputs(7102)) or (layer0_outputs(3966));
    outputs(5975) <= layer0_outputs(6903);
    outputs(5976) <= (layer0_outputs(6051)) and not (layer0_outputs(2724));
    outputs(5977) <= layer0_outputs(6753);
    outputs(5978) <= layer0_outputs(3944);
    outputs(5979) <= not(layer0_outputs(4885));
    outputs(5980) <= (layer0_outputs(6241)) xor (layer0_outputs(6952));
    outputs(5981) <= not(layer0_outputs(6141));
    outputs(5982) <= (layer0_outputs(376)) and not (layer0_outputs(4713));
    outputs(5983) <= layer0_outputs(5215);
    outputs(5984) <= not((layer0_outputs(1883)) or (layer0_outputs(3844)));
    outputs(5985) <= not((layer0_outputs(3927)) and (layer0_outputs(1994)));
    outputs(5986) <= (layer0_outputs(2468)) and (layer0_outputs(7530));
    outputs(5987) <= (layer0_outputs(2024)) and (layer0_outputs(1112));
    outputs(5988) <= (layer0_outputs(2066)) and not (layer0_outputs(3506));
    outputs(5989) <= (layer0_outputs(2481)) and not (layer0_outputs(5045));
    outputs(5990) <= not((layer0_outputs(7277)) xor (layer0_outputs(1706)));
    outputs(5991) <= not(layer0_outputs(1017));
    outputs(5992) <= (layer0_outputs(7454)) and not (layer0_outputs(3323));
    outputs(5993) <= layer0_outputs(4258);
    outputs(5994) <= layer0_outputs(1965);
    outputs(5995) <= layer0_outputs(5735);
    outputs(5996) <= not(layer0_outputs(3470));
    outputs(5997) <= layer0_outputs(5108);
    outputs(5998) <= (layer0_outputs(601)) and (layer0_outputs(5470));
    outputs(5999) <= layer0_outputs(2949);
    outputs(6000) <= not(layer0_outputs(2679)) or (layer0_outputs(1085));
    outputs(6001) <= layer0_outputs(7352);
    outputs(6002) <= (layer0_outputs(1904)) and not (layer0_outputs(6278));
    outputs(6003) <= (layer0_outputs(1019)) and not (layer0_outputs(2722));
    outputs(6004) <= (layer0_outputs(7003)) xor (layer0_outputs(2405));
    outputs(6005) <= (layer0_outputs(3446)) and (layer0_outputs(1698));
    outputs(6006) <= (layer0_outputs(2415)) and not (layer0_outputs(1400));
    outputs(6007) <= (layer0_outputs(2448)) and (layer0_outputs(3252));
    outputs(6008) <= not((layer0_outputs(2412)) and (layer0_outputs(1715)));
    outputs(6009) <= (layer0_outputs(314)) and not (layer0_outputs(5284));
    outputs(6010) <= not((layer0_outputs(5491)) xor (layer0_outputs(5933)));
    outputs(6011) <= (layer0_outputs(5462)) xor (layer0_outputs(6290));
    outputs(6012) <= layer0_outputs(6277);
    outputs(6013) <= (layer0_outputs(4597)) and (layer0_outputs(1687));
    outputs(6014) <= (layer0_outputs(379)) and not (layer0_outputs(3327));
    outputs(6015) <= (layer0_outputs(3296)) and not (layer0_outputs(7475));
    outputs(6016) <= layer0_outputs(5122);
    outputs(6017) <= layer0_outputs(2896);
    outputs(6018) <= not(layer0_outputs(1184));
    outputs(6019) <= not((layer0_outputs(1834)) xor (layer0_outputs(4122)));
    outputs(6020) <= layer0_outputs(6862);
    outputs(6021) <= not(layer0_outputs(5488));
    outputs(6022) <= not(layer0_outputs(2214));
    outputs(6023) <= layer0_outputs(2185);
    outputs(6024) <= layer0_outputs(3787);
    outputs(6025) <= not((layer0_outputs(5282)) xor (layer0_outputs(2296)));
    outputs(6026) <= not(layer0_outputs(489)) or (layer0_outputs(317));
    outputs(6027) <= (layer0_outputs(2540)) and not (layer0_outputs(3052));
    outputs(6028) <= layer0_outputs(2263);
    outputs(6029) <= layer0_outputs(6899);
    outputs(6030) <= layer0_outputs(4951);
    outputs(6031) <= (layer0_outputs(6158)) and (layer0_outputs(2832));
    outputs(6032) <= not(layer0_outputs(204));
    outputs(6033) <= not(layer0_outputs(921));
    outputs(6034) <= not(layer0_outputs(3578));
    outputs(6035) <= not((layer0_outputs(2707)) xor (layer0_outputs(4545)));
    outputs(6036) <= not((layer0_outputs(6207)) xor (layer0_outputs(553)));
    outputs(6037) <= (layer0_outputs(7299)) and not (layer0_outputs(3073));
    outputs(6038) <= (layer0_outputs(6276)) and not (layer0_outputs(1016));
    outputs(6039) <= not((layer0_outputs(6141)) xor (layer0_outputs(5577)));
    outputs(6040) <= not(layer0_outputs(6443));
    outputs(6041) <= (layer0_outputs(988)) and not (layer0_outputs(854));
    outputs(6042) <= not((layer0_outputs(1717)) xor (layer0_outputs(4362)));
    outputs(6043) <= not((layer0_outputs(6700)) and (layer0_outputs(4877)));
    outputs(6044) <= layer0_outputs(5800);
    outputs(6045) <= layer0_outputs(5815);
    outputs(6046) <= not(layer0_outputs(5222));
    outputs(6047) <= layer0_outputs(6839);
    outputs(6048) <= (layer0_outputs(1799)) and (layer0_outputs(1735));
    outputs(6049) <= not(layer0_outputs(4723));
    outputs(6050) <= layer0_outputs(3090);
    outputs(6051) <= (layer0_outputs(3098)) and not (layer0_outputs(2550));
    outputs(6052) <= (layer0_outputs(5120)) and not (layer0_outputs(1688));
    outputs(6053) <= layer0_outputs(2148);
    outputs(6054) <= (layer0_outputs(7273)) xor (layer0_outputs(3575));
    outputs(6055) <= (layer0_outputs(3818)) and (layer0_outputs(1419));
    outputs(6056) <= (layer0_outputs(6510)) and not (layer0_outputs(4992));
    outputs(6057) <= (layer0_outputs(5745)) xor (layer0_outputs(5883));
    outputs(6058) <= not(layer0_outputs(1061));
    outputs(6059) <= not((layer0_outputs(1974)) and (layer0_outputs(870)));
    outputs(6060) <= not(layer0_outputs(1782));
    outputs(6061) <= not(layer0_outputs(2612));
    outputs(6062) <= layer0_outputs(2280);
    outputs(6063) <= (layer0_outputs(3313)) xor (layer0_outputs(5805));
    outputs(6064) <= (layer0_outputs(518)) and (layer0_outputs(242));
    outputs(6065) <= not(layer0_outputs(3302));
    outputs(6066) <= (layer0_outputs(2620)) xor (layer0_outputs(6281));
    outputs(6067) <= (layer0_outputs(5027)) and not (layer0_outputs(5798));
    outputs(6068) <= layer0_outputs(2240);
    outputs(6069) <= layer0_outputs(2338);
    outputs(6070) <= not((layer0_outputs(1141)) xor (layer0_outputs(650)));
    outputs(6071) <= layer0_outputs(175);
    outputs(6072) <= not(layer0_outputs(3408));
    outputs(6073) <= not((layer0_outputs(5932)) xor (layer0_outputs(3549)));
    outputs(6074) <= not(layer0_outputs(1744));
    outputs(6075) <= (layer0_outputs(3920)) xor (layer0_outputs(3486));
    outputs(6076) <= layer0_outputs(2247);
    outputs(6077) <= not(layer0_outputs(2124));
    outputs(6078) <= (layer0_outputs(4876)) xor (layer0_outputs(6238));
    outputs(6079) <= not((layer0_outputs(727)) xor (layer0_outputs(2123)));
    outputs(6080) <= (layer0_outputs(4166)) xor (layer0_outputs(5435));
    outputs(6081) <= (layer0_outputs(7364)) and not (layer0_outputs(7254));
    outputs(6082) <= not((layer0_outputs(2986)) or (layer0_outputs(5605)));
    outputs(6083) <= layer0_outputs(4064);
    outputs(6084) <= not(layer0_outputs(667));
    outputs(6085) <= not(layer0_outputs(4818));
    outputs(6086) <= not(layer0_outputs(4709));
    outputs(6087) <= (layer0_outputs(3972)) xor (layer0_outputs(1600));
    outputs(6088) <= not(layer0_outputs(7460));
    outputs(6089) <= (layer0_outputs(7328)) or (layer0_outputs(7518));
    outputs(6090) <= not((layer0_outputs(7617)) xor (layer0_outputs(1861)));
    outputs(6091) <= layer0_outputs(5219);
    outputs(6092) <= not((layer0_outputs(5289)) and (layer0_outputs(3169)));
    outputs(6093) <= layer0_outputs(5167);
    outputs(6094) <= not((layer0_outputs(3801)) or (layer0_outputs(4424)));
    outputs(6095) <= not(layer0_outputs(923));
    outputs(6096) <= (layer0_outputs(2346)) xor (layer0_outputs(851));
    outputs(6097) <= (layer0_outputs(4772)) and not (layer0_outputs(509));
    outputs(6098) <= (layer0_outputs(5522)) xor (layer0_outputs(7456));
    outputs(6099) <= (layer0_outputs(5334)) and not (layer0_outputs(4913));
    outputs(6100) <= not((layer0_outputs(4949)) xor (layer0_outputs(3897)));
    outputs(6101) <= not((layer0_outputs(2428)) or (layer0_outputs(2192)));
    outputs(6102) <= (layer0_outputs(3513)) or (layer0_outputs(1510));
    outputs(6103) <= not(layer0_outputs(5525)) or (layer0_outputs(2390));
    outputs(6104) <= not(layer0_outputs(3914));
    outputs(6105) <= (layer0_outputs(4892)) and not (layer0_outputs(3169));
    outputs(6106) <= not(layer0_outputs(7057));
    outputs(6107) <= layer0_outputs(1363);
    outputs(6108) <= not(layer0_outputs(6239));
    outputs(6109) <= not((layer0_outputs(5776)) xor (layer0_outputs(1264)));
    outputs(6110) <= not((layer0_outputs(5743)) or (layer0_outputs(2860)));
    outputs(6111) <= '0';
    outputs(6112) <= layer0_outputs(1803);
    outputs(6113) <= (layer0_outputs(1219)) and not (layer0_outputs(6421));
    outputs(6114) <= layer0_outputs(7227);
    outputs(6115) <= (layer0_outputs(194)) or (layer0_outputs(6089));
    outputs(6116) <= not(layer0_outputs(6441)) or (layer0_outputs(1115));
    outputs(6117) <= layer0_outputs(2976);
    outputs(6118) <= (layer0_outputs(6874)) and (layer0_outputs(1337));
    outputs(6119) <= not(layer0_outputs(801));
    outputs(6120) <= (layer0_outputs(4988)) xor (layer0_outputs(643));
    outputs(6121) <= not((layer0_outputs(7339)) xor (layer0_outputs(220)));
    outputs(6122) <= not(layer0_outputs(3225));
    outputs(6123) <= not((layer0_outputs(1534)) and (layer0_outputs(396)));
    outputs(6124) <= not(layer0_outputs(5752));
    outputs(6125) <= not(layer0_outputs(2345));
    outputs(6126) <= not(layer0_outputs(4585));
    outputs(6127) <= '0';
    outputs(6128) <= not((layer0_outputs(4701)) or (layer0_outputs(1852)));
    outputs(6129) <= not((layer0_outputs(5466)) xor (layer0_outputs(5921)));
    outputs(6130) <= (layer0_outputs(1850)) and (layer0_outputs(6422));
    outputs(6131) <= (layer0_outputs(2784)) and (layer0_outputs(1528));
    outputs(6132) <= layer0_outputs(4218);
    outputs(6133) <= not((layer0_outputs(6597)) or (layer0_outputs(4497)));
    outputs(6134) <= (layer0_outputs(2204)) xor (layer0_outputs(5086));
    outputs(6135) <= layer0_outputs(302);
    outputs(6136) <= not((layer0_outputs(5299)) xor (layer0_outputs(7469)));
    outputs(6137) <= not((layer0_outputs(6180)) or (layer0_outputs(3538)));
    outputs(6138) <= not(layer0_outputs(4551));
    outputs(6139) <= (layer0_outputs(7117)) or (layer0_outputs(176));
    outputs(6140) <= (layer0_outputs(6932)) and not (layer0_outputs(2173));
    outputs(6141) <= layer0_outputs(3971);
    outputs(6142) <= not(layer0_outputs(4981)) or (layer0_outputs(7333));
    outputs(6143) <= (layer0_outputs(760)) xor (layer0_outputs(5302));
    outputs(6144) <= layer0_outputs(2829);
    outputs(6145) <= not((layer0_outputs(4984)) xor (layer0_outputs(6394)));
    outputs(6146) <= not((layer0_outputs(6950)) or (layer0_outputs(4574)));
    outputs(6147) <= (layer0_outputs(4651)) and (layer0_outputs(4251));
    outputs(6148) <= (layer0_outputs(4719)) and not (layer0_outputs(4715));
    outputs(6149) <= (layer0_outputs(1706)) xor (layer0_outputs(1378));
    outputs(6150) <= (layer0_outputs(3468)) xor (layer0_outputs(3185));
    outputs(6151) <= not((layer0_outputs(2627)) xor (layer0_outputs(4163)));
    outputs(6152) <= (layer0_outputs(2305)) and not (layer0_outputs(5472));
    outputs(6153) <= not((layer0_outputs(3680)) xor (layer0_outputs(1678)));
    outputs(6154) <= not(layer0_outputs(7200));
    outputs(6155) <= (layer0_outputs(5770)) and not (layer0_outputs(1473));
    outputs(6156) <= (layer0_outputs(3835)) xor (layer0_outputs(2367));
    outputs(6157) <= layer0_outputs(2743);
    outputs(6158) <= not(layer0_outputs(7011)) or (layer0_outputs(1607));
    outputs(6159) <= (layer0_outputs(5419)) xor (layer0_outputs(257));
    outputs(6160) <= not(layer0_outputs(6869));
    outputs(6161) <= layer0_outputs(705);
    outputs(6162) <= not(layer0_outputs(5226));
    outputs(6163) <= (layer0_outputs(3352)) and not (layer0_outputs(6142));
    outputs(6164) <= (layer0_outputs(5030)) xor (layer0_outputs(1587));
    outputs(6165) <= layer0_outputs(765);
    outputs(6166) <= not(layer0_outputs(1667));
    outputs(6167) <= layer0_outputs(4676);
    outputs(6168) <= (layer0_outputs(591)) or (layer0_outputs(6836));
    outputs(6169) <= layer0_outputs(6);
    outputs(6170) <= (layer0_outputs(6983)) xor (layer0_outputs(47));
    outputs(6171) <= not(layer0_outputs(7314));
    outputs(6172) <= not((layer0_outputs(6084)) xor (layer0_outputs(5272)));
    outputs(6173) <= (layer0_outputs(7332)) and not (layer0_outputs(4353));
    outputs(6174) <= layer0_outputs(5958);
    outputs(6175) <= (layer0_outputs(3777)) xor (layer0_outputs(6017));
    outputs(6176) <= layer0_outputs(703);
    outputs(6177) <= not(layer0_outputs(6293));
    outputs(6178) <= not(layer0_outputs(5140)) or (layer0_outputs(388));
    outputs(6179) <= not(layer0_outputs(2667));
    outputs(6180) <= not(layer0_outputs(6848));
    outputs(6181) <= (layer0_outputs(6852)) and not (layer0_outputs(3793));
    outputs(6182) <= not((layer0_outputs(2970)) or (layer0_outputs(929)));
    outputs(6183) <= (layer0_outputs(3577)) xor (layer0_outputs(7428));
    outputs(6184) <= not(layer0_outputs(6435));
    outputs(6185) <= layer0_outputs(6412);
    outputs(6186) <= not((layer0_outputs(5210)) xor (layer0_outputs(3023)));
    outputs(6187) <= (layer0_outputs(5343)) and (layer0_outputs(4596));
    outputs(6188) <= (layer0_outputs(2318)) xor (layer0_outputs(6106));
    outputs(6189) <= (layer0_outputs(4816)) xor (layer0_outputs(6451));
    outputs(6190) <= layer0_outputs(7232);
    outputs(6191) <= (layer0_outputs(687)) and not (layer0_outputs(2566));
    outputs(6192) <= (layer0_outputs(426)) and not (layer0_outputs(5420));
    outputs(6193) <= layer0_outputs(6522);
    outputs(6194) <= (layer0_outputs(1140)) xor (layer0_outputs(1931));
    outputs(6195) <= not(layer0_outputs(588));
    outputs(6196) <= not((layer0_outputs(4940)) and (layer0_outputs(853)));
    outputs(6197) <= not(layer0_outputs(225));
    outputs(6198) <= layer0_outputs(4860);
    outputs(6199) <= not(layer0_outputs(4788));
    outputs(6200) <= (layer0_outputs(1460)) xor (layer0_outputs(968));
    outputs(6201) <= (layer0_outputs(2293)) or (layer0_outputs(2023));
    outputs(6202) <= not(layer0_outputs(1332));
    outputs(6203) <= not(layer0_outputs(6331));
    outputs(6204) <= not(layer0_outputs(2107));
    outputs(6205) <= (layer0_outputs(3863)) and (layer0_outputs(748));
    outputs(6206) <= (layer0_outputs(7405)) xor (layer0_outputs(3272));
    outputs(6207) <= layer0_outputs(2002);
    outputs(6208) <= not((layer0_outputs(5547)) xor (layer0_outputs(5841)));
    outputs(6209) <= (layer0_outputs(2238)) and not (layer0_outputs(1885));
    outputs(6210) <= not(layer0_outputs(6902)) or (layer0_outputs(4599));
    outputs(6211) <= not((layer0_outputs(559)) xor (layer0_outputs(6002)));
    outputs(6212) <= layer0_outputs(3439);
    outputs(6213) <= (layer0_outputs(6114)) xor (layer0_outputs(1169));
    outputs(6214) <= not(layer0_outputs(2932)) or (layer0_outputs(3688));
    outputs(6215) <= not((layer0_outputs(1723)) xor (layer0_outputs(5302)));
    outputs(6216) <= not((layer0_outputs(4223)) xor (layer0_outputs(1555)));
    outputs(6217) <= layer0_outputs(76);
    outputs(6218) <= not(layer0_outputs(3675)) or (layer0_outputs(2559));
    outputs(6219) <= not(layer0_outputs(1066));
    outputs(6220) <= not((layer0_outputs(5356)) xor (layer0_outputs(6172)));
    outputs(6221) <= not(layer0_outputs(2973)) or (layer0_outputs(4589));
    outputs(6222) <= not(layer0_outputs(1253));
    outputs(6223) <= not(layer0_outputs(4733)) or (layer0_outputs(5610));
    outputs(6224) <= not(layer0_outputs(3151));
    outputs(6225) <= not(layer0_outputs(6559)) or (layer0_outputs(5023));
    outputs(6226) <= (layer0_outputs(5700)) and not (layer0_outputs(6201));
    outputs(6227) <= (layer0_outputs(1731)) and not (layer0_outputs(5270));
    outputs(6228) <= not(layer0_outputs(4787));
    outputs(6229) <= (layer0_outputs(3722)) and (layer0_outputs(4285));
    outputs(6230) <= not((layer0_outputs(5369)) xor (layer0_outputs(6381)));
    outputs(6231) <= '1';
    outputs(6232) <= layer0_outputs(2353);
    outputs(6233) <= not(layer0_outputs(6839));
    outputs(6234) <= not((layer0_outputs(1064)) xor (layer0_outputs(3497)));
    outputs(6235) <= (layer0_outputs(1584)) xor (layer0_outputs(1672));
    outputs(6236) <= (layer0_outputs(4700)) xor (layer0_outputs(6427));
    outputs(6237) <= (layer0_outputs(5317)) and not (layer0_outputs(737));
    outputs(6238) <= not(layer0_outputs(876)) or (layer0_outputs(7539));
    outputs(6239) <= not((layer0_outputs(6018)) xor (layer0_outputs(7587)));
    outputs(6240) <= layer0_outputs(7677);
    outputs(6241) <= (layer0_outputs(6995)) xor (layer0_outputs(5337));
    outputs(6242) <= not(layer0_outputs(6934)) or (layer0_outputs(2768));
    outputs(6243) <= not(layer0_outputs(2782));
    outputs(6244) <= (layer0_outputs(6307)) xor (layer0_outputs(2111));
    outputs(6245) <= not(layer0_outputs(450));
    outputs(6246) <= layer0_outputs(2177);
    outputs(6247) <= not(layer0_outputs(3007));
    outputs(6248) <= layer0_outputs(6800);
    outputs(6249) <= not(layer0_outputs(4728)) or (layer0_outputs(1666));
    outputs(6250) <= layer0_outputs(7030);
    outputs(6251) <= not(layer0_outputs(5820)) or (layer0_outputs(5327));
    outputs(6252) <= not(layer0_outputs(7506)) or (layer0_outputs(6195));
    outputs(6253) <= not(layer0_outputs(136));
    outputs(6254) <= (layer0_outputs(720)) xor (layer0_outputs(3601));
    outputs(6255) <= not(layer0_outputs(113));
    outputs(6256) <= not((layer0_outputs(7052)) and (layer0_outputs(1252)));
    outputs(6257) <= (layer0_outputs(788)) and not (layer0_outputs(3242));
    outputs(6258) <= not(layer0_outputs(5487)) or (layer0_outputs(1338));
    outputs(6259) <= '1';
    outputs(6260) <= layer0_outputs(2971);
    outputs(6261) <= (layer0_outputs(1264)) or (layer0_outputs(6191));
    outputs(6262) <= not(layer0_outputs(3875));
    outputs(6263) <= layer0_outputs(1106);
    outputs(6264) <= not((layer0_outputs(3027)) xor (layer0_outputs(2016)));
    outputs(6265) <= not((layer0_outputs(349)) xor (layer0_outputs(7605)));
    outputs(6266) <= layer0_outputs(5974);
    outputs(6267) <= not(layer0_outputs(6388));
    outputs(6268) <= layer0_outputs(987);
    outputs(6269) <= not(layer0_outputs(1282));
    outputs(6270) <= layer0_outputs(688);
    outputs(6271) <= (layer0_outputs(1401)) xor (layer0_outputs(1156));
    outputs(6272) <= not(layer0_outputs(5537));
    outputs(6273) <= (layer0_outputs(107)) and not (layer0_outputs(1301));
    outputs(6274) <= layer0_outputs(5886);
    outputs(6275) <= not(layer0_outputs(1434));
    outputs(6276) <= layer0_outputs(2020);
    outputs(6277) <= (layer0_outputs(5996)) xor (layer0_outputs(2234));
    outputs(6278) <= not(layer0_outputs(1019));
    outputs(6279) <= not((layer0_outputs(6755)) and (layer0_outputs(3257)));
    outputs(6280) <= (layer0_outputs(1274)) and (layer0_outputs(7054));
    outputs(6281) <= not(layer0_outputs(6811)) or (layer0_outputs(4792));
    outputs(6282) <= not(layer0_outputs(6459));
    outputs(6283) <= not((layer0_outputs(3463)) and (layer0_outputs(782)));
    outputs(6284) <= not((layer0_outputs(1670)) xor (layer0_outputs(3432)));
    outputs(6285) <= (layer0_outputs(6477)) xor (layer0_outputs(4564));
    outputs(6286) <= not((layer0_outputs(3145)) or (layer0_outputs(764)));
    outputs(6287) <= layer0_outputs(6742);
    outputs(6288) <= not((layer0_outputs(7273)) xor (layer0_outputs(5894)));
    outputs(6289) <= not(layer0_outputs(7254)) or (layer0_outputs(5608));
    outputs(6290) <= not(layer0_outputs(162));
    outputs(6291) <= not(layer0_outputs(4460)) or (layer0_outputs(1988));
    outputs(6292) <= (layer0_outputs(1522)) xor (layer0_outputs(776));
    outputs(6293) <= not(layer0_outputs(365));
    outputs(6294) <= (layer0_outputs(6350)) xor (layer0_outputs(797));
    outputs(6295) <= not(layer0_outputs(5316));
    outputs(6296) <= (layer0_outputs(7146)) xor (layer0_outputs(287));
    outputs(6297) <= not((layer0_outputs(7554)) and (layer0_outputs(7181)));
    outputs(6298) <= not(layer0_outputs(3217));
    outputs(6299) <= layer0_outputs(1612);
    outputs(6300) <= (layer0_outputs(3402)) and not (layer0_outputs(311));
    outputs(6301) <= (layer0_outputs(3279)) and not (layer0_outputs(7177));
    outputs(6302) <= '1';
    outputs(6303) <= (layer0_outputs(5616)) and (layer0_outputs(232));
    outputs(6304) <= layer0_outputs(4151);
    outputs(6305) <= not((layer0_outputs(4508)) xor (layer0_outputs(4946)));
    outputs(6306) <= (layer0_outputs(3039)) or (layer0_outputs(1691));
    outputs(6307) <= not((layer0_outputs(2908)) or (layer0_outputs(1116)));
    outputs(6308) <= not((layer0_outputs(62)) xor (layer0_outputs(5466)));
    outputs(6309) <= not((layer0_outputs(6622)) xor (layer0_outputs(3657)));
    outputs(6310) <= (layer0_outputs(5882)) xor (layer0_outputs(1914));
    outputs(6311) <= not(layer0_outputs(361));
    outputs(6312) <= layer0_outputs(6251);
    outputs(6313) <= layer0_outputs(4974);
    outputs(6314) <= not((layer0_outputs(5139)) xor (layer0_outputs(3493)));
    outputs(6315) <= not(layer0_outputs(3343));
    outputs(6316) <= layer0_outputs(4148);
    outputs(6317) <= (layer0_outputs(518)) and not (layer0_outputs(798));
    outputs(6318) <= not((layer0_outputs(937)) or (layer0_outputs(2282)));
    outputs(6319) <= (layer0_outputs(6739)) xor (layer0_outputs(5075));
    outputs(6320) <= layer0_outputs(6315);
    outputs(6321) <= not(layer0_outputs(4900));
    outputs(6322) <= layer0_outputs(4719);
    outputs(6323) <= (layer0_outputs(6042)) xor (layer0_outputs(693));
    outputs(6324) <= layer0_outputs(7027);
    outputs(6325) <= (layer0_outputs(14)) and (layer0_outputs(1771));
    outputs(6326) <= layer0_outputs(3076);
    outputs(6327) <= not((layer0_outputs(6199)) xor (layer0_outputs(4794)));
    outputs(6328) <= not(layer0_outputs(1951));
    outputs(6329) <= not(layer0_outputs(2659));
    outputs(6330) <= layer0_outputs(1211);
    outputs(6331) <= (layer0_outputs(3641)) or (layer0_outputs(5018));
    outputs(6332) <= layer0_outputs(4965);
    outputs(6333) <= layer0_outputs(2792);
    outputs(6334) <= (layer0_outputs(1547)) or (layer0_outputs(3859));
    outputs(6335) <= not(layer0_outputs(6763)) or (layer0_outputs(1133));
    outputs(6336) <= layer0_outputs(6567);
    outputs(6337) <= (layer0_outputs(3190)) and not (layer0_outputs(3911));
    outputs(6338) <= layer0_outputs(6843);
    outputs(6339) <= not(layer0_outputs(2022));
    outputs(6340) <= not(layer0_outputs(3891));
    outputs(6341) <= not((layer0_outputs(1433)) xor (layer0_outputs(5121)));
    outputs(6342) <= (layer0_outputs(1880)) or (layer0_outputs(6488));
    outputs(6343) <= not((layer0_outputs(7168)) xor (layer0_outputs(7416)));
    outputs(6344) <= layer0_outputs(147);
    outputs(6345) <= not((layer0_outputs(2794)) xor (layer0_outputs(1602)));
    outputs(6346) <= not(layer0_outputs(3010));
    outputs(6347) <= (layer0_outputs(4904)) xor (layer0_outputs(5427));
    outputs(6348) <= not((layer0_outputs(609)) xor (layer0_outputs(7574)));
    outputs(6349) <= layer0_outputs(3545);
    outputs(6350) <= not(layer0_outputs(4643));
    outputs(6351) <= (layer0_outputs(1999)) and not (layer0_outputs(2982));
    outputs(6352) <= (layer0_outputs(3600)) xor (layer0_outputs(3679));
    outputs(6353) <= not(layer0_outputs(623));
    outputs(6354) <= layer0_outputs(977);
    outputs(6355) <= not((layer0_outputs(3265)) xor (layer0_outputs(3844)));
    outputs(6356) <= not((layer0_outputs(693)) and (layer0_outputs(2358)));
    outputs(6357) <= layer0_outputs(2178);
    outputs(6358) <= not(layer0_outputs(1256)) or (layer0_outputs(4101));
    outputs(6359) <= (layer0_outputs(5369)) and not (layer0_outputs(6547));
    outputs(6360) <= (layer0_outputs(4255)) xor (layer0_outputs(3752));
    outputs(6361) <= (layer0_outputs(104)) xor (layer0_outputs(6065));
    outputs(6362) <= (layer0_outputs(681)) xor (layer0_outputs(5382));
    outputs(6363) <= (layer0_outputs(4716)) and (layer0_outputs(3508));
    outputs(6364) <= layer0_outputs(1883);
    outputs(6365) <= not(layer0_outputs(2325)) or (layer0_outputs(3012));
    outputs(6366) <= '1';
    outputs(6367) <= layer0_outputs(5409);
    outputs(6368) <= (layer0_outputs(112)) and not (layer0_outputs(3176));
    outputs(6369) <= not((layer0_outputs(3526)) xor (layer0_outputs(4050)));
    outputs(6370) <= (layer0_outputs(5631)) xor (layer0_outputs(3292));
    outputs(6371) <= (layer0_outputs(1154)) xor (layer0_outputs(3812));
    outputs(6372) <= layer0_outputs(2602);
    outputs(6373) <= layer0_outputs(5325);
    outputs(6374) <= not(layer0_outputs(3401));
    outputs(6375) <= not((layer0_outputs(7441)) and (layer0_outputs(7113)));
    outputs(6376) <= layer0_outputs(4503);
    outputs(6377) <= not(layer0_outputs(6531)) or (layer0_outputs(4046));
    outputs(6378) <= layer0_outputs(1781);
    outputs(6379) <= layer0_outputs(607);
    outputs(6380) <= not(layer0_outputs(6799));
    outputs(6381) <= layer0_outputs(4955);
    outputs(6382) <= not(layer0_outputs(5467));
    outputs(6383) <= (layer0_outputs(6165)) and (layer0_outputs(4280));
    outputs(6384) <= (layer0_outputs(4743)) xor (layer0_outputs(6031));
    outputs(6385) <= layer0_outputs(2113);
    outputs(6386) <= not(layer0_outputs(7327));
    outputs(6387) <= layer0_outputs(2627);
    outputs(6388) <= not((layer0_outputs(761)) xor (layer0_outputs(3695)));
    outputs(6389) <= not(layer0_outputs(150));
    outputs(6390) <= (layer0_outputs(5983)) xor (layer0_outputs(3568));
    outputs(6391) <= not((layer0_outputs(3979)) or (layer0_outputs(1462)));
    outputs(6392) <= (layer0_outputs(6648)) xor (layer0_outputs(4306));
    outputs(6393) <= not(layer0_outputs(7308));
    outputs(6394) <= layer0_outputs(5604);
    outputs(6395) <= not(layer0_outputs(1398));
    outputs(6396) <= (layer0_outputs(3151)) xor (layer0_outputs(1506));
    outputs(6397) <= (layer0_outputs(4138)) and not (layer0_outputs(4057));
    outputs(6398) <= not(layer0_outputs(675));
    outputs(6399) <= (layer0_outputs(7326)) and (layer0_outputs(3933));
    outputs(6400) <= not(layer0_outputs(6153));
    outputs(6401) <= not((layer0_outputs(1926)) or (layer0_outputs(7455)));
    outputs(6402) <= not(layer0_outputs(2879));
    outputs(6403) <= not(layer0_outputs(1778)) or (layer0_outputs(5975));
    outputs(6404) <= not(layer0_outputs(701)) or (layer0_outputs(4641));
    outputs(6405) <= not((layer0_outputs(2835)) xor (layer0_outputs(886)));
    outputs(6406) <= layer0_outputs(1224);
    outputs(6407) <= not((layer0_outputs(1823)) xor (layer0_outputs(643)));
    outputs(6408) <= (layer0_outputs(1651)) and not (layer0_outputs(5718));
    outputs(6409) <= (layer0_outputs(2702)) xor (layer0_outputs(3292));
    outputs(6410) <= not(layer0_outputs(5339));
    outputs(6411) <= '1';
    outputs(6412) <= layer0_outputs(7651);
    outputs(6413) <= (layer0_outputs(1707)) xor (layer0_outputs(924));
    outputs(6414) <= layer0_outputs(670);
    outputs(6415) <= not(layer0_outputs(4609));
    outputs(6416) <= (layer0_outputs(5881)) xor (layer0_outputs(6450));
    outputs(6417) <= (layer0_outputs(6064)) and not (layer0_outputs(5323));
    outputs(6418) <= not((layer0_outputs(7009)) and (layer0_outputs(3334)));
    outputs(6419) <= not(layer0_outputs(4941));
    outputs(6420) <= not(layer0_outputs(6539));
    outputs(6421) <= not(layer0_outputs(2446));
    outputs(6422) <= not(layer0_outputs(3201));
    outputs(6423) <= not(layer0_outputs(473));
    outputs(6424) <= layer0_outputs(6025);
    outputs(6425) <= layer0_outputs(5132);
    outputs(6426) <= not(layer0_outputs(2475));
    outputs(6427) <= not((layer0_outputs(1040)) xor (layer0_outputs(2278)));
    outputs(6428) <= (layer0_outputs(6822)) and not (layer0_outputs(3534));
    outputs(6429) <= (layer0_outputs(1623)) and (layer0_outputs(2570));
    outputs(6430) <= layer0_outputs(472);
    outputs(6431) <= not((layer0_outputs(355)) or (layer0_outputs(893)));
    outputs(6432) <= not(layer0_outputs(3855));
    outputs(6433) <= not((layer0_outputs(6312)) and (layer0_outputs(6927)));
    outputs(6434) <= (layer0_outputs(1439)) xor (layer0_outputs(1413));
    outputs(6435) <= (layer0_outputs(1393)) xor (layer0_outputs(7385));
    outputs(6436) <= not(layer0_outputs(4173)) or (layer0_outputs(716));
    outputs(6437) <= (layer0_outputs(7257)) xor (layer0_outputs(1108));
    outputs(6438) <= layer0_outputs(418);
    outputs(6439) <= (layer0_outputs(3269)) xor (layer0_outputs(4780));
    outputs(6440) <= (layer0_outputs(4392)) and not (layer0_outputs(2186));
    outputs(6441) <= not(layer0_outputs(7367));
    outputs(6442) <= not(layer0_outputs(341));
    outputs(6443) <= layer0_outputs(3976);
    outputs(6444) <= (layer0_outputs(7001)) xor (layer0_outputs(4022));
    outputs(6445) <= not(layer0_outputs(2647)) or (layer0_outputs(1785));
    outputs(6446) <= (layer0_outputs(6736)) xor (layer0_outputs(1854));
    outputs(6447) <= not((layer0_outputs(3404)) xor (layer0_outputs(6885)));
    outputs(6448) <= not((layer0_outputs(6993)) xor (layer0_outputs(6586)));
    outputs(6449) <= (layer0_outputs(4066)) or (layer0_outputs(6957));
    outputs(6450) <= layer0_outputs(5110);
    outputs(6451) <= (layer0_outputs(1720)) and not (layer0_outputs(1358));
    outputs(6452) <= not((layer0_outputs(2955)) xor (layer0_outputs(7062)));
    outputs(6453) <= (layer0_outputs(1844)) and not (layer0_outputs(5524));
    outputs(6454) <= (layer0_outputs(6627)) and not (layer0_outputs(7464));
    outputs(6455) <= not(layer0_outputs(408));
    outputs(6456) <= not(layer0_outputs(4781)) or (layer0_outputs(3771));
    outputs(6457) <= not((layer0_outputs(2723)) xor (layer0_outputs(5582)));
    outputs(6458) <= layer0_outputs(6361);
    outputs(6459) <= '1';
    outputs(6460) <= layer0_outputs(2077);
    outputs(6461) <= (layer0_outputs(2843)) and (layer0_outputs(5761));
    outputs(6462) <= not((layer0_outputs(1514)) and (layer0_outputs(3063)));
    outputs(6463) <= (layer0_outputs(2569)) and not (layer0_outputs(4264));
    outputs(6464) <= not(layer0_outputs(1258));
    outputs(6465) <= (layer0_outputs(2191)) or (layer0_outputs(2961));
    outputs(6466) <= not((layer0_outputs(6156)) or (layer0_outputs(5456)));
    outputs(6467) <= (layer0_outputs(5499)) and not (layer0_outputs(6370));
    outputs(6468) <= (layer0_outputs(5336)) or (layer0_outputs(3030));
    outputs(6469) <= (layer0_outputs(1167)) xor (layer0_outputs(4297));
    outputs(6470) <= layer0_outputs(6561);
    outputs(6471) <= not(layer0_outputs(1415)) or (layer0_outputs(7581));
    outputs(6472) <= layer0_outputs(5111);
    outputs(6473) <= (layer0_outputs(6419)) xor (layer0_outputs(7013));
    outputs(6474) <= layer0_outputs(2832);
    outputs(6475) <= (layer0_outputs(531)) xor (layer0_outputs(3877));
    outputs(6476) <= not(layer0_outputs(7578));
    outputs(6477) <= (layer0_outputs(6097)) and not (layer0_outputs(7412));
    outputs(6478) <= not(layer0_outputs(1703)) or (layer0_outputs(2959));
    outputs(6479) <= layer0_outputs(5040);
    outputs(6480) <= not((layer0_outputs(5731)) xor (layer0_outputs(4559)));
    outputs(6481) <= (layer0_outputs(1762)) xor (layer0_outputs(7378));
    outputs(6482) <= not((layer0_outputs(2351)) xor (layer0_outputs(1929)));
    outputs(6483) <= layer0_outputs(4101);
    outputs(6484) <= not(layer0_outputs(1118));
    outputs(6485) <= not(layer0_outputs(5758)) or (layer0_outputs(1536));
    outputs(6486) <= (layer0_outputs(6701)) or (layer0_outputs(6889));
    outputs(6487) <= (layer0_outputs(1748)) xor (layer0_outputs(4421));
    outputs(6488) <= (layer0_outputs(28)) xor (layer0_outputs(7243));
    outputs(6489) <= (layer0_outputs(1012)) xor (layer0_outputs(461));
    outputs(6490) <= not(layer0_outputs(3410)) or (layer0_outputs(5257));
    outputs(6491) <= layer0_outputs(2500);
    outputs(6492) <= not(layer0_outputs(7580));
    outputs(6493) <= (layer0_outputs(1760)) xor (layer0_outputs(6093));
    outputs(6494) <= not(layer0_outputs(3989)) or (layer0_outputs(5408));
    outputs(6495) <= not((layer0_outputs(1479)) xor (layer0_outputs(5114)));
    outputs(6496) <= (layer0_outputs(3024)) and not (layer0_outputs(7438));
    outputs(6497) <= (layer0_outputs(7193)) xor (layer0_outputs(5667));
    outputs(6498) <= (layer0_outputs(1637)) xor (layer0_outputs(3111));
    outputs(6499) <= not(layer0_outputs(7330));
    outputs(6500) <= not(layer0_outputs(5104));
    outputs(6501) <= not((layer0_outputs(7636)) xor (layer0_outputs(2061)));
    outputs(6502) <= layer0_outputs(603);
    outputs(6503) <= not(layer0_outputs(7594));
    outputs(6504) <= (layer0_outputs(2636)) xor (layer0_outputs(2639));
    outputs(6505) <= not(layer0_outputs(1868));
    outputs(6506) <= (layer0_outputs(6879)) and (layer0_outputs(7283));
    outputs(6507) <= layer0_outputs(7486);
    outputs(6508) <= (layer0_outputs(3188)) xor (layer0_outputs(1617));
    outputs(6509) <= not((layer0_outputs(5279)) and (layer0_outputs(7174)));
    outputs(6510) <= not((layer0_outputs(6961)) and (layer0_outputs(3079)));
    outputs(6511) <= not((layer0_outputs(327)) xor (layer0_outputs(7046)));
    outputs(6512) <= not((layer0_outputs(1745)) xor (layer0_outputs(5704)));
    outputs(6513) <= layer0_outputs(3503);
    outputs(6514) <= (layer0_outputs(4455)) or (layer0_outputs(1879));
    outputs(6515) <= (layer0_outputs(79)) xor (layer0_outputs(6162));
    outputs(6516) <= not(layer0_outputs(4315));
    outputs(6517) <= not((layer0_outputs(5421)) xor (layer0_outputs(7343)));
    outputs(6518) <= not(layer0_outputs(2994));
    outputs(6519) <= layer0_outputs(6257);
    outputs(6520) <= layer0_outputs(1895);
    outputs(6521) <= layer0_outputs(2512);
    outputs(6522) <= not(layer0_outputs(4556));
    outputs(6523) <= not((layer0_outputs(2525)) xor (layer0_outputs(2055)));
    outputs(6524) <= not(layer0_outputs(1023));
    outputs(6525) <= (layer0_outputs(6163)) xor (layer0_outputs(6267));
    outputs(6526) <= not(layer0_outputs(7500));
    outputs(6527) <= (layer0_outputs(7643)) xor (layer0_outputs(3815));
    outputs(6528) <= (layer0_outputs(2603)) xor (layer0_outputs(4385));
    outputs(6529) <= not(layer0_outputs(6575)) or (layer0_outputs(4140));
    outputs(6530) <= layer0_outputs(129);
    outputs(6531) <= layer0_outputs(6056);
    outputs(6532) <= not(layer0_outputs(6757));
    outputs(6533) <= layer0_outputs(678);
    outputs(6534) <= layer0_outputs(5850);
    outputs(6535) <= (layer0_outputs(1824)) xor (layer0_outputs(4944));
    outputs(6536) <= not(layer0_outputs(1657));
    outputs(6537) <= layer0_outputs(2988);
    outputs(6538) <= layer0_outputs(4485);
    outputs(6539) <= not(layer0_outputs(2920)) or (layer0_outputs(6729));
    outputs(6540) <= layer0_outputs(2795);
    outputs(6541) <= (layer0_outputs(3143)) and (layer0_outputs(402));
    outputs(6542) <= not(layer0_outputs(1303));
    outputs(6543) <= layer0_outputs(5766);
    outputs(6544) <= not((layer0_outputs(5232)) xor (layer0_outputs(1792)));
    outputs(6545) <= not(layer0_outputs(3613));
    outputs(6546) <= not(layer0_outputs(1575));
    outputs(6547) <= not((layer0_outputs(6680)) and (layer0_outputs(1332)));
    outputs(6548) <= layer0_outputs(1344);
    outputs(6549) <= layer0_outputs(950);
    outputs(6550) <= (layer0_outputs(3234)) xor (layer0_outputs(2201));
    outputs(6551) <= (layer0_outputs(5613)) xor (layer0_outputs(4413));
    outputs(6552) <= (layer0_outputs(3457)) or (layer0_outputs(4605));
    outputs(6553) <= not(layer0_outputs(290));
    outputs(6554) <= not(layer0_outputs(1693));
    outputs(6555) <= not(layer0_outputs(2993)) or (layer0_outputs(4055));
    outputs(6556) <= not(layer0_outputs(6478));
    outputs(6557) <= (layer0_outputs(5184)) xor (layer0_outputs(3295));
    outputs(6558) <= (layer0_outputs(138)) and not (layer0_outputs(195));
    outputs(6559) <= not(layer0_outputs(3792));
    outputs(6560) <= not((layer0_outputs(4694)) xor (layer0_outputs(4569)));
    outputs(6561) <= not((layer0_outputs(4788)) or (layer0_outputs(3785)));
    outputs(6562) <= not((layer0_outputs(5786)) and (layer0_outputs(1893)));
    outputs(6563) <= layer0_outputs(54);
    outputs(6564) <= not(layer0_outputs(1923));
    outputs(6565) <= not((layer0_outputs(844)) xor (layer0_outputs(5903)));
    outputs(6566) <= not((layer0_outputs(6634)) or (layer0_outputs(7255)));
    outputs(6567) <= layer0_outputs(3156);
    outputs(6568) <= not(layer0_outputs(6362));
    outputs(6569) <= layer0_outputs(4211);
    outputs(6570) <= layer0_outputs(3061);
    outputs(6571) <= not(layer0_outputs(4495));
    outputs(6572) <= not(layer0_outputs(2440));
    outputs(6573) <= (layer0_outputs(2740)) xor (layer0_outputs(1378));
    outputs(6574) <= not((layer0_outputs(6805)) xor (layer0_outputs(6813)));
    outputs(6575) <= not(layer0_outputs(1265)) or (layer0_outputs(7515));
    outputs(6576) <= not(layer0_outputs(5803));
    outputs(6577) <= not((layer0_outputs(2225)) and (layer0_outputs(2527)));
    outputs(6578) <= not((layer0_outputs(5263)) xor (layer0_outputs(3048)));
    outputs(6579) <= (layer0_outputs(5121)) xor (layer0_outputs(6228));
    outputs(6580) <= not((layer0_outputs(2882)) xor (layer0_outputs(6125)));
    outputs(6581) <= not(layer0_outputs(3523));
    outputs(6582) <= not(layer0_outputs(7199));
    outputs(6583) <= '1';
    outputs(6584) <= layer0_outputs(567);
    outputs(6585) <= not(layer0_outputs(6229));
    outputs(6586) <= not((layer0_outputs(4731)) xor (layer0_outputs(6715)));
    outputs(6587) <= not((layer0_outputs(7110)) xor (layer0_outputs(6718)));
    outputs(6588) <= not((layer0_outputs(34)) xor (layer0_outputs(5180)));
    outputs(6589) <= (layer0_outputs(5732)) xor (layer0_outputs(4626));
    outputs(6590) <= not(layer0_outputs(336));
    outputs(6591) <= not(layer0_outputs(5152)) or (layer0_outputs(2560));
    outputs(6592) <= not((layer0_outputs(4766)) and (layer0_outputs(7307)));
    outputs(6593) <= not(layer0_outputs(7297));
    outputs(6594) <= layer0_outputs(1560);
    outputs(6595) <= (layer0_outputs(7459)) and not (layer0_outputs(4658));
    outputs(6596) <= layer0_outputs(340);
    outputs(6597) <= not(layer0_outputs(646)) or (layer0_outputs(4189));
    outputs(6598) <= not(layer0_outputs(4932));
    outputs(6599) <= layer0_outputs(4061);
    outputs(6600) <= not(layer0_outputs(5177)) or (layer0_outputs(7253));
    outputs(6601) <= (layer0_outputs(7578)) xor (layer0_outputs(273));
    outputs(6602) <= (layer0_outputs(4016)) xor (layer0_outputs(3524));
    outputs(6603) <= not((layer0_outputs(6754)) xor (layer0_outputs(2353)));
    outputs(6604) <= layer0_outputs(493);
    outputs(6605) <= layer0_outputs(580);
    outputs(6606) <= (layer0_outputs(5383)) xor (layer0_outputs(4523));
    outputs(6607) <= not(layer0_outputs(4288));
    outputs(6608) <= layer0_outputs(3444);
    outputs(6609) <= (layer0_outputs(2891)) xor (layer0_outputs(3110));
    outputs(6610) <= layer0_outputs(2143);
    outputs(6611) <= not(layer0_outputs(3952));
    outputs(6612) <= not((layer0_outputs(4648)) xor (layer0_outputs(6583)));
    outputs(6613) <= not((layer0_outputs(4715)) or (layer0_outputs(1297)));
    outputs(6614) <= (layer0_outputs(4274)) and (layer0_outputs(3166));
    outputs(6615) <= (layer0_outputs(1653)) and not (layer0_outputs(2032));
    outputs(6616) <= not((layer0_outputs(5362)) xor (layer0_outputs(50)));
    outputs(6617) <= not(layer0_outputs(5144)) or (layer0_outputs(1833));
    outputs(6618) <= (layer0_outputs(6832)) xor (layer0_outputs(6603));
    outputs(6619) <= (layer0_outputs(4361)) xor (layer0_outputs(2945));
    outputs(6620) <= not(layer0_outputs(7502));
    outputs(6621) <= layer0_outputs(3449);
    outputs(6622) <= not(layer0_outputs(7549)) or (layer0_outputs(2943));
    outputs(6623) <= not(layer0_outputs(6588));
    outputs(6624) <= not(layer0_outputs(5436)) or (layer0_outputs(2454));
    outputs(6625) <= (layer0_outputs(1435)) xor (layer0_outputs(4945));
    outputs(6626) <= (layer0_outputs(1726)) and not (layer0_outputs(4229));
    outputs(6627) <= not((layer0_outputs(6247)) or (layer0_outputs(4297)));
    outputs(6628) <= not(layer0_outputs(7476));
    outputs(6629) <= not(layer0_outputs(993));
    outputs(6630) <= not(layer0_outputs(6543));
    outputs(6631) <= not((layer0_outputs(3929)) or (layer0_outputs(5577)));
    outputs(6632) <= (layer0_outputs(4337)) and not (layer0_outputs(6291));
    outputs(6633) <= layer0_outputs(2460);
    outputs(6634) <= not(layer0_outputs(2551));
    outputs(6635) <= (layer0_outputs(6572)) and not (layer0_outputs(4202));
    outputs(6636) <= not(layer0_outputs(683)) or (layer0_outputs(5201));
    outputs(6637) <= layer0_outputs(2664);
    outputs(6638) <= not(layer0_outputs(6644)) or (layer0_outputs(1709));
    outputs(6639) <= not((layer0_outputs(667)) xor (layer0_outputs(2678)));
    outputs(6640) <= not(layer0_outputs(4526));
    outputs(6641) <= layer0_outputs(2632);
    outputs(6642) <= not((layer0_outputs(1567)) xor (layer0_outputs(1539)));
    outputs(6643) <= (layer0_outputs(7662)) or (layer0_outputs(2470));
    outputs(6644) <= not(layer0_outputs(474));
    outputs(6645) <= not((layer0_outputs(1871)) xor (layer0_outputs(5797)));
    outputs(6646) <= not(layer0_outputs(1078)) or (layer0_outputs(3370));
    outputs(6647) <= not((layer0_outputs(6213)) xor (layer0_outputs(5972)));
    outputs(6648) <= not(layer0_outputs(3421));
    outputs(6649) <= not(layer0_outputs(3234)) or (layer0_outputs(4199));
    outputs(6650) <= (layer0_outputs(6301)) xor (layer0_outputs(7525));
    outputs(6651) <= not((layer0_outputs(3942)) xor (layer0_outputs(5926)));
    outputs(6652) <= not(layer0_outputs(4329));
    outputs(6653) <= (layer0_outputs(6932)) and not (layer0_outputs(148));
    outputs(6654) <= (layer0_outputs(3928)) and not (layer0_outputs(1566));
    outputs(6655) <= not((layer0_outputs(1464)) or (layer0_outputs(1139)));
    outputs(6656) <= not((layer0_outputs(4756)) xor (layer0_outputs(5759)));
    outputs(6657) <= not((layer0_outputs(5280)) xor (layer0_outputs(6226)));
    outputs(6658) <= not(layer0_outputs(5191));
    outputs(6659) <= (layer0_outputs(5152)) xor (layer0_outputs(4368));
    outputs(6660) <= not((layer0_outputs(4490)) xor (layer0_outputs(2728)));
    outputs(6661) <= layer0_outputs(1928);
    outputs(6662) <= layer0_outputs(3870);
    outputs(6663) <= not((layer0_outputs(1128)) xor (layer0_outputs(4019)));
    outputs(6664) <= not(layer0_outputs(1373)) or (layer0_outputs(2014));
    outputs(6665) <= not((layer0_outputs(2538)) xor (layer0_outputs(552)));
    outputs(6666) <= (layer0_outputs(591)) or (layer0_outputs(4521));
    outputs(6667) <= not(layer0_outputs(941));
    outputs(6668) <= not((layer0_outputs(1806)) xor (layer0_outputs(168)));
    outputs(6669) <= not(layer0_outputs(5657));
    outputs(6670) <= (layer0_outputs(2343)) xor (layer0_outputs(7343));
    outputs(6671) <= not((layer0_outputs(3922)) xor (layer0_outputs(6288)));
    outputs(6672) <= '1';
    outputs(6673) <= not(layer0_outputs(190));
    outputs(6674) <= layer0_outputs(5372);
    outputs(6675) <= (layer0_outputs(3115)) and (layer0_outputs(1858));
    outputs(6676) <= not((layer0_outputs(3088)) or (layer0_outputs(1507)));
    outputs(6677) <= (layer0_outputs(7614)) xor (layer0_outputs(6701));
    outputs(6678) <= (layer0_outputs(4541)) or (layer0_outputs(6294));
    outputs(6679) <= layer0_outputs(4192);
    outputs(6680) <= not((layer0_outputs(3827)) xor (layer0_outputs(4916)));
    outputs(6681) <= not(layer0_outputs(4432)) or (layer0_outputs(2067));
    outputs(6682) <= not(layer0_outputs(6896));
    outputs(6683) <= not((layer0_outputs(200)) xor (layer0_outputs(864)));
    outputs(6684) <= (layer0_outputs(1097)) and not (layer0_outputs(453));
    outputs(6685) <= not(layer0_outputs(7618)) or (layer0_outputs(5739));
    outputs(6686) <= layer0_outputs(5182);
    outputs(6687) <= layer0_outputs(5565);
    outputs(6688) <= not((layer0_outputs(5870)) xor (layer0_outputs(4408)));
    outputs(6689) <= not((layer0_outputs(5142)) xor (layer0_outputs(4309)));
    outputs(6690) <= (layer0_outputs(4576)) xor (layer0_outputs(5651));
    outputs(6691) <= layer0_outputs(1144);
    outputs(6692) <= layer0_outputs(1669);
    outputs(6693) <= not(layer0_outputs(2909));
    outputs(6694) <= (layer0_outputs(6200)) and (layer0_outputs(1174));
    outputs(6695) <= not(layer0_outputs(7601));
    outputs(6696) <= layer0_outputs(850);
    outputs(6697) <= not(layer0_outputs(7571));
    outputs(6698) <= (layer0_outputs(4100)) and (layer0_outputs(4581));
    outputs(6699) <= (layer0_outputs(5734)) xor (layer0_outputs(1276));
    outputs(6700) <= (layer0_outputs(281)) and not (layer0_outputs(5387));
    outputs(6701) <= (layer0_outputs(2435)) or (layer0_outputs(1699));
    outputs(6702) <= not(layer0_outputs(4893));
    outputs(6703) <= not((layer0_outputs(3400)) xor (layer0_outputs(3239)));
    outputs(6704) <= (layer0_outputs(6403)) or (layer0_outputs(4529));
    outputs(6705) <= (layer0_outputs(6652)) xor (layer0_outputs(3509));
    outputs(6706) <= (layer0_outputs(3153)) xor (layer0_outputs(4310));
    outputs(6707) <= (layer0_outputs(2294)) xor (layer0_outputs(3091));
    outputs(6708) <= layer0_outputs(846);
    outputs(6709) <= not(layer0_outputs(685));
    outputs(6710) <= not((layer0_outputs(1571)) xor (layer0_outputs(2719)));
    outputs(6711) <= not(layer0_outputs(516));
    outputs(6712) <= (layer0_outputs(347)) and not (layer0_outputs(1249));
    outputs(6713) <= layer0_outputs(1465);
    outputs(6714) <= (layer0_outputs(6733)) and (layer0_outputs(698));
    outputs(6715) <= layer0_outputs(7499);
    outputs(6716) <= not(layer0_outputs(3329)) or (layer0_outputs(1149));
    outputs(6717) <= (layer0_outputs(3955)) and (layer0_outputs(6406));
    outputs(6718) <= (layer0_outputs(3029)) xor (layer0_outputs(5009));
    outputs(6719) <= (layer0_outputs(5664)) and not (layer0_outputs(3219));
    outputs(6720) <= layer0_outputs(7096);
    outputs(6721) <= not((layer0_outputs(1342)) xor (layer0_outputs(2418)));
    outputs(6722) <= not(layer0_outputs(6421)) or (layer0_outputs(4638));
    outputs(6723) <= (layer0_outputs(3882)) xor (layer0_outputs(5723));
    outputs(6724) <= layer0_outputs(888);
    outputs(6725) <= not((layer0_outputs(4958)) xor (layer0_outputs(3230)));
    outputs(6726) <= not(layer0_outputs(6277));
    outputs(6727) <= not((layer0_outputs(6710)) xor (layer0_outputs(4894)));
    outputs(6728) <= not(layer0_outputs(4689));
    outputs(6729) <= not((layer0_outputs(721)) and (layer0_outputs(1402)));
    outputs(6730) <= layer0_outputs(6596);
    outputs(6731) <= not(layer0_outputs(7659)) or (layer0_outputs(7664));
    outputs(6732) <= not(layer0_outputs(4097));
    outputs(6733) <= (layer0_outputs(6957)) or (layer0_outputs(2488));
    outputs(6734) <= not(layer0_outputs(3158));
    outputs(6735) <= not((layer0_outputs(4076)) and (layer0_outputs(5424)));
    outputs(6736) <= (layer0_outputs(3380)) and not (layer0_outputs(6207));
    outputs(6737) <= (layer0_outputs(548)) xor (layer0_outputs(1757));
    outputs(6738) <= layer0_outputs(5441);
    outputs(6739) <= not(layer0_outputs(5100));
    outputs(6740) <= (layer0_outputs(4379)) and not (layer0_outputs(4159));
    outputs(6741) <= '1';
    outputs(6742) <= (layer0_outputs(3444)) or (layer0_outputs(6766));
    outputs(6743) <= not(layer0_outputs(7585));
    outputs(6744) <= layer0_outputs(6918);
    outputs(6745) <= (layer0_outputs(5793)) xor (layer0_outputs(5370));
    outputs(6746) <= (layer0_outputs(1167)) xor (layer0_outputs(3744));
    outputs(6747) <= not(layer0_outputs(2660));
    outputs(6748) <= not((layer0_outputs(3709)) xor (layer0_outputs(823)));
    outputs(6749) <= not(layer0_outputs(1188));
    outputs(6750) <= not(layer0_outputs(648)) or (layer0_outputs(7065));
    outputs(6751) <= layer0_outputs(1418);
    outputs(6752) <= layer0_outputs(6081);
    outputs(6753) <= not((layer0_outputs(5094)) xor (layer0_outputs(2167)));
    outputs(6754) <= not((layer0_outputs(6192)) xor (layer0_outputs(3674)));
    outputs(6755) <= layer0_outputs(2451);
    outputs(6756) <= not(layer0_outputs(7264));
    outputs(6757) <= layer0_outputs(5865);
    outputs(6758) <= (layer0_outputs(1717)) xor (layer0_outputs(1570));
    outputs(6759) <= (layer0_outputs(834)) or (layer0_outputs(6996));
    outputs(6760) <= (layer0_outputs(3785)) xor (layer0_outputs(2329));
    outputs(6761) <= (layer0_outputs(5831)) xor (layer0_outputs(5273));
    outputs(6762) <= not((layer0_outputs(6948)) xor (layer0_outputs(660)));
    outputs(6763) <= not(layer0_outputs(5544)) or (layer0_outputs(2784));
    outputs(6764) <= (layer0_outputs(7528)) xor (layer0_outputs(242));
    outputs(6765) <= not(layer0_outputs(157));
    outputs(6766) <= not((layer0_outputs(6926)) xor (layer0_outputs(5987)));
    outputs(6767) <= layer0_outputs(6810);
    outputs(6768) <= not((layer0_outputs(1581)) xor (layer0_outputs(1847)));
    outputs(6769) <= not(layer0_outputs(2738));
    outputs(6770) <= not((layer0_outputs(4997)) and (layer0_outputs(4316)));
    outputs(6771) <= not(layer0_outputs(1802));
    outputs(6772) <= layer0_outputs(5257);
    outputs(6773) <= not(layer0_outputs(1716));
    outputs(6774) <= not((layer0_outputs(6411)) xor (layer0_outputs(6358)));
    outputs(6775) <= layer0_outputs(6251);
    outputs(6776) <= (layer0_outputs(2684)) or (layer0_outputs(4425));
    outputs(6777) <= not(layer0_outputs(5711));
    outputs(6778) <= layer0_outputs(3207);
    outputs(6779) <= (layer0_outputs(84)) xor (layer0_outputs(3609));
    outputs(6780) <= (layer0_outputs(7276)) and not (layer0_outputs(6121));
    outputs(6781) <= layer0_outputs(1242);
    outputs(6782) <= not((layer0_outputs(7345)) and (layer0_outputs(5318)));
    outputs(6783) <= (layer0_outputs(3756)) xor (layer0_outputs(6353));
    outputs(6784) <= layer0_outputs(2803);
    outputs(6785) <= (layer0_outputs(6534)) xor (layer0_outputs(6700));
    outputs(6786) <= (layer0_outputs(16)) xor (layer0_outputs(2791));
    outputs(6787) <= not((layer0_outputs(3845)) xor (layer0_outputs(7565)));
    outputs(6788) <= not((layer0_outputs(1291)) xor (layer0_outputs(439)));
    outputs(6789) <= layer0_outputs(7267);
    outputs(6790) <= (layer0_outputs(530)) or (layer0_outputs(1207));
    outputs(6791) <= not(layer0_outputs(4667));
    outputs(6792) <= not((layer0_outputs(2894)) xor (layer0_outputs(1780)));
    outputs(6793) <= layer0_outputs(1365);
    outputs(6794) <= not(layer0_outputs(754));
    outputs(6795) <= (layer0_outputs(7275)) and (layer0_outputs(2488));
    outputs(6796) <= not((layer0_outputs(6419)) or (layer0_outputs(3224)));
    outputs(6797) <= (layer0_outputs(2363)) and not (layer0_outputs(3354));
    outputs(6798) <= not(layer0_outputs(6246));
    outputs(6799) <= not(layer0_outputs(6893)) or (layer0_outputs(5945));
    outputs(6800) <= layer0_outputs(4808);
    outputs(6801) <= (layer0_outputs(2762)) and not (layer0_outputs(1716));
    outputs(6802) <= not((layer0_outputs(2181)) xor (layer0_outputs(5008)));
    outputs(6803) <= not(layer0_outputs(4045)) or (layer0_outputs(1978));
    outputs(6804) <= layer0_outputs(590);
    outputs(6805) <= layer0_outputs(3521);
    outputs(6806) <= (layer0_outputs(5397)) xor (layer0_outputs(1616));
    outputs(6807) <= not(layer0_outputs(3216));
    outputs(6808) <= (layer0_outputs(7143)) xor (layer0_outputs(2779));
    outputs(6809) <= layer0_outputs(5530);
    outputs(6810) <= layer0_outputs(1991);
    outputs(6811) <= (layer0_outputs(5664)) and (layer0_outputs(1468));
    outputs(6812) <= not(layer0_outputs(3805));
    outputs(6813) <= layer0_outputs(1970);
    outputs(6814) <= not((layer0_outputs(6901)) xor (layer0_outputs(169)));
    outputs(6815) <= (layer0_outputs(5567)) xor (layer0_outputs(3808));
    outputs(6816) <= layer0_outputs(5599);
    outputs(6817) <= not(layer0_outputs(3137)) or (layer0_outputs(3089));
    outputs(6818) <= layer0_outputs(2861);
    outputs(6819) <= not(layer0_outputs(2839)) or (layer0_outputs(119));
    outputs(6820) <= (layer0_outputs(1524)) xor (layer0_outputs(6779));
    outputs(6821) <= (layer0_outputs(3178)) or (layer0_outputs(3450));
    outputs(6822) <= layer0_outputs(38);
    outputs(6823) <= not(layer0_outputs(1368));
    outputs(6824) <= not((layer0_outputs(3686)) xor (layer0_outputs(4680)));
    outputs(6825) <= not((layer0_outputs(7113)) xor (layer0_outputs(1483)));
    outputs(6826) <= layer0_outputs(626);
    outputs(6827) <= (layer0_outputs(1250)) xor (layer0_outputs(5966));
    outputs(6828) <= not((layer0_outputs(3564)) or (layer0_outputs(1086)));
    outputs(6829) <= (layer0_outputs(6433)) xor (layer0_outputs(3688));
    outputs(6830) <= layer0_outputs(2019);
    outputs(6831) <= not(layer0_outputs(1814));
    outputs(6832) <= layer0_outputs(6674);
    outputs(6833) <= layer0_outputs(524);
    outputs(6834) <= (layer0_outputs(1831)) and not (layer0_outputs(6467));
    outputs(6835) <= layer0_outputs(1138);
    outputs(6836) <= layer0_outputs(7077);
    outputs(6837) <= layer0_outputs(5204);
    outputs(6838) <= layer0_outputs(2499);
    outputs(6839) <= (layer0_outputs(6100)) and not (layer0_outputs(7624));
    outputs(6840) <= layer0_outputs(4996);
    outputs(6841) <= (layer0_outputs(6346)) or (layer0_outputs(4665));
    outputs(6842) <= layer0_outputs(5031);
    outputs(6843) <= (layer0_outputs(2926)) or (layer0_outputs(1702));
    outputs(6844) <= not(layer0_outputs(6076)) or (layer0_outputs(1289));
    outputs(6845) <= not((layer0_outputs(6731)) xor (layer0_outputs(4502)));
    outputs(6846) <= (layer0_outputs(3819)) and not (layer0_outputs(4098));
    outputs(6847) <= (layer0_outputs(7223)) and not (layer0_outputs(695));
    outputs(6848) <= layer0_outputs(1003);
    outputs(6849) <= not(layer0_outputs(2994));
    outputs(6850) <= (layer0_outputs(6703)) xor (layer0_outputs(5092));
    outputs(6851) <= (layer0_outputs(5873)) or (layer0_outputs(5899));
    outputs(6852) <= (layer0_outputs(1430)) xor (layer0_outputs(3591));
    outputs(6853) <= layer0_outputs(1347);
    outputs(6854) <= (layer0_outputs(151)) xor (layer0_outputs(4607));
    outputs(6855) <= (layer0_outputs(165)) and not (layer0_outputs(4450));
    outputs(6856) <= (layer0_outputs(141)) and not (layer0_outputs(1626));
    outputs(6857) <= (layer0_outputs(2267)) xor (layer0_outputs(2720));
    outputs(6858) <= (layer0_outputs(4110)) and not (layer0_outputs(2290));
    outputs(6859) <= not(layer0_outputs(1960)) or (layer0_outputs(4250));
    outputs(6860) <= (layer0_outputs(1478)) xor (layer0_outputs(6582));
    outputs(6861) <= (layer0_outputs(2060)) xor (layer0_outputs(4089));
    outputs(6862) <= not((layer0_outputs(1408)) or (layer0_outputs(7293)));
    outputs(6863) <= layer0_outputs(3274);
    outputs(6864) <= not(layer0_outputs(4461));
    outputs(6865) <= not(layer0_outputs(462)) or (layer0_outputs(4500));
    outputs(6866) <= (layer0_outputs(7008)) xor (layer0_outputs(292));
    outputs(6867) <= not(layer0_outputs(4727)) or (layer0_outputs(1559));
    outputs(6868) <= not((layer0_outputs(2964)) or (layer0_outputs(7129)));
    outputs(6869) <= layer0_outputs(935);
    outputs(6870) <= layer0_outputs(7219);
    outputs(6871) <= not(layer0_outputs(570));
    outputs(6872) <= (layer0_outputs(3187)) and (layer0_outputs(2740));
    outputs(6873) <= not(layer0_outputs(4790));
    outputs(6874) <= not((layer0_outputs(1922)) and (layer0_outputs(4345)));
    outputs(6875) <= layer0_outputs(5166);
    outputs(6876) <= not(layer0_outputs(199)) or (layer0_outputs(4217));
    outputs(6877) <= not((layer0_outputs(5740)) xor (layer0_outputs(228)));
    outputs(6878) <= (layer0_outputs(5129)) xor (layer0_outputs(3661));
    outputs(6879) <= not(layer0_outputs(3911));
    outputs(6880) <= not((layer0_outputs(4702)) and (layer0_outputs(7032)));
    outputs(6881) <= not((layer0_outputs(3947)) xor (layer0_outputs(3107)));
    outputs(6882) <= (layer0_outputs(1421)) xor (layer0_outputs(7047));
    outputs(6883) <= (layer0_outputs(1789)) xor (layer0_outputs(471));
    outputs(6884) <= (layer0_outputs(3126)) or (layer0_outputs(1611));
    outputs(6885) <= not(layer0_outputs(3502)) or (layer0_outputs(1704));
    outputs(6886) <= layer0_outputs(6254);
    outputs(6887) <= layer0_outputs(6411);
    outputs(6888) <= not((layer0_outputs(1030)) or (layer0_outputs(1590)));
    outputs(6889) <= not(layer0_outputs(4620)) or (layer0_outputs(5266));
    outputs(6890) <= (layer0_outputs(4988)) or (layer0_outputs(6177));
    outputs(6891) <= not((layer0_outputs(4884)) or (layer0_outputs(2312)));
    outputs(6892) <= not(layer0_outputs(1098));
    outputs(6893) <= not(layer0_outputs(2901));
    outputs(6894) <= layer0_outputs(2194);
    outputs(6895) <= (layer0_outputs(869)) xor (layer0_outputs(4135));
    outputs(6896) <= (layer0_outputs(6897)) and not (layer0_outputs(4314));
    outputs(6897) <= not((layer0_outputs(7629)) xor (layer0_outputs(2892)));
    outputs(6898) <= (layer0_outputs(3813)) or (layer0_outputs(2266));
    outputs(6899) <= not(layer0_outputs(2995));
    outputs(6900) <= not(layer0_outputs(5615));
    outputs(6901) <= (layer0_outputs(6619)) xor (layer0_outputs(7263));
    outputs(6902) <= (layer0_outputs(5288)) xor (layer0_outputs(914));
    outputs(6903) <= layer0_outputs(1535);
    outputs(6904) <= not((layer0_outputs(3734)) and (layer0_outputs(1374)));
    outputs(6905) <= (layer0_outputs(4486)) xor (layer0_outputs(5159));
    outputs(6906) <= (layer0_outputs(2139)) and (layer0_outputs(6930));
    outputs(6907) <= not(layer0_outputs(4003));
    outputs(6908) <= layer0_outputs(4160);
    outputs(6909) <= not(layer0_outputs(6366)) or (layer0_outputs(7178));
    outputs(6910) <= not((layer0_outputs(7456)) xor (layer0_outputs(1601)));
    outputs(6911) <= layer0_outputs(3479);
    outputs(6912) <= (layer0_outputs(5619)) and not (layer0_outputs(2232));
    outputs(6913) <= not((layer0_outputs(5304)) xor (layer0_outputs(5458)));
    outputs(6914) <= layer0_outputs(1210);
    outputs(6915) <= not(layer0_outputs(2324));
    outputs(6916) <= not(layer0_outputs(6884));
    outputs(6917) <= (layer0_outputs(7152)) and not (layer0_outputs(4090));
    outputs(6918) <= not(layer0_outputs(4532));
    outputs(6919) <= not(layer0_outputs(6217));
    outputs(6920) <= layer0_outputs(5947);
    outputs(6921) <= (layer0_outputs(4429)) and not (layer0_outputs(4103));
    outputs(6922) <= (layer0_outputs(1597)) and (layer0_outputs(1101));
    outputs(6923) <= (layer0_outputs(903)) and not (layer0_outputs(2239));
    outputs(6924) <= not(layer0_outputs(6534));
    outputs(6925) <= (layer0_outputs(4265)) xor (layer0_outputs(1212));
    outputs(6926) <= (layer0_outputs(519)) xor (layer0_outputs(441));
    outputs(6927) <= (layer0_outputs(2736)) and not (layer0_outputs(2696));
    outputs(6928) <= layer0_outputs(6882);
    outputs(6929) <= not((layer0_outputs(5216)) or (layer0_outputs(4950)));
    outputs(6930) <= not(layer0_outputs(5812));
    outputs(6931) <= not((layer0_outputs(3633)) xor (layer0_outputs(7383)));
    outputs(6932) <= not((layer0_outputs(7069)) or (layer0_outputs(6144)));
    outputs(6933) <= not(layer0_outputs(5980));
    outputs(6934) <= (layer0_outputs(1009)) and not (layer0_outputs(5156));
    outputs(6935) <= not(layer0_outputs(6788));
    outputs(6936) <= layer0_outputs(5070);
    outputs(6937) <= (layer0_outputs(6465)) and not (layer0_outputs(4074));
    outputs(6938) <= not((layer0_outputs(5333)) xor (layer0_outputs(133)));
    outputs(6939) <= not((layer0_outputs(1354)) and (layer0_outputs(3782)));
    outputs(6940) <= not(layer0_outputs(3740));
    outputs(6941) <= layer0_outputs(6902);
    outputs(6942) <= (layer0_outputs(6237)) and not (layer0_outputs(5510));
    outputs(6943) <= not(layer0_outputs(4257));
    outputs(6944) <= layer0_outputs(6662);
    outputs(6945) <= not(layer0_outputs(7398));
    outputs(6946) <= layer0_outputs(379);
    outputs(6947) <= (layer0_outputs(913)) xor (layer0_outputs(4775));
    outputs(6948) <= (layer0_outputs(1935)) or (layer0_outputs(1838));
    outputs(6949) <= layer0_outputs(763);
    outputs(6950) <= not(layer0_outputs(7544));
    outputs(6951) <= not((layer0_outputs(569)) or (layer0_outputs(4807)));
    outputs(6952) <= (layer0_outputs(2314)) xor (layer0_outputs(7553));
    outputs(6953) <= (layer0_outputs(7482)) and (layer0_outputs(2182));
    outputs(6954) <= layer0_outputs(1002);
    outputs(6955) <= '0';
    outputs(6956) <= not(layer0_outputs(4911));
    outputs(6957) <= (layer0_outputs(6599)) xor (layer0_outputs(1176));
    outputs(6958) <= (layer0_outputs(3112)) and not (layer0_outputs(7555));
    outputs(6959) <= not((layer0_outputs(2534)) xor (layer0_outputs(3780)));
    outputs(6960) <= not(layer0_outputs(7411)) or (layer0_outputs(7631));
    outputs(6961) <= not(layer0_outputs(3864)) or (layer0_outputs(2987));
    outputs(6962) <= layer0_outputs(1820);
    outputs(6963) <= (layer0_outputs(5115)) and (layer0_outputs(3398));
    outputs(6964) <= (layer0_outputs(5637)) and not (layer0_outputs(5418));
    outputs(6965) <= (layer0_outputs(1389)) and not (layer0_outputs(2257));
    outputs(6966) <= (layer0_outputs(782)) and not (layer0_outputs(6693));
    outputs(6967) <= (layer0_outputs(4049)) xor (layer0_outputs(4389));
    outputs(6968) <= not((layer0_outputs(7216)) xor (layer0_outputs(3932)));
    outputs(6969) <= (layer0_outputs(300)) xor (layer0_outputs(5583));
    outputs(6970) <= '0';
    outputs(6971) <= layer0_outputs(7648);
    outputs(6972) <= layer0_outputs(2937);
    outputs(6973) <= not(layer0_outputs(3754));
    outputs(6974) <= layer0_outputs(4482);
    outputs(6975) <= not(layer0_outputs(2912));
    outputs(6976) <= (layer0_outputs(4044)) and (layer0_outputs(7557));
    outputs(6977) <= layer0_outputs(2377);
    outputs(6978) <= layer0_outputs(3121);
    outputs(6979) <= not(layer0_outputs(1109));
    outputs(6980) <= (layer0_outputs(5918)) xor (layer0_outputs(3773));
    outputs(6981) <= (layer0_outputs(3441)) and not (layer0_outputs(2923));
    outputs(6982) <= layer0_outputs(2911);
    outputs(6983) <= not((layer0_outputs(5149)) xor (layer0_outputs(5436)));
    outputs(6984) <= (layer0_outputs(6430)) and (layer0_outputs(2720));
    outputs(6985) <= not((layer0_outputs(872)) or (layer0_outputs(801)));
    outputs(6986) <= (layer0_outputs(3879)) xor (layer0_outputs(1629));
    outputs(6987) <= not(layer0_outputs(4997)) or (layer0_outputs(6787));
    outputs(6988) <= not((layer0_outputs(3094)) or (layer0_outputs(2578)));
    outputs(6989) <= (layer0_outputs(6995)) and not (layer0_outputs(72));
    outputs(6990) <= (layer0_outputs(2758)) xor (layer0_outputs(3126));
    outputs(6991) <= not((layer0_outputs(3127)) or (layer0_outputs(133)));
    outputs(6992) <= layer0_outputs(1043);
    outputs(6993) <= '0';
    outputs(6994) <= layer0_outputs(2579);
    outputs(6995) <= not((layer0_outputs(5413)) xor (layer0_outputs(871)));
    outputs(6996) <= (layer0_outputs(2170)) and not (layer0_outputs(7384));
    outputs(6997) <= not(layer0_outputs(880));
    outputs(6998) <= not(layer0_outputs(2392));
    outputs(6999) <= layer0_outputs(2012);
    outputs(7000) <= layer0_outputs(5896);
    outputs(7001) <= (layer0_outputs(2857)) and not (layer0_outputs(6191));
    outputs(7002) <= not(layer0_outputs(5629));
    outputs(7003) <= (layer0_outputs(1526)) xor (layer0_outputs(4697));
    outputs(7004) <= not((layer0_outputs(354)) or (layer0_outputs(1049)));
    outputs(7005) <= (layer0_outputs(5481)) and not (layer0_outputs(5823));
    outputs(7006) <= not(layer0_outputs(4521));
    outputs(7007) <= not(layer0_outputs(7237));
    outputs(7008) <= (layer0_outputs(4079)) and not (layer0_outputs(0));
    outputs(7009) <= not(layer0_outputs(2157));
    outputs(7010) <= (layer0_outputs(7452)) and (layer0_outputs(6575));
    outputs(7011) <= not(layer0_outputs(1964));
    outputs(7012) <= layer0_outputs(3588);
    outputs(7013) <= not(layer0_outputs(7201)) or (layer0_outputs(7626));
    outputs(7014) <= not((layer0_outputs(2278)) xor (layer0_outputs(3318)));
    outputs(7015) <= not(layer0_outputs(3465));
    outputs(7016) <= not((layer0_outputs(4599)) or (layer0_outputs(6287)));
    outputs(7017) <= not(layer0_outputs(2533));
    outputs(7018) <= layer0_outputs(134);
    outputs(7019) <= (layer0_outputs(2407)) xor (layer0_outputs(478));
    outputs(7020) <= not(layer0_outputs(3770));
    outputs(7021) <= (layer0_outputs(3267)) xor (layer0_outputs(1526));
    outputs(7022) <= (layer0_outputs(2209)) and (layer0_outputs(4249));
    outputs(7023) <= not(layer0_outputs(1349));
    outputs(7024) <= not((layer0_outputs(6953)) or (layer0_outputs(1426)));
    outputs(7025) <= not(layer0_outputs(4393));
    outputs(7026) <= not(layer0_outputs(5371));
    outputs(7027) <= not((layer0_outputs(4804)) xor (layer0_outputs(1233)));
    outputs(7028) <= not((layer0_outputs(5339)) xor (layer0_outputs(4350)));
    outputs(7029) <= not(layer0_outputs(2883));
    outputs(7030) <= (layer0_outputs(5461)) and not (layer0_outputs(5475));
    outputs(7031) <= not(layer0_outputs(745));
    outputs(7032) <= not((layer0_outputs(3378)) xor (layer0_outputs(6666)));
    outputs(7033) <= '1';
    outputs(7034) <= layer0_outputs(6733);
    outputs(7035) <= (layer0_outputs(3964)) and not (layer0_outputs(3771));
    outputs(7036) <= not((layer0_outputs(4105)) or (layer0_outputs(4169)));
    outputs(7037) <= not((layer0_outputs(931)) xor (layer0_outputs(6250)));
    outputs(7038) <= layer0_outputs(2844);
    outputs(7039) <= layer0_outputs(365);
    outputs(7040) <= layer0_outputs(2847);
    outputs(7041) <= not((layer0_outputs(7064)) and (layer0_outputs(5324)));
    outputs(7042) <= not((layer0_outputs(3187)) xor (layer0_outputs(7043)));
    outputs(7043) <= not(layer0_outputs(5283));
    outputs(7044) <= not(layer0_outputs(2884));
    outputs(7045) <= (layer0_outputs(161)) xor (layer0_outputs(7679));
    outputs(7046) <= (layer0_outputs(3162)) and not (layer0_outputs(53));
    outputs(7047) <= not((layer0_outputs(7347)) or (layer0_outputs(6571)));
    outputs(7048) <= layer0_outputs(4416);
    outputs(7049) <= (layer0_outputs(3592)) and not (layer0_outputs(3903));
    outputs(7050) <= layer0_outputs(4277);
    outputs(7051) <= not(layer0_outputs(3373));
    outputs(7052) <= (layer0_outputs(3297)) and not (layer0_outputs(819));
    outputs(7053) <= (layer0_outputs(1892)) or (layer0_outputs(4366));
    outputs(7054) <= '0';
    outputs(7055) <= not(layer0_outputs(5924));
    outputs(7056) <= layer0_outputs(5784);
    outputs(7057) <= not(layer0_outputs(7592));
    outputs(7058) <= (layer0_outputs(1582)) and (layer0_outputs(18));
    outputs(7059) <= not(layer0_outputs(3655));
    outputs(7060) <= not(layer0_outputs(1385));
    outputs(7061) <= (layer0_outputs(1220)) xor (layer0_outputs(6331));
    outputs(7062) <= (layer0_outputs(3948)) xor (layer0_outputs(33));
    outputs(7063) <= not(layer0_outputs(7353));
    outputs(7064) <= not(layer0_outputs(2956));
    outputs(7065) <= not(layer0_outputs(26));
    outputs(7066) <= not(layer0_outputs(556));
    outputs(7067) <= (layer0_outputs(1311)) and not (layer0_outputs(6591));
    outputs(7068) <= (layer0_outputs(1910)) and not (layer0_outputs(652));
    outputs(7069) <= layer0_outputs(6230);
    outputs(7070) <= not((layer0_outputs(7635)) and (layer0_outputs(756)));
    outputs(7071) <= layer0_outputs(973);
    outputs(7072) <= layer0_outputs(2225);
    outputs(7073) <= (layer0_outputs(986)) and not (layer0_outputs(6035));
    outputs(7074) <= not(layer0_outputs(5773));
    outputs(7075) <= (layer0_outputs(6755)) and not (layer0_outputs(3556));
    outputs(7076) <= not(layer0_outputs(6062));
    outputs(7077) <= not(layer0_outputs(1474)) or (layer0_outputs(7567));
    outputs(7078) <= not((layer0_outputs(6328)) or (layer0_outputs(2800)));
    outputs(7079) <= not(layer0_outputs(4216)) or (layer0_outputs(2984));
    outputs(7080) <= (layer0_outputs(6925)) and (layer0_outputs(6673));
    outputs(7081) <= not(layer0_outputs(4349));
    outputs(7082) <= (layer0_outputs(3372)) xor (layer0_outputs(508));
    outputs(7083) <= not((layer0_outputs(7452)) and (layer0_outputs(5829)));
    outputs(7084) <= not((layer0_outputs(7247)) or (layer0_outputs(2697)));
    outputs(7085) <= (layer0_outputs(5150)) and (layer0_outputs(1830));
    outputs(7086) <= layer0_outputs(7402);
    outputs(7087) <= not(layer0_outputs(3558)) or (layer0_outputs(445));
    outputs(7088) <= (layer0_outputs(4275)) and not (layer0_outputs(2659));
    outputs(7089) <= not(layer0_outputs(2653)) or (layer0_outputs(5089));
    outputs(7090) <= (layer0_outputs(6455)) and not (layer0_outputs(5818));
    outputs(7091) <= not(layer0_outputs(7646)) or (layer0_outputs(5500));
    outputs(7092) <= (layer0_outputs(5195)) xor (layer0_outputs(7623));
    outputs(7093) <= layer0_outputs(6782);
    outputs(7094) <= not(layer0_outputs(5779));
    outputs(7095) <= (layer0_outputs(7302)) and (layer0_outputs(2048));
    outputs(7096) <= not((layer0_outputs(6871)) xor (layer0_outputs(115)));
    outputs(7097) <= layer0_outputs(3900);
    outputs(7098) <= layer0_outputs(3261);
    outputs(7099) <= (layer0_outputs(4016)) and not (layer0_outputs(894));
    outputs(7100) <= layer0_outputs(3905);
    outputs(7101) <= layer0_outputs(697);
    outputs(7102) <= layer0_outputs(7612);
    outputs(7103) <= (layer0_outputs(1373)) xor (layer0_outputs(1677));
    outputs(7104) <= layer0_outputs(5966);
    outputs(7105) <= not((layer0_outputs(2354)) xor (layer0_outputs(2866)));
    outputs(7106) <= (layer0_outputs(6909)) xor (layer0_outputs(1983));
    outputs(7107) <= not(layer0_outputs(6487));
    outputs(7108) <= layer0_outputs(5813);
    outputs(7109) <= not((layer0_outputs(2355)) and (layer0_outputs(6639)));
    outputs(7110) <= not((layer0_outputs(4787)) and (layer0_outputs(3026)));
    outputs(7111) <= (layer0_outputs(88)) and not (layer0_outputs(3053));
    outputs(7112) <= (layer0_outputs(7324)) xor (layer0_outputs(2833));
    outputs(7113) <= not(layer0_outputs(3848));
    outputs(7114) <= not(layer0_outputs(6992));
    outputs(7115) <= not((layer0_outputs(4068)) xor (layer0_outputs(3685)));
    outputs(7116) <= (layer0_outputs(2931)) and not (layer0_outputs(1690));
    outputs(7117) <= (layer0_outputs(2811)) and not (layer0_outputs(1145));
    outputs(7118) <= layer0_outputs(1712);
    outputs(7119) <= not(layer0_outputs(654));
    outputs(7120) <= layer0_outputs(2963);
    outputs(7121) <= not((layer0_outputs(2675)) and (layer0_outputs(6765)));
    outputs(7122) <= not(layer0_outputs(3847));
    outputs(7123) <= not((layer0_outputs(6937)) xor (layer0_outputs(1295)));
    outputs(7124) <= layer0_outputs(5332);
    outputs(7125) <= layer0_outputs(4433);
    outputs(7126) <= (layer0_outputs(2638)) and not (layer0_outputs(5832));
    outputs(7127) <= not(layer0_outputs(6990));
    outputs(7128) <= not(layer0_outputs(3166));
    outputs(7129) <= not(layer0_outputs(2884));
    outputs(7130) <= not(layer0_outputs(6329)) or (layer0_outputs(2654));
    outputs(7131) <= not((layer0_outputs(3120)) or (layer0_outputs(3326)));
    outputs(7132) <= (layer0_outputs(321)) or (layer0_outputs(2200));
    outputs(7133) <= not(layer0_outputs(2307)) or (layer0_outputs(135));
    outputs(7134) <= not((layer0_outputs(4125)) or (layer0_outputs(924)));
    outputs(7135) <= not(layer0_outputs(1202));
    outputs(7136) <= not(layer0_outputs(3336));
    outputs(7137) <= layer0_outputs(7392);
    outputs(7138) <= not(layer0_outputs(7342));
    outputs(7139) <= not((layer0_outputs(2867)) xor (layer0_outputs(2830)));
    outputs(7140) <= (layer0_outputs(5939)) and (layer0_outputs(5951));
    outputs(7141) <= not(layer0_outputs(4922));
    outputs(7142) <= not((layer0_outputs(2292)) or (layer0_outputs(4778)));
    outputs(7143) <= (layer0_outputs(262)) xor (layer0_outputs(7555));
    outputs(7144) <= (layer0_outputs(4801)) and (layer0_outputs(2867));
    outputs(7145) <= (layer0_outputs(425)) and not (layer0_outputs(3196));
    outputs(7146) <= layer0_outputs(5003);
    outputs(7147) <= not((layer0_outputs(296)) or (layer0_outputs(2808)));
    outputs(7148) <= not((layer0_outputs(2328)) or (layer0_outputs(6033)));
    outputs(7149) <= (layer0_outputs(1357)) and not (layer0_outputs(3445));
    outputs(7150) <= (layer0_outputs(2015)) and not (layer0_outputs(6862));
    outputs(7151) <= not(layer0_outputs(6062)) or (layer0_outputs(6857));
    outputs(7152) <= (layer0_outputs(4897)) and not (layer0_outputs(1384));
    outputs(7153) <= not(layer0_outputs(1170)) or (layer0_outputs(771));
    outputs(7154) <= not((layer0_outputs(1551)) xor (layer0_outputs(2521)));
    outputs(7155) <= not((layer0_outputs(2342)) xor (layer0_outputs(7429)));
    outputs(7156) <= not(layer0_outputs(3114));
    outputs(7157) <= '0';
    outputs(7158) <= layer0_outputs(2362);
    outputs(7159) <= not(layer0_outputs(5479));
    outputs(7160) <= (layer0_outputs(5544)) and not (layer0_outputs(5668));
    outputs(7161) <= not(layer0_outputs(5312));
    outputs(7162) <= layer0_outputs(85);
    outputs(7163) <= (layer0_outputs(273)) and (layer0_outputs(4928));
    outputs(7164) <= (layer0_outputs(4514)) and not (layer0_outputs(7248));
    outputs(7165) <= layer0_outputs(1818);
    outputs(7166) <= layer0_outputs(6096);
    outputs(7167) <= layer0_outputs(178);
    outputs(7168) <= (layer0_outputs(4458)) and not (layer0_outputs(378));
    outputs(7169) <= not((layer0_outputs(5404)) and (layer0_outputs(615)));
    outputs(7170) <= (layer0_outputs(5019)) and (layer0_outputs(551));
    outputs(7171) <= (layer0_outputs(3258)) xor (layer0_outputs(7221));
    outputs(7172) <= not(layer0_outputs(5715));
    outputs(7173) <= not(layer0_outputs(7493));
    outputs(7174) <= layer0_outputs(795);
    outputs(7175) <= not(layer0_outputs(201));
    outputs(7176) <= not((layer0_outputs(5197)) or (layer0_outputs(6572)));
    outputs(7177) <= not((layer0_outputs(4348)) xor (layer0_outputs(5317)));
    outputs(7178) <= not(layer0_outputs(1324));
    outputs(7179) <= (layer0_outputs(384)) and not (layer0_outputs(2298));
    outputs(7180) <= not(layer0_outputs(4037));
    outputs(7181) <= not((layer0_outputs(922)) or (layer0_outputs(5693)));
    outputs(7182) <= '0';
    outputs(7183) <= (layer0_outputs(935)) xor (layer0_outputs(7160));
    outputs(7184) <= (layer0_outputs(4453)) or (layer0_outputs(6460));
    outputs(7185) <= not(layer0_outputs(2873));
    outputs(7186) <= not(layer0_outputs(5570)) or (layer0_outputs(4220));
    outputs(7187) <= (layer0_outputs(4738)) or (layer0_outputs(4209));
    outputs(7188) <= not((layer0_outputs(4)) or (layer0_outputs(6552)));
    outputs(7189) <= not(layer0_outputs(7602));
    outputs(7190) <= not((layer0_outputs(1024)) xor (layer0_outputs(6958)));
    outputs(7191) <= (layer0_outputs(2304)) xor (layer0_outputs(4378));
    outputs(7192) <= not(layer0_outputs(872));
    outputs(7193) <= not((layer0_outputs(128)) or (layer0_outputs(3772)));
    outputs(7194) <= not((layer0_outputs(4386)) xor (layer0_outputs(4294)));
    outputs(7195) <= layer0_outputs(5200);
    outputs(7196) <= layer0_outputs(126);
    outputs(7197) <= layer0_outputs(2796);
    outputs(7198) <= (layer0_outputs(6344)) xor (layer0_outputs(1989));
    outputs(7199) <= not((layer0_outputs(5511)) xor (layer0_outputs(23)));
    outputs(7200) <= (layer0_outputs(2478)) xor (layer0_outputs(1267));
    outputs(7201) <= not(layer0_outputs(3727));
    outputs(7202) <= (layer0_outputs(6068)) and not (layer0_outputs(3689));
    outputs(7203) <= (layer0_outputs(3563)) and (layer0_outputs(5349));
    outputs(7204) <= (layer0_outputs(4359)) xor (layer0_outputs(1231));
    outputs(7205) <= (layer0_outputs(2033)) and not (layer0_outputs(6126));
    outputs(7206) <= (layer0_outputs(2040)) xor (layer0_outputs(6974));
    outputs(7207) <= not(layer0_outputs(2334));
    outputs(7208) <= (layer0_outputs(3105)) and not (layer0_outputs(512));
    outputs(7209) <= (layer0_outputs(1997)) xor (layer0_outputs(1867));
    outputs(7210) <= layer0_outputs(2915);
    outputs(7211) <= (layer0_outputs(4777)) and not (layer0_outputs(4837));
    outputs(7212) <= not((layer0_outputs(7602)) or (layer0_outputs(2862)));
    outputs(7213) <= not((layer0_outputs(7436)) or (layer0_outputs(769)));
    outputs(7214) <= (layer0_outputs(3874)) or (layer0_outputs(7465));
    outputs(7215) <= not(layer0_outputs(6069));
    outputs(7216) <= layer0_outputs(74);
    outputs(7217) <= not((layer0_outputs(1336)) xor (layer0_outputs(2443)));
    outputs(7218) <= not(layer0_outputs(7657));
    outputs(7219) <= (layer0_outputs(2050)) and not (layer0_outputs(6479));
    outputs(7220) <= not((layer0_outputs(1036)) xor (layer0_outputs(6978)));
    outputs(7221) <= (layer0_outputs(420)) xor (layer0_outputs(1032));
    outputs(7222) <= layer0_outputs(4356);
    outputs(7223) <= layer0_outputs(5893);
    outputs(7224) <= not((layer0_outputs(2946)) or (layer0_outputs(309)));
    outputs(7225) <= layer0_outputs(3360);
    outputs(7226) <= not(layer0_outputs(558));
    outputs(7227) <= layer0_outputs(7325);
    outputs(7228) <= not((layer0_outputs(3820)) xor (layer0_outputs(1226)));
    outputs(7229) <= (layer0_outputs(507)) xor (layer0_outputs(6595));
    outputs(7230) <= (layer0_outputs(1450)) and not (layer0_outputs(4538));
    outputs(7231) <= not((layer0_outputs(4417)) or (layer0_outputs(6834)));
    outputs(7232) <= not(layer0_outputs(6272));
    outputs(7233) <= not(layer0_outputs(3018));
    outputs(7234) <= (layer0_outputs(2454)) xor (layer0_outputs(2466));
    outputs(7235) <= (layer0_outputs(6826)) xor (layer0_outputs(1773));
    outputs(7236) <= not(layer0_outputs(7375));
    outputs(7237) <= not(layer0_outputs(6497)) or (layer0_outputs(2893));
    outputs(7238) <= (layer0_outputs(2503)) and not (layer0_outputs(3854));
    outputs(7239) <= not(layer0_outputs(284));
    outputs(7240) <= (layer0_outputs(2542)) and not (layer0_outputs(1142));
    outputs(7241) <= not((layer0_outputs(6891)) xor (layer0_outputs(4861)));
    outputs(7242) <= not(layer0_outputs(991));
    outputs(7243) <= not(layer0_outputs(2303));
    outputs(7244) <= layer0_outputs(6815);
    outputs(7245) <= not((layer0_outputs(1179)) xor (layer0_outputs(5672)));
    outputs(7246) <= not((layer0_outputs(1684)) or (layer0_outputs(3462)));
    outputs(7247) <= (layer0_outputs(424)) and (layer0_outputs(4285));
    outputs(7248) <= not(layer0_outputs(6205));
    outputs(7249) <= layer0_outputs(2963);
    outputs(7250) <= layer0_outputs(3365);
    outputs(7251) <= not((layer0_outputs(360)) xor (layer0_outputs(4185)));
    outputs(7252) <= not(layer0_outputs(6435));
    outputs(7253) <= not(layer0_outputs(4169));
    outputs(7254) <= (layer0_outputs(4055)) xor (layer0_outputs(1241));
    outputs(7255) <= (layer0_outputs(7311)) xor (layer0_outputs(6846));
    outputs(7256) <= not((layer0_outputs(2366)) xor (layer0_outputs(1670)));
    outputs(7257) <= (layer0_outputs(1761)) xor (layer0_outputs(4908));
    outputs(7258) <= (layer0_outputs(6548)) and not (layer0_outputs(6443));
    outputs(7259) <= (layer0_outputs(339)) xor (layer0_outputs(1438));
    outputs(7260) <= (layer0_outputs(4958)) xor (layer0_outputs(443));
    outputs(7261) <= not((layer0_outputs(132)) or (layer0_outputs(6414)));
    outputs(7262) <= not((layer0_outputs(5174)) xor (layer0_outputs(4661)));
    outputs(7263) <= (layer0_outputs(5394)) and not (layer0_outputs(4783));
    outputs(7264) <= (layer0_outputs(190)) and (layer0_outputs(2287));
    outputs(7265) <= not(layer0_outputs(1202)) or (layer0_outputs(2011));
    outputs(7266) <= (layer0_outputs(6023)) and (layer0_outputs(3426));
    outputs(7267) <= layer0_outputs(162);
    outputs(7268) <= not(layer0_outputs(2828)) or (layer0_outputs(6264));
    outputs(7269) <= layer0_outputs(3971);
    outputs(7270) <= not(layer0_outputs(81));
    outputs(7271) <= not((layer0_outputs(2404)) or (layer0_outputs(5768)));
    outputs(7272) <= not(layer0_outputs(1719)) or (layer0_outputs(1560));
    outputs(7273) <= layer0_outputs(2275);
    outputs(7274) <= (layer0_outputs(3247)) and not (layer0_outputs(3780));
    outputs(7275) <= layer0_outputs(1611);
    outputs(7276) <= layer0_outputs(3732);
    outputs(7277) <= (layer0_outputs(7319)) and not (layer0_outputs(4154));
    outputs(7278) <= not(layer0_outputs(2258)) or (layer0_outputs(6083));
    outputs(7279) <= (layer0_outputs(3389)) and (layer0_outputs(1901));
    outputs(7280) <= not(layer0_outputs(1913)) or (layer0_outputs(3724));
    outputs(7281) <= layer0_outputs(3414);
    outputs(7282) <= not((layer0_outputs(815)) xor (layer0_outputs(3478)));
    outputs(7283) <= layer0_outputs(6523);
    outputs(7284) <= not(layer0_outputs(1842));
    outputs(7285) <= not(layer0_outputs(6069));
    outputs(7286) <= layer0_outputs(1031);
    outputs(7287) <= layer0_outputs(4636);
    outputs(7288) <= (layer0_outputs(5435)) and (layer0_outputs(4382));
    outputs(7289) <= '0';
    outputs(7290) <= not(layer0_outputs(2203));
    outputs(7291) <= not((layer0_outputs(1669)) xor (layer0_outputs(7280)));
    outputs(7292) <= not((layer0_outputs(2862)) or (layer0_outputs(4899)));
    outputs(7293) <= not(layer0_outputs(6265)) or (layer0_outputs(6294));
    outputs(7294) <= not(layer0_outputs(5124));
    outputs(7295) <= not(layer0_outputs(3097)) or (layer0_outputs(5161));
    outputs(7296) <= (layer0_outputs(4299)) and (layer0_outputs(2351));
    outputs(7297) <= (layer0_outputs(3891)) and not (layer0_outputs(6423));
    outputs(7298) <= (layer0_outputs(6038)) and not (layer0_outputs(2810));
    outputs(7299) <= not((layer0_outputs(1671)) or (layer0_outputs(5094)));
    outputs(7300) <= not((layer0_outputs(6205)) or (layer0_outputs(2845)));
    outputs(7301) <= layer0_outputs(6314);
    outputs(7302) <= layer0_outputs(539);
    outputs(7303) <= not(layer0_outputs(4228));
    outputs(7304) <= not((layer0_outputs(3628)) xor (layer0_outputs(4375)));
    outputs(7305) <= layer0_outputs(3483);
    outputs(7306) <= (layer0_outputs(1490)) or (layer0_outputs(470));
    outputs(7307) <= (layer0_outputs(5989)) and not (layer0_outputs(1609));
    outputs(7308) <= (layer0_outputs(2421)) and not (layer0_outputs(500));
    outputs(7309) <= (layer0_outputs(2777)) xor (layer0_outputs(3710));
    outputs(7310) <= (layer0_outputs(7446)) and (layer0_outputs(4855));
    outputs(7311) <= not((layer0_outputs(6497)) or (layer0_outputs(2568)));
    outputs(7312) <= not(layer0_outputs(1549));
    outputs(7313) <= (layer0_outputs(5707)) and not (layer0_outputs(56));
    outputs(7314) <= (layer0_outputs(7258)) and not (layer0_outputs(890));
    outputs(7315) <= not(layer0_outputs(1961));
    outputs(7316) <= layer0_outputs(5753);
    outputs(7317) <= not(layer0_outputs(2157));
    outputs(7318) <= not((layer0_outputs(3958)) or (layer0_outputs(6829)));
    outputs(7319) <= not((layer0_outputs(3629)) xor (layer0_outputs(5571)));
    outputs(7320) <= layer0_outputs(1280);
    outputs(7321) <= (layer0_outputs(3881)) xor (layer0_outputs(2343));
    outputs(7322) <= not((layer0_outputs(2126)) and (layer0_outputs(2734)));
    outputs(7323) <= layer0_outputs(1520);
    outputs(7324) <= layer0_outputs(5993);
    outputs(7325) <= not(layer0_outputs(7244));
    outputs(7326) <= (layer0_outputs(6713)) or (layer0_outputs(6219));
    outputs(7327) <= layer0_outputs(7420);
    outputs(7328) <= layer0_outputs(5931);
    outputs(7329) <= (layer0_outputs(4699)) and (layer0_outputs(905));
    outputs(7330) <= (layer0_outputs(604)) xor (layer0_outputs(6323));
    outputs(7331) <= (layer0_outputs(3122)) and not (layer0_outputs(5879));
    outputs(7332) <= layer0_outputs(1058);
    outputs(7333) <= (layer0_outputs(2877)) and not (layer0_outputs(1123));
    outputs(7334) <= (layer0_outputs(2494)) and not (layer0_outputs(1695));
    outputs(7335) <= not(layer0_outputs(7485)) or (layer0_outputs(4436));
    outputs(7336) <= not((layer0_outputs(4488)) xor (layer0_outputs(5196)));
    outputs(7337) <= not(layer0_outputs(6036));
    outputs(7338) <= not((layer0_outputs(7639)) xor (layer0_outputs(2395)));
    outputs(7339) <= (layer0_outputs(4017)) and not (layer0_outputs(5296));
    outputs(7340) <= not(layer0_outputs(1781));
    outputs(7341) <= not(layer0_outputs(153));
    outputs(7342) <= (layer0_outputs(1245)) xor (layer0_outputs(2147));
    outputs(7343) <= not(layer0_outputs(7440)) or (layer0_outputs(1339));
    outputs(7344) <= not((layer0_outputs(2373)) or (layer0_outputs(6457)));
    outputs(7345) <= layer0_outputs(1313);
    outputs(7346) <= layer0_outputs(363);
    outputs(7347) <= not(layer0_outputs(1681));
    outputs(7348) <= (layer0_outputs(6863)) and (layer0_outputs(7195));
    outputs(7349) <= not((layer0_outputs(6011)) or (layer0_outputs(5172)));
    outputs(7350) <= (layer0_outputs(4655)) xor (layer0_outputs(5887));
    outputs(7351) <= (layer0_outputs(5954)) xor (layer0_outputs(5529));
    outputs(7352) <= (layer0_outputs(3645)) and not (layer0_outputs(4210));
    outputs(7353) <= not((layer0_outputs(6149)) or (layer0_outputs(1485)));
    outputs(7354) <= (layer0_outputs(1583)) and (layer0_outputs(6088));
    outputs(7355) <= (layer0_outputs(2427)) and not (layer0_outputs(269));
    outputs(7356) <= not((layer0_outputs(6354)) or (layer0_outputs(1636)));
    outputs(7357) <= layer0_outputs(4834);
    outputs(7358) <= not((layer0_outputs(1363)) or (layer0_outputs(3386)));
    outputs(7359) <= (layer0_outputs(1036)) and (layer0_outputs(3550));
    outputs(7360) <= (layer0_outputs(3476)) and (layer0_outputs(3389));
    outputs(7361) <= (layer0_outputs(7434)) and not (layer0_outputs(5846));
    outputs(7362) <= (layer0_outputs(6222)) and not (layer0_outputs(4380));
    outputs(7363) <= (layer0_outputs(3899)) and not (layer0_outputs(6215));
    outputs(7364) <= not(layer0_outputs(833));
    outputs(7365) <= (layer0_outputs(3560)) and (layer0_outputs(8));
    outputs(7366) <= (layer0_outputs(6493)) xor (layer0_outputs(4657));
    outputs(7367) <= layer0_outputs(4678);
    outputs(7368) <= not(layer0_outputs(1229));
    outputs(7369) <= not((layer0_outputs(7118)) xor (layer0_outputs(6679)));
    outputs(7370) <= not(layer0_outputs(2004));
    outputs(7371) <= layer0_outputs(5231);
    outputs(7372) <= (layer0_outputs(4434)) xor (layer0_outputs(2344));
    outputs(7373) <= not(layer0_outputs(6193)) or (layer0_outputs(1139));
    outputs(7374) <= layer0_outputs(1911);
    outputs(7375) <= layer0_outputs(5029);
    outputs(7376) <= not(layer0_outputs(2699));
    outputs(7377) <= (layer0_outputs(2840)) and not (layer0_outputs(4295));
    outputs(7378) <= (layer0_outputs(7668)) xor (layer0_outputs(7500));
    outputs(7379) <= layer0_outputs(2196);
    outputs(7380) <= (layer0_outputs(2966)) and (layer0_outputs(6777));
    outputs(7381) <= layer0_outputs(3460);
    outputs(7382) <= not((layer0_outputs(2467)) xor (layer0_outputs(1028)));
    outputs(7383) <= not(layer0_outputs(250));
    outputs(7384) <= not(layer0_outputs(3067));
    outputs(7385) <= (layer0_outputs(6984)) and not (layer0_outputs(1115));
    outputs(7386) <= not((layer0_outputs(7028)) xor (layer0_outputs(3860)));
    outputs(7387) <= (layer0_outputs(2608)) or (layer0_outputs(2246));
    outputs(7388) <= (layer0_outputs(1484)) and not (layer0_outputs(4383));
    outputs(7389) <= (layer0_outputs(3676)) and (layer0_outputs(6530));
    outputs(7390) <= not(layer0_outputs(2233));
    outputs(7391) <= (layer0_outputs(6595)) and not (layer0_outputs(3644));
    outputs(7392) <= not((layer0_outputs(2939)) xor (layer0_outputs(1303)));
    outputs(7393) <= not(layer0_outputs(6317));
    outputs(7394) <= layer0_outputs(5795);
    outputs(7395) <= not(layer0_outputs(5297));
    outputs(7396) <= (layer0_outputs(6998)) xor (layer0_outputs(3116));
    outputs(7397) <= (layer0_outputs(7086)) and (layer0_outputs(3135));
    outputs(7398) <= not(layer0_outputs(504));
    outputs(7399) <= layer0_outputs(6769);
    outputs(7400) <= not(layer0_outputs(6206));
    outputs(7401) <= layer0_outputs(3557);
    outputs(7402) <= (layer0_outputs(3387)) and (layer0_outputs(3352));
    outputs(7403) <= (layer0_outputs(4668)) and not (layer0_outputs(3520));
    outputs(7404) <= (layer0_outputs(642)) xor (layer0_outputs(6797));
    outputs(7405) <= layer0_outputs(3353);
    outputs(7406) <= not(layer0_outputs(2771));
    outputs(7407) <= (layer0_outputs(1687)) and (layer0_outputs(1039));
    outputs(7408) <= not((layer0_outputs(4848)) or (layer0_outputs(1106)));
    outputs(7409) <= not(layer0_outputs(7007)) or (layer0_outputs(6925));
    outputs(7410) <= (layer0_outputs(4440)) and not (layer0_outputs(336));
    outputs(7411) <= layer0_outputs(3475);
    outputs(7412) <= not(layer0_outputs(2289)) or (layer0_outputs(4130));
    outputs(7413) <= not((layer0_outputs(526)) xor (layer0_outputs(5932)));
    outputs(7414) <= not(layer0_outputs(4136));
    outputs(7415) <= (layer0_outputs(1310)) xor (layer0_outputs(3860));
    outputs(7416) <= layer0_outputs(2935);
    outputs(7417) <= not(layer0_outputs(1495));
    outputs(7418) <= layer0_outputs(694);
    outputs(7419) <= layer0_outputs(7155);
    outputs(7420) <= not(layer0_outputs(7044));
    outputs(7421) <= not(layer0_outputs(7559));
    outputs(7422) <= not((layer0_outputs(389)) xor (layer0_outputs(2778)));
    outputs(7423) <= layer0_outputs(5804);
    outputs(7424) <= (layer0_outputs(5016)) and (layer0_outputs(4072));
    outputs(7425) <= not(layer0_outputs(2926));
    outputs(7426) <= not(layer0_outputs(955));
    outputs(7427) <= not((layer0_outputs(2053)) and (layer0_outputs(1585)));
    outputs(7428) <= layer0_outputs(7406);
    outputs(7429) <= not(layer0_outputs(4853)) or (layer0_outputs(5558));
    outputs(7430) <= not(layer0_outputs(7484));
    outputs(7431) <= not((layer0_outputs(1942)) xor (layer0_outputs(350)));
    outputs(7432) <= not(layer0_outputs(4963));
    outputs(7433) <= (layer0_outputs(572)) xor (layer0_outputs(6010));
    outputs(7434) <= not(layer0_outputs(1825));
    outputs(7435) <= layer0_outputs(3837);
    outputs(7436) <= '0';
    outputs(7437) <= layer0_outputs(2618);
    outputs(7438) <= layer0_outputs(7194);
    outputs(7439) <= not(layer0_outputs(656));
    outputs(7440) <= layer0_outputs(5806);
    outputs(7441) <= (layer0_outputs(2998)) and (layer0_outputs(5871));
    outputs(7442) <= not((layer0_outputs(7219)) or (layer0_outputs(121)));
    outputs(7443) <= (layer0_outputs(7383)) and not (layer0_outputs(1157));
    outputs(7444) <= (layer0_outputs(381)) and not (layer0_outputs(6827));
    outputs(7445) <= not((layer0_outputs(4333)) and (layer0_outputs(5053)));
    outputs(7446) <= (layer0_outputs(7214)) xor (layer0_outputs(1261));
    outputs(7447) <= not(layer0_outputs(2118));
    outputs(7448) <= layer0_outputs(1367);
    outputs(7449) <= (layer0_outputs(4478)) xor (layer0_outputs(5658));
    outputs(7450) <= (layer0_outputs(5141)) and not (layer0_outputs(7610));
    outputs(7451) <= (layer0_outputs(7585)) and (layer0_outputs(896));
    outputs(7452) <= not(layer0_outputs(4127));
    outputs(7453) <= not(layer0_outputs(4783));
    outputs(7454) <= (layer0_outputs(1089)) or (layer0_outputs(6801));
    outputs(7455) <= (layer0_outputs(6602)) and (layer0_outputs(3888));
    outputs(7456) <= not(layer0_outputs(2447));
    outputs(7457) <= not((layer0_outputs(2295)) or (layer0_outputs(3683)));
    outputs(7458) <= layer0_outputs(753);
    outputs(7459) <= not(layer0_outputs(7109));
    outputs(7460) <= layer0_outputs(1447);
    outputs(7461) <= (layer0_outputs(118)) and not (layer0_outputs(3275));
    outputs(7462) <= layer0_outputs(5686);
    outputs(7463) <= (layer0_outputs(249)) and not (layer0_outputs(403));
    outputs(7464) <= not((layer0_outputs(5400)) xor (layer0_outputs(4093)));
    outputs(7465) <= layer0_outputs(6858);
    outputs(7466) <= (layer0_outputs(4422)) and not (layer0_outputs(7629));
    outputs(7467) <= not(layer0_outputs(6116)) or (layer0_outputs(7558));
    outputs(7468) <= (layer0_outputs(4622)) and not (layer0_outputs(2558));
    outputs(7469) <= not((layer0_outputs(3230)) or (layer0_outputs(4492)));
    outputs(7470) <= (layer0_outputs(2975)) and not (layer0_outputs(2692));
    outputs(7471) <= (layer0_outputs(3397)) and not (layer0_outputs(3015));
    outputs(7472) <= (layer0_outputs(171)) xor (layer0_outputs(1544));
    outputs(7473) <= not(layer0_outputs(1364));
    outputs(7474) <= (layer0_outputs(4498)) xor (layer0_outputs(4256));
    outputs(7475) <= not((layer0_outputs(6295)) xor (layer0_outputs(3540)));
    outputs(7476) <= not(layer0_outputs(5388)) or (layer0_outputs(1513));
    outputs(7477) <= layer0_outputs(1328);
    outputs(7478) <= layer0_outputs(3548);
    outputs(7479) <= (layer0_outputs(6654)) and not (layer0_outputs(3117));
    outputs(7480) <= (layer0_outputs(7530)) xor (layer0_outputs(1291));
    outputs(7481) <= not((layer0_outputs(5179)) or (layer0_outputs(5961)));
    outputs(7482) <= not((layer0_outputs(1565)) or (layer0_outputs(1012)));
    outputs(7483) <= (layer0_outputs(544)) and not (layer0_outputs(5043));
    outputs(7484) <= (layer0_outputs(4381)) xor (layer0_outputs(1501));
    outputs(7485) <= layer0_outputs(6179);
    outputs(7486) <= not((layer0_outputs(6568)) xor (layer0_outputs(7102)));
    outputs(7487) <= not(layer0_outputs(4276)) or (layer0_outputs(1228));
    outputs(7488) <= not((layer0_outputs(7621)) or (layer0_outputs(3565)));
    outputs(7489) <= layer0_outputs(2054);
    outputs(7490) <= layer0_outputs(4694);
    outputs(7491) <= not((layer0_outputs(1123)) or (layer0_outputs(5507)));
    outputs(7492) <= not(layer0_outputs(7552));
    outputs(7493) <= layer0_outputs(3185);
    outputs(7494) <= (layer0_outputs(4317)) and not (layer0_outputs(1416));
    outputs(7495) <= (layer0_outputs(6018)) and not (layer0_outputs(5402));
    outputs(7496) <= (layer0_outputs(2133)) and not (layer0_outputs(4986));
    outputs(7497) <= (layer0_outputs(898)) xor (layer0_outputs(1683));
    outputs(7498) <= layer0_outputs(5576);
    outputs(7499) <= (layer0_outputs(2070)) and (layer0_outputs(5962));
    outputs(7500) <= (layer0_outputs(4587)) xor (layer0_outputs(1765));
    outputs(7501) <= (layer0_outputs(2196)) and not (layer0_outputs(1650));
    outputs(7502) <= not((layer0_outputs(7487)) xor (layer0_outputs(3909)));
    outputs(7503) <= not(layer0_outputs(6210)) or (layer0_outputs(1212));
    outputs(7504) <= not(layer0_outputs(989));
    outputs(7505) <= layer0_outputs(1769);
    outputs(7506) <= not(layer0_outputs(2248)) or (layer0_outputs(4874));
    outputs(7507) <= not((layer0_outputs(527)) or (layer0_outputs(746)));
    outputs(7508) <= not((layer0_outputs(6910)) xor (layer0_outputs(4150)));
    outputs(7509) <= (layer0_outputs(2904)) and (layer0_outputs(2317));
    outputs(7510) <= not(layer0_outputs(3317));
    outputs(7511) <= layer0_outputs(3714);
    outputs(7512) <= not(layer0_outputs(4625));
    outputs(7513) <= not((layer0_outputs(4426)) xor (layer0_outputs(3710)));
    outputs(7514) <= (layer0_outputs(793)) xor (layer0_outputs(5561));
    outputs(7515) <= not((layer0_outputs(2583)) or (layer0_outputs(2330)));
    outputs(7516) <= not(layer0_outputs(2836));
    outputs(7517) <= layer0_outputs(4330);
    outputs(7518) <= not((layer0_outputs(2293)) xor (layer0_outputs(6465)));
    outputs(7519) <= (layer0_outputs(3335)) xor (layer0_outputs(4670));
    outputs(7520) <= not((layer0_outputs(4969)) xor (layer0_outputs(6084)));
    outputs(7521) <= (layer0_outputs(18)) and not (layer0_outputs(4233));
    outputs(7522) <= layer0_outputs(167);
    outputs(7523) <= (layer0_outputs(5653)) and (layer0_outputs(5794));
    outputs(7524) <= layer0_outputs(1288);
    outputs(7525) <= not((layer0_outputs(6658)) and (layer0_outputs(3324)));
    outputs(7526) <= not(layer0_outputs(5728));
    outputs(7527) <= (layer0_outputs(3978)) and (layer0_outputs(5070));
    outputs(7528) <= (layer0_outputs(5865)) and not (layer0_outputs(5569));
    outputs(7529) <= (layer0_outputs(3382)) and (layer0_outputs(265));
    outputs(7530) <= (layer0_outputs(1668)) and not (layer0_outputs(761));
    outputs(7531) <= (layer0_outputs(4529)) and not (layer0_outputs(5897));
    outputs(7532) <= not((layer0_outputs(2455)) or (layer0_outputs(93)));
    outputs(7533) <= not(layer0_outputs(4117));
    outputs(7534) <= not((layer0_outputs(1680)) xor (layer0_outputs(1632)));
    outputs(7535) <= (layer0_outputs(4659)) and not (layer0_outputs(753));
    outputs(7536) <= not((layer0_outputs(944)) or (layer0_outputs(3220)));
    outputs(7537) <= layer0_outputs(4586);
    outputs(7538) <= (layer0_outputs(3598)) and not (layer0_outputs(486));
    outputs(7539) <= layer0_outputs(3350);
    outputs(7540) <= layer0_outputs(5373);
    outputs(7541) <= '0';
    outputs(7542) <= (layer0_outputs(4690)) and not (layer0_outputs(1741));
    outputs(7543) <= not((layer0_outputs(3614)) or (layer0_outputs(6416)));
    outputs(7544) <= not(layer0_outputs(6834));
    outputs(7545) <= (layer0_outputs(6901)) and (layer0_outputs(767));
    outputs(7546) <= not((layer0_outputs(2127)) xor (layer0_outputs(4895)));
    outputs(7547) <= not(layer0_outputs(7154));
    outputs(7548) <= not((layer0_outputs(1041)) or (layer0_outputs(5169)));
    outputs(7549) <= (layer0_outputs(326)) and not (layer0_outputs(6989));
    outputs(7550) <= (layer0_outputs(4308)) and not (layer0_outputs(4343));
    outputs(7551) <= not(layer0_outputs(3005));
    outputs(7552) <= (layer0_outputs(487)) and not (layer0_outputs(6752));
    outputs(7553) <= (layer0_outputs(2748)) and (layer0_outputs(6016));
    outputs(7554) <= layer0_outputs(4328);
    outputs(7555) <= (layer0_outputs(2081)) and not (layer0_outputs(3033));
    outputs(7556) <= (layer0_outputs(147)) xor (layer0_outputs(5024));
    outputs(7557) <= layer0_outputs(1346);
    outputs(7558) <= (layer0_outputs(4059)) xor (layer0_outputs(166));
    outputs(7559) <= not(layer0_outputs(6983));
    outputs(7560) <= not(layer0_outputs(1677));
    outputs(7561) <= (layer0_outputs(4662)) and not (layer0_outputs(6550));
    outputs(7562) <= not((layer0_outputs(4517)) and (layer0_outputs(2674)));
    outputs(7563) <= (layer0_outputs(3676)) and (layer0_outputs(3630));
    outputs(7564) <= layer0_outputs(6080);
    outputs(7565) <= (layer0_outputs(1610)) xor (layer0_outputs(2648));
    outputs(7566) <= not(layer0_outputs(3361));
    outputs(7567) <= not((layer0_outputs(5582)) xor (layer0_outputs(3092)));
    outputs(7568) <= not(layer0_outputs(1654));
    outputs(7569) <= not((layer0_outputs(5900)) and (layer0_outputs(6670)));
    outputs(7570) <= (layer0_outputs(2575)) or (layer0_outputs(948));
    outputs(7571) <= not(layer0_outputs(468));
    outputs(7572) <= (layer0_outputs(505)) xor (layer0_outputs(6606));
    outputs(7573) <= layer0_outputs(3422);
    outputs(7574) <= not(layer0_outputs(5092));
    outputs(7575) <= not((layer0_outputs(2250)) and (layer0_outputs(680)));
    outputs(7576) <= (layer0_outputs(4548)) and not (layer0_outputs(4053));
    outputs(7577) <= layer0_outputs(4447);
    outputs(7578) <= layer0_outputs(4070);
    outputs(7579) <= not(layer0_outputs(6780));
    outputs(7580) <= not((layer0_outputs(2262)) and (layer0_outputs(81)));
    outputs(7581) <= (layer0_outputs(1600)) and not (layer0_outputs(7285));
    outputs(7582) <= (layer0_outputs(1972)) and (layer0_outputs(2088));
    outputs(7583) <= not(layer0_outputs(4280));
    outputs(7584) <= not(layer0_outputs(5241));
    outputs(7585) <= not(layer0_outputs(3337));
    outputs(7586) <= (layer0_outputs(4029)) and not (layer0_outputs(770));
    outputs(7587) <= not((layer0_outputs(4752)) xor (layer0_outputs(4673)));
    outputs(7588) <= not((layer0_outputs(7622)) xor (layer0_outputs(7180)));
    outputs(7589) <= (layer0_outputs(5051)) and (layer0_outputs(5784));
    outputs(7590) <= not((layer0_outputs(2094)) xor (layer0_outputs(5138)));
    outputs(7591) <= '1';
    outputs(7592) <= layer0_outputs(1818);
    outputs(7593) <= not(layer0_outputs(3813));
    outputs(7594) <= not(layer0_outputs(149));
    outputs(7595) <= (layer0_outputs(3893)) and (layer0_outputs(4942));
    outputs(7596) <= layer0_outputs(2275);
    outputs(7597) <= not(layer0_outputs(2272));
    outputs(7598) <= not((layer0_outputs(5006)) xor (layer0_outputs(4226)));
    outputs(7599) <= not(layer0_outputs(2721));
    outputs(7600) <= not(layer0_outputs(4934));
    outputs(7601) <= not((layer0_outputs(179)) xor (layer0_outputs(2820)));
    outputs(7602) <= not(layer0_outputs(270));
    outputs(7603) <= layer0_outputs(4038);
    outputs(7604) <= not(layer0_outputs(1563));
    outputs(7605) <= layer0_outputs(539);
    outputs(7606) <= (layer0_outputs(740)) and not (layer0_outputs(4908));
    outputs(7607) <= not(layer0_outputs(7607));
    outputs(7608) <= not((layer0_outputs(4029)) xor (layer0_outputs(6747)));
    outputs(7609) <= layer0_outputs(3238);
    outputs(7610) <= layer0_outputs(2636);
    outputs(7611) <= not((layer0_outputs(1454)) and (layer0_outputs(6154)));
    outputs(7612) <= (layer0_outputs(5042)) and (layer0_outputs(4968));
    outputs(7613) <= not((layer0_outputs(5077)) xor (layer0_outputs(5687)));
    outputs(7614) <= (layer0_outputs(344)) or (layer0_outputs(3820));
    outputs(7615) <= (layer0_outputs(7183)) and not (layer0_outputs(6938));
    outputs(7616) <= not(layer0_outputs(7647)) or (layer0_outputs(6139));
    outputs(7617) <= (layer0_outputs(4725)) xor (layer0_outputs(2755));
    outputs(7618) <= not(layer0_outputs(3167));
    outputs(7619) <= layer0_outputs(1562);
    outputs(7620) <= layer0_outputs(1127);
    outputs(7621) <= (layer0_outputs(6019)) xor (layer0_outputs(2596));
    outputs(7622) <= not((layer0_outputs(6551)) and (layer0_outputs(5357)));
    outputs(7623) <= not((layer0_outputs(2288)) or (layer0_outputs(2629)));
    outputs(7624) <= (layer0_outputs(2745)) xor (layer0_outputs(3191));
    outputs(7625) <= (layer0_outputs(17)) and not (layer0_outputs(3291));
    outputs(7626) <= not(layer0_outputs(1648));
    outputs(7627) <= (layer0_outputs(1027)) and not (layer0_outputs(2955));
    outputs(7628) <= (layer0_outputs(393)) xor (layer0_outputs(5994));
    outputs(7629) <= (layer0_outputs(2474)) and (layer0_outputs(2074));
    outputs(7630) <= not(layer0_outputs(5788));
    outputs(7631) <= not((layer0_outputs(4111)) or (layer0_outputs(3241)));
    outputs(7632) <= (layer0_outputs(6874)) and (layer0_outputs(1696));
    outputs(7633) <= not((layer0_outputs(6386)) or (layer0_outputs(2785)));
    outputs(7634) <= (layer0_outputs(4662)) and not (layer0_outputs(3114));
    outputs(7635) <= (layer0_outputs(3348)) xor (layer0_outputs(1561));
    outputs(7636) <= layer0_outputs(4562);
    outputs(7637) <= (layer0_outputs(4696)) xor (layer0_outputs(4171));
    outputs(7638) <= not((layer0_outputs(6741)) or (layer0_outputs(5452)));
    outputs(7639) <= (layer0_outputs(1369)) and not (layer0_outputs(3925));
    outputs(7640) <= not(layer0_outputs(1423)) or (layer0_outputs(598));
    outputs(7641) <= layer0_outputs(1704);
    outputs(7642) <= (layer0_outputs(6483)) xor (layer0_outputs(3232));
    outputs(7643) <= not((layer0_outputs(7495)) or (layer0_outputs(6124)));
    outputs(7644) <= (layer0_outputs(4753)) or (layer0_outputs(7628));
    outputs(7645) <= not((layer0_outputs(4750)) xor (layer0_outputs(6662)));
    outputs(7646) <= (layer0_outputs(6883)) and not (layer0_outputs(7495));
    outputs(7647) <= not(layer0_outputs(221));
    outputs(7648) <= layer0_outputs(217);
    outputs(7649) <= (layer0_outputs(3088)) and (layer0_outputs(2621));
    outputs(7650) <= (layer0_outputs(261)) and not (layer0_outputs(3180));
    outputs(7651) <= (layer0_outputs(2795)) and not (layer0_outputs(5291));
    outputs(7652) <= (layer0_outputs(3490)) and not (layer0_outputs(657));
    outputs(7653) <= (layer0_outputs(6468)) and (layer0_outputs(2315));
    outputs(7654) <= not(layer0_outputs(1860));
    outputs(7655) <= (layer0_outputs(6866)) and not (layer0_outputs(5186));
    outputs(7656) <= (layer0_outputs(4729)) and not (layer0_outputs(7407));
    outputs(7657) <= (layer0_outputs(5808)) xor (layer0_outputs(7261));
    outputs(7658) <= (layer0_outputs(3681)) and (layer0_outputs(4937));
    outputs(7659) <= not(layer0_outputs(4962));
    outputs(7660) <= not((layer0_outputs(1962)) xor (layer0_outputs(2313)));
    outputs(7661) <= (layer0_outputs(689)) and not (layer0_outputs(7589));
    outputs(7662) <= layer0_outputs(3954);
    outputs(7663) <= (layer0_outputs(7381)) and (layer0_outputs(1404));
    outputs(7664) <= not(layer0_outputs(3035));
    outputs(7665) <= (layer0_outputs(5146)) and (layer0_outputs(4163));
    outputs(7666) <= not(layer0_outputs(5568));
    outputs(7667) <= layer0_outputs(4387);
    outputs(7668) <= not(layer0_outputs(2304));
    outputs(7669) <= not((layer0_outputs(1523)) or (layer0_outputs(554)));
    outputs(7670) <= layer0_outputs(3577);
    outputs(7671) <= (layer0_outputs(6444)) and not (layer0_outputs(52));
    outputs(7672) <= not(layer0_outputs(2028));
    outputs(7673) <= layer0_outputs(103);
    outputs(7674) <= layer0_outputs(1);
    outputs(7675) <= (layer0_outputs(2104)) and not (layer0_outputs(885));
    outputs(7676) <= (layer0_outputs(714)) and not (layer0_outputs(2948));
    outputs(7677) <= (layer0_outputs(5208)) and (layer0_outputs(5875));
    outputs(7678) <= (layer0_outputs(5068)) or (layer0_outputs(4474));
    outputs(7679) <= (layer0_outputs(5721)) and (layer0_outputs(1655));

end Behavioral;
