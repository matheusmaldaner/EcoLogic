library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(12799 downto 0);
    signal layer1_outputs: std_logic_vector(12799 downto 0);
    signal layer2_outputs: std_logic_vector(12799 downto 0);
    signal layer3_outputs: std_logic_vector(12799 downto 0);
    signal layer4_outputs: std_logic_vector(12799 downto 0);
    signal layer5_outputs: std_logic_vector(12799 downto 0);
    signal layer6_outputs: std_logic_vector(12799 downto 0);

begin
    layer0_outputs(0) <= not b;
    layer0_outputs(1) <= '1';
    layer0_outputs(2) <= b and not a;
    layer0_outputs(3) <= b and not a;
    layer0_outputs(4) <= '0';
    layer0_outputs(5) <= '0';
    layer0_outputs(6) <= not (a or b);
    layer0_outputs(7) <= a xor b;
    layer0_outputs(8) <= a or b;
    layer0_outputs(9) <= not a;
    layer0_outputs(10) <= not b;
    layer0_outputs(11) <= a;
    layer0_outputs(12) <= '0';
    layer0_outputs(13) <= not b or a;
    layer0_outputs(14) <= not a;
    layer0_outputs(15) <= a or b;
    layer0_outputs(16) <= a or b;
    layer0_outputs(17) <= not (a xor b);
    layer0_outputs(18) <= not (a xor b);
    layer0_outputs(19) <= not (a or b);
    layer0_outputs(20) <= a xor b;
    layer0_outputs(21) <= b;
    layer0_outputs(22) <= b and not a;
    layer0_outputs(23) <= not b;
    layer0_outputs(24) <= '0';
    layer0_outputs(25) <= a and not b;
    layer0_outputs(26) <= not a;
    layer0_outputs(27) <= '0';
    layer0_outputs(28) <= not b;
    layer0_outputs(29) <= b;
    layer0_outputs(30) <= '1';
    layer0_outputs(31) <= a;
    layer0_outputs(32) <= a or b;
    layer0_outputs(33) <= not a or b;
    layer0_outputs(34) <= a and b;
    layer0_outputs(35) <= a xor b;
    layer0_outputs(36) <= a xor b;
    layer0_outputs(37) <= a xor b;
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= b and not a;
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= a;
    layer0_outputs(42) <= not (a or b);
    layer0_outputs(43) <= b and not a;
    layer0_outputs(44) <= not b;
    layer0_outputs(45) <= not (a xor b);
    layer0_outputs(46) <= b;
    layer0_outputs(47) <= not b;
    layer0_outputs(48) <= a and not b;
    layer0_outputs(49) <= not (a and b);
    layer0_outputs(50) <= not b;
    layer0_outputs(51) <= a and not b;
    layer0_outputs(52) <= '0';
    layer0_outputs(53) <= not b;
    layer0_outputs(54) <= not (a or b);
    layer0_outputs(55) <= not (a or b);
    layer0_outputs(56) <= b;
    layer0_outputs(57) <= a or b;
    layer0_outputs(58) <= b and not a;
    layer0_outputs(59) <= not b or a;
    layer0_outputs(60) <= a;
    layer0_outputs(61) <= not a or b;
    layer0_outputs(62) <= a;
    layer0_outputs(63) <= b;
    layer0_outputs(64) <= a and b;
    layer0_outputs(65) <= b and not a;
    layer0_outputs(66) <= not b or a;
    layer0_outputs(67) <= a xor b;
    layer0_outputs(68) <= b and not a;
    layer0_outputs(69) <= a and b;
    layer0_outputs(70) <= not (a and b);
    layer0_outputs(71) <= not b or a;
    layer0_outputs(72) <= not a or b;
    layer0_outputs(73) <= not b or a;
    layer0_outputs(74) <= not a or b;
    layer0_outputs(75) <= '1';
    layer0_outputs(76) <= b;
    layer0_outputs(77) <= '1';
    layer0_outputs(78) <= b;
    layer0_outputs(79) <= b and not a;
    layer0_outputs(80) <= a xor b;
    layer0_outputs(81) <= a and not b;
    layer0_outputs(82) <= not a or b;
    layer0_outputs(83) <= not a or b;
    layer0_outputs(84) <= not b or a;
    layer0_outputs(85) <= not a;
    layer0_outputs(86) <= a xor b;
    layer0_outputs(87) <= '0';
    layer0_outputs(88) <= a and b;
    layer0_outputs(89) <= b;
    layer0_outputs(90) <= not a or b;
    layer0_outputs(91) <= not a;
    layer0_outputs(92) <= a and b;
    layer0_outputs(93) <= a and b;
    layer0_outputs(94) <= '0';
    layer0_outputs(95) <= a or b;
    layer0_outputs(96) <= a or b;
    layer0_outputs(97) <= a and not b;
    layer0_outputs(98) <= '1';
    layer0_outputs(99) <= b;
    layer0_outputs(100) <= a and not b;
    layer0_outputs(101) <= not (a or b);
    layer0_outputs(102) <= b;
    layer0_outputs(103) <= a or b;
    layer0_outputs(104) <= not b or a;
    layer0_outputs(105) <= not a or b;
    layer0_outputs(106) <= not (a or b);
    layer0_outputs(107) <= not a or b;
    layer0_outputs(108) <= not (a xor b);
    layer0_outputs(109) <= a or b;
    layer0_outputs(110) <= not b or a;
    layer0_outputs(111) <= not a;
    layer0_outputs(112) <= not (a or b);
    layer0_outputs(113) <= a or b;
    layer0_outputs(114) <= a and not b;
    layer0_outputs(115) <= not (a xor b);
    layer0_outputs(116) <= '1';
    layer0_outputs(117) <= b;
    layer0_outputs(118) <= not (a and b);
    layer0_outputs(119) <= not (a or b);
    layer0_outputs(120) <= a;
    layer0_outputs(121) <= a or b;
    layer0_outputs(122) <= a or b;
    layer0_outputs(123) <= a;
    layer0_outputs(124) <= a or b;
    layer0_outputs(125) <= a and not b;
    layer0_outputs(126) <= a;
    layer0_outputs(127) <= a xor b;
    layer0_outputs(128) <= not b;
    layer0_outputs(129) <= not b;
    layer0_outputs(130) <= '1';
    layer0_outputs(131) <= b and not a;
    layer0_outputs(132) <= a and b;
    layer0_outputs(133) <= a xor b;
    layer0_outputs(134) <= not (a xor b);
    layer0_outputs(135) <= not a or b;
    layer0_outputs(136) <= b;
    layer0_outputs(137) <= a and not b;
    layer0_outputs(138) <= a and b;
    layer0_outputs(139) <= b and not a;
    layer0_outputs(140) <= not a;
    layer0_outputs(141) <= not (a or b);
    layer0_outputs(142) <= b;
    layer0_outputs(143) <= not (a or b);
    layer0_outputs(144) <= a and not b;
    layer0_outputs(145) <= not (a and b);
    layer0_outputs(146) <= b;
    layer0_outputs(147) <= a and not b;
    layer0_outputs(148) <= '1';
    layer0_outputs(149) <= not a;
    layer0_outputs(150) <= not b or a;
    layer0_outputs(151) <= not b or a;
    layer0_outputs(152) <= not b or a;
    layer0_outputs(153) <= not a or b;
    layer0_outputs(154) <= a or b;
    layer0_outputs(155) <= a xor b;
    layer0_outputs(156) <= not (a or b);
    layer0_outputs(157) <= a;
    layer0_outputs(158) <= b;
    layer0_outputs(159) <= b and not a;
    layer0_outputs(160) <= a xor b;
    layer0_outputs(161) <= not (a xor b);
    layer0_outputs(162) <= a;
    layer0_outputs(163) <= a xor b;
    layer0_outputs(164) <= '1';
    layer0_outputs(165) <= b;
    layer0_outputs(166) <= b;
    layer0_outputs(167) <= not (a or b);
    layer0_outputs(168) <= not (a or b);
    layer0_outputs(169) <= not (a or b);
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= not (a and b);
    layer0_outputs(172) <= a and not b;
    layer0_outputs(173) <= a or b;
    layer0_outputs(174) <= not a;
    layer0_outputs(175) <= not (a and b);
    layer0_outputs(176) <= a;
    layer0_outputs(177) <= b;
    layer0_outputs(178) <= a or b;
    layer0_outputs(179) <= b;
    layer0_outputs(180) <= not b or a;
    layer0_outputs(181) <= b;
    layer0_outputs(182) <= '0';
    layer0_outputs(183) <= not (a xor b);
    layer0_outputs(184) <= a or b;
    layer0_outputs(185) <= not (a and b);
    layer0_outputs(186) <= not b or a;
    layer0_outputs(187) <= not a;
    layer0_outputs(188) <= not a;
    layer0_outputs(189) <= a and not b;
    layer0_outputs(190) <= a xor b;
    layer0_outputs(191) <= '0';
    layer0_outputs(192) <= a and not b;
    layer0_outputs(193) <= a;
    layer0_outputs(194) <= a or b;
    layer0_outputs(195) <= '0';
    layer0_outputs(196) <= not b;
    layer0_outputs(197) <= b and not a;
    layer0_outputs(198) <= not b;
    layer0_outputs(199) <= a and not b;
    layer0_outputs(200) <= not b;
    layer0_outputs(201) <= b and not a;
    layer0_outputs(202) <= not (a xor b);
    layer0_outputs(203) <= a or b;
    layer0_outputs(204) <= a;
    layer0_outputs(205) <= not (a xor b);
    layer0_outputs(206) <= a xor b;
    layer0_outputs(207) <= a xor b;
    layer0_outputs(208) <= not (a and b);
    layer0_outputs(209) <= not (a and b);
    layer0_outputs(210) <= b;
    layer0_outputs(211) <= b;
    layer0_outputs(212) <= a and b;
    layer0_outputs(213) <= b;
    layer0_outputs(214) <= b and not a;
    layer0_outputs(215) <= not (a or b);
    layer0_outputs(216) <= a or b;
    layer0_outputs(217) <= not b;
    layer0_outputs(218) <= a or b;
    layer0_outputs(219) <= not a;
    layer0_outputs(220) <= not a;
    layer0_outputs(221) <= '1';
    layer0_outputs(222) <= not (a xor b);
    layer0_outputs(223) <= a xor b;
    layer0_outputs(224) <= not b;
    layer0_outputs(225) <= a or b;
    layer0_outputs(226) <= not (a and b);
    layer0_outputs(227) <= b and not a;
    layer0_outputs(228) <= a and b;
    layer0_outputs(229) <= not a or b;
    layer0_outputs(230) <= not (a or b);
    layer0_outputs(231) <= b and not a;
    layer0_outputs(232) <= not b or a;
    layer0_outputs(233) <= not b;
    layer0_outputs(234) <= not a or b;
    layer0_outputs(235) <= not (a and b);
    layer0_outputs(236) <= a and b;
    layer0_outputs(237) <= not b or a;
    layer0_outputs(238) <= a and not b;
    layer0_outputs(239) <= not a;
    layer0_outputs(240) <= not (a xor b);
    layer0_outputs(241) <= not a or b;
    layer0_outputs(242) <= not a;
    layer0_outputs(243) <= not b or a;
    layer0_outputs(244) <= a and not b;
    layer0_outputs(245) <= b;
    layer0_outputs(246) <= not a;
    layer0_outputs(247) <= not (a xor b);
    layer0_outputs(248) <= a and b;
    layer0_outputs(249) <= a or b;
    layer0_outputs(250) <= not (a or b);
    layer0_outputs(251) <= a or b;
    layer0_outputs(252) <= not b or a;
    layer0_outputs(253) <= a and not b;
    layer0_outputs(254) <= a or b;
    layer0_outputs(255) <= not a;
    layer0_outputs(256) <= not (a xor b);
    layer0_outputs(257) <= not a or b;
    layer0_outputs(258) <= a xor b;
    layer0_outputs(259) <= a xor b;
    layer0_outputs(260) <= not b or a;
    layer0_outputs(261) <= not (a or b);
    layer0_outputs(262) <= a;
    layer0_outputs(263) <= b and not a;
    layer0_outputs(264) <= not (a xor b);
    layer0_outputs(265) <= '0';
    layer0_outputs(266) <= not a;
    layer0_outputs(267) <= '1';
    layer0_outputs(268) <= not b;
    layer0_outputs(269) <= a and not b;
    layer0_outputs(270) <= '1';
    layer0_outputs(271) <= not a;
    layer0_outputs(272) <= a or b;
    layer0_outputs(273) <= not a;
    layer0_outputs(274) <= '1';
    layer0_outputs(275) <= a or b;
    layer0_outputs(276) <= a;
    layer0_outputs(277) <= not b;
    layer0_outputs(278) <= not (a xor b);
    layer0_outputs(279) <= not b or a;
    layer0_outputs(280) <= b;
    layer0_outputs(281) <= not a;
    layer0_outputs(282) <= not b or a;
    layer0_outputs(283) <= not (a xor b);
    layer0_outputs(284) <= not b or a;
    layer0_outputs(285) <= not a or b;
    layer0_outputs(286) <= not a;
    layer0_outputs(287) <= not a;
    layer0_outputs(288) <= a xor b;
    layer0_outputs(289) <= not a;
    layer0_outputs(290) <= '0';
    layer0_outputs(291) <= a;
    layer0_outputs(292) <= not (a xor b);
    layer0_outputs(293) <= not (a xor b);
    layer0_outputs(294) <= b and not a;
    layer0_outputs(295) <= not (a xor b);
    layer0_outputs(296) <= b;
    layer0_outputs(297) <= not b;
    layer0_outputs(298) <= a;
    layer0_outputs(299) <= not (a or b);
    layer0_outputs(300) <= not a;
    layer0_outputs(301) <= b;
    layer0_outputs(302) <= not b;
    layer0_outputs(303) <= b and not a;
    layer0_outputs(304) <= not b;
    layer0_outputs(305) <= a xor b;
    layer0_outputs(306) <= not (a and b);
    layer0_outputs(307) <= not b or a;
    layer0_outputs(308) <= a or b;
    layer0_outputs(309) <= a or b;
    layer0_outputs(310) <= a and b;
    layer0_outputs(311) <= a or b;
    layer0_outputs(312) <= a xor b;
    layer0_outputs(313) <= a and not b;
    layer0_outputs(314) <= not b;
    layer0_outputs(315) <= not b or a;
    layer0_outputs(316) <= a or b;
    layer0_outputs(317) <= '0';
    layer0_outputs(318) <= not (a or b);
    layer0_outputs(319) <= not (a and b);
    layer0_outputs(320) <= b;
    layer0_outputs(321) <= a xor b;
    layer0_outputs(322) <= not (a or b);
    layer0_outputs(323) <= '0';
    layer0_outputs(324) <= not a;
    layer0_outputs(325) <= not (a or b);
    layer0_outputs(326) <= '1';
    layer0_outputs(327) <= b;
    layer0_outputs(328) <= not (a or b);
    layer0_outputs(329) <= not a;
    layer0_outputs(330) <= a;
    layer0_outputs(331) <= b;
    layer0_outputs(332) <= a;
    layer0_outputs(333) <= not (a and b);
    layer0_outputs(334) <= not (a xor b);
    layer0_outputs(335) <= not (a and b);
    layer0_outputs(336) <= b;
    layer0_outputs(337) <= a and b;
    layer0_outputs(338) <= b and not a;
    layer0_outputs(339) <= '1';
    layer0_outputs(340) <= not b or a;
    layer0_outputs(341) <= a or b;
    layer0_outputs(342) <= not b or a;
    layer0_outputs(343) <= not (a xor b);
    layer0_outputs(344) <= '0';
    layer0_outputs(345) <= '0';
    layer0_outputs(346) <= b and not a;
    layer0_outputs(347) <= a xor b;
    layer0_outputs(348) <= b;
    layer0_outputs(349) <= not a or b;
    layer0_outputs(350) <= not b;
    layer0_outputs(351) <= b and not a;
    layer0_outputs(352) <= a and not b;
    layer0_outputs(353) <= a or b;
    layer0_outputs(354) <= '1';
    layer0_outputs(355) <= '1';
    layer0_outputs(356) <= a and not b;
    layer0_outputs(357) <= b;
    layer0_outputs(358) <= a and b;
    layer0_outputs(359) <= not (a and b);
    layer0_outputs(360) <= not (a or b);
    layer0_outputs(361) <= a xor b;
    layer0_outputs(362) <= b and not a;
    layer0_outputs(363) <= not (a and b);
    layer0_outputs(364) <= b;
    layer0_outputs(365) <= not b;
    layer0_outputs(366) <= b and not a;
    layer0_outputs(367) <= a xor b;
    layer0_outputs(368) <= '1';
    layer0_outputs(369) <= b and not a;
    layer0_outputs(370) <= not (a or b);
    layer0_outputs(371) <= a and b;
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= not a;
    layer0_outputs(374) <= a or b;
    layer0_outputs(375) <= not b or a;
    layer0_outputs(376) <= a and not b;
    layer0_outputs(377) <= b;
    layer0_outputs(378) <= not a or b;
    layer0_outputs(379) <= not b;
    layer0_outputs(380) <= not a;
    layer0_outputs(381) <= not a;
    layer0_outputs(382) <= not (a or b);
    layer0_outputs(383) <= not (a or b);
    layer0_outputs(384) <= a and not b;
    layer0_outputs(385) <= b;
    layer0_outputs(386) <= not a;
    layer0_outputs(387) <= '0';
    layer0_outputs(388) <= not (a and b);
    layer0_outputs(389) <= '1';
    layer0_outputs(390) <= a;
    layer0_outputs(391) <= b;
    layer0_outputs(392) <= a or b;
    layer0_outputs(393) <= a and b;
    layer0_outputs(394) <= not a or b;
    layer0_outputs(395) <= not (a xor b);
    layer0_outputs(396) <= b and not a;
    layer0_outputs(397) <= not a;
    layer0_outputs(398) <= not a or b;
    layer0_outputs(399) <= a and b;
    layer0_outputs(400) <= b and not a;
    layer0_outputs(401) <= a and not b;
    layer0_outputs(402) <= a and not b;
    layer0_outputs(403) <= b;
    layer0_outputs(404) <= b;
    layer0_outputs(405) <= not (a and b);
    layer0_outputs(406) <= '1';
    layer0_outputs(407) <= b;
    layer0_outputs(408) <= not (a or b);
    layer0_outputs(409) <= not a;
    layer0_outputs(410) <= not a or b;
    layer0_outputs(411) <= a and not b;
    layer0_outputs(412) <= not b;
    layer0_outputs(413) <= '1';
    layer0_outputs(414) <= a and not b;
    layer0_outputs(415) <= '0';
    layer0_outputs(416) <= b;
    layer0_outputs(417) <= '1';
    layer0_outputs(418) <= a and not b;
    layer0_outputs(419) <= not a;
    layer0_outputs(420) <= b and not a;
    layer0_outputs(421) <= not (a or b);
    layer0_outputs(422) <= b;
    layer0_outputs(423) <= not b or a;
    layer0_outputs(424) <= not b or a;
    layer0_outputs(425) <= not (a or b);
    layer0_outputs(426) <= a or b;
    layer0_outputs(427) <= not a;
    layer0_outputs(428) <= b;
    layer0_outputs(429) <= b and not a;
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= b and not a;
    layer0_outputs(432) <= not (a or b);
    layer0_outputs(433) <= a or b;
    layer0_outputs(434) <= a or b;
    layer0_outputs(435) <= a;
    layer0_outputs(436) <= b;
    layer0_outputs(437) <= a;
    layer0_outputs(438) <= not (a and b);
    layer0_outputs(439) <= b;
    layer0_outputs(440) <= not (a xor b);
    layer0_outputs(441) <= b;
    layer0_outputs(442) <= a or b;
    layer0_outputs(443) <= not (a or b);
    layer0_outputs(444) <= not (a or b);
    layer0_outputs(445) <= not (a or b);
    layer0_outputs(446) <= '0';
    layer0_outputs(447) <= b and not a;
    layer0_outputs(448) <= a or b;
    layer0_outputs(449) <= not b or a;
    layer0_outputs(450) <= not a;
    layer0_outputs(451) <= a;
    layer0_outputs(452) <= a and b;
    layer0_outputs(453) <= not a or b;
    layer0_outputs(454) <= not b;
    layer0_outputs(455) <= a or b;
    layer0_outputs(456) <= a or b;
    layer0_outputs(457) <= a and b;
    layer0_outputs(458) <= not a;
    layer0_outputs(459) <= not b;
    layer0_outputs(460) <= a or b;
    layer0_outputs(461) <= a;
    layer0_outputs(462) <= not (a or b);
    layer0_outputs(463) <= b and not a;
    layer0_outputs(464) <= a;
    layer0_outputs(465) <= not b;
    layer0_outputs(466) <= a xor b;
    layer0_outputs(467) <= not a;
    layer0_outputs(468) <= '1';
    layer0_outputs(469) <= a xor b;
    layer0_outputs(470) <= not (a xor b);
    layer0_outputs(471) <= a;
    layer0_outputs(472) <= not (a xor b);
    layer0_outputs(473) <= '0';
    layer0_outputs(474) <= b and not a;
    layer0_outputs(475) <= not (a or b);
    layer0_outputs(476) <= not a or b;
    layer0_outputs(477) <= not (a or b);
    layer0_outputs(478) <= a;
    layer0_outputs(479) <= not a or b;
    layer0_outputs(480) <= b;
    layer0_outputs(481) <= not (a and b);
    layer0_outputs(482) <= a and not b;
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= b;
    layer0_outputs(485) <= '0';
    layer0_outputs(486) <= not a;
    layer0_outputs(487) <= not b or a;
    layer0_outputs(488) <= not (a or b);
    layer0_outputs(489) <= '1';
    layer0_outputs(490) <= not a or b;
    layer0_outputs(491) <= not (a and b);
    layer0_outputs(492) <= a or b;
    layer0_outputs(493) <= not a;
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= a or b;
    layer0_outputs(496) <= a or b;
    layer0_outputs(497) <= b and not a;
    layer0_outputs(498) <= not b or a;
    layer0_outputs(499) <= not a or b;
    layer0_outputs(500) <= a xor b;
    layer0_outputs(501) <= not (a xor b);
    layer0_outputs(502) <= b;
    layer0_outputs(503) <= a and b;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= not a;
    layer0_outputs(506) <= not (a and b);
    layer0_outputs(507) <= not a or b;
    layer0_outputs(508) <= not (a and b);
    layer0_outputs(509) <= not (a xor b);
    layer0_outputs(510) <= not (a xor b);
    layer0_outputs(511) <= not (a or b);
    layer0_outputs(512) <= not b;
    layer0_outputs(513) <= a xor b;
    layer0_outputs(514) <= not b or a;
    layer0_outputs(515) <= b;
    layer0_outputs(516) <= not a;
    layer0_outputs(517) <= not (a xor b);
    layer0_outputs(518) <= b and not a;
    layer0_outputs(519) <= not (a and b);
    layer0_outputs(520) <= a or b;
    layer0_outputs(521) <= '0';
    layer0_outputs(522) <= not a;
    layer0_outputs(523) <= b and not a;
    layer0_outputs(524) <= b;
    layer0_outputs(525) <= a and not b;
    layer0_outputs(526) <= not (a and b);
    layer0_outputs(527) <= not (a or b);
    layer0_outputs(528) <= not (a and b);
    layer0_outputs(529) <= a xor b;
    layer0_outputs(530) <= a;
    layer0_outputs(531) <= a and not b;
    layer0_outputs(532) <= a and b;
    layer0_outputs(533) <= b and not a;
    layer0_outputs(534) <= not (a xor b);
    layer0_outputs(535) <= a and not b;
    layer0_outputs(536) <= a xor b;
    layer0_outputs(537) <= not b or a;
    layer0_outputs(538) <= not (a or b);
    layer0_outputs(539) <= '0';
    layer0_outputs(540) <= not a;
    layer0_outputs(541) <= '0';
    layer0_outputs(542) <= a and b;
    layer0_outputs(543) <= not a;
    layer0_outputs(544) <= not b;
    layer0_outputs(545) <= not b;
    layer0_outputs(546) <= a;
    layer0_outputs(547) <= not (a or b);
    layer0_outputs(548) <= '1';
    layer0_outputs(549) <= not b;
    layer0_outputs(550) <= not a or b;
    layer0_outputs(551) <= not a;
    layer0_outputs(552) <= a and b;
    layer0_outputs(553) <= not a;
    layer0_outputs(554) <= '1';
    layer0_outputs(555) <= not b;
    layer0_outputs(556) <= not (a or b);
    layer0_outputs(557) <= not b;
    layer0_outputs(558) <= not (a and b);
    layer0_outputs(559) <= a and not b;
    layer0_outputs(560) <= not b;
    layer0_outputs(561) <= not b;
    layer0_outputs(562) <= b;
    layer0_outputs(563) <= a and not b;
    layer0_outputs(564) <= not a or b;
    layer0_outputs(565) <= '0';
    layer0_outputs(566) <= b and not a;
    layer0_outputs(567) <= not b;
    layer0_outputs(568) <= not b or a;
    layer0_outputs(569) <= not a;
    layer0_outputs(570) <= a or b;
    layer0_outputs(571) <= not b;
    layer0_outputs(572) <= b;
    layer0_outputs(573) <= b and not a;
    layer0_outputs(574) <= not b;
    layer0_outputs(575) <= b;
    layer0_outputs(576) <= not b or a;
    layer0_outputs(577) <= not (a or b);
    layer0_outputs(578) <= a xor b;
    layer0_outputs(579) <= not a;
    layer0_outputs(580) <= a xor b;
    layer0_outputs(581) <= not a;
    layer0_outputs(582) <= not a;
    layer0_outputs(583) <= a;
    layer0_outputs(584) <= b and not a;
    layer0_outputs(585) <= not b or a;
    layer0_outputs(586) <= a xor b;
    layer0_outputs(587) <= not a or b;
    layer0_outputs(588) <= not a or b;
    layer0_outputs(589) <= '1';
    layer0_outputs(590) <= not b or a;
    layer0_outputs(591) <= a or b;
    layer0_outputs(592) <= not (a and b);
    layer0_outputs(593) <= a and b;
    layer0_outputs(594) <= a;
    layer0_outputs(595) <= b;
    layer0_outputs(596) <= not a;
    layer0_outputs(597) <= not (a or b);
    layer0_outputs(598) <= b;
    layer0_outputs(599) <= not (a xor b);
    layer0_outputs(600) <= '1';
    layer0_outputs(601) <= a xor b;
    layer0_outputs(602) <= not a or b;
    layer0_outputs(603) <= not b or a;
    layer0_outputs(604) <= a or b;
    layer0_outputs(605) <= not a or b;
    layer0_outputs(606) <= a and b;
    layer0_outputs(607) <= not b or a;
    layer0_outputs(608) <= a or b;
    layer0_outputs(609) <= a xor b;
    layer0_outputs(610) <= a or b;
    layer0_outputs(611) <= not b or a;
    layer0_outputs(612) <= a;
    layer0_outputs(613) <= not a;
    layer0_outputs(614) <= not (a and b);
    layer0_outputs(615) <= not a or b;
    layer0_outputs(616) <= not b or a;
    layer0_outputs(617) <= not (a xor b);
    layer0_outputs(618) <= b;
    layer0_outputs(619) <= not a or b;
    layer0_outputs(620) <= a xor b;
    layer0_outputs(621) <= a or b;
    layer0_outputs(622) <= a xor b;
    layer0_outputs(623) <= b and not a;
    layer0_outputs(624) <= '0';
    layer0_outputs(625) <= a;
    layer0_outputs(626) <= a and b;
    layer0_outputs(627) <= a;
    layer0_outputs(628) <= a or b;
    layer0_outputs(629) <= '1';
    layer0_outputs(630) <= a xor b;
    layer0_outputs(631) <= a or b;
    layer0_outputs(632) <= a and b;
    layer0_outputs(633) <= a;
    layer0_outputs(634) <= a and not b;
    layer0_outputs(635) <= not (a and b);
    layer0_outputs(636) <= not b or a;
    layer0_outputs(637) <= not (a and b);
    layer0_outputs(638) <= not a;
    layer0_outputs(639) <= b and not a;
    layer0_outputs(640) <= not a;
    layer0_outputs(641) <= not a or b;
    layer0_outputs(642) <= '0';
    layer0_outputs(643) <= not (a xor b);
    layer0_outputs(644) <= a or b;
    layer0_outputs(645) <= not a or b;
    layer0_outputs(646) <= not b;
    layer0_outputs(647) <= a or b;
    layer0_outputs(648) <= b and not a;
    layer0_outputs(649) <= not (a xor b);
    layer0_outputs(650) <= not b;
    layer0_outputs(651) <= '1';
    layer0_outputs(652) <= a or b;
    layer0_outputs(653) <= a and b;
    layer0_outputs(654) <= a and b;
    layer0_outputs(655) <= not (a or b);
    layer0_outputs(656) <= '0';
    layer0_outputs(657) <= not (a xor b);
    layer0_outputs(658) <= not (a or b);
    layer0_outputs(659) <= not a;
    layer0_outputs(660) <= a;
    layer0_outputs(661) <= not a;
    layer0_outputs(662) <= not a or b;
    layer0_outputs(663) <= not a or b;
    layer0_outputs(664) <= b;
    layer0_outputs(665) <= '0';
    layer0_outputs(666) <= a;
    layer0_outputs(667) <= a xor b;
    layer0_outputs(668) <= a or b;
    layer0_outputs(669) <= not (a and b);
    layer0_outputs(670) <= not (a and b);
    layer0_outputs(671) <= '0';
    layer0_outputs(672) <= b;
    layer0_outputs(673) <= a or b;
    layer0_outputs(674) <= a and not b;
    layer0_outputs(675) <= not (a and b);
    layer0_outputs(676) <= a and not b;
    layer0_outputs(677) <= not (a or b);
    layer0_outputs(678) <= not (a and b);
    layer0_outputs(679) <= a xor b;
    layer0_outputs(680) <= not (a xor b);
    layer0_outputs(681) <= '0';
    layer0_outputs(682) <= not a or b;
    layer0_outputs(683) <= b;
    layer0_outputs(684) <= not b;
    layer0_outputs(685) <= b;
    layer0_outputs(686) <= not (a xor b);
    layer0_outputs(687) <= '1';
    layer0_outputs(688) <= a;
    layer0_outputs(689) <= a and b;
    layer0_outputs(690) <= not b or a;
    layer0_outputs(691) <= not b or a;
    layer0_outputs(692) <= a or b;
    layer0_outputs(693) <= not a;
    layer0_outputs(694) <= a and b;
    layer0_outputs(695) <= not b or a;
    layer0_outputs(696) <= '1';
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= b and not a;
    layer0_outputs(699) <= not a;
    layer0_outputs(700) <= not a;
    layer0_outputs(701) <= not (a or b);
    layer0_outputs(702) <= not (a and b);
    layer0_outputs(703) <= a and not b;
    layer0_outputs(704) <= '0';
    layer0_outputs(705) <= b and not a;
    layer0_outputs(706) <= not b;
    layer0_outputs(707) <= not a or b;
    layer0_outputs(708) <= not (a or b);
    layer0_outputs(709) <= '0';
    layer0_outputs(710) <= a and not b;
    layer0_outputs(711) <= a and not b;
    layer0_outputs(712) <= not b or a;
    layer0_outputs(713) <= a and not b;
    layer0_outputs(714) <= not (a or b);
    layer0_outputs(715) <= a or b;
    layer0_outputs(716) <= '1';
    layer0_outputs(717) <= not (a or b);
    layer0_outputs(718) <= a and b;
    layer0_outputs(719) <= b;
    layer0_outputs(720) <= not (a and b);
    layer0_outputs(721) <= not b;
    layer0_outputs(722) <= a and not b;
    layer0_outputs(723) <= a or b;
    layer0_outputs(724) <= not a or b;
    layer0_outputs(725) <= not a or b;
    layer0_outputs(726) <= not (a and b);
    layer0_outputs(727) <= '0';
    layer0_outputs(728) <= b;
    layer0_outputs(729) <= b;
    layer0_outputs(730) <= not a;
    layer0_outputs(731) <= a and not b;
    layer0_outputs(732) <= b and not a;
    layer0_outputs(733) <= not b;
    layer0_outputs(734) <= '0';
    layer0_outputs(735) <= not (a or b);
    layer0_outputs(736) <= a;
    layer0_outputs(737) <= not a or b;
    layer0_outputs(738) <= b and not a;
    layer0_outputs(739) <= not b or a;
    layer0_outputs(740) <= not b;
    layer0_outputs(741) <= a and not b;
    layer0_outputs(742) <= a xor b;
    layer0_outputs(743) <= not b or a;
    layer0_outputs(744) <= not b;
    layer0_outputs(745) <= not (a xor b);
    layer0_outputs(746) <= b;
    layer0_outputs(747) <= a and not b;
    layer0_outputs(748) <= not (a xor b);
    layer0_outputs(749) <= a;
    layer0_outputs(750) <= b and not a;
    layer0_outputs(751) <= not a or b;
    layer0_outputs(752) <= b and not a;
    layer0_outputs(753) <= '1';
    layer0_outputs(754) <= a or b;
    layer0_outputs(755) <= '0';
    layer0_outputs(756) <= not a or b;
    layer0_outputs(757) <= b and not a;
    layer0_outputs(758) <= not a or b;
    layer0_outputs(759) <= not b or a;
    layer0_outputs(760) <= b;
    layer0_outputs(761) <= a;
    layer0_outputs(762) <= not (a xor b);
    layer0_outputs(763) <= not a or b;
    layer0_outputs(764) <= a;
    layer0_outputs(765) <= b;
    layer0_outputs(766) <= a;
    layer0_outputs(767) <= a or b;
    layer0_outputs(768) <= not b;
    layer0_outputs(769) <= '1';
    layer0_outputs(770) <= not (a or b);
    layer0_outputs(771) <= not (a and b);
    layer0_outputs(772) <= not b or a;
    layer0_outputs(773) <= '1';
    layer0_outputs(774) <= a or b;
    layer0_outputs(775) <= not (a xor b);
    layer0_outputs(776) <= '0';
    layer0_outputs(777) <= a and not b;
    layer0_outputs(778) <= a and b;
    layer0_outputs(779) <= a xor b;
    layer0_outputs(780) <= not b or a;
    layer0_outputs(781) <= not (a xor b);
    layer0_outputs(782) <= b;
    layer0_outputs(783) <= a xor b;
    layer0_outputs(784) <= not (a or b);
    layer0_outputs(785) <= a or b;
    layer0_outputs(786) <= not (a xor b);
    layer0_outputs(787) <= not (a or b);
    layer0_outputs(788) <= a and b;
    layer0_outputs(789) <= '1';
    layer0_outputs(790) <= not b;
    layer0_outputs(791) <= a;
    layer0_outputs(792) <= a;
    layer0_outputs(793) <= b;
    layer0_outputs(794) <= not (a xor b);
    layer0_outputs(795) <= not a;
    layer0_outputs(796) <= not a;
    layer0_outputs(797) <= not b;
    layer0_outputs(798) <= not a or b;
    layer0_outputs(799) <= not (a and b);
    layer0_outputs(800) <= not (a and b);
    layer0_outputs(801) <= a or b;
    layer0_outputs(802) <= '1';
    layer0_outputs(803) <= a and not b;
    layer0_outputs(804) <= not (a or b);
    layer0_outputs(805) <= not (a xor b);
    layer0_outputs(806) <= a;
    layer0_outputs(807) <= not a;
    layer0_outputs(808) <= a;
    layer0_outputs(809) <= a and not b;
    layer0_outputs(810) <= not b or a;
    layer0_outputs(811) <= not a;
    layer0_outputs(812) <= not b;
    layer0_outputs(813) <= not a or b;
    layer0_outputs(814) <= not a or b;
    layer0_outputs(815) <= a or b;
    layer0_outputs(816) <= a and b;
    layer0_outputs(817) <= not b or a;
    layer0_outputs(818) <= a;
    layer0_outputs(819) <= not b;
    layer0_outputs(820) <= a or b;
    layer0_outputs(821) <= not (a or b);
    layer0_outputs(822) <= not a or b;
    layer0_outputs(823) <= not (a xor b);
    layer0_outputs(824) <= b and not a;
    layer0_outputs(825) <= not b or a;
    layer0_outputs(826) <= a;
    layer0_outputs(827) <= not a or b;
    layer0_outputs(828) <= a and not b;
    layer0_outputs(829) <= not b;
    layer0_outputs(830) <= not (a or b);
    layer0_outputs(831) <= a and not b;
    layer0_outputs(832) <= a and not b;
    layer0_outputs(833) <= not (a or b);
    layer0_outputs(834) <= not (a or b);
    layer0_outputs(835) <= a;
    layer0_outputs(836) <= b;
    layer0_outputs(837) <= b and not a;
    layer0_outputs(838) <= a;
    layer0_outputs(839) <= not a or b;
    layer0_outputs(840) <= '0';
    layer0_outputs(841) <= a or b;
    layer0_outputs(842) <= not a or b;
    layer0_outputs(843) <= a xor b;
    layer0_outputs(844) <= a xor b;
    layer0_outputs(845) <= a or b;
    layer0_outputs(846) <= not a or b;
    layer0_outputs(847) <= b;
    layer0_outputs(848) <= not (a and b);
    layer0_outputs(849) <= b;
    layer0_outputs(850) <= not b or a;
    layer0_outputs(851) <= a and not b;
    layer0_outputs(852) <= not (a xor b);
    layer0_outputs(853) <= not (a and b);
    layer0_outputs(854) <= not b;
    layer0_outputs(855) <= a xor b;
    layer0_outputs(856) <= a;
    layer0_outputs(857) <= b and not a;
    layer0_outputs(858) <= a;
    layer0_outputs(859) <= not b or a;
    layer0_outputs(860) <= '0';
    layer0_outputs(861) <= not a;
    layer0_outputs(862) <= a and not b;
    layer0_outputs(863) <= a;
    layer0_outputs(864) <= not a or b;
    layer0_outputs(865) <= '0';
    layer0_outputs(866) <= a and b;
    layer0_outputs(867) <= not (a and b);
    layer0_outputs(868) <= b;
    layer0_outputs(869) <= b and not a;
    layer0_outputs(870) <= not a;
    layer0_outputs(871) <= not (a xor b);
    layer0_outputs(872) <= not (a or b);
    layer0_outputs(873) <= '1';
    layer0_outputs(874) <= '0';
    layer0_outputs(875) <= not a or b;
    layer0_outputs(876) <= a and not b;
    layer0_outputs(877) <= b;
    layer0_outputs(878) <= not (a and b);
    layer0_outputs(879) <= not b;
    layer0_outputs(880) <= a and not b;
    layer0_outputs(881) <= a and not b;
    layer0_outputs(882) <= not a;
    layer0_outputs(883) <= not b or a;
    layer0_outputs(884) <= not (a or b);
    layer0_outputs(885) <= b and not a;
    layer0_outputs(886) <= a;
    layer0_outputs(887) <= not (a and b);
    layer0_outputs(888) <= b and not a;
    layer0_outputs(889) <= a and not b;
    layer0_outputs(890) <= a and not b;
    layer0_outputs(891) <= b;
    layer0_outputs(892) <= b;
    layer0_outputs(893) <= not a or b;
    layer0_outputs(894) <= not (a or b);
    layer0_outputs(895) <= not (a and b);
    layer0_outputs(896) <= b;
    layer0_outputs(897) <= not (a xor b);
    layer0_outputs(898) <= not a;
    layer0_outputs(899) <= not b or a;
    layer0_outputs(900) <= not a;
    layer0_outputs(901) <= not (a or b);
    layer0_outputs(902) <= not a;
    layer0_outputs(903) <= a and not b;
    layer0_outputs(904) <= not b or a;
    layer0_outputs(905) <= a or b;
    layer0_outputs(906) <= a and not b;
    layer0_outputs(907) <= '0';
    layer0_outputs(908) <= b and not a;
    layer0_outputs(909) <= a and b;
    layer0_outputs(910) <= not (a or b);
    layer0_outputs(911) <= a or b;
    layer0_outputs(912) <= b and not a;
    layer0_outputs(913) <= not (a xor b);
    layer0_outputs(914) <= b;
    layer0_outputs(915) <= not b;
    layer0_outputs(916) <= not a;
    layer0_outputs(917) <= a or b;
    layer0_outputs(918) <= not (a or b);
    layer0_outputs(919) <= not b;
    layer0_outputs(920) <= not a;
    layer0_outputs(921) <= not b;
    layer0_outputs(922) <= not a or b;
    layer0_outputs(923) <= not (a and b);
    layer0_outputs(924) <= a;
    layer0_outputs(925) <= not b;
    layer0_outputs(926) <= a and b;
    layer0_outputs(927) <= '1';
    layer0_outputs(928) <= not (a or b);
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= b;
    layer0_outputs(931) <= a and b;
    layer0_outputs(932) <= b and not a;
    layer0_outputs(933) <= a or b;
    layer0_outputs(934) <= a and b;
    layer0_outputs(935) <= not b or a;
    layer0_outputs(936) <= not (a or b);
    layer0_outputs(937) <= not (a and b);
    layer0_outputs(938) <= '0';
    layer0_outputs(939) <= not (a xor b);
    layer0_outputs(940) <= not b or a;
    layer0_outputs(941) <= a and not b;
    layer0_outputs(942) <= a xor b;
    layer0_outputs(943) <= b and not a;
    layer0_outputs(944) <= not (a xor b);
    layer0_outputs(945) <= not (a or b);
    layer0_outputs(946) <= not (a or b);
    layer0_outputs(947) <= b and not a;
    layer0_outputs(948) <= b and not a;
    layer0_outputs(949) <= a or b;
    layer0_outputs(950) <= '1';
    layer0_outputs(951) <= '0';
    layer0_outputs(952) <= not b;
    layer0_outputs(953) <= not (a xor b);
    layer0_outputs(954) <= not a or b;
    layer0_outputs(955) <= not (a xor b);
    layer0_outputs(956) <= b;
    layer0_outputs(957) <= a and not b;
    layer0_outputs(958) <= not (a xor b);
    layer0_outputs(959) <= not b or a;
    layer0_outputs(960) <= not a;
    layer0_outputs(961) <= not a or b;
    layer0_outputs(962) <= b;
    layer0_outputs(963) <= not a;
    layer0_outputs(964) <= '1';
    layer0_outputs(965) <= not b or a;
    layer0_outputs(966) <= '0';
    layer0_outputs(967) <= a or b;
    layer0_outputs(968) <= not a or b;
    layer0_outputs(969) <= a or b;
    layer0_outputs(970) <= b;
    layer0_outputs(971) <= not a;
    layer0_outputs(972) <= not (a or b);
    layer0_outputs(973) <= not b;
    layer0_outputs(974) <= not a;
    layer0_outputs(975) <= not (a or b);
    layer0_outputs(976) <= not b;
    layer0_outputs(977) <= not (a xor b);
    layer0_outputs(978) <= not (a xor b);
    layer0_outputs(979) <= a;
    layer0_outputs(980) <= '1';
    layer0_outputs(981) <= not a;
    layer0_outputs(982) <= '0';
    layer0_outputs(983) <= not a;
    layer0_outputs(984) <= a or b;
    layer0_outputs(985) <= not (a and b);
    layer0_outputs(986) <= b;
    layer0_outputs(987) <= b;
    layer0_outputs(988) <= not (a or b);
    layer0_outputs(989) <= not b;
    layer0_outputs(990) <= a;
    layer0_outputs(991) <= a;
    layer0_outputs(992) <= '0';
    layer0_outputs(993) <= a xor b;
    layer0_outputs(994) <= a xor b;
    layer0_outputs(995) <= '1';
    layer0_outputs(996) <= b;
    layer0_outputs(997) <= a and b;
    layer0_outputs(998) <= not (a or b);
    layer0_outputs(999) <= a xor b;
    layer0_outputs(1000) <= a or b;
    layer0_outputs(1001) <= b and not a;
    layer0_outputs(1002) <= '1';
    layer0_outputs(1003) <= a or b;
    layer0_outputs(1004) <= a xor b;
    layer0_outputs(1005) <= a and not b;
    layer0_outputs(1006) <= '1';
    layer0_outputs(1007) <= a;
    layer0_outputs(1008) <= '1';
    layer0_outputs(1009) <= a;
    layer0_outputs(1010) <= not b;
    layer0_outputs(1011) <= not (a or b);
    layer0_outputs(1012) <= not (a xor b);
    layer0_outputs(1013) <= not (a xor b);
    layer0_outputs(1014) <= b and not a;
    layer0_outputs(1015) <= b;
    layer0_outputs(1016) <= a and not b;
    layer0_outputs(1017) <= '1';
    layer0_outputs(1018) <= not (a or b);
    layer0_outputs(1019) <= b;
    layer0_outputs(1020) <= b and not a;
    layer0_outputs(1021) <= not b or a;
    layer0_outputs(1022) <= '1';
    layer0_outputs(1023) <= not a;
    layer0_outputs(1024) <= a or b;
    layer0_outputs(1025) <= '1';
    layer0_outputs(1026) <= not b;
    layer0_outputs(1027) <= b and not a;
    layer0_outputs(1028) <= not (a and b);
    layer0_outputs(1029) <= b;
    layer0_outputs(1030) <= not (a xor b);
    layer0_outputs(1031) <= not (a or b);
    layer0_outputs(1032) <= a xor b;
    layer0_outputs(1033) <= not b;
    layer0_outputs(1034) <= a and b;
    layer0_outputs(1035) <= not a;
    layer0_outputs(1036) <= a and b;
    layer0_outputs(1037) <= not a or b;
    layer0_outputs(1038) <= a xor b;
    layer0_outputs(1039) <= a;
    layer0_outputs(1040) <= '0';
    layer0_outputs(1041) <= a xor b;
    layer0_outputs(1042) <= b;
    layer0_outputs(1043) <= not (a and b);
    layer0_outputs(1044) <= a and not b;
    layer0_outputs(1045) <= not a;
    layer0_outputs(1046) <= not a;
    layer0_outputs(1047) <= not a;
    layer0_outputs(1048) <= b;
    layer0_outputs(1049) <= '0';
    layer0_outputs(1050) <= b and not a;
    layer0_outputs(1051) <= a;
    layer0_outputs(1052) <= not b;
    layer0_outputs(1053) <= not (a or b);
    layer0_outputs(1054) <= a and not b;
    layer0_outputs(1055) <= a xor b;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= not b or a;
    layer0_outputs(1058) <= not (a or b);
    layer0_outputs(1059) <= '0';
    layer0_outputs(1060) <= b;
    layer0_outputs(1061) <= not (a xor b);
    layer0_outputs(1062) <= a;
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= not (a and b);
    layer0_outputs(1065) <= b and not a;
    layer0_outputs(1066) <= not b;
    layer0_outputs(1067) <= not (a or b);
    layer0_outputs(1068) <= a and b;
    layer0_outputs(1069) <= not (a or b);
    layer0_outputs(1070) <= a;
    layer0_outputs(1071) <= not a;
    layer0_outputs(1072) <= not (a xor b);
    layer0_outputs(1073) <= not (a xor b);
    layer0_outputs(1074) <= a;
    layer0_outputs(1075) <= b and not a;
    layer0_outputs(1076) <= a and b;
    layer0_outputs(1077) <= b;
    layer0_outputs(1078) <= a or b;
    layer0_outputs(1079) <= not (a xor b);
    layer0_outputs(1080) <= a xor b;
    layer0_outputs(1081) <= '0';
    layer0_outputs(1082) <= not b;
    layer0_outputs(1083) <= b;
    layer0_outputs(1084) <= not (a and b);
    layer0_outputs(1085) <= a and not b;
    layer0_outputs(1086) <= a;
    layer0_outputs(1087) <= a or b;
    layer0_outputs(1088) <= '1';
    layer0_outputs(1089) <= not (a and b);
    layer0_outputs(1090) <= a;
    layer0_outputs(1091) <= b and not a;
    layer0_outputs(1092) <= '0';
    layer0_outputs(1093) <= a;
    layer0_outputs(1094) <= a or b;
    layer0_outputs(1095) <= not (a xor b);
    layer0_outputs(1096) <= a and b;
    layer0_outputs(1097) <= a and not b;
    layer0_outputs(1098) <= not a;
    layer0_outputs(1099) <= not a or b;
    layer0_outputs(1100) <= b and not a;
    layer0_outputs(1101) <= a;
    layer0_outputs(1102) <= b and not a;
    layer0_outputs(1103) <= not b;
    layer0_outputs(1104) <= a and b;
    layer0_outputs(1105) <= b and not a;
    layer0_outputs(1106) <= a and not b;
    layer0_outputs(1107) <= not b or a;
    layer0_outputs(1108) <= a or b;
    layer0_outputs(1109) <= b and not a;
    layer0_outputs(1110) <= '0';
    layer0_outputs(1111) <= a;
    layer0_outputs(1112) <= not b or a;
    layer0_outputs(1113) <= a xor b;
    layer0_outputs(1114) <= '0';
    layer0_outputs(1115) <= not (a xor b);
    layer0_outputs(1116) <= not b or a;
    layer0_outputs(1117) <= a and b;
    layer0_outputs(1118) <= a or b;
    layer0_outputs(1119) <= a and b;
    layer0_outputs(1120) <= a or b;
    layer0_outputs(1121) <= b;
    layer0_outputs(1122) <= a and not b;
    layer0_outputs(1123) <= a or b;
    layer0_outputs(1124) <= '1';
    layer0_outputs(1125) <= b;
    layer0_outputs(1126) <= not a;
    layer0_outputs(1127) <= not (a or b);
    layer0_outputs(1128) <= b;
    layer0_outputs(1129) <= not (a and b);
    layer0_outputs(1130) <= not a;
    layer0_outputs(1131) <= '0';
    layer0_outputs(1132) <= b and not a;
    layer0_outputs(1133) <= not a;
    layer0_outputs(1134) <= not (a or b);
    layer0_outputs(1135) <= not (a or b);
    layer0_outputs(1136) <= a;
    layer0_outputs(1137) <= a;
    layer0_outputs(1138) <= a and b;
    layer0_outputs(1139) <= not (a and b);
    layer0_outputs(1140) <= a;
    layer0_outputs(1141) <= not a;
    layer0_outputs(1142) <= a and b;
    layer0_outputs(1143) <= '1';
    layer0_outputs(1144) <= '1';
    layer0_outputs(1145) <= a and b;
    layer0_outputs(1146) <= a and b;
    layer0_outputs(1147) <= not b or a;
    layer0_outputs(1148) <= not (a xor b);
    layer0_outputs(1149) <= not b;
    layer0_outputs(1150) <= a xor b;
    layer0_outputs(1151) <= b;
    layer0_outputs(1152) <= not (a or b);
    layer0_outputs(1153) <= not (a or b);
    layer0_outputs(1154) <= not a or b;
    layer0_outputs(1155) <= b;
    layer0_outputs(1156) <= not a;
    layer0_outputs(1157) <= not (a xor b);
    layer0_outputs(1158) <= not a;
    layer0_outputs(1159) <= a and b;
    layer0_outputs(1160) <= b;
    layer0_outputs(1161) <= '1';
    layer0_outputs(1162) <= not (a or b);
    layer0_outputs(1163) <= a xor b;
    layer0_outputs(1164) <= not (a or b);
    layer0_outputs(1165) <= not b or a;
    layer0_outputs(1166) <= '1';
    layer0_outputs(1167) <= b and not a;
    layer0_outputs(1168) <= not (a or b);
    layer0_outputs(1169) <= not b;
    layer0_outputs(1170) <= not a;
    layer0_outputs(1171) <= not (a or b);
    layer0_outputs(1172) <= b;
    layer0_outputs(1173) <= '1';
    layer0_outputs(1174) <= a and b;
    layer0_outputs(1175) <= not a;
    layer0_outputs(1176) <= a;
    layer0_outputs(1177) <= not (a or b);
    layer0_outputs(1178) <= '0';
    layer0_outputs(1179) <= not b or a;
    layer0_outputs(1180) <= not a or b;
    layer0_outputs(1181) <= not (a and b);
    layer0_outputs(1182) <= not (a or b);
    layer0_outputs(1183) <= not (a xor b);
    layer0_outputs(1184) <= not a or b;
    layer0_outputs(1185) <= a or b;
    layer0_outputs(1186) <= '1';
    layer0_outputs(1187) <= b and not a;
    layer0_outputs(1188) <= a or b;
    layer0_outputs(1189) <= not b;
    layer0_outputs(1190) <= not (a xor b);
    layer0_outputs(1191) <= not (a and b);
    layer0_outputs(1192) <= not (a or b);
    layer0_outputs(1193) <= not a;
    layer0_outputs(1194) <= a and not b;
    layer0_outputs(1195) <= not (a or b);
    layer0_outputs(1196) <= not a or b;
    layer0_outputs(1197) <= not (a or b);
    layer0_outputs(1198) <= not (a or b);
    layer0_outputs(1199) <= b and not a;
    layer0_outputs(1200) <= not a;
    layer0_outputs(1201) <= not a;
    layer0_outputs(1202) <= not (a xor b);
    layer0_outputs(1203) <= not (a or b);
    layer0_outputs(1204) <= a and b;
    layer0_outputs(1205) <= '0';
    layer0_outputs(1206) <= a and b;
    layer0_outputs(1207) <= not a;
    layer0_outputs(1208) <= '1';
    layer0_outputs(1209) <= not a or b;
    layer0_outputs(1210) <= not (a or b);
    layer0_outputs(1211) <= not (a xor b);
    layer0_outputs(1212) <= '0';
    layer0_outputs(1213) <= not (a or b);
    layer0_outputs(1214) <= b;
    layer0_outputs(1215) <= a or b;
    layer0_outputs(1216) <= not b;
    layer0_outputs(1217) <= not b;
    layer0_outputs(1218) <= a or b;
    layer0_outputs(1219) <= not (a and b);
    layer0_outputs(1220) <= b;
    layer0_outputs(1221) <= a or b;
    layer0_outputs(1222) <= a and not b;
    layer0_outputs(1223) <= a and not b;
    layer0_outputs(1224) <= not (a or b);
    layer0_outputs(1225) <= not (a and b);
    layer0_outputs(1226) <= b and not a;
    layer0_outputs(1227) <= not a or b;
    layer0_outputs(1228) <= b and not a;
    layer0_outputs(1229) <= not a;
    layer0_outputs(1230) <= '0';
    layer0_outputs(1231) <= not b;
    layer0_outputs(1232) <= a or b;
    layer0_outputs(1233) <= a and not b;
    layer0_outputs(1234) <= not b or a;
    layer0_outputs(1235) <= '0';
    layer0_outputs(1236) <= a or b;
    layer0_outputs(1237) <= a and b;
    layer0_outputs(1238) <= not (a xor b);
    layer0_outputs(1239) <= not b;
    layer0_outputs(1240) <= not b or a;
    layer0_outputs(1241) <= a;
    layer0_outputs(1242) <= a xor b;
    layer0_outputs(1243) <= b;
    layer0_outputs(1244) <= not b or a;
    layer0_outputs(1245) <= not a;
    layer0_outputs(1246) <= not a or b;
    layer0_outputs(1247) <= '0';
    layer0_outputs(1248) <= not a or b;
    layer0_outputs(1249) <= not (a or b);
    layer0_outputs(1250) <= a and not b;
    layer0_outputs(1251) <= a or b;
    layer0_outputs(1252) <= a and b;
    layer0_outputs(1253) <= a xor b;
    layer0_outputs(1254) <= b and not a;
    layer0_outputs(1255) <= b;
    layer0_outputs(1256) <= not (a and b);
    layer0_outputs(1257) <= not a;
    layer0_outputs(1258) <= not (a or b);
    layer0_outputs(1259) <= not (a or b);
    layer0_outputs(1260) <= not a or b;
    layer0_outputs(1261) <= a and not b;
    layer0_outputs(1262) <= not (a xor b);
    layer0_outputs(1263) <= a;
    layer0_outputs(1264) <= a and b;
    layer0_outputs(1265) <= not (a or b);
    layer0_outputs(1266) <= a and b;
    layer0_outputs(1267) <= a or b;
    layer0_outputs(1268) <= b;
    layer0_outputs(1269) <= '1';
    layer0_outputs(1270) <= not b;
    layer0_outputs(1271) <= not (a and b);
    layer0_outputs(1272) <= a or b;
    layer0_outputs(1273) <= a and not b;
    layer0_outputs(1274) <= not a or b;
    layer0_outputs(1275) <= not (a and b);
    layer0_outputs(1276) <= not a or b;
    layer0_outputs(1277) <= not a or b;
    layer0_outputs(1278) <= not b or a;
    layer0_outputs(1279) <= b and not a;
    layer0_outputs(1280) <= b and not a;
    layer0_outputs(1281) <= not b or a;
    layer0_outputs(1282) <= '0';
    layer0_outputs(1283) <= not a;
    layer0_outputs(1284) <= not (a or b);
    layer0_outputs(1285) <= not a or b;
    layer0_outputs(1286) <= b and not a;
    layer0_outputs(1287) <= a xor b;
    layer0_outputs(1288) <= a and not b;
    layer0_outputs(1289) <= not a;
    layer0_outputs(1290) <= a xor b;
    layer0_outputs(1291) <= a;
    layer0_outputs(1292) <= not (a and b);
    layer0_outputs(1293) <= b and not a;
    layer0_outputs(1294) <= not a or b;
    layer0_outputs(1295) <= a and b;
    layer0_outputs(1296) <= b and not a;
    layer0_outputs(1297) <= not a;
    layer0_outputs(1298) <= a;
    layer0_outputs(1299) <= a and b;
    layer0_outputs(1300) <= not (a and b);
    layer0_outputs(1301) <= a and b;
    layer0_outputs(1302) <= b and not a;
    layer0_outputs(1303) <= b and not a;
    layer0_outputs(1304) <= not (a or b);
    layer0_outputs(1305) <= not b or a;
    layer0_outputs(1306) <= not (a and b);
    layer0_outputs(1307) <= not b;
    layer0_outputs(1308) <= not (a or b);
    layer0_outputs(1309) <= '0';
    layer0_outputs(1310) <= a or b;
    layer0_outputs(1311) <= not (a and b);
    layer0_outputs(1312) <= not b;
    layer0_outputs(1313) <= a;
    layer0_outputs(1314) <= not b;
    layer0_outputs(1315) <= not b or a;
    layer0_outputs(1316) <= a or b;
    layer0_outputs(1317) <= not a;
    layer0_outputs(1318) <= not a;
    layer0_outputs(1319) <= b and not a;
    layer0_outputs(1320) <= not b;
    layer0_outputs(1321) <= a xor b;
    layer0_outputs(1322) <= not (a or b);
    layer0_outputs(1323) <= a and not b;
    layer0_outputs(1324) <= not a or b;
    layer0_outputs(1325) <= not b;
    layer0_outputs(1326) <= not a;
    layer0_outputs(1327) <= a xor b;
    layer0_outputs(1328) <= a or b;
    layer0_outputs(1329) <= a or b;
    layer0_outputs(1330) <= not (a and b);
    layer0_outputs(1331) <= a;
    layer0_outputs(1332) <= not a or b;
    layer0_outputs(1333) <= not b;
    layer0_outputs(1334) <= not a;
    layer0_outputs(1335) <= not b;
    layer0_outputs(1336) <= not (a xor b);
    layer0_outputs(1337) <= not b or a;
    layer0_outputs(1338) <= a xor b;
    layer0_outputs(1339) <= '0';
    layer0_outputs(1340) <= not b or a;
    layer0_outputs(1341) <= a or b;
    layer0_outputs(1342) <= a and b;
    layer0_outputs(1343) <= a or b;
    layer0_outputs(1344) <= a or b;
    layer0_outputs(1345) <= a and b;
    layer0_outputs(1346) <= not b;
    layer0_outputs(1347) <= b;
    layer0_outputs(1348) <= '1';
    layer0_outputs(1349) <= a or b;
    layer0_outputs(1350) <= not b;
    layer0_outputs(1351) <= not (a xor b);
    layer0_outputs(1352) <= not a or b;
    layer0_outputs(1353) <= not (a and b);
    layer0_outputs(1354) <= not (a xor b);
    layer0_outputs(1355) <= a or b;
    layer0_outputs(1356) <= '1';
    layer0_outputs(1357) <= not (a or b);
    layer0_outputs(1358) <= not (a and b);
    layer0_outputs(1359) <= not b;
    layer0_outputs(1360) <= a and b;
    layer0_outputs(1361) <= a;
    layer0_outputs(1362) <= a or b;
    layer0_outputs(1363) <= a xor b;
    layer0_outputs(1364) <= '0';
    layer0_outputs(1365) <= not (a and b);
    layer0_outputs(1366) <= b;
    layer0_outputs(1367) <= not (a or b);
    layer0_outputs(1368) <= b and not a;
    layer0_outputs(1369) <= not (a xor b);
    layer0_outputs(1370) <= not (a xor b);
    layer0_outputs(1371) <= not (a xor b);
    layer0_outputs(1372) <= a or b;
    layer0_outputs(1373) <= not b or a;
    layer0_outputs(1374) <= b and not a;
    layer0_outputs(1375) <= '1';
    layer0_outputs(1376) <= not (a xor b);
    layer0_outputs(1377) <= not a;
    layer0_outputs(1378) <= '1';
    layer0_outputs(1379) <= not a;
    layer0_outputs(1380) <= a;
    layer0_outputs(1381) <= not b;
    layer0_outputs(1382) <= b and not a;
    layer0_outputs(1383) <= not (a and b);
    layer0_outputs(1384) <= not (a xor b);
    layer0_outputs(1385) <= not (a and b);
    layer0_outputs(1386) <= b and not a;
    layer0_outputs(1387) <= not (a or b);
    layer0_outputs(1388) <= not b or a;
    layer0_outputs(1389) <= a xor b;
    layer0_outputs(1390) <= a;
    layer0_outputs(1391) <= not b or a;
    layer0_outputs(1392) <= a or b;
    layer0_outputs(1393) <= a and not b;
    layer0_outputs(1394) <= not (a xor b);
    layer0_outputs(1395) <= a xor b;
    layer0_outputs(1396) <= not b or a;
    layer0_outputs(1397) <= '1';
    layer0_outputs(1398) <= not (a or b);
    layer0_outputs(1399) <= not b;
    layer0_outputs(1400) <= not b or a;
    layer0_outputs(1401) <= not (a or b);
    layer0_outputs(1402) <= not a;
    layer0_outputs(1403) <= b and not a;
    layer0_outputs(1404) <= not b or a;
    layer0_outputs(1405) <= not b;
    layer0_outputs(1406) <= a and not b;
    layer0_outputs(1407) <= b;
    layer0_outputs(1408) <= not a or b;
    layer0_outputs(1409) <= a and not b;
    layer0_outputs(1410) <= not b or a;
    layer0_outputs(1411) <= a and not b;
    layer0_outputs(1412) <= not b;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= a and b;
    layer0_outputs(1415) <= not a or b;
    layer0_outputs(1416) <= a and not b;
    layer0_outputs(1417) <= not (a xor b);
    layer0_outputs(1418) <= not b or a;
    layer0_outputs(1419) <= not a;
    layer0_outputs(1420) <= b and not a;
    layer0_outputs(1421) <= a or b;
    layer0_outputs(1422) <= '0';
    layer0_outputs(1423) <= not b;
    layer0_outputs(1424) <= a;
    layer0_outputs(1425) <= not a or b;
    layer0_outputs(1426) <= not a or b;
    layer0_outputs(1427) <= not a;
    layer0_outputs(1428) <= not b;
    layer0_outputs(1429) <= b and not a;
    layer0_outputs(1430) <= not b or a;
    layer0_outputs(1431) <= b and not a;
    layer0_outputs(1432) <= not b;
    layer0_outputs(1433) <= not a;
    layer0_outputs(1434) <= b;
    layer0_outputs(1435) <= not b or a;
    layer0_outputs(1436) <= not (a and b);
    layer0_outputs(1437) <= not (a or b);
    layer0_outputs(1438) <= a or b;
    layer0_outputs(1439) <= not a or b;
    layer0_outputs(1440) <= not a or b;
    layer0_outputs(1441) <= a or b;
    layer0_outputs(1442) <= a and b;
    layer0_outputs(1443) <= not b;
    layer0_outputs(1444) <= not b or a;
    layer0_outputs(1445) <= a or b;
    layer0_outputs(1446) <= '1';
    layer0_outputs(1447) <= b and not a;
    layer0_outputs(1448) <= b;
    layer0_outputs(1449) <= not (a or b);
    layer0_outputs(1450) <= a;
    layer0_outputs(1451) <= not (a and b);
    layer0_outputs(1452) <= not (a or b);
    layer0_outputs(1453) <= '1';
    layer0_outputs(1454) <= a and not b;
    layer0_outputs(1455) <= not (a or b);
    layer0_outputs(1456) <= not b;
    layer0_outputs(1457) <= a;
    layer0_outputs(1458) <= not (a or b);
    layer0_outputs(1459) <= not (a or b);
    layer0_outputs(1460) <= not (a or b);
    layer0_outputs(1461) <= a;
    layer0_outputs(1462) <= not (a or b);
    layer0_outputs(1463) <= not a or b;
    layer0_outputs(1464) <= a or b;
    layer0_outputs(1465) <= not a or b;
    layer0_outputs(1466) <= not (a xor b);
    layer0_outputs(1467) <= b;
    layer0_outputs(1468) <= a and b;
    layer0_outputs(1469) <= not b;
    layer0_outputs(1470) <= '0';
    layer0_outputs(1471) <= '1';
    layer0_outputs(1472) <= not a or b;
    layer0_outputs(1473) <= not b or a;
    layer0_outputs(1474) <= not (a xor b);
    layer0_outputs(1475) <= not a;
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= not (a xor b);
    layer0_outputs(1478) <= a or b;
    layer0_outputs(1479) <= a xor b;
    layer0_outputs(1480) <= not (a and b);
    layer0_outputs(1481) <= not b or a;
    layer0_outputs(1482) <= a xor b;
    layer0_outputs(1483) <= not (a or b);
    layer0_outputs(1484) <= not (a and b);
    layer0_outputs(1485) <= not (a and b);
    layer0_outputs(1486) <= not b;
    layer0_outputs(1487) <= not a;
    layer0_outputs(1488) <= '1';
    layer0_outputs(1489) <= not a;
    layer0_outputs(1490) <= not (a xor b);
    layer0_outputs(1491) <= not (a xor b);
    layer0_outputs(1492) <= not (a xor b);
    layer0_outputs(1493) <= a xor b;
    layer0_outputs(1494) <= not b or a;
    layer0_outputs(1495) <= not b;
    layer0_outputs(1496) <= not (a or b);
    layer0_outputs(1497) <= not (a or b);
    layer0_outputs(1498) <= not a;
    layer0_outputs(1499) <= not a or b;
    layer0_outputs(1500) <= b and not a;
    layer0_outputs(1501) <= a or b;
    layer0_outputs(1502) <= a or b;
    layer0_outputs(1503) <= not b;
    layer0_outputs(1504) <= b;
    layer0_outputs(1505) <= not a or b;
    layer0_outputs(1506) <= a and not b;
    layer0_outputs(1507) <= not b;
    layer0_outputs(1508) <= not b or a;
    layer0_outputs(1509) <= not a or b;
    layer0_outputs(1510) <= a or b;
    layer0_outputs(1511) <= not (a or b);
    layer0_outputs(1512) <= not (a xor b);
    layer0_outputs(1513) <= not b;
    layer0_outputs(1514) <= a xor b;
    layer0_outputs(1515) <= not (a or b);
    layer0_outputs(1516) <= '1';
    layer0_outputs(1517) <= not a;
    layer0_outputs(1518) <= a or b;
    layer0_outputs(1519) <= b;
    layer0_outputs(1520) <= b and not a;
    layer0_outputs(1521) <= not b;
    layer0_outputs(1522) <= not b;
    layer0_outputs(1523) <= a or b;
    layer0_outputs(1524) <= a or b;
    layer0_outputs(1525) <= not a;
    layer0_outputs(1526) <= not b;
    layer0_outputs(1527) <= not b;
    layer0_outputs(1528) <= not b;
    layer0_outputs(1529) <= '0';
    layer0_outputs(1530) <= a or b;
    layer0_outputs(1531) <= '1';
    layer0_outputs(1532) <= a;
    layer0_outputs(1533) <= not (a or b);
    layer0_outputs(1534) <= '0';
    layer0_outputs(1535) <= not a;
    layer0_outputs(1536) <= '1';
    layer0_outputs(1537) <= not b or a;
    layer0_outputs(1538) <= a and not b;
    layer0_outputs(1539) <= not a;
    layer0_outputs(1540) <= not b;
    layer0_outputs(1541) <= not a;
    layer0_outputs(1542) <= '1';
    layer0_outputs(1543) <= '1';
    layer0_outputs(1544) <= a and not b;
    layer0_outputs(1545) <= a or b;
    layer0_outputs(1546) <= not a;
    layer0_outputs(1547) <= not (a xor b);
    layer0_outputs(1548) <= not (a xor b);
    layer0_outputs(1549) <= not a;
    layer0_outputs(1550) <= b and not a;
    layer0_outputs(1551) <= '0';
    layer0_outputs(1552) <= a or b;
    layer0_outputs(1553) <= b;
    layer0_outputs(1554) <= not (a and b);
    layer0_outputs(1555) <= not b or a;
    layer0_outputs(1556) <= not (a or b);
    layer0_outputs(1557) <= not a;
    layer0_outputs(1558) <= not a;
    layer0_outputs(1559) <= not (a and b);
    layer0_outputs(1560) <= not a;
    layer0_outputs(1561) <= a;
    layer0_outputs(1562) <= not b or a;
    layer0_outputs(1563) <= a and not b;
    layer0_outputs(1564) <= a;
    layer0_outputs(1565) <= a or b;
    layer0_outputs(1566) <= not b or a;
    layer0_outputs(1567) <= not b or a;
    layer0_outputs(1568) <= not a or b;
    layer0_outputs(1569) <= not b;
    layer0_outputs(1570) <= a and b;
    layer0_outputs(1571) <= not b or a;
    layer0_outputs(1572) <= a and not b;
    layer0_outputs(1573) <= b;
    layer0_outputs(1574) <= a and b;
    layer0_outputs(1575) <= not b;
    layer0_outputs(1576) <= not b or a;
    layer0_outputs(1577) <= not (a xor b);
    layer0_outputs(1578) <= '1';
    layer0_outputs(1579) <= not b;
    layer0_outputs(1580) <= a and b;
    layer0_outputs(1581) <= a and not b;
    layer0_outputs(1582) <= not b;
    layer0_outputs(1583) <= a xor b;
    layer0_outputs(1584) <= a xor b;
    layer0_outputs(1585) <= a or b;
    layer0_outputs(1586) <= a;
    layer0_outputs(1587) <= not b;
    layer0_outputs(1588) <= not (a xor b);
    layer0_outputs(1589) <= b and not a;
    layer0_outputs(1590) <= b and not a;
    layer0_outputs(1591) <= '1';
    layer0_outputs(1592) <= b and not a;
    layer0_outputs(1593) <= not a;
    layer0_outputs(1594) <= not b or a;
    layer0_outputs(1595) <= not b;
    layer0_outputs(1596) <= a and b;
    layer0_outputs(1597) <= not b;
    layer0_outputs(1598) <= b;
    layer0_outputs(1599) <= b and not a;
    layer0_outputs(1600) <= a and b;
    layer0_outputs(1601) <= b;
    layer0_outputs(1602) <= not (a or b);
    layer0_outputs(1603) <= not b or a;
    layer0_outputs(1604) <= a or b;
    layer0_outputs(1605) <= not b or a;
    layer0_outputs(1606) <= a and not b;
    layer0_outputs(1607) <= not b or a;
    layer0_outputs(1608) <= b and not a;
    layer0_outputs(1609) <= not (a xor b);
    layer0_outputs(1610) <= b and not a;
    layer0_outputs(1611) <= '0';
    layer0_outputs(1612) <= not (a and b);
    layer0_outputs(1613) <= not (a or b);
    layer0_outputs(1614) <= not a or b;
    layer0_outputs(1615) <= not (a or b);
    layer0_outputs(1616) <= a and b;
    layer0_outputs(1617) <= not b or a;
    layer0_outputs(1618) <= not b;
    layer0_outputs(1619) <= not (a and b);
    layer0_outputs(1620) <= not (a xor b);
    layer0_outputs(1621) <= a or b;
    layer0_outputs(1622) <= not a;
    layer0_outputs(1623) <= not (a or b);
    layer0_outputs(1624) <= not a;
    layer0_outputs(1625) <= a or b;
    layer0_outputs(1626) <= '0';
    layer0_outputs(1627) <= b;
    layer0_outputs(1628) <= not (a xor b);
    layer0_outputs(1629) <= not b or a;
    layer0_outputs(1630) <= '0';
    layer0_outputs(1631) <= '1';
    layer0_outputs(1632) <= '1';
    layer0_outputs(1633) <= a xor b;
    layer0_outputs(1634) <= not a;
    layer0_outputs(1635) <= not a or b;
    layer0_outputs(1636) <= b;
    layer0_outputs(1637) <= not (a xor b);
    layer0_outputs(1638) <= a and not b;
    layer0_outputs(1639) <= not b;
    layer0_outputs(1640) <= a or b;
    layer0_outputs(1641) <= b;
    layer0_outputs(1642) <= not (a or b);
    layer0_outputs(1643) <= a;
    layer0_outputs(1644) <= not a or b;
    layer0_outputs(1645) <= a or b;
    layer0_outputs(1646) <= a;
    layer0_outputs(1647) <= not a;
    layer0_outputs(1648) <= a;
    layer0_outputs(1649) <= a;
    layer0_outputs(1650) <= '1';
    layer0_outputs(1651) <= not b or a;
    layer0_outputs(1652) <= a and not b;
    layer0_outputs(1653) <= a xor b;
    layer0_outputs(1654) <= a and b;
    layer0_outputs(1655) <= not (a or b);
    layer0_outputs(1656) <= not a;
    layer0_outputs(1657) <= not a;
    layer0_outputs(1658) <= b;
    layer0_outputs(1659) <= not b;
    layer0_outputs(1660) <= a xor b;
    layer0_outputs(1661) <= not (a xor b);
    layer0_outputs(1662) <= a or b;
    layer0_outputs(1663) <= not b or a;
    layer0_outputs(1664) <= not (a and b);
    layer0_outputs(1665) <= b;
    layer0_outputs(1666) <= a xor b;
    layer0_outputs(1667) <= b and not a;
    layer0_outputs(1668) <= a and not b;
    layer0_outputs(1669) <= b and not a;
    layer0_outputs(1670) <= a or b;
    layer0_outputs(1671) <= not b;
    layer0_outputs(1672) <= b;
    layer0_outputs(1673) <= not b;
    layer0_outputs(1674) <= not b;
    layer0_outputs(1675) <= a xor b;
    layer0_outputs(1676) <= not (a or b);
    layer0_outputs(1677) <= not a or b;
    layer0_outputs(1678) <= b and not a;
    layer0_outputs(1679) <= a and b;
    layer0_outputs(1680) <= a and not b;
    layer0_outputs(1681) <= '0';
    layer0_outputs(1682) <= a and b;
    layer0_outputs(1683) <= not a or b;
    layer0_outputs(1684) <= a xor b;
    layer0_outputs(1685) <= '1';
    layer0_outputs(1686) <= not a;
    layer0_outputs(1687) <= not b or a;
    layer0_outputs(1688) <= a and b;
    layer0_outputs(1689) <= b and not a;
    layer0_outputs(1690) <= not b or a;
    layer0_outputs(1691) <= a and b;
    layer0_outputs(1692) <= a or b;
    layer0_outputs(1693) <= a and not b;
    layer0_outputs(1694) <= a and b;
    layer0_outputs(1695) <= not b;
    layer0_outputs(1696) <= not (a xor b);
    layer0_outputs(1697) <= not (a xor b);
    layer0_outputs(1698) <= not (a xor b);
    layer0_outputs(1699) <= not a or b;
    layer0_outputs(1700) <= not a or b;
    layer0_outputs(1701) <= not b;
    layer0_outputs(1702) <= not a or b;
    layer0_outputs(1703) <= '1';
    layer0_outputs(1704) <= b and not a;
    layer0_outputs(1705) <= not a or b;
    layer0_outputs(1706) <= not (a or b);
    layer0_outputs(1707) <= not b or a;
    layer0_outputs(1708) <= a and not b;
    layer0_outputs(1709) <= not (a and b);
    layer0_outputs(1710) <= a xor b;
    layer0_outputs(1711) <= a xor b;
    layer0_outputs(1712) <= not (a or b);
    layer0_outputs(1713) <= not (a or b);
    layer0_outputs(1714) <= not (a xor b);
    layer0_outputs(1715) <= b;
    layer0_outputs(1716) <= a xor b;
    layer0_outputs(1717) <= a and b;
    layer0_outputs(1718) <= not (a or b);
    layer0_outputs(1719) <= '1';
    layer0_outputs(1720) <= a xor b;
    layer0_outputs(1721) <= a or b;
    layer0_outputs(1722) <= b;
    layer0_outputs(1723) <= a or b;
    layer0_outputs(1724) <= not (a or b);
    layer0_outputs(1725) <= not (a or b);
    layer0_outputs(1726) <= a xor b;
    layer0_outputs(1727) <= '1';
    layer0_outputs(1728) <= not b or a;
    layer0_outputs(1729) <= not (a xor b);
    layer0_outputs(1730) <= a and b;
    layer0_outputs(1731) <= a;
    layer0_outputs(1732) <= not (a xor b);
    layer0_outputs(1733) <= b;
    layer0_outputs(1734) <= b and not a;
    layer0_outputs(1735) <= a and not b;
    layer0_outputs(1736) <= not b;
    layer0_outputs(1737) <= a and not b;
    layer0_outputs(1738) <= b;
    layer0_outputs(1739) <= b;
    layer0_outputs(1740) <= b;
    layer0_outputs(1741) <= a or b;
    layer0_outputs(1742) <= not b or a;
    layer0_outputs(1743) <= not (a and b);
    layer0_outputs(1744) <= not b;
    layer0_outputs(1745) <= not (a xor b);
    layer0_outputs(1746) <= a;
    layer0_outputs(1747) <= a or b;
    layer0_outputs(1748) <= b;
    layer0_outputs(1749) <= a and b;
    layer0_outputs(1750) <= not b or a;
    layer0_outputs(1751) <= not b;
    layer0_outputs(1752) <= not (a xor b);
    layer0_outputs(1753) <= b and not a;
    layer0_outputs(1754) <= a and not b;
    layer0_outputs(1755) <= a and b;
    layer0_outputs(1756) <= '0';
    layer0_outputs(1757) <= not a or b;
    layer0_outputs(1758) <= b;
    layer0_outputs(1759) <= not b;
    layer0_outputs(1760) <= a and not b;
    layer0_outputs(1761) <= a or b;
    layer0_outputs(1762) <= not a;
    layer0_outputs(1763) <= b;
    layer0_outputs(1764) <= not a;
    layer0_outputs(1765) <= not a or b;
    layer0_outputs(1766) <= a;
    layer0_outputs(1767) <= not a;
    layer0_outputs(1768) <= not a or b;
    layer0_outputs(1769) <= '0';
    layer0_outputs(1770) <= not b;
    layer0_outputs(1771) <= not b or a;
    layer0_outputs(1772) <= b and not a;
    layer0_outputs(1773) <= a;
    layer0_outputs(1774) <= not (a and b);
    layer0_outputs(1775) <= a xor b;
    layer0_outputs(1776) <= not a or b;
    layer0_outputs(1777) <= not b or a;
    layer0_outputs(1778) <= '0';
    layer0_outputs(1779) <= not a;
    layer0_outputs(1780) <= '1';
    layer0_outputs(1781) <= b;
    layer0_outputs(1782) <= a or b;
    layer0_outputs(1783) <= a and b;
    layer0_outputs(1784) <= a xor b;
    layer0_outputs(1785) <= a and b;
    layer0_outputs(1786) <= not b;
    layer0_outputs(1787) <= b;
    layer0_outputs(1788) <= b;
    layer0_outputs(1789) <= not a;
    layer0_outputs(1790) <= a xor b;
    layer0_outputs(1791) <= not (a or b);
    layer0_outputs(1792) <= not (a or b);
    layer0_outputs(1793) <= a and b;
    layer0_outputs(1794) <= not a or b;
    layer0_outputs(1795) <= '0';
    layer0_outputs(1796) <= not b;
    layer0_outputs(1797) <= not a;
    layer0_outputs(1798) <= not a or b;
    layer0_outputs(1799) <= not (a xor b);
    layer0_outputs(1800) <= not (a or b);
    layer0_outputs(1801) <= not b;
    layer0_outputs(1802) <= a or b;
    layer0_outputs(1803) <= '0';
    layer0_outputs(1804) <= b;
    layer0_outputs(1805) <= not (a and b);
    layer0_outputs(1806) <= b;
    layer0_outputs(1807) <= a and b;
    layer0_outputs(1808) <= b and not a;
    layer0_outputs(1809) <= a;
    layer0_outputs(1810) <= not a or b;
    layer0_outputs(1811) <= not (a and b);
    layer0_outputs(1812) <= a;
    layer0_outputs(1813) <= not a or b;
    layer0_outputs(1814) <= a and b;
    layer0_outputs(1815) <= '0';
    layer0_outputs(1816) <= '1';
    layer0_outputs(1817) <= not a;
    layer0_outputs(1818) <= not b;
    layer0_outputs(1819) <= not (a xor b);
    layer0_outputs(1820) <= b and not a;
    layer0_outputs(1821) <= a;
    layer0_outputs(1822) <= '1';
    layer0_outputs(1823) <= '0';
    layer0_outputs(1824) <= not (a xor b);
    layer0_outputs(1825) <= a and b;
    layer0_outputs(1826) <= a or b;
    layer0_outputs(1827) <= not a;
    layer0_outputs(1828) <= a xor b;
    layer0_outputs(1829) <= '1';
    layer0_outputs(1830) <= not b;
    layer0_outputs(1831) <= a or b;
    layer0_outputs(1832) <= a or b;
    layer0_outputs(1833) <= not a or b;
    layer0_outputs(1834) <= not (a xor b);
    layer0_outputs(1835) <= a and not b;
    layer0_outputs(1836) <= a or b;
    layer0_outputs(1837) <= not b;
    layer0_outputs(1838) <= a and not b;
    layer0_outputs(1839) <= b and not a;
    layer0_outputs(1840) <= '1';
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= a and not b;
    layer0_outputs(1843) <= a and not b;
    layer0_outputs(1844) <= '0';
    layer0_outputs(1845) <= a;
    layer0_outputs(1846) <= '1';
    layer0_outputs(1847) <= not b;
    layer0_outputs(1848) <= not (a and b);
    layer0_outputs(1849) <= not b or a;
    layer0_outputs(1850) <= a;
    layer0_outputs(1851) <= not a;
    layer0_outputs(1852) <= b;
    layer0_outputs(1853) <= '0';
    layer0_outputs(1854) <= a xor b;
    layer0_outputs(1855) <= not (a xor b);
    layer0_outputs(1856) <= not a or b;
    layer0_outputs(1857) <= not (a xor b);
    layer0_outputs(1858) <= not a or b;
    layer0_outputs(1859) <= a or b;
    layer0_outputs(1860) <= a or b;
    layer0_outputs(1861) <= not b or a;
    layer0_outputs(1862) <= a and not b;
    layer0_outputs(1863) <= a;
    layer0_outputs(1864) <= not b;
    layer0_outputs(1865) <= not (a xor b);
    layer0_outputs(1866) <= not b or a;
    layer0_outputs(1867) <= b;
    layer0_outputs(1868) <= b;
    layer0_outputs(1869) <= not (a xor b);
    layer0_outputs(1870) <= a or b;
    layer0_outputs(1871) <= not (a or b);
    layer0_outputs(1872) <= not (a and b);
    layer0_outputs(1873) <= a xor b;
    layer0_outputs(1874) <= b and not a;
    layer0_outputs(1875) <= a xor b;
    layer0_outputs(1876) <= a xor b;
    layer0_outputs(1877) <= '1';
    layer0_outputs(1878) <= a xor b;
    layer0_outputs(1879) <= not (a and b);
    layer0_outputs(1880) <= a and b;
    layer0_outputs(1881) <= not (a xor b);
    layer0_outputs(1882) <= not b;
    layer0_outputs(1883) <= b and not a;
    layer0_outputs(1884) <= not b or a;
    layer0_outputs(1885) <= a or b;
    layer0_outputs(1886) <= a;
    layer0_outputs(1887) <= not b or a;
    layer0_outputs(1888) <= not b;
    layer0_outputs(1889) <= not b or a;
    layer0_outputs(1890) <= a or b;
    layer0_outputs(1891) <= not a or b;
    layer0_outputs(1892) <= not b or a;
    layer0_outputs(1893) <= not (a xor b);
    layer0_outputs(1894) <= a xor b;
    layer0_outputs(1895) <= not (a xor b);
    layer0_outputs(1896) <= b and not a;
    layer0_outputs(1897) <= a and b;
    layer0_outputs(1898) <= a;
    layer0_outputs(1899) <= a and not b;
    layer0_outputs(1900) <= a;
    layer0_outputs(1901) <= a xor b;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= not b;
    layer0_outputs(1904) <= b;
    layer0_outputs(1905) <= b;
    layer0_outputs(1906) <= not b or a;
    layer0_outputs(1907) <= not (a and b);
    layer0_outputs(1908) <= '0';
    layer0_outputs(1909) <= b;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= a;
    layer0_outputs(1912) <= '0';
    layer0_outputs(1913) <= not a or b;
    layer0_outputs(1914) <= '1';
    layer0_outputs(1915) <= not (a and b);
    layer0_outputs(1916) <= not b or a;
    layer0_outputs(1917) <= a or b;
    layer0_outputs(1918) <= not (a and b);
    layer0_outputs(1919) <= not (a xor b);
    layer0_outputs(1920) <= a or b;
    layer0_outputs(1921) <= not b;
    layer0_outputs(1922) <= b and not a;
    layer0_outputs(1923) <= not a or b;
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= not b;
    layer0_outputs(1926) <= not (a xor b);
    layer0_outputs(1927) <= not a;
    layer0_outputs(1928) <= not (a or b);
    layer0_outputs(1929) <= a and b;
    layer0_outputs(1930) <= a and not b;
    layer0_outputs(1931) <= b and not a;
    layer0_outputs(1932) <= a and not b;
    layer0_outputs(1933) <= b;
    layer0_outputs(1934) <= a or b;
    layer0_outputs(1935) <= a;
    layer0_outputs(1936) <= not a or b;
    layer0_outputs(1937) <= a and b;
    layer0_outputs(1938) <= '1';
    layer0_outputs(1939) <= not (a or b);
    layer0_outputs(1940) <= not b or a;
    layer0_outputs(1941) <= a and not b;
    layer0_outputs(1942) <= a;
    layer0_outputs(1943) <= b and not a;
    layer0_outputs(1944) <= a or b;
    layer0_outputs(1945) <= a and b;
    layer0_outputs(1946) <= a xor b;
    layer0_outputs(1947) <= not (a or b);
    layer0_outputs(1948) <= not a;
    layer0_outputs(1949) <= not a or b;
    layer0_outputs(1950) <= '1';
    layer0_outputs(1951) <= b and not a;
    layer0_outputs(1952) <= not (a or b);
    layer0_outputs(1953) <= not b or a;
    layer0_outputs(1954) <= not b or a;
    layer0_outputs(1955) <= a and not b;
    layer0_outputs(1956) <= not b;
    layer0_outputs(1957) <= a xor b;
    layer0_outputs(1958) <= '1';
    layer0_outputs(1959) <= not a;
    layer0_outputs(1960) <= '1';
    layer0_outputs(1961) <= not a or b;
    layer0_outputs(1962) <= not a or b;
    layer0_outputs(1963) <= a and b;
    layer0_outputs(1964) <= not a;
    layer0_outputs(1965) <= b and not a;
    layer0_outputs(1966) <= not a or b;
    layer0_outputs(1967) <= '1';
    layer0_outputs(1968) <= a and b;
    layer0_outputs(1969) <= b and not a;
    layer0_outputs(1970) <= '0';
    layer0_outputs(1971) <= not (a and b);
    layer0_outputs(1972) <= not b;
    layer0_outputs(1973) <= not b or a;
    layer0_outputs(1974) <= '1';
    layer0_outputs(1975) <= not (a and b);
    layer0_outputs(1976) <= a or b;
    layer0_outputs(1977) <= not a;
    layer0_outputs(1978) <= a;
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a and b;
    layer0_outputs(1981) <= '1';
    layer0_outputs(1982) <= not (a or b);
    layer0_outputs(1983) <= a and b;
    layer0_outputs(1984) <= a or b;
    layer0_outputs(1985) <= '0';
    layer0_outputs(1986) <= a and not b;
    layer0_outputs(1987) <= b;
    layer0_outputs(1988) <= b;
    layer0_outputs(1989) <= a or b;
    layer0_outputs(1990) <= not b or a;
    layer0_outputs(1991) <= a or b;
    layer0_outputs(1992) <= a and not b;
    layer0_outputs(1993) <= not a or b;
    layer0_outputs(1994) <= not b or a;
    layer0_outputs(1995) <= '0';
    layer0_outputs(1996) <= '0';
    layer0_outputs(1997) <= not a or b;
    layer0_outputs(1998) <= '0';
    layer0_outputs(1999) <= a and not b;
    layer0_outputs(2000) <= a or b;
    layer0_outputs(2001) <= b;
    layer0_outputs(2002) <= b;
    layer0_outputs(2003) <= not b or a;
    layer0_outputs(2004) <= a or b;
    layer0_outputs(2005) <= not (a xor b);
    layer0_outputs(2006) <= b;
    layer0_outputs(2007) <= a;
    layer0_outputs(2008) <= a and not b;
    layer0_outputs(2009) <= b;
    layer0_outputs(2010) <= not b;
    layer0_outputs(2011) <= a or b;
    layer0_outputs(2012) <= not b;
    layer0_outputs(2013) <= not b or a;
    layer0_outputs(2014) <= not (a xor b);
    layer0_outputs(2015) <= not a or b;
    layer0_outputs(2016) <= a and b;
    layer0_outputs(2017) <= not (a and b);
    layer0_outputs(2018) <= not (a and b);
    layer0_outputs(2019) <= b;
    layer0_outputs(2020) <= not (a and b);
    layer0_outputs(2021) <= not a;
    layer0_outputs(2022) <= not a;
    layer0_outputs(2023) <= not b or a;
    layer0_outputs(2024) <= a and not b;
    layer0_outputs(2025) <= not (a or b);
    layer0_outputs(2026) <= not a;
    layer0_outputs(2027) <= not a or b;
    layer0_outputs(2028) <= not (a and b);
    layer0_outputs(2029) <= not b or a;
    layer0_outputs(2030) <= b and not a;
    layer0_outputs(2031) <= not (a xor b);
    layer0_outputs(2032) <= not a;
    layer0_outputs(2033) <= a xor b;
    layer0_outputs(2034) <= not a;
    layer0_outputs(2035) <= not a or b;
    layer0_outputs(2036) <= not a;
    layer0_outputs(2037) <= '1';
    layer0_outputs(2038) <= '0';
    layer0_outputs(2039) <= not (a and b);
    layer0_outputs(2040) <= not a;
    layer0_outputs(2041) <= a;
    layer0_outputs(2042) <= a and not b;
    layer0_outputs(2043) <= a;
    layer0_outputs(2044) <= not (a or b);
    layer0_outputs(2045) <= not (a and b);
    layer0_outputs(2046) <= not b or a;
    layer0_outputs(2047) <= not (a or b);
    layer0_outputs(2048) <= not b;
    layer0_outputs(2049) <= a or b;
    layer0_outputs(2050) <= not (a and b);
    layer0_outputs(2051) <= '1';
    layer0_outputs(2052) <= a and not b;
    layer0_outputs(2053) <= a and b;
    layer0_outputs(2054) <= '0';
    layer0_outputs(2055) <= not (a or b);
    layer0_outputs(2056) <= not (a or b);
    layer0_outputs(2057) <= not (a or b);
    layer0_outputs(2058) <= not (a or b);
    layer0_outputs(2059) <= a xor b;
    layer0_outputs(2060) <= b and not a;
    layer0_outputs(2061) <= not (a xor b);
    layer0_outputs(2062) <= b and not a;
    layer0_outputs(2063) <= not (a xor b);
    layer0_outputs(2064) <= not b or a;
    layer0_outputs(2065) <= not (a or b);
    layer0_outputs(2066) <= not a or b;
    layer0_outputs(2067) <= not a;
    layer0_outputs(2068) <= not b;
    layer0_outputs(2069) <= not (a or b);
    layer0_outputs(2070) <= not (a or b);
    layer0_outputs(2071) <= b and not a;
    layer0_outputs(2072) <= '0';
    layer0_outputs(2073) <= b;
    layer0_outputs(2074) <= not (a and b);
    layer0_outputs(2075) <= not a;
    layer0_outputs(2076) <= not a or b;
    layer0_outputs(2077) <= a and not b;
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= not (a xor b);
    layer0_outputs(2080) <= a or b;
    layer0_outputs(2081) <= not a;
    layer0_outputs(2082) <= not (a and b);
    layer0_outputs(2083) <= a and not b;
    layer0_outputs(2084) <= not b or a;
    layer0_outputs(2085) <= not a;
    layer0_outputs(2086) <= a xor b;
    layer0_outputs(2087) <= a xor b;
    layer0_outputs(2088) <= not (a or b);
    layer0_outputs(2089) <= not (a and b);
    layer0_outputs(2090) <= not b or a;
    layer0_outputs(2091) <= not (a xor b);
    layer0_outputs(2092) <= not b;
    layer0_outputs(2093) <= b and not a;
    layer0_outputs(2094) <= a or b;
    layer0_outputs(2095) <= a and not b;
    layer0_outputs(2096) <= a or b;
    layer0_outputs(2097) <= not a;
    layer0_outputs(2098) <= b and not a;
    layer0_outputs(2099) <= not b;
    layer0_outputs(2100) <= a and b;
    layer0_outputs(2101) <= a;
    layer0_outputs(2102) <= a and b;
    layer0_outputs(2103) <= '0';
    layer0_outputs(2104) <= a and b;
    layer0_outputs(2105) <= a and b;
    layer0_outputs(2106) <= not (a or b);
    layer0_outputs(2107) <= not a;
    layer0_outputs(2108) <= a and not b;
    layer0_outputs(2109) <= not (a or b);
    layer0_outputs(2110) <= a;
    layer0_outputs(2111) <= a and b;
    layer0_outputs(2112) <= not b;
    layer0_outputs(2113) <= a or b;
    layer0_outputs(2114) <= a xor b;
    layer0_outputs(2115) <= a xor b;
    layer0_outputs(2116) <= not (a or b);
    layer0_outputs(2117) <= not b;
    layer0_outputs(2118) <= b;
    layer0_outputs(2119) <= b and not a;
    layer0_outputs(2120) <= b;
    layer0_outputs(2121) <= b;
    layer0_outputs(2122) <= a and not b;
    layer0_outputs(2123) <= '0';
    layer0_outputs(2124) <= not a or b;
    layer0_outputs(2125) <= '0';
    layer0_outputs(2126) <= not b;
    layer0_outputs(2127) <= not (a and b);
    layer0_outputs(2128) <= a or b;
    layer0_outputs(2129) <= b and not a;
    layer0_outputs(2130) <= not a or b;
    layer0_outputs(2131) <= not a or b;
    layer0_outputs(2132) <= not b or a;
    layer0_outputs(2133) <= not (a and b);
    layer0_outputs(2134) <= not a or b;
    layer0_outputs(2135) <= a and not b;
    layer0_outputs(2136) <= a and b;
    layer0_outputs(2137) <= not b;
    layer0_outputs(2138) <= not a or b;
    layer0_outputs(2139) <= a and not b;
    layer0_outputs(2140) <= not a;
    layer0_outputs(2141) <= not (a or b);
    layer0_outputs(2142) <= a or b;
    layer0_outputs(2143) <= not (a or b);
    layer0_outputs(2144) <= b and not a;
    layer0_outputs(2145) <= not (a and b);
    layer0_outputs(2146) <= '1';
    layer0_outputs(2147) <= b and not a;
    layer0_outputs(2148) <= not b or a;
    layer0_outputs(2149) <= b;
    layer0_outputs(2150) <= b;
    layer0_outputs(2151) <= '1';
    layer0_outputs(2152) <= not a;
    layer0_outputs(2153) <= not (a and b);
    layer0_outputs(2154) <= a and not b;
    layer0_outputs(2155) <= a and b;
    layer0_outputs(2156) <= a;
    layer0_outputs(2157) <= b and not a;
    layer0_outputs(2158) <= a and b;
    layer0_outputs(2159) <= a;
    layer0_outputs(2160) <= not b;
    layer0_outputs(2161) <= not b;
    layer0_outputs(2162) <= not (a xor b);
    layer0_outputs(2163) <= b and not a;
    layer0_outputs(2164) <= b;
    layer0_outputs(2165) <= not (a or b);
    layer0_outputs(2166) <= not a;
    layer0_outputs(2167) <= not b or a;
    layer0_outputs(2168) <= not a or b;
    layer0_outputs(2169) <= a;
    layer0_outputs(2170) <= not (a or b);
    layer0_outputs(2171) <= a and not b;
    layer0_outputs(2172) <= b and not a;
    layer0_outputs(2173) <= not b;
    layer0_outputs(2174) <= not a or b;
    layer0_outputs(2175) <= not a or b;
    layer0_outputs(2176) <= a;
    layer0_outputs(2177) <= a and b;
    layer0_outputs(2178) <= '0';
    layer0_outputs(2179) <= not (a and b);
    layer0_outputs(2180) <= not b or a;
    layer0_outputs(2181) <= a and not b;
    layer0_outputs(2182) <= a;
    layer0_outputs(2183) <= not b or a;
    layer0_outputs(2184) <= a and not b;
    layer0_outputs(2185) <= a xor b;
    layer0_outputs(2186) <= b and not a;
    layer0_outputs(2187) <= a and not b;
    layer0_outputs(2188) <= a and not b;
    layer0_outputs(2189) <= '1';
    layer0_outputs(2190) <= a or b;
    layer0_outputs(2191) <= not (a and b);
    layer0_outputs(2192) <= '0';
    layer0_outputs(2193) <= not a;
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= a or b;
    layer0_outputs(2196) <= not (a and b);
    layer0_outputs(2197) <= a or b;
    layer0_outputs(2198) <= not (a xor b);
    layer0_outputs(2199) <= a and not b;
    layer0_outputs(2200) <= not (a or b);
    layer0_outputs(2201) <= a and b;
    layer0_outputs(2202) <= not b;
    layer0_outputs(2203) <= not (a and b);
    layer0_outputs(2204) <= not (a and b);
    layer0_outputs(2205) <= b;
    layer0_outputs(2206) <= not a;
    layer0_outputs(2207) <= a and not b;
    layer0_outputs(2208) <= '0';
    layer0_outputs(2209) <= a or b;
    layer0_outputs(2210) <= not (a or b);
    layer0_outputs(2211) <= not (a and b);
    layer0_outputs(2212) <= a;
    layer0_outputs(2213) <= a;
    layer0_outputs(2214) <= b and not a;
    layer0_outputs(2215) <= a and b;
    layer0_outputs(2216) <= b;
    layer0_outputs(2217) <= '1';
    layer0_outputs(2218) <= not (a and b);
    layer0_outputs(2219) <= not b;
    layer0_outputs(2220) <= not b;
    layer0_outputs(2221) <= a and not b;
    layer0_outputs(2222) <= b;
    layer0_outputs(2223) <= a and b;
    layer0_outputs(2224) <= not b;
    layer0_outputs(2225) <= a and not b;
    layer0_outputs(2226) <= a;
    layer0_outputs(2227) <= a and b;
    layer0_outputs(2228) <= '1';
    layer0_outputs(2229) <= not a;
    layer0_outputs(2230) <= b;
    layer0_outputs(2231) <= b and not a;
    layer0_outputs(2232) <= not (a xor b);
    layer0_outputs(2233) <= not b or a;
    layer0_outputs(2234) <= not (a xor b);
    layer0_outputs(2235) <= not a;
    layer0_outputs(2236) <= not (a xor b);
    layer0_outputs(2237) <= not a;
    layer0_outputs(2238) <= not b;
    layer0_outputs(2239) <= b and not a;
    layer0_outputs(2240) <= a and not b;
    layer0_outputs(2241) <= not (a xor b);
    layer0_outputs(2242) <= '1';
    layer0_outputs(2243) <= a xor b;
    layer0_outputs(2244) <= not b;
    layer0_outputs(2245) <= b;
    layer0_outputs(2246) <= not (a xor b);
    layer0_outputs(2247) <= not a or b;
    layer0_outputs(2248) <= not (a and b);
    layer0_outputs(2249) <= not b or a;
    layer0_outputs(2250) <= not (a xor b);
    layer0_outputs(2251) <= not (a or b);
    layer0_outputs(2252) <= '1';
    layer0_outputs(2253) <= '1';
    layer0_outputs(2254) <= b;
    layer0_outputs(2255) <= not (a xor b);
    layer0_outputs(2256) <= b and not a;
    layer0_outputs(2257) <= b;
    layer0_outputs(2258) <= not b or a;
    layer0_outputs(2259) <= a and not b;
    layer0_outputs(2260) <= not a or b;
    layer0_outputs(2261) <= a xor b;
    layer0_outputs(2262) <= a or b;
    layer0_outputs(2263) <= not (a or b);
    layer0_outputs(2264) <= not (a xor b);
    layer0_outputs(2265) <= not b or a;
    layer0_outputs(2266) <= not b;
    layer0_outputs(2267) <= a or b;
    layer0_outputs(2268) <= not a;
    layer0_outputs(2269) <= not (a xor b);
    layer0_outputs(2270) <= not a or b;
    layer0_outputs(2271) <= a or b;
    layer0_outputs(2272) <= a;
    layer0_outputs(2273) <= not a or b;
    layer0_outputs(2274) <= not (a xor b);
    layer0_outputs(2275) <= not b or a;
    layer0_outputs(2276) <= '0';
    layer0_outputs(2277) <= not (a and b);
    layer0_outputs(2278) <= not (a xor b);
    layer0_outputs(2279) <= not (a xor b);
    layer0_outputs(2280) <= not (a and b);
    layer0_outputs(2281) <= a and not b;
    layer0_outputs(2282) <= b and not a;
    layer0_outputs(2283) <= a and not b;
    layer0_outputs(2284) <= not a or b;
    layer0_outputs(2285) <= '1';
    layer0_outputs(2286) <= not b;
    layer0_outputs(2287) <= b;
    layer0_outputs(2288) <= b and not a;
    layer0_outputs(2289) <= not a or b;
    layer0_outputs(2290) <= '1';
    layer0_outputs(2291) <= b;
    layer0_outputs(2292) <= '0';
    layer0_outputs(2293) <= '0';
    layer0_outputs(2294) <= not (a or b);
    layer0_outputs(2295) <= not (a xor b);
    layer0_outputs(2296) <= not a or b;
    layer0_outputs(2297) <= not b or a;
    layer0_outputs(2298) <= b and not a;
    layer0_outputs(2299) <= '1';
    layer0_outputs(2300) <= not b;
    layer0_outputs(2301) <= not (a xor b);
    layer0_outputs(2302) <= not b;
    layer0_outputs(2303) <= not (a xor b);
    layer0_outputs(2304) <= not (a or b);
    layer0_outputs(2305) <= a xor b;
    layer0_outputs(2306) <= a;
    layer0_outputs(2307) <= b and not a;
    layer0_outputs(2308) <= not (a or b);
    layer0_outputs(2309) <= '0';
    layer0_outputs(2310) <= not a or b;
    layer0_outputs(2311) <= not (a or b);
    layer0_outputs(2312) <= a;
    layer0_outputs(2313) <= a or b;
    layer0_outputs(2314) <= not (a or b);
    layer0_outputs(2315) <= not b or a;
    layer0_outputs(2316) <= not (a xor b);
    layer0_outputs(2317) <= not a or b;
    layer0_outputs(2318) <= a xor b;
    layer0_outputs(2319) <= a;
    layer0_outputs(2320) <= not a;
    layer0_outputs(2321) <= a or b;
    layer0_outputs(2322) <= b;
    layer0_outputs(2323) <= not a or b;
    layer0_outputs(2324) <= a and not b;
    layer0_outputs(2325) <= a or b;
    layer0_outputs(2326) <= not b;
    layer0_outputs(2327) <= not (a or b);
    layer0_outputs(2328) <= a and not b;
    layer0_outputs(2329) <= a or b;
    layer0_outputs(2330) <= not (a or b);
    layer0_outputs(2331) <= not (a xor b);
    layer0_outputs(2332) <= a and not b;
    layer0_outputs(2333) <= not (a or b);
    layer0_outputs(2334) <= not (a and b);
    layer0_outputs(2335) <= not b;
    layer0_outputs(2336) <= not b;
    layer0_outputs(2337) <= '1';
    layer0_outputs(2338) <= not b or a;
    layer0_outputs(2339) <= b;
    layer0_outputs(2340) <= not (a xor b);
    layer0_outputs(2341) <= not (a or b);
    layer0_outputs(2342) <= not a;
    layer0_outputs(2343) <= not b;
    layer0_outputs(2344) <= not (a or b);
    layer0_outputs(2345) <= a and not b;
    layer0_outputs(2346) <= a;
    layer0_outputs(2347) <= a;
    layer0_outputs(2348) <= a;
    layer0_outputs(2349) <= a or b;
    layer0_outputs(2350) <= '0';
    layer0_outputs(2351) <= b and not a;
    layer0_outputs(2352) <= not b or a;
    layer0_outputs(2353) <= not (a and b);
    layer0_outputs(2354) <= '1';
    layer0_outputs(2355) <= not (a xor b);
    layer0_outputs(2356) <= not a or b;
    layer0_outputs(2357) <= a;
    layer0_outputs(2358) <= not (a or b);
    layer0_outputs(2359) <= a and not b;
    layer0_outputs(2360) <= b;
    layer0_outputs(2361) <= not a or b;
    layer0_outputs(2362) <= b and not a;
    layer0_outputs(2363) <= b;
    layer0_outputs(2364) <= not b;
    layer0_outputs(2365) <= not a;
    layer0_outputs(2366) <= not (a or b);
    layer0_outputs(2367) <= b and not a;
    layer0_outputs(2368) <= a and b;
    layer0_outputs(2369) <= not a;
    layer0_outputs(2370) <= not b;
    layer0_outputs(2371) <= a;
    layer0_outputs(2372) <= not b or a;
    layer0_outputs(2373) <= not a or b;
    layer0_outputs(2374) <= not b or a;
    layer0_outputs(2375) <= b and not a;
    layer0_outputs(2376) <= a and not b;
    layer0_outputs(2377) <= not a or b;
    layer0_outputs(2378) <= a xor b;
    layer0_outputs(2379) <= a;
    layer0_outputs(2380) <= a xor b;
    layer0_outputs(2381) <= a and not b;
    layer0_outputs(2382) <= '0';
    layer0_outputs(2383) <= b;
    layer0_outputs(2384) <= not (a xor b);
    layer0_outputs(2385) <= a;
    layer0_outputs(2386) <= not (a xor b);
    layer0_outputs(2387) <= a or b;
    layer0_outputs(2388) <= '0';
    layer0_outputs(2389) <= a or b;
    layer0_outputs(2390) <= not (a and b);
    layer0_outputs(2391) <= b;
    layer0_outputs(2392) <= a and not b;
    layer0_outputs(2393) <= a or b;
    layer0_outputs(2394) <= b;
    layer0_outputs(2395) <= a and not b;
    layer0_outputs(2396) <= '0';
    layer0_outputs(2397) <= a or b;
    layer0_outputs(2398) <= not (a and b);
    layer0_outputs(2399) <= b;
    layer0_outputs(2400) <= a or b;
    layer0_outputs(2401) <= not a or b;
    layer0_outputs(2402) <= a xor b;
    layer0_outputs(2403) <= not a;
    layer0_outputs(2404) <= not (a or b);
    layer0_outputs(2405) <= '0';
    layer0_outputs(2406) <= a;
    layer0_outputs(2407) <= b and not a;
    layer0_outputs(2408) <= a and not b;
    layer0_outputs(2409) <= a or b;
    layer0_outputs(2410) <= not b or a;
    layer0_outputs(2411) <= not b;
    layer0_outputs(2412) <= b and not a;
    layer0_outputs(2413) <= not b or a;
    layer0_outputs(2414) <= not (a xor b);
    layer0_outputs(2415) <= a and not b;
    layer0_outputs(2416) <= '1';
    layer0_outputs(2417) <= b;
    layer0_outputs(2418) <= a and not b;
    layer0_outputs(2419) <= b and not a;
    layer0_outputs(2420) <= b and not a;
    layer0_outputs(2421) <= not b or a;
    layer0_outputs(2422) <= not a;
    layer0_outputs(2423) <= '0';
    layer0_outputs(2424) <= b;
    layer0_outputs(2425) <= b and not a;
    layer0_outputs(2426) <= b;
    layer0_outputs(2427) <= a or b;
    layer0_outputs(2428) <= a xor b;
    layer0_outputs(2429) <= a;
    layer0_outputs(2430) <= b;
    layer0_outputs(2431) <= not a or b;
    layer0_outputs(2432) <= b;
    layer0_outputs(2433) <= b and not a;
    layer0_outputs(2434) <= a and not b;
    layer0_outputs(2435) <= not a;
    layer0_outputs(2436) <= a;
    layer0_outputs(2437) <= a or b;
    layer0_outputs(2438) <= a or b;
    layer0_outputs(2439) <= not b;
    layer0_outputs(2440) <= not (a and b);
    layer0_outputs(2441) <= not a;
    layer0_outputs(2442) <= a or b;
    layer0_outputs(2443) <= b;
    layer0_outputs(2444) <= not (a xor b);
    layer0_outputs(2445) <= not (a or b);
    layer0_outputs(2446) <= a;
    layer0_outputs(2447) <= not (a and b);
    layer0_outputs(2448) <= not a or b;
    layer0_outputs(2449) <= b and not a;
    layer0_outputs(2450) <= a;
    layer0_outputs(2451) <= b and not a;
    layer0_outputs(2452) <= b;
    layer0_outputs(2453) <= not (a and b);
    layer0_outputs(2454) <= a;
    layer0_outputs(2455) <= a or b;
    layer0_outputs(2456) <= not (a or b);
    layer0_outputs(2457) <= b and not a;
    layer0_outputs(2458) <= not (a xor b);
    layer0_outputs(2459) <= not (a or b);
    layer0_outputs(2460) <= not a;
    layer0_outputs(2461) <= a;
    layer0_outputs(2462) <= a or b;
    layer0_outputs(2463) <= not b;
    layer0_outputs(2464) <= not a;
    layer0_outputs(2465) <= not (a xor b);
    layer0_outputs(2466) <= not (a and b);
    layer0_outputs(2467) <= a and not b;
    layer0_outputs(2468) <= not (a or b);
    layer0_outputs(2469) <= a xor b;
    layer0_outputs(2470) <= '0';
    layer0_outputs(2471) <= not (a xor b);
    layer0_outputs(2472) <= b;
    layer0_outputs(2473) <= not a;
    layer0_outputs(2474) <= not a;
    layer0_outputs(2475) <= a;
    layer0_outputs(2476) <= a;
    layer0_outputs(2477) <= b;
    layer0_outputs(2478) <= not a;
    layer0_outputs(2479) <= a and not b;
    layer0_outputs(2480) <= not b;
    layer0_outputs(2481) <= b;
    layer0_outputs(2482) <= a xor b;
    layer0_outputs(2483) <= '1';
    layer0_outputs(2484) <= a and b;
    layer0_outputs(2485) <= not (a or b);
    layer0_outputs(2486) <= b;
    layer0_outputs(2487) <= a or b;
    layer0_outputs(2488) <= not b;
    layer0_outputs(2489) <= not (a xor b);
    layer0_outputs(2490) <= not (a xor b);
    layer0_outputs(2491) <= not a;
    layer0_outputs(2492) <= '0';
    layer0_outputs(2493) <= '0';
    layer0_outputs(2494) <= a and b;
    layer0_outputs(2495) <= not (a or b);
    layer0_outputs(2496) <= a xor b;
    layer0_outputs(2497) <= a xor b;
    layer0_outputs(2498) <= a or b;
    layer0_outputs(2499) <= not b;
    layer0_outputs(2500) <= not a or b;
    layer0_outputs(2501) <= a;
    layer0_outputs(2502) <= '1';
    layer0_outputs(2503) <= not (a xor b);
    layer0_outputs(2504) <= a or b;
    layer0_outputs(2505) <= not (a xor b);
    layer0_outputs(2506) <= not a or b;
    layer0_outputs(2507) <= not (a or b);
    layer0_outputs(2508) <= not b;
    layer0_outputs(2509) <= not b or a;
    layer0_outputs(2510) <= '0';
    layer0_outputs(2511) <= '0';
    layer0_outputs(2512) <= a or b;
    layer0_outputs(2513) <= not a;
    layer0_outputs(2514) <= '0';
    layer0_outputs(2515) <= not b or a;
    layer0_outputs(2516) <= a or b;
    layer0_outputs(2517) <= a xor b;
    layer0_outputs(2518) <= b and not a;
    layer0_outputs(2519) <= a and not b;
    layer0_outputs(2520) <= not b;
    layer0_outputs(2521) <= b and not a;
    layer0_outputs(2522) <= b and not a;
    layer0_outputs(2523) <= not a;
    layer0_outputs(2524) <= not (a xor b);
    layer0_outputs(2525) <= not b;
    layer0_outputs(2526) <= a and b;
    layer0_outputs(2527) <= b;
    layer0_outputs(2528) <= '1';
    layer0_outputs(2529) <= a;
    layer0_outputs(2530) <= a;
    layer0_outputs(2531) <= not a or b;
    layer0_outputs(2532) <= not (a or b);
    layer0_outputs(2533) <= not (a xor b);
    layer0_outputs(2534) <= '0';
    layer0_outputs(2535) <= not a;
    layer0_outputs(2536) <= not b or a;
    layer0_outputs(2537) <= not b;
    layer0_outputs(2538) <= a or b;
    layer0_outputs(2539) <= b;
    layer0_outputs(2540) <= not (a and b);
    layer0_outputs(2541) <= a xor b;
    layer0_outputs(2542) <= not a;
    layer0_outputs(2543) <= a and not b;
    layer0_outputs(2544) <= not (a xor b);
    layer0_outputs(2545) <= a;
    layer0_outputs(2546) <= not a;
    layer0_outputs(2547) <= a and b;
    layer0_outputs(2548) <= not (a or b);
    layer0_outputs(2549) <= b;
    layer0_outputs(2550) <= not a;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= b and not a;
    layer0_outputs(2553) <= a;
    layer0_outputs(2554) <= b;
    layer0_outputs(2555) <= a;
    layer0_outputs(2556) <= '1';
    layer0_outputs(2557) <= '0';
    layer0_outputs(2558) <= not a or b;
    layer0_outputs(2559) <= b;
    layer0_outputs(2560) <= not a;
    layer0_outputs(2561) <= a and not b;
    layer0_outputs(2562) <= not b;
    layer0_outputs(2563) <= b;
    layer0_outputs(2564) <= a;
    layer0_outputs(2565) <= a and not b;
    layer0_outputs(2566) <= a;
    layer0_outputs(2567) <= b and not a;
    layer0_outputs(2568) <= not b or a;
    layer0_outputs(2569) <= a or b;
    layer0_outputs(2570) <= a and b;
    layer0_outputs(2571) <= a and b;
    layer0_outputs(2572) <= not b or a;
    layer0_outputs(2573) <= a and b;
    layer0_outputs(2574) <= not (a xor b);
    layer0_outputs(2575) <= a or b;
    layer0_outputs(2576) <= a and not b;
    layer0_outputs(2577) <= b;
    layer0_outputs(2578) <= not b or a;
    layer0_outputs(2579) <= a xor b;
    layer0_outputs(2580) <= not a;
    layer0_outputs(2581) <= '0';
    layer0_outputs(2582) <= not (a or b);
    layer0_outputs(2583) <= a and not b;
    layer0_outputs(2584) <= '0';
    layer0_outputs(2585) <= not (a or b);
    layer0_outputs(2586) <= not (a or b);
    layer0_outputs(2587) <= not (a and b);
    layer0_outputs(2588) <= a;
    layer0_outputs(2589) <= not b;
    layer0_outputs(2590) <= a;
    layer0_outputs(2591) <= '0';
    layer0_outputs(2592) <= not b or a;
    layer0_outputs(2593) <= a or b;
    layer0_outputs(2594) <= a or b;
    layer0_outputs(2595) <= a and b;
    layer0_outputs(2596) <= not (a or b);
    layer0_outputs(2597) <= not b;
    layer0_outputs(2598) <= '1';
    layer0_outputs(2599) <= b and not a;
    layer0_outputs(2600) <= '0';
    layer0_outputs(2601) <= a xor b;
    layer0_outputs(2602) <= b and not a;
    layer0_outputs(2603) <= not (a and b);
    layer0_outputs(2604) <= not a;
    layer0_outputs(2605) <= not (a or b);
    layer0_outputs(2606) <= not (a or b);
    layer0_outputs(2607) <= a;
    layer0_outputs(2608) <= not b;
    layer0_outputs(2609) <= a;
    layer0_outputs(2610) <= a and b;
    layer0_outputs(2611) <= b and not a;
    layer0_outputs(2612) <= b and not a;
    layer0_outputs(2613) <= not (a and b);
    layer0_outputs(2614) <= not (a xor b);
    layer0_outputs(2615) <= a and not b;
    layer0_outputs(2616) <= not (a or b);
    layer0_outputs(2617) <= not a;
    layer0_outputs(2618) <= a and b;
    layer0_outputs(2619) <= a;
    layer0_outputs(2620) <= not a or b;
    layer0_outputs(2621) <= not a;
    layer0_outputs(2622) <= not b or a;
    layer0_outputs(2623) <= b;
    layer0_outputs(2624) <= not a;
    layer0_outputs(2625) <= b;
    layer0_outputs(2626) <= not b or a;
    layer0_outputs(2627) <= a and not b;
    layer0_outputs(2628) <= a xor b;
    layer0_outputs(2629) <= a xor b;
    layer0_outputs(2630) <= not b or a;
    layer0_outputs(2631) <= a and b;
    layer0_outputs(2632) <= a and not b;
    layer0_outputs(2633) <= not a;
    layer0_outputs(2634) <= a xor b;
    layer0_outputs(2635) <= not b;
    layer0_outputs(2636) <= not a;
    layer0_outputs(2637) <= not a;
    layer0_outputs(2638) <= b;
    layer0_outputs(2639) <= not a;
    layer0_outputs(2640) <= a and not b;
    layer0_outputs(2641) <= a and not b;
    layer0_outputs(2642) <= not (a and b);
    layer0_outputs(2643) <= a and b;
    layer0_outputs(2644) <= a;
    layer0_outputs(2645) <= a and b;
    layer0_outputs(2646) <= b and not a;
    layer0_outputs(2647) <= not b or a;
    layer0_outputs(2648) <= not b or a;
    layer0_outputs(2649) <= b;
    layer0_outputs(2650) <= a;
    layer0_outputs(2651) <= '1';
    layer0_outputs(2652) <= not b;
    layer0_outputs(2653) <= a or b;
    layer0_outputs(2654) <= a;
    layer0_outputs(2655) <= not a or b;
    layer0_outputs(2656) <= not a;
    layer0_outputs(2657) <= b and not a;
    layer0_outputs(2658) <= '1';
    layer0_outputs(2659) <= b;
    layer0_outputs(2660) <= a or b;
    layer0_outputs(2661) <= not b;
    layer0_outputs(2662) <= not a;
    layer0_outputs(2663) <= not b or a;
    layer0_outputs(2664) <= b and not a;
    layer0_outputs(2665) <= not a;
    layer0_outputs(2666) <= a;
    layer0_outputs(2667) <= not (a and b);
    layer0_outputs(2668) <= b and not a;
    layer0_outputs(2669) <= not (a or b);
    layer0_outputs(2670) <= not b;
    layer0_outputs(2671) <= not (a or b);
    layer0_outputs(2672) <= b;
    layer0_outputs(2673) <= b;
    layer0_outputs(2674) <= not a or b;
    layer0_outputs(2675) <= not a;
    layer0_outputs(2676) <= not a;
    layer0_outputs(2677) <= not (a xor b);
    layer0_outputs(2678) <= a and not b;
    layer0_outputs(2679) <= not a or b;
    layer0_outputs(2680) <= not (a xor b);
    layer0_outputs(2681) <= not (a xor b);
    layer0_outputs(2682) <= b;
    layer0_outputs(2683) <= not (a xor b);
    layer0_outputs(2684) <= not b;
    layer0_outputs(2685) <= a xor b;
    layer0_outputs(2686) <= a xor b;
    layer0_outputs(2687) <= not (a or b);
    layer0_outputs(2688) <= '0';
    layer0_outputs(2689) <= a xor b;
    layer0_outputs(2690) <= not (a xor b);
    layer0_outputs(2691) <= b;
    layer0_outputs(2692) <= a and not b;
    layer0_outputs(2693) <= a or b;
    layer0_outputs(2694) <= not a or b;
    layer0_outputs(2695) <= not (a xor b);
    layer0_outputs(2696) <= not a;
    layer0_outputs(2697) <= '1';
    layer0_outputs(2698) <= not b;
    layer0_outputs(2699) <= a or b;
    layer0_outputs(2700) <= a or b;
    layer0_outputs(2701) <= b;
    layer0_outputs(2702) <= b;
    layer0_outputs(2703) <= '1';
    layer0_outputs(2704) <= not a or b;
    layer0_outputs(2705) <= b and not a;
    layer0_outputs(2706) <= not (a or b);
    layer0_outputs(2707) <= a and not b;
    layer0_outputs(2708) <= not a;
    layer0_outputs(2709) <= not (a and b);
    layer0_outputs(2710) <= '0';
    layer0_outputs(2711) <= a xor b;
    layer0_outputs(2712) <= a and not b;
    layer0_outputs(2713) <= not a;
    layer0_outputs(2714) <= '0';
    layer0_outputs(2715) <= b;
    layer0_outputs(2716) <= b and not a;
    layer0_outputs(2717) <= a xor b;
    layer0_outputs(2718) <= '0';
    layer0_outputs(2719) <= a or b;
    layer0_outputs(2720) <= a or b;
    layer0_outputs(2721) <= a;
    layer0_outputs(2722) <= not a;
    layer0_outputs(2723) <= not b;
    layer0_outputs(2724) <= a;
    layer0_outputs(2725) <= not (a or b);
    layer0_outputs(2726) <= b;
    layer0_outputs(2727) <= not (a xor b);
    layer0_outputs(2728) <= a and b;
    layer0_outputs(2729) <= not (a or b);
    layer0_outputs(2730) <= b;
    layer0_outputs(2731) <= not (a xor b);
    layer0_outputs(2732) <= not a or b;
    layer0_outputs(2733) <= not (a xor b);
    layer0_outputs(2734) <= not (a or b);
    layer0_outputs(2735) <= b;
    layer0_outputs(2736) <= '0';
    layer0_outputs(2737) <= not (a or b);
    layer0_outputs(2738) <= not (a or b);
    layer0_outputs(2739) <= a and b;
    layer0_outputs(2740) <= not b or a;
    layer0_outputs(2741) <= not a or b;
    layer0_outputs(2742) <= not b;
    layer0_outputs(2743) <= '1';
    layer0_outputs(2744) <= not a;
    layer0_outputs(2745) <= a or b;
    layer0_outputs(2746) <= '1';
    layer0_outputs(2747) <= not a;
    layer0_outputs(2748) <= '1';
    layer0_outputs(2749) <= not b;
    layer0_outputs(2750) <= not (a and b);
    layer0_outputs(2751) <= not (a xor b);
    layer0_outputs(2752) <= a xor b;
    layer0_outputs(2753) <= '1';
    layer0_outputs(2754) <= a or b;
    layer0_outputs(2755) <= b and not a;
    layer0_outputs(2756) <= not (a xor b);
    layer0_outputs(2757) <= a;
    layer0_outputs(2758) <= a and not b;
    layer0_outputs(2759) <= a xor b;
    layer0_outputs(2760) <= '0';
    layer0_outputs(2761) <= a;
    layer0_outputs(2762) <= a or b;
    layer0_outputs(2763) <= not (a and b);
    layer0_outputs(2764) <= a;
    layer0_outputs(2765) <= not a or b;
    layer0_outputs(2766) <= a or b;
    layer0_outputs(2767) <= a and not b;
    layer0_outputs(2768) <= a;
    layer0_outputs(2769) <= b;
    layer0_outputs(2770) <= not (a and b);
    layer0_outputs(2771) <= not b;
    layer0_outputs(2772) <= a and b;
    layer0_outputs(2773) <= not (a xor b);
    layer0_outputs(2774) <= not b or a;
    layer0_outputs(2775) <= not a;
    layer0_outputs(2776) <= not a or b;
    layer0_outputs(2777) <= not (a or b);
    layer0_outputs(2778) <= a or b;
    layer0_outputs(2779) <= not (a and b);
    layer0_outputs(2780) <= a and not b;
    layer0_outputs(2781) <= '0';
    layer0_outputs(2782) <= a and b;
    layer0_outputs(2783) <= b and not a;
    layer0_outputs(2784) <= '1';
    layer0_outputs(2785) <= not a;
    layer0_outputs(2786) <= not a or b;
    layer0_outputs(2787) <= not (a and b);
    layer0_outputs(2788) <= b and not a;
    layer0_outputs(2789) <= a xor b;
    layer0_outputs(2790) <= not (a and b);
    layer0_outputs(2791) <= a or b;
    layer0_outputs(2792) <= a and b;
    layer0_outputs(2793) <= not (a xor b);
    layer0_outputs(2794) <= not a;
    layer0_outputs(2795) <= a;
    layer0_outputs(2796) <= a and b;
    layer0_outputs(2797) <= not b;
    layer0_outputs(2798) <= a or b;
    layer0_outputs(2799) <= not a;
    layer0_outputs(2800) <= not (a xor b);
    layer0_outputs(2801) <= not a;
    layer0_outputs(2802) <= a and b;
    layer0_outputs(2803) <= not (a xor b);
    layer0_outputs(2804) <= '1';
    layer0_outputs(2805) <= b;
    layer0_outputs(2806) <= a or b;
    layer0_outputs(2807) <= not b;
    layer0_outputs(2808) <= not (a and b);
    layer0_outputs(2809) <= '0';
    layer0_outputs(2810) <= not b;
    layer0_outputs(2811) <= b and not a;
    layer0_outputs(2812) <= b and not a;
    layer0_outputs(2813) <= '1';
    layer0_outputs(2814) <= b;
    layer0_outputs(2815) <= not a or b;
    layer0_outputs(2816) <= a and b;
    layer0_outputs(2817) <= b;
    layer0_outputs(2818) <= a xor b;
    layer0_outputs(2819) <= b and not a;
    layer0_outputs(2820) <= not a;
    layer0_outputs(2821) <= not a or b;
    layer0_outputs(2822) <= a and b;
    layer0_outputs(2823) <= not b;
    layer0_outputs(2824) <= a and b;
    layer0_outputs(2825) <= '0';
    layer0_outputs(2826) <= b;
    layer0_outputs(2827) <= a and b;
    layer0_outputs(2828) <= a and not b;
    layer0_outputs(2829) <= '0';
    layer0_outputs(2830) <= not b;
    layer0_outputs(2831) <= not b or a;
    layer0_outputs(2832) <= not a or b;
    layer0_outputs(2833) <= not b or a;
    layer0_outputs(2834) <= not b;
    layer0_outputs(2835) <= '0';
    layer0_outputs(2836) <= b and not a;
    layer0_outputs(2837) <= not (a xor b);
    layer0_outputs(2838) <= not (a and b);
    layer0_outputs(2839) <= a or b;
    layer0_outputs(2840) <= a and b;
    layer0_outputs(2841) <= not b or a;
    layer0_outputs(2842) <= not (a or b);
    layer0_outputs(2843) <= a;
    layer0_outputs(2844) <= a;
    layer0_outputs(2845) <= not (a or b);
    layer0_outputs(2846) <= a xor b;
    layer0_outputs(2847) <= a xor b;
    layer0_outputs(2848) <= not a;
    layer0_outputs(2849) <= a or b;
    layer0_outputs(2850) <= '1';
    layer0_outputs(2851) <= b and not a;
    layer0_outputs(2852) <= not (a or b);
    layer0_outputs(2853) <= '1';
    layer0_outputs(2854) <= not a or b;
    layer0_outputs(2855) <= a and not b;
    layer0_outputs(2856) <= a and not b;
    layer0_outputs(2857) <= not (a or b);
    layer0_outputs(2858) <= not a or b;
    layer0_outputs(2859) <= b;
    layer0_outputs(2860) <= a and not b;
    layer0_outputs(2861) <= a xor b;
    layer0_outputs(2862) <= b and not a;
    layer0_outputs(2863) <= '0';
    layer0_outputs(2864) <= '0';
    layer0_outputs(2865) <= a xor b;
    layer0_outputs(2866) <= a;
    layer0_outputs(2867) <= b;
    layer0_outputs(2868) <= not a;
    layer0_outputs(2869) <= not (a or b);
    layer0_outputs(2870) <= b and not a;
    layer0_outputs(2871) <= not b or a;
    layer0_outputs(2872) <= a or b;
    layer0_outputs(2873) <= not (a xor b);
    layer0_outputs(2874) <= a or b;
    layer0_outputs(2875) <= not a;
    layer0_outputs(2876) <= a or b;
    layer0_outputs(2877) <= not b or a;
    layer0_outputs(2878) <= not b;
    layer0_outputs(2879) <= not b;
    layer0_outputs(2880) <= a;
    layer0_outputs(2881) <= '0';
    layer0_outputs(2882) <= not a;
    layer0_outputs(2883) <= not a or b;
    layer0_outputs(2884) <= not (a xor b);
    layer0_outputs(2885) <= a and not b;
    layer0_outputs(2886) <= a or b;
    layer0_outputs(2887) <= b;
    layer0_outputs(2888) <= a or b;
    layer0_outputs(2889) <= a xor b;
    layer0_outputs(2890) <= not b;
    layer0_outputs(2891) <= b;
    layer0_outputs(2892) <= not (a xor b);
    layer0_outputs(2893) <= a or b;
    layer0_outputs(2894) <= not (a xor b);
    layer0_outputs(2895) <= not (a or b);
    layer0_outputs(2896) <= not b or a;
    layer0_outputs(2897) <= a and not b;
    layer0_outputs(2898) <= b;
    layer0_outputs(2899) <= a and not b;
    layer0_outputs(2900) <= not b or a;
    layer0_outputs(2901) <= a or b;
    layer0_outputs(2902) <= not (a or b);
    layer0_outputs(2903) <= not (a or b);
    layer0_outputs(2904) <= not b or a;
    layer0_outputs(2905) <= b;
    layer0_outputs(2906) <= a and b;
    layer0_outputs(2907) <= not b or a;
    layer0_outputs(2908) <= not (a and b);
    layer0_outputs(2909) <= not b;
    layer0_outputs(2910) <= not b;
    layer0_outputs(2911) <= not b;
    layer0_outputs(2912) <= not a;
    layer0_outputs(2913) <= not (a xor b);
    layer0_outputs(2914) <= not a or b;
    layer0_outputs(2915) <= not (a xor b);
    layer0_outputs(2916) <= a and b;
    layer0_outputs(2917) <= not b;
    layer0_outputs(2918) <= '0';
    layer0_outputs(2919) <= a and not b;
    layer0_outputs(2920) <= a and b;
    layer0_outputs(2921) <= a or b;
    layer0_outputs(2922) <= a xor b;
    layer0_outputs(2923) <= not a;
    layer0_outputs(2924) <= b and not a;
    layer0_outputs(2925) <= a and b;
    layer0_outputs(2926) <= not (a or b);
    layer0_outputs(2927) <= not (a and b);
    layer0_outputs(2928) <= not a or b;
    layer0_outputs(2929) <= a;
    layer0_outputs(2930) <= not b or a;
    layer0_outputs(2931) <= a or b;
    layer0_outputs(2932) <= not a or b;
    layer0_outputs(2933) <= not a or b;
    layer0_outputs(2934) <= a and b;
    layer0_outputs(2935) <= not (a or b);
    layer0_outputs(2936) <= not (a or b);
    layer0_outputs(2937) <= b;
    layer0_outputs(2938) <= not b;
    layer0_outputs(2939) <= not b or a;
    layer0_outputs(2940) <= a or b;
    layer0_outputs(2941) <= not (a and b);
    layer0_outputs(2942) <= not a or b;
    layer0_outputs(2943) <= b;
    layer0_outputs(2944) <= a;
    layer0_outputs(2945) <= a and b;
    layer0_outputs(2946) <= not a or b;
    layer0_outputs(2947) <= not b;
    layer0_outputs(2948) <= not b or a;
    layer0_outputs(2949) <= b;
    layer0_outputs(2950) <= a;
    layer0_outputs(2951) <= not (a or b);
    layer0_outputs(2952) <= b and not a;
    layer0_outputs(2953) <= not (a or b);
    layer0_outputs(2954) <= not (a xor b);
    layer0_outputs(2955) <= not (a xor b);
    layer0_outputs(2956) <= not (a and b);
    layer0_outputs(2957) <= b;
    layer0_outputs(2958) <= '0';
    layer0_outputs(2959) <= not (a or b);
    layer0_outputs(2960) <= not a or b;
    layer0_outputs(2961) <= a or b;
    layer0_outputs(2962) <= '1';
    layer0_outputs(2963) <= a and b;
    layer0_outputs(2964) <= a xor b;
    layer0_outputs(2965) <= not b or a;
    layer0_outputs(2966) <= b and not a;
    layer0_outputs(2967) <= not a or b;
    layer0_outputs(2968) <= a or b;
    layer0_outputs(2969) <= '1';
    layer0_outputs(2970) <= not a or b;
    layer0_outputs(2971) <= a xor b;
    layer0_outputs(2972) <= not b;
    layer0_outputs(2973) <= a and not b;
    layer0_outputs(2974) <= not (a or b);
    layer0_outputs(2975) <= '1';
    layer0_outputs(2976) <= not (a xor b);
    layer0_outputs(2977) <= a and b;
    layer0_outputs(2978) <= a xor b;
    layer0_outputs(2979) <= a;
    layer0_outputs(2980) <= not b or a;
    layer0_outputs(2981) <= not b;
    layer0_outputs(2982) <= not (a or b);
    layer0_outputs(2983) <= b;
    layer0_outputs(2984) <= not b or a;
    layer0_outputs(2985) <= a and not b;
    layer0_outputs(2986) <= '0';
    layer0_outputs(2987) <= '0';
    layer0_outputs(2988) <= b and not a;
    layer0_outputs(2989) <= not b or a;
    layer0_outputs(2990) <= not b;
    layer0_outputs(2991) <= not a or b;
    layer0_outputs(2992) <= a xor b;
    layer0_outputs(2993) <= b;
    layer0_outputs(2994) <= not (a or b);
    layer0_outputs(2995) <= not (a xor b);
    layer0_outputs(2996) <= b;
    layer0_outputs(2997) <= '1';
    layer0_outputs(2998) <= '0';
    layer0_outputs(2999) <= not b or a;
    layer0_outputs(3000) <= a;
    layer0_outputs(3001) <= a;
    layer0_outputs(3002) <= a and b;
    layer0_outputs(3003) <= not (a or b);
    layer0_outputs(3004) <= a;
    layer0_outputs(3005) <= not (a xor b);
    layer0_outputs(3006) <= a or b;
    layer0_outputs(3007) <= '0';
    layer0_outputs(3008) <= not a;
    layer0_outputs(3009) <= a xor b;
    layer0_outputs(3010) <= not (a and b);
    layer0_outputs(3011) <= a and not b;
    layer0_outputs(3012) <= a xor b;
    layer0_outputs(3013) <= b and not a;
    layer0_outputs(3014) <= '1';
    layer0_outputs(3015) <= not b or a;
    layer0_outputs(3016) <= a and not b;
    layer0_outputs(3017) <= not a or b;
    layer0_outputs(3018) <= not (a xor b);
    layer0_outputs(3019) <= not b;
    layer0_outputs(3020) <= not a;
    layer0_outputs(3021) <= a;
    layer0_outputs(3022) <= not (a and b);
    layer0_outputs(3023) <= not b;
    layer0_outputs(3024) <= not a;
    layer0_outputs(3025) <= b and not a;
    layer0_outputs(3026) <= '1';
    layer0_outputs(3027) <= a or b;
    layer0_outputs(3028) <= b and not a;
    layer0_outputs(3029) <= a and not b;
    layer0_outputs(3030) <= a xor b;
    layer0_outputs(3031) <= b and not a;
    layer0_outputs(3032) <= not b or a;
    layer0_outputs(3033) <= b and not a;
    layer0_outputs(3034) <= not b;
    layer0_outputs(3035) <= b;
    layer0_outputs(3036) <= b;
    layer0_outputs(3037) <= not (a xor b);
    layer0_outputs(3038) <= a;
    layer0_outputs(3039) <= not a or b;
    layer0_outputs(3040) <= not b;
    layer0_outputs(3041) <= '1';
    layer0_outputs(3042) <= not b or a;
    layer0_outputs(3043) <= '0';
    layer0_outputs(3044) <= b and not a;
    layer0_outputs(3045) <= '0';
    layer0_outputs(3046) <= not (a and b);
    layer0_outputs(3047) <= a xor b;
    layer0_outputs(3048) <= a or b;
    layer0_outputs(3049) <= not a;
    layer0_outputs(3050) <= not a;
    layer0_outputs(3051) <= not a or b;
    layer0_outputs(3052) <= a xor b;
    layer0_outputs(3053) <= not b or a;
    layer0_outputs(3054) <= not (a or b);
    layer0_outputs(3055) <= not (a and b);
    layer0_outputs(3056) <= a and b;
    layer0_outputs(3057) <= not a or b;
    layer0_outputs(3058) <= a;
    layer0_outputs(3059) <= a;
    layer0_outputs(3060) <= not (a or b);
    layer0_outputs(3061) <= a and not b;
    layer0_outputs(3062) <= not a or b;
    layer0_outputs(3063) <= not b or a;
    layer0_outputs(3064) <= not a or b;
    layer0_outputs(3065) <= b;
    layer0_outputs(3066) <= not b;
    layer0_outputs(3067) <= a and b;
    layer0_outputs(3068) <= a or b;
    layer0_outputs(3069) <= b and not a;
    layer0_outputs(3070) <= a or b;
    layer0_outputs(3071) <= not (a or b);
    layer0_outputs(3072) <= b and not a;
    layer0_outputs(3073) <= not a or b;
    layer0_outputs(3074) <= b;
    layer0_outputs(3075) <= a and b;
    layer0_outputs(3076) <= a;
    layer0_outputs(3077) <= not a or b;
    layer0_outputs(3078) <= not b or a;
    layer0_outputs(3079) <= '0';
    layer0_outputs(3080) <= '0';
    layer0_outputs(3081) <= '1';
    layer0_outputs(3082) <= not a;
    layer0_outputs(3083) <= a and b;
    layer0_outputs(3084) <= b;
    layer0_outputs(3085) <= a or b;
    layer0_outputs(3086) <= not a;
    layer0_outputs(3087) <= not b;
    layer0_outputs(3088) <= a;
    layer0_outputs(3089) <= a and not b;
    layer0_outputs(3090) <= a xor b;
    layer0_outputs(3091) <= not b;
    layer0_outputs(3092) <= not a or b;
    layer0_outputs(3093) <= not b or a;
    layer0_outputs(3094) <= a and b;
    layer0_outputs(3095) <= a or b;
    layer0_outputs(3096) <= not (a or b);
    layer0_outputs(3097) <= '0';
    layer0_outputs(3098) <= a and not b;
    layer0_outputs(3099) <= '1';
    layer0_outputs(3100) <= a or b;
    layer0_outputs(3101) <= a and not b;
    layer0_outputs(3102) <= a xor b;
    layer0_outputs(3103) <= not b or a;
    layer0_outputs(3104) <= a;
    layer0_outputs(3105) <= a or b;
    layer0_outputs(3106) <= a or b;
    layer0_outputs(3107) <= b and not a;
    layer0_outputs(3108) <= b;
    layer0_outputs(3109) <= b;
    layer0_outputs(3110) <= a xor b;
    layer0_outputs(3111) <= a and not b;
    layer0_outputs(3112) <= a and not b;
    layer0_outputs(3113) <= not (a xor b);
    layer0_outputs(3114) <= a or b;
    layer0_outputs(3115) <= not (a or b);
    layer0_outputs(3116) <= b;
    layer0_outputs(3117) <= not a;
    layer0_outputs(3118) <= a and not b;
    layer0_outputs(3119) <= a and b;
    layer0_outputs(3120) <= a or b;
    layer0_outputs(3121) <= a or b;
    layer0_outputs(3122) <= '0';
    layer0_outputs(3123) <= not b;
    layer0_outputs(3124) <= a and not b;
    layer0_outputs(3125) <= a or b;
    layer0_outputs(3126) <= a xor b;
    layer0_outputs(3127) <= a and not b;
    layer0_outputs(3128) <= b and not a;
    layer0_outputs(3129) <= a xor b;
    layer0_outputs(3130) <= '1';
    layer0_outputs(3131) <= not b;
    layer0_outputs(3132) <= b and not a;
    layer0_outputs(3133) <= a;
    layer0_outputs(3134) <= a or b;
    layer0_outputs(3135) <= b and not a;
    layer0_outputs(3136) <= not a;
    layer0_outputs(3137) <= not a or b;
    layer0_outputs(3138) <= a and not b;
    layer0_outputs(3139) <= a and b;
    layer0_outputs(3140) <= not (a or b);
    layer0_outputs(3141) <= '0';
    layer0_outputs(3142) <= not b;
    layer0_outputs(3143) <= not (a or b);
    layer0_outputs(3144) <= a or b;
    layer0_outputs(3145) <= '0';
    layer0_outputs(3146) <= not b or a;
    layer0_outputs(3147) <= not b;
    layer0_outputs(3148) <= not b or a;
    layer0_outputs(3149) <= '1';
    layer0_outputs(3150) <= b;
    layer0_outputs(3151) <= a;
    layer0_outputs(3152) <= not b;
    layer0_outputs(3153) <= a xor b;
    layer0_outputs(3154) <= not a;
    layer0_outputs(3155) <= '0';
    layer0_outputs(3156) <= b and not a;
    layer0_outputs(3157) <= not b;
    layer0_outputs(3158) <= '0';
    layer0_outputs(3159) <= not b or a;
    layer0_outputs(3160) <= not b or a;
    layer0_outputs(3161) <= not (a or b);
    layer0_outputs(3162) <= not b;
    layer0_outputs(3163) <= '0';
    layer0_outputs(3164) <= '1';
    layer0_outputs(3165) <= '1';
    layer0_outputs(3166) <= not a;
    layer0_outputs(3167) <= a and not b;
    layer0_outputs(3168) <= '0';
    layer0_outputs(3169) <= not b;
    layer0_outputs(3170) <= a or b;
    layer0_outputs(3171) <= not b or a;
    layer0_outputs(3172) <= not b;
    layer0_outputs(3173) <= not a;
    layer0_outputs(3174) <= '0';
    layer0_outputs(3175) <= not a or b;
    layer0_outputs(3176) <= not (a xor b);
    layer0_outputs(3177) <= not b or a;
    layer0_outputs(3178) <= a or b;
    layer0_outputs(3179) <= not b or a;
    layer0_outputs(3180) <= not a or b;
    layer0_outputs(3181) <= b and not a;
    layer0_outputs(3182) <= not b or a;
    layer0_outputs(3183) <= a or b;
    layer0_outputs(3184) <= a and b;
    layer0_outputs(3185) <= '0';
    layer0_outputs(3186) <= a;
    layer0_outputs(3187) <= not (a and b);
    layer0_outputs(3188) <= not b;
    layer0_outputs(3189) <= b;
    layer0_outputs(3190) <= not b or a;
    layer0_outputs(3191) <= '1';
    layer0_outputs(3192) <= '1';
    layer0_outputs(3193) <= not b;
    layer0_outputs(3194) <= a or b;
    layer0_outputs(3195) <= a or b;
    layer0_outputs(3196) <= not b or a;
    layer0_outputs(3197) <= a or b;
    layer0_outputs(3198) <= '1';
    layer0_outputs(3199) <= a or b;
    layer0_outputs(3200) <= '1';
    layer0_outputs(3201) <= not b;
    layer0_outputs(3202) <= not b;
    layer0_outputs(3203) <= not (a or b);
    layer0_outputs(3204) <= '1';
    layer0_outputs(3205) <= not b or a;
    layer0_outputs(3206) <= not (a or b);
    layer0_outputs(3207) <= not a;
    layer0_outputs(3208) <= not b;
    layer0_outputs(3209) <= '1';
    layer0_outputs(3210) <= not (a xor b);
    layer0_outputs(3211) <= not a or b;
    layer0_outputs(3212) <= a and b;
    layer0_outputs(3213) <= not (a xor b);
    layer0_outputs(3214) <= not b;
    layer0_outputs(3215) <= '1';
    layer0_outputs(3216) <= a and b;
    layer0_outputs(3217) <= b;
    layer0_outputs(3218) <= a;
    layer0_outputs(3219) <= a;
    layer0_outputs(3220) <= not (a or b);
    layer0_outputs(3221) <= b;
    layer0_outputs(3222) <= a;
    layer0_outputs(3223) <= a xor b;
    layer0_outputs(3224) <= a;
    layer0_outputs(3225) <= a or b;
    layer0_outputs(3226) <= not (a xor b);
    layer0_outputs(3227) <= not b;
    layer0_outputs(3228) <= a and b;
    layer0_outputs(3229) <= not b or a;
    layer0_outputs(3230) <= not (a xor b);
    layer0_outputs(3231) <= a or b;
    layer0_outputs(3232) <= '0';
    layer0_outputs(3233) <= '0';
    layer0_outputs(3234) <= not (a or b);
    layer0_outputs(3235) <= '0';
    layer0_outputs(3236) <= b;
    layer0_outputs(3237) <= not a;
    layer0_outputs(3238) <= not (a xor b);
    layer0_outputs(3239) <= not (a and b);
    layer0_outputs(3240) <= b;
    layer0_outputs(3241) <= not (a or b);
    layer0_outputs(3242) <= b;
    layer0_outputs(3243) <= b and not a;
    layer0_outputs(3244) <= not (a and b);
    layer0_outputs(3245) <= b and not a;
    layer0_outputs(3246) <= not (a and b);
    layer0_outputs(3247) <= b and not a;
    layer0_outputs(3248) <= a;
    layer0_outputs(3249) <= a or b;
    layer0_outputs(3250) <= not b;
    layer0_outputs(3251) <= not (a xor b);
    layer0_outputs(3252) <= not (a or b);
    layer0_outputs(3253) <= b;
    layer0_outputs(3254) <= not a;
    layer0_outputs(3255) <= '1';
    layer0_outputs(3256) <= a xor b;
    layer0_outputs(3257) <= a or b;
    layer0_outputs(3258) <= a xor b;
    layer0_outputs(3259) <= not (a xor b);
    layer0_outputs(3260) <= not b;
    layer0_outputs(3261) <= not b or a;
    layer0_outputs(3262) <= not (a xor b);
    layer0_outputs(3263) <= not a;
    layer0_outputs(3264) <= not a;
    layer0_outputs(3265) <= not (a xor b);
    layer0_outputs(3266) <= a xor b;
    layer0_outputs(3267) <= '0';
    layer0_outputs(3268) <= a xor b;
    layer0_outputs(3269) <= not (a xor b);
    layer0_outputs(3270) <= b and not a;
    layer0_outputs(3271) <= not b or a;
    layer0_outputs(3272) <= not b or a;
    layer0_outputs(3273) <= a and not b;
    layer0_outputs(3274) <= a and not b;
    layer0_outputs(3275) <= b;
    layer0_outputs(3276) <= not a;
    layer0_outputs(3277) <= a or b;
    layer0_outputs(3278) <= a and b;
    layer0_outputs(3279) <= a or b;
    layer0_outputs(3280) <= '1';
    layer0_outputs(3281) <= not (a or b);
    layer0_outputs(3282) <= a xor b;
    layer0_outputs(3283) <= a or b;
    layer0_outputs(3284) <= b and not a;
    layer0_outputs(3285) <= a and b;
    layer0_outputs(3286) <= a or b;
    layer0_outputs(3287) <= a and b;
    layer0_outputs(3288) <= a xor b;
    layer0_outputs(3289) <= not a;
    layer0_outputs(3290) <= not (a or b);
    layer0_outputs(3291) <= b and not a;
    layer0_outputs(3292) <= not (a or b);
    layer0_outputs(3293) <= b;
    layer0_outputs(3294) <= '1';
    layer0_outputs(3295) <= not b;
    layer0_outputs(3296) <= b and not a;
    layer0_outputs(3297) <= a or b;
    layer0_outputs(3298) <= a and not b;
    layer0_outputs(3299) <= a and not b;
    layer0_outputs(3300) <= not b;
    layer0_outputs(3301) <= a or b;
    layer0_outputs(3302) <= a or b;
    layer0_outputs(3303) <= not a;
    layer0_outputs(3304) <= b and not a;
    layer0_outputs(3305) <= '1';
    layer0_outputs(3306) <= not b or a;
    layer0_outputs(3307) <= not (a xor b);
    layer0_outputs(3308) <= a;
    layer0_outputs(3309) <= b;
    layer0_outputs(3310) <= not a;
    layer0_outputs(3311) <= a xor b;
    layer0_outputs(3312) <= a or b;
    layer0_outputs(3313) <= not (a and b);
    layer0_outputs(3314) <= not (a xor b);
    layer0_outputs(3315) <= not b;
    layer0_outputs(3316) <= not a;
    layer0_outputs(3317) <= b;
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= b;
    layer0_outputs(3320) <= b;
    layer0_outputs(3321) <= a xor b;
    layer0_outputs(3322) <= not b or a;
    layer0_outputs(3323) <= a or b;
    layer0_outputs(3324) <= a and not b;
    layer0_outputs(3325) <= a or b;
    layer0_outputs(3326) <= b and not a;
    layer0_outputs(3327) <= not (a or b);
    layer0_outputs(3328) <= not b;
    layer0_outputs(3329) <= b;
    layer0_outputs(3330) <= not a or b;
    layer0_outputs(3331) <= not (a or b);
    layer0_outputs(3332) <= not a or b;
    layer0_outputs(3333) <= a or b;
    layer0_outputs(3334) <= a and not b;
    layer0_outputs(3335) <= '1';
    layer0_outputs(3336) <= not b;
    layer0_outputs(3337) <= b and not a;
    layer0_outputs(3338) <= not b or a;
    layer0_outputs(3339) <= not (a and b);
    layer0_outputs(3340) <= not b or a;
    layer0_outputs(3341) <= a;
    layer0_outputs(3342) <= not a or b;
    layer0_outputs(3343) <= a xor b;
    layer0_outputs(3344) <= not (a or b);
    layer0_outputs(3345) <= a and not b;
    layer0_outputs(3346) <= '1';
    layer0_outputs(3347) <= not b;
    layer0_outputs(3348) <= a or b;
    layer0_outputs(3349) <= a xor b;
    layer0_outputs(3350) <= a and not b;
    layer0_outputs(3351) <= a or b;
    layer0_outputs(3352) <= a;
    layer0_outputs(3353) <= '0';
    layer0_outputs(3354) <= a xor b;
    layer0_outputs(3355) <= a and not b;
    layer0_outputs(3356) <= not a or b;
    layer0_outputs(3357) <= a and not b;
    layer0_outputs(3358) <= a and not b;
    layer0_outputs(3359) <= not (a or b);
    layer0_outputs(3360) <= not (a and b);
    layer0_outputs(3361) <= b and not a;
    layer0_outputs(3362) <= a;
    layer0_outputs(3363) <= not a or b;
    layer0_outputs(3364) <= a;
    layer0_outputs(3365) <= a xor b;
    layer0_outputs(3366) <= not (a and b);
    layer0_outputs(3367) <= b and not a;
    layer0_outputs(3368) <= b;
    layer0_outputs(3369) <= a and not b;
    layer0_outputs(3370) <= not a or b;
    layer0_outputs(3371) <= not b or a;
    layer0_outputs(3372) <= a xor b;
    layer0_outputs(3373) <= a or b;
    layer0_outputs(3374) <= '1';
    layer0_outputs(3375) <= not b or a;
    layer0_outputs(3376) <= not (a or b);
    layer0_outputs(3377) <= not (a or b);
    layer0_outputs(3378) <= a and b;
    layer0_outputs(3379) <= not b;
    layer0_outputs(3380) <= a;
    layer0_outputs(3381) <= a and not b;
    layer0_outputs(3382) <= a or b;
    layer0_outputs(3383) <= not b or a;
    layer0_outputs(3384) <= not a or b;
    layer0_outputs(3385) <= not b or a;
    layer0_outputs(3386) <= a;
    layer0_outputs(3387) <= not (a or b);
    layer0_outputs(3388) <= not (a xor b);
    layer0_outputs(3389) <= a and b;
    layer0_outputs(3390) <= b;
    layer0_outputs(3391) <= a and b;
    layer0_outputs(3392) <= a xor b;
    layer0_outputs(3393) <= not a or b;
    layer0_outputs(3394) <= '0';
    layer0_outputs(3395) <= a xor b;
    layer0_outputs(3396) <= a or b;
    layer0_outputs(3397) <= a or b;
    layer0_outputs(3398) <= a;
    layer0_outputs(3399) <= not (a xor b);
    layer0_outputs(3400) <= not (a or b);
    layer0_outputs(3401) <= not b;
    layer0_outputs(3402) <= a xor b;
    layer0_outputs(3403) <= not a or b;
    layer0_outputs(3404) <= a;
    layer0_outputs(3405) <= not (a or b);
    layer0_outputs(3406) <= b;
    layer0_outputs(3407) <= '1';
    layer0_outputs(3408) <= not a;
    layer0_outputs(3409) <= not (a and b);
    layer0_outputs(3410) <= not (a or b);
    layer0_outputs(3411) <= not (a or b);
    layer0_outputs(3412) <= '0';
    layer0_outputs(3413) <= not (a xor b);
    layer0_outputs(3414) <= not a or b;
    layer0_outputs(3415) <= not (a xor b);
    layer0_outputs(3416) <= not a or b;
    layer0_outputs(3417) <= not (a or b);
    layer0_outputs(3418) <= a or b;
    layer0_outputs(3419) <= a;
    layer0_outputs(3420) <= a and not b;
    layer0_outputs(3421) <= a or b;
    layer0_outputs(3422) <= a xor b;
    layer0_outputs(3423) <= a and not b;
    layer0_outputs(3424) <= '1';
    layer0_outputs(3425) <= not (a and b);
    layer0_outputs(3426) <= not b;
    layer0_outputs(3427) <= not (a and b);
    layer0_outputs(3428) <= '1';
    layer0_outputs(3429) <= '0';
    layer0_outputs(3430) <= a or b;
    layer0_outputs(3431) <= a and b;
    layer0_outputs(3432) <= not a or b;
    layer0_outputs(3433) <= b;
    layer0_outputs(3434) <= '1';
    layer0_outputs(3435) <= not b;
    layer0_outputs(3436) <= not a;
    layer0_outputs(3437) <= not (a and b);
    layer0_outputs(3438) <= a and b;
    layer0_outputs(3439) <= b and not a;
    layer0_outputs(3440) <= not a or b;
    layer0_outputs(3441) <= b;
    layer0_outputs(3442) <= a or b;
    layer0_outputs(3443) <= not a or b;
    layer0_outputs(3444) <= b and not a;
    layer0_outputs(3445) <= not (a xor b);
    layer0_outputs(3446) <= a xor b;
    layer0_outputs(3447) <= not b;
    layer0_outputs(3448) <= not (a xor b);
    layer0_outputs(3449) <= b;
    layer0_outputs(3450) <= a or b;
    layer0_outputs(3451) <= a;
    layer0_outputs(3452) <= b;
    layer0_outputs(3453) <= not (a or b);
    layer0_outputs(3454) <= not (a xor b);
    layer0_outputs(3455) <= '1';
    layer0_outputs(3456) <= a or b;
    layer0_outputs(3457) <= '0';
    layer0_outputs(3458) <= a or b;
    layer0_outputs(3459) <= not a;
    layer0_outputs(3460) <= not b;
    layer0_outputs(3461) <= b;
    layer0_outputs(3462) <= not (a and b);
    layer0_outputs(3463) <= not (a xor b);
    layer0_outputs(3464) <= not a;
    layer0_outputs(3465) <= a;
    layer0_outputs(3466) <= not (a and b);
    layer0_outputs(3467) <= '1';
    layer0_outputs(3468) <= a or b;
    layer0_outputs(3469) <= b;
    layer0_outputs(3470) <= b and not a;
    layer0_outputs(3471) <= not (a and b);
    layer0_outputs(3472) <= a xor b;
    layer0_outputs(3473) <= a or b;
    layer0_outputs(3474) <= b;
    layer0_outputs(3475) <= '0';
    layer0_outputs(3476) <= a and b;
    layer0_outputs(3477) <= a and b;
    layer0_outputs(3478) <= not b;
    layer0_outputs(3479) <= not a or b;
    layer0_outputs(3480) <= not b or a;
    layer0_outputs(3481) <= a xor b;
    layer0_outputs(3482) <= not a;
    layer0_outputs(3483) <= a or b;
    layer0_outputs(3484) <= a or b;
    layer0_outputs(3485) <= not a;
    layer0_outputs(3486) <= a and b;
    layer0_outputs(3487) <= '1';
    layer0_outputs(3488) <= not (a or b);
    layer0_outputs(3489) <= not b;
    layer0_outputs(3490) <= '1';
    layer0_outputs(3491) <= a or b;
    layer0_outputs(3492) <= a xor b;
    layer0_outputs(3493) <= b;
    layer0_outputs(3494) <= a and b;
    layer0_outputs(3495) <= a and b;
    layer0_outputs(3496) <= a and b;
    layer0_outputs(3497) <= not a;
    layer0_outputs(3498) <= b and not a;
    layer0_outputs(3499) <= b;
    layer0_outputs(3500) <= not b;
    layer0_outputs(3501) <= b;
    layer0_outputs(3502) <= not (a or b);
    layer0_outputs(3503) <= not a;
    layer0_outputs(3504) <= not b;
    layer0_outputs(3505) <= not (a or b);
    layer0_outputs(3506) <= a;
    layer0_outputs(3507) <= a and not b;
    layer0_outputs(3508) <= not b;
    layer0_outputs(3509) <= a and not b;
    layer0_outputs(3510) <= not (a xor b);
    layer0_outputs(3511) <= not (a and b);
    layer0_outputs(3512) <= a and b;
    layer0_outputs(3513) <= a or b;
    layer0_outputs(3514) <= not (a or b);
    layer0_outputs(3515) <= a or b;
    layer0_outputs(3516) <= b and not a;
    layer0_outputs(3517) <= not (a or b);
    layer0_outputs(3518) <= not b or a;
    layer0_outputs(3519) <= not (a and b);
    layer0_outputs(3520) <= not a or b;
    layer0_outputs(3521) <= not a or b;
    layer0_outputs(3522) <= not a or b;
    layer0_outputs(3523) <= not a or b;
    layer0_outputs(3524) <= not b;
    layer0_outputs(3525) <= '0';
    layer0_outputs(3526) <= a and b;
    layer0_outputs(3527) <= '1';
    layer0_outputs(3528) <= not (a or b);
    layer0_outputs(3529) <= '0';
    layer0_outputs(3530) <= a or b;
    layer0_outputs(3531) <= a and not b;
    layer0_outputs(3532) <= a or b;
    layer0_outputs(3533) <= b;
    layer0_outputs(3534) <= '1';
    layer0_outputs(3535) <= '1';
    layer0_outputs(3536) <= not a;
    layer0_outputs(3537) <= not a;
    layer0_outputs(3538) <= a and b;
    layer0_outputs(3539) <= not (a and b);
    layer0_outputs(3540) <= not (a and b);
    layer0_outputs(3541) <= not (a or b);
    layer0_outputs(3542) <= a;
    layer0_outputs(3543) <= not (a or b);
    layer0_outputs(3544) <= not a;
    layer0_outputs(3545) <= not b;
    layer0_outputs(3546) <= not b;
    layer0_outputs(3547) <= not (a xor b);
    layer0_outputs(3548) <= not b or a;
    layer0_outputs(3549) <= not (a xor b);
    layer0_outputs(3550) <= a and b;
    layer0_outputs(3551) <= not (a or b);
    layer0_outputs(3552) <= not b;
    layer0_outputs(3553) <= not a or b;
    layer0_outputs(3554) <= not a;
    layer0_outputs(3555) <= not a;
    layer0_outputs(3556) <= a xor b;
    layer0_outputs(3557) <= '1';
    layer0_outputs(3558) <= not (a and b);
    layer0_outputs(3559) <= not (a or b);
    layer0_outputs(3560) <= a;
    layer0_outputs(3561) <= not a or b;
    layer0_outputs(3562) <= not (a or b);
    layer0_outputs(3563) <= a;
    layer0_outputs(3564) <= not (a xor b);
    layer0_outputs(3565) <= a or b;
    layer0_outputs(3566) <= a or b;
    layer0_outputs(3567) <= a;
    layer0_outputs(3568) <= a;
    layer0_outputs(3569) <= a xor b;
    layer0_outputs(3570) <= not a;
    layer0_outputs(3571) <= a or b;
    layer0_outputs(3572) <= a or b;
    layer0_outputs(3573) <= not a;
    layer0_outputs(3574) <= a and not b;
    layer0_outputs(3575) <= a and b;
    layer0_outputs(3576) <= a xor b;
    layer0_outputs(3577) <= '0';
    layer0_outputs(3578) <= not b or a;
    layer0_outputs(3579) <= a and b;
    layer0_outputs(3580) <= '0';
    layer0_outputs(3581) <= a and not b;
    layer0_outputs(3582) <= b and not a;
    layer0_outputs(3583) <= not a or b;
    layer0_outputs(3584) <= b;
    layer0_outputs(3585) <= a and not b;
    layer0_outputs(3586) <= '1';
    layer0_outputs(3587) <= a;
    layer0_outputs(3588) <= not (a xor b);
    layer0_outputs(3589) <= b and not a;
    layer0_outputs(3590) <= not (a or b);
    layer0_outputs(3591) <= a xor b;
    layer0_outputs(3592) <= '0';
    layer0_outputs(3593) <= b;
    layer0_outputs(3594) <= not a or b;
    layer0_outputs(3595) <= '0';
    layer0_outputs(3596) <= not (a or b);
    layer0_outputs(3597) <= not a;
    layer0_outputs(3598) <= not b;
    layer0_outputs(3599) <= not b or a;
    layer0_outputs(3600) <= not (a or b);
    layer0_outputs(3601) <= not (a or b);
    layer0_outputs(3602) <= a xor b;
    layer0_outputs(3603) <= '1';
    layer0_outputs(3604) <= a;
    layer0_outputs(3605) <= not b or a;
    layer0_outputs(3606) <= a or b;
    layer0_outputs(3607) <= b;
    layer0_outputs(3608) <= not (a or b);
    layer0_outputs(3609) <= not (a or b);
    layer0_outputs(3610) <= a or b;
    layer0_outputs(3611) <= not b;
    layer0_outputs(3612) <= not a;
    layer0_outputs(3613) <= not (a xor b);
    layer0_outputs(3614) <= b;
    layer0_outputs(3615) <= not (a and b);
    layer0_outputs(3616) <= '1';
    layer0_outputs(3617) <= not b;
    layer0_outputs(3618) <= not b;
    layer0_outputs(3619) <= b and not a;
    layer0_outputs(3620) <= not a;
    layer0_outputs(3621) <= a;
    layer0_outputs(3622) <= a xor b;
    layer0_outputs(3623) <= '1';
    layer0_outputs(3624) <= b;
    layer0_outputs(3625) <= not a or b;
    layer0_outputs(3626) <= not a;
    layer0_outputs(3627) <= b and not a;
    layer0_outputs(3628) <= not (a or b);
    layer0_outputs(3629) <= '1';
    layer0_outputs(3630) <= a xor b;
    layer0_outputs(3631) <= not a;
    layer0_outputs(3632) <= a;
    layer0_outputs(3633) <= b;
    layer0_outputs(3634) <= a and not b;
    layer0_outputs(3635) <= a or b;
    layer0_outputs(3636) <= a;
    layer0_outputs(3637) <= not a or b;
    layer0_outputs(3638) <= not b;
    layer0_outputs(3639) <= not a or b;
    layer0_outputs(3640) <= not (a and b);
    layer0_outputs(3641) <= a;
    layer0_outputs(3642) <= not a;
    layer0_outputs(3643) <= '0';
    layer0_outputs(3644) <= not (a xor b);
    layer0_outputs(3645) <= not b;
    layer0_outputs(3646) <= not a;
    layer0_outputs(3647) <= b and not a;
    layer0_outputs(3648) <= a;
    layer0_outputs(3649) <= b and not a;
    layer0_outputs(3650) <= a or b;
    layer0_outputs(3651) <= a and not b;
    layer0_outputs(3652) <= not b or a;
    layer0_outputs(3653) <= b and not a;
    layer0_outputs(3654) <= not a;
    layer0_outputs(3655) <= a or b;
    layer0_outputs(3656) <= not a or b;
    layer0_outputs(3657) <= not b;
    layer0_outputs(3658) <= not (a or b);
    layer0_outputs(3659) <= a and b;
    layer0_outputs(3660) <= b;
    layer0_outputs(3661) <= not (a xor b);
    layer0_outputs(3662) <= not (a or b);
    layer0_outputs(3663) <= a xor b;
    layer0_outputs(3664) <= not (a and b);
    layer0_outputs(3665) <= not a;
    layer0_outputs(3666) <= not a or b;
    layer0_outputs(3667) <= not (a or b);
    layer0_outputs(3668) <= a or b;
    layer0_outputs(3669) <= not a;
    layer0_outputs(3670) <= a and not b;
    layer0_outputs(3671) <= not a or b;
    layer0_outputs(3672) <= b;
    layer0_outputs(3673) <= not a or b;
    layer0_outputs(3674) <= a and b;
    layer0_outputs(3675) <= not (a or b);
    layer0_outputs(3676) <= a;
    layer0_outputs(3677) <= not (a or b);
    layer0_outputs(3678) <= b and not a;
    layer0_outputs(3679) <= b and not a;
    layer0_outputs(3680) <= b and not a;
    layer0_outputs(3681) <= not (a or b);
    layer0_outputs(3682) <= not b or a;
    layer0_outputs(3683) <= a xor b;
    layer0_outputs(3684) <= a and b;
    layer0_outputs(3685) <= a;
    layer0_outputs(3686) <= a;
    layer0_outputs(3687) <= '0';
    layer0_outputs(3688) <= b;
    layer0_outputs(3689) <= not a;
    layer0_outputs(3690) <= not b or a;
    layer0_outputs(3691) <= '0';
    layer0_outputs(3692) <= not b;
    layer0_outputs(3693) <= not (a or b);
    layer0_outputs(3694) <= not (a xor b);
    layer0_outputs(3695) <= not a or b;
    layer0_outputs(3696) <= not a;
    layer0_outputs(3697) <= not (a and b);
    layer0_outputs(3698) <= not a or b;
    layer0_outputs(3699) <= not a;
    layer0_outputs(3700) <= a;
    layer0_outputs(3701) <= a and b;
    layer0_outputs(3702) <= a;
    layer0_outputs(3703) <= a and not b;
    layer0_outputs(3704) <= a or b;
    layer0_outputs(3705) <= not b;
    layer0_outputs(3706) <= b;
    layer0_outputs(3707) <= a;
    layer0_outputs(3708) <= not (a or b);
    layer0_outputs(3709) <= not a or b;
    layer0_outputs(3710) <= b and not a;
    layer0_outputs(3711) <= not (a or b);
    layer0_outputs(3712) <= a or b;
    layer0_outputs(3713) <= '0';
    layer0_outputs(3714) <= a or b;
    layer0_outputs(3715) <= not (a and b);
    layer0_outputs(3716) <= not (a and b);
    layer0_outputs(3717) <= b;
    layer0_outputs(3718) <= b;
    layer0_outputs(3719) <= not (a xor b);
    layer0_outputs(3720) <= not (a xor b);
    layer0_outputs(3721) <= not b;
    layer0_outputs(3722) <= '0';
    layer0_outputs(3723) <= not a or b;
    layer0_outputs(3724) <= a or b;
    layer0_outputs(3725) <= not (a or b);
    layer0_outputs(3726) <= not b;
    layer0_outputs(3727) <= a;
    layer0_outputs(3728) <= a;
    layer0_outputs(3729) <= a or b;
    layer0_outputs(3730) <= b;
    layer0_outputs(3731) <= b and not a;
    layer0_outputs(3732) <= not a;
    layer0_outputs(3733) <= not b or a;
    layer0_outputs(3734) <= not (a xor b);
    layer0_outputs(3735) <= a or b;
    layer0_outputs(3736) <= not a or b;
    layer0_outputs(3737) <= a or b;
    layer0_outputs(3738) <= not b;
    layer0_outputs(3739) <= a;
    layer0_outputs(3740) <= '1';
    layer0_outputs(3741) <= not (a or b);
    layer0_outputs(3742) <= '0';
    layer0_outputs(3743) <= a or b;
    layer0_outputs(3744) <= a or b;
    layer0_outputs(3745) <= a or b;
    layer0_outputs(3746) <= a;
    layer0_outputs(3747) <= not b or a;
    layer0_outputs(3748) <= b and not a;
    layer0_outputs(3749) <= a;
    layer0_outputs(3750) <= not (a and b);
    layer0_outputs(3751) <= not (a or b);
    layer0_outputs(3752) <= a and b;
    layer0_outputs(3753) <= b and not a;
    layer0_outputs(3754) <= b;
    layer0_outputs(3755) <= not b;
    layer0_outputs(3756) <= not b;
    layer0_outputs(3757) <= not (a xor b);
    layer0_outputs(3758) <= a or b;
    layer0_outputs(3759) <= not (a or b);
    layer0_outputs(3760) <= '0';
    layer0_outputs(3761) <= '1';
    layer0_outputs(3762) <= a or b;
    layer0_outputs(3763) <= not a;
    layer0_outputs(3764) <= a;
    layer0_outputs(3765) <= not (a or b);
    layer0_outputs(3766) <= a or b;
    layer0_outputs(3767) <= not (a or b);
    layer0_outputs(3768) <= not (a and b);
    layer0_outputs(3769) <= a xor b;
    layer0_outputs(3770) <= not a or b;
    layer0_outputs(3771) <= not b or a;
    layer0_outputs(3772) <= a and b;
    layer0_outputs(3773) <= not (a and b);
    layer0_outputs(3774) <= not (a or b);
    layer0_outputs(3775) <= not (a or b);
    layer0_outputs(3776) <= not b or a;
    layer0_outputs(3777) <= '0';
    layer0_outputs(3778) <= b;
    layer0_outputs(3779) <= b and not a;
    layer0_outputs(3780) <= '0';
    layer0_outputs(3781) <= b;
    layer0_outputs(3782) <= not b or a;
    layer0_outputs(3783) <= a or b;
    layer0_outputs(3784) <= a xor b;
    layer0_outputs(3785) <= not b;
    layer0_outputs(3786) <= b;
    layer0_outputs(3787) <= not b;
    layer0_outputs(3788) <= a xor b;
    layer0_outputs(3789) <= a or b;
    layer0_outputs(3790) <= a;
    layer0_outputs(3791) <= not (a or b);
    layer0_outputs(3792) <= a or b;
    layer0_outputs(3793) <= not (a or b);
    layer0_outputs(3794) <= not (a and b);
    layer0_outputs(3795) <= a xor b;
    layer0_outputs(3796) <= not a;
    layer0_outputs(3797) <= not b;
    layer0_outputs(3798) <= b and not a;
    layer0_outputs(3799) <= not (a or b);
    layer0_outputs(3800) <= not b or a;
    layer0_outputs(3801) <= '0';
    layer0_outputs(3802) <= not (a or b);
    layer0_outputs(3803) <= a and not b;
    layer0_outputs(3804) <= not b;
    layer0_outputs(3805) <= not b or a;
    layer0_outputs(3806) <= a and not b;
    layer0_outputs(3807) <= a and not b;
    layer0_outputs(3808) <= a and not b;
    layer0_outputs(3809) <= not (a or b);
    layer0_outputs(3810) <= not (a xor b);
    layer0_outputs(3811) <= not b;
    layer0_outputs(3812) <= a or b;
    layer0_outputs(3813) <= a;
    layer0_outputs(3814) <= '0';
    layer0_outputs(3815) <= a;
    layer0_outputs(3816) <= b;
    layer0_outputs(3817) <= not a;
    layer0_outputs(3818) <= b;
    layer0_outputs(3819) <= not b or a;
    layer0_outputs(3820) <= not a or b;
    layer0_outputs(3821) <= not b or a;
    layer0_outputs(3822) <= a xor b;
    layer0_outputs(3823) <= b and not a;
    layer0_outputs(3824) <= a and b;
    layer0_outputs(3825) <= b and not a;
    layer0_outputs(3826) <= not (a xor b);
    layer0_outputs(3827) <= b and not a;
    layer0_outputs(3828) <= not a;
    layer0_outputs(3829) <= not a or b;
    layer0_outputs(3830) <= b;
    layer0_outputs(3831) <= not (a or b);
    layer0_outputs(3832) <= b and not a;
    layer0_outputs(3833) <= not b;
    layer0_outputs(3834) <= not b or a;
    layer0_outputs(3835) <= a or b;
    layer0_outputs(3836) <= '1';
    layer0_outputs(3837) <= not (a or b);
    layer0_outputs(3838) <= not (a or b);
    layer0_outputs(3839) <= not b or a;
    layer0_outputs(3840) <= b;
    layer0_outputs(3841) <= a;
    layer0_outputs(3842) <= '0';
    layer0_outputs(3843) <= not a or b;
    layer0_outputs(3844) <= not (a and b);
    layer0_outputs(3845) <= not (a xor b);
    layer0_outputs(3846) <= not b or a;
    layer0_outputs(3847) <= a or b;
    layer0_outputs(3848) <= not b;
    layer0_outputs(3849) <= '1';
    layer0_outputs(3850) <= not b or a;
    layer0_outputs(3851) <= '0';
    layer0_outputs(3852) <= not a;
    layer0_outputs(3853) <= not b or a;
    layer0_outputs(3854) <= not (a xor b);
    layer0_outputs(3855) <= not (a xor b);
    layer0_outputs(3856) <= '1';
    layer0_outputs(3857) <= a;
    layer0_outputs(3858) <= a;
    layer0_outputs(3859) <= not b;
    layer0_outputs(3860) <= b;
    layer0_outputs(3861) <= not (a or b);
    layer0_outputs(3862) <= not (a or b);
    layer0_outputs(3863) <= not a or b;
    layer0_outputs(3864) <= not b;
    layer0_outputs(3865) <= a xor b;
    layer0_outputs(3866) <= a xor b;
    layer0_outputs(3867) <= not a;
    layer0_outputs(3868) <= b and not a;
    layer0_outputs(3869) <= a or b;
    layer0_outputs(3870) <= not b;
    layer0_outputs(3871) <= not (a and b);
    layer0_outputs(3872) <= not a or b;
    layer0_outputs(3873) <= '0';
    layer0_outputs(3874) <= not a;
    layer0_outputs(3875) <= not b or a;
    layer0_outputs(3876) <= not b;
    layer0_outputs(3877) <= b and not a;
    layer0_outputs(3878) <= not b or a;
    layer0_outputs(3879) <= b;
    layer0_outputs(3880) <= not a or b;
    layer0_outputs(3881) <= not a or b;
    layer0_outputs(3882) <= not (a or b);
    layer0_outputs(3883) <= not b;
    layer0_outputs(3884) <= not a;
    layer0_outputs(3885) <= not (a xor b);
    layer0_outputs(3886) <= not (a and b);
    layer0_outputs(3887) <= not b or a;
    layer0_outputs(3888) <= not (a and b);
    layer0_outputs(3889) <= b and not a;
    layer0_outputs(3890) <= not a;
    layer0_outputs(3891) <= not b;
    layer0_outputs(3892) <= a and not b;
    layer0_outputs(3893) <= a or b;
    layer0_outputs(3894) <= b;
    layer0_outputs(3895) <= not b;
    layer0_outputs(3896) <= a and not b;
    layer0_outputs(3897) <= not (a xor b);
    layer0_outputs(3898) <= '1';
    layer0_outputs(3899) <= not (a or b);
    layer0_outputs(3900) <= a or b;
    layer0_outputs(3901) <= a and b;
    layer0_outputs(3902) <= not (a xor b);
    layer0_outputs(3903) <= not a;
    layer0_outputs(3904) <= not (a xor b);
    layer0_outputs(3905) <= a and b;
    layer0_outputs(3906) <= not a;
    layer0_outputs(3907) <= not a or b;
    layer0_outputs(3908) <= not (a xor b);
    layer0_outputs(3909) <= '0';
    layer0_outputs(3910) <= not (a xor b);
    layer0_outputs(3911) <= a xor b;
    layer0_outputs(3912) <= a and b;
    layer0_outputs(3913) <= not (a or b);
    layer0_outputs(3914) <= not (a or b);
    layer0_outputs(3915) <= a and not b;
    layer0_outputs(3916) <= a or b;
    layer0_outputs(3917) <= not a;
    layer0_outputs(3918) <= not (a or b);
    layer0_outputs(3919) <= not a or b;
    layer0_outputs(3920) <= not (a or b);
    layer0_outputs(3921) <= b;
    layer0_outputs(3922) <= not b;
    layer0_outputs(3923) <= not a;
    layer0_outputs(3924) <= a or b;
    layer0_outputs(3925) <= not b;
    layer0_outputs(3926) <= a and b;
    layer0_outputs(3927) <= not (a or b);
    layer0_outputs(3928) <= a or b;
    layer0_outputs(3929) <= not (a xor b);
    layer0_outputs(3930) <= b;
    layer0_outputs(3931) <= not b or a;
    layer0_outputs(3932) <= a and not b;
    layer0_outputs(3933) <= a;
    layer0_outputs(3934) <= not (a xor b);
    layer0_outputs(3935) <= '1';
    layer0_outputs(3936) <= a;
    layer0_outputs(3937) <= '0';
    layer0_outputs(3938) <= not (a xor b);
    layer0_outputs(3939) <= not b or a;
    layer0_outputs(3940) <= not a;
    layer0_outputs(3941) <= not (a xor b);
    layer0_outputs(3942) <= not b;
    layer0_outputs(3943) <= '0';
    layer0_outputs(3944) <= not a;
    layer0_outputs(3945) <= b;
    layer0_outputs(3946) <= '1';
    layer0_outputs(3947) <= '1';
    layer0_outputs(3948) <= not b;
    layer0_outputs(3949) <= b and not a;
    layer0_outputs(3950) <= a;
    layer0_outputs(3951) <= not (a xor b);
    layer0_outputs(3952) <= '0';
    layer0_outputs(3953) <= b;
    layer0_outputs(3954) <= a;
    layer0_outputs(3955) <= not (a and b);
    layer0_outputs(3956) <= b;
    layer0_outputs(3957) <= a and b;
    layer0_outputs(3958) <= a and not b;
    layer0_outputs(3959) <= not a or b;
    layer0_outputs(3960) <= not a;
    layer0_outputs(3961) <= not b;
    layer0_outputs(3962) <= '1';
    layer0_outputs(3963) <= a xor b;
    layer0_outputs(3964) <= not a;
    layer0_outputs(3965) <= '0';
    layer0_outputs(3966) <= not (a or b);
    layer0_outputs(3967) <= not a;
    layer0_outputs(3968) <= not (a xor b);
    layer0_outputs(3969) <= '1';
    layer0_outputs(3970) <= b and not a;
    layer0_outputs(3971) <= a or b;
    layer0_outputs(3972) <= not b;
    layer0_outputs(3973) <= not (a or b);
    layer0_outputs(3974) <= '1';
    layer0_outputs(3975) <= '0';
    layer0_outputs(3976) <= a and b;
    layer0_outputs(3977) <= b and not a;
    layer0_outputs(3978) <= a or b;
    layer0_outputs(3979) <= a or b;
    layer0_outputs(3980) <= not a or b;
    layer0_outputs(3981) <= not b;
    layer0_outputs(3982) <= not a or b;
    layer0_outputs(3983) <= not a;
    layer0_outputs(3984) <= not (a xor b);
    layer0_outputs(3985) <= a or b;
    layer0_outputs(3986) <= b and not a;
    layer0_outputs(3987) <= '1';
    layer0_outputs(3988) <= not b;
    layer0_outputs(3989) <= a xor b;
    layer0_outputs(3990) <= a;
    layer0_outputs(3991) <= not a or b;
    layer0_outputs(3992) <= b and not a;
    layer0_outputs(3993) <= a xor b;
    layer0_outputs(3994) <= a;
    layer0_outputs(3995) <= b;
    layer0_outputs(3996) <= a and not b;
    layer0_outputs(3997) <= a xor b;
    layer0_outputs(3998) <= not b;
    layer0_outputs(3999) <= a and not b;
    layer0_outputs(4000) <= '1';
    layer0_outputs(4001) <= a and b;
    layer0_outputs(4002) <= not a or b;
    layer0_outputs(4003) <= b and not a;
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= not (a xor b);
    layer0_outputs(4006) <= not a;
    layer0_outputs(4007) <= a or b;
    layer0_outputs(4008) <= not b;
    layer0_outputs(4009) <= not (a or b);
    layer0_outputs(4010) <= not (a and b);
    layer0_outputs(4011) <= a and not b;
    layer0_outputs(4012) <= not a or b;
    layer0_outputs(4013) <= '1';
    layer0_outputs(4014) <= not (a or b);
    layer0_outputs(4015) <= not (a or b);
    layer0_outputs(4016) <= not a;
    layer0_outputs(4017) <= not b;
    layer0_outputs(4018) <= '0';
    layer0_outputs(4019) <= b and not a;
    layer0_outputs(4020) <= a and b;
    layer0_outputs(4021) <= a;
    layer0_outputs(4022) <= b and not a;
    layer0_outputs(4023) <= '1';
    layer0_outputs(4024) <= b and not a;
    layer0_outputs(4025) <= not a or b;
    layer0_outputs(4026) <= not b or a;
    layer0_outputs(4027) <= not b or a;
    layer0_outputs(4028) <= a;
    layer0_outputs(4029) <= not b;
    layer0_outputs(4030) <= b and not a;
    layer0_outputs(4031) <= not (a or b);
    layer0_outputs(4032) <= not a or b;
    layer0_outputs(4033) <= a or b;
    layer0_outputs(4034) <= not b or a;
    layer0_outputs(4035) <= a and b;
    layer0_outputs(4036) <= not b;
    layer0_outputs(4037) <= b and not a;
    layer0_outputs(4038) <= not a or b;
    layer0_outputs(4039) <= not b or a;
    layer0_outputs(4040) <= not (a xor b);
    layer0_outputs(4041) <= not (a xor b);
    layer0_outputs(4042) <= a and not b;
    layer0_outputs(4043) <= b and not a;
    layer0_outputs(4044) <= a;
    layer0_outputs(4045) <= b;
    layer0_outputs(4046) <= a xor b;
    layer0_outputs(4047) <= not (a xor b);
    layer0_outputs(4048) <= not b;
    layer0_outputs(4049) <= a and not b;
    layer0_outputs(4050) <= not b;
    layer0_outputs(4051) <= not a;
    layer0_outputs(4052) <= b and not a;
    layer0_outputs(4053) <= not (a xor b);
    layer0_outputs(4054) <= not b;
    layer0_outputs(4055) <= b and not a;
    layer0_outputs(4056) <= a or b;
    layer0_outputs(4057) <= a;
    layer0_outputs(4058) <= b;
    layer0_outputs(4059) <= not b;
    layer0_outputs(4060) <= b;
    layer0_outputs(4061) <= not b or a;
    layer0_outputs(4062) <= b;
    layer0_outputs(4063) <= not (a and b);
    layer0_outputs(4064) <= not (a or b);
    layer0_outputs(4065) <= b and not a;
    layer0_outputs(4066) <= '0';
    layer0_outputs(4067) <= not (a or b);
    layer0_outputs(4068) <= not a;
    layer0_outputs(4069) <= b and not a;
    layer0_outputs(4070) <= a or b;
    layer0_outputs(4071) <= a and not b;
    layer0_outputs(4072) <= '1';
    layer0_outputs(4073) <= b;
    layer0_outputs(4074) <= not a or b;
    layer0_outputs(4075) <= not a;
    layer0_outputs(4076) <= not b or a;
    layer0_outputs(4077) <= not a;
    layer0_outputs(4078) <= not b;
    layer0_outputs(4079) <= a and not b;
    layer0_outputs(4080) <= a xor b;
    layer0_outputs(4081) <= '1';
    layer0_outputs(4082) <= a or b;
    layer0_outputs(4083) <= a xor b;
    layer0_outputs(4084) <= not a or b;
    layer0_outputs(4085) <= not (a or b);
    layer0_outputs(4086) <= a or b;
    layer0_outputs(4087) <= not b;
    layer0_outputs(4088) <= not b;
    layer0_outputs(4089) <= not (a and b);
    layer0_outputs(4090) <= '0';
    layer0_outputs(4091) <= not (a xor b);
    layer0_outputs(4092) <= a;
    layer0_outputs(4093) <= '1';
    layer0_outputs(4094) <= a or b;
    layer0_outputs(4095) <= a and not b;
    layer0_outputs(4096) <= b;
    layer0_outputs(4097) <= not (a or b);
    layer0_outputs(4098) <= not b;
    layer0_outputs(4099) <= '0';
    layer0_outputs(4100) <= not b;
    layer0_outputs(4101) <= not b;
    layer0_outputs(4102) <= a xor b;
    layer0_outputs(4103) <= not b or a;
    layer0_outputs(4104) <= a and not b;
    layer0_outputs(4105) <= not b or a;
    layer0_outputs(4106) <= a and not b;
    layer0_outputs(4107) <= a;
    layer0_outputs(4108) <= a xor b;
    layer0_outputs(4109) <= not b;
    layer0_outputs(4110) <= not (a xor b);
    layer0_outputs(4111) <= not (a or b);
    layer0_outputs(4112) <= a xor b;
    layer0_outputs(4113) <= not b;
    layer0_outputs(4114) <= a and not b;
    layer0_outputs(4115) <= a or b;
    layer0_outputs(4116) <= a or b;
    layer0_outputs(4117) <= a and b;
    layer0_outputs(4118) <= a or b;
    layer0_outputs(4119) <= a xor b;
    layer0_outputs(4120) <= b;
    layer0_outputs(4121) <= not a or b;
    layer0_outputs(4122) <= a and b;
    layer0_outputs(4123) <= a and b;
    layer0_outputs(4124) <= not a or b;
    layer0_outputs(4125) <= a or b;
    layer0_outputs(4126) <= not (a or b);
    layer0_outputs(4127) <= a;
    layer0_outputs(4128) <= not a;
    layer0_outputs(4129) <= not a or b;
    layer0_outputs(4130) <= a or b;
    layer0_outputs(4131) <= not (a xor b);
    layer0_outputs(4132) <= not (a xor b);
    layer0_outputs(4133) <= b;
    layer0_outputs(4134) <= not b or a;
    layer0_outputs(4135) <= not b;
    layer0_outputs(4136) <= b and not a;
    layer0_outputs(4137) <= not (a or b);
    layer0_outputs(4138) <= a;
    layer0_outputs(4139) <= a or b;
    layer0_outputs(4140) <= not b;
    layer0_outputs(4141) <= a and b;
    layer0_outputs(4142) <= a xor b;
    layer0_outputs(4143) <= not (a xor b);
    layer0_outputs(4144) <= a and b;
    layer0_outputs(4145) <= not (a xor b);
    layer0_outputs(4146) <= not a;
    layer0_outputs(4147) <= not (a xor b);
    layer0_outputs(4148) <= not b or a;
    layer0_outputs(4149) <= b;
    layer0_outputs(4150) <= not (a xor b);
    layer0_outputs(4151) <= not (a xor b);
    layer0_outputs(4152) <= b;
    layer0_outputs(4153) <= a;
    layer0_outputs(4154) <= a;
    layer0_outputs(4155) <= not a or b;
    layer0_outputs(4156) <= not a;
    layer0_outputs(4157) <= not a or b;
    layer0_outputs(4158) <= a;
    layer0_outputs(4159) <= b;
    layer0_outputs(4160) <= a or b;
    layer0_outputs(4161) <= not b or a;
    layer0_outputs(4162) <= a or b;
    layer0_outputs(4163) <= not (a xor b);
    layer0_outputs(4164) <= not a or b;
    layer0_outputs(4165) <= '1';
    layer0_outputs(4166) <= not (a or b);
    layer0_outputs(4167) <= not (a or b);
    layer0_outputs(4168) <= not b;
    layer0_outputs(4169) <= '1';
    layer0_outputs(4170) <= not (a or b);
    layer0_outputs(4171) <= not a;
    layer0_outputs(4172) <= a or b;
    layer0_outputs(4173) <= a xor b;
    layer0_outputs(4174) <= '0';
    layer0_outputs(4175) <= not a or b;
    layer0_outputs(4176) <= not (a or b);
    layer0_outputs(4177) <= not b;
    layer0_outputs(4178) <= '1';
    layer0_outputs(4179) <= a;
    layer0_outputs(4180) <= not a;
    layer0_outputs(4181) <= a and not b;
    layer0_outputs(4182) <= a or b;
    layer0_outputs(4183) <= a and b;
    layer0_outputs(4184) <= a and not b;
    layer0_outputs(4185) <= b and not a;
    layer0_outputs(4186) <= a xor b;
    layer0_outputs(4187) <= not (a and b);
    layer0_outputs(4188) <= not b or a;
    layer0_outputs(4189) <= not (a or b);
    layer0_outputs(4190) <= '0';
    layer0_outputs(4191) <= not b or a;
    layer0_outputs(4192) <= not a or b;
    layer0_outputs(4193) <= a and not b;
    layer0_outputs(4194) <= '1';
    layer0_outputs(4195) <= not a;
    layer0_outputs(4196) <= not a;
    layer0_outputs(4197) <= '1';
    layer0_outputs(4198) <= b;
    layer0_outputs(4199) <= a and b;
    layer0_outputs(4200) <= a or b;
    layer0_outputs(4201) <= a;
    layer0_outputs(4202) <= '0';
    layer0_outputs(4203) <= not (a xor b);
    layer0_outputs(4204) <= a;
    layer0_outputs(4205) <= not (a or b);
    layer0_outputs(4206) <= not a;
    layer0_outputs(4207) <= a or b;
    layer0_outputs(4208) <= not (a or b);
    layer0_outputs(4209) <= a and not b;
    layer0_outputs(4210) <= '1';
    layer0_outputs(4211) <= a xor b;
    layer0_outputs(4212) <= a or b;
    layer0_outputs(4213) <= a or b;
    layer0_outputs(4214) <= a xor b;
    layer0_outputs(4215) <= not (a xor b);
    layer0_outputs(4216) <= not (a or b);
    layer0_outputs(4217) <= a or b;
    layer0_outputs(4218) <= a;
    layer0_outputs(4219) <= '0';
    layer0_outputs(4220) <= a and not b;
    layer0_outputs(4221) <= a and b;
    layer0_outputs(4222) <= not (a or b);
    layer0_outputs(4223) <= '0';
    layer0_outputs(4224) <= not (a xor b);
    layer0_outputs(4225) <= b and not a;
    layer0_outputs(4226) <= not b;
    layer0_outputs(4227) <= not b;
    layer0_outputs(4228) <= '0';
    layer0_outputs(4229) <= not a;
    layer0_outputs(4230) <= a;
    layer0_outputs(4231) <= a or b;
    layer0_outputs(4232) <= b;
    layer0_outputs(4233) <= not a;
    layer0_outputs(4234) <= '0';
    layer0_outputs(4235) <= a or b;
    layer0_outputs(4236) <= not a or b;
    layer0_outputs(4237) <= not b;
    layer0_outputs(4238) <= not (a xor b);
    layer0_outputs(4239) <= not a;
    layer0_outputs(4240) <= b and not a;
    layer0_outputs(4241) <= not b or a;
    layer0_outputs(4242) <= not b or a;
    layer0_outputs(4243) <= not b;
    layer0_outputs(4244) <= '1';
    layer0_outputs(4245) <= not a;
    layer0_outputs(4246) <= a and not b;
    layer0_outputs(4247) <= not b or a;
    layer0_outputs(4248) <= not a;
    layer0_outputs(4249) <= not (a or b);
    layer0_outputs(4250) <= '1';
    layer0_outputs(4251) <= not a or b;
    layer0_outputs(4252) <= a or b;
    layer0_outputs(4253) <= a;
    layer0_outputs(4254) <= a;
    layer0_outputs(4255) <= '0';
    layer0_outputs(4256) <= not (a and b);
    layer0_outputs(4257) <= a and not b;
    layer0_outputs(4258) <= not a or b;
    layer0_outputs(4259) <= not a or b;
    layer0_outputs(4260) <= not (a and b);
    layer0_outputs(4261) <= a;
    layer0_outputs(4262) <= not (a xor b);
    layer0_outputs(4263) <= '1';
    layer0_outputs(4264) <= not (a or b);
    layer0_outputs(4265) <= '0';
    layer0_outputs(4266) <= not (a or b);
    layer0_outputs(4267) <= not b;
    layer0_outputs(4268) <= not b or a;
    layer0_outputs(4269) <= a;
    layer0_outputs(4270) <= not (a xor b);
    layer0_outputs(4271) <= '0';
    layer0_outputs(4272) <= b;
    layer0_outputs(4273) <= a xor b;
    layer0_outputs(4274) <= '0';
    layer0_outputs(4275) <= b and not a;
    layer0_outputs(4276) <= a and b;
    layer0_outputs(4277) <= '0';
    layer0_outputs(4278) <= '0';
    layer0_outputs(4279) <= b and not a;
    layer0_outputs(4280) <= a or b;
    layer0_outputs(4281) <= not (a and b);
    layer0_outputs(4282) <= not b or a;
    layer0_outputs(4283) <= a xor b;
    layer0_outputs(4284) <= not a;
    layer0_outputs(4285) <= not a;
    layer0_outputs(4286) <= '1';
    layer0_outputs(4287) <= a xor b;
    layer0_outputs(4288) <= b and not a;
    layer0_outputs(4289) <= '1';
    layer0_outputs(4290) <= b;
    layer0_outputs(4291) <= a or b;
    layer0_outputs(4292) <= a or b;
    layer0_outputs(4293) <= not (a xor b);
    layer0_outputs(4294) <= a xor b;
    layer0_outputs(4295) <= b;
    layer0_outputs(4296) <= not a;
    layer0_outputs(4297) <= a or b;
    layer0_outputs(4298) <= not (a xor b);
    layer0_outputs(4299) <= not a;
    layer0_outputs(4300) <= not (a xor b);
    layer0_outputs(4301) <= not b;
    layer0_outputs(4302) <= not (a or b);
    layer0_outputs(4303) <= '1';
    layer0_outputs(4304) <= '0';
    layer0_outputs(4305) <= b;
    layer0_outputs(4306) <= not a;
    layer0_outputs(4307) <= not b or a;
    layer0_outputs(4308) <= b;
    layer0_outputs(4309) <= a and not b;
    layer0_outputs(4310) <= '0';
    layer0_outputs(4311) <= not b;
    layer0_outputs(4312) <= not b;
    layer0_outputs(4313) <= a;
    layer0_outputs(4314) <= not b or a;
    layer0_outputs(4315) <= a and not b;
    layer0_outputs(4316) <= a and b;
    layer0_outputs(4317) <= not (a xor b);
    layer0_outputs(4318) <= not a or b;
    layer0_outputs(4319) <= not (a xor b);
    layer0_outputs(4320) <= a and not b;
    layer0_outputs(4321) <= a or b;
    layer0_outputs(4322) <= a or b;
    layer0_outputs(4323) <= '1';
    layer0_outputs(4324) <= not b;
    layer0_outputs(4325) <= '1';
    layer0_outputs(4326) <= not (a or b);
    layer0_outputs(4327) <= not a or b;
    layer0_outputs(4328) <= b and not a;
    layer0_outputs(4329) <= not (a and b);
    layer0_outputs(4330) <= not b;
    layer0_outputs(4331) <= '0';
    layer0_outputs(4332) <= not a or b;
    layer0_outputs(4333) <= a xor b;
    layer0_outputs(4334) <= not a;
    layer0_outputs(4335) <= not (a and b);
    layer0_outputs(4336) <= not (a or b);
    layer0_outputs(4337) <= b;
    layer0_outputs(4338) <= a and b;
    layer0_outputs(4339) <= a and b;
    layer0_outputs(4340) <= a and b;
    layer0_outputs(4341) <= not b;
    layer0_outputs(4342) <= a xor b;
    layer0_outputs(4343) <= not (a xor b);
    layer0_outputs(4344) <= a and b;
    layer0_outputs(4345) <= not b;
    layer0_outputs(4346) <= a;
    layer0_outputs(4347) <= a;
    layer0_outputs(4348) <= a or b;
    layer0_outputs(4349) <= not (a xor b);
    layer0_outputs(4350) <= a and not b;
    layer0_outputs(4351) <= not (a and b);
    layer0_outputs(4352) <= a;
    layer0_outputs(4353) <= a xor b;
    layer0_outputs(4354) <= a and b;
    layer0_outputs(4355) <= a and b;
    layer0_outputs(4356) <= a and not b;
    layer0_outputs(4357) <= a and b;
    layer0_outputs(4358) <= not (a or b);
    layer0_outputs(4359) <= b and not a;
    layer0_outputs(4360) <= not (a or b);
    layer0_outputs(4361) <= a or b;
    layer0_outputs(4362) <= a;
    layer0_outputs(4363) <= '0';
    layer0_outputs(4364) <= b and not a;
    layer0_outputs(4365) <= a and not b;
    layer0_outputs(4366) <= not (a or b);
    layer0_outputs(4367) <= not a or b;
    layer0_outputs(4368) <= '1';
    layer0_outputs(4369) <= a or b;
    layer0_outputs(4370) <= a and b;
    layer0_outputs(4371) <= b;
    layer0_outputs(4372) <= not (a or b);
    layer0_outputs(4373) <= not (a xor b);
    layer0_outputs(4374) <= b;
    layer0_outputs(4375) <= not a or b;
    layer0_outputs(4376) <= not b;
    layer0_outputs(4377) <= not (a or b);
    layer0_outputs(4378) <= '1';
    layer0_outputs(4379) <= a;
    layer0_outputs(4380) <= b and not a;
    layer0_outputs(4381) <= b;
    layer0_outputs(4382) <= a or b;
    layer0_outputs(4383) <= a or b;
    layer0_outputs(4384) <= not b;
    layer0_outputs(4385) <= a;
    layer0_outputs(4386) <= not b;
    layer0_outputs(4387) <= not a;
    layer0_outputs(4388) <= a xor b;
    layer0_outputs(4389) <= '0';
    layer0_outputs(4390) <= not (a or b);
    layer0_outputs(4391) <= a and not b;
    layer0_outputs(4392) <= '1';
    layer0_outputs(4393) <= not a;
    layer0_outputs(4394) <= not b or a;
    layer0_outputs(4395) <= not b or a;
    layer0_outputs(4396) <= a and b;
    layer0_outputs(4397) <= a xor b;
    layer0_outputs(4398) <= not (a or b);
    layer0_outputs(4399) <= not (a xor b);
    layer0_outputs(4400) <= not (a and b);
    layer0_outputs(4401) <= not (a xor b);
    layer0_outputs(4402) <= a and not b;
    layer0_outputs(4403) <= not b or a;
    layer0_outputs(4404) <= not b;
    layer0_outputs(4405) <= a and b;
    layer0_outputs(4406) <= '0';
    layer0_outputs(4407) <= not b or a;
    layer0_outputs(4408) <= b and not a;
    layer0_outputs(4409) <= not a;
    layer0_outputs(4410) <= not b;
    layer0_outputs(4411) <= not (a or b);
    layer0_outputs(4412) <= not (a xor b);
    layer0_outputs(4413) <= not b;
    layer0_outputs(4414) <= not (a or b);
    layer0_outputs(4415) <= a or b;
    layer0_outputs(4416) <= a or b;
    layer0_outputs(4417) <= a and not b;
    layer0_outputs(4418) <= not b;
    layer0_outputs(4419) <= '1';
    layer0_outputs(4420) <= a;
    layer0_outputs(4421) <= not a or b;
    layer0_outputs(4422) <= a xor b;
    layer0_outputs(4423) <= b and not a;
    layer0_outputs(4424) <= a or b;
    layer0_outputs(4425) <= a or b;
    layer0_outputs(4426) <= b and not a;
    layer0_outputs(4427) <= b and not a;
    layer0_outputs(4428) <= not a or b;
    layer0_outputs(4429) <= a and b;
    layer0_outputs(4430) <= a and not b;
    layer0_outputs(4431) <= not (a or b);
    layer0_outputs(4432) <= b;
    layer0_outputs(4433) <= not (a or b);
    layer0_outputs(4434) <= a;
    layer0_outputs(4435) <= a xor b;
    layer0_outputs(4436) <= a or b;
    layer0_outputs(4437) <= a or b;
    layer0_outputs(4438) <= not (a and b);
    layer0_outputs(4439) <= b;
    layer0_outputs(4440) <= not b;
    layer0_outputs(4441) <= a and not b;
    layer0_outputs(4442) <= b and not a;
    layer0_outputs(4443) <= a;
    layer0_outputs(4444) <= a xor b;
    layer0_outputs(4445) <= a or b;
    layer0_outputs(4446) <= b and not a;
    layer0_outputs(4447) <= a or b;
    layer0_outputs(4448) <= not b;
    layer0_outputs(4449) <= not a;
    layer0_outputs(4450) <= not b or a;
    layer0_outputs(4451) <= not b or a;
    layer0_outputs(4452) <= a and b;
    layer0_outputs(4453) <= a or b;
    layer0_outputs(4454) <= a xor b;
    layer0_outputs(4455) <= '1';
    layer0_outputs(4456) <= not b;
    layer0_outputs(4457) <= a;
    layer0_outputs(4458) <= '1';
    layer0_outputs(4459) <= not b;
    layer0_outputs(4460) <= not (a and b);
    layer0_outputs(4461) <= '0';
    layer0_outputs(4462) <= not b;
    layer0_outputs(4463) <= not b or a;
    layer0_outputs(4464) <= not (a and b);
    layer0_outputs(4465) <= not b or a;
    layer0_outputs(4466) <= b;
    layer0_outputs(4467) <= a;
    layer0_outputs(4468) <= not b;
    layer0_outputs(4469) <= a or b;
    layer0_outputs(4470) <= b;
    layer0_outputs(4471) <= not a;
    layer0_outputs(4472) <= not (a xor b);
    layer0_outputs(4473) <= '1';
    layer0_outputs(4474) <= not a;
    layer0_outputs(4475) <= not a;
    layer0_outputs(4476) <= a or b;
    layer0_outputs(4477) <= a xor b;
    layer0_outputs(4478) <= b and not a;
    layer0_outputs(4479) <= a or b;
    layer0_outputs(4480) <= not b;
    layer0_outputs(4481) <= a and not b;
    layer0_outputs(4482) <= not (a and b);
    layer0_outputs(4483) <= a xor b;
    layer0_outputs(4484) <= '0';
    layer0_outputs(4485) <= not (a and b);
    layer0_outputs(4486) <= not a or b;
    layer0_outputs(4487) <= a or b;
    layer0_outputs(4488) <= not (a or b);
    layer0_outputs(4489) <= not (a or b);
    layer0_outputs(4490) <= '1';
    layer0_outputs(4491) <= a and not b;
    layer0_outputs(4492) <= not (a or b);
    layer0_outputs(4493) <= not a;
    layer0_outputs(4494) <= not b;
    layer0_outputs(4495) <= '0';
    layer0_outputs(4496) <= b and not a;
    layer0_outputs(4497) <= a and not b;
    layer0_outputs(4498) <= a;
    layer0_outputs(4499) <= not b;
    layer0_outputs(4500) <= a and b;
    layer0_outputs(4501) <= b and not a;
    layer0_outputs(4502) <= a or b;
    layer0_outputs(4503) <= a and not b;
    layer0_outputs(4504) <= not a;
    layer0_outputs(4505) <= b;
    layer0_outputs(4506) <= not (a or b);
    layer0_outputs(4507) <= a and not b;
    layer0_outputs(4508) <= b;
    layer0_outputs(4509) <= not (a and b);
    layer0_outputs(4510) <= a or b;
    layer0_outputs(4511) <= a or b;
    layer0_outputs(4512) <= not a or b;
    layer0_outputs(4513) <= not a or b;
    layer0_outputs(4514) <= not a or b;
    layer0_outputs(4515) <= a;
    layer0_outputs(4516) <= a and not b;
    layer0_outputs(4517) <= not b;
    layer0_outputs(4518) <= not a or b;
    layer0_outputs(4519) <= not a;
    layer0_outputs(4520) <= not (a xor b);
    layer0_outputs(4521) <= not a or b;
    layer0_outputs(4522) <= b;
    layer0_outputs(4523) <= a or b;
    layer0_outputs(4524) <= not (a xor b);
    layer0_outputs(4525) <= not b or a;
    layer0_outputs(4526) <= b and not a;
    layer0_outputs(4527) <= not (a xor b);
    layer0_outputs(4528) <= a;
    layer0_outputs(4529) <= not (a xor b);
    layer0_outputs(4530) <= not (a xor b);
    layer0_outputs(4531) <= '0';
    layer0_outputs(4532) <= a and b;
    layer0_outputs(4533) <= not b;
    layer0_outputs(4534) <= a and b;
    layer0_outputs(4535) <= a;
    layer0_outputs(4536) <= a;
    layer0_outputs(4537) <= not (a or b);
    layer0_outputs(4538) <= not (a and b);
    layer0_outputs(4539) <= not (a or b);
    layer0_outputs(4540) <= b and not a;
    layer0_outputs(4541) <= a;
    layer0_outputs(4542) <= a or b;
    layer0_outputs(4543) <= '1';
    layer0_outputs(4544) <= b and not a;
    layer0_outputs(4545) <= a and not b;
    layer0_outputs(4546) <= not (a and b);
    layer0_outputs(4547) <= not b or a;
    layer0_outputs(4548) <= a;
    layer0_outputs(4549) <= '0';
    layer0_outputs(4550) <= not b;
    layer0_outputs(4551) <= '1';
    layer0_outputs(4552) <= not b or a;
    layer0_outputs(4553) <= a xor b;
    layer0_outputs(4554) <= a and b;
    layer0_outputs(4555) <= b;
    layer0_outputs(4556) <= a or b;
    layer0_outputs(4557) <= not b;
    layer0_outputs(4558) <= not a or b;
    layer0_outputs(4559) <= a or b;
    layer0_outputs(4560) <= not b;
    layer0_outputs(4561) <= not a or b;
    layer0_outputs(4562) <= '0';
    layer0_outputs(4563) <= a xor b;
    layer0_outputs(4564) <= a;
    layer0_outputs(4565) <= not (a or b);
    layer0_outputs(4566) <= not a;
    layer0_outputs(4567) <= a;
    layer0_outputs(4568) <= not a or b;
    layer0_outputs(4569) <= a or b;
    layer0_outputs(4570) <= b and not a;
    layer0_outputs(4571) <= not a or b;
    layer0_outputs(4572) <= not a or b;
    layer0_outputs(4573) <= not b;
    layer0_outputs(4574) <= not b or a;
    layer0_outputs(4575) <= a and b;
    layer0_outputs(4576) <= not a;
    layer0_outputs(4577) <= not b;
    layer0_outputs(4578) <= not (a or b);
    layer0_outputs(4579) <= not (a or b);
    layer0_outputs(4580) <= a;
    layer0_outputs(4581) <= '0';
    layer0_outputs(4582) <= not (a and b);
    layer0_outputs(4583) <= a;
    layer0_outputs(4584) <= not (a or b);
    layer0_outputs(4585) <= not b;
    layer0_outputs(4586) <= a or b;
    layer0_outputs(4587) <= not (a and b);
    layer0_outputs(4588) <= not b;
    layer0_outputs(4589) <= not (a or b);
    layer0_outputs(4590) <= not a or b;
    layer0_outputs(4591) <= a and b;
    layer0_outputs(4592) <= a or b;
    layer0_outputs(4593) <= '1';
    layer0_outputs(4594) <= a or b;
    layer0_outputs(4595) <= b;
    layer0_outputs(4596) <= a and not b;
    layer0_outputs(4597) <= a and b;
    layer0_outputs(4598) <= a xor b;
    layer0_outputs(4599) <= a xor b;
    layer0_outputs(4600) <= b and not a;
    layer0_outputs(4601) <= '0';
    layer0_outputs(4602) <= not b;
    layer0_outputs(4603) <= '0';
    layer0_outputs(4604) <= not (a or b);
    layer0_outputs(4605) <= not (a xor b);
    layer0_outputs(4606) <= a and not b;
    layer0_outputs(4607) <= b;
    layer0_outputs(4608) <= a xor b;
    layer0_outputs(4609) <= not a;
    layer0_outputs(4610) <= b;
    layer0_outputs(4611) <= not a or b;
    layer0_outputs(4612) <= not a or b;
    layer0_outputs(4613) <= a or b;
    layer0_outputs(4614) <= b and not a;
    layer0_outputs(4615) <= not (a xor b);
    layer0_outputs(4616) <= not b or a;
    layer0_outputs(4617) <= b and not a;
    layer0_outputs(4618) <= a;
    layer0_outputs(4619) <= not a;
    layer0_outputs(4620) <= a and not b;
    layer0_outputs(4621) <= not (a xor b);
    layer0_outputs(4622) <= not b or a;
    layer0_outputs(4623) <= '1';
    layer0_outputs(4624) <= not b or a;
    layer0_outputs(4625) <= a or b;
    layer0_outputs(4626) <= not a;
    layer0_outputs(4627) <= not a or b;
    layer0_outputs(4628) <= a and not b;
    layer0_outputs(4629) <= not b or a;
    layer0_outputs(4630) <= b;
    layer0_outputs(4631) <= b and not a;
    layer0_outputs(4632) <= a;
    layer0_outputs(4633) <= a and not b;
    layer0_outputs(4634) <= not (a xor b);
    layer0_outputs(4635) <= b;
    layer0_outputs(4636) <= not (a xor b);
    layer0_outputs(4637) <= b;
    layer0_outputs(4638) <= not b;
    layer0_outputs(4639) <= not (a and b);
    layer0_outputs(4640) <= a xor b;
    layer0_outputs(4641) <= a and b;
    layer0_outputs(4642) <= not b or a;
    layer0_outputs(4643) <= a and not b;
    layer0_outputs(4644) <= a;
    layer0_outputs(4645) <= not (a or b);
    layer0_outputs(4646) <= a xor b;
    layer0_outputs(4647) <= not (a or b);
    layer0_outputs(4648) <= a and b;
    layer0_outputs(4649) <= b and not a;
    layer0_outputs(4650) <= b and not a;
    layer0_outputs(4651) <= not a or b;
    layer0_outputs(4652) <= not (a and b);
    layer0_outputs(4653) <= a and b;
    layer0_outputs(4654) <= b and not a;
    layer0_outputs(4655) <= not (a or b);
    layer0_outputs(4656) <= not b or a;
    layer0_outputs(4657) <= not b or a;
    layer0_outputs(4658) <= a and b;
    layer0_outputs(4659) <= not (a and b);
    layer0_outputs(4660) <= not a;
    layer0_outputs(4661) <= not (a xor b);
    layer0_outputs(4662) <= '0';
    layer0_outputs(4663) <= a xor b;
    layer0_outputs(4664) <= not a;
    layer0_outputs(4665) <= not b or a;
    layer0_outputs(4666) <= a xor b;
    layer0_outputs(4667) <= b and not a;
    layer0_outputs(4668) <= not (a and b);
    layer0_outputs(4669) <= b;
    layer0_outputs(4670) <= b;
    layer0_outputs(4671) <= not (a or b);
    layer0_outputs(4672) <= not b;
    layer0_outputs(4673) <= a xor b;
    layer0_outputs(4674) <= a or b;
    layer0_outputs(4675) <= '0';
    layer0_outputs(4676) <= a xor b;
    layer0_outputs(4677) <= not (a xor b);
    layer0_outputs(4678) <= '0';
    layer0_outputs(4679) <= '1';
    layer0_outputs(4680) <= not (a and b);
    layer0_outputs(4681) <= not (a and b);
    layer0_outputs(4682) <= not (a or b);
    layer0_outputs(4683) <= a;
    layer0_outputs(4684) <= not b or a;
    layer0_outputs(4685) <= a and b;
    layer0_outputs(4686) <= not a;
    layer0_outputs(4687) <= b and not a;
    layer0_outputs(4688) <= b and not a;
    layer0_outputs(4689) <= a and not b;
    layer0_outputs(4690) <= not (a or b);
    layer0_outputs(4691) <= a or b;
    layer0_outputs(4692) <= a;
    layer0_outputs(4693) <= a;
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= a xor b;
    layer0_outputs(4696) <= '0';
    layer0_outputs(4697) <= '0';
    layer0_outputs(4698) <= not b or a;
    layer0_outputs(4699) <= a xor b;
    layer0_outputs(4700) <= not (a or b);
    layer0_outputs(4701) <= a;
    layer0_outputs(4702) <= not (a or b);
    layer0_outputs(4703) <= a or b;
    layer0_outputs(4704) <= a and not b;
    layer0_outputs(4705) <= b;
    layer0_outputs(4706) <= a xor b;
    layer0_outputs(4707) <= b and not a;
    layer0_outputs(4708) <= not (a and b);
    layer0_outputs(4709) <= a;
    layer0_outputs(4710) <= not a;
    layer0_outputs(4711) <= not a or b;
    layer0_outputs(4712) <= '1';
    layer0_outputs(4713) <= not (a xor b);
    layer0_outputs(4714) <= a or b;
    layer0_outputs(4715) <= a xor b;
    layer0_outputs(4716) <= b and not a;
    layer0_outputs(4717) <= not a or b;
    layer0_outputs(4718) <= not a or b;
    layer0_outputs(4719) <= '0';
    layer0_outputs(4720) <= not (a and b);
    layer0_outputs(4721) <= b;
    layer0_outputs(4722) <= not a or b;
    layer0_outputs(4723) <= not b or a;
    layer0_outputs(4724) <= not b;
    layer0_outputs(4725) <= not (a or b);
    layer0_outputs(4726) <= not (a xor b);
    layer0_outputs(4727) <= a xor b;
    layer0_outputs(4728) <= '1';
    layer0_outputs(4729) <= not (a or b);
    layer0_outputs(4730) <= not a or b;
    layer0_outputs(4731) <= b and not a;
    layer0_outputs(4732) <= not (a xor b);
    layer0_outputs(4733) <= not (a xor b);
    layer0_outputs(4734) <= not b or a;
    layer0_outputs(4735) <= '0';
    layer0_outputs(4736) <= not (a or b);
    layer0_outputs(4737) <= b;
    layer0_outputs(4738) <= b;
    layer0_outputs(4739) <= a and b;
    layer0_outputs(4740) <= a and b;
    layer0_outputs(4741) <= b;
    layer0_outputs(4742) <= not (a or b);
    layer0_outputs(4743) <= not (a xor b);
    layer0_outputs(4744) <= b and not a;
    layer0_outputs(4745) <= not (a or b);
    layer0_outputs(4746) <= a and not b;
    layer0_outputs(4747) <= not a or b;
    layer0_outputs(4748) <= b;
    layer0_outputs(4749) <= not (a and b);
    layer0_outputs(4750) <= not (a or b);
    layer0_outputs(4751) <= not (a and b);
    layer0_outputs(4752) <= b;
    layer0_outputs(4753) <= b and not a;
    layer0_outputs(4754) <= a;
    layer0_outputs(4755) <= b;
    layer0_outputs(4756) <= a;
    layer0_outputs(4757) <= a;
    layer0_outputs(4758) <= not a or b;
    layer0_outputs(4759) <= not (a or b);
    layer0_outputs(4760) <= b;
    layer0_outputs(4761) <= '1';
    layer0_outputs(4762) <= not (a or b);
    layer0_outputs(4763) <= not b or a;
    layer0_outputs(4764) <= not (a or b);
    layer0_outputs(4765) <= '0';
    layer0_outputs(4766) <= a and not b;
    layer0_outputs(4767) <= '1';
    layer0_outputs(4768) <= not a or b;
    layer0_outputs(4769) <= '1';
    layer0_outputs(4770) <= b and not a;
    layer0_outputs(4771) <= not a;
    layer0_outputs(4772) <= not (a or b);
    layer0_outputs(4773) <= not a or b;
    layer0_outputs(4774) <= a;
    layer0_outputs(4775) <= not (a and b);
    layer0_outputs(4776) <= not (a xor b);
    layer0_outputs(4777) <= a;
    layer0_outputs(4778) <= not b or a;
    layer0_outputs(4779) <= '0';
    layer0_outputs(4780) <= a and b;
    layer0_outputs(4781) <= a xor b;
    layer0_outputs(4782) <= b;
    layer0_outputs(4783) <= '1';
    layer0_outputs(4784) <= a and b;
    layer0_outputs(4785) <= a xor b;
    layer0_outputs(4786) <= a or b;
    layer0_outputs(4787) <= not b or a;
    layer0_outputs(4788) <= not b;
    layer0_outputs(4789) <= not a or b;
    layer0_outputs(4790) <= not a;
    layer0_outputs(4791) <= '0';
    layer0_outputs(4792) <= b and not a;
    layer0_outputs(4793) <= a and b;
    layer0_outputs(4794) <= not (a xor b);
    layer0_outputs(4795) <= a and not b;
    layer0_outputs(4796) <= a;
    layer0_outputs(4797) <= not a;
    layer0_outputs(4798) <= '0';
    layer0_outputs(4799) <= a;
    layer0_outputs(4800) <= a or b;
    layer0_outputs(4801) <= a or b;
    layer0_outputs(4802) <= a xor b;
    layer0_outputs(4803) <= not b or a;
    layer0_outputs(4804) <= a and not b;
    layer0_outputs(4805) <= not (a xor b);
    layer0_outputs(4806) <= '0';
    layer0_outputs(4807) <= b;
    layer0_outputs(4808) <= a and not b;
    layer0_outputs(4809) <= '0';
    layer0_outputs(4810) <= not a or b;
    layer0_outputs(4811) <= a or b;
    layer0_outputs(4812) <= a and not b;
    layer0_outputs(4813) <= not a;
    layer0_outputs(4814) <= not a;
    layer0_outputs(4815) <= not (a or b);
    layer0_outputs(4816) <= '0';
    layer0_outputs(4817) <= a and b;
    layer0_outputs(4818) <= not a;
    layer0_outputs(4819) <= b and not a;
    layer0_outputs(4820) <= b and not a;
    layer0_outputs(4821) <= not (a or b);
    layer0_outputs(4822) <= not a;
    layer0_outputs(4823) <= not a or b;
    layer0_outputs(4824) <= not (a and b);
    layer0_outputs(4825) <= b;
    layer0_outputs(4826) <= not (a xor b);
    layer0_outputs(4827) <= a and not b;
    layer0_outputs(4828) <= a xor b;
    layer0_outputs(4829) <= not a or b;
    layer0_outputs(4830) <= not b;
    layer0_outputs(4831) <= a or b;
    layer0_outputs(4832) <= b and not a;
    layer0_outputs(4833) <= a xor b;
    layer0_outputs(4834) <= a and b;
    layer0_outputs(4835) <= b and not a;
    layer0_outputs(4836) <= not b;
    layer0_outputs(4837) <= a and not b;
    layer0_outputs(4838) <= a and b;
    layer0_outputs(4839) <= a or b;
    layer0_outputs(4840) <= not b or a;
    layer0_outputs(4841) <= a or b;
    layer0_outputs(4842) <= not b;
    layer0_outputs(4843) <= b;
    layer0_outputs(4844) <= a and b;
    layer0_outputs(4845) <= b and not a;
    layer0_outputs(4846) <= b;
    layer0_outputs(4847) <= b;
    layer0_outputs(4848) <= a and b;
    layer0_outputs(4849) <= a xor b;
    layer0_outputs(4850) <= b and not a;
    layer0_outputs(4851) <= '0';
    layer0_outputs(4852) <= not (a or b);
    layer0_outputs(4853) <= not b;
    layer0_outputs(4854) <= a or b;
    layer0_outputs(4855) <= a or b;
    layer0_outputs(4856) <= a or b;
    layer0_outputs(4857) <= not b or a;
    layer0_outputs(4858) <= not (a or b);
    layer0_outputs(4859) <= a xor b;
    layer0_outputs(4860) <= not b;
    layer0_outputs(4861) <= not a;
    layer0_outputs(4862) <= not (a xor b);
    layer0_outputs(4863) <= '0';
    layer0_outputs(4864) <= b;
    layer0_outputs(4865) <= '1';
    layer0_outputs(4866) <= not (a or b);
    layer0_outputs(4867) <= a;
    layer0_outputs(4868) <= not (a xor b);
    layer0_outputs(4869) <= b;
    layer0_outputs(4870) <= not a or b;
    layer0_outputs(4871) <= a and not b;
    layer0_outputs(4872) <= not b or a;
    layer0_outputs(4873) <= not a;
    layer0_outputs(4874) <= not (a or b);
    layer0_outputs(4875) <= not a or b;
    layer0_outputs(4876) <= not (a and b);
    layer0_outputs(4877) <= a and b;
    layer0_outputs(4878) <= a or b;
    layer0_outputs(4879) <= a and not b;
    layer0_outputs(4880) <= not a;
    layer0_outputs(4881) <= not a or b;
    layer0_outputs(4882) <= not b;
    layer0_outputs(4883) <= b and not a;
    layer0_outputs(4884) <= b;
    layer0_outputs(4885) <= not (a or b);
    layer0_outputs(4886) <= not (a xor b);
    layer0_outputs(4887) <= not (a xor b);
    layer0_outputs(4888) <= b and not a;
    layer0_outputs(4889) <= a and not b;
    layer0_outputs(4890) <= '0';
    layer0_outputs(4891) <= not (a xor b);
    layer0_outputs(4892) <= a and not b;
    layer0_outputs(4893) <= a and not b;
    layer0_outputs(4894) <= b;
    layer0_outputs(4895) <= b;
    layer0_outputs(4896) <= a xor b;
    layer0_outputs(4897) <= not (a and b);
    layer0_outputs(4898) <= a and not b;
    layer0_outputs(4899) <= '1';
    layer0_outputs(4900) <= a or b;
    layer0_outputs(4901) <= a;
    layer0_outputs(4902) <= not (a xor b);
    layer0_outputs(4903) <= '0';
    layer0_outputs(4904) <= not a;
    layer0_outputs(4905) <= b;
    layer0_outputs(4906) <= not (a xor b);
    layer0_outputs(4907) <= b and not a;
    layer0_outputs(4908) <= not b;
    layer0_outputs(4909) <= not a or b;
    layer0_outputs(4910) <= b;
    layer0_outputs(4911) <= not b;
    layer0_outputs(4912) <= not (a or b);
    layer0_outputs(4913) <= a or b;
    layer0_outputs(4914) <= b and not a;
    layer0_outputs(4915) <= not a or b;
    layer0_outputs(4916) <= a xor b;
    layer0_outputs(4917) <= a xor b;
    layer0_outputs(4918) <= not b;
    layer0_outputs(4919) <= a;
    layer0_outputs(4920) <= a;
    layer0_outputs(4921) <= b and not a;
    layer0_outputs(4922) <= not (a or b);
    layer0_outputs(4923) <= a xor b;
    layer0_outputs(4924) <= a;
    layer0_outputs(4925) <= a or b;
    layer0_outputs(4926) <= a xor b;
    layer0_outputs(4927) <= a and b;
    layer0_outputs(4928) <= '1';
    layer0_outputs(4929) <= a or b;
    layer0_outputs(4930) <= not a;
    layer0_outputs(4931) <= not b or a;
    layer0_outputs(4932) <= a and not b;
    layer0_outputs(4933) <= not a or b;
    layer0_outputs(4934) <= a or b;
    layer0_outputs(4935) <= a or b;
    layer0_outputs(4936) <= not (a or b);
    layer0_outputs(4937) <= b and not a;
    layer0_outputs(4938) <= a xor b;
    layer0_outputs(4939) <= a and not b;
    layer0_outputs(4940) <= not a or b;
    layer0_outputs(4941) <= '1';
    layer0_outputs(4942) <= not b;
    layer0_outputs(4943) <= not a;
    layer0_outputs(4944) <= a and not b;
    layer0_outputs(4945) <= not b;
    layer0_outputs(4946) <= b;
    layer0_outputs(4947) <= not (a or b);
    layer0_outputs(4948) <= b;
    layer0_outputs(4949) <= not a or b;
    layer0_outputs(4950) <= not (a or b);
    layer0_outputs(4951) <= '0';
    layer0_outputs(4952) <= not b;
    layer0_outputs(4953) <= b;
    layer0_outputs(4954) <= b;
    layer0_outputs(4955) <= '0';
    layer0_outputs(4956) <= not (a or b);
    layer0_outputs(4957) <= '1';
    layer0_outputs(4958) <= a and not b;
    layer0_outputs(4959) <= a or b;
    layer0_outputs(4960) <= not (a xor b);
    layer0_outputs(4961) <= not (a or b);
    layer0_outputs(4962) <= a and b;
    layer0_outputs(4963) <= not a or b;
    layer0_outputs(4964) <= not a;
    layer0_outputs(4965) <= a or b;
    layer0_outputs(4966) <= '0';
    layer0_outputs(4967) <= not a;
    layer0_outputs(4968) <= not a;
    layer0_outputs(4969) <= not a;
    layer0_outputs(4970) <= not b or a;
    layer0_outputs(4971) <= not b or a;
    layer0_outputs(4972) <= a and b;
    layer0_outputs(4973) <= not b;
    layer0_outputs(4974) <= b;
    layer0_outputs(4975) <= '1';
    layer0_outputs(4976) <= a;
    layer0_outputs(4977) <= b and not a;
    layer0_outputs(4978) <= b and not a;
    layer0_outputs(4979) <= a or b;
    layer0_outputs(4980) <= not b;
    layer0_outputs(4981) <= a and b;
    layer0_outputs(4982) <= not b or a;
    layer0_outputs(4983) <= '1';
    layer0_outputs(4984) <= b and not a;
    layer0_outputs(4985) <= '0';
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= a;
    layer0_outputs(4988) <= not (a xor b);
    layer0_outputs(4989) <= not b;
    layer0_outputs(4990) <= a or b;
    layer0_outputs(4991) <= not a;
    layer0_outputs(4992) <= a;
    layer0_outputs(4993) <= not a;
    layer0_outputs(4994) <= not (a or b);
    layer0_outputs(4995) <= not b or a;
    layer0_outputs(4996) <= a and b;
    layer0_outputs(4997) <= a or b;
    layer0_outputs(4998) <= not a or b;
    layer0_outputs(4999) <= a;
    layer0_outputs(5000) <= not (a and b);
    layer0_outputs(5001) <= not (a and b);
    layer0_outputs(5002) <= a or b;
    layer0_outputs(5003) <= not a or b;
    layer0_outputs(5004) <= '0';
    layer0_outputs(5005) <= a or b;
    layer0_outputs(5006) <= not b or a;
    layer0_outputs(5007) <= not b;
    layer0_outputs(5008) <= not b or a;
    layer0_outputs(5009) <= not a or b;
    layer0_outputs(5010) <= '1';
    layer0_outputs(5011) <= a or b;
    layer0_outputs(5012) <= a or b;
    layer0_outputs(5013) <= b;
    layer0_outputs(5014) <= not (a or b);
    layer0_outputs(5015) <= not b or a;
    layer0_outputs(5016) <= not b or a;
    layer0_outputs(5017) <= not (a and b);
    layer0_outputs(5018) <= a and b;
    layer0_outputs(5019) <= a;
    layer0_outputs(5020) <= not b;
    layer0_outputs(5021) <= b and not a;
    layer0_outputs(5022) <= a xor b;
    layer0_outputs(5023) <= not a or b;
    layer0_outputs(5024) <= a xor b;
    layer0_outputs(5025) <= not a;
    layer0_outputs(5026) <= a and not b;
    layer0_outputs(5027) <= not a or b;
    layer0_outputs(5028) <= a;
    layer0_outputs(5029) <= not (a and b);
    layer0_outputs(5030) <= not (a xor b);
    layer0_outputs(5031) <= b;
    layer0_outputs(5032) <= a and not b;
    layer0_outputs(5033) <= not (a or b);
    layer0_outputs(5034) <= b;
    layer0_outputs(5035) <= not (a xor b);
    layer0_outputs(5036) <= not (a and b);
    layer0_outputs(5037) <= a or b;
    layer0_outputs(5038) <= not (a or b);
    layer0_outputs(5039) <= b and not a;
    layer0_outputs(5040) <= not a;
    layer0_outputs(5041) <= a or b;
    layer0_outputs(5042) <= not b or a;
    layer0_outputs(5043) <= a xor b;
    layer0_outputs(5044) <= not a or b;
    layer0_outputs(5045) <= not (a xor b);
    layer0_outputs(5046) <= b;
    layer0_outputs(5047) <= a and b;
    layer0_outputs(5048) <= not (a or b);
    layer0_outputs(5049) <= not (a or b);
    layer0_outputs(5050) <= not b;
    layer0_outputs(5051) <= a xor b;
    layer0_outputs(5052) <= not (a or b);
    layer0_outputs(5053) <= b;
    layer0_outputs(5054) <= not b or a;
    layer0_outputs(5055) <= a;
    layer0_outputs(5056) <= a and b;
    layer0_outputs(5057) <= b;
    layer0_outputs(5058) <= not b;
    layer0_outputs(5059) <= '1';
    layer0_outputs(5060) <= a or b;
    layer0_outputs(5061) <= not a or b;
    layer0_outputs(5062) <= '1';
    layer0_outputs(5063) <= '0';
    layer0_outputs(5064) <= b;
    layer0_outputs(5065) <= a or b;
    layer0_outputs(5066) <= a and not b;
    layer0_outputs(5067) <= '0';
    layer0_outputs(5068) <= a;
    layer0_outputs(5069) <= a xor b;
    layer0_outputs(5070) <= not (a or b);
    layer0_outputs(5071) <= not (a xor b);
    layer0_outputs(5072) <= not (a xor b);
    layer0_outputs(5073) <= '1';
    layer0_outputs(5074) <= not b;
    layer0_outputs(5075) <= b;
    layer0_outputs(5076) <= a;
    layer0_outputs(5077) <= not a;
    layer0_outputs(5078) <= not (a xor b);
    layer0_outputs(5079) <= '0';
    layer0_outputs(5080) <= not a or b;
    layer0_outputs(5081) <= not (a xor b);
    layer0_outputs(5082) <= not (a xor b);
    layer0_outputs(5083) <= a;
    layer0_outputs(5084) <= not (a xor b);
    layer0_outputs(5085) <= a;
    layer0_outputs(5086) <= a xor b;
    layer0_outputs(5087) <= a or b;
    layer0_outputs(5088) <= b and not a;
    layer0_outputs(5089) <= a xor b;
    layer0_outputs(5090) <= not a or b;
    layer0_outputs(5091) <= b;
    layer0_outputs(5092) <= a and b;
    layer0_outputs(5093) <= not (a xor b);
    layer0_outputs(5094) <= b;
    layer0_outputs(5095) <= b;
    layer0_outputs(5096) <= not (a and b);
    layer0_outputs(5097) <= a;
    layer0_outputs(5098) <= b;
    layer0_outputs(5099) <= a or b;
    layer0_outputs(5100) <= a or b;
    layer0_outputs(5101) <= '0';
    layer0_outputs(5102) <= not a or b;
    layer0_outputs(5103) <= not b or a;
    layer0_outputs(5104) <= not (a or b);
    layer0_outputs(5105) <= not b or a;
    layer0_outputs(5106) <= a xor b;
    layer0_outputs(5107) <= not b;
    layer0_outputs(5108) <= a and b;
    layer0_outputs(5109) <= a;
    layer0_outputs(5110) <= '1';
    layer0_outputs(5111) <= not b;
    layer0_outputs(5112) <= not b or a;
    layer0_outputs(5113) <= not a or b;
    layer0_outputs(5114) <= not a or b;
    layer0_outputs(5115) <= a xor b;
    layer0_outputs(5116) <= not b or a;
    layer0_outputs(5117) <= a;
    layer0_outputs(5118) <= a or b;
    layer0_outputs(5119) <= not b;
    layer0_outputs(5120) <= a;
    layer0_outputs(5121) <= not (a and b);
    layer0_outputs(5122) <= '0';
    layer0_outputs(5123) <= not b;
    layer0_outputs(5124) <= not b;
    layer0_outputs(5125) <= not a;
    layer0_outputs(5126) <= '1';
    layer0_outputs(5127) <= not (a and b);
    layer0_outputs(5128) <= not (a and b);
    layer0_outputs(5129) <= b;
    layer0_outputs(5130) <= b and not a;
    layer0_outputs(5131) <= not a or b;
    layer0_outputs(5132) <= not (a or b);
    layer0_outputs(5133) <= a or b;
    layer0_outputs(5134) <= not b or a;
    layer0_outputs(5135) <= a xor b;
    layer0_outputs(5136) <= b and not a;
    layer0_outputs(5137) <= not a;
    layer0_outputs(5138) <= not a or b;
    layer0_outputs(5139) <= not b or a;
    layer0_outputs(5140) <= '1';
    layer0_outputs(5141) <= '0';
    layer0_outputs(5142) <= a and b;
    layer0_outputs(5143) <= not (a xor b);
    layer0_outputs(5144) <= a;
    layer0_outputs(5145) <= a or b;
    layer0_outputs(5146) <= not a or b;
    layer0_outputs(5147) <= a;
    layer0_outputs(5148) <= a;
    layer0_outputs(5149) <= b;
    layer0_outputs(5150) <= a and not b;
    layer0_outputs(5151) <= not b or a;
    layer0_outputs(5152) <= a and b;
    layer0_outputs(5153) <= a;
    layer0_outputs(5154) <= not (a and b);
    layer0_outputs(5155) <= a or b;
    layer0_outputs(5156) <= a and b;
    layer0_outputs(5157) <= not a or b;
    layer0_outputs(5158) <= not a;
    layer0_outputs(5159) <= a or b;
    layer0_outputs(5160) <= a and not b;
    layer0_outputs(5161) <= not a;
    layer0_outputs(5162) <= b;
    layer0_outputs(5163) <= not (a and b);
    layer0_outputs(5164) <= not (a or b);
    layer0_outputs(5165) <= a;
    layer0_outputs(5166) <= b;
    layer0_outputs(5167) <= a xor b;
    layer0_outputs(5168) <= a or b;
    layer0_outputs(5169) <= b;
    layer0_outputs(5170) <= a and b;
    layer0_outputs(5171) <= not (a or b);
    layer0_outputs(5172) <= a or b;
    layer0_outputs(5173) <= not b or a;
    layer0_outputs(5174) <= not (a or b);
    layer0_outputs(5175) <= '1';
    layer0_outputs(5176) <= a;
    layer0_outputs(5177) <= '1';
    layer0_outputs(5178) <= b and not a;
    layer0_outputs(5179) <= '1';
    layer0_outputs(5180) <= a;
    layer0_outputs(5181) <= a;
    layer0_outputs(5182) <= a and not b;
    layer0_outputs(5183) <= a and b;
    layer0_outputs(5184) <= a xor b;
    layer0_outputs(5185) <= a xor b;
    layer0_outputs(5186) <= a and not b;
    layer0_outputs(5187) <= not a;
    layer0_outputs(5188) <= '0';
    layer0_outputs(5189) <= a or b;
    layer0_outputs(5190) <= '1';
    layer0_outputs(5191) <= b;
    layer0_outputs(5192) <= not b;
    layer0_outputs(5193) <= not a;
    layer0_outputs(5194) <= a xor b;
    layer0_outputs(5195) <= b;
    layer0_outputs(5196) <= not a;
    layer0_outputs(5197) <= not (a or b);
    layer0_outputs(5198) <= a xor b;
    layer0_outputs(5199) <= a or b;
    layer0_outputs(5200) <= b;
    layer0_outputs(5201) <= not (a or b);
    layer0_outputs(5202) <= a and not b;
    layer0_outputs(5203) <= '0';
    layer0_outputs(5204) <= a;
    layer0_outputs(5205) <= '0';
    layer0_outputs(5206) <= not a or b;
    layer0_outputs(5207) <= '0';
    layer0_outputs(5208) <= b;
    layer0_outputs(5209) <= a;
    layer0_outputs(5210) <= a or b;
    layer0_outputs(5211) <= a and b;
    layer0_outputs(5212) <= b and not a;
    layer0_outputs(5213) <= '0';
    layer0_outputs(5214) <= a xor b;
    layer0_outputs(5215) <= a;
    layer0_outputs(5216) <= a or b;
    layer0_outputs(5217) <= a or b;
    layer0_outputs(5218) <= not b;
    layer0_outputs(5219) <= a and b;
    layer0_outputs(5220) <= b and not a;
    layer0_outputs(5221) <= a and not b;
    layer0_outputs(5222) <= not b or a;
    layer0_outputs(5223) <= a or b;
    layer0_outputs(5224) <= a or b;
    layer0_outputs(5225) <= not (a or b);
    layer0_outputs(5226) <= a and b;
    layer0_outputs(5227) <= '0';
    layer0_outputs(5228) <= b and not a;
    layer0_outputs(5229) <= a and not b;
    layer0_outputs(5230) <= not b;
    layer0_outputs(5231) <= not a or b;
    layer0_outputs(5232) <= not b or a;
    layer0_outputs(5233) <= not (a or b);
    layer0_outputs(5234) <= b and not a;
    layer0_outputs(5235) <= b and not a;
    layer0_outputs(5236) <= a xor b;
    layer0_outputs(5237) <= not (a or b);
    layer0_outputs(5238) <= a or b;
    layer0_outputs(5239) <= not (a or b);
    layer0_outputs(5240) <= not b or a;
    layer0_outputs(5241) <= a;
    layer0_outputs(5242) <= a;
    layer0_outputs(5243) <= not b;
    layer0_outputs(5244) <= a and b;
    layer0_outputs(5245) <= a;
    layer0_outputs(5246) <= a and not b;
    layer0_outputs(5247) <= not b or a;
    layer0_outputs(5248) <= a and b;
    layer0_outputs(5249) <= a xor b;
    layer0_outputs(5250) <= not b;
    layer0_outputs(5251) <= not (a and b);
    layer0_outputs(5252) <= b;
    layer0_outputs(5253) <= not b or a;
    layer0_outputs(5254) <= b and not a;
    layer0_outputs(5255) <= b;
    layer0_outputs(5256) <= b;
    layer0_outputs(5257) <= not (a and b);
    layer0_outputs(5258) <= b;
    layer0_outputs(5259) <= '0';
    layer0_outputs(5260) <= not (a xor b);
    layer0_outputs(5261) <= '0';
    layer0_outputs(5262) <= not (a or b);
    layer0_outputs(5263) <= not (a or b);
    layer0_outputs(5264) <= a and not b;
    layer0_outputs(5265) <= a or b;
    layer0_outputs(5266) <= not b;
    layer0_outputs(5267) <= b and not a;
    layer0_outputs(5268) <= not b;
    layer0_outputs(5269) <= not (a and b);
    layer0_outputs(5270) <= a or b;
    layer0_outputs(5271) <= a and not b;
    layer0_outputs(5272) <= not a or b;
    layer0_outputs(5273) <= '1';
    layer0_outputs(5274) <= not (a or b);
    layer0_outputs(5275) <= a xor b;
    layer0_outputs(5276) <= not (a and b);
    layer0_outputs(5277) <= not b or a;
    layer0_outputs(5278) <= not a or b;
    layer0_outputs(5279) <= not (a xor b);
    layer0_outputs(5280) <= '0';
    layer0_outputs(5281) <= not (a and b);
    layer0_outputs(5282) <= b;
    layer0_outputs(5283) <= b;
    layer0_outputs(5284) <= not (a and b);
    layer0_outputs(5285) <= b and not a;
    layer0_outputs(5286) <= b;
    layer0_outputs(5287) <= not (a or b);
    layer0_outputs(5288) <= not (a or b);
    layer0_outputs(5289) <= not a or b;
    layer0_outputs(5290) <= a or b;
    layer0_outputs(5291) <= a and not b;
    layer0_outputs(5292) <= '0';
    layer0_outputs(5293) <= a and not b;
    layer0_outputs(5294) <= a xor b;
    layer0_outputs(5295) <= not (a xor b);
    layer0_outputs(5296) <= not b or a;
    layer0_outputs(5297) <= not (a or b);
    layer0_outputs(5298) <= not a or b;
    layer0_outputs(5299) <= not b;
    layer0_outputs(5300) <= b;
    layer0_outputs(5301) <= '0';
    layer0_outputs(5302) <= a;
    layer0_outputs(5303) <= '0';
    layer0_outputs(5304) <= a and not b;
    layer0_outputs(5305) <= not a or b;
    layer0_outputs(5306) <= b and not a;
    layer0_outputs(5307) <= a xor b;
    layer0_outputs(5308) <= a or b;
    layer0_outputs(5309) <= a;
    layer0_outputs(5310) <= not b;
    layer0_outputs(5311) <= not a;
    layer0_outputs(5312) <= not (a or b);
    layer0_outputs(5313) <= a or b;
    layer0_outputs(5314) <= not (a and b);
    layer0_outputs(5315) <= not a or b;
    layer0_outputs(5316) <= not a or b;
    layer0_outputs(5317) <= a or b;
    layer0_outputs(5318) <= a xor b;
    layer0_outputs(5319) <= '1';
    layer0_outputs(5320) <= a and not b;
    layer0_outputs(5321) <= not a or b;
    layer0_outputs(5322) <= a and b;
    layer0_outputs(5323) <= not (a or b);
    layer0_outputs(5324) <= b;
    layer0_outputs(5325) <= '0';
    layer0_outputs(5326) <= not b;
    layer0_outputs(5327) <= b;
    layer0_outputs(5328) <= not (a or b);
    layer0_outputs(5329) <= '1';
    layer0_outputs(5330) <= a;
    layer0_outputs(5331) <= a or b;
    layer0_outputs(5332) <= a and not b;
    layer0_outputs(5333) <= a xor b;
    layer0_outputs(5334) <= '1';
    layer0_outputs(5335) <= not a or b;
    layer0_outputs(5336) <= not a or b;
    layer0_outputs(5337) <= not (a xor b);
    layer0_outputs(5338) <= a or b;
    layer0_outputs(5339) <= b and not a;
    layer0_outputs(5340) <= a;
    layer0_outputs(5341) <= not b or a;
    layer0_outputs(5342) <= not (a and b);
    layer0_outputs(5343) <= not (a and b);
    layer0_outputs(5344) <= a or b;
    layer0_outputs(5345) <= '1';
    layer0_outputs(5346) <= a or b;
    layer0_outputs(5347) <= a and b;
    layer0_outputs(5348) <= a and b;
    layer0_outputs(5349) <= a or b;
    layer0_outputs(5350) <= b;
    layer0_outputs(5351) <= not (a and b);
    layer0_outputs(5352) <= '0';
    layer0_outputs(5353) <= a and b;
    layer0_outputs(5354) <= b;
    layer0_outputs(5355) <= not (a or b);
    layer0_outputs(5356) <= a;
    layer0_outputs(5357) <= not (a or b);
    layer0_outputs(5358) <= not (a xor b);
    layer0_outputs(5359) <= not (a or b);
    layer0_outputs(5360) <= '0';
    layer0_outputs(5361) <= not b;
    layer0_outputs(5362) <= not (a xor b);
    layer0_outputs(5363) <= not a;
    layer0_outputs(5364) <= not (a xor b);
    layer0_outputs(5365) <= not (a xor b);
    layer0_outputs(5366) <= '1';
    layer0_outputs(5367) <= not b or a;
    layer0_outputs(5368) <= a xor b;
    layer0_outputs(5369) <= not a or b;
    layer0_outputs(5370) <= not b;
    layer0_outputs(5371) <= not a;
    layer0_outputs(5372) <= not (a or b);
    layer0_outputs(5373) <= not (a and b);
    layer0_outputs(5374) <= '0';
    layer0_outputs(5375) <= not (a xor b);
    layer0_outputs(5376) <= a or b;
    layer0_outputs(5377) <= not (a or b);
    layer0_outputs(5378) <= '1';
    layer0_outputs(5379) <= not b;
    layer0_outputs(5380) <= '0';
    layer0_outputs(5381) <= not b or a;
    layer0_outputs(5382) <= a;
    layer0_outputs(5383) <= not b;
    layer0_outputs(5384) <= not a or b;
    layer0_outputs(5385) <= b and not a;
    layer0_outputs(5386) <= a xor b;
    layer0_outputs(5387) <= not a;
    layer0_outputs(5388) <= not (a or b);
    layer0_outputs(5389) <= b and not a;
    layer0_outputs(5390) <= a and b;
    layer0_outputs(5391) <= a;
    layer0_outputs(5392) <= a xor b;
    layer0_outputs(5393) <= not (a and b);
    layer0_outputs(5394) <= not a or b;
    layer0_outputs(5395) <= a and not b;
    layer0_outputs(5396) <= b and not a;
    layer0_outputs(5397) <= a xor b;
    layer0_outputs(5398) <= b;
    layer0_outputs(5399) <= not a;
    layer0_outputs(5400) <= b;
    layer0_outputs(5401) <= not b or a;
    layer0_outputs(5402) <= a or b;
    layer0_outputs(5403) <= b and not a;
    layer0_outputs(5404) <= not (a and b);
    layer0_outputs(5405) <= not (a and b);
    layer0_outputs(5406) <= a xor b;
    layer0_outputs(5407) <= a xor b;
    layer0_outputs(5408) <= b;
    layer0_outputs(5409) <= a or b;
    layer0_outputs(5410) <= not b;
    layer0_outputs(5411) <= b;
    layer0_outputs(5412) <= not b or a;
    layer0_outputs(5413) <= not (a and b);
    layer0_outputs(5414) <= '0';
    layer0_outputs(5415) <= a or b;
    layer0_outputs(5416) <= a or b;
    layer0_outputs(5417) <= a and b;
    layer0_outputs(5418) <= not (a and b);
    layer0_outputs(5419) <= a or b;
    layer0_outputs(5420) <= not (a xor b);
    layer0_outputs(5421) <= not b or a;
    layer0_outputs(5422) <= not b or a;
    layer0_outputs(5423) <= a and not b;
    layer0_outputs(5424) <= not (a or b);
    layer0_outputs(5425) <= not b or a;
    layer0_outputs(5426) <= not b or a;
    layer0_outputs(5427) <= b and not a;
    layer0_outputs(5428) <= b;
    layer0_outputs(5429) <= not b;
    layer0_outputs(5430) <= not (a or b);
    layer0_outputs(5431) <= not b;
    layer0_outputs(5432) <= a;
    layer0_outputs(5433) <= a and b;
    layer0_outputs(5434) <= not b;
    layer0_outputs(5435) <= a or b;
    layer0_outputs(5436) <= not a;
    layer0_outputs(5437) <= not b or a;
    layer0_outputs(5438) <= a;
    layer0_outputs(5439) <= b;
    layer0_outputs(5440) <= '0';
    layer0_outputs(5441) <= a or b;
    layer0_outputs(5442) <= not (a xor b);
    layer0_outputs(5443) <= not b or a;
    layer0_outputs(5444) <= not a or b;
    layer0_outputs(5445) <= not b;
    layer0_outputs(5446) <= not b or a;
    layer0_outputs(5447) <= not b;
    layer0_outputs(5448) <= not b;
    layer0_outputs(5449) <= not (a and b);
    layer0_outputs(5450) <= a;
    layer0_outputs(5451) <= not a;
    layer0_outputs(5452) <= a and b;
    layer0_outputs(5453) <= b;
    layer0_outputs(5454) <= not (a and b);
    layer0_outputs(5455) <= a or b;
    layer0_outputs(5456) <= not (a or b);
    layer0_outputs(5457) <= not (a or b);
    layer0_outputs(5458) <= not a;
    layer0_outputs(5459) <= a or b;
    layer0_outputs(5460) <= not (a and b);
    layer0_outputs(5461) <= b;
    layer0_outputs(5462) <= not (a and b);
    layer0_outputs(5463) <= not b;
    layer0_outputs(5464) <= a and not b;
    layer0_outputs(5465) <= a and not b;
    layer0_outputs(5466) <= not (a xor b);
    layer0_outputs(5467) <= a and b;
    layer0_outputs(5468) <= not (a and b);
    layer0_outputs(5469) <= not (a and b);
    layer0_outputs(5470) <= b;
    layer0_outputs(5471) <= a xor b;
    layer0_outputs(5472) <= a or b;
    layer0_outputs(5473) <= not (a and b);
    layer0_outputs(5474) <= a and not b;
    layer0_outputs(5475) <= a or b;
    layer0_outputs(5476) <= a xor b;
    layer0_outputs(5477) <= a and b;
    layer0_outputs(5478) <= b and not a;
    layer0_outputs(5479) <= a and not b;
    layer0_outputs(5480) <= b and not a;
    layer0_outputs(5481) <= b and not a;
    layer0_outputs(5482) <= not b;
    layer0_outputs(5483) <= not a;
    layer0_outputs(5484) <= not a;
    layer0_outputs(5485) <= '1';
    layer0_outputs(5486) <= not b or a;
    layer0_outputs(5487) <= a or b;
    layer0_outputs(5488) <= not b;
    layer0_outputs(5489) <= not a;
    layer0_outputs(5490) <= a or b;
    layer0_outputs(5491) <= a and not b;
    layer0_outputs(5492) <= not b;
    layer0_outputs(5493) <= a and not b;
    layer0_outputs(5494) <= not a;
    layer0_outputs(5495) <= not (a and b);
    layer0_outputs(5496) <= not b;
    layer0_outputs(5497) <= not a or b;
    layer0_outputs(5498) <= b and not a;
    layer0_outputs(5499) <= '1';
    layer0_outputs(5500) <= '0';
    layer0_outputs(5501) <= not (a xor b);
    layer0_outputs(5502) <= '1';
    layer0_outputs(5503) <= not a;
    layer0_outputs(5504) <= not b;
    layer0_outputs(5505) <= b and not a;
    layer0_outputs(5506) <= not (a or b);
    layer0_outputs(5507) <= a and b;
    layer0_outputs(5508) <= a and not b;
    layer0_outputs(5509) <= not b or a;
    layer0_outputs(5510) <= not (a or b);
    layer0_outputs(5511) <= a;
    layer0_outputs(5512) <= not a;
    layer0_outputs(5513) <= a;
    layer0_outputs(5514) <= a;
    layer0_outputs(5515) <= not (a or b);
    layer0_outputs(5516) <= a or b;
    layer0_outputs(5517) <= a or b;
    layer0_outputs(5518) <= a and not b;
    layer0_outputs(5519) <= not (a xor b);
    layer0_outputs(5520) <= a and not b;
    layer0_outputs(5521) <= b;
    layer0_outputs(5522) <= a and b;
    layer0_outputs(5523) <= not a;
    layer0_outputs(5524) <= a xor b;
    layer0_outputs(5525) <= not a;
    layer0_outputs(5526) <= not (a or b);
    layer0_outputs(5527) <= a;
    layer0_outputs(5528) <= a xor b;
    layer0_outputs(5529) <= not (a or b);
    layer0_outputs(5530) <= not b;
    layer0_outputs(5531) <= not a or b;
    layer0_outputs(5532) <= b and not a;
    layer0_outputs(5533) <= '0';
    layer0_outputs(5534) <= not a or b;
    layer0_outputs(5535) <= not a or b;
    layer0_outputs(5536) <= not (a and b);
    layer0_outputs(5537) <= b;
    layer0_outputs(5538) <= a and b;
    layer0_outputs(5539) <= a or b;
    layer0_outputs(5540) <= not a or b;
    layer0_outputs(5541) <= a or b;
    layer0_outputs(5542) <= not b or a;
    layer0_outputs(5543) <= not b or a;
    layer0_outputs(5544) <= not (a or b);
    layer0_outputs(5545) <= '0';
    layer0_outputs(5546) <= not a or b;
    layer0_outputs(5547) <= not b;
    layer0_outputs(5548) <= not b or a;
    layer0_outputs(5549) <= not b or a;
    layer0_outputs(5550) <= '0';
    layer0_outputs(5551) <= a or b;
    layer0_outputs(5552) <= '0';
    layer0_outputs(5553) <= '1';
    layer0_outputs(5554) <= not b;
    layer0_outputs(5555) <= a and not b;
    layer0_outputs(5556) <= a;
    layer0_outputs(5557) <= a;
    layer0_outputs(5558) <= '0';
    layer0_outputs(5559) <= b and not a;
    layer0_outputs(5560) <= not a;
    layer0_outputs(5561) <= a xor b;
    layer0_outputs(5562) <= not b;
    layer0_outputs(5563) <= not b or a;
    layer0_outputs(5564) <= not (a xor b);
    layer0_outputs(5565) <= b;
    layer0_outputs(5566) <= a xor b;
    layer0_outputs(5567) <= b;
    layer0_outputs(5568) <= a;
    layer0_outputs(5569) <= not a or b;
    layer0_outputs(5570) <= a and not b;
    layer0_outputs(5571) <= b;
    layer0_outputs(5572) <= not (a xor b);
    layer0_outputs(5573) <= b and not a;
    layer0_outputs(5574) <= a xor b;
    layer0_outputs(5575) <= not (a or b);
    layer0_outputs(5576) <= not (a xor b);
    layer0_outputs(5577) <= not (a or b);
    layer0_outputs(5578) <= a;
    layer0_outputs(5579) <= not (a xor b);
    layer0_outputs(5580) <= a and not b;
    layer0_outputs(5581) <= a and not b;
    layer0_outputs(5582) <= b;
    layer0_outputs(5583) <= a and b;
    layer0_outputs(5584) <= not a;
    layer0_outputs(5585) <= b;
    layer0_outputs(5586) <= b;
    layer0_outputs(5587) <= not b or a;
    layer0_outputs(5588) <= a and b;
    layer0_outputs(5589) <= not a or b;
    layer0_outputs(5590) <= not b;
    layer0_outputs(5591) <= a xor b;
    layer0_outputs(5592) <= not a or b;
    layer0_outputs(5593) <= a and b;
    layer0_outputs(5594) <= not (a or b);
    layer0_outputs(5595) <= b and not a;
    layer0_outputs(5596) <= a;
    layer0_outputs(5597) <= not a or b;
    layer0_outputs(5598) <= not a or b;
    layer0_outputs(5599) <= '0';
    layer0_outputs(5600) <= a or b;
    layer0_outputs(5601) <= a;
    layer0_outputs(5602) <= '1';
    layer0_outputs(5603) <= not (a and b);
    layer0_outputs(5604) <= b and not a;
    layer0_outputs(5605) <= a;
    layer0_outputs(5606) <= b;
    layer0_outputs(5607) <= not (a xor b);
    layer0_outputs(5608) <= not (a xor b);
    layer0_outputs(5609) <= not (a and b);
    layer0_outputs(5610) <= b and not a;
    layer0_outputs(5611) <= not b or a;
    layer0_outputs(5612) <= not a or b;
    layer0_outputs(5613) <= not b;
    layer0_outputs(5614) <= '1';
    layer0_outputs(5615) <= not b;
    layer0_outputs(5616) <= a and not b;
    layer0_outputs(5617) <= a;
    layer0_outputs(5618) <= '1';
    layer0_outputs(5619) <= '1';
    layer0_outputs(5620) <= not (a xor b);
    layer0_outputs(5621) <= a or b;
    layer0_outputs(5622) <= a or b;
    layer0_outputs(5623) <= not b or a;
    layer0_outputs(5624) <= not a or b;
    layer0_outputs(5625) <= a and not b;
    layer0_outputs(5626) <= '0';
    layer0_outputs(5627) <= not b;
    layer0_outputs(5628) <= a and b;
    layer0_outputs(5629) <= b and not a;
    layer0_outputs(5630) <= not a;
    layer0_outputs(5631) <= a and b;
    layer0_outputs(5632) <= not a or b;
    layer0_outputs(5633) <= not a;
    layer0_outputs(5634) <= '0';
    layer0_outputs(5635) <= b;
    layer0_outputs(5636) <= not (a xor b);
    layer0_outputs(5637) <= a and not b;
    layer0_outputs(5638) <= not (a xor b);
    layer0_outputs(5639) <= not a or b;
    layer0_outputs(5640) <= '0';
    layer0_outputs(5641) <= '1';
    layer0_outputs(5642) <= not (a or b);
    layer0_outputs(5643) <= not b;
    layer0_outputs(5644) <= a;
    layer0_outputs(5645) <= a xor b;
    layer0_outputs(5646) <= a;
    layer0_outputs(5647) <= b;
    layer0_outputs(5648) <= a xor b;
    layer0_outputs(5649) <= not (a or b);
    layer0_outputs(5650) <= not (a or b);
    layer0_outputs(5651) <= '0';
    layer0_outputs(5652) <= a or b;
    layer0_outputs(5653) <= a xor b;
    layer0_outputs(5654) <= not a;
    layer0_outputs(5655) <= a xor b;
    layer0_outputs(5656) <= not a;
    layer0_outputs(5657) <= not b;
    layer0_outputs(5658) <= '1';
    layer0_outputs(5659) <= b and not a;
    layer0_outputs(5660) <= '1';
    layer0_outputs(5661) <= not (a or b);
    layer0_outputs(5662) <= not a;
    layer0_outputs(5663) <= '1';
    layer0_outputs(5664) <= not (a xor b);
    layer0_outputs(5665) <= a and not b;
    layer0_outputs(5666) <= a;
    layer0_outputs(5667) <= not b or a;
    layer0_outputs(5668) <= not (a and b);
    layer0_outputs(5669) <= a and not b;
    layer0_outputs(5670) <= b and not a;
    layer0_outputs(5671) <= not (a or b);
    layer0_outputs(5672) <= not (a and b);
    layer0_outputs(5673) <= not (a or b);
    layer0_outputs(5674) <= b and not a;
    layer0_outputs(5675) <= b and not a;
    layer0_outputs(5676) <= not (a xor b);
    layer0_outputs(5677) <= not b;
    layer0_outputs(5678) <= not b or a;
    layer0_outputs(5679) <= not a;
    layer0_outputs(5680) <= not a;
    layer0_outputs(5681) <= not b;
    layer0_outputs(5682) <= a and b;
    layer0_outputs(5683) <= not a or b;
    layer0_outputs(5684) <= '0';
    layer0_outputs(5685) <= not a or b;
    layer0_outputs(5686) <= not a;
    layer0_outputs(5687) <= not (a or b);
    layer0_outputs(5688) <= b;
    layer0_outputs(5689) <= a and not b;
    layer0_outputs(5690) <= a;
    layer0_outputs(5691) <= not a;
    layer0_outputs(5692) <= a and not b;
    layer0_outputs(5693) <= a or b;
    layer0_outputs(5694) <= a xor b;
    layer0_outputs(5695) <= not (a xor b);
    layer0_outputs(5696) <= not (a or b);
    layer0_outputs(5697) <= not (a xor b);
    layer0_outputs(5698) <= a xor b;
    layer0_outputs(5699) <= a;
    layer0_outputs(5700) <= not (a or b);
    layer0_outputs(5701) <= a and not b;
    layer0_outputs(5702) <= a;
    layer0_outputs(5703) <= b and not a;
    layer0_outputs(5704) <= b and not a;
    layer0_outputs(5705) <= not (a xor b);
    layer0_outputs(5706) <= a or b;
    layer0_outputs(5707) <= a and not b;
    layer0_outputs(5708) <= not (a and b);
    layer0_outputs(5709) <= a and b;
    layer0_outputs(5710) <= a;
    layer0_outputs(5711) <= '1';
    layer0_outputs(5712) <= a or b;
    layer0_outputs(5713) <= a or b;
    layer0_outputs(5714) <= a xor b;
    layer0_outputs(5715) <= not a or b;
    layer0_outputs(5716) <= not (a or b);
    layer0_outputs(5717) <= not a;
    layer0_outputs(5718) <= not a or b;
    layer0_outputs(5719) <= a or b;
    layer0_outputs(5720) <= a xor b;
    layer0_outputs(5721) <= a or b;
    layer0_outputs(5722) <= '1';
    layer0_outputs(5723) <= a and b;
    layer0_outputs(5724) <= a;
    layer0_outputs(5725) <= a;
    layer0_outputs(5726) <= b;
    layer0_outputs(5727) <= a and not b;
    layer0_outputs(5728) <= not a;
    layer0_outputs(5729) <= not (a xor b);
    layer0_outputs(5730) <= not (a xor b);
    layer0_outputs(5731) <= not (a or b);
    layer0_outputs(5732) <= b and not a;
    layer0_outputs(5733) <= a and b;
    layer0_outputs(5734) <= not b;
    layer0_outputs(5735) <= not b;
    layer0_outputs(5736) <= a and not b;
    layer0_outputs(5737) <= a or b;
    layer0_outputs(5738) <= '1';
    layer0_outputs(5739) <= '0';
    layer0_outputs(5740) <= a and b;
    layer0_outputs(5741) <= a;
    layer0_outputs(5742) <= not a or b;
    layer0_outputs(5743) <= not b or a;
    layer0_outputs(5744) <= not (a or b);
    layer0_outputs(5745) <= not b or a;
    layer0_outputs(5746) <= not a or b;
    layer0_outputs(5747) <= not b;
    layer0_outputs(5748) <= a or b;
    layer0_outputs(5749) <= a and not b;
    layer0_outputs(5750) <= not (a and b);
    layer0_outputs(5751) <= a or b;
    layer0_outputs(5752) <= b;
    layer0_outputs(5753) <= '1';
    layer0_outputs(5754) <= not a;
    layer0_outputs(5755) <= a;
    layer0_outputs(5756) <= a;
    layer0_outputs(5757) <= not (a xor b);
    layer0_outputs(5758) <= not a or b;
    layer0_outputs(5759) <= not (a or b);
    layer0_outputs(5760) <= not (a or b);
    layer0_outputs(5761) <= not a;
    layer0_outputs(5762) <= b and not a;
    layer0_outputs(5763) <= a and not b;
    layer0_outputs(5764) <= b and not a;
    layer0_outputs(5765) <= '0';
    layer0_outputs(5766) <= a and b;
    layer0_outputs(5767) <= a and not b;
    layer0_outputs(5768) <= not a or b;
    layer0_outputs(5769) <= b;
    layer0_outputs(5770) <= '1';
    layer0_outputs(5771) <= a and not b;
    layer0_outputs(5772) <= a or b;
    layer0_outputs(5773) <= not (a or b);
    layer0_outputs(5774) <= not a or b;
    layer0_outputs(5775) <= not (a or b);
    layer0_outputs(5776) <= a and b;
    layer0_outputs(5777) <= a xor b;
    layer0_outputs(5778) <= not b;
    layer0_outputs(5779) <= a and b;
    layer0_outputs(5780) <= a xor b;
    layer0_outputs(5781) <= not (a xor b);
    layer0_outputs(5782) <= not (a xor b);
    layer0_outputs(5783) <= a or b;
    layer0_outputs(5784) <= a xor b;
    layer0_outputs(5785) <= not (a xor b);
    layer0_outputs(5786) <= not (a xor b);
    layer0_outputs(5787) <= not b;
    layer0_outputs(5788) <= a and not b;
    layer0_outputs(5789) <= b and not a;
    layer0_outputs(5790) <= not (a xor b);
    layer0_outputs(5791) <= b;
    layer0_outputs(5792) <= not b;
    layer0_outputs(5793) <= a;
    layer0_outputs(5794) <= a and b;
    layer0_outputs(5795) <= not a or b;
    layer0_outputs(5796) <= b and not a;
    layer0_outputs(5797) <= a and b;
    layer0_outputs(5798) <= a xor b;
    layer0_outputs(5799) <= a and not b;
    layer0_outputs(5800) <= a xor b;
    layer0_outputs(5801) <= not b;
    layer0_outputs(5802) <= a;
    layer0_outputs(5803) <= '0';
    layer0_outputs(5804) <= not b;
    layer0_outputs(5805) <= not (a or b);
    layer0_outputs(5806) <= a or b;
    layer0_outputs(5807) <= not (a xor b);
    layer0_outputs(5808) <= not b;
    layer0_outputs(5809) <= b;
    layer0_outputs(5810) <= a or b;
    layer0_outputs(5811) <= not b;
    layer0_outputs(5812) <= b;
    layer0_outputs(5813) <= a;
    layer0_outputs(5814) <= b;
    layer0_outputs(5815) <= b;
    layer0_outputs(5816) <= a and b;
    layer0_outputs(5817) <= not b or a;
    layer0_outputs(5818) <= not (a xor b);
    layer0_outputs(5819) <= not b;
    layer0_outputs(5820) <= b;
    layer0_outputs(5821) <= not (a xor b);
    layer0_outputs(5822) <= b;
    layer0_outputs(5823) <= a;
    layer0_outputs(5824) <= a;
    layer0_outputs(5825) <= not a or b;
    layer0_outputs(5826) <= a xor b;
    layer0_outputs(5827) <= a and b;
    layer0_outputs(5828) <= b;
    layer0_outputs(5829) <= a and b;
    layer0_outputs(5830) <= not a or b;
    layer0_outputs(5831) <= b and not a;
    layer0_outputs(5832) <= b;
    layer0_outputs(5833) <= '0';
    layer0_outputs(5834) <= not (a or b);
    layer0_outputs(5835) <= not (a or b);
    layer0_outputs(5836) <= b;
    layer0_outputs(5837) <= a and not b;
    layer0_outputs(5838) <= b;
    layer0_outputs(5839) <= not a or b;
    layer0_outputs(5840) <= not (a and b);
    layer0_outputs(5841) <= not (a and b);
    layer0_outputs(5842) <= not b;
    layer0_outputs(5843) <= not b;
    layer0_outputs(5844) <= a xor b;
    layer0_outputs(5845) <= not (a and b);
    layer0_outputs(5846) <= not b or a;
    layer0_outputs(5847) <= a or b;
    layer0_outputs(5848) <= not a;
    layer0_outputs(5849) <= not (a or b);
    layer0_outputs(5850) <= not b;
    layer0_outputs(5851) <= '0';
    layer0_outputs(5852) <= not (a xor b);
    layer0_outputs(5853) <= not (a and b);
    layer0_outputs(5854) <= not (a or b);
    layer0_outputs(5855) <= b and not a;
    layer0_outputs(5856) <= '0';
    layer0_outputs(5857) <= not b;
    layer0_outputs(5858) <= b;
    layer0_outputs(5859) <= a;
    layer0_outputs(5860) <= '0';
    layer0_outputs(5861) <= not b;
    layer0_outputs(5862) <= not b or a;
    layer0_outputs(5863) <= not b;
    layer0_outputs(5864) <= '1';
    layer0_outputs(5865) <= a or b;
    layer0_outputs(5866) <= not b or a;
    layer0_outputs(5867) <= a xor b;
    layer0_outputs(5868) <= not (a xor b);
    layer0_outputs(5869) <= not b or a;
    layer0_outputs(5870) <= not (a xor b);
    layer0_outputs(5871) <= '1';
    layer0_outputs(5872) <= not a;
    layer0_outputs(5873) <= '1';
    layer0_outputs(5874) <= not b;
    layer0_outputs(5875) <= not a or b;
    layer0_outputs(5876) <= a and not b;
    layer0_outputs(5877) <= b;
    layer0_outputs(5878) <= a xor b;
    layer0_outputs(5879) <= not (a xor b);
    layer0_outputs(5880) <= not (a or b);
    layer0_outputs(5881) <= a;
    layer0_outputs(5882) <= b and not a;
    layer0_outputs(5883) <= a and not b;
    layer0_outputs(5884) <= b and not a;
    layer0_outputs(5885) <= a and not b;
    layer0_outputs(5886) <= a;
    layer0_outputs(5887) <= a xor b;
    layer0_outputs(5888) <= not a or b;
    layer0_outputs(5889) <= a and not b;
    layer0_outputs(5890) <= '1';
    layer0_outputs(5891) <= b;
    layer0_outputs(5892) <= '0';
    layer0_outputs(5893) <= not a or b;
    layer0_outputs(5894) <= a and not b;
    layer0_outputs(5895) <= not b or a;
    layer0_outputs(5896) <= not (a or b);
    layer0_outputs(5897) <= a or b;
    layer0_outputs(5898) <= not a or b;
    layer0_outputs(5899) <= b;
    layer0_outputs(5900) <= not (a and b);
    layer0_outputs(5901) <= not (a xor b);
    layer0_outputs(5902) <= not b or a;
    layer0_outputs(5903) <= a xor b;
    layer0_outputs(5904) <= not (a or b);
    layer0_outputs(5905) <= not a;
    layer0_outputs(5906) <= not a;
    layer0_outputs(5907) <= a or b;
    layer0_outputs(5908) <= a xor b;
    layer0_outputs(5909) <= not (a xor b);
    layer0_outputs(5910) <= '0';
    layer0_outputs(5911) <= not (a or b);
    layer0_outputs(5912) <= '0';
    layer0_outputs(5913) <= a and b;
    layer0_outputs(5914) <= not a or b;
    layer0_outputs(5915) <= not b or a;
    layer0_outputs(5916) <= a;
    layer0_outputs(5917) <= not (a xor b);
    layer0_outputs(5918) <= not b or a;
    layer0_outputs(5919) <= not (a or b);
    layer0_outputs(5920) <= not a or b;
    layer0_outputs(5921) <= not (a or b);
    layer0_outputs(5922) <= not (a xor b);
    layer0_outputs(5923) <= '0';
    layer0_outputs(5924) <= a;
    layer0_outputs(5925) <= '0';
    layer0_outputs(5926) <= not (a or b);
    layer0_outputs(5927) <= a and not b;
    layer0_outputs(5928) <= b;
    layer0_outputs(5929) <= not (a or b);
    layer0_outputs(5930) <= not b or a;
    layer0_outputs(5931) <= not a or b;
    layer0_outputs(5932) <= a;
    layer0_outputs(5933) <= a or b;
    layer0_outputs(5934) <= b and not a;
    layer0_outputs(5935) <= a xor b;
    layer0_outputs(5936) <= a;
    layer0_outputs(5937) <= not (a and b);
    layer0_outputs(5938) <= a and not b;
    layer0_outputs(5939) <= not a;
    layer0_outputs(5940) <= a or b;
    layer0_outputs(5941) <= a and not b;
    layer0_outputs(5942) <= a xor b;
    layer0_outputs(5943) <= a;
    layer0_outputs(5944) <= b;
    layer0_outputs(5945) <= not b;
    layer0_outputs(5946) <= not (a and b);
    layer0_outputs(5947) <= b;
    layer0_outputs(5948) <= not a or b;
    layer0_outputs(5949) <= '1';
    layer0_outputs(5950) <= not b;
    layer0_outputs(5951) <= a or b;
    layer0_outputs(5952) <= a and b;
    layer0_outputs(5953) <= b and not a;
    layer0_outputs(5954) <= '0';
    layer0_outputs(5955) <= a or b;
    layer0_outputs(5956) <= not (a xor b);
    layer0_outputs(5957) <= not (a and b);
    layer0_outputs(5958) <= not (a or b);
    layer0_outputs(5959) <= a xor b;
    layer0_outputs(5960) <= not (a or b);
    layer0_outputs(5961) <= a or b;
    layer0_outputs(5962) <= a;
    layer0_outputs(5963) <= a or b;
    layer0_outputs(5964) <= not a or b;
    layer0_outputs(5965) <= a;
    layer0_outputs(5966) <= a xor b;
    layer0_outputs(5967) <= not a;
    layer0_outputs(5968) <= not a or b;
    layer0_outputs(5969) <= not b or a;
    layer0_outputs(5970) <= a;
    layer0_outputs(5971) <= not (a xor b);
    layer0_outputs(5972) <= b and not a;
    layer0_outputs(5973) <= b and not a;
    layer0_outputs(5974) <= a and b;
    layer0_outputs(5975) <= a and not b;
    layer0_outputs(5976) <= a and not b;
    layer0_outputs(5977) <= not (a xor b);
    layer0_outputs(5978) <= '0';
    layer0_outputs(5979) <= not b or a;
    layer0_outputs(5980) <= not (a xor b);
    layer0_outputs(5981) <= not a;
    layer0_outputs(5982) <= '0';
    layer0_outputs(5983) <= '0';
    layer0_outputs(5984) <= not (a and b);
    layer0_outputs(5985) <= a and not b;
    layer0_outputs(5986) <= not a;
    layer0_outputs(5987) <= not a or b;
    layer0_outputs(5988) <= a and not b;
    layer0_outputs(5989) <= not (a or b);
    layer0_outputs(5990) <= b;
    layer0_outputs(5991) <= not (a or b);
    layer0_outputs(5992) <= a and not b;
    layer0_outputs(5993) <= b;
    layer0_outputs(5994) <= a;
    layer0_outputs(5995) <= '0';
    layer0_outputs(5996) <= '0';
    layer0_outputs(5997) <= a and not b;
    layer0_outputs(5998) <= not (a or b);
    layer0_outputs(5999) <= '1';
    layer0_outputs(6000) <= not (a or b);
    layer0_outputs(6001) <= not (a xor b);
    layer0_outputs(6002) <= a or b;
    layer0_outputs(6003) <= b;
    layer0_outputs(6004) <= '1';
    layer0_outputs(6005) <= not (a and b);
    layer0_outputs(6006) <= not (a xor b);
    layer0_outputs(6007) <= b;
    layer0_outputs(6008) <= not (a and b);
    layer0_outputs(6009) <= not b;
    layer0_outputs(6010) <= '1';
    layer0_outputs(6011) <= not (a or b);
    layer0_outputs(6012) <= a xor b;
    layer0_outputs(6013) <= a and not b;
    layer0_outputs(6014) <= '1';
    layer0_outputs(6015) <= not (a and b);
    layer0_outputs(6016) <= b;
    layer0_outputs(6017) <= a or b;
    layer0_outputs(6018) <= a;
    layer0_outputs(6019) <= a and not b;
    layer0_outputs(6020) <= a;
    layer0_outputs(6021) <= a xor b;
    layer0_outputs(6022) <= '1';
    layer0_outputs(6023) <= b;
    layer0_outputs(6024) <= not b or a;
    layer0_outputs(6025) <= not (a or b);
    layer0_outputs(6026) <= a;
    layer0_outputs(6027) <= '0';
    layer0_outputs(6028) <= '1';
    layer0_outputs(6029) <= not (a or b);
    layer0_outputs(6030) <= b and not a;
    layer0_outputs(6031) <= b and not a;
    layer0_outputs(6032) <= '0';
    layer0_outputs(6033) <= not (a xor b);
    layer0_outputs(6034) <= a xor b;
    layer0_outputs(6035) <= not a;
    layer0_outputs(6036) <= a or b;
    layer0_outputs(6037) <= a or b;
    layer0_outputs(6038) <= a or b;
    layer0_outputs(6039) <= not a;
    layer0_outputs(6040) <= a xor b;
    layer0_outputs(6041) <= not (a or b);
    layer0_outputs(6042) <= not b or a;
    layer0_outputs(6043) <= a xor b;
    layer0_outputs(6044) <= b;
    layer0_outputs(6045) <= not (a xor b);
    layer0_outputs(6046) <= a xor b;
    layer0_outputs(6047) <= b and not a;
    layer0_outputs(6048) <= not b;
    layer0_outputs(6049) <= not (a or b);
    layer0_outputs(6050) <= a or b;
    layer0_outputs(6051) <= not a or b;
    layer0_outputs(6052) <= not b or a;
    layer0_outputs(6053) <= not a;
    layer0_outputs(6054) <= not (a or b);
    layer0_outputs(6055) <= not (a xor b);
    layer0_outputs(6056) <= b and not a;
    layer0_outputs(6057) <= a;
    layer0_outputs(6058) <= not a;
    layer0_outputs(6059) <= a and b;
    layer0_outputs(6060) <= '1';
    layer0_outputs(6061) <= not a or b;
    layer0_outputs(6062) <= not a or b;
    layer0_outputs(6063) <= not a or b;
    layer0_outputs(6064) <= a xor b;
    layer0_outputs(6065) <= a xor b;
    layer0_outputs(6066) <= not a;
    layer0_outputs(6067) <= not (a xor b);
    layer0_outputs(6068) <= not (a and b);
    layer0_outputs(6069) <= '1';
    layer0_outputs(6070) <= a and not b;
    layer0_outputs(6071) <= a or b;
    layer0_outputs(6072) <= a and not b;
    layer0_outputs(6073) <= not (a or b);
    layer0_outputs(6074) <= a xor b;
    layer0_outputs(6075) <= not a;
    layer0_outputs(6076) <= b;
    layer0_outputs(6077) <= a xor b;
    layer0_outputs(6078) <= not a or b;
    layer0_outputs(6079) <= not b or a;
    layer0_outputs(6080) <= '0';
    layer0_outputs(6081) <= b and not a;
    layer0_outputs(6082) <= not (a or b);
    layer0_outputs(6083) <= not b or a;
    layer0_outputs(6084) <= not (a xor b);
    layer0_outputs(6085) <= not (a or b);
    layer0_outputs(6086) <= not (a or b);
    layer0_outputs(6087) <= a and not b;
    layer0_outputs(6088) <= not b or a;
    layer0_outputs(6089) <= not a;
    layer0_outputs(6090) <= a;
    layer0_outputs(6091) <= b and not a;
    layer0_outputs(6092) <= not (a or b);
    layer0_outputs(6093) <= a;
    layer0_outputs(6094) <= not (a or b);
    layer0_outputs(6095) <= not (a and b);
    layer0_outputs(6096) <= not (a and b);
    layer0_outputs(6097) <= not (a and b);
    layer0_outputs(6098) <= b and not a;
    layer0_outputs(6099) <= b;
    layer0_outputs(6100) <= a or b;
    layer0_outputs(6101) <= not a;
    layer0_outputs(6102) <= a;
    layer0_outputs(6103) <= not a or b;
    layer0_outputs(6104) <= '1';
    layer0_outputs(6105) <= '0';
    layer0_outputs(6106) <= a or b;
    layer0_outputs(6107) <= not a or b;
    layer0_outputs(6108) <= not (a or b);
    layer0_outputs(6109) <= a and not b;
    layer0_outputs(6110) <= b;
    layer0_outputs(6111) <= not (a and b);
    layer0_outputs(6112) <= not a;
    layer0_outputs(6113) <= a;
    layer0_outputs(6114) <= '1';
    layer0_outputs(6115) <= a;
    layer0_outputs(6116) <= '1';
    layer0_outputs(6117) <= a and not b;
    layer0_outputs(6118) <= not (a and b);
    layer0_outputs(6119) <= not (a xor b);
    layer0_outputs(6120) <= not a or b;
    layer0_outputs(6121) <= not (a xor b);
    layer0_outputs(6122) <= a xor b;
    layer0_outputs(6123) <= a;
    layer0_outputs(6124) <= not a;
    layer0_outputs(6125) <= b;
    layer0_outputs(6126) <= a and not b;
    layer0_outputs(6127) <= not (a or b);
    layer0_outputs(6128) <= b and not a;
    layer0_outputs(6129) <= not (a xor b);
    layer0_outputs(6130) <= not a;
    layer0_outputs(6131) <= b and not a;
    layer0_outputs(6132) <= not (a and b);
    layer0_outputs(6133) <= a;
    layer0_outputs(6134) <= not (a or b);
    layer0_outputs(6135) <= not a or b;
    layer0_outputs(6136) <= a;
    layer0_outputs(6137) <= not (a xor b);
    layer0_outputs(6138) <= a and b;
    layer0_outputs(6139) <= '0';
    layer0_outputs(6140) <= not (a xor b);
    layer0_outputs(6141) <= not (a xor b);
    layer0_outputs(6142) <= a and b;
    layer0_outputs(6143) <= '0';
    layer0_outputs(6144) <= a and not b;
    layer0_outputs(6145) <= a or b;
    layer0_outputs(6146) <= b;
    layer0_outputs(6147) <= a;
    layer0_outputs(6148) <= a and not b;
    layer0_outputs(6149) <= '1';
    layer0_outputs(6150) <= a or b;
    layer0_outputs(6151) <= not a;
    layer0_outputs(6152) <= not (a or b);
    layer0_outputs(6153) <= a and b;
    layer0_outputs(6154) <= a xor b;
    layer0_outputs(6155) <= not a or b;
    layer0_outputs(6156) <= not b;
    layer0_outputs(6157) <= not a;
    layer0_outputs(6158) <= not a;
    layer0_outputs(6159) <= a;
    layer0_outputs(6160) <= not b or a;
    layer0_outputs(6161) <= b and not a;
    layer0_outputs(6162) <= '0';
    layer0_outputs(6163) <= b;
    layer0_outputs(6164) <= a and b;
    layer0_outputs(6165) <= a or b;
    layer0_outputs(6166) <= not a or b;
    layer0_outputs(6167) <= a or b;
    layer0_outputs(6168) <= b and not a;
    layer0_outputs(6169) <= b and not a;
    layer0_outputs(6170) <= not (a and b);
    layer0_outputs(6171) <= not b;
    layer0_outputs(6172) <= a;
    layer0_outputs(6173) <= a and not b;
    layer0_outputs(6174) <= b and not a;
    layer0_outputs(6175) <= not b;
    layer0_outputs(6176) <= a xor b;
    layer0_outputs(6177) <= a or b;
    layer0_outputs(6178) <= b;
    layer0_outputs(6179) <= not b;
    layer0_outputs(6180) <= '0';
    layer0_outputs(6181) <= not (a xor b);
    layer0_outputs(6182) <= a xor b;
    layer0_outputs(6183) <= a or b;
    layer0_outputs(6184) <= not (a and b);
    layer0_outputs(6185) <= not (a or b);
    layer0_outputs(6186) <= a or b;
    layer0_outputs(6187) <= not a;
    layer0_outputs(6188) <= b and not a;
    layer0_outputs(6189) <= a and b;
    layer0_outputs(6190) <= not (a xor b);
    layer0_outputs(6191) <= b;
    layer0_outputs(6192) <= a xor b;
    layer0_outputs(6193) <= '0';
    layer0_outputs(6194) <= not a or b;
    layer0_outputs(6195) <= not a or b;
    layer0_outputs(6196) <= not a or b;
    layer0_outputs(6197) <= a or b;
    layer0_outputs(6198) <= a and b;
    layer0_outputs(6199) <= '0';
    layer0_outputs(6200) <= not (a xor b);
    layer0_outputs(6201) <= not a;
    layer0_outputs(6202) <= not b or a;
    layer0_outputs(6203) <= a xor b;
    layer0_outputs(6204) <= a and not b;
    layer0_outputs(6205) <= a xor b;
    layer0_outputs(6206) <= a and b;
    layer0_outputs(6207) <= a xor b;
    layer0_outputs(6208) <= not a or b;
    layer0_outputs(6209) <= b and not a;
    layer0_outputs(6210) <= b and not a;
    layer0_outputs(6211) <= not b;
    layer0_outputs(6212) <= not (a and b);
    layer0_outputs(6213) <= not a;
    layer0_outputs(6214) <= a and not b;
    layer0_outputs(6215) <= b;
    layer0_outputs(6216) <= not (a and b);
    layer0_outputs(6217) <= a xor b;
    layer0_outputs(6218) <= not (a or b);
    layer0_outputs(6219) <= a or b;
    layer0_outputs(6220) <= a or b;
    layer0_outputs(6221) <= a xor b;
    layer0_outputs(6222) <= a or b;
    layer0_outputs(6223) <= not (a xor b);
    layer0_outputs(6224) <= b and not a;
    layer0_outputs(6225) <= not b;
    layer0_outputs(6226) <= '0';
    layer0_outputs(6227) <= not (a and b);
    layer0_outputs(6228) <= not (a and b);
    layer0_outputs(6229) <= not (a or b);
    layer0_outputs(6230) <= a xor b;
    layer0_outputs(6231) <= not a;
    layer0_outputs(6232) <= a;
    layer0_outputs(6233) <= not a or b;
    layer0_outputs(6234) <= not b or a;
    layer0_outputs(6235) <= b and not a;
    layer0_outputs(6236) <= a;
    layer0_outputs(6237) <= not b;
    layer0_outputs(6238) <= not a;
    layer0_outputs(6239) <= b and not a;
    layer0_outputs(6240) <= a;
    layer0_outputs(6241) <= not (a xor b);
    layer0_outputs(6242) <= not b or a;
    layer0_outputs(6243) <= not (a and b);
    layer0_outputs(6244) <= not (a xor b);
    layer0_outputs(6245) <= not a;
    layer0_outputs(6246) <= not a or b;
    layer0_outputs(6247) <= not b;
    layer0_outputs(6248) <= not b;
    layer0_outputs(6249) <= '0';
    layer0_outputs(6250) <= a or b;
    layer0_outputs(6251) <= a xor b;
    layer0_outputs(6252) <= b;
    layer0_outputs(6253) <= b and not a;
    layer0_outputs(6254) <= a and not b;
    layer0_outputs(6255) <= a and b;
    layer0_outputs(6256) <= a xor b;
    layer0_outputs(6257) <= a;
    layer0_outputs(6258) <= not a;
    layer0_outputs(6259) <= not (a and b);
    layer0_outputs(6260) <= not b or a;
    layer0_outputs(6261) <= a and b;
    layer0_outputs(6262) <= a and b;
    layer0_outputs(6263) <= b;
    layer0_outputs(6264) <= not b;
    layer0_outputs(6265) <= not a or b;
    layer0_outputs(6266) <= b and not a;
    layer0_outputs(6267) <= not (a xor b);
    layer0_outputs(6268) <= not a or b;
    layer0_outputs(6269) <= b;
    layer0_outputs(6270) <= '1';
    layer0_outputs(6271) <= '0';
    layer0_outputs(6272) <= not b or a;
    layer0_outputs(6273) <= not a or b;
    layer0_outputs(6274) <= a and b;
    layer0_outputs(6275) <= not (a or b);
    layer0_outputs(6276) <= not a or b;
    layer0_outputs(6277) <= a xor b;
    layer0_outputs(6278) <= a and not b;
    layer0_outputs(6279) <= not (a or b);
    layer0_outputs(6280) <= a or b;
    layer0_outputs(6281) <= not b or a;
    layer0_outputs(6282) <= a and not b;
    layer0_outputs(6283) <= not (a or b);
    layer0_outputs(6284) <= b;
    layer0_outputs(6285) <= not (a and b);
    layer0_outputs(6286) <= a or b;
    layer0_outputs(6287) <= a xor b;
    layer0_outputs(6288) <= '0';
    layer0_outputs(6289) <= not a or b;
    layer0_outputs(6290) <= not (a or b);
    layer0_outputs(6291) <= not (a or b);
    layer0_outputs(6292) <= '1';
    layer0_outputs(6293) <= a xor b;
    layer0_outputs(6294) <= not (a xor b);
    layer0_outputs(6295) <= a;
    layer0_outputs(6296) <= not (a xor b);
    layer0_outputs(6297) <= '0';
    layer0_outputs(6298) <= a xor b;
    layer0_outputs(6299) <= not (a xor b);
    layer0_outputs(6300) <= not b;
    layer0_outputs(6301) <= a and not b;
    layer0_outputs(6302) <= a or b;
    layer0_outputs(6303) <= a or b;
    layer0_outputs(6304) <= a or b;
    layer0_outputs(6305) <= not b;
    layer0_outputs(6306) <= a and b;
    layer0_outputs(6307) <= a and b;
    layer0_outputs(6308) <= not a;
    layer0_outputs(6309) <= a and not b;
    layer0_outputs(6310) <= b;
    layer0_outputs(6311) <= a xor b;
    layer0_outputs(6312) <= not b;
    layer0_outputs(6313) <= a xor b;
    layer0_outputs(6314) <= a or b;
    layer0_outputs(6315) <= not (a or b);
    layer0_outputs(6316) <= b;
    layer0_outputs(6317) <= a and b;
    layer0_outputs(6318) <= not a or b;
    layer0_outputs(6319) <= not a or b;
    layer0_outputs(6320) <= not a or b;
    layer0_outputs(6321) <= a xor b;
    layer0_outputs(6322) <= '0';
    layer0_outputs(6323) <= a xor b;
    layer0_outputs(6324) <= '0';
    layer0_outputs(6325) <= not b;
    layer0_outputs(6326) <= not b or a;
    layer0_outputs(6327) <= not (a or b);
    layer0_outputs(6328) <= not a;
    layer0_outputs(6329) <= b and not a;
    layer0_outputs(6330) <= b and not a;
    layer0_outputs(6331) <= b;
    layer0_outputs(6332) <= not b;
    layer0_outputs(6333) <= not (a and b);
    layer0_outputs(6334) <= not b or a;
    layer0_outputs(6335) <= b;
    layer0_outputs(6336) <= b;
    layer0_outputs(6337) <= not b;
    layer0_outputs(6338) <= b;
    layer0_outputs(6339) <= not (a or b);
    layer0_outputs(6340) <= '1';
    layer0_outputs(6341) <= a and b;
    layer0_outputs(6342) <= a;
    layer0_outputs(6343) <= a or b;
    layer0_outputs(6344) <= a or b;
    layer0_outputs(6345) <= not a;
    layer0_outputs(6346) <= a;
    layer0_outputs(6347) <= b and not a;
    layer0_outputs(6348) <= b and not a;
    layer0_outputs(6349) <= a and not b;
    layer0_outputs(6350) <= not a;
    layer0_outputs(6351) <= a xor b;
    layer0_outputs(6352) <= a and not b;
    layer0_outputs(6353) <= not (a and b);
    layer0_outputs(6354) <= a and not b;
    layer0_outputs(6355) <= '0';
    layer0_outputs(6356) <= '0';
    layer0_outputs(6357) <= not b;
    layer0_outputs(6358) <= a;
    layer0_outputs(6359) <= not (a xor b);
    layer0_outputs(6360) <= a and not b;
    layer0_outputs(6361) <= '1';
    layer0_outputs(6362) <= not b or a;
    layer0_outputs(6363) <= not (a and b);
    layer0_outputs(6364) <= not a;
    layer0_outputs(6365) <= not b;
    layer0_outputs(6366) <= not (a xor b);
    layer0_outputs(6367) <= not b or a;
    layer0_outputs(6368) <= '0';
    layer0_outputs(6369) <= not (a or b);
    layer0_outputs(6370) <= not a or b;
    layer0_outputs(6371) <= not a;
    layer0_outputs(6372) <= '0';
    layer0_outputs(6373) <= a and b;
    layer0_outputs(6374) <= not (a xor b);
    layer0_outputs(6375) <= not b or a;
    layer0_outputs(6376) <= a or b;
    layer0_outputs(6377) <= not b or a;
    layer0_outputs(6378) <= not b;
    layer0_outputs(6379) <= not b or a;
    layer0_outputs(6380) <= a xor b;
    layer0_outputs(6381) <= a or b;
    layer0_outputs(6382) <= b and not a;
    layer0_outputs(6383) <= a and not b;
    layer0_outputs(6384) <= a;
    layer0_outputs(6385) <= not a or b;
    layer0_outputs(6386) <= b;
    layer0_outputs(6387) <= a;
    layer0_outputs(6388) <= a and not b;
    layer0_outputs(6389) <= a;
    layer0_outputs(6390) <= not b;
    layer0_outputs(6391) <= a xor b;
    layer0_outputs(6392) <= not (a xor b);
    layer0_outputs(6393) <= not b;
    layer0_outputs(6394) <= not b;
    layer0_outputs(6395) <= b;
    layer0_outputs(6396) <= not (a and b);
    layer0_outputs(6397) <= a and b;
    layer0_outputs(6398) <= b and not a;
    layer0_outputs(6399) <= not a or b;
    layer0_outputs(6400) <= a or b;
    layer0_outputs(6401) <= not b;
    layer0_outputs(6402) <= not b or a;
    layer0_outputs(6403) <= not a;
    layer0_outputs(6404) <= a xor b;
    layer0_outputs(6405) <= not a or b;
    layer0_outputs(6406) <= not (a or b);
    layer0_outputs(6407) <= not b or a;
    layer0_outputs(6408) <= not b;
    layer0_outputs(6409) <= b;
    layer0_outputs(6410) <= a or b;
    layer0_outputs(6411) <= b and not a;
    layer0_outputs(6412) <= not b;
    layer0_outputs(6413) <= b and not a;
    layer0_outputs(6414) <= not a;
    layer0_outputs(6415) <= not b or a;
    layer0_outputs(6416) <= '0';
    layer0_outputs(6417) <= not a;
    layer0_outputs(6418) <= not a;
    layer0_outputs(6419) <= b;
    layer0_outputs(6420) <= b and not a;
    layer0_outputs(6421) <= b and not a;
    layer0_outputs(6422) <= a or b;
    layer0_outputs(6423) <= not (a and b);
    layer0_outputs(6424) <= not b;
    layer0_outputs(6425) <= not (a and b);
    layer0_outputs(6426) <= not (a or b);
    layer0_outputs(6427) <= '0';
    layer0_outputs(6428) <= '1';
    layer0_outputs(6429) <= a xor b;
    layer0_outputs(6430) <= a or b;
    layer0_outputs(6431) <= not (a or b);
    layer0_outputs(6432) <= a and not b;
    layer0_outputs(6433) <= not a;
    layer0_outputs(6434) <= a;
    layer0_outputs(6435) <= not a;
    layer0_outputs(6436) <= not b;
    layer0_outputs(6437) <= '0';
    layer0_outputs(6438) <= b and not a;
    layer0_outputs(6439) <= a and not b;
    layer0_outputs(6440) <= b;
    layer0_outputs(6441) <= not a;
    layer0_outputs(6442) <= a;
    layer0_outputs(6443) <= b;
    layer0_outputs(6444) <= '1';
    layer0_outputs(6445) <= not a;
    layer0_outputs(6446) <= a xor b;
    layer0_outputs(6447) <= a or b;
    layer0_outputs(6448) <= b;
    layer0_outputs(6449) <= not (a or b);
    layer0_outputs(6450) <= a and not b;
    layer0_outputs(6451) <= '0';
    layer0_outputs(6452) <= not a;
    layer0_outputs(6453) <= b;
    layer0_outputs(6454) <= not (a and b);
    layer0_outputs(6455) <= not b or a;
    layer0_outputs(6456) <= a;
    layer0_outputs(6457) <= b;
    layer0_outputs(6458) <= not b or a;
    layer0_outputs(6459) <= '1';
    layer0_outputs(6460) <= not (a or b);
    layer0_outputs(6461) <= '1';
    layer0_outputs(6462) <= not (a xor b);
    layer0_outputs(6463) <= not (a or b);
    layer0_outputs(6464) <= not a or b;
    layer0_outputs(6465) <= not a or b;
    layer0_outputs(6466) <= not (a and b);
    layer0_outputs(6467) <= a or b;
    layer0_outputs(6468) <= a;
    layer0_outputs(6469) <= not (a or b);
    layer0_outputs(6470) <= b;
    layer0_outputs(6471) <= not b or a;
    layer0_outputs(6472) <= not (a or b);
    layer0_outputs(6473) <= a and b;
    layer0_outputs(6474) <= not (a xor b);
    layer0_outputs(6475) <= a;
    layer0_outputs(6476) <= b and not a;
    layer0_outputs(6477) <= a or b;
    layer0_outputs(6478) <= not a;
    layer0_outputs(6479) <= not (a xor b);
    layer0_outputs(6480) <= a and not b;
    layer0_outputs(6481) <= not a;
    layer0_outputs(6482) <= '0';
    layer0_outputs(6483) <= a or b;
    layer0_outputs(6484) <= not (a or b);
    layer0_outputs(6485) <= not (a xor b);
    layer0_outputs(6486) <= a;
    layer0_outputs(6487) <= a and not b;
    layer0_outputs(6488) <= a and not b;
    layer0_outputs(6489) <= a;
    layer0_outputs(6490) <= b and not a;
    layer0_outputs(6491) <= not b;
    layer0_outputs(6492) <= not b or a;
    layer0_outputs(6493) <= not (a xor b);
    layer0_outputs(6494) <= not (a xor b);
    layer0_outputs(6495) <= not b or a;
    layer0_outputs(6496) <= not a or b;
    layer0_outputs(6497) <= not b or a;
    layer0_outputs(6498) <= not b;
    layer0_outputs(6499) <= not (a or b);
    layer0_outputs(6500) <= a and b;
    layer0_outputs(6501) <= a;
    layer0_outputs(6502) <= a;
    layer0_outputs(6503) <= not (a and b);
    layer0_outputs(6504) <= not a;
    layer0_outputs(6505) <= not (a or b);
    layer0_outputs(6506) <= not b or a;
    layer0_outputs(6507) <= '0';
    layer0_outputs(6508) <= a or b;
    layer0_outputs(6509) <= not (a and b);
    layer0_outputs(6510) <= b;
    layer0_outputs(6511) <= a and b;
    layer0_outputs(6512) <= not a;
    layer0_outputs(6513) <= not (a or b);
    layer0_outputs(6514) <= b and not a;
    layer0_outputs(6515) <= not a;
    layer0_outputs(6516) <= a or b;
    layer0_outputs(6517) <= a or b;
    layer0_outputs(6518) <= not b;
    layer0_outputs(6519) <= a or b;
    layer0_outputs(6520) <= not (a or b);
    layer0_outputs(6521) <= a;
    layer0_outputs(6522) <= a xor b;
    layer0_outputs(6523) <= not a;
    layer0_outputs(6524) <= b;
    layer0_outputs(6525) <= b;
    layer0_outputs(6526) <= b and not a;
    layer0_outputs(6527) <= b;
    layer0_outputs(6528) <= not b or a;
    layer0_outputs(6529) <= a;
    layer0_outputs(6530) <= not (a and b);
    layer0_outputs(6531) <= not a or b;
    layer0_outputs(6532) <= not (a xor b);
    layer0_outputs(6533) <= a and not b;
    layer0_outputs(6534) <= not b;
    layer0_outputs(6535) <= a and not b;
    layer0_outputs(6536) <= not a;
    layer0_outputs(6537) <= b;
    layer0_outputs(6538) <= a or b;
    layer0_outputs(6539) <= a or b;
    layer0_outputs(6540) <= '0';
    layer0_outputs(6541) <= b;
    layer0_outputs(6542) <= b and not a;
    layer0_outputs(6543) <= not b or a;
    layer0_outputs(6544) <= b;
    layer0_outputs(6545) <= not (a xor b);
    layer0_outputs(6546) <= not b;
    layer0_outputs(6547) <= b;
    layer0_outputs(6548) <= not a;
    layer0_outputs(6549) <= a xor b;
    layer0_outputs(6550) <= not b or a;
    layer0_outputs(6551) <= a or b;
    layer0_outputs(6552) <= a and b;
    layer0_outputs(6553) <= not (a xor b);
    layer0_outputs(6554) <= not b;
    layer0_outputs(6555) <= not b;
    layer0_outputs(6556) <= not (a or b);
    layer0_outputs(6557) <= a and b;
    layer0_outputs(6558) <= '1';
    layer0_outputs(6559) <= not a;
    layer0_outputs(6560) <= a xor b;
    layer0_outputs(6561) <= a;
    layer0_outputs(6562) <= a and b;
    layer0_outputs(6563) <= not (a or b);
    layer0_outputs(6564) <= b;
    layer0_outputs(6565) <= not (a and b);
    layer0_outputs(6566) <= b;
    layer0_outputs(6567) <= a;
    layer0_outputs(6568) <= not b or a;
    layer0_outputs(6569) <= not b;
    layer0_outputs(6570) <= b and not a;
    layer0_outputs(6571) <= not (a or b);
    layer0_outputs(6572) <= not a or b;
    layer0_outputs(6573) <= not a;
    layer0_outputs(6574) <= a;
    layer0_outputs(6575) <= a or b;
    layer0_outputs(6576) <= a and not b;
    layer0_outputs(6577) <= not b;
    layer0_outputs(6578) <= a and not b;
    layer0_outputs(6579) <= b;
    layer0_outputs(6580) <= a or b;
    layer0_outputs(6581) <= b and not a;
    layer0_outputs(6582) <= not b;
    layer0_outputs(6583) <= a xor b;
    layer0_outputs(6584) <= a and b;
    layer0_outputs(6585) <= a xor b;
    layer0_outputs(6586) <= not b;
    layer0_outputs(6587) <= '1';
    layer0_outputs(6588) <= not (a xor b);
    layer0_outputs(6589) <= '0';
    layer0_outputs(6590) <= '1';
    layer0_outputs(6591) <= '0';
    layer0_outputs(6592) <= not b or a;
    layer0_outputs(6593) <= b and not a;
    layer0_outputs(6594) <= not (a and b);
    layer0_outputs(6595) <= not b;
    layer0_outputs(6596) <= a;
    layer0_outputs(6597) <= not b or a;
    layer0_outputs(6598) <= a and not b;
    layer0_outputs(6599) <= a or b;
    layer0_outputs(6600) <= a or b;
    layer0_outputs(6601) <= b;
    layer0_outputs(6602) <= not b or a;
    layer0_outputs(6603) <= a;
    layer0_outputs(6604) <= a xor b;
    layer0_outputs(6605) <= a;
    layer0_outputs(6606) <= a;
    layer0_outputs(6607) <= not b or a;
    layer0_outputs(6608) <= not (a xor b);
    layer0_outputs(6609) <= not a or b;
    layer0_outputs(6610) <= b and not a;
    layer0_outputs(6611) <= '0';
    layer0_outputs(6612) <= a and b;
    layer0_outputs(6613) <= a xor b;
    layer0_outputs(6614) <= not a or b;
    layer0_outputs(6615) <= a and not b;
    layer0_outputs(6616) <= a and b;
    layer0_outputs(6617) <= not (a xor b);
    layer0_outputs(6618) <= not (a xor b);
    layer0_outputs(6619) <= not b;
    layer0_outputs(6620) <= not a or b;
    layer0_outputs(6621) <= not a;
    layer0_outputs(6622) <= b and not a;
    layer0_outputs(6623) <= b and not a;
    layer0_outputs(6624) <= '0';
    layer0_outputs(6625) <= a or b;
    layer0_outputs(6626) <= '0';
    layer0_outputs(6627) <= not a or b;
    layer0_outputs(6628) <= not b or a;
    layer0_outputs(6629) <= a and not b;
    layer0_outputs(6630) <= not b;
    layer0_outputs(6631) <= b and not a;
    layer0_outputs(6632) <= not a or b;
    layer0_outputs(6633) <= a or b;
    layer0_outputs(6634) <= a and not b;
    layer0_outputs(6635) <= a and not b;
    layer0_outputs(6636) <= b and not a;
    layer0_outputs(6637) <= not a;
    layer0_outputs(6638) <= a and b;
    layer0_outputs(6639) <= not (a or b);
    layer0_outputs(6640) <= not (a and b);
    layer0_outputs(6641) <= not a;
    layer0_outputs(6642) <= not b;
    layer0_outputs(6643) <= a and b;
    layer0_outputs(6644) <= not (a xor b);
    layer0_outputs(6645) <= not (a and b);
    layer0_outputs(6646) <= not b or a;
    layer0_outputs(6647) <= b and not a;
    layer0_outputs(6648) <= not b;
    layer0_outputs(6649) <= not a;
    layer0_outputs(6650) <= a and b;
    layer0_outputs(6651) <= b;
    layer0_outputs(6652) <= a xor b;
    layer0_outputs(6653) <= not b;
    layer0_outputs(6654) <= a xor b;
    layer0_outputs(6655) <= a xor b;
    layer0_outputs(6656) <= not (a or b);
    layer0_outputs(6657) <= a xor b;
    layer0_outputs(6658) <= not (a xor b);
    layer0_outputs(6659) <= a or b;
    layer0_outputs(6660) <= not a;
    layer0_outputs(6661) <= '0';
    layer0_outputs(6662) <= a or b;
    layer0_outputs(6663) <= b;
    layer0_outputs(6664) <= b;
    layer0_outputs(6665) <= not (a xor b);
    layer0_outputs(6666) <= not a or b;
    layer0_outputs(6667) <= not (a xor b);
    layer0_outputs(6668) <= b;
    layer0_outputs(6669) <= b;
    layer0_outputs(6670) <= a and b;
    layer0_outputs(6671) <= not b or a;
    layer0_outputs(6672) <= b and not a;
    layer0_outputs(6673) <= b;
    layer0_outputs(6674) <= a or b;
    layer0_outputs(6675) <= b and not a;
    layer0_outputs(6676) <= '1';
    layer0_outputs(6677) <= b;
    layer0_outputs(6678) <= not (a xor b);
    layer0_outputs(6679) <= not (a xor b);
    layer0_outputs(6680) <= a and not b;
    layer0_outputs(6681) <= not (a and b);
    layer0_outputs(6682) <= a xor b;
    layer0_outputs(6683) <= not (a xor b);
    layer0_outputs(6684) <= a xor b;
    layer0_outputs(6685) <= not a;
    layer0_outputs(6686) <= b;
    layer0_outputs(6687) <= not (a or b);
    layer0_outputs(6688) <= a or b;
    layer0_outputs(6689) <= not (a or b);
    layer0_outputs(6690) <= a and b;
    layer0_outputs(6691) <= not a or b;
    layer0_outputs(6692) <= not a;
    layer0_outputs(6693) <= a or b;
    layer0_outputs(6694) <= b and not a;
    layer0_outputs(6695) <= not (a xor b);
    layer0_outputs(6696) <= b and not a;
    layer0_outputs(6697) <= not b or a;
    layer0_outputs(6698) <= not b;
    layer0_outputs(6699) <= not b or a;
    layer0_outputs(6700) <= not (a or b);
    layer0_outputs(6701) <= not a;
    layer0_outputs(6702) <= b;
    layer0_outputs(6703) <= a and b;
    layer0_outputs(6704) <= a or b;
    layer0_outputs(6705) <= a and b;
    layer0_outputs(6706) <= a xor b;
    layer0_outputs(6707) <= not (a or b);
    layer0_outputs(6708) <= not (a or b);
    layer0_outputs(6709) <= b;
    layer0_outputs(6710) <= b;
    layer0_outputs(6711) <= '0';
    layer0_outputs(6712) <= not a or b;
    layer0_outputs(6713) <= not a or b;
    layer0_outputs(6714) <= b;
    layer0_outputs(6715) <= a and b;
    layer0_outputs(6716) <= not b;
    layer0_outputs(6717) <= not b;
    layer0_outputs(6718) <= not (a xor b);
    layer0_outputs(6719) <= not b;
    layer0_outputs(6720) <= '1';
    layer0_outputs(6721) <= '0';
    layer0_outputs(6722) <= b and not a;
    layer0_outputs(6723) <= b;
    layer0_outputs(6724) <= a and not b;
    layer0_outputs(6725) <= not b or a;
    layer0_outputs(6726) <= not a;
    layer0_outputs(6727) <= b;
    layer0_outputs(6728) <= not b or a;
    layer0_outputs(6729) <= a xor b;
    layer0_outputs(6730) <= b;
    layer0_outputs(6731) <= a or b;
    layer0_outputs(6732) <= a;
    layer0_outputs(6733) <= a or b;
    layer0_outputs(6734) <= not (a and b);
    layer0_outputs(6735) <= a;
    layer0_outputs(6736) <= not (a or b);
    layer0_outputs(6737) <= a or b;
    layer0_outputs(6738) <= not (a xor b);
    layer0_outputs(6739) <= a;
    layer0_outputs(6740) <= a or b;
    layer0_outputs(6741) <= not a;
    layer0_outputs(6742) <= a xor b;
    layer0_outputs(6743) <= not a or b;
    layer0_outputs(6744) <= not (a or b);
    layer0_outputs(6745) <= '0';
    layer0_outputs(6746) <= not a;
    layer0_outputs(6747) <= not (a or b);
    layer0_outputs(6748) <= a or b;
    layer0_outputs(6749) <= a and b;
    layer0_outputs(6750) <= a and b;
    layer0_outputs(6751) <= '1';
    layer0_outputs(6752) <= '1';
    layer0_outputs(6753) <= not (a xor b);
    layer0_outputs(6754) <= a and b;
    layer0_outputs(6755) <= not a;
    layer0_outputs(6756) <= a or b;
    layer0_outputs(6757) <= a or b;
    layer0_outputs(6758) <= a or b;
    layer0_outputs(6759) <= not (a xor b);
    layer0_outputs(6760) <= a;
    layer0_outputs(6761) <= not (a or b);
    layer0_outputs(6762) <= b;
    layer0_outputs(6763) <= not a or b;
    layer0_outputs(6764) <= not b;
    layer0_outputs(6765) <= not (a or b);
    layer0_outputs(6766) <= not (a or b);
    layer0_outputs(6767) <= not a or b;
    layer0_outputs(6768) <= a or b;
    layer0_outputs(6769) <= b and not a;
    layer0_outputs(6770) <= not a;
    layer0_outputs(6771) <= '1';
    layer0_outputs(6772) <= not (a and b);
    layer0_outputs(6773) <= not (a and b);
    layer0_outputs(6774) <= not a;
    layer0_outputs(6775) <= b;
    layer0_outputs(6776) <= a and not b;
    layer0_outputs(6777) <= not (a and b);
    layer0_outputs(6778) <= a xor b;
    layer0_outputs(6779) <= '0';
    layer0_outputs(6780) <= '1';
    layer0_outputs(6781) <= b;
    layer0_outputs(6782) <= not a or b;
    layer0_outputs(6783) <= a;
    layer0_outputs(6784) <= a xor b;
    layer0_outputs(6785) <= a xor b;
    layer0_outputs(6786) <= not (a or b);
    layer0_outputs(6787) <= '1';
    layer0_outputs(6788) <= not a;
    layer0_outputs(6789) <= a and not b;
    layer0_outputs(6790) <= a and b;
    layer0_outputs(6791) <= a xor b;
    layer0_outputs(6792) <= a or b;
    layer0_outputs(6793) <= '0';
    layer0_outputs(6794) <= not (a xor b);
    layer0_outputs(6795) <= not (a xor b);
    layer0_outputs(6796) <= not a or b;
    layer0_outputs(6797) <= not a or b;
    layer0_outputs(6798) <= b;
    layer0_outputs(6799) <= a;
    layer0_outputs(6800) <= a;
    layer0_outputs(6801) <= '0';
    layer0_outputs(6802) <= not (a or b);
    layer0_outputs(6803) <= b;
    layer0_outputs(6804) <= not b;
    layer0_outputs(6805) <= b and not a;
    layer0_outputs(6806) <= b;
    layer0_outputs(6807) <= '0';
    layer0_outputs(6808) <= not a;
    layer0_outputs(6809) <= b and not a;
    layer0_outputs(6810) <= a;
    layer0_outputs(6811) <= not (a and b);
    layer0_outputs(6812) <= a xor b;
    layer0_outputs(6813) <= not b or a;
    layer0_outputs(6814) <= '0';
    layer0_outputs(6815) <= '1';
    layer0_outputs(6816) <= not a;
    layer0_outputs(6817) <= b and not a;
    layer0_outputs(6818) <= b;
    layer0_outputs(6819) <= b;
    layer0_outputs(6820) <= not b or a;
    layer0_outputs(6821) <= b;
    layer0_outputs(6822) <= a;
    layer0_outputs(6823) <= not a;
    layer0_outputs(6824) <= '0';
    layer0_outputs(6825) <= not a;
    layer0_outputs(6826) <= a;
    layer0_outputs(6827) <= b and not a;
    layer0_outputs(6828) <= not a or b;
    layer0_outputs(6829) <= not (a or b);
    layer0_outputs(6830) <= not (a and b);
    layer0_outputs(6831) <= not b or a;
    layer0_outputs(6832) <= not b;
    layer0_outputs(6833) <= '1';
    layer0_outputs(6834) <= a xor b;
    layer0_outputs(6835) <= a or b;
    layer0_outputs(6836) <= not b;
    layer0_outputs(6837) <= not (a and b);
    layer0_outputs(6838) <= not b;
    layer0_outputs(6839) <= b;
    layer0_outputs(6840) <= not b;
    layer0_outputs(6841) <= a and not b;
    layer0_outputs(6842) <= not a;
    layer0_outputs(6843) <= not (a or b);
    layer0_outputs(6844) <= a or b;
    layer0_outputs(6845) <= b;
    layer0_outputs(6846) <= a xor b;
    layer0_outputs(6847) <= a and b;
    layer0_outputs(6848) <= a;
    layer0_outputs(6849) <= not b or a;
    layer0_outputs(6850) <= '1';
    layer0_outputs(6851) <= '1';
    layer0_outputs(6852) <= not b;
    layer0_outputs(6853) <= not (a or b);
    layer0_outputs(6854) <= a xor b;
    layer0_outputs(6855) <= b;
    layer0_outputs(6856) <= b;
    layer0_outputs(6857) <= not (a xor b);
    layer0_outputs(6858) <= b;
    layer0_outputs(6859) <= a xor b;
    layer0_outputs(6860) <= not (a and b);
    layer0_outputs(6861) <= not a or b;
    layer0_outputs(6862) <= not (a and b);
    layer0_outputs(6863) <= not a or b;
    layer0_outputs(6864) <= not a;
    layer0_outputs(6865) <= a xor b;
    layer0_outputs(6866) <= not b;
    layer0_outputs(6867) <= '0';
    layer0_outputs(6868) <= not b;
    layer0_outputs(6869) <= not (a xor b);
    layer0_outputs(6870) <= a and not b;
    layer0_outputs(6871) <= not (a and b);
    layer0_outputs(6872) <= not a;
    layer0_outputs(6873) <= not b;
    layer0_outputs(6874) <= a;
    layer0_outputs(6875) <= a xor b;
    layer0_outputs(6876) <= a xor b;
    layer0_outputs(6877) <= a;
    layer0_outputs(6878) <= not (a xor b);
    layer0_outputs(6879) <= not (a xor b);
    layer0_outputs(6880) <= not a or b;
    layer0_outputs(6881) <= b and not a;
    layer0_outputs(6882) <= a or b;
    layer0_outputs(6883) <= a;
    layer0_outputs(6884) <= not b;
    layer0_outputs(6885) <= a and not b;
    layer0_outputs(6886) <= not b or a;
    layer0_outputs(6887) <= not a;
    layer0_outputs(6888) <= a and b;
    layer0_outputs(6889) <= not b or a;
    layer0_outputs(6890) <= b;
    layer0_outputs(6891) <= not a;
    layer0_outputs(6892) <= not b;
    layer0_outputs(6893) <= a or b;
    layer0_outputs(6894) <= a;
    layer0_outputs(6895) <= a and b;
    layer0_outputs(6896) <= a or b;
    layer0_outputs(6897) <= not b;
    layer0_outputs(6898) <= a or b;
    layer0_outputs(6899) <= a or b;
    layer0_outputs(6900) <= not (a or b);
    layer0_outputs(6901) <= not b or a;
    layer0_outputs(6902) <= a or b;
    layer0_outputs(6903) <= not b;
    layer0_outputs(6904) <= not a;
    layer0_outputs(6905) <= a;
    layer0_outputs(6906) <= not b or a;
    layer0_outputs(6907) <= a and not b;
    layer0_outputs(6908) <= not b or a;
    layer0_outputs(6909) <= a xor b;
    layer0_outputs(6910) <= a and b;
    layer0_outputs(6911) <= not (a xor b);
    layer0_outputs(6912) <= not b or a;
    layer0_outputs(6913) <= not b or a;
    layer0_outputs(6914) <= not (a and b);
    layer0_outputs(6915) <= a;
    layer0_outputs(6916) <= a and not b;
    layer0_outputs(6917) <= not a or b;
    layer0_outputs(6918) <= '0';
    layer0_outputs(6919) <= not a;
    layer0_outputs(6920) <= a;
    layer0_outputs(6921) <= b;
    layer0_outputs(6922) <= a or b;
    layer0_outputs(6923) <= b and not a;
    layer0_outputs(6924) <= a or b;
    layer0_outputs(6925) <= a or b;
    layer0_outputs(6926) <= not a or b;
    layer0_outputs(6927) <= '0';
    layer0_outputs(6928) <= a or b;
    layer0_outputs(6929) <= not a;
    layer0_outputs(6930) <= a;
    layer0_outputs(6931) <= a and b;
    layer0_outputs(6932) <= not (a xor b);
    layer0_outputs(6933) <= '0';
    layer0_outputs(6934) <= not a;
    layer0_outputs(6935) <= not b;
    layer0_outputs(6936) <= not a;
    layer0_outputs(6937) <= a xor b;
    layer0_outputs(6938) <= not b or a;
    layer0_outputs(6939) <= '1';
    layer0_outputs(6940) <= not (a or b);
    layer0_outputs(6941) <= a xor b;
    layer0_outputs(6942) <= '0';
    layer0_outputs(6943) <= not a or b;
    layer0_outputs(6944) <= not b;
    layer0_outputs(6945) <= not b or a;
    layer0_outputs(6946) <= a or b;
    layer0_outputs(6947) <= a and b;
    layer0_outputs(6948) <= not a;
    layer0_outputs(6949) <= not b or a;
    layer0_outputs(6950) <= not (a or b);
    layer0_outputs(6951) <= not b;
    layer0_outputs(6952) <= '0';
    layer0_outputs(6953) <= a and not b;
    layer0_outputs(6954) <= a xor b;
    layer0_outputs(6955) <= a and not b;
    layer0_outputs(6956) <= a or b;
    layer0_outputs(6957) <= '1';
    layer0_outputs(6958) <= not a or b;
    layer0_outputs(6959) <= not (a xor b);
    layer0_outputs(6960) <= b;
    layer0_outputs(6961) <= a or b;
    layer0_outputs(6962) <= a and b;
    layer0_outputs(6963) <= not b;
    layer0_outputs(6964) <= not b or a;
    layer0_outputs(6965) <= a or b;
    layer0_outputs(6966) <= a;
    layer0_outputs(6967) <= '0';
    layer0_outputs(6968) <= b and not a;
    layer0_outputs(6969) <= a xor b;
    layer0_outputs(6970) <= '1';
    layer0_outputs(6971) <= '0';
    layer0_outputs(6972) <= not b;
    layer0_outputs(6973) <= not a;
    layer0_outputs(6974) <= b and not a;
    layer0_outputs(6975) <= '1';
    layer0_outputs(6976) <= a or b;
    layer0_outputs(6977) <= not (a xor b);
    layer0_outputs(6978) <= a or b;
    layer0_outputs(6979) <= not b or a;
    layer0_outputs(6980) <= not (a xor b);
    layer0_outputs(6981) <= b;
    layer0_outputs(6982) <= b and not a;
    layer0_outputs(6983) <= a xor b;
    layer0_outputs(6984) <= '0';
    layer0_outputs(6985) <= not (a or b);
    layer0_outputs(6986) <= b;
    layer0_outputs(6987) <= not (a or b);
    layer0_outputs(6988) <= a and b;
    layer0_outputs(6989) <= a and not b;
    layer0_outputs(6990) <= not b or a;
    layer0_outputs(6991) <= not b or a;
    layer0_outputs(6992) <= b and not a;
    layer0_outputs(6993) <= a;
    layer0_outputs(6994) <= b;
    layer0_outputs(6995) <= '1';
    layer0_outputs(6996) <= not b or a;
    layer0_outputs(6997) <= b and not a;
    layer0_outputs(6998) <= a;
    layer0_outputs(6999) <= not (a xor b);
    layer0_outputs(7000) <= not (a and b);
    layer0_outputs(7001) <= not a;
    layer0_outputs(7002) <= not b or a;
    layer0_outputs(7003) <= not (a and b);
    layer0_outputs(7004) <= not a;
    layer0_outputs(7005) <= '1';
    layer0_outputs(7006) <= not b;
    layer0_outputs(7007) <= not b or a;
    layer0_outputs(7008) <= a xor b;
    layer0_outputs(7009) <= not a;
    layer0_outputs(7010) <= not a;
    layer0_outputs(7011) <= not (a or b);
    layer0_outputs(7012) <= a and b;
    layer0_outputs(7013) <= not (a or b);
    layer0_outputs(7014) <= not a or b;
    layer0_outputs(7015) <= a and not b;
    layer0_outputs(7016) <= not b;
    layer0_outputs(7017) <= b;
    layer0_outputs(7018) <= '1';
    layer0_outputs(7019) <= a and not b;
    layer0_outputs(7020) <= b and not a;
    layer0_outputs(7021) <= b and not a;
    layer0_outputs(7022) <= a and not b;
    layer0_outputs(7023) <= not a;
    layer0_outputs(7024) <= not (a xor b);
    layer0_outputs(7025) <= b and not a;
    layer0_outputs(7026) <= not (a and b);
    layer0_outputs(7027) <= a or b;
    layer0_outputs(7028) <= not (a or b);
    layer0_outputs(7029) <= b;
    layer0_outputs(7030) <= not a or b;
    layer0_outputs(7031) <= a and not b;
    layer0_outputs(7032) <= a xor b;
    layer0_outputs(7033) <= not b or a;
    layer0_outputs(7034) <= '1';
    layer0_outputs(7035) <= a and b;
    layer0_outputs(7036) <= not b;
    layer0_outputs(7037) <= not (a and b);
    layer0_outputs(7038) <= not (a or b);
    layer0_outputs(7039) <= not (a or b);
    layer0_outputs(7040) <= a and b;
    layer0_outputs(7041) <= not b;
    layer0_outputs(7042) <= '1';
    layer0_outputs(7043) <= b;
    layer0_outputs(7044) <= not b or a;
    layer0_outputs(7045) <= '1';
    layer0_outputs(7046) <= b;
    layer0_outputs(7047) <= not (a xor b);
    layer0_outputs(7048) <= not a or b;
    layer0_outputs(7049) <= '0';
    layer0_outputs(7050) <= '1';
    layer0_outputs(7051) <= b;
    layer0_outputs(7052) <= not a;
    layer0_outputs(7053) <= not (a and b);
    layer0_outputs(7054) <= b and not a;
    layer0_outputs(7055) <= '1';
    layer0_outputs(7056) <= not a or b;
    layer0_outputs(7057) <= not b;
    layer0_outputs(7058) <= '0';
    layer0_outputs(7059) <= a xor b;
    layer0_outputs(7060) <= b;
    layer0_outputs(7061) <= a and not b;
    layer0_outputs(7062) <= b;
    layer0_outputs(7063) <= not (a xor b);
    layer0_outputs(7064) <= not b or a;
    layer0_outputs(7065) <= a xor b;
    layer0_outputs(7066) <= '1';
    layer0_outputs(7067) <= not a;
    layer0_outputs(7068) <= b and not a;
    layer0_outputs(7069) <= not (a xor b);
    layer0_outputs(7070) <= a or b;
    layer0_outputs(7071) <= '0';
    layer0_outputs(7072) <= a and b;
    layer0_outputs(7073) <= not b;
    layer0_outputs(7074) <= not (a and b);
    layer0_outputs(7075) <= not (a and b);
    layer0_outputs(7076) <= a xor b;
    layer0_outputs(7077) <= not (a and b);
    layer0_outputs(7078) <= b and not a;
    layer0_outputs(7079) <= not (a or b);
    layer0_outputs(7080) <= b;
    layer0_outputs(7081) <= a;
    layer0_outputs(7082) <= not b or a;
    layer0_outputs(7083) <= a;
    layer0_outputs(7084) <= not b;
    layer0_outputs(7085) <= a xor b;
    layer0_outputs(7086) <= a xor b;
    layer0_outputs(7087) <= a;
    layer0_outputs(7088) <= not a or b;
    layer0_outputs(7089) <= '1';
    layer0_outputs(7090) <= not (a or b);
    layer0_outputs(7091) <= b;
    layer0_outputs(7092) <= not b or a;
    layer0_outputs(7093) <= a xor b;
    layer0_outputs(7094) <= not b;
    layer0_outputs(7095) <= a xor b;
    layer0_outputs(7096) <= not a;
    layer0_outputs(7097) <= not (a xor b);
    layer0_outputs(7098) <= not b;
    layer0_outputs(7099) <= not b;
    layer0_outputs(7100) <= not b;
    layer0_outputs(7101) <= not b;
    layer0_outputs(7102) <= not b;
    layer0_outputs(7103) <= not b or a;
    layer0_outputs(7104) <= not (a or b);
    layer0_outputs(7105) <= a;
    layer0_outputs(7106) <= not a or b;
    layer0_outputs(7107) <= not b;
    layer0_outputs(7108) <= a or b;
    layer0_outputs(7109) <= a and b;
    layer0_outputs(7110) <= a or b;
    layer0_outputs(7111) <= a and not b;
    layer0_outputs(7112) <= a and not b;
    layer0_outputs(7113) <= a or b;
    layer0_outputs(7114) <= not (a xor b);
    layer0_outputs(7115) <= a or b;
    layer0_outputs(7116) <= a and not b;
    layer0_outputs(7117) <= not a or b;
    layer0_outputs(7118) <= not b or a;
    layer0_outputs(7119) <= a and b;
    layer0_outputs(7120) <= a xor b;
    layer0_outputs(7121) <= '0';
    layer0_outputs(7122) <= a and not b;
    layer0_outputs(7123) <= not a;
    layer0_outputs(7124) <= not (a xor b);
    layer0_outputs(7125) <= a and b;
    layer0_outputs(7126) <= a and not b;
    layer0_outputs(7127) <= not b;
    layer0_outputs(7128) <= a xor b;
    layer0_outputs(7129) <= not b or a;
    layer0_outputs(7130) <= a and not b;
    layer0_outputs(7131) <= '1';
    layer0_outputs(7132) <= b;
    layer0_outputs(7133) <= not (a or b);
    layer0_outputs(7134) <= not b;
    layer0_outputs(7135) <= not a;
    layer0_outputs(7136) <= a and b;
    layer0_outputs(7137) <= not (a xor b);
    layer0_outputs(7138) <= not (a and b);
    layer0_outputs(7139) <= a xor b;
    layer0_outputs(7140) <= not b;
    layer0_outputs(7141) <= not b or a;
    layer0_outputs(7142) <= not (a xor b);
    layer0_outputs(7143) <= a and b;
    layer0_outputs(7144) <= b;
    layer0_outputs(7145) <= not b;
    layer0_outputs(7146) <= not a;
    layer0_outputs(7147) <= not a;
    layer0_outputs(7148) <= not b;
    layer0_outputs(7149) <= a;
    layer0_outputs(7150) <= not b or a;
    layer0_outputs(7151) <= not (a and b);
    layer0_outputs(7152) <= '1';
    layer0_outputs(7153) <= a;
    layer0_outputs(7154) <= b and not a;
    layer0_outputs(7155) <= not b;
    layer0_outputs(7156) <= '1';
    layer0_outputs(7157) <= '0';
    layer0_outputs(7158) <= a;
    layer0_outputs(7159) <= a and b;
    layer0_outputs(7160) <= not b or a;
    layer0_outputs(7161) <= not b;
    layer0_outputs(7162) <= not (a xor b);
    layer0_outputs(7163) <= not (a or b);
    layer0_outputs(7164) <= not a or b;
    layer0_outputs(7165) <= not b;
    layer0_outputs(7166) <= not b or a;
    layer0_outputs(7167) <= a xor b;
    layer0_outputs(7168) <= not a or b;
    layer0_outputs(7169) <= a and b;
    layer0_outputs(7170) <= b;
    layer0_outputs(7171) <= b and not a;
    layer0_outputs(7172) <= a;
    layer0_outputs(7173) <= not b;
    layer0_outputs(7174) <= not b or a;
    layer0_outputs(7175) <= a and b;
    layer0_outputs(7176) <= a;
    layer0_outputs(7177) <= not (a or b);
    layer0_outputs(7178) <= not (a xor b);
    layer0_outputs(7179) <= not b or a;
    layer0_outputs(7180) <= not a or b;
    layer0_outputs(7181) <= '1';
    layer0_outputs(7182) <= b and not a;
    layer0_outputs(7183) <= not (a xor b);
    layer0_outputs(7184) <= not b;
    layer0_outputs(7185) <= not a;
    layer0_outputs(7186) <= not (a and b);
    layer0_outputs(7187) <= not a;
    layer0_outputs(7188) <= a xor b;
    layer0_outputs(7189) <= b and not a;
    layer0_outputs(7190) <= not a or b;
    layer0_outputs(7191) <= a;
    layer0_outputs(7192) <= b;
    layer0_outputs(7193) <= not a or b;
    layer0_outputs(7194) <= not (a or b);
    layer0_outputs(7195) <= not a;
    layer0_outputs(7196) <= not (a xor b);
    layer0_outputs(7197) <= not b;
    layer0_outputs(7198) <= a xor b;
    layer0_outputs(7199) <= not a;
    layer0_outputs(7200) <= '1';
    layer0_outputs(7201) <= not b;
    layer0_outputs(7202) <= a;
    layer0_outputs(7203) <= '1';
    layer0_outputs(7204) <= a and b;
    layer0_outputs(7205) <= '0';
    layer0_outputs(7206) <= b and not a;
    layer0_outputs(7207) <= a and not b;
    layer0_outputs(7208) <= a;
    layer0_outputs(7209) <= not a;
    layer0_outputs(7210) <= b;
    layer0_outputs(7211) <= a and not b;
    layer0_outputs(7212) <= a;
    layer0_outputs(7213) <= not a;
    layer0_outputs(7214) <= '1';
    layer0_outputs(7215) <= not (a or b);
    layer0_outputs(7216) <= not (a or b);
    layer0_outputs(7217) <= not a or b;
    layer0_outputs(7218) <= '1';
    layer0_outputs(7219) <= a and b;
    layer0_outputs(7220) <= not (a xor b);
    layer0_outputs(7221) <= b;
    layer0_outputs(7222) <= not a;
    layer0_outputs(7223) <= '1';
    layer0_outputs(7224) <= a or b;
    layer0_outputs(7225) <= not (a and b);
    layer0_outputs(7226) <= not (a and b);
    layer0_outputs(7227) <= a or b;
    layer0_outputs(7228) <= a xor b;
    layer0_outputs(7229) <= not (a or b);
    layer0_outputs(7230) <= a;
    layer0_outputs(7231) <= '1';
    layer0_outputs(7232) <= not a;
    layer0_outputs(7233) <= not (a xor b);
    layer0_outputs(7234) <= b and not a;
    layer0_outputs(7235) <= not a or b;
    layer0_outputs(7236) <= a and not b;
    layer0_outputs(7237) <= not (a xor b);
    layer0_outputs(7238) <= not (a and b);
    layer0_outputs(7239) <= not (a and b);
    layer0_outputs(7240) <= not b;
    layer0_outputs(7241) <= '1';
    layer0_outputs(7242) <= not (a and b);
    layer0_outputs(7243) <= a or b;
    layer0_outputs(7244) <= not a;
    layer0_outputs(7245) <= b and not a;
    layer0_outputs(7246) <= '1';
    layer0_outputs(7247) <= not (a or b);
    layer0_outputs(7248) <= b;
    layer0_outputs(7249) <= b and not a;
    layer0_outputs(7250) <= not (a xor b);
    layer0_outputs(7251) <= '1';
    layer0_outputs(7252) <= b and not a;
    layer0_outputs(7253) <= '1';
    layer0_outputs(7254) <= not (a or b);
    layer0_outputs(7255) <= a;
    layer0_outputs(7256) <= not b;
    layer0_outputs(7257) <= not b;
    layer0_outputs(7258) <= not (a or b);
    layer0_outputs(7259) <= not b;
    layer0_outputs(7260) <= not (a or b);
    layer0_outputs(7261) <= not (a or b);
    layer0_outputs(7262) <= a;
    layer0_outputs(7263) <= not a or b;
    layer0_outputs(7264) <= not (a xor b);
    layer0_outputs(7265) <= not (a or b);
    layer0_outputs(7266) <= not a;
    layer0_outputs(7267) <= not (a or b);
    layer0_outputs(7268) <= not (a or b);
    layer0_outputs(7269) <= a and b;
    layer0_outputs(7270) <= a and b;
    layer0_outputs(7271) <= not b;
    layer0_outputs(7272) <= not a or b;
    layer0_outputs(7273) <= not a;
    layer0_outputs(7274) <= b;
    layer0_outputs(7275) <= not b or a;
    layer0_outputs(7276) <= not (a or b);
    layer0_outputs(7277) <= not a;
    layer0_outputs(7278) <= a and not b;
    layer0_outputs(7279) <= not (a or b);
    layer0_outputs(7280) <= not b;
    layer0_outputs(7281) <= '0';
    layer0_outputs(7282) <= a and not b;
    layer0_outputs(7283) <= not a or b;
    layer0_outputs(7284) <= '0';
    layer0_outputs(7285) <= a;
    layer0_outputs(7286) <= a or b;
    layer0_outputs(7287) <= b;
    layer0_outputs(7288) <= a xor b;
    layer0_outputs(7289) <= b and not a;
    layer0_outputs(7290) <= not b or a;
    layer0_outputs(7291) <= a and b;
    layer0_outputs(7292) <= b and not a;
    layer0_outputs(7293) <= not (a and b);
    layer0_outputs(7294) <= not (a or b);
    layer0_outputs(7295) <= a and b;
    layer0_outputs(7296) <= not a;
    layer0_outputs(7297) <= '0';
    layer0_outputs(7298) <= not (a and b);
    layer0_outputs(7299) <= a and not b;
    layer0_outputs(7300) <= not b;
    layer0_outputs(7301) <= b;
    layer0_outputs(7302) <= a xor b;
    layer0_outputs(7303) <= a;
    layer0_outputs(7304) <= not a or b;
    layer0_outputs(7305) <= not (a or b);
    layer0_outputs(7306) <= not (a and b);
    layer0_outputs(7307) <= not (a xor b);
    layer0_outputs(7308) <= a;
    layer0_outputs(7309) <= not (a or b);
    layer0_outputs(7310) <= a or b;
    layer0_outputs(7311) <= not a;
    layer0_outputs(7312) <= a and not b;
    layer0_outputs(7313) <= not (a xor b);
    layer0_outputs(7314) <= b;
    layer0_outputs(7315) <= not a;
    layer0_outputs(7316) <= b;
    layer0_outputs(7317) <= not a;
    layer0_outputs(7318) <= a xor b;
    layer0_outputs(7319) <= a;
    layer0_outputs(7320) <= not (a xor b);
    layer0_outputs(7321) <= '1';
    layer0_outputs(7322) <= b and not a;
    layer0_outputs(7323) <= a or b;
    layer0_outputs(7324) <= not a;
    layer0_outputs(7325) <= a and b;
    layer0_outputs(7326) <= b;
    layer0_outputs(7327) <= '1';
    layer0_outputs(7328) <= not a or b;
    layer0_outputs(7329) <= a or b;
    layer0_outputs(7330) <= a or b;
    layer0_outputs(7331) <= not a;
    layer0_outputs(7332) <= not (a and b);
    layer0_outputs(7333) <= not (a and b);
    layer0_outputs(7334) <= not a or b;
    layer0_outputs(7335) <= a or b;
    layer0_outputs(7336) <= a or b;
    layer0_outputs(7337) <= a and not b;
    layer0_outputs(7338) <= b;
    layer0_outputs(7339) <= a and not b;
    layer0_outputs(7340) <= a or b;
    layer0_outputs(7341) <= not (a and b);
    layer0_outputs(7342) <= not a;
    layer0_outputs(7343) <= not a or b;
    layer0_outputs(7344) <= not b;
    layer0_outputs(7345) <= not b or a;
    layer0_outputs(7346) <= a;
    layer0_outputs(7347) <= not a;
    layer0_outputs(7348) <= '1';
    layer0_outputs(7349) <= b;
    layer0_outputs(7350) <= not (a or b);
    layer0_outputs(7351) <= a;
    layer0_outputs(7352) <= not b or a;
    layer0_outputs(7353) <= not b;
    layer0_outputs(7354) <= not (a and b);
    layer0_outputs(7355) <= a;
    layer0_outputs(7356) <= not (a xor b);
    layer0_outputs(7357) <= not b;
    layer0_outputs(7358) <= not a or b;
    layer0_outputs(7359) <= a or b;
    layer0_outputs(7360) <= '0';
    layer0_outputs(7361) <= b;
    layer0_outputs(7362) <= not a or b;
    layer0_outputs(7363) <= not b;
    layer0_outputs(7364) <= a and b;
    layer0_outputs(7365) <= a or b;
    layer0_outputs(7366) <= a;
    layer0_outputs(7367) <= not a or b;
    layer0_outputs(7368) <= b;
    layer0_outputs(7369) <= not (a or b);
    layer0_outputs(7370) <= not (a and b);
    layer0_outputs(7371) <= not a;
    layer0_outputs(7372) <= not (a or b);
    layer0_outputs(7373) <= not b;
    layer0_outputs(7374) <= not a;
    layer0_outputs(7375) <= not b;
    layer0_outputs(7376) <= not (a or b);
    layer0_outputs(7377) <= not b;
    layer0_outputs(7378) <= '1';
    layer0_outputs(7379) <= a;
    layer0_outputs(7380) <= b and not a;
    layer0_outputs(7381) <= not (a and b);
    layer0_outputs(7382) <= not b or a;
    layer0_outputs(7383) <= b and not a;
    layer0_outputs(7384) <= a and not b;
    layer0_outputs(7385) <= a and b;
    layer0_outputs(7386) <= b and not a;
    layer0_outputs(7387) <= a and b;
    layer0_outputs(7388) <= not a or b;
    layer0_outputs(7389) <= a;
    layer0_outputs(7390) <= a and b;
    layer0_outputs(7391) <= a;
    layer0_outputs(7392) <= b;
    layer0_outputs(7393) <= not b;
    layer0_outputs(7394) <= b and not a;
    layer0_outputs(7395) <= a or b;
    layer0_outputs(7396) <= '0';
    layer0_outputs(7397) <= not (a and b);
    layer0_outputs(7398) <= not (a or b);
    layer0_outputs(7399) <= not (a and b);
    layer0_outputs(7400) <= a xor b;
    layer0_outputs(7401) <= a;
    layer0_outputs(7402) <= a and b;
    layer0_outputs(7403) <= a;
    layer0_outputs(7404) <= not b or a;
    layer0_outputs(7405) <= not (a or b);
    layer0_outputs(7406) <= not (a and b);
    layer0_outputs(7407) <= '0';
    layer0_outputs(7408) <= not (a or b);
    layer0_outputs(7409) <= not b or a;
    layer0_outputs(7410) <= a or b;
    layer0_outputs(7411) <= a and b;
    layer0_outputs(7412) <= not (a xor b);
    layer0_outputs(7413) <= a and not b;
    layer0_outputs(7414) <= a and b;
    layer0_outputs(7415) <= not (a xor b);
    layer0_outputs(7416) <= '1';
    layer0_outputs(7417) <= b and not a;
    layer0_outputs(7418) <= not (a or b);
    layer0_outputs(7419) <= a;
    layer0_outputs(7420) <= not b;
    layer0_outputs(7421) <= b and not a;
    layer0_outputs(7422) <= a or b;
    layer0_outputs(7423) <= not a;
    layer0_outputs(7424) <= not b or a;
    layer0_outputs(7425) <= a;
    layer0_outputs(7426) <= b;
    layer0_outputs(7427) <= not a;
    layer0_outputs(7428) <= a;
    layer0_outputs(7429) <= b and not a;
    layer0_outputs(7430) <= not a or b;
    layer0_outputs(7431) <= not (a or b);
    layer0_outputs(7432) <= not a or b;
    layer0_outputs(7433) <= not (a xor b);
    layer0_outputs(7434) <= a;
    layer0_outputs(7435) <= a and b;
    layer0_outputs(7436) <= a or b;
    layer0_outputs(7437) <= a and not b;
    layer0_outputs(7438) <= not b;
    layer0_outputs(7439) <= a and not b;
    layer0_outputs(7440) <= a xor b;
    layer0_outputs(7441) <= a and not b;
    layer0_outputs(7442) <= not b;
    layer0_outputs(7443) <= not a or b;
    layer0_outputs(7444) <= not a;
    layer0_outputs(7445) <= not (a xor b);
    layer0_outputs(7446) <= not (a or b);
    layer0_outputs(7447) <= '1';
    layer0_outputs(7448) <= not b or a;
    layer0_outputs(7449) <= not (a and b);
    layer0_outputs(7450) <= b and not a;
    layer0_outputs(7451) <= not (a and b);
    layer0_outputs(7452) <= a or b;
    layer0_outputs(7453) <= a xor b;
    layer0_outputs(7454) <= a xor b;
    layer0_outputs(7455) <= not (a or b);
    layer0_outputs(7456) <= a or b;
    layer0_outputs(7457) <= a or b;
    layer0_outputs(7458) <= not (a and b);
    layer0_outputs(7459) <= a and b;
    layer0_outputs(7460) <= a;
    layer0_outputs(7461) <= a;
    layer0_outputs(7462) <= not (a and b);
    layer0_outputs(7463) <= not (a or b);
    layer0_outputs(7464) <= not b or a;
    layer0_outputs(7465) <= b and not a;
    layer0_outputs(7466) <= a or b;
    layer0_outputs(7467) <= a or b;
    layer0_outputs(7468) <= a and not b;
    layer0_outputs(7469) <= b and not a;
    layer0_outputs(7470) <= not (a or b);
    layer0_outputs(7471) <= a and b;
    layer0_outputs(7472) <= a or b;
    layer0_outputs(7473) <= not b or a;
    layer0_outputs(7474) <= not (a or b);
    layer0_outputs(7475) <= b;
    layer0_outputs(7476) <= not a;
    layer0_outputs(7477) <= a or b;
    layer0_outputs(7478) <= a or b;
    layer0_outputs(7479) <= not (a or b);
    layer0_outputs(7480) <= a and b;
    layer0_outputs(7481) <= not a;
    layer0_outputs(7482) <= a and not b;
    layer0_outputs(7483) <= a or b;
    layer0_outputs(7484) <= not (a xor b);
    layer0_outputs(7485) <= not a;
    layer0_outputs(7486) <= not (a xor b);
    layer0_outputs(7487) <= not (a or b);
    layer0_outputs(7488) <= '0';
    layer0_outputs(7489) <= b and not a;
    layer0_outputs(7490) <= a;
    layer0_outputs(7491) <= a;
    layer0_outputs(7492) <= not a;
    layer0_outputs(7493) <= a and not b;
    layer0_outputs(7494) <= not b;
    layer0_outputs(7495) <= not b or a;
    layer0_outputs(7496) <= a and b;
    layer0_outputs(7497) <= not a;
    layer0_outputs(7498) <= a xor b;
    layer0_outputs(7499) <= '0';
    layer0_outputs(7500) <= not (a and b);
    layer0_outputs(7501) <= not a or b;
    layer0_outputs(7502) <= '0';
    layer0_outputs(7503) <= '1';
    layer0_outputs(7504) <= not a;
    layer0_outputs(7505) <= a or b;
    layer0_outputs(7506) <= a xor b;
    layer0_outputs(7507) <= a xor b;
    layer0_outputs(7508) <= '0';
    layer0_outputs(7509) <= not (a or b);
    layer0_outputs(7510) <= not b;
    layer0_outputs(7511) <= b and not a;
    layer0_outputs(7512) <= b and not a;
    layer0_outputs(7513) <= a;
    layer0_outputs(7514) <= b;
    layer0_outputs(7515) <= '1';
    layer0_outputs(7516) <= not a or b;
    layer0_outputs(7517) <= b;
    layer0_outputs(7518) <= a and not b;
    layer0_outputs(7519) <= not a;
    layer0_outputs(7520) <= not b or a;
    layer0_outputs(7521) <= '1';
    layer0_outputs(7522) <= b;
    layer0_outputs(7523) <= b and not a;
    layer0_outputs(7524) <= a and not b;
    layer0_outputs(7525) <= a and b;
    layer0_outputs(7526) <= not (a xor b);
    layer0_outputs(7527) <= a and not b;
    layer0_outputs(7528) <= '1';
    layer0_outputs(7529) <= not (a or b);
    layer0_outputs(7530) <= a or b;
    layer0_outputs(7531) <= b;
    layer0_outputs(7532) <= a;
    layer0_outputs(7533) <= not (a or b);
    layer0_outputs(7534) <= b;
    layer0_outputs(7535) <= a or b;
    layer0_outputs(7536) <= not (a or b);
    layer0_outputs(7537) <= '1';
    layer0_outputs(7538) <= a xor b;
    layer0_outputs(7539) <= not a;
    layer0_outputs(7540) <= '1';
    layer0_outputs(7541) <= a and not b;
    layer0_outputs(7542) <= '0';
    layer0_outputs(7543) <= not a;
    layer0_outputs(7544) <= a;
    layer0_outputs(7545) <= not (a and b);
    layer0_outputs(7546) <= a;
    layer0_outputs(7547) <= not a or b;
    layer0_outputs(7548) <= not a;
    layer0_outputs(7549) <= not a or b;
    layer0_outputs(7550) <= not b or a;
    layer0_outputs(7551) <= not b;
    layer0_outputs(7552) <= not b;
    layer0_outputs(7553) <= not b;
    layer0_outputs(7554) <= a or b;
    layer0_outputs(7555) <= not a or b;
    layer0_outputs(7556) <= not b or a;
    layer0_outputs(7557) <= not b;
    layer0_outputs(7558) <= a xor b;
    layer0_outputs(7559) <= b and not a;
    layer0_outputs(7560) <= a or b;
    layer0_outputs(7561) <= b;
    layer0_outputs(7562) <= b;
    layer0_outputs(7563) <= '0';
    layer0_outputs(7564) <= not (a and b);
    layer0_outputs(7565) <= a and b;
    layer0_outputs(7566) <= b;
    layer0_outputs(7567) <= a or b;
    layer0_outputs(7568) <= '1';
    layer0_outputs(7569) <= not (a xor b);
    layer0_outputs(7570) <= a xor b;
    layer0_outputs(7571) <= a or b;
    layer0_outputs(7572) <= a xor b;
    layer0_outputs(7573) <= '1';
    layer0_outputs(7574) <= not b;
    layer0_outputs(7575) <= not (a or b);
    layer0_outputs(7576) <= a or b;
    layer0_outputs(7577) <= a or b;
    layer0_outputs(7578) <= a or b;
    layer0_outputs(7579) <= not (a or b);
    layer0_outputs(7580) <= not (a or b);
    layer0_outputs(7581) <= a and b;
    layer0_outputs(7582) <= a and not b;
    layer0_outputs(7583) <= a and not b;
    layer0_outputs(7584) <= not b or a;
    layer0_outputs(7585) <= a or b;
    layer0_outputs(7586) <= not b;
    layer0_outputs(7587) <= b and not a;
    layer0_outputs(7588) <= a and not b;
    layer0_outputs(7589) <= not b;
    layer0_outputs(7590) <= b;
    layer0_outputs(7591) <= a and b;
    layer0_outputs(7592) <= not b or a;
    layer0_outputs(7593) <= '0';
    layer0_outputs(7594) <= b;
    layer0_outputs(7595) <= '1';
    layer0_outputs(7596) <= not b or a;
    layer0_outputs(7597) <= not (a or b);
    layer0_outputs(7598) <= b and not a;
    layer0_outputs(7599) <= not b or a;
    layer0_outputs(7600) <= a and b;
    layer0_outputs(7601) <= not a;
    layer0_outputs(7602) <= a;
    layer0_outputs(7603) <= not (a or b);
    layer0_outputs(7604) <= not (a xor b);
    layer0_outputs(7605) <= not (a or b);
    layer0_outputs(7606) <= a xor b;
    layer0_outputs(7607) <= a xor b;
    layer0_outputs(7608) <= a and not b;
    layer0_outputs(7609) <= a;
    layer0_outputs(7610) <= a or b;
    layer0_outputs(7611) <= a xor b;
    layer0_outputs(7612) <= a or b;
    layer0_outputs(7613) <= a and not b;
    layer0_outputs(7614) <= a or b;
    layer0_outputs(7615) <= not (a and b);
    layer0_outputs(7616) <= not a or b;
    layer0_outputs(7617) <= a xor b;
    layer0_outputs(7618) <= '0';
    layer0_outputs(7619) <= not b or a;
    layer0_outputs(7620) <= b and not a;
    layer0_outputs(7621) <= not (a and b);
    layer0_outputs(7622) <= not (a and b);
    layer0_outputs(7623) <= a and not b;
    layer0_outputs(7624) <= not a or b;
    layer0_outputs(7625) <= not b or a;
    layer0_outputs(7626) <= not (a or b);
    layer0_outputs(7627) <= not a or b;
    layer0_outputs(7628) <= not b;
    layer0_outputs(7629) <= b and not a;
    layer0_outputs(7630) <= a;
    layer0_outputs(7631) <= b and not a;
    layer0_outputs(7632) <= not a;
    layer0_outputs(7633) <= a;
    layer0_outputs(7634) <= a and not b;
    layer0_outputs(7635) <= not b;
    layer0_outputs(7636) <= not a or b;
    layer0_outputs(7637) <= '1';
    layer0_outputs(7638) <= not (a or b);
    layer0_outputs(7639) <= a or b;
    layer0_outputs(7640) <= '0';
    layer0_outputs(7641) <= not a or b;
    layer0_outputs(7642) <= not b or a;
    layer0_outputs(7643) <= b;
    layer0_outputs(7644) <= a xor b;
    layer0_outputs(7645) <= a;
    layer0_outputs(7646) <= not a or b;
    layer0_outputs(7647) <= a or b;
    layer0_outputs(7648) <= a xor b;
    layer0_outputs(7649) <= not b or a;
    layer0_outputs(7650) <= '0';
    layer0_outputs(7651) <= a and not b;
    layer0_outputs(7652) <= a or b;
    layer0_outputs(7653) <= not (a or b);
    layer0_outputs(7654) <= a and not b;
    layer0_outputs(7655) <= not a or b;
    layer0_outputs(7656) <= not (a and b);
    layer0_outputs(7657) <= not (a or b);
    layer0_outputs(7658) <= not a;
    layer0_outputs(7659) <= a;
    layer0_outputs(7660) <= not b or a;
    layer0_outputs(7661) <= a or b;
    layer0_outputs(7662) <= a or b;
    layer0_outputs(7663) <= a or b;
    layer0_outputs(7664) <= '0';
    layer0_outputs(7665) <= a xor b;
    layer0_outputs(7666) <= a or b;
    layer0_outputs(7667) <= '1';
    layer0_outputs(7668) <= b;
    layer0_outputs(7669) <= not a;
    layer0_outputs(7670) <= b and not a;
    layer0_outputs(7671) <= not (a xor b);
    layer0_outputs(7672) <= not b;
    layer0_outputs(7673) <= b and not a;
    layer0_outputs(7674) <= a xor b;
    layer0_outputs(7675) <= not a or b;
    layer0_outputs(7676) <= not (a xor b);
    layer0_outputs(7677) <= b;
    layer0_outputs(7678) <= a;
    layer0_outputs(7679) <= a or b;
    layer0_outputs(7680) <= not b;
    layer0_outputs(7681) <= not (a xor b);
    layer0_outputs(7682) <= not a or b;
    layer0_outputs(7683) <= a;
    layer0_outputs(7684) <= '1';
    layer0_outputs(7685) <= not (a or b);
    layer0_outputs(7686) <= b;
    layer0_outputs(7687) <= '0';
    layer0_outputs(7688) <= b and not a;
    layer0_outputs(7689) <= not a or b;
    layer0_outputs(7690) <= not a or b;
    layer0_outputs(7691) <= not (a or b);
    layer0_outputs(7692) <= not (a or b);
    layer0_outputs(7693) <= not (a xor b);
    layer0_outputs(7694) <= not a;
    layer0_outputs(7695) <= not (a xor b);
    layer0_outputs(7696) <= '0';
    layer0_outputs(7697) <= not b or a;
    layer0_outputs(7698) <= b and not a;
    layer0_outputs(7699) <= b;
    layer0_outputs(7700) <= a and not b;
    layer0_outputs(7701) <= b;
    layer0_outputs(7702) <= not a or b;
    layer0_outputs(7703) <= '1';
    layer0_outputs(7704) <= not b or a;
    layer0_outputs(7705) <= not (a xor b);
    layer0_outputs(7706) <= not a or b;
    layer0_outputs(7707) <= not a;
    layer0_outputs(7708) <= not a or b;
    layer0_outputs(7709) <= a;
    layer0_outputs(7710) <= a or b;
    layer0_outputs(7711) <= a xor b;
    layer0_outputs(7712) <= not b;
    layer0_outputs(7713) <= b and not a;
    layer0_outputs(7714) <= not a or b;
    layer0_outputs(7715) <= '1';
    layer0_outputs(7716) <= a xor b;
    layer0_outputs(7717) <= a;
    layer0_outputs(7718) <= a;
    layer0_outputs(7719) <= a and b;
    layer0_outputs(7720) <= not a;
    layer0_outputs(7721) <= '0';
    layer0_outputs(7722) <= not a or b;
    layer0_outputs(7723) <= not (a xor b);
    layer0_outputs(7724) <= a and not b;
    layer0_outputs(7725) <= a or b;
    layer0_outputs(7726) <= not (a xor b);
    layer0_outputs(7727) <= a or b;
    layer0_outputs(7728) <= not a or b;
    layer0_outputs(7729) <= not b or a;
    layer0_outputs(7730) <= not b or a;
    layer0_outputs(7731) <= not (a and b);
    layer0_outputs(7732) <= a;
    layer0_outputs(7733) <= not b or a;
    layer0_outputs(7734) <= a xor b;
    layer0_outputs(7735) <= not a or b;
    layer0_outputs(7736) <= not b or a;
    layer0_outputs(7737) <= '1';
    layer0_outputs(7738) <= a xor b;
    layer0_outputs(7739) <= not (a or b);
    layer0_outputs(7740) <= not a;
    layer0_outputs(7741) <= not (a or b);
    layer0_outputs(7742) <= a and not b;
    layer0_outputs(7743) <= a;
    layer0_outputs(7744) <= '1';
    layer0_outputs(7745) <= '1';
    layer0_outputs(7746) <= '1';
    layer0_outputs(7747) <= a;
    layer0_outputs(7748) <= a or b;
    layer0_outputs(7749) <= a and not b;
    layer0_outputs(7750) <= not a;
    layer0_outputs(7751) <= a and b;
    layer0_outputs(7752) <= not (a or b);
    layer0_outputs(7753) <= a or b;
    layer0_outputs(7754) <= a or b;
    layer0_outputs(7755) <= a or b;
    layer0_outputs(7756) <= a;
    layer0_outputs(7757) <= '1';
    layer0_outputs(7758) <= b and not a;
    layer0_outputs(7759) <= not (a xor b);
    layer0_outputs(7760) <= a or b;
    layer0_outputs(7761) <= not (a or b);
    layer0_outputs(7762) <= b and not a;
    layer0_outputs(7763) <= not a;
    layer0_outputs(7764) <= not (a and b);
    layer0_outputs(7765) <= not a;
    layer0_outputs(7766) <= a;
    layer0_outputs(7767) <= a xor b;
    layer0_outputs(7768) <= b and not a;
    layer0_outputs(7769) <= not (a and b);
    layer0_outputs(7770) <= not a;
    layer0_outputs(7771) <= not (a xor b);
    layer0_outputs(7772) <= not b;
    layer0_outputs(7773) <= not (a or b);
    layer0_outputs(7774) <= a or b;
    layer0_outputs(7775) <= a;
    layer0_outputs(7776) <= '0';
    layer0_outputs(7777) <= not (a or b);
    layer0_outputs(7778) <= not (a or b);
    layer0_outputs(7779) <= not a or b;
    layer0_outputs(7780) <= a and b;
    layer0_outputs(7781) <= not (a and b);
    layer0_outputs(7782) <= a or b;
    layer0_outputs(7783) <= not (a xor b);
    layer0_outputs(7784) <= b;
    layer0_outputs(7785) <= not (a xor b);
    layer0_outputs(7786) <= not a;
    layer0_outputs(7787) <= not a or b;
    layer0_outputs(7788) <= b and not a;
    layer0_outputs(7789) <= not b;
    layer0_outputs(7790) <= not a or b;
    layer0_outputs(7791) <= not a or b;
    layer0_outputs(7792) <= a or b;
    layer0_outputs(7793) <= b;
    layer0_outputs(7794) <= b;
    layer0_outputs(7795) <= not (a xor b);
    layer0_outputs(7796) <= not (a or b);
    layer0_outputs(7797) <= not a or b;
    layer0_outputs(7798) <= not (a xor b);
    layer0_outputs(7799) <= '1';
    layer0_outputs(7800) <= not a;
    layer0_outputs(7801) <= a or b;
    layer0_outputs(7802) <= '0';
    layer0_outputs(7803) <= not b;
    layer0_outputs(7804) <= not b;
    layer0_outputs(7805) <= a or b;
    layer0_outputs(7806) <= b and not a;
    layer0_outputs(7807) <= not (a or b);
    layer0_outputs(7808) <= not b or a;
    layer0_outputs(7809) <= not (a or b);
    layer0_outputs(7810) <= b and not a;
    layer0_outputs(7811) <= not (a and b);
    layer0_outputs(7812) <= a and b;
    layer0_outputs(7813) <= '0';
    layer0_outputs(7814) <= not b or a;
    layer0_outputs(7815) <= b;
    layer0_outputs(7816) <= not (a or b);
    layer0_outputs(7817) <= b;
    layer0_outputs(7818) <= not (a and b);
    layer0_outputs(7819) <= not (a and b);
    layer0_outputs(7820) <= a and not b;
    layer0_outputs(7821) <= b and not a;
    layer0_outputs(7822) <= not a;
    layer0_outputs(7823) <= not b or a;
    layer0_outputs(7824) <= a;
    layer0_outputs(7825) <= not (a and b);
    layer0_outputs(7826) <= not (a xor b);
    layer0_outputs(7827) <= a or b;
    layer0_outputs(7828) <= a xor b;
    layer0_outputs(7829) <= b;
    layer0_outputs(7830) <= b and not a;
    layer0_outputs(7831) <= not a or b;
    layer0_outputs(7832) <= not b;
    layer0_outputs(7833) <= a;
    layer0_outputs(7834) <= not b;
    layer0_outputs(7835) <= a xor b;
    layer0_outputs(7836) <= a;
    layer0_outputs(7837) <= a or b;
    layer0_outputs(7838) <= not b;
    layer0_outputs(7839) <= not a or b;
    layer0_outputs(7840) <= not b or a;
    layer0_outputs(7841) <= b and not a;
    layer0_outputs(7842) <= not (a xor b);
    layer0_outputs(7843) <= a;
    layer0_outputs(7844) <= a xor b;
    layer0_outputs(7845) <= not a or b;
    layer0_outputs(7846) <= a and b;
    layer0_outputs(7847) <= not (a xor b);
    layer0_outputs(7848) <= '1';
    layer0_outputs(7849) <= a and b;
    layer0_outputs(7850) <= a;
    layer0_outputs(7851) <= a and b;
    layer0_outputs(7852) <= a;
    layer0_outputs(7853) <= a xor b;
    layer0_outputs(7854) <= not a;
    layer0_outputs(7855) <= not b or a;
    layer0_outputs(7856) <= not (a or b);
    layer0_outputs(7857) <= not a or b;
    layer0_outputs(7858) <= not a or b;
    layer0_outputs(7859) <= not (a or b);
    layer0_outputs(7860) <= a;
    layer0_outputs(7861) <= a or b;
    layer0_outputs(7862) <= not a or b;
    layer0_outputs(7863) <= b;
    layer0_outputs(7864) <= not (a or b);
    layer0_outputs(7865) <= a and b;
    layer0_outputs(7866) <= not (a or b);
    layer0_outputs(7867) <= b and not a;
    layer0_outputs(7868) <= not b;
    layer0_outputs(7869) <= not (a or b);
    layer0_outputs(7870) <= not (a and b);
    layer0_outputs(7871) <= not b;
    layer0_outputs(7872) <= not a;
    layer0_outputs(7873) <= b;
    layer0_outputs(7874) <= a xor b;
    layer0_outputs(7875) <= a;
    layer0_outputs(7876) <= not a;
    layer0_outputs(7877) <= not (a xor b);
    layer0_outputs(7878) <= '0';
    layer0_outputs(7879) <= a or b;
    layer0_outputs(7880) <= a or b;
    layer0_outputs(7881) <= a xor b;
    layer0_outputs(7882) <= not b or a;
    layer0_outputs(7883) <= not (a xor b);
    layer0_outputs(7884) <= a or b;
    layer0_outputs(7885) <= b;
    layer0_outputs(7886) <= a and not b;
    layer0_outputs(7887) <= a or b;
    layer0_outputs(7888) <= not a or b;
    layer0_outputs(7889) <= a and b;
    layer0_outputs(7890) <= not (a xor b);
    layer0_outputs(7891) <= a xor b;
    layer0_outputs(7892) <= a;
    layer0_outputs(7893) <= not (a xor b);
    layer0_outputs(7894) <= a and b;
    layer0_outputs(7895) <= a and not b;
    layer0_outputs(7896) <= a or b;
    layer0_outputs(7897) <= not a or b;
    layer0_outputs(7898) <= '1';
    layer0_outputs(7899) <= not b or a;
    layer0_outputs(7900) <= a and b;
    layer0_outputs(7901) <= not b or a;
    layer0_outputs(7902) <= not b;
    layer0_outputs(7903) <= not b;
    layer0_outputs(7904) <= not a or b;
    layer0_outputs(7905) <= a and not b;
    layer0_outputs(7906) <= '1';
    layer0_outputs(7907) <= '1';
    layer0_outputs(7908) <= '1';
    layer0_outputs(7909) <= b and not a;
    layer0_outputs(7910) <= a and b;
    layer0_outputs(7911) <= '0';
    layer0_outputs(7912) <= a;
    layer0_outputs(7913) <= a or b;
    layer0_outputs(7914) <= a and not b;
    layer0_outputs(7915) <= '1';
    layer0_outputs(7916) <= a xor b;
    layer0_outputs(7917) <= not b;
    layer0_outputs(7918) <= a or b;
    layer0_outputs(7919) <= a and not b;
    layer0_outputs(7920) <= not b or a;
    layer0_outputs(7921) <= a or b;
    layer0_outputs(7922) <= '0';
    layer0_outputs(7923) <= a or b;
    layer0_outputs(7924) <= b;
    layer0_outputs(7925) <= a or b;
    layer0_outputs(7926) <= a or b;
    layer0_outputs(7927) <= a and not b;
    layer0_outputs(7928) <= a and b;
    layer0_outputs(7929) <= '1';
    layer0_outputs(7930) <= b;
    layer0_outputs(7931) <= '1';
    layer0_outputs(7932) <= b;
    layer0_outputs(7933) <= not b;
    layer0_outputs(7934) <= '0';
    layer0_outputs(7935) <= b and not a;
    layer0_outputs(7936) <= a;
    layer0_outputs(7937) <= not b;
    layer0_outputs(7938) <= a and not b;
    layer0_outputs(7939) <= not (a or b);
    layer0_outputs(7940) <= not a;
    layer0_outputs(7941) <= not a;
    layer0_outputs(7942) <= not b or a;
    layer0_outputs(7943) <= a xor b;
    layer0_outputs(7944) <= a and not b;
    layer0_outputs(7945) <= not a;
    layer0_outputs(7946) <= not (a or b);
    layer0_outputs(7947) <= a xor b;
    layer0_outputs(7948) <= not (a or b);
    layer0_outputs(7949) <= a or b;
    layer0_outputs(7950) <= b;
    layer0_outputs(7951) <= not (a and b);
    layer0_outputs(7952) <= a xor b;
    layer0_outputs(7953) <= not a;
    layer0_outputs(7954) <= a;
    layer0_outputs(7955) <= a;
    layer0_outputs(7956) <= not (a or b);
    layer0_outputs(7957) <= not (a or b);
    layer0_outputs(7958) <= not (a or b);
    layer0_outputs(7959) <= a xor b;
    layer0_outputs(7960) <= b and not a;
    layer0_outputs(7961) <= not b;
    layer0_outputs(7962) <= not a;
    layer0_outputs(7963) <= '0';
    layer0_outputs(7964) <= not a;
    layer0_outputs(7965) <= not (a or b);
    layer0_outputs(7966) <= not a;
    layer0_outputs(7967) <= '0';
    layer0_outputs(7968) <= b;
    layer0_outputs(7969) <= a or b;
    layer0_outputs(7970) <= not (a and b);
    layer0_outputs(7971) <= a xor b;
    layer0_outputs(7972) <= not (a or b);
    layer0_outputs(7973) <= not b or a;
    layer0_outputs(7974) <= '1';
    layer0_outputs(7975) <= a or b;
    layer0_outputs(7976) <= a or b;
    layer0_outputs(7977) <= b;
    layer0_outputs(7978) <= a and b;
    layer0_outputs(7979) <= not (a xor b);
    layer0_outputs(7980) <= a;
    layer0_outputs(7981) <= a;
    layer0_outputs(7982) <= a or b;
    layer0_outputs(7983) <= a or b;
    layer0_outputs(7984) <= not a;
    layer0_outputs(7985) <= not b;
    layer0_outputs(7986) <= not b or a;
    layer0_outputs(7987) <= b;
    layer0_outputs(7988) <= a xor b;
    layer0_outputs(7989) <= not b;
    layer0_outputs(7990) <= '0';
    layer0_outputs(7991) <= not (a xor b);
    layer0_outputs(7992) <= '1';
    layer0_outputs(7993) <= a and b;
    layer0_outputs(7994) <= not (a and b);
    layer0_outputs(7995) <= a xor b;
    layer0_outputs(7996) <= not (a or b);
    layer0_outputs(7997) <= b and not a;
    layer0_outputs(7998) <= not (a and b);
    layer0_outputs(7999) <= not (a or b);
    layer0_outputs(8000) <= not (a xor b);
    layer0_outputs(8001) <= not a or b;
    layer0_outputs(8002) <= a and b;
    layer0_outputs(8003) <= not a or b;
    layer0_outputs(8004) <= a xor b;
    layer0_outputs(8005) <= not b;
    layer0_outputs(8006) <= not a;
    layer0_outputs(8007) <= '0';
    layer0_outputs(8008) <= a;
    layer0_outputs(8009) <= a;
    layer0_outputs(8010) <= '0';
    layer0_outputs(8011) <= not a;
    layer0_outputs(8012) <= not a or b;
    layer0_outputs(8013) <= b;
    layer0_outputs(8014) <= not (a and b);
    layer0_outputs(8015) <= a;
    layer0_outputs(8016) <= not a or b;
    layer0_outputs(8017) <= b;
    layer0_outputs(8018) <= a and not b;
    layer0_outputs(8019) <= not (a xor b);
    layer0_outputs(8020) <= a and b;
    layer0_outputs(8021) <= a and not b;
    layer0_outputs(8022) <= b and not a;
    layer0_outputs(8023) <= a or b;
    layer0_outputs(8024) <= '1';
    layer0_outputs(8025) <= not a or b;
    layer0_outputs(8026) <= a or b;
    layer0_outputs(8027) <= a;
    layer0_outputs(8028) <= '1';
    layer0_outputs(8029) <= a xor b;
    layer0_outputs(8030) <= a xor b;
    layer0_outputs(8031) <= not b;
    layer0_outputs(8032) <= not (a or b);
    layer0_outputs(8033) <= a and b;
    layer0_outputs(8034) <= not (a or b);
    layer0_outputs(8035) <= not (a xor b);
    layer0_outputs(8036) <= b and not a;
    layer0_outputs(8037) <= '0';
    layer0_outputs(8038) <= not (a or b);
    layer0_outputs(8039) <= not b or a;
    layer0_outputs(8040) <= '1';
    layer0_outputs(8041) <= a or b;
    layer0_outputs(8042) <= not a;
    layer0_outputs(8043) <= not a;
    layer0_outputs(8044) <= a;
    layer0_outputs(8045) <= a xor b;
    layer0_outputs(8046) <= not a or b;
    layer0_outputs(8047) <= not (a or b);
    layer0_outputs(8048) <= a;
    layer0_outputs(8049) <= a xor b;
    layer0_outputs(8050) <= not (a or b);
    layer0_outputs(8051) <= a;
    layer0_outputs(8052) <= not b;
    layer0_outputs(8053) <= a xor b;
    layer0_outputs(8054) <= not (a and b);
    layer0_outputs(8055) <= not (a or b);
    layer0_outputs(8056) <= not b;
    layer0_outputs(8057) <= not a or b;
    layer0_outputs(8058) <= a and not b;
    layer0_outputs(8059) <= a or b;
    layer0_outputs(8060) <= a and not b;
    layer0_outputs(8061) <= not b;
    layer0_outputs(8062) <= '1';
    layer0_outputs(8063) <= a and b;
    layer0_outputs(8064) <= b and not a;
    layer0_outputs(8065) <= a or b;
    layer0_outputs(8066) <= a and not b;
    layer0_outputs(8067) <= '0';
    layer0_outputs(8068) <= '1';
    layer0_outputs(8069) <= b;
    layer0_outputs(8070) <= not b;
    layer0_outputs(8071) <= a;
    layer0_outputs(8072) <= not (a xor b);
    layer0_outputs(8073) <= not (a xor b);
    layer0_outputs(8074) <= a and b;
    layer0_outputs(8075) <= a;
    layer0_outputs(8076) <= not b;
    layer0_outputs(8077) <= not a;
    layer0_outputs(8078) <= a;
    layer0_outputs(8079) <= a;
    layer0_outputs(8080) <= a;
    layer0_outputs(8081) <= a and not b;
    layer0_outputs(8082) <= a and b;
    layer0_outputs(8083) <= b and not a;
    layer0_outputs(8084) <= a;
    layer0_outputs(8085) <= not (a xor b);
    layer0_outputs(8086) <= not (a and b);
    layer0_outputs(8087) <= a;
    layer0_outputs(8088) <= not b;
    layer0_outputs(8089) <= a or b;
    layer0_outputs(8090) <= b;
    layer0_outputs(8091) <= not a or b;
    layer0_outputs(8092) <= not b;
    layer0_outputs(8093) <= not (a or b);
    layer0_outputs(8094) <= not (a or b);
    layer0_outputs(8095) <= a and not b;
    layer0_outputs(8096) <= '1';
    layer0_outputs(8097) <= a;
    layer0_outputs(8098) <= '0';
    layer0_outputs(8099) <= not (a xor b);
    layer0_outputs(8100) <= b;
    layer0_outputs(8101) <= not b or a;
    layer0_outputs(8102) <= b and not a;
    layer0_outputs(8103) <= not b or a;
    layer0_outputs(8104) <= a;
    layer0_outputs(8105) <= not b;
    layer0_outputs(8106) <= not b or a;
    layer0_outputs(8107) <= not (a xor b);
    layer0_outputs(8108) <= a;
    layer0_outputs(8109) <= b;
    layer0_outputs(8110) <= b;
    layer0_outputs(8111) <= '1';
    layer0_outputs(8112) <= a xor b;
    layer0_outputs(8113) <= b;
    layer0_outputs(8114) <= a xor b;
    layer0_outputs(8115) <= a or b;
    layer0_outputs(8116) <= not b;
    layer0_outputs(8117) <= '1';
    layer0_outputs(8118) <= not (a and b);
    layer0_outputs(8119) <= '1';
    layer0_outputs(8120) <= not a or b;
    layer0_outputs(8121) <= not b;
    layer0_outputs(8122) <= not (a or b);
    layer0_outputs(8123) <= a xor b;
    layer0_outputs(8124) <= not (a xor b);
    layer0_outputs(8125) <= a and not b;
    layer0_outputs(8126) <= b and not a;
    layer0_outputs(8127) <= a or b;
    layer0_outputs(8128) <= '0';
    layer0_outputs(8129) <= b;
    layer0_outputs(8130) <= b and not a;
    layer0_outputs(8131) <= a and b;
    layer0_outputs(8132) <= a;
    layer0_outputs(8133) <= a and not b;
    layer0_outputs(8134) <= a xor b;
    layer0_outputs(8135) <= '1';
    layer0_outputs(8136) <= not (a or b);
    layer0_outputs(8137) <= b and not a;
    layer0_outputs(8138) <= not (a or b);
    layer0_outputs(8139) <= a;
    layer0_outputs(8140) <= a and b;
    layer0_outputs(8141) <= '0';
    layer0_outputs(8142) <= not (a or b);
    layer0_outputs(8143) <= b;
    layer0_outputs(8144) <= b and not a;
    layer0_outputs(8145) <= a or b;
    layer0_outputs(8146) <= a or b;
    layer0_outputs(8147) <= b;
    layer0_outputs(8148) <= not b;
    layer0_outputs(8149) <= b;
    layer0_outputs(8150) <= not (a xor b);
    layer0_outputs(8151) <= '0';
    layer0_outputs(8152) <= not b or a;
    layer0_outputs(8153) <= a;
    layer0_outputs(8154) <= a and b;
    layer0_outputs(8155) <= '1';
    layer0_outputs(8156) <= a xor b;
    layer0_outputs(8157) <= a xor b;
    layer0_outputs(8158) <= not a or b;
    layer0_outputs(8159) <= not a;
    layer0_outputs(8160) <= a;
    layer0_outputs(8161) <= not a;
    layer0_outputs(8162) <= a or b;
    layer0_outputs(8163) <= not (a xor b);
    layer0_outputs(8164) <= not b or a;
    layer0_outputs(8165) <= a and not b;
    layer0_outputs(8166) <= a and b;
    layer0_outputs(8167) <= a xor b;
    layer0_outputs(8168) <= '0';
    layer0_outputs(8169) <= a and b;
    layer0_outputs(8170) <= not a or b;
    layer0_outputs(8171) <= not b;
    layer0_outputs(8172) <= a and not b;
    layer0_outputs(8173) <= a or b;
    layer0_outputs(8174) <= not (a and b);
    layer0_outputs(8175) <= not (a xor b);
    layer0_outputs(8176) <= not a or b;
    layer0_outputs(8177) <= a or b;
    layer0_outputs(8178) <= not b;
    layer0_outputs(8179) <= not a;
    layer0_outputs(8180) <= b;
    layer0_outputs(8181) <= not a;
    layer0_outputs(8182) <= '1';
    layer0_outputs(8183) <= not b;
    layer0_outputs(8184) <= not b;
    layer0_outputs(8185) <= not b;
    layer0_outputs(8186) <= a or b;
    layer0_outputs(8187) <= not a or b;
    layer0_outputs(8188) <= b;
    layer0_outputs(8189) <= b;
    layer0_outputs(8190) <= not (a or b);
    layer0_outputs(8191) <= '0';
    layer0_outputs(8192) <= not b or a;
    layer0_outputs(8193) <= '1';
    layer0_outputs(8194) <= b and not a;
    layer0_outputs(8195) <= a and b;
    layer0_outputs(8196) <= not (a xor b);
    layer0_outputs(8197) <= a and not b;
    layer0_outputs(8198) <= not (a xor b);
    layer0_outputs(8199) <= a or b;
    layer0_outputs(8200) <= not (a or b);
    layer0_outputs(8201) <= not b or a;
    layer0_outputs(8202) <= not (a and b);
    layer0_outputs(8203) <= not (a and b);
    layer0_outputs(8204) <= a and not b;
    layer0_outputs(8205) <= not b or a;
    layer0_outputs(8206) <= a xor b;
    layer0_outputs(8207) <= a and not b;
    layer0_outputs(8208) <= not b or a;
    layer0_outputs(8209) <= not b or a;
    layer0_outputs(8210) <= b;
    layer0_outputs(8211) <= a or b;
    layer0_outputs(8212) <= not a;
    layer0_outputs(8213) <= not a;
    layer0_outputs(8214) <= not (a or b);
    layer0_outputs(8215) <= a xor b;
    layer0_outputs(8216) <= not (a and b);
    layer0_outputs(8217) <= not b;
    layer0_outputs(8218) <= a or b;
    layer0_outputs(8219) <= a xor b;
    layer0_outputs(8220) <= a xor b;
    layer0_outputs(8221) <= not a or b;
    layer0_outputs(8222) <= a and b;
    layer0_outputs(8223) <= '0';
    layer0_outputs(8224) <= not b or a;
    layer0_outputs(8225) <= a and b;
    layer0_outputs(8226) <= '1';
    layer0_outputs(8227) <= '0';
    layer0_outputs(8228) <= b;
    layer0_outputs(8229) <= b and not a;
    layer0_outputs(8230) <= not b;
    layer0_outputs(8231) <= b;
    layer0_outputs(8232) <= b and not a;
    layer0_outputs(8233) <= '1';
    layer0_outputs(8234) <= not b;
    layer0_outputs(8235) <= a and not b;
    layer0_outputs(8236) <= a or b;
    layer0_outputs(8237) <= '1';
    layer0_outputs(8238) <= b and not a;
    layer0_outputs(8239) <= not a;
    layer0_outputs(8240) <= not (a or b);
    layer0_outputs(8241) <= not b or a;
    layer0_outputs(8242) <= '0';
    layer0_outputs(8243) <= b and not a;
    layer0_outputs(8244) <= '0';
    layer0_outputs(8245) <= a or b;
    layer0_outputs(8246) <= b;
    layer0_outputs(8247) <= a or b;
    layer0_outputs(8248) <= b and not a;
    layer0_outputs(8249) <= b;
    layer0_outputs(8250) <= not b or a;
    layer0_outputs(8251) <= '1';
    layer0_outputs(8252) <= not (a and b);
    layer0_outputs(8253) <= not a or b;
    layer0_outputs(8254) <= not b;
    layer0_outputs(8255) <= '0';
    layer0_outputs(8256) <= a and b;
    layer0_outputs(8257) <= not b or a;
    layer0_outputs(8258) <= a and not b;
    layer0_outputs(8259) <= a and not b;
    layer0_outputs(8260) <= a;
    layer0_outputs(8261) <= not b;
    layer0_outputs(8262) <= not a;
    layer0_outputs(8263) <= a xor b;
    layer0_outputs(8264) <= not (a xor b);
    layer0_outputs(8265) <= '1';
    layer0_outputs(8266) <= not a;
    layer0_outputs(8267) <= a and not b;
    layer0_outputs(8268) <= not b or a;
    layer0_outputs(8269) <= b;
    layer0_outputs(8270) <= not (a and b);
    layer0_outputs(8271) <= not a;
    layer0_outputs(8272) <= a and b;
    layer0_outputs(8273) <= not a or b;
    layer0_outputs(8274) <= a or b;
    layer0_outputs(8275) <= a;
    layer0_outputs(8276) <= not b or a;
    layer0_outputs(8277) <= a or b;
    layer0_outputs(8278) <= not (a or b);
    layer0_outputs(8279) <= a and not b;
    layer0_outputs(8280) <= not b;
    layer0_outputs(8281) <= '1';
    layer0_outputs(8282) <= b;
    layer0_outputs(8283) <= a;
    layer0_outputs(8284) <= a xor b;
    layer0_outputs(8285) <= '1';
    layer0_outputs(8286) <= a;
    layer0_outputs(8287) <= not (a and b);
    layer0_outputs(8288) <= a;
    layer0_outputs(8289) <= a or b;
    layer0_outputs(8290) <= not a;
    layer0_outputs(8291) <= not (a or b);
    layer0_outputs(8292) <= b and not a;
    layer0_outputs(8293) <= a or b;
    layer0_outputs(8294) <= '0';
    layer0_outputs(8295) <= not b;
    layer0_outputs(8296) <= not b;
    layer0_outputs(8297) <= '0';
    layer0_outputs(8298) <= '1';
    layer0_outputs(8299) <= not (a and b);
    layer0_outputs(8300) <= a or b;
    layer0_outputs(8301) <= not b or a;
    layer0_outputs(8302) <= a or b;
    layer0_outputs(8303) <= not b;
    layer0_outputs(8304) <= a;
    layer0_outputs(8305) <= b;
    layer0_outputs(8306) <= not b or a;
    layer0_outputs(8307) <= a and b;
    layer0_outputs(8308) <= not a;
    layer0_outputs(8309) <= not a or b;
    layer0_outputs(8310) <= not (a xor b);
    layer0_outputs(8311) <= a or b;
    layer0_outputs(8312) <= not (a xor b);
    layer0_outputs(8313) <= b and not a;
    layer0_outputs(8314) <= a and b;
    layer0_outputs(8315) <= '0';
    layer0_outputs(8316) <= a and b;
    layer0_outputs(8317) <= b;
    layer0_outputs(8318) <= a;
    layer0_outputs(8319) <= a and b;
    layer0_outputs(8320) <= not a or b;
    layer0_outputs(8321) <= b and not a;
    layer0_outputs(8322) <= not a;
    layer0_outputs(8323) <= '1';
    layer0_outputs(8324) <= a and not b;
    layer0_outputs(8325) <= not b;
    layer0_outputs(8326) <= not (a xor b);
    layer0_outputs(8327) <= not a or b;
    layer0_outputs(8328) <= not (a or b);
    layer0_outputs(8329) <= b and not a;
    layer0_outputs(8330) <= not (a xor b);
    layer0_outputs(8331) <= not a;
    layer0_outputs(8332) <= not (a or b);
    layer0_outputs(8333) <= not b;
    layer0_outputs(8334) <= a;
    layer0_outputs(8335) <= not (a and b);
    layer0_outputs(8336) <= not b or a;
    layer0_outputs(8337) <= '0';
    layer0_outputs(8338) <= a and b;
    layer0_outputs(8339) <= a and not b;
    layer0_outputs(8340) <= a or b;
    layer0_outputs(8341) <= not a or b;
    layer0_outputs(8342) <= a or b;
    layer0_outputs(8343) <= not (a or b);
    layer0_outputs(8344) <= not b;
    layer0_outputs(8345) <= not a;
    layer0_outputs(8346) <= a and not b;
    layer0_outputs(8347) <= b;
    layer0_outputs(8348) <= b;
    layer0_outputs(8349) <= a and b;
    layer0_outputs(8350) <= not a;
    layer0_outputs(8351) <= not a;
    layer0_outputs(8352) <= not b or a;
    layer0_outputs(8353) <= not b;
    layer0_outputs(8354) <= not (a and b);
    layer0_outputs(8355) <= not b;
    layer0_outputs(8356) <= b;
    layer0_outputs(8357) <= a xor b;
    layer0_outputs(8358) <= a or b;
    layer0_outputs(8359) <= a xor b;
    layer0_outputs(8360) <= not a;
    layer0_outputs(8361) <= not a;
    layer0_outputs(8362) <= not (a or b);
    layer0_outputs(8363) <= not (a or b);
    layer0_outputs(8364) <= not b or a;
    layer0_outputs(8365) <= b;
    layer0_outputs(8366) <= b;
    layer0_outputs(8367) <= a and not b;
    layer0_outputs(8368) <= not a;
    layer0_outputs(8369) <= b and not a;
    layer0_outputs(8370) <= not b or a;
    layer0_outputs(8371) <= b and not a;
    layer0_outputs(8372) <= not b;
    layer0_outputs(8373) <= not a;
    layer0_outputs(8374) <= b;
    layer0_outputs(8375) <= a and not b;
    layer0_outputs(8376) <= a or b;
    layer0_outputs(8377) <= b;
    layer0_outputs(8378) <= a and b;
    layer0_outputs(8379) <= a and b;
    layer0_outputs(8380) <= b and not a;
    layer0_outputs(8381) <= not b or a;
    layer0_outputs(8382) <= not a or b;
    layer0_outputs(8383) <= not (a or b);
    layer0_outputs(8384) <= not b or a;
    layer0_outputs(8385) <= not (a and b);
    layer0_outputs(8386) <= b and not a;
    layer0_outputs(8387) <= not (a and b);
    layer0_outputs(8388) <= a xor b;
    layer0_outputs(8389) <= not a or b;
    layer0_outputs(8390) <= b;
    layer0_outputs(8391) <= a and b;
    layer0_outputs(8392) <= a xor b;
    layer0_outputs(8393) <= not b or a;
    layer0_outputs(8394) <= not a;
    layer0_outputs(8395) <= a and not b;
    layer0_outputs(8396) <= b and not a;
    layer0_outputs(8397) <= not a or b;
    layer0_outputs(8398) <= '1';
    layer0_outputs(8399) <= not b;
    layer0_outputs(8400) <= not a;
    layer0_outputs(8401) <= '0';
    layer0_outputs(8402) <= b and not a;
    layer0_outputs(8403) <= not a;
    layer0_outputs(8404) <= not a or b;
    layer0_outputs(8405) <= a;
    layer0_outputs(8406) <= a xor b;
    layer0_outputs(8407) <= not a;
    layer0_outputs(8408) <= a xor b;
    layer0_outputs(8409) <= not (a xor b);
    layer0_outputs(8410) <= '0';
    layer0_outputs(8411) <= '1';
    layer0_outputs(8412) <= not b or a;
    layer0_outputs(8413) <= not (a and b);
    layer0_outputs(8414) <= a;
    layer0_outputs(8415) <= not b;
    layer0_outputs(8416) <= a or b;
    layer0_outputs(8417) <= a or b;
    layer0_outputs(8418) <= not a;
    layer0_outputs(8419) <= '0';
    layer0_outputs(8420) <= '0';
    layer0_outputs(8421) <= a and not b;
    layer0_outputs(8422) <= a and not b;
    layer0_outputs(8423) <= a or b;
    layer0_outputs(8424) <= not b;
    layer0_outputs(8425) <= a;
    layer0_outputs(8426) <= not (a or b);
    layer0_outputs(8427) <= not (a or b);
    layer0_outputs(8428) <= b and not a;
    layer0_outputs(8429) <= a xor b;
    layer0_outputs(8430) <= b;
    layer0_outputs(8431) <= not (a xor b);
    layer0_outputs(8432) <= a and b;
    layer0_outputs(8433) <= not a or b;
    layer0_outputs(8434) <= a and not b;
    layer0_outputs(8435) <= a and b;
    layer0_outputs(8436) <= not (a or b);
    layer0_outputs(8437) <= not b;
    layer0_outputs(8438) <= a;
    layer0_outputs(8439) <= a and not b;
    layer0_outputs(8440) <= a and b;
    layer0_outputs(8441) <= not (a or b);
    layer0_outputs(8442) <= not b or a;
    layer0_outputs(8443) <= not b or a;
    layer0_outputs(8444) <= '0';
    layer0_outputs(8445) <= '1';
    layer0_outputs(8446) <= not a or b;
    layer0_outputs(8447) <= b and not a;
    layer0_outputs(8448) <= a and not b;
    layer0_outputs(8449) <= a and not b;
    layer0_outputs(8450) <= a or b;
    layer0_outputs(8451) <= a xor b;
    layer0_outputs(8452) <= not (a or b);
    layer0_outputs(8453) <= a xor b;
    layer0_outputs(8454) <= not (a and b);
    layer0_outputs(8455) <= '0';
    layer0_outputs(8456) <= not (a and b);
    layer0_outputs(8457) <= b and not a;
    layer0_outputs(8458) <= a;
    layer0_outputs(8459) <= b and not a;
    layer0_outputs(8460) <= a or b;
    layer0_outputs(8461) <= not (a or b);
    layer0_outputs(8462) <= b;
    layer0_outputs(8463) <= not (a or b);
    layer0_outputs(8464) <= a;
    layer0_outputs(8465) <= not (a and b);
    layer0_outputs(8466) <= b and not a;
    layer0_outputs(8467) <= '0';
    layer0_outputs(8468) <= not a or b;
    layer0_outputs(8469) <= not a;
    layer0_outputs(8470) <= a xor b;
    layer0_outputs(8471) <= not (a and b);
    layer0_outputs(8472) <= not b or a;
    layer0_outputs(8473) <= b;
    layer0_outputs(8474) <= '0';
    layer0_outputs(8475) <= '0';
    layer0_outputs(8476) <= b;
    layer0_outputs(8477) <= a and not b;
    layer0_outputs(8478) <= not a or b;
    layer0_outputs(8479) <= not (a and b);
    layer0_outputs(8480) <= a and b;
    layer0_outputs(8481) <= not b;
    layer0_outputs(8482) <= a and not b;
    layer0_outputs(8483) <= not b or a;
    layer0_outputs(8484) <= not (a xor b);
    layer0_outputs(8485) <= b;
    layer0_outputs(8486) <= a and not b;
    layer0_outputs(8487) <= not a or b;
    layer0_outputs(8488) <= b;
    layer0_outputs(8489) <= a and b;
    layer0_outputs(8490) <= a and not b;
    layer0_outputs(8491) <= not (a xor b);
    layer0_outputs(8492) <= '1';
    layer0_outputs(8493) <= not a;
    layer0_outputs(8494) <= not a;
    layer0_outputs(8495) <= not (a or b);
    layer0_outputs(8496) <= not (a xor b);
    layer0_outputs(8497) <= a xor b;
    layer0_outputs(8498) <= not b;
    layer0_outputs(8499) <= a or b;
    layer0_outputs(8500) <= a xor b;
    layer0_outputs(8501) <= a or b;
    layer0_outputs(8502) <= not b;
    layer0_outputs(8503) <= '0';
    layer0_outputs(8504) <= a;
    layer0_outputs(8505) <= a xor b;
    layer0_outputs(8506) <= not (a and b);
    layer0_outputs(8507) <= a xor b;
    layer0_outputs(8508) <= a or b;
    layer0_outputs(8509) <= not a;
    layer0_outputs(8510) <= not (a or b);
    layer0_outputs(8511) <= b;
    layer0_outputs(8512) <= a and b;
    layer0_outputs(8513) <= b;
    layer0_outputs(8514) <= not a or b;
    layer0_outputs(8515) <= a or b;
    layer0_outputs(8516) <= not (a xor b);
    layer0_outputs(8517) <= not b or a;
    layer0_outputs(8518) <= b;
    layer0_outputs(8519) <= not a;
    layer0_outputs(8520) <= not b;
    layer0_outputs(8521) <= a xor b;
    layer0_outputs(8522) <= not (a or b);
    layer0_outputs(8523) <= a xor b;
    layer0_outputs(8524) <= not a or b;
    layer0_outputs(8525) <= a xor b;
    layer0_outputs(8526) <= not b;
    layer0_outputs(8527) <= b;
    layer0_outputs(8528) <= not (a and b);
    layer0_outputs(8529) <= a;
    layer0_outputs(8530) <= b and not a;
    layer0_outputs(8531) <= not b or a;
    layer0_outputs(8532) <= b and not a;
    layer0_outputs(8533) <= not b or a;
    layer0_outputs(8534) <= not b;
    layer0_outputs(8535) <= not a or b;
    layer0_outputs(8536) <= a or b;
    layer0_outputs(8537) <= '0';
    layer0_outputs(8538) <= b and not a;
    layer0_outputs(8539) <= b;
    layer0_outputs(8540) <= b;
    layer0_outputs(8541) <= not (a and b);
    layer0_outputs(8542) <= a;
    layer0_outputs(8543) <= b and not a;
    layer0_outputs(8544) <= a;
    layer0_outputs(8545) <= '1';
    layer0_outputs(8546) <= not (a xor b);
    layer0_outputs(8547) <= a and not b;
    layer0_outputs(8548) <= a and not b;
    layer0_outputs(8549) <= '0';
    layer0_outputs(8550) <= not (a or b);
    layer0_outputs(8551) <= a or b;
    layer0_outputs(8552) <= a or b;
    layer0_outputs(8553) <= not a;
    layer0_outputs(8554) <= not (a and b);
    layer0_outputs(8555) <= not (a or b);
    layer0_outputs(8556) <= '1';
    layer0_outputs(8557) <= a xor b;
    layer0_outputs(8558) <= not b;
    layer0_outputs(8559) <= b;
    layer0_outputs(8560) <= b and not a;
    layer0_outputs(8561) <= not b;
    layer0_outputs(8562) <= a or b;
    layer0_outputs(8563) <= not a or b;
    layer0_outputs(8564) <= b and not a;
    layer0_outputs(8565) <= b;
    layer0_outputs(8566) <= '0';
    layer0_outputs(8567) <= a and not b;
    layer0_outputs(8568) <= a and not b;
    layer0_outputs(8569) <= not (a xor b);
    layer0_outputs(8570) <= a or b;
    layer0_outputs(8571) <= a xor b;
    layer0_outputs(8572) <= a;
    layer0_outputs(8573) <= b and not a;
    layer0_outputs(8574) <= b and not a;
    layer0_outputs(8575) <= a and b;
    layer0_outputs(8576) <= not (a or b);
    layer0_outputs(8577) <= not a;
    layer0_outputs(8578) <= not b or a;
    layer0_outputs(8579) <= a xor b;
    layer0_outputs(8580) <= a or b;
    layer0_outputs(8581) <= not a or b;
    layer0_outputs(8582) <= a and not b;
    layer0_outputs(8583) <= a or b;
    layer0_outputs(8584) <= not (a or b);
    layer0_outputs(8585) <= a;
    layer0_outputs(8586) <= not (a or b);
    layer0_outputs(8587) <= not (a and b);
    layer0_outputs(8588) <= not a;
    layer0_outputs(8589) <= a;
    layer0_outputs(8590) <= a and b;
    layer0_outputs(8591) <= '1';
    layer0_outputs(8592) <= not b;
    layer0_outputs(8593) <= b and not a;
    layer0_outputs(8594) <= a or b;
    layer0_outputs(8595) <= a;
    layer0_outputs(8596) <= a or b;
    layer0_outputs(8597) <= a and not b;
    layer0_outputs(8598) <= a xor b;
    layer0_outputs(8599) <= b;
    layer0_outputs(8600) <= not (a and b);
    layer0_outputs(8601) <= not a;
    layer0_outputs(8602) <= not b;
    layer0_outputs(8603) <= not (a or b);
    layer0_outputs(8604) <= a;
    layer0_outputs(8605) <= a xor b;
    layer0_outputs(8606) <= a;
    layer0_outputs(8607) <= '1';
    layer0_outputs(8608) <= not a or b;
    layer0_outputs(8609) <= not (a and b);
    layer0_outputs(8610) <= a or b;
    layer0_outputs(8611) <= not (a or b);
    layer0_outputs(8612) <= not a or b;
    layer0_outputs(8613) <= a and not b;
    layer0_outputs(8614) <= a xor b;
    layer0_outputs(8615) <= b;
    layer0_outputs(8616) <= not a or b;
    layer0_outputs(8617) <= a;
    layer0_outputs(8618) <= not (a xor b);
    layer0_outputs(8619) <= not (a xor b);
    layer0_outputs(8620) <= '0';
    layer0_outputs(8621) <= a xor b;
    layer0_outputs(8622) <= '0';
    layer0_outputs(8623) <= a or b;
    layer0_outputs(8624) <= not b;
    layer0_outputs(8625) <= b and not a;
    layer0_outputs(8626) <= b;
    layer0_outputs(8627) <= a and not b;
    layer0_outputs(8628) <= b;
    layer0_outputs(8629) <= a;
    layer0_outputs(8630) <= not b;
    layer0_outputs(8631) <= a and b;
    layer0_outputs(8632) <= not a or b;
    layer0_outputs(8633) <= a or b;
    layer0_outputs(8634) <= a or b;
    layer0_outputs(8635) <= not b;
    layer0_outputs(8636) <= a and b;
    layer0_outputs(8637) <= a xor b;
    layer0_outputs(8638) <= not (a xor b);
    layer0_outputs(8639) <= '1';
    layer0_outputs(8640) <= not b;
    layer0_outputs(8641) <= a and b;
    layer0_outputs(8642) <= not (a and b);
    layer0_outputs(8643) <= a;
    layer0_outputs(8644) <= '1';
    layer0_outputs(8645) <= b;
    layer0_outputs(8646) <= a or b;
    layer0_outputs(8647) <= a and not b;
    layer0_outputs(8648) <= '1';
    layer0_outputs(8649) <= not (a or b);
    layer0_outputs(8650) <= a and not b;
    layer0_outputs(8651) <= b and not a;
    layer0_outputs(8652) <= '0';
    layer0_outputs(8653) <= not a;
    layer0_outputs(8654) <= b and not a;
    layer0_outputs(8655) <= not a;
    layer0_outputs(8656) <= not b;
    layer0_outputs(8657) <= '1';
    layer0_outputs(8658) <= b;
    layer0_outputs(8659) <= a and not b;
    layer0_outputs(8660) <= not a;
    layer0_outputs(8661) <= '1';
    layer0_outputs(8662) <= a or b;
    layer0_outputs(8663) <= a or b;
    layer0_outputs(8664) <= not b or a;
    layer0_outputs(8665) <= a;
    layer0_outputs(8666) <= '0';
    layer0_outputs(8667) <= not a;
    layer0_outputs(8668) <= not a;
    layer0_outputs(8669) <= '1';
    layer0_outputs(8670) <= b;
    layer0_outputs(8671) <= a and b;
    layer0_outputs(8672) <= not a;
    layer0_outputs(8673) <= not a or b;
    layer0_outputs(8674) <= '1';
    layer0_outputs(8675) <= not a;
    layer0_outputs(8676) <= b and not a;
    layer0_outputs(8677) <= a or b;
    layer0_outputs(8678) <= b and not a;
    layer0_outputs(8679) <= a xor b;
    layer0_outputs(8680) <= not b;
    layer0_outputs(8681) <= not (a and b);
    layer0_outputs(8682) <= not (a or b);
    layer0_outputs(8683) <= not (a xor b);
    layer0_outputs(8684) <= a xor b;
    layer0_outputs(8685) <= '1';
    layer0_outputs(8686) <= a;
    layer0_outputs(8687) <= not (a or b);
    layer0_outputs(8688) <= a and not b;
    layer0_outputs(8689) <= not b or a;
    layer0_outputs(8690) <= not (a xor b);
    layer0_outputs(8691) <= not b or a;
    layer0_outputs(8692) <= not (a and b);
    layer0_outputs(8693) <= not (a or b);
    layer0_outputs(8694) <= '1';
    layer0_outputs(8695) <= not (a and b);
    layer0_outputs(8696) <= not b;
    layer0_outputs(8697) <= '1';
    layer0_outputs(8698) <= a;
    layer0_outputs(8699) <= not b;
    layer0_outputs(8700) <= a or b;
    layer0_outputs(8701) <= '1';
    layer0_outputs(8702) <= b;
    layer0_outputs(8703) <= a or b;
    layer0_outputs(8704) <= '1';
    layer0_outputs(8705) <= a and not b;
    layer0_outputs(8706) <= a or b;
    layer0_outputs(8707) <= not b;
    layer0_outputs(8708) <= a and not b;
    layer0_outputs(8709) <= not (a or b);
    layer0_outputs(8710) <= not b;
    layer0_outputs(8711) <= '1';
    layer0_outputs(8712) <= not (a xor b);
    layer0_outputs(8713) <= b and not a;
    layer0_outputs(8714) <= not (a or b);
    layer0_outputs(8715) <= not a;
    layer0_outputs(8716) <= b;
    layer0_outputs(8717) <= not (a xor b);
    layer0_outputs(8718) <= '1';
    layer0_outputs(8719) <= not a;
    layer0_outputs(8720) <= a and not b;
    layer0_outputs(8721) <= not b;
    layer0_outputs(8722) <= a;
    layer0_outputs(8723) <= not (a or b);
    layer0_outputs(8724) <= '1';
    layer0_outputs(8725) <= a and not b;
    layer0_outputs(8726) <= b;
    layer0_outputs(8727) <= not a;
    layer0_outputs(8728) <= a or b;
    layer0_outputs(8729) <= not (a xor b);
    layer0_outputs(8730) <= a or b;
    layer0_outputs(8731) <= a xor b;
    layer0_outputs(8732) <= not a or b;
    layer0_outputs(8733) <= '0';
    layer0_outputs(8734) <= a xor b;
    layer0_outputs(8735) <= not a;
    layer0_outputs(8736) <= a and b;
    layer0_outputs(8737) <= not a;
    layer0_outputs(8738) <= '0';
    layer0_outputs(8739) <= not b;
    layer0_outputs(8740) <= '0';
    layer0_outputs(8741) <= not a;
    layer0_outputs(8742) <= a;
    layer0_outputs(8743) <= not a;
    layer0_outputs(8744) <= a xor b;
    layer0_outputs(8745) <= not a;
    layer0_outputs(8746) <= a xor b;
    layer0_outputs(8747) <= a or b;
    layer0_outputs(8748) <= not b or a;
    layer0_outputs(8749) <= b;
    layer0_outputs(8750) <= not (a and b);
    layer0_outputs(8751) <= not (a and b);
    layer0_outputs(8752) <= not (a or b);
    layer0_outputs(8753) <= not (a xor b);
    layer0_outputs(8754) <= '0';
    layer0_outputs(8755) <= not b or a;
    layer0_outputs(8756) <= a xor b;
    layer0_outputs(8757) <= b and not a;
    layer0_outputs(8758) <= not a;
    layer0_outputs(8759) <= b;
    layer0_outputs(8760) <= not (a or b);
    layer0_outputs(8761) <= not b;
    layer0_outputs(8762) <= not a;
    layer0_outputs(8763) <= a or b;
    layer0_outputs(8764) <= not (a or b);
    layer0_outputs(8765) <= not (a xor b);
    layer0_outputs(8766) <= a;
    layer0_outputs(8767) <= a and b;
    layer0_outputs(8768) <= '1';
    layer0_outputs(8769) <= not (a and b);
    layer0_outputs(8770) <= not (a or b);
    layer0_outputs(8771) <= a or b;
    layer0_outputs(8772) <= not a or b;
    layer0_outputs(8773) <= b;
    layer0_outputs(8774) <= not a or b;
    layer0_outputs(8775) <= a and not b;
    layer0_outputs(8776) <= b;
    layer0_outputs(8777) <= not (a xor b);
    layer0_outputs(8778) <= not a or b;
    layer0_outputs(8779) <= not b;
    layer0_outputs(8780) <= a xor b;
    layer0_outputs(8781) <= not (a and b);
    layer0_outputs(8782) <= b and not a;
    layer0_outputs(8783) <= not a;
    layer0_outputs(8784) <= not b;
    layer0_outputs(8785) <= a and not b;
    layer0_outputs(8786) <= a and b;
    layer0_outputs(8787) <= not (a and b);
    layer0_outputs(8788) <= a and b;
    layer0_outputs(8789) <= a or b;
    layer0_outputs(8790) <= not b or a;
    layer0_outputs(8791) <= not b or a;
    layer0_outputs(8792) <= not a or b;
    layer0_outputs(8793) <= not a;
    layer0_outputs(8794) <= a xor b;
    layer0_outputs(8795) <= b;
    layer0_outputs(8796) <= a;
    layer0_outputs(8797) <= a and not b;
    layer0_outputs(8798) <= '1';
    layer0_outputs(8799) <= not a or b;
    layer0_outputs(8800) <= not (a or b);
    layer0_outputs(8801) <= a and not b;
    layer0_outputs(8802) <= a or b;
    layer0_outputs(8803) <= not (a or b);
    layer0_outputs(8804) <= '1';
    layer0_outputs(8805) <= a;
    layer0_outputs(8806) <= b and not a;
    layer0_outputs(8807) <= not a;
    layer0_outputs(8808) <= not (a and b);
    layer0_outputs(8809) <= b;
    layer0_outputs(8810) <= a;
    layer0_outputs(8811) <= '0';
    layer0_outputs(8812) <= b and not a;
    layer0_outputs(8813) <= a and b;
    layer0_outputs(8814) <= b;
    layer0_outputs(8815) <= a;
    layer0_outputs(8816) <= not a;
    layer0_outputs(8817) <= not b or a;
    layer0_outputs(8818) <= a and not b;
    layer0_outputs(8819) <= a and not b;
    layer0_outputs(8820) <= a xor b;
    layer0_outputs(8821) <= a or b;
    layer0_outputs(8822) <= b and not a;
    layer0_outputs(8823) <= '1';
    layer0_outputs(8824) <= a and not b;
    layer0_outputs(8825) <= b and not a;
    layer0_outputs(8826) <= a or b;
    layer0_outputs(8827) <= not (a and b);
    layer0_outputs(8828) <= b;
    layer0_outputs(8829) <= not b or a;
    layer0_outputs(8830) <= not b;
    layer0_outputs(8831) <= not a or b;
    layer0_outputs(8832) <= b;
    layer0_outputs(8833) <= '1';
    layer0_outputs(8834) <= a and not b;
    layer0_outputs(8835) <= not b or a;
    layer0_outputs(8836) <= '1';
    layer0_outputs(8837) <= not b;
    layer0_outputs(8838) <= not b;
    layer0_outputs(8839) <= a and not b;
    layer0_outputs(8840) <= a or b;
    layer0_outputs(8841) <= not a or b;
    layer0_outputs(8842) <= '0';
    layer0_outputs(8843) <= a;
    layer0_outputs(8844) <= not a or b;
    layer0_outputs(8845) <= a or b;
    layer0_outputs(8846) <= not b;
    layer0_outputs(8847) <= b;
    layer0_outputs(8848) <= not a or b;
    layer0_outputs(8849) <= '0';
    layer0_outputs(8850) <= a;
    layer0_outputs(8851) <= a;
    layer0_outputs(8852) <= b;
    layer0_outputs(8853) <= '0';
    layer0_outputs(8854) <= not b or a;
    layer0_outputs(8855) <= a and not b;
    layer0_outputs(8856) <= not a or b;
    layer0_outputs(8857) <= a and b;
    layer0_outputs(8858) <= a or b;
    layer0_outputs(8859) <= b;
    layer0_outputs(8860) <= not a or b;
    layer0_outputs(8861) <= not a or b;
    layer0_outputs(8862) <= a;
    layer0_outputs(8863) <= '0';
    layer0_outputs(8864) <= not (a or b);
    layer0_outputs(8865) <= a and b;
    layer0_outputs(8866) <= a xor b;
    layer0_outputs(8867) <= not a or b;
    layer0_outputs(8868) <= not b or a;
    layer0_outputs(8869) <= not (a and b);
    layer0_outputs(8870) <= a and b;
    layer0_outputs(8871) <= '1';
    layer0_outputs(8872) <= a and b;
    layer0_outputs(8873) <= not a;
    layer0_outputs(8874) <= a or b;
    layer0_outputs(8875) <= b;
    layer0_outputs(8876) <= not a;
    layer0_outputs(8877) <= not b;
    layer0_outputs(8878) <= a and not b;
    layer0_outputs(8879) <= a or b;
    layer0_outputs(8880) <= not (a and b);
    layer0_outputs(8881) <= not b or a;
    layer0_outputs(8882) <= not (a and b);
    layer0_outputs(8883) <= not a or b;
    layer0_outputs(8884) <= '0';
    layer0_outputs(8885) <= a;
    layer0_outputs(8886) <= a;
    layer0_outputs(8887) <= a and not b;
    layer0_outputs(8888) <= not (a or b);
    layer0_outputs(8889) <= not (a xor b);
    layer0_outputs(8890) <= not a;
    layer0_outputs(8891) <= a;
    layer0_outputs(8892) <= not a;
    layer0_outputs(8893) <= a xor b;
    layer0_outputs(8894) <= b and not a;
    layer0_outputs(8895) <= not (a and b);
    layer0_outputs(8896) <= not b or a;
    layer0_outputs(8897) <= not (a or b);
    layer0_outputs(8898) <= '1';
    layer0_outputs(8899) <= not a or b;
    layer0_outputs(8900) <= not a;
    layer0_outputs(8901) <= not (a or b);
    layer0_outputs(8902) <= not a or b;
    layer0_outputs(8903) <= not b or a;
    layer0_outputs(8904) <= not (a or b);
    layer0_outputs(8905) <= a xor b;
    layer0_outputs(8906) <= not a or b;
    layer0_outputs(8907) <= not a;
    layer0_outputs(8908) <= a and b;
    layer0_outputs(8909) <= not a;
    layer0_outputs(8910) <= not (a xor b);
    layer0_outputs(8911) <= b;
    layer0_outputs(8912) <= not b;
    layer0_outputs(8913) <= a;
    layer0_outputs(8914) <= a and b;
    layer0_outputs(8915) <= '0';
    layer0_outputs(8916) <= b;
    layer0_outputs(8917) <= not a or b;
    layer0_outputs(8918) <= b and not a;
    layer0_outputs(8919) <= a or b;
    layer0_outputs(8920) <= b and not a;
    layer0_outputs(8921) <= a or b;
    layer0_outputs(8922) <= not b;
    layer0_outputs(8923) <= a or b;
    layer0_outputs(8924) <= not (a or b);
    layer0_outputs(8925) <= not (a xor b);
    layer0_outputs(8926) <= not a;
    layer0_outputs(8927) <= a;
    layer0_outputs(8928) <= not b;
    layer0_outputs(8929) <= a;
    layer0_outputs(8930) <= not (a and b);
    layer0_outputs(8931) <= a and not b;
    layer0_outputs(8932) <= a or b;
    layer0_outputs(8933) <= a and b;
    layer0_outputs(8934) <= a xor b;
    layer0_outputs(8935) <= not b or a;
    layer0_outputs(8936) <= a and not b;
    layer0_outputs(8937) <= not b;
    layer0_outputs(8938) <= a and not b;
    layer0_outputs(8939) <= not a;
    layer0_outputs(8940) <= '1';
    layer0_outputs(8941) <= b;
    layer0_outputs(8942) <= not a or b;
    layer0_outputs(8943) <= not (a or b);
    layer0_outputs(8944) <= not (a or b);
    layer0_outputs(8945) <= not (a and b);
    layer0_outputs(8946) <= '0';
    layer0_outputs(8947) <= a or b;
    layer0_outputs(8948) <= a and b;
    layer0_outputs(8949) <= not a;
    layer0_outputs(8950) <= '0';
    layer0_outputs(8951) <= a or b;
    layer0_outputs(8952) <= not b;
    layer0_outputs(8953) <= a;
    layer0_outputs(8954) <= a or b;
    layer0_outputs(8955) <= not (a and b);
    layer0_outputs(8956) <= not (a and b);
    layer0_outputs(8957) <= '0';
    layer0_outputs(8958) <= not a or b;
    layer0_outputs(8959) <= not b or a;
    layer0_outputs(8960) <= a and not b;
    layer0_outputs(8961) <= '0';
    layer0_outputs(8962) <= a or b;
    layer0_outputs(8963) <= a and not b;
    layer0_outputs(8964) <= b and not a;
    layer0_outputs(8965) <= not b;
    layer0_outputs(8966) <= a and b;
    layer0_outputs(8967) <= a xor b;
    layer0_outputs(8968) <= a xor b;
    layer0_outputs(8969) <= not (a xor b);
    layer0_outputs(8970) <= '1';
    layer0_outputs(8971) <= b and not a;
    layer0_outputs(8972) <= a and not b;
    layer0_outputs(8973) <= not (a and b);
    layer0_outputs(8974) <= not (a or b);
    layer0_outputs(8975) <= a xor b;
    layer0_outputs(8976) <= not (a or b);
    layer0_outputs(8977) <= not a or b;
    layer0_outputs(8978) <= '0';
    layer0_outputs(8979) <= a;
    layer0_outputs(8980) <= a xor b;
    layer0_outputs(8981) <= '1';
    layer0_outputs(8982) <= '1';
    layer0_outputs(8983) <= b;
    layer0_outputs(8984) <= a and not b;
    layer0_outputs(8985) <= not (a or b);
    layer0_outputs(8986) <= not (a or b);
    layer0_outputs(8987) <= a and not b;
    layer0_outputs(8988) <= not (a or b);
    layer0_outputs(8989) <= not (a or b);
    layer0_outputs(8990) <= b and not a;
    layer0_outputs(8991) <= a xor b;
    layer0_outputs(8992) <= not b or a;
    layer0_outputs(8993) <= not (a xor b);
    layer0_outputs(8994) <= a or b;
    layer0_outputs(8995) <= a;
    layer0_outputs(8996) <= not (a and b);
    layer0_outputs(8997) <= not a;
    layer0_outputs(8998) <= a and not b;
    layer0_outputs(8999) <= a;
    layer0_outputs(9000) <= a or b;
    layer0_outputs(9001) <= not a;
    layer0_outputs(9002) <= not (a xor b);
    layer0_outputs(9003) <= a;
    layer0_outputs(9004) <= not a;
    layer0_outputs(9005) <= a;
    layer0_outputs(9006) <= a and not b;
    layer0_outputs(9007) <= b;
    layer0_outputs(9008) <= a and b;
    layer0_outputs(9009) <= not b;
    layer0_outputs(9010) <= not (a xor b);
    layer0_outputs(9011) <= b;
    layer0_outputs(9012) <= not (a xor b);
    layer0_outputs(9013) <= not b;
    layer0_outputs(9014) <= not (a and b);
    layer0_outputs(9015) <= b and not a;
    layer0_outputs(9016) <= not (a xor b);
    layer0_outputs(9017) <= a and not b;
    layer0_outputs(9018) <= a or b;
    layer0_outputs(9019) <= a;
    layer0_outputs(9020) <= not a;
    layer0_outputs(9021) <= not (a or b);
    layer0_outputs(9022) <= a xor b;
    layer0_outputs(9023) <= a and not b;
    layer0_outputs(9024) <= a and not b;
    layer0_outputs(9025) <= not a;
    layer0_outputs(9026) <= not a;
    layer0_outputs(9027) <= not (a or b);
    layer0_outputs(9028) <= b and not a;
    layer0_outputs(9029) <= a and not b;
    layer0_outputs(9030) <= not a or b;
    layer0_outputs(9031) <= a or b;
    layer0_outputs(9032) <= not b;
    layer0_outputs(9033) <= '1';
    layer0_outputs(9034) <= '0';
    layer0_outputs(9035) <= not b or a;
    layer0_outputs(9036) <= not a;
    layer0_outputs(9037) <= a or b;
    layer0_outputs(9038) <= '0';
    layer0_outputs(9039) <= not a or b;
    layer0_outputs(9040) <= not (a or b);
    layer0_outputs(9041) <= not (a or b);
    layer0_outputs(9042) <= not a or b;
    layer0_outputs(9043) <= b;
    layer0_outputs(9044) <= a xor b;
    layer0_outputs(9045) <= not a or b;
    layer0_outputs(9046) <= not a;
    layer0_outputs(9047) <= b and not a;
    layer0_outputs(9048) <= a xor b;
    layer0_outputs(9049) <= b and not a;
    layer0_outputs(9050) <= a or b;
    layer0_outputs(9051) <= '1';
    layer0_outputs(9052) <= a or b;
    layer0_outputs(9053) <= b;
    layer0_outputs(9054) <= a or b;
    layer0_outputs(9055) <= not a;
    layer0_outputs(9056) <= b and not a;
    layer0_outputs(9057) <= a and b;
    layer0_outputs(9058) <= not b or a;
    layer0_outputs(9059) <= '1';
    layer0_outputs(9060) <= not (a or b);
    layer0_outputs(9061) <= not b;
    layer0_outputs(9062) <= not b or a;
    layer0_outputs(9063) <= not (a and b);
    layer0_outputs(9064) <= a and not b;
    layer0_outputs(9065) <= not b;
    layer0_outputs(9066) <= a xor b;
    layer0_outputs(9067) <= not a or b;
    layer0_outputs(9068) <= '1';
    layer0_outputs(9069) <= not (a xor b);
    layer0_outputs(9070) <= a;
    layer0_outputs(9071) <= a and b;
    layer0_outputs(9072) <= b and not a;
    layer0_outputs(9073) <= not a or b;
    layer0_outputs(9074) <= not (a xor b);
    layer0_outputs(9075) <= a;
    layer0_outputs(9076) <= not (a and b);
    layer0_outputs(9077) <= not (a or b);
    layer0_outputs(9078) <= not b or a;
    layer0_outputs(9079) <= not (a and b);
    layer0_outputs(9080) <= not b;
    layer0_outputs(9081) <= not a;
    layer0_outputs(9082) <= not (a xor b);
    layer0_outputs(9083) <= b;
    layer0_outputs(9084) <= not a;
    layer0_outputs(9085) <= '0';
    layer0_outputs(9086) <= '1';
    layer0_outputs(9087) <= not (a or b);
    layer0_outputs(9088) <= a xor b;
    layer0_outputs(9089) <= not b or a;
    layer0_outputs(9090) <= not b;
    layer0_outputs(9091) <= a and b;
    layer0_outputs(9092) <= not (a or b);
    layer0_outputs(9093) <= a;
    layer0_outputs(9094) <= not b;
    layer0_outputs(9095) <= not b or a;
    layer0_outputs(9096) <= b;
    layer0_outputs(9097) <= b and not a;
    layer0_outputs(9098) <= '1';
    layer0_outputs(9099) <= a;
    layer0_outputs(9100) <= not a or b;
    layer0_outputs(9101) <= not a;
    layer0_outputs(9102) <= a xor b;
    layer0_outputs(9103) <= b;
    layer0_outputs(9104) <= not a or b;
    layer0_outputs(9105) <= '0';
    layer0_outputs(9106) <= not b or a;
    layer0_outputs(9107) <= not a;
    layer0_outputs(9108) <= not b or a;
    layer0_outputs(9109) <= b and not a;
    layer0_outputs(9110) <= a xor b;
    layer0_outputs(9111) <= not b;
    layer0_outputs(9112) <= not (a xor b);
    layer0_outputs(9113) <= b;
    layer0_outputs(9114) <= a and not b;
    layer0_outputs(9115) <= not b or a;
    layer0_outputs(9116) <= a or b;
    layer0_outputs(9117) <= not (a and b);
    layer0_outputs(9118) <= not (a and b);
    layer0_outputs(9119) <= '0';
    layer0_outputs(9120) <= a and not b;
    layer0_outputs(9121) <= a or b;
    layer0_outputs(9122) <= a xor b;
    layer0_outputs(9123) <= a or b;
    layer0_outputs(9124) <= not a;
    layer0_outputs(9125) <= not (a xor b);
    layer0_outputs(9126) <= not (a xor b);
    layer0_outputs(9127) <= not a or b;
    layer0_outputs(9128) <= not b;
    layer0_outputs(9129) <= not a or b;
    layer0_outputs(9130) <= a;
    layer0_outputs(9131) <= a or b;
    layer0_outputs(9132) <= not b or a;
    layer0_outputs(9133) <= b and not a;
    layer0_outputs(9134) <= a or b;
    layer0_outputs(9135) <= b;
    layer0_outputs(9136) <= b;
    layer0_outputs(9137) <= a and b;
    layer0_outputs(9138) <= not a or b;
    layer0_outputs(9139) <= a;
    layer0_outputs(9140) <= a xor b;
    layer0_outputs(9141) <= b and not a;
    layer0_outputs(9142) <= a and not b;
    layer0_outputs(9143) <= not b;
    layer0_outputs(9144) <= not (a or b);
    layer0_outputs(9145) <= a and not b;
    layer0_outputs(9146) <= a and b;
    layer0_outputs(9147) <= not b;
    layer0_outputs(9148) <= b and not a;
    layer0_outputs(9149) <= a and not b;
    layer0_outputs(9150) <= a xor b;
    layer0_outputs(9151) <= not b or a;
    layer0_outputs(9152) <= '1';
    layer0_outputs(9153) <= not a or b;
    layer0_outputs(9154) <= b;
    layer0_outputs(9155) <= a;
    layer0_outputs(9156) <= b;
    layer0_outputs(9157) <= not a;
    layer0_outputs(9158) <= '0';
    layer0_outputs(9159) <= b;
    layer0_outputs(9160) <= a and b;
    layer0_outputs(9161) <= not a;
    layer0_outputs(9162) <= a and not b;
    layer0_outputs(9163) <= not (a or b);
    layer0_outputs(9164) <= not b;
    layer0_outputs(9165) <= a;
    layer0_outputs(9166) <= a and not b;
    layer0_outputs(9167) <= not a or b;
    layer0_outputs(9168) <= a and b;
    layer0_outputs(9169) <= a;
    layer0_outputs(9170) <= a and not b;
    layer0_outputs(9171) <= '0';
    layer0_outputs(9172) <= not (a xor b);
    layer0_outputs(9173) <= a and b;
    layer0_outputs(9174) <= not b or a;
    layer0_outputs(9175) <= not b;
    layer0_outputs(9176) <= not b;
    layer0_outputs(9177) <= not b;
    layer0_outputs(9178) <= a;
    layer0_outputs(9179) <= b;
    layer0_outputs(9180) <= not a or b;
    layer0_outputs(9181) <= b;
    layer0_outputs(9182) <= a;
    layer0_outputs(9183) <= a and b;
    layer0_outputs(9184) <= a;
    layer0_outputs(9185) <= b;
    layer0_outputs(9186) <= not (a xor b);
    layer0_outputs(9187) <= not (a and b);
    layer0_outputs(9188) <= not (a and b);
    layer0_outputs(9189) <= b and not a;
    layer0_outputs(9190) <= a;
    layer0_outputs(9191) <= a xor b;
    layer0_outputs(9192) <= not b or a;
    layer0_outputs(9193) <= not (a xor b);
    layer0_outputs(9194) <= b and not a;
    layer0_outputs(9195) <= not b;
    layer0_outputs(9196) <= a and b;
    layer0_outputs(9197) <= not b;
    layer0_outputs(9198) <= not (a or b);
    layer0_outputs(9199) <= b;
    layer0_outputs(9200) <= a or b;
    layer0_outputs(9201) <= not a or b;
    layer0_outputs(9202) <= not b or a;
    layer0_outputs(9203) <= a and not b;
    layer0_outputs(9204) <= not b;
    layer0_outputs(9205) <= a or b;
    layer0_outputs(9206) <= '1';
    layer0_outputs(9207) <= a xor b;
    layer0_outputs(9208) <= b and not a;
    layer0_outputs(9209) <= a;
    layer0_outputs(9210) <= not (a and b);
    layer0_outputs(9211) <= a;
    layer0_outputs(9212) <= not (a and b);
    layer0_outputs(9213) <= a or b;
    layer0_outputs(9214) <= a and b;
    layer0_outputs(9215) <= a or b;
    layer0_outputs(9216) <= not (a xor b);
    layer0_outputs(9217) <= not b;
    layer0_outputs(9218) <= a;
    layer0_outputs(9219) <= not b;
    layer0_outputs(9220) <= not a;
    layer0_outputs(9221) <= not (a xor b);
    layer0_outputs(9222) <= a;
    layer0_outputs(9223) <= b and not a;
    layer0_outputs(9224) <= a;
    layer0_outputs(9225) <= not (a or b);
    layer0_outputs(9226) <= not a;
    layer0_outputs(9227) <= b;
    layer0_outputs(9228) <= a and not b;
    layer0_outputs(9229) <= not b or a;
    layer0_outputs(9230) <= not a;
    layer0_outputs(9231) <= b;
    layer0_outputs(9232) <= b;
    layer0_outputs(9233) <= a;
    layer0_outputs(9234) <= a and not b;
    layer0_outputs(9235) <= a and b;
    layer0_outputs(9236) <= b;
    layer0_outputs(9237) <= not (a xor b);
    layer0_outputs(9238) <= not b;
    layer0_outputs(9239) <= a and not b;
    layer0_outputs(9240) <= not b;
    layer0_outputs(9241) <= not (a or b);
    layer0_outputs(9242) <= a and not b;
    layer0_outputs(9243) <= a or b;
    layer0_outputs(9244) <= not b or a;
    layer0_outputs(9245) <= not (a xor b);
    layer0_outputs(9246) <= '1';
    layer0_outputs(9247) <= b;
    layer0_outputs(9248) <= b;
    layer0_outputs(9249) <= not a or b;
    layer0_outputs(9250) <= b;
    layer0_outputs(9251) <= not (a or b);
    layer0_outputs(9252) <= not (a and b);
    layer0_outputs(9253) <= '0';
    layer0_outputs(9254) <= '1';
    layer0_outputs(9255) <= '0';
    layer0_outputs(9256) <= a xor b;
    layer0_outputs(9257) <= '1';
    layer0_outputs(9258) <= not a;
    layer0_outputs(9259) <= a and b;
    layer0_outputs(9260) <= a;
    layer0_outputs(9261) <= a xor b;
    layer0_outputs(9262) <= a or b;
    layer0_outputs(9263) <= a;
    layer0_outputs(9264) <= '0';
    layer0_outputs(9265) <= a;
    layer0_outputs(9266) <= not (a or b);
    layer0_outputs(9267) <= b;
    layer0_outputs(9268) <= not b or a;
    layer0_outputs(9269) <= b and not a;
    layer0_outputs(9270) <= not (a xor b);
    layer0_outputs(9271) <= not (a or b);
    layer0_outputs(9272) <= not a or b;
    layer0_outputs(9273) <= a and not b;
    layer0_outputs(9274) <= not a;
    layer0_outputs(9275) <= a;
    layer0_outputs(9276) <= not a or b;
    layer0_outputs(9277) <= not (a and b);
    layer0_outputs(9278) <= not b;
    layer0_outputs(9279) <= a xor b;
    layer0_outputs(9280) <= '0';
    layer0_outputs(9281) <= not a;
    layer0_outputs(9282) <= a and not b;
    layer0_outputs(9283) <= not b or a;
    layer0_outputs(9284) <= not b;
    layer0_outputs(9285) <= a and b;
    layer0_outputs(9286) <= b;
    layer0_outputs(9287) <= not (a and b);
    layer0_outputs(9288) <= b and not a;
    layer0_outputs(9289) <= not (a xor b);
    layer0_outputs(9290) <= not (a or b);
    layer0_outputs(9291) <= not a;
    layer0_outputs(9292) <= not a;
    layer0_outputs(9293) <= not b;
    layer0_outputs(9294) <= not (a xor b);
    layer0_outputs(9295) <= not b or a;
    layer0_outputs(9296) <= a xor b;
    layer0_outputs(9297) <= '1';
    layer0_outputs(9298) <= not (a and b);
    layer0_outputs(9299) <= a and not b;
    layer0_outputs(9300) <= a and not b;
    layer0_outputs(9301) <= not b or a;
    layer0_outputs(9302) <= not a or b;
    layer0_outputs(9303) <= not (a or b);
    layer0_outputs(9304) <= not (a or b);
    layer0_outputs(9305) <= a or b;
    layer0_outputs(9306) <= b;
    layer0_outputs(9307) <= not a;
    layer0_outputs(9308) <= not a or b;
    layer0_outputs(9309) <= a;
    layer0_outputs(9310) <= '0';
    layer0_outputs(9311) <= a and not b;
    layer0_outputs(9312) <= a xor b;
    layer0_outputs(9313) <= not a or b;
    layer0_outputs(9314) <= not (a or b);
    layer0_outputs(9315) <= not b or a;
    layer0_outputs(9316) <= b and not a;
    layer0_outputs(9317) <= b and not a;
    layer0_outputs(9318) <= not (a or b);
    layer0_outputs(9319) <= a and b;
    layer0_outputs(9320) <= a xor b;
    layer0_outputs(9321) <= not b or a;
    layer0_outputs(9322) <= not (a or b);
    layer0_outputs(9323) <= '0';
    layer0_outputs(9324) <= '0';
    layer0_outputs(9325) <= b;
    layer0_outputs(9326) <= not a or b;
    layer0_outputs(9327) <= a and b;
    layer0_outputs(9328) <= a or b;
    layer0_outputs(9329) <= a;
    layer0_outputs(9330) <= a xor b;
    layer0_outputs(9331) <= a or b;
    layer0_outputs(9332) <= '0';
    layer0_outputs(9333) <= not (a xor b);
    layer0_outputs(9334) <= not b or a;
    layer0_outputs(9335) <= a and not b;
    layer0_outputs(9336) <= not (a xor b);
    layer0_outputs(9337) <= not b or a;
    layer0_outputs(9338) <= not (a xor b);
    layer0_outputs(9339) <= not (a or b);
    layer0_outputs(9340) <= a and not b;
    layer0_outputs(9341) <= not (a or b);
    layer0_outputs(9342) <= not a or b;
    layer0_outputs(9343) <= not b;
    layer0_outputs(9344) <= a and not b;
    layer0_outputs(9345) <= not b or a;
    layer0_outputs(9346) <= a and b;
    layer0_outputs(9347) <= a or b;
    layer0_outputs(9348) <= not b or a;
    layer0_outputs(9349) <= not b;
    layer0_outputs(9350) <= not b;
    layer0_outputs(9351) <= not a or b;
    layer0_outputs(9352) <= not (a xor b);
    layer0_outputs(9353) <= b and not a;
    layer0_outputs(9354) <= a xor b;
    layer0_outputs(9355) <= b;
    layer0_outputs(9356) <= a xor b;
    layer0_outputs(9357) <= not (a xor b);
    layer0_outputs(9358) <= not (a xor b);
    layer0_outputs(9359) <= a or b;
    layer0_outputs(9360) <= not b or a;
    layer0_outputs(9361) <= '0';
    layer0_outputs(9362) <= b;
    layer0_outputs(9363) <= a and not b;
    layer0_outputs(9364) <= b;
    layer0_outputs(9365) <= not (a or b);
    layer0_outputs(9366) <= a or b;
    layer0_outputs(9367) <= a and not b;
    layer0_outputs(9368) <= '1';
    layer0_outputs(9369) <= a;
    layer0_outputs(9370) <= not (a xor b);
    layer0_outputs(9371) <= a and not b;
    layer0_outputs(9372) <= not b;
    layer0_outputs(9373) <= a and not b;
    layer0_outputs(9374) <= a or b;
    layer0_outputs(9375) <= a and not b;
    layer0_outputs(9376) <= not b or a;
    layer0_outputs(9377) <= not a or b;
    layer0_outputs(9378) <= a xor b;
    layer0_outputs(9379) <= '1';
    layer0_outputs(9380) <= a and not b;
    layer0_outputs(9381) <= not (a or b);
    layer0_outputs(9382) <= a;
    layer0_outputs(9383) <= a and not b;
    layer0_outputs(9384) <= '0';
    layer0_outputs(9385) <= a and b;
    layer0_outputs(9386) <= not a;
    layer0_outputs(9387) <= not a;
    layer0_outputs(9388) <= not (a or b);
    layer0_outputs(9389) <= '1';
    layer0_outputs(9390) <= not (a or b);
    layer0_outputs(9391) <= b;
    layer0_outputs(9392) <= not a;
    layer0_outputs(9393) <= not b;
    layer0_outputs(9394) <= a xor b;
    layer0_outputs(9395) <= a or b;
    layer0_outputs(9396) <= a or b;
    layer0_outputs(9397) <= not a;
    layer0_outputs(9398) <= a xor b;
    layer0_outputs(9399) <= a and not b;
    layer0_outputs(9400) <= not (a or b);
    layer0_outputs(9401) <= not a;
    layer0_outputs(9402) <= a and b;
    layer0_outputs(9403) <= b;
    layer0_outputs(9404) <= b;
    layer0_outputs(9405) <= b and not a;
    layer0_outputs(9406) <= not a or b;
    layer0_outputs(9407) <= not b;
    layer0_outputs(9408) <= '0';
    layer0_outputs(9409) <= a xor b;
    layer0_outputs(9410) <= a xor b;
    layer0_outputs(9411) <= '1';
    layer0_outputs(9412) <= a;
    layer0_outputs(9413) <= '0';
    layer0_outputs(9414) <= a and b;
    layer0_outputs(9415) <= not b;
    layer0_outputs(9416) <= not b or a;
    layer0_outputs(9417) <= not a;
    layer0_outputs(9418) <= not b or a;
    layer0_outputs(9419) <= not a;
    layer0_outputs(9420) <= not (a and b);
    layer0_outputs(9421) <= not b;
    layer0_outputs(9422) <= not (a or b);
    layer0_outputs(9423) <= not b;
    layer0_outputs(9424) <= a and not b;
    layer0_outputs(9425) <= not (a or b);
    layer0_outputs(9426) <= a or b;
    layer0_outputs(9427) <= not a;
    layer0_outputs(9428) <= not a or b;
    layer0_outputs(9429) <= b;
    layer0_outputs(9430) <= b and not a;
    layer0_outputs(9431) <= not (a xor b);
    layer0_outputs(9432) <= a xor b;
    layer0_outputs(9433) <= a and not b;
    layer0_outputs(9434) <= not b or a;
    layer0_outputs(9435) <= not b;
    layer0_outputs(9436) <= a;
    layer0_outputs(9437) <= a and b;
    layer0_outputs(9438) <= not (a xor b);
    layer0_outputs(9439) <= a;
    layer0_outputs(9440) <= not a or b;
    layer0_outputs(9441) <= a or b;
    layer0_outputs(9442) <= not (a and b);
    layer0_outputs(9443) <= not (a or b);
    layer0_outputs(9444) <= not (a or b);
    layer0_outputs(9445) <= b and not a;
    layer0_outputs(9446) <= not a or b;
    layer0_outputs(9447) <= a xor b;
    layer0_outputs(9448) <= a or b;
    layer0_outputs(9449) <= not b;
    layer0_outputs(9450) <= not (a xor b);
    layer0_outputs(9451) <= not (a xor b);
    layer0_outputs(9452) <= not (a or b);
    layer0_outputs(9453) <= not (a and b);
    layer0_outputs(9454) <= a xor b;
    layer0_outputs(9455) <= b and not a;
    layer0_outputs(9456) <= a or b;
    layer0_outputs(9457) <= not (a xor b);
    layer0_outputs(9458) <= not a or b;
    layer0_outputs(9459) <= b;
    layer0_outputs(9460) <= a;
    layer0_outputs(9461) <= '1';
    layer0_outputs(9462) <= not b or a;
    layer0_outputs(9463) <= not b;
    layer0_outputs(9464) <= not (a xor b);
    layer0_outputs(9465) <= b;
    layer0_outputs(9466) <= a and not b;
    layer0_outputs(9467) <= a or b;
    layer0_outputs(9468) <= a or b;
    layer0_outputs(9469) <= not (a xor b);
    layer0_outputs(9470) <= not a;
    layer0_outputs(9471) <= not b;
    layer0_outputs(9472) <= not (a and b);
    layer0_outputs(9473) <= not (a or b);
    layer0_outputs(9474) <= b;
    layer0_outputs(9475) <= b;
    layer0_outputs(9476) <= not b;
    layer0_outputs(9477) <= not b;
    layer0_outputs(9478) <= a or b;
    layer0_outputs(9479) <= a xor b;
    layer0_outputs(9480) <= not (a and b);
    layer0_outputs(9481) <= not b;
    layer0_outputs(9482) <= '0';
    layer0_outputs(9483) <= not b;
    layer0_outputs(9484) <= not (a or b);
    layer0_outputs(9485) <= not (a or b);
    layer0_outputs(9486) <= not b;
    layer0_outputs(9487) <= not a or b;
    layer0_outputs(9488) <= not a or b;
    layer0_outputs(9489) <= '1';
    layer0_outputs(9490) <= a and b;
    layer0_outputs(9491) <= a or b;
    layer0_outputs(9492) <= a or b;
    layer0_outputs(9493) <= '0';
    layer0_outputs(9494) <= not (a xor b);
    layer0_outputs(9495) <= not a;
    layer0_outputs(9496) <= not a;
    layer0_outputs(9497) <= b and not a;
    layer0_outputs(9498) <= b;
    layer0_outputs(9499) <= not a;
    layer0_outputs(9500) <= not a;
    layer0_outputs(9501) <= a or b;
    layer0_outputs(9502) <= not (a or b);
    layer0_outputs(9503) <= not b or a;
    layer0_outputs(9504) <= not (a xor b);
    layer0_outputs(9505) <= a and not b;
    layer0_outputs(9506) <= not a or b;
    layer0_outputs(9507) <= a xor b;
    layer0_outputs(9508) <= not (a or b);
    layer0_outputs(9509) <= a or b;
    layer0_outputs(9510) <= not a or b;
    layer0_outputs(9511) <= not (a or b);
    layer0_outputs(9512) <= b and not a;
    layer0_outputs(9513) <= not (a or b);
    layer0_outputs(9514) <= b and not a;
    layer0_outputs(9515) <= not (a and b);
    layer0_outputs(9516) <= a or b;
    layer0_outputs(9517) <= a xor b;
    layer0_outputs(9518) <= b;
    layer0_outputs(9519) <= a xor b;
    layer0_outputs(9520) <= not (a and b);
    layer0_outputs(9521) <= not b or a;
    layer0_outputs(9522) <= not (a xor b);
    layer0_outputs(9523) <= not b or a;
    layer0_outputs(9524) <= b;
    layer0_outputs(9525) <= '1';
    layer0_outputs(9526) <= a and b;
    layer0_outputs(9527) <= '0';
    layer0_outputs(9528) <= not b or a;
    layer0_outputs(9529) <= not (a xor b);
    layer0_outputs(9530) <= not b or a;
    layer0_outputs(9531) <= not (a or b);
    layer0_outputs(9532) <= not (a and b);
    layer0_outputs(9533) <= b;
    layer0_outputs(9534) <= not b;
    layer0_outputs(9535) <= not (a xor b);
    layer0_outputs(9536) <= not a;
    layer0_outputs(9537) <= not b or a;
    layer0_outputs(9538) <= b;
    layer0_outputs(9539) <= not (a xor b);
    layer0_outputs(9540) <= not b;
    layer0_outputs(9541) <= a;
    layer0_outputs(9542) <= a;
    layer0_outputs(9543) <= '1';
    layer0_outputs(9544) <= a xor b;
    layer0_outputs(9545) <= not a;
    layer0_outputs(9546) <= a and b;
    layer0_outputs(9547) <= b;
    layer0_outputs(9548) <= b and not a;
    layer0_outputs(9549) <= '0';
    layer0_outputs(9550) <= not b or a;
    layer0_outputs(9551) <= not a;
    layer0_outputs(9552) <= not a or b;
    layer0_outputs(9553) <= not (a xor b);
    layer0_outputs(9554) <= a and not b;
    layer0_outputs(9555) <= a or b;
    layer0_outputs(9556) <= '0';
    layer0_outputs(9557) <= not (a xor b);
    layer0_outputs(9558) <= not (a or b);
    layer0_outputs(9559) <= not a or b;
    layer0_outputs(9560) <= a;
    layer0_outputs(9561) <= b;
    layer0_outputs(9562) <= not a or b;
    layer0_outputs(9563) <= not (a xor b);
    layer0_outputs(9564) <= a and not b;
    layer0_outputs(9565) <= '1';
    layer0_outputs(9566) <= b;
    layer0_outputs(9567) <= a;
    layer0_outputs(9568) <= not b;
    layer0_outputs(9569) <= a xor b;
    layer0_outputs(9570) <= b and not a;
    layer0_outputs(9571) <= not b;
    layer0_outputs(9572) <= not (a or b);
    layer0_outputs(9573) <= b and not a;
    layer0_outputs(9574) <= '1';
    layer0_outputs(9575) <= a and b;
    layer0_outputs(9576) <= '0';
    layer0_outputs(9577) <= not a or b;
    layer0_outputs(9578) <= not (a and b);
    layer0_outputs(9579) <= b and not a;
    layer0_outputs(9580) <= not b;
    layer0_outputs(9581) <= a and b;
    layer0_outputs(9582) <= not (a or b);
    layer0_outputs(9583) <= a or b;
    layer0_outputs(9584) <= a and not b;
    layer0_outputs(9585) <= a and not b;
    layer0_outputs(9586) <= not (a or b);
    layer0_outputs(9587) <= not a;
    layer0_outputs(9588) <= '0';
    layer0_outputs(9589) <= not b;
    layer0_outputs(9590) <= not a or b;
    layer0_outputs(9591) <= not a or b;
    layer0_outputs(9592) <= a and b;
    layer0_outputs(9593) <= a or b;
    layer0_outputs(9594) <= a and b;
    layer0_outputs(9595) <= not b or a;
    layer0_outputs(9596) <= not (a or b);
    layer0_outputs(9597) <= not b;
    layer0_outputs(9598) <= '1';
    layer0_outputs(9599) <= a;
    layer0_outputs(9600) <= a or b;
    layer0_outputs(9601) <= a or b;
    layer0_outputs(9602) <= a;
    layer0_outputs(9603) <= not (a and b);
    layer0_outputs(9604) <= not b or a;
    layer0_outputs(9605) <= not (a xor b);
    layer0_outputs(9606) <= a xor b;
    layer0_outputs(9607) <= '1';
    layer0_outputs(9608) <= a and b;
    layer0_outputs(9609) <= not b;
    layer0_outputs(9610) <= '0';
    layer0_outputs(9611) <= a xor b;
    layer0_outputs(9612) <= not b or a;
    layer0_outputs(9613) <= not b or a;
    layer0_outputs(9614) <= a xor b;
    layer0_outputs(9615) <= not b or a;
    layer0_outputs(9616) <= not (a xor b);
    layer0_outputs(9617) <= not (a xor b);
    layer0_outputs(9618) <= not a;
    layer0_outputs(9619) <= b and not a;
    layer0_outputs(9620) <= a or b;
    layer0_outputs(9621) <= a or b;
    layer0_outputs(9622) <= not (a xor b);
    layer0_outputs(9623) <= '1';
    layer0_outputs(9624) <= a xor b;
    layer0_outputs(9625) <= a and not b;
    layer0_outputs(9626) <= b and not a;
    layer0_outputs(9627) <= b and not a;
    layer0_outputs(9628) <= a or b;
    layer0_outputs(9629) <= not (a and b);
    layer0_outputs(9630) <= not (a or b);
    layer0_outputs(9631) <= not (a or b);
    layer0_outputs(9632) <= a and not b;
    layer0_outputs(9633) <= a or b;
    layer0_outputs(9634) <= not a;
    layer0_outputs(9635) <= a;
    layer0_outputs(9636) <= '0';
    layer0_outputs(9637) <= '0';
    layer0_outputs(9638) <= a;
    layer0_outputs(9639) <= b;
    layer0_outputs(9640) <= b and not a;
    layer0_outputs(9641) <= not (a or b);
    layer0_outputs(9642) <= b and not a;
    layer0_outputs(9643) <= not b;
    layer0_outputs(9644) <= '1';
    layer0_outputs(9645) <= not a;
    layer0_outputs(9646) <= not b;
    layer0_outputs(9647) <= not (a or b);
    layer0_outputs(9648) <= '1';
    layer0_outputs(9649) <= a and b;
    layer0_outputs(9650) <= b;
    layer0_outputs(9651) <= a xor b;
    layer0_outputs(9652) <= not b or a;
    layer0_outputs(9653) <= not (a or b);
    layer0_outputs(9654) <= a or b;
    layer0_outputs(9655) <= a xor b;
    layer0_outputs(9656) <= a or b;
    layer0_outputs(9657) <= not b;
    layer0_outputs(9658) <= not b or a;
    layer0_outputs(9659) <= not b or a;
    layer0_outputs(9660) <= not b;
    layer0_outputs(9661) <= not (a and b);
    layer0_outputs(9662) <= not a;
    layer0_outputs(9663) <= '0';
    layer0_outputs(9664) <= not (a or b);
    layer0_outputs(9665) <= not (a and b);
    layer0_outputs(9666) <= not (a xor b);
    layer0_outputs(9667) <= not a;
    layer0_outputs(9668) <= a;
    layer0_outputs(9669) <= '0';
    layer0_outputs(9670) <= a;
    layer0_outputs(9671) <= b and not a;
    layer0_outputs(9672) <= a or b;
    layer0_outputs(9673) <= not (a or b);
    layer0_outputs(9674) <= b and not a;
    layer0_outputs(9675) <= a and not b;
    layer0_outputs(9676) <= not (a or b);
    layer0_outputs(9677) <= a xor b;
    layer0_outputs(9678) <= not (a or b);
    layer0_outputs(9679) <= '1';
    layer0_outputs(9680) <= a and b;
    layer0_outputs(9681) <= a;
    layer0_outputs(9682) <= a;
    layer0_outputs(9683) <= b;
    layer0_outputs(9684) <= a;
    layer0_outputs(9685) <= not a;
    layer0_outputs(9686) <= a and b;
    layer0_outputs(9687) <= '0';
    layer0_outputs(9688) <= a and not b;
    layer0_outputs(9689) <= a;
    layer0_outputs(9690) <= not a;
    layer0_outputs(9691) <= '0';
    layer0_outputs(9692) <= not a;
    layer0_outputs(9693) <= not b;
    layer0_outputs(9694) <= not b;
    layer0_outputs(9695) <= a xor b;
    layer0_outputs(9696) <= b and not a;
    layer0_outputs(9697) <= not (a and b);
    layer0_outputs(9698) <= a and b;
    layer0_outputs(9699) <= a and not b;
    layer0_outputs(9700) <= '0';
    layer0_outputs(9701) <= a or b;
    layer0_outputs(9702) <= b;
    layer0_outputs(9703) <= not a;
    layer0_outputs(9704) <= a or b;
    layer0_outputs(9705) <= not b;
    layer0_outputs(9706) <= a xor b;
    layer0_outputs(9707) <= not (a and b);
    layer0_outputs(9708) <= b;
    layer0_outputs(9709) <= a;
    layer0_outputs(9710) <= a and not b;
    layer0_outputs(9711) <= not a;
    layer0_outputs(9712) <= not b;
    layer0_outputs(9713) <= b;
    layer0_outputs(9714) <= a or b;
    layer0_outputs(9715) <= not a;
    layer0_outputs(9716) <= a and not b;
    layer0_outputs(9717) <= '0';
    layer0_outputs(9718) <= not (a and b);
    layer0_outputs(9719) <= not a or b;
    layer0_outputs(9720) <= not b or a;
    layer0_outputs(9721) <= a;
    layer0_outputs(9722) <= a;
    layer0_outputs(9723) <= b and not a;
    layer0_outputs(9724) <= '0';
    layer0_outputs(9725) <= not (a or b);
    layer0_outputs(9726) <= not a or b;
    layer0_outputs(9727) <= b;
    layer0_outputs(9728) <= b and not a;
    layer0_outputs(9729) <= a and not b;
    layer0_outputs(9730) <= b;
    layer0_outputs(9731) <= b;
    layer0_outputs(9732) <= b;
    layer0_outputs(9733) <= b;
    layer0_outputs(9734) <= b;
    layer0_outputs(9735) <= a or b;
    layer0_outputs(9736) <= not (a or b);
    layer0_outputs(9737) <= a xor b;
    layer0_outputs(9738) <= not b;
    layer0_outputs(9739) <= not (a xor b);
    layer0_outputs(9740) <= a xor b;
    layer0_outputs(9741) <= not (a or b);
    layer0_outputs(9742) <= not (a xor b);
    layer0_outputs(9743) <= not a or b;
    layer0_outputs(9744) <= a or b;
    layer0_outputs(9745) <= a xor b;
    layer0_outputs(9746) <= a;
    layer0_outputs(9747) <= a or b;
    layer0_outputs(9748) <= a;
    layer0_outputs(9749) <= b;
    layer0_outputs(9750) <= b;
    layer0_outputs(9751) <= '0';
    layer0_outputs(9752) <= not a or b;
    layer0_outputs(9753) <= not a or b;
    layer0_outputs(9754) <= '1';
    layer0_outputs(9755) <= not (a xor b);
    layer0_outputs(9756) <= a and b;
    layer0_outputs(9757) <= a or b;
    layer0_outputs(9758) <= a xor b;
    layer0_outputs(9759) <= a and not b;
    layer0_outputs(9760) <= a;
    layer0_outputs(9761) <= a or b;
    layer0_outputs(9762) <= a and b;
    layer0_outputs(9763) <= a xor b;
    layer0_outputs(9764) <= a;
    layer0_outputs(9765) <= not a or b;
    layer0_outputs(9766) <= not (a and b);
    layer0_outputs(9767) <= not (a or b);
    layer0_outputs(9768) <= not (a xor b);
    layer0_outputs(9769) <= not a;
    layer0_outputs(9770) <= a;
    layer0_outputs(9771) <= not a;
    layer0_outputs(9772) <= not a or b;
    layer0_outputs(9773) <= a;
    layer0_outputs(9774) <= b and not a;
    layer0_outputs(9775) <= not (a or b);
    layer0_outputs(9776) <= a;
    layer0_outputs(9777) <= a or b;
    layer0_outputs(9778) <= b;
    layer0_outputs(9779) <= a;
    layer0_outputs(9780) <= a or b;
    layer0_outputs(9781) <= not b;
    layer0_outputs(9782) <= a and not b;
    layer0_outputs(9783) <= a and b;
    layer0_outputs(9784) <= a or b;
    layer0_outputs(9785) <= '0';
    layer0_outputs(9786) <= not (a or b);
    layer0_outputs(9787) <= b;
    layer0_outputs(9788) <= not (a xor b);
    layer0_outputs(9789) <= '1';
    layer0_outputs(9790) <= not a or b;
    layer0_outputs(9791) <= b and not a;
    layer0_outputs(9792) <= not (a or b);
    layer0_outputs(9793) <= a xor b;
    layer0_outputs(9794) <= a or b;
    layer0_outputs(9795) <= not (a or b);
    layer0_outputs(9796) <= not (a or b);
    layer0_outputs(9797) <= not (a and b);
    layer0_outputs(9798) <= b;
    layer0_outputs(9799) <= not (a and b);
    layer0_outputs(9800) <= a or b;
    layer0_outputs(9801) <= '0';
    layer0_outputs(9802) <= b;
    layer0_outputs(9803) <= b and not a;
    layer0_outputs(9804) <= not (a xor b);
    layer0_outputs(9805) <= not a;
    layer0_outputs(9806) <= a and b;
    layer0_outputs(9807) <= '1';
    layer0_outputs(9808) <= not b or a;
    layer0_outputs(9809) <= a;
    layer0_outputs(9810) <= not (a or b);
    layer0_outputs(9811) <= a;
    layer0_outputs(9812) <= b;
    layer0_outputs(9813) <= a or b;
    layer0_outputs(9814) <= not (a or b);
    layer0_outputs(9815) <= a xor b;
    layer0_outputs(9816) <= not (a and b);
    layer0_outputs(9817) <= b;
    layer0_outputs(9818) <= a or b;
    layer0_outputs(9819) <= '0';
    layer0_outputs(9820) <= not (a xor b);
    layer0_outputs(9821) <= a and b;
    layer0_outputs(9822) <= b and not a;
    layer0_outputs(9823) <= not b or a;
    layer0_outputs(9824) <= '0';
    layer0_outputs(9825) <= not (a xor b);
    layer0_outputs(9826) <= not b;
    layer0_outputs(9827) <= not a or b;
    layer0_outputs(9828) <= b;
    layer0_outputs(9829) <= b and not a;
    layer0_outputs(9830) <= b;
    layer0_outputs(9831) <= a and not b;
    layer0_outputs(9832) <= not (a or b);
    layer0_outputs(9833) <= b;
    layer0_outputs(9834) <= not (a xor b);
    layer0_outputs(9835) <= not (a or b);
    layer0_outputs(9836) <= a or b;
    layer0_outputs(9837) <= a or b;
    layer0_outputs(9838) <= b and not a;
    layer0_outputs(9839) <= not b or a;
    layer0_outputs(9840) <= not b;
    layer0_outputs(9841) <= a or b;
    layer0_outputs(9842) <= a and not b;
    layer0_outputs(9843) <= not b;
    layer0_outputs(9844) <= a or b;
    layer0_outputs(9845) <= not b or a;
    layer0_outputs(9846) <= a xor b;
    layer0_outputs(9847) <= not (a or b);
    layer0_outputs(9848) <= not (a or b);
    layer0_outputs(9849) <= not (a and b);
    layer0_outputs(9850) <= a;
    layer0_outputs(9851) <= b;
    layer0_outputs(9852) <= not (a and b);
    layer0_outputs(9853) <= b;
    layer0_outputs(9854) <= not a;
    layer0_outputs(9855) <= not b or a;
    layer0_outputs(9856) <= b and not a;
    layer0_outputs(9857) <= not a or b;
    layer0_outputs(9858) <= not (a and b);
    layer0_outputs(9859) <= a and b;
    layer0_outputs(9860) <= '0';
    layer0_outputs(9861) <= not a or b;
    layer0_outputs(9862) <= not b or a;
    layer0_outputs(9863) <= not b or a;
    layer0_outputs(9864) <= not a;
    layer0_outputs(9865) <= a or b;
    layer0_outputs(9866) <= a and not b;
    layer0_outputs(9867) <= not b or a;
    layer0_outputs(9868) <= not (a or b);
    layer0_outputs(9869) <= not (a or b);
    layer0_outputs(9870) <= not a or b;
    layer0_outputs(9871) <= not b;
    layer0_outputs(9872) <= not b;
    layer0_outputs(9873) <= not b;
    layer0_outputs(9874) <= a or b;
    layer0_outputs(9875) <= a;
    layer0_outputs(9876) <= not (a or b);
    layer0_outputs(9877) <= not (a xor b);
    layer0_outputs(9878) <= b;
    layer0_outputs(9879) <= a and not b;
    layer0_outputs(9880) <= not (a xor b);
    layer0_outputs(9881) <= not (a xor b);
    layer0_outputs(9882) <= a and not b;
    layer0_outputs(9883) <= not b;
    layer0_outputs(9884) <= '0';
    layer0_outputs(9885) <= b and not a;
    layer0_outputs(9886) <= '0';
    layer0_outputs(9887) <= not (a xor b);
    layer0_outputs(9888) <= not (a xor b);
    layer0_outputs(9889) <= a and not b;
    layer0_outputs(9890) <= not b;
    layer0_outputs(9891) <= '1';
    layer0_outputs(9892) <= a and not b;
    layer0_outputs(9893) <= '1';
    layer0_outputs(9894) <= not b or a;
    layer0_outputs(9895) <= '0';
    layer0_outputs(9896) <= a and not b;
    layer0_outputs(9897) <= not a or b;
    layer0_outputs(9898) <= a and not b;
    layer0_outputs(9899) <= b;
    layer0_outputs(9900) <= a;
    layer0_outputs(9901) <= not a;
    layer0_outputs(9902) <= not (a and b);
    layer0_outputs(9903) <= not b;
    layer0_outputs(9904) <= a;
    layer0_outputs(9905) <= a xor b;
    layer0_outputs(9906) <= not a or b;
    layer0_outputs(9907) <= a or b;
    layer0_outputs(9908) <= not (a or b);
    layer0_outputs(9909) <= a and not b;
    layer0_outputs(9910) <= not (a and b);
    layer0_outputs(9911) <= not (a and b);
    layer0_outputs(9912) <= a and not b;
    layer0_outputs(9913) <= b;
    layer0_outputs(9914) <= a;
    layer0_outputs(9915) <= b and not a;
    layer0_outputs(9916) <= not (a xor b);
    layer0_outputs(9917) <= not a;
    layer0_outputs(9918) <= b;
    layer0_outputs(9919) <= not (a or b);
    layer0_outputs(9920) <= not b or a;
    layer0_outputs(9921) <= b;
    layer0_outputs(9922) <= not (a or b);
    layer0_outputs(9923) <= not (a or b);
    layer0_outputs(9924) <= not a or b;
    layer0_outputs(9925) <= not a;
    layer0_outputs(9926) <= a;
    layer0_outputs(9927) <= a;
    layer0_outputs(9928) <= a;
    layer0_outputs(9929) <= a and not b;
    layer0_outputs(9930) <= not (a xor b);
    layer0_outputs(9931) <= a or b;
    layer0_outputs(9932) <= not b or a;
    layer0_outputs(9933) <= a and not b;
    layer0_outputs(9934) <= not (a and b);
    layer0_outputs(9935) <= b and not a;
    layer0_outputs(9936) <= not b;
    layer0_outputs(9937) <= b;
    layer0_outputs(9938) <= a or b;
    layer0_outputs(9939) <= not a;
    layer0_outputs(9940) <= not (a and b);
    layer0_outputs(9941) <= a and not b;
    layer0_outputs(9942) <= b and not a;
    layer0_outputs(9943) <= not b;
    layer0_outputs(9944) <= not (a and b);
    layer0_outputs(9945) <= b and not a;
    layer0_outputs(9946) <= not (a and b);
    layer0_outputs(9947) <= not b or a;
    layer0_outputs(9948) <= not (a xor b);
    layer0_outputs(9949) <= '0';
    layer0_outputs(9950) <= not b or a;
    layer0_outputs(9951) <= not (a and b);
    layer0_outputs(9952) <= a xor b;
    layer0_outputs(9953) <= not b or a;
    layer0_outputs(9954) <= not a;
    layer0_outputs(9955) <= not a or b;
    layer0_outputs(9956) <= '0';
    layer0_outputs(9957) <= a and not b;
    layer0_outputs(9958) <= b and not a;
    layer0_outputs(9959) <= a or b;
    layer0_outputs(9960) <= '1';
    layer0_outputs(9961) <= not (a and b);
    layer0_outputs(9962) <= a and not b;
    layer0_outputs(9963) <= a and not b;
    layer0_outputs(9964) <= not (a xor b);
    layer0_outputs(9965) <= '0';
    layer0_outputs(9966) <= b and not a;
    layer0_outputs(9967) <= a or b;
    layer0_outputs(9968) <= not a or b;
    layer0_outputs(9969) <= not (a xor b);
    layer0_outputs(9970) <= not a;
    layer0_outputs(9971) <= a and not b;
    layer0_outputs(9972) <= a and not b;
    layer0_outputs(9973) <= a;
    layer0_outputs(9974) <= '0';
    layer0_outputs(9975) <= a or b;
    layer0_outputs(9976) <= not (a and b);
    layer0_outputs(9977) <= a and b;
    layer0_outputs(9978) <= a;
    layer0_outputs(9979) <= a and not b;
    layer0_outputs(9980) <= a or b;
    layer0_outputs(9981) <= '1';
    layer0_outputs(9982) <= not a or b;
    layer0_outputs(9983) <= a or b;
    layer0_outputs(9984) <= a and b;
    layer0_outputs(9985) <= not a or b;
    layer0_outputs(9986) <= not b or a;
    layer0_outputs(9987) <= '0';
    layer0_outputs(9988) <= not b or a;
    layer0_outputs(9989) <= b;
    layer0_outputs(9990) <= not (a or b);
    layer0_outputs(9991) <= a;
    layer0_outputs(9992) <= a and not b;
    layer0_outputs(9993) <= not a or b;
    layer0_outputs(9994) <= not a;
    layer0_outputs(9995) <= not a;
    layer0_outputs(9996) <= a or b;
    layer0_outputs(9997) <= not a;
    layer0_outputs(9998) <= a or b;
    layer0_outputs(9999) <= '1';
    layer0_outputs(10000) <= not (a or b);
    layer0_outputs(10001) <= b and not a;
    layer0_outputs(10002) <= b;
    layer0_outputs(10003) <= a and b;
    layer0_outputs(10004) <= not a;
    layer0_outputs(10005) <= not (a or b);
    layer0_outputs(10006) <= not b;
    layer0_outputs(10007) <= not a or b;
    layer0_outputs(10008) <= not (a and b);
    layer0_outputs(10009) <= not (a and b);
    layer0_outputs(10010) <= a;
    layer0_outputs(10011) <= a and b;
    layer0_outputs(10012) <= not (a and b);
    layer0_outputs(10013) <= a and b;
    layer0_outputs(10014) <= not b;
    layer0_outputs(10015) <= not b;
    layer0_outputs(10016) <= a xor b;
    layer0_outputs(10017) <= a and not b;
    layer0_outputs(10018) <= a;
    layer0_outputs(10019) <= a xor b;
    layer0_outputs(10020) <= not (a or b);
    layer0_outputs(10021) <= '1';
    layer0_outputs(10022) <= not b;
    layer0_outputs(10023) <= b;
    layer0_outputs(10024) <= a or b;
    layer0_outputs(10025) <= not a or b;
    layer0_outputs(10026) <= not (a and b);
    layer0_outputs(10027) <= a;
    layer0_outputs(10028) <= b and not a;
    layer0_outputs(10029) <= not b or a;
    layer0_outputs(10030) <= '0';
    layer0_outputs(10031) <= not a or b;
    layer0_outputs(10032) <= b and not a;
    layer0_outputs(10033) <= not b;
    layer0_outputs(10034) <= a;
    layer0_outputs(10035) <= a xor b;
    layer0_outputs(10036) <= b and not a;
    layer0_outputs(10037) <= not b;
    layer0_outputs(10038) <= not (a and b);
    layer0_outputs(10039) <= b and not a;
    layer0_outputs(10040) <= a;
    layer0_outputs(10041) <= not b;
    layer0_outputs(10042) <= a and b;
    layer0_outputs(10043) <= not a or b;
    layer0_outputs(10044) <= not (a xor b);
    layer0_outputs(10045) <= not a;
    layer0_outputs(10046) <= not a;
    layer0_outputs(10047) <= not a or b;
    layer0_outputs(10048) <= '1';
    layer0_outputs(10049) <= b and not a;
    layer0_outputs(10050) <= not b or a;
    layer0_outputs(10051) <= not b;
    layer0_outputs(10052) <= a or b;
    layer0_outputs(10053) <= b;
    layer0_outputs(10054) <= not (a and b);
    layer0_outputs(10055) <= b;
    layer0_outputs(10056) <= b;
    layer0_outputs(10057) <= a and not b;
    layer0_outputs(10058) <= not (a xor b);
    layer0_outputs(10059) <= '0';
    layer0_outputs(10060) <= not b;
    layer0_outputs(10061) <= '1';
    layer0_outputs(10062) <= '1';
    layer0_outputs(10063) <= b;
    layer0_outputs(10064) <= b;
    layer0_outputs(10065) <= b;
    layer0_outputs(10066) <= a;
    layer0_outputs(10067) <= not b or a;
    layer0_outputs(10068) <= a and b;
    layer0_outputs(10069) <= not b or a;
    layer0_outputs(10070) <= not (a and b);
    layer0_outputs(10071) <= '1';
    layer0_outputs(10072) <= b;
    layer0_outputs(10073) <= not a;
    layer0_outputs(10074) <= '0';
    layer0_outputs(10075) <= not a;
    layer0_outputs(10076) <= a;
    layer0_outputs(10077) <= '1';
    layer0_outputs(10078) <= not b;
    layer0_outputs(10079) <= a;
    layer0_outputs(10080) <= not b or a;
    layer0_outputs(10081) <= '1';
    layer0_outputs(10082) <= a or b;
    layer0_outputs(10083) <= a xor b;
    layer0_outputs(10084) <= not (a and b);
    layer0_outputs(10085) <= not a;
    layer0_outputs(10086) <= not b;
    layer0_outputs(10087) <= b and not a;
    layer0_outputs(10088) <= '1';
    layer0_outputs(10089) <= not a;
    layer0_outputs(10090) <= not a or b;
    layer0_outputs(10091) <= not a or b;
    layer0_outputs(10092) <= a and b;
    layer0_outputs(10093) <= a xor b;
    layer0_outputs(10094) <= not a or b;
    layer0_outputs(10095) <= a;
    layer0_outputs(10096) <= b and not a;
    layer0_outputs(10097) <= a;
    layer0_outputs(10098) <= '0';
    layer0_outputs(10099) <= not (a xor b);
    layer0_outputs(10100) <= not (a xor b);
    layer0_outputs(10101) <= not a;
    layer0_outputs(10102) <= a and not b;
    layer0_outputs(10103) <= b;
    layer0_outputs(10104) <= not a;
    layer0_outputs(10105) <= a or b;
    layer0_outputs(10106) <= not a;
    layer0_outputs(10107) <= not b;
    layer0_outputs(10108) <= not b;
    layer0_outputs(10109) <= not b;
    layer0_outputs(10110) <= a and not b;
    layer0_outputs(10111) <= '1';
    layer0_outputs(10112) <= not (a and b);
    layer0_outputs(10113) <= a and not b;
    layer0_outputs(10114) <= not b or a;
    layer0_outputs(10115) <= a and b;
    layer0_outputs(10116) <= a and not b;
    layer0_outputs(10117) <= b and not a;
    layer0_outputs(10118) <= not (a and b);
    layer0_outputs(10119) <= not (a or b);
    layer0_outputs(10120) <= b;
    layer0_outputs(10121) <= not a or b;
    layer0_outputs(10122) <= not b or a;
    layer0_outputs(10123) <= a and not b;
    layer0_outputs(10124) <= a or b;
    layer0_outputs(10125) <= a and not b;
    layer0_outputs(10126) <= b;
    layer0_outputs(10127) <= not (a xor b);
    layer0_outputs(10128) <= a;
    layer0_outputs(10129) <= '1';
    layer0_outputs(10130) <= a and b;
    layer0_outputs(10131) <= a or b;
    layer0_outputs(10132) <= not a;
    layer0_outputs(10133) <= a or b;
    layer0_outputs(10134) <= b and not a;
    layer0_outputs(10135) <= b;
    layer0_outputs(10136) <= a and b;
    layer0_outputs(10137) <= b;
    layer0_outputs(10138) <= a or b;
    layer0_outputs(10139) <= not (a and b);
    layer0_outputs(10140) <= not b or a;
    layer0_outputs(10141) <= not a;
    layer0_outputs(10142) <= '1';
    layer0_outputs(10143) <= a and b;
    layer0_outputs(10144) <= a;
    layer0_outputs(10145) <= not b or a;
    layer0_outputs(10146) <= not b;
    layer0_outputs(10147) <= b and not a;
    layer0_outputs(10148) <= not b;
    layer0_outputs(10149) <= '0';
    layer0_outputs(10150) <= not a;
    layer0_outputs(10151) <= not (a or b);
    layer0_outputs(10152) <= not (a and b);
    layer0_outputs(10153) <= '1';
    layer0_outputs(10154) <= '0';
    layer0_outputs(10155) <= not (a or b);
    layer0_outputs(10156) <= a and not b;
    layer0_outputs(10157) <= not a or b;
    layer0_outputs(10158) <= a xor b;
    layer0_outputs(10159) <= a;
    layer0_outputs(10160) <= a and not b;
    layer0_outputs(10161) <= a or b;
    layer0_outputs(10162) <= not (a or b);
    layer0_outputs(10163) <= not b or a;
    layer0_outputs(10164) <= not (a xor b);
    layer0_outputs(10165) <= not b;
    layer0_outputs(10166) <= a xor b;
    layer0_outputs(10167) <= not a;
    layer0_outputs(10168) <= not a;
    layer0_outputs(10169) <= not (a or b);
    layer0_outputs(10170) <= '0';
    layer0_outputs(10171) <= not b or a;
    layer0_outputs(10172) <= '0';
    layer0_outputs(10173) <= not a or b;
    layer0_outputs(10174) <= '0';
    layer0_outputs(10175) <= not (a and b);
    layer0_outputs(10176) <= a;
    layer0_outputs(10177) <= a xor b;
    layer0_outputs(10178) <= not a;
    layer0_outputs(10179) <= not (a and b);
    layer0_outputs(10180) <= a or b;
    layer0_outputs(10181) <= not a or b;
    layer0_outputs(10182) <= not b or a;
    layer0_outputs(10183) <= a and not b;
    layer0_outputs(10184) <= a xor b;
    layer0_outputs(10185) <= b and not a;
    layer0_outputs(10186) <= '0';
    layer0_outputs(10187) <= not a;
    layer0_outputs(10188) <= a or b;
    layer0_outputs(10189) <= a or b;
    layer0_outputs(10190) <= not a;
    layer0_outputs(10191) <= not (a and b);
    layer0_outputs(10192) <= not (a or b);
    layer0_outputs(10193) <= a and not b;
    layer0_outputs(10194) <= not a or b;
    layer0_outputs(10195) <= not b;
    layer0_outputs(10196) <= not b;
    layer0_outputs(10197) <= not (a xor b);
    layer0_outputs(10198) <= not a or b;
    layer0_outputs(10199) <= not (a and b);
    layer0_outputs(10200) <= a or b;
    layer0_outputs(10201) <= a and not b;
    layer0_outputs(10202) <= not b or a;
    layer0_outputs(10203) <= a;
    layer0_outputs(10204) <= '1';
    layer0_outputs(10205) <= '0';
    layer0_outputs(10206) <= not a or b;
    layer0_outputs(10207) <= a xor b;
    layer0_outputs(10208) <= a xor b;
    layer0_outputs(10209) <= '0';
    layer0_outputs(10210) <= not b;
    layer0_outputs(10211) <= not (a or b);
    layer0_outputs(10212) <= b;
    layer0_outputs(10213) <= not a or b;
    layer0_outputs(10214) <= a xor b;
    layer0_outputs(10215) <= a and b;
    layer0_outputs(10216) <= not (a xor b);
    layer0_outputs(10217) <= a and b;
    layer0_outputs(10218) <= a or b;
    layer0_outputs(10219) <= b;
    layer0_outputs(10220) <= not a or b;
    layer0_outputs(10221) <= '1';
    layer0_outputs(10222) <= not b or a;
    layer0_outputs(10223) <= a xor b;
    layer0_outputs(10224) <= '0';
    layer0_outputs(10225) <= a or b;
    layer0_outputs(10226) <= not a;
    layer0_outputs(10227) <= not a;
    layer0_outputs(10228) <= b;
    layer0_outputs(10229) <= b;
    layer0_outputs(10230) <= not (a and b);
    layer0_outputs(10231) <= b;
    layer0_outputs(10232) <= not b or a;
    layer0_outputs(10233) <= not (a xor b);
    layer0_outputs(10234) <= '0';
    layer0_outputs(10235) <= not a or b;
    layer0_outputs(10236) <= not a or b;
    layer0_outputs(10237) <= not (a or b);
    layer0_outputs(10238) <= not b;
    layer0_outputs(10239) <= a or b;
    layer0_outputs(10240) <= not a;
    layer0_outputs(10241) <= not (a xor b);
    layer0_outputs(10242) <= not (a xor b);
    layer0_outputs(10243) <= not (a and b);
    layer0_outputs(10244) <= not (a or b);
    layer0_outputs(10245) <= not b;
    layer0_outputs(10246) <= a and b;
    layer0_outputs(10247) <= a;
    layer0_outputs(10248) <= '1';
    layer0_outputs(10249) <= not b;
    layer0_outputs(10250) <= not b or a;
    layer0_outputs(10251) <= a xor b;
    layer0_outputs(10252) <= '0';
    layer0_outputs(10253) <= b and not a;
    layer0_outputs(10254) <= not b or a;
    layer0_outputs(10255) <= not (a xor b);
    layer0_outputs(10256) <= not b;
    layer0_outputs(10257) <= b;
    layer0_outputs(10258) <= '0';
    layer0_outputs(10259) <= not b;
    layer0_outputs(10260) <= not (a xor b);
    layer0_outputs(10261) <= b;
    layer0_outputs(10262) <= a and not b;
    layer0_outputs(10263) <= not (a or b);
    layer0_outputs(10264) <= a and not b;
    layer0_outputs(10265) <= not a or b;
    layer0_outputs(10266) <= a;
    layer0_outputs(10267) <= b;
    layer0_outputs(10268) <= b and not a;
    layer0_outputs(10269) <= '1';
    layer0_outputs(10270) <= not (a xor b);
    layer0_outputs(10271) <= b;
    layer0_outputs(10272) <= a or b;
    layer0_outputs(10273) <= not a or b;
    layer0_outputs(10274) <= not (a or b);
    layer0_outputs(10275) <= a or b;
    layer0_outputs(10276) <= a xor b;
    layer0_outputs(10277) <= b and not a;
    layer0_outputs(10278) <= not (a xor b);
    layer0_outputs(10279) <= a;
    layer0_outputs(10280) <= a;
    layer0_outputs(10281) <= not (a or b);
    layer0_outputs(10282) <= a or b;
    layer0_outputs(10283) <= '0';
    layer0_outputs(10284) <= not a;
    layer0_outputs(10285) <= '1';
    layer0_outputs(10286) <= not a or b;
    layer0_outputs(10287) <= not b;
    layer0_outputs(10288) <= b;
    layer0_outputs(10289) <= a and not b;
    layer0_outputs(10290) <= b and not a;
    layer0_outputs(10291) <= not (a or b);
    layer0_outputs(10292) <= a xor b;
    layer0_outputs(10293) <= a;
    layer0_outputs(10294) <= not (a or b);
    layer0_outputs(10295) <= not (a and b);
    layer0_outputs(10296) <= not a or b;
    layer0_outputs(10297) <= a and b;
    layer0_outputs(10298) <= a xor b;
    layer0_outputs(10299) <= a or b;
    layer0_outputs(10300) <= a xor b;
    layer0_outputs(10301) <= not b or a;
    layer0_outputs(10302) <= a and not b;
    layer0_outputs(10303) <= not a;
    layer0_outputs(10304) <= a and not b;
    layer0_outputs(10305) <= a;
    layer0_outputs(10306) <= not (a or b);
    layer0_outputs(10307) <= a xor b;
    layer0_outputs(10308) <= not (a or b);
    layer0_outputs(10309) <= a and not b;
    layer0_outputs(10310) <= a and b;
    layer0_outputs(10311) <= a;
    layer0_outputs(10312) <= not (a xor b);
    layer0_outputs(10313) <= not (a and b);
    layer0_outputs(10314) <= a and not b;
    layer0_outputs(10315) <= not (a or b);
    layer0_outputs(10316) <= not b;
    layer0_outputs(10317) <= a or b;
    layer0_outputs(10318) <= b;
    layer0_outputs(10319) <= not a or b;
    layer0_outputs(10320) <= a or b;
    layer0_outputs(10321) <= not b or a;
    layer0_outputs(10322) <= a or b;
    layer0_outputs(10323) <= a or b;
    layer0_outputs(10324) <= not b or a;
    layer0_outputs(10325) <= a and b;
    layer0_outputs(10326) <= '0';
    layer0_outputs(10327) <= not b;
    layer0_outputs(10328) <= not (a or b);
    layer0_outputs(10329) <= b;
    layer0_outputs(10330) <= '1';
    layer0_outputs(10331) <= not a or b;
    layer0_outputs(10332) <= '0';
    layer0_outputs(10333) <= not b;
    layer0_outputs(10334) <= not (a and b);
    layer0_outputs(10335) <= not a or b;
    layer0_outputs(10336) <= '1';
    layer0_outputs(10337) <= b;
    layer0_outputs(10338) <= b and not a;
    layer0_outputs(10339) <= a xor b;
    layer0_outputs(10340) <= b;
    layer0_outputs(10341) <= a and b;
    layer0_outputs(10342) <= b and not a;
    layer0_outputs(10343) <= not (a xor b);
    layer0_outputs(10344) <= b and not a;
    layer0_outputs(10345) <= '0';
    layer0_outputs(10346) <= '0';
    layer0_outputs(10347) <= b;
    layer0_outputs(10348) <= not b;
    layer0_outputs(10349) <= not (a xor b);
    layer0_outputs(10350) <= not (a or b);
    layer0_outputs(10351) <= not a;
    layer0_outputs(10352) <= not a or b;
    layer0_outputs(10353) <= '1';
    layer0_outputs(10354) <= '1';
    layer0_outputs(10355) <= a;
    layer0_outputs(10356) <= not a or b;
    layer0_outputs(10357) <= not (a xor b);
    layer0_outputs(10358) <= a and b;
    layer0_outputs(10359) <= a or b;
    layer0_outputs(10360) <= not b or a;
    layer0_outputs(10361) <= not a;
    layer0_outputs(10362) <= not b or a;
    layer0_outputs(10363) <= not a;
    layer0_outputs(10364) <= b and not a;
    layer0_outputs(10365) <= a or b;
    layer0_outputs(10366) <= '0';
    layer0_outputs(10367) <= a;
    layer0_outputs(10368) <= a;
    layer0_outputs(10369) <= b and not a;
    layer0_outputs(10370) <= b and not a;
    layer0_outputs(10371) <= not (a and b);
    layer0_outputs(10372) <= not (a and b);
    layer0_outputs(10373) <= not a;
    layer0_outputs(10374) <= a and b;
    layer0_outputs(10375) <= a and not b;
    layer0_outputs(10376) <= not (a xor b);
    layer0_outputs(10377) <= b and not a;
    layer0_outputs(10378) <= not b;
    layer0_outputs(10379) <= '1';
    layer0_outputs(10380) <= not a;
    layer0_outputs(10381) <= a or b;
    layer0_outputs(10382) <= not a;
    layer0_outputs(10383) <= a;
    layer0_outputs(10384) <= b;
    layer0_outputs(10385) <= not (a xor b);
    layer0_outputs(10386) <= a xor b;
    layer0_outputs(10387) <= a and b;
    layer0_outputs(10388) <= a and not b;
    layer0_outputs(10389) <= not b or a;
    layer0_outputs(10390) <= a;
    layer0_outputs(10391) <= b;
    layer0_outputs(10392) <= a and b;
    layer0_outputs(10393) <= not (a and b);
    layer0_outputs(10394) <= a;
    layer0_outputs(10395) <= '0';
    layer0_outputs(10396) <= a and not b;
    layer0_outputs(10397) <= a or b;
    layer0_outputs(10398) <= a xor b;
    layer0_outputs(10399) <= a;
    layer0_outputs(10400) <= a or b;
    layer0_outputs(10401) <= not b or a;
    layer0_outputs(10402) <= a xor b;
    layer0_outputs(10403) <= not (a and b);
    layer0_outputs(10404) <= a and not b;
    layer0_outputs(10405) <= not a;
    layer0_outputs(10406) <= not (a or b);
    layer0_outputs(10407) <= not b;
    layer0_outputs(10408) <= '0';
    layer0_outputs(10409) <= not (a xor b);
    layer0_outputs(10410) <= b and not a;
    layer0_outputs(10411) <= a xor b;
    layer0_outputs(10412) <= not (a or b);
    layer0_outputs(10413) <= not b;
    layer0_outputs(10414) <= b and not a;
    layer0_outputs(10415) <= a or b;
    layer0_outputs(10416) <= not a or b;
    layer0_outputs(10417) <= not b or a;
    layer0_outputs(10418) <= a;
    layer0_outputs(10419) <= a or b;
    layer0_outputs(10420) <= not a or b;
    layer0_outputs(10421) <= b;
    layer0_outputs(10422) <= not b;
    layer0_outputs(10423) <= not b or a;
    layer0_outputs(10424) <= not a or b;
    layer0_outputs(10425) <= not (a xor b);
    layer0_outputs(10426) <= a;
    layer0_outputs(10427) <= b and not a;
    layer0_outputs(10428) <= a;
    layer0_outputs(10429) <= not (a xor b);
    layer0_outputs(10430) <= not a;
    layer0_outputs(10431) <= not b or a;
    layer0_outputs(10432) <= a;
    layer0_outputs(10433) <= not (a xor b);
    layer0_outputs(10434) <= not b or a;
    layer0_outputs(10435) <= b and not a;
    layer0_outputs(10436) <= not (a or b);
    layer0_outputs(10437) <= not (a and b);
    layer0_outputs(10438) <= not (a and b);
    layer0_outputs(10439) <= a;
    layer0_outputs(10440) <= a;
    layer0_outputs(10441) <= b;
    layer0_outputs(10442) <= not a or b;
    layer0_outputs(10443) <= b;
    layer0_outputs(10444) <= not a or b;
    layer0_outputs(10445) <= not a or b;
    layer0_outputs(10446) <= not (a xor b);
    layer0_outputs(10447) <= not b;
    layer0_outputs(10448) <= not (a or b);
    layer0_outputs(10449) <= not a;
    layer0_outputs(10450) <= b;
    layer0_outputs(10451) <= b;
    layer0_outputs(10452) <= not (a and b);
    layer0_outputs(10453) <= not a;
    layer0_outputs(10454) <= b;
    layer0_outputs(10455) <= not (a xor b);
    layer0_outputs(10456) <= not b or a;
    layer0_outputs(10457) <= a or b;
    layer0_outputs(10458) <= b and not a;
    layer0_outputs(10459) <= not b or a;
    layer0_outputs(10460) <= '1';
    layer0_outputs(10461) <= not a or b;
    layer0_outputs(10462) <= not b or a;
    layer0_outputs(10463) <= a and not b;
    layer0_outputs(10464) <= not (a or b);
    layer0_outputs(10465) <= not b or a;
    layer0_outputs(10466) <= not b or a;
    layer0_outputs(10467) <= not (a or b);
    layer0_outputs(10468) <= not a;
    layer0_outputs(10469) <= '1';
    layer0_outputs(10470) <= a and b;
    layer0_outputs(10471) <= not (a or b);
    layer0_outputs(10472) <= '0';
    layer0_outputs(10473) <= a or b;
    layer0_outputs(10474) <= '0';
    layer0_outputs(10475) <= not b;
    layer0_outputs(10476) <= a and not b;
    layer0_outputs(10477) <= not b;
    layer0_outputs(10478) <= not b;
    layer0_outputs(10479) <= a;
    layer0_outputs(10480) <= not b or a;
    layer0_outputs(10481) <= a and b;
    layer0_outputs(10482) <= not (a or b);
    layer0_outputs(10483) <= not (a or b);
    layer0_outputs(10484) <= not a or b;
    layer0_outputs(10485) <= not a or b;
    layer0_outputs(10486) <= not (a xor b);
    layer0_outputs(10487) <= not (a or b);
    layer0_outputs(10488) <= not (a or b);
    layer0_outputs(10489) <= '0';
    layer0_outputs(10490) <= a and b;
    layer0_outputs(10491) <= not a;
    layer0_outputs(10492) <= not a;
    layer0_outputs(10493) <= not (a or b);
    layer0_outputs(10494) <= not a;
    layer0_outputs(10495) <= a or b;
    layer0_outputs(10496) <= a xor b;
    layer0_outputs(10497) <= a;
    layer0_outputs(10498) <= not b or a;
    layer0_outputs(10499) <= a;
    layer0_outputs(10500) <= a and not b;
    layer0_outputs(10501) <= b and not a;
    layer0_outputs(10502) <= not b or a;
    layer0_outputs(10503) <= not b;
    layer0_outputs(10504) <= not a or b;
    layer0_outputs(10505) <= not b;
    layer0_outputs(10506) <= a xor b;
    layer0_outputs(10507) <= '1';
    layer0_outputs(10508) <= b;
    layer0_outputs(10509) <= not b or a;
    layer0_outputs(10510) <= not a;
    layer0_outputs(10511) <= not (a xor b);
    layer0_outputs(10512) <= not (a and b);
    layer0_outputs(10513) <= b and not a;
    layer0_outputs(10514) <= b and not a;
    layer0_outputs(10515) <= a;
    layer0_outputs(10516) <= not a;
    layer0_outputs(10517) <= not b or a;
    layer0_outputs(10518) <= '0';
    layer0_outputs(10519) <= b;
    layer0_outputs(10520) <= not a;
    layer0_outputs(10521) <= not b;
    layer0_outputs(10522) <= not b or a;
    layer0_outputs(10523) <= not b or a;
    layer0_outputs(10524) <= not (a or b);
    layer0_outputs(10525) <= not (a xor b);
    layer0_outputs(10526) <= not (a and b);
    layer0_outputs(10527) <= a or b;
    layer0_outputs(10528) <= not a;
    layer0_outputs(10529) <= a or b;
    layer0_outputs(10530) <= not b;
    layer0_outputs(10531) <= a;
    layer0_outputs(10532) <= not a;
    layer0_outputs(10533) <= not (a xor b);
    layer0_outputs(10534) <= not a;
    layer0_outputs(10535) <= a xor b;
    layer0_outputs(10536) <= not a;
    layer0_outputs(10537) <= b;
    layer0_outputs(10538) <= a or b;
    layer0_outputs(10539) <= not (a and b);
    layer0_outputs(10540) <= not a;
    layer0_outputs(10541) <= not (a xor b);
    layer0_outputs(10542) <= b and not a;
    layer0_outputs(10543) <= not (a and b);
    layer0_outputs(10544) <= not (a or b);
    layer0_outputs(10545) <= not b;
    layer0_outputs(10546) <= b;
    layer0_outputs(10547) <= not (a or b);
    layer0_outputs(10548) <= a and not b;
    layer0_outputs(10549) <= a or b;
    layer0_outputs(10550) <= not (a or b);
    layer0_outputs(10551) <= a or b;
    layer0_outputs(10552) <= b and not a;
    layer0_outputs(10553) <= not (a or b);
    layer0_outputs(10554) <= not b;
    layer0_outputs(10555) <= not b;
    layer0_outputs(10556) <= not a or b;
    layer0_outputs(10557) <= a or b;
    layer0_outputs(10558) <= a or b;
    layer0_outputs(10559) <= not a or b;
    layer0_outputs(10560) <= b;
    layer0_outputs(10561) <= not b;
    layer0_outputs(10562) <= a xor b;
    layer0_outputs(10563) <= not b or a;
    layer0_outputs(10564) <= a;
    layer0_outputs(10565) <= not b or a;
    layer0_outputs(10566) <= not (a or b);
    layer0_outputs(10567) <= b;
    layer0_outputs(10568) <= b and not a;
    layer0_outputs(10569) <= '1';
    layer0_outputs(10570) <= '0';
    layer0_outputs(10571) <= b and not a;
    layer0_outputs(10572) <= not (a and b);
    layer0_outputs(10573) <= '1';
    layer0_outputs(10574) <= b;
    layer0_outputs(10575) <= not b or a;
    layer0_outputs(10576) <= not (a or b);
    layer0_outputs(10577) <= '1';
    layer0_outputs(10578) <= a and not b;
    layer0_outputs(10579) <= b;
    layer0_outputs(10580) <= not (a or b);
    layer0_outputs(10581) <= not (a xor b);
    layer0_outputs(10582) <= not (a xor b);
    layer0_outputs(10583) <= not a or b;
    layer0_outputs(10584) <= a or b;
    layer0_outputs(10585) <= b;
    layer0_outputs(10586) <= not (a or b);
    layer0_outputs(10587) <= a and not b;
    layer0_outputs(10588) <= not a or b;
    layer0_outputs(10589) <= not (a or b);
    layer0_outputs(10590) <= not (a and b);
    layer0_outputs(10591) <= not (a xor b);
    layer0_outputs(10592) <= a or b;
    layer0_outputs(10593) <= a and not b;
    layer0_outputs(10594) <= a;
    layer0_outputs(10595) <= a or b;
    layer0_outputs(10596) <= a or b;
    layer0_outputs(10597) <= '1';
    layer0_outputs(10598) <= not a;
    layer0_outputs(10599) <= a xor b;
    layer0_outputs(10600) <= b and not a;
    layer0_outputs(10601) <= a and b;
    layer0_outputs(10602) <= '1';
    layer0_outputs(10603) <= not (a xor b);
    layer0_outputs(10604) <= a xor b;
    layer0_outputs(10605) <= not (a and b);
    layer0_outputs(10606) <= b and not a;
    layer0_outputs(10607) <= a xor b;
    layer0_outputs(10608) <= not (a or b);
    layer0_outputs(10609) <= b;
    layer0_outputs(10610) <= a and b;
    layer0_outputs(10611) <= a and not b;
    layer0_outputs(10612) <= b;
    layer0_outputs(10613) <= not (a or b);
    layer0_outputs(10614) <= not a or b;
    layer0_outputs(10615) <= b;
    layer0_outputs(10616) <= not a or b;
    layer0_outputs(10617) <= a xor b;
    layer0_outputs(10618) <= not a or b;
    layer0_outputs(10619) <= a or b;
    layer0_outputs(10620) <= not (a or b);
    layer0_outputs(10621) <= a and b;
    layer0_outputs(10622) <= a xor b;
    layer0_outputs(10623) <= a or b;
    layer0_outputs(10624) <= a and b;
    layer0_outputs(10625) <= '0';
    layer0_outputs(10626) <= not (a and b);
    layer0_outputs(10627) <= a;
    layer0_outputs(10628) <= not b or a;
    layer0_outputs(10629) <= not (a xor b);
    layer0_outputs(10630) <= a and not b;
    layer0_outputs(10631) <= a and b;
    layer0_outputs(10632) <= a xor b;
    layer0_outputs(10633) <= a and not b;
    layer0_outputs(10634) <= not b;
    layer0_outputs(10635) <= a;
    layer0_outputs(10636) <= a;
    layer0_outputs(10637) <= not b;
    layer0_outputs(10638) <= b and not a;
    layer0_outputs(10639) <= not (a or b);
    layer0_outputs(10640) <= b and not a;
    layer0_outputs(10641) <= not (a xor b);
    layer0_outputs(10642) <= not b;
    layer0_outputs(10643) <= not (a and b);
    layer0_outputs(10644) <= not (a or b);
    layer0_outputs(10645) <= not (a or b);
    layer0_outputs(10646) <= not (a or b);
    layer0_outputs(10647) <= a and not b;
    layer0_outputs(10648) <= a xor b;
    layer0_outputs(10649) <= '1';
    layer0_outputs(10650) <= not b or a;
    layer0_outputs(10651) <= a or b;
    layer0_outputs(10652) <= not a;
    layer0_outputs(10653) <= '1';
    layer0_outputs(10654) <= a or b;
    layer0_outputs(10655) <= not (a xor b);
    layer0_outputs(10656) <= '0';
    layer0_outputs(10657) <= b and not a;
    layer0_outputs(10658) <= b;
    layer0_outputs(10659) <= not b or a;
    layer0_outputs(10660) <= not b or a;
    layer0_outputs(10661) <= '0';
    layer0_outputs(10662) <= a xor b;
    layer0_outputs(10663) <= not (a or b);
    layer0_outputs(10664) <= a;
    layer0_outputs(10665) <= a;
    layer0_outputs(10666) <= not b or a;
    layer0_outputs(10667) <= not b;
    layer0_outputs(10668) <= b and not a;
    layer0_outputs(10669) <= not (a or b);
    layer0_outputs(10670) <= '0';
    layer0_outputs(10671) <= '0';
    layer0_outputs(10672) <= b and not a;
    layer0_outputs(10673) <= a or b;
    layer0_outputs(10674) <= not (a or b);
    layer0_outputs(10675) <= '0';
    layer0_outputs(10676) <= not a;
    layer0_outputs(10677) <= '0';
    layer0_outputs(10678) <= '1';
    layer0_outputs(10679) <= a and not b;
    layer0_outputs(10680) <= not b;
    layer0_outputs(10681) <= a and b;
    layer0_outputs(10682) <= '0';
    layer0_outputs(10683) <= not (a or b);
    layer0_outputs(10684) <= b;
    layer0_outputs(10685) <= a and not b;
    layer0_outputs(10686) <= a;
    layer0_outputs(10687) <= '0';
    layer0_outputs(10688) <= a;
    layer0_outputs(10689) <= not (a xor b);
    layer0_outputs(10690) <= not b or a;
    layer0_outputs(10691) <= not b or a;
    layer0_outputs(10692) <= a and not b;
    layer0_outputs(10693) <= not (a or b);
    layer0_outputs(10694) <= a and not b;
    layer0_outputs(10695) <= not (a xor b);
    layer0_outputs(10696) <= '0';
    layer0_outputs(10697) <= not (a xor b);
    layer0_outputs(10698) <= not (a or b);
    layer0_outputs(10699) <= b;
    layer0_outputs(10700) <= a xor b;
    layer0_outputs(10701) <= not a;
    layer0_outputs(10702) <= a;
    layer0_outputs(10703) <= a and not b;
    layer0_outputs(10704) <= '0';
    layer0_outputs(10705) <= a or b;
    layer0_outputs(10706) <= '0';
    layer0_outputs(10707) <= a and b;
    layer0_outputs(10708) <= not (a xor b);
    layer0_outputs(10709) <= not (a and b);
    layer0_outputs(10710) <= b and not a;
    layer0_outputs(10711) <= '0';
    layer0_outputs(10712) <= a;
    layer0_outputs(10713) <= not (a xor b);
    layer0_outputs(10714) <= '1';
    layer0_outputs(10715) <= '0';
    layer0_outputs(10716) <= not (a xor b);
    layer0_outputs(10717) <= '0';
    layer0_outputs(10718) <= '0';
    layer0_outputs(10719) <= '0';
    layer0_outputs(10720) <= a and b;
    layer0_outputs(10721) <= b;
    layer0_outputs(10722) <= not (a or b);
    layer0_outputs(10723) <= a or b;
    layer0_outputs(10724) <= a and b;
    layer0_outputs(10725) <= a xor b;
    layer0_outputs(10726) <= '1';
    layer0_outputs(10727) <= not (a and b);
    layer0_outputs(10728) <= a and b;
    layer0_outputs(10729) <= not (a and b);
    layer0_outputs(10730) <= not (a and b);
    layer0_outputs(10731) <= '0';
    layer0_outputs(10732) <= b and not a;
    layer0_outputs(10733) <= b;
    layer0_outputs(10734) <= a or b;
    layer0_outputs(10735) <= a or b;
    layer0_outputs(10736) <= b;
    layer0_outputs(10737) <= not b or a;
    layer0_outputs(10738) <= not (a or b);
    layer0_outputs(10739) <= not a or b;
    layer0_outputs(10740) <= not b;
    layer0_outputs(10741) <= not a or b;
    layer0_outputs(10742) <= a and b;
    layer0_outputs(10743) <= not (a xor b);
    layer0_outputs(10744) <= not (a xor b);
    layer0_outputs(10745) <= not (a xor b);
    layer0_outputs(10746) <= b and not a;
    layer0_outputs(10747) <= not (a or b);
    layer0_outputs(10748) <= not (a and b);
    layer0_outputs(10749) <= b;
    layer0_outputs(10750) <= a;
    layer0_outputs(10751) <= not (a or b);
    layer0_outputs(10752) <= '0';
    layer0_outputs(10753) <= not (a or b);
    layer0_outputs(10754) <= a or b;
    layer0_outputs(10755) <= a;
    layer0_outputs(10756) <= '0';
    layer0_outputs(10757) <= not a or b;
    layer0_outputs(10758) <= a and b;
    layer0_outputs(10759) <= a;
    layer0_outputs(10760) <= not a;
    layer0_outputs(10761) <= not b;
    layer0_outputs(10762) <= b and not a;
    layer0_outputs(10763) <= b;
    layer0_outputs(10764) <= not b or a;
    layer0_outputs(10765) <= '1';
    layer0_outputs(10766) <= b and not a;
    layer0_outputs(10767) <= not a;
    layer0_outputs(10768) <= not a;
    layer0_outputs(10769) <= not (a and b);
    layer0_outputs(10770) <= not (a or b);
    layer0_outputs(10771) <= not a;
    layer0_outputs(10772) <= a or b;
    layer0_outputs(10773) <= b and not a;
    layer0_outputs(10774) <= not (a or b);
    layer0_outputs(10775) <= a xor b;
    layer0_outputs(10776) <= b;
    layer0_outputs(10777) <= a and b;
    layer0_outputs(10778) <= a or b;
    layer0_outputs(10779) <= not a or b;
    layer0_outputs(10780) <= a and not b;
    layer0_outputs(10781) <= not b;
    layer0_outputs(10782) <= '0';
    layer0_outputs(10783) <= not b;
    layer0_outputs(10784) <= not b or a;
    layer0_outputs(10785) <= a xor b;
    layer0_outputs(10786) <= not b;
    layer0_outputs(10787) <= not a;
    layer0_outputs(10788) <= a or b;
    layer0_outputs(10789) <= not b;
    layer0_outputs(10790) <= a xor b;
    layer0_outputs(10791) <= not b or a;
    layer0_outputs(10792) <= not (a or b);
    layer0_outputs(10793) <= not (a xor b);
    layer0_outputs(10794) <= a and not b;
    layer0_outputs(10795) <= not a or b;
    layer0_outputs(10796) <= b and not a;
    layer0_outputs(10797) <= not a;
    layer0_outputs(10798) <= a and b;
    layer0_outputs(10799) <= '0';
    layer0_outputs(10800) <= not (a or b);
    layer0_outputs(10801) <= a or b;
    layer0_outputs(10802) <= not (a or b);
    layer0_outputs(10803) <= not b;
    layer0_outputs(10804) <= a;
    layer0_outputs(10805) <= not (a or b);
    layer0_outputs(10806) <= b;
    layer0_outputs(10807) <= not b;
    layer0_outputs(10808) <= a and not b;
    layer0_outputs(10809) <= not (a or b);
    layer0_outputs(10810) <= not (a or b);
    layer0_outputs(10811) <= '0';
    layer0_outputs(10812) <= not a or b;
    layer0_outputs(10813) <= not b or a;
    layer0_outputs(10814) <= not b;
    layer0_outputs(10815) <= a or b;
    layer0_outputs(10816) <= a and not b;
    layer0_outputs(10817) <= a;
    layer0_outputs(10818) <= a xor b;
    layer0_outputs(10819) <= not (a or b);
    layer0_outputs(10820) <= not a or b;
    layer0_outputs(10821) <= not (a or b);
    layer0_outputs(10822) <= a and not b;
    layer0_outputs(10823) <= not a or b;
    layer0_outputs(10824) <= a or b;
    layer0_outputs(10825) <= not a;
    layer0_outputs(10826) <= not a or b;
    layer0_outputs(10827) <= not a or b;
    layer0_outputs(10828) <= a xor b;
    layer0_outputs(10829) <= b and not a;
    layer0_outputs(10830) <= a;
    layer0_outputs(10831) <= not (a xor b);
    layer0_outputs(10832) <= not (a xor b);
    layer0_outputs(10833) <= a and b;
    layer0_outputs(10834) <= a and not b;
    layer0_outputs(10835) <= not a;
    layer0_outputs(10836) <= a;
    layer0_outputs(10837) <= a or b;
    layer0_outputs(10838) <= '0';
    layer0_outputs(10839) <= '1';
    layer0_outputs(10840) <= a;
    layer0_outputs(10841) <= not a;
    layer0_outputs(10842) <= not (a xor b);
    layer0_outputs(10843) <= not (a xor b);
    layer0_outputs(10844) <= b;
    layer0_outputs(10845) <= a or b;
    layer0_outputs(10846) <= a xor b;
    layer0_outputs(10847) <= not (a and b);
    layer0_outputs(10848) <= '0';
    layer0_outputs(10849) <= b and not a;
    layer0_outputs(10850) <= a or b;
    layer0_outputs(10851) <= a xor b;
    layer0_outputs(10852) <= not b;
    layer0_outputs(10853) <= a or b;
    layer0_outputs(10854) <= a and b;
    layer0_outputs(10855) <= not a or b;
    layer0_outputs(10856) <= a and b;
    layer0_outputs(10857) <= not b or a;
    layer0_outputs(10858) <= a xor b;
    layer0_outputs(10859) <= b and not a;
    layer0_outputs(10860) <= not b or a;
    layer0_outputs(10861) <= not a;
    layer0_outputs(10862) <= not (a and b);
    layer0_outputs(10863) <= not (a or b);
    layer0_outputs(10864) <= a or b;
    layer0_outputs(10865) <= not b or a;
    layer0_outputs(10866) <= not (a and b);
    layer0_outputs(10867) <= '1';
    layer0_outputs(10868) <= not (a or b);
    layer0_outputs(10869) <= not (a or b);
    layer0_outputs(10870) <= not b or a;
    layer0_outputs(10871) <= not (a or b);
    layer0_outputs(10872) <= not (a xor b);
    layer0_outputs(10873) <= a;
    layer0_outputs(10874) <= a;
    layer0_outputs(10875) <= not b;
    layer0_outputs(10876) <= not a or b;
    layer0_outputs(10877) <= not a or b;
    layer0_outputs(10878) <= a and b;
    layer0_outputs(10879) <= not (a xor b);
    layer0_outputs(10880) <= a and not b;
    layer0_outputs(10881) <= a xor b;
    layer0_outputs(10882) <= a;
    layer0_outputs(10883) <= not a or b;
    layer0_outputs(10884) <= not b;
    layer0_outputs(10885) <= '1';
    layer0_outputs(10886) <= a;
    layer0_outputs(10887) <= not b;
    layer0_outputs(10888) <= not (a xor b);
    layer0_outputs(10889) <= not a or b;
    layer0_outputs(10890) <= not (a xor b);
    layer0_outputs(10891) <= a or b;
    layer0_outputs(10892) <= a or b;
    layer0_outputs(10893) <= b and not a;
    layer0_outputs(10894) <= not a;
    layer0_outputs(10895) <= not (a xor b);
    layer0_outputs(10896) <= b and not a;
    layer0_outputs(10897) <= not b;
    layer0_outputs(10898) <= a or b;
    layer0_outputs(10899) <= a and not b;
    layer0_outputs(10900) <= a;
    layer0_outputs(10901) <= b;
    layer0_outputs(10902) <= b and not a;
    layer0_outputs(10903) <= not (a or b);
    layer0_outputs(10904) <= not a;
    layer0_outputs(10905) <= b and not a;
    layer0_outputs(10906) <= not a;
    layer0_outputs(10907) <= not b;
    layer0_outputs(10908) <= b;
    layer0_outputs(10909) <= not b;
    layer0_outputs(10910) <= not (a xor b);
    layer0_outputs(10911) <= not (a or b);
    layer0_outputs(10912) <= not a;
    layer0_outputs(10913) <= '0';
    layer0_outputs(10914) <= b and not a;
    layer0_outputs(10915) <= a and not b;
    layer0_outputs(10916) <= not a or b;
    layer0_outputs(10917) <= a or b;
    layer0_outputs(10918) <= b;
    layer0_outputs(10919) <= '0';
    layer0_outputs(10920) <= a or b;
    layer0_outputs(10921) <= b;
    layer0_outputs(10922) <= not b;
    layer0_outputs(10923) <= not a or b;
    layer0_outputs(10924) <= not a or b;
    layer0_outputs(10925) <= not b;
    layer0_outputs(10926) <= not b or a;
    layer0_outputs(10927) <= not b;
    layer0_outputs(10928) <= a;
    layer0_outputs(10929) <= a or b;
    layer0_outputs(10930) <= not (a and b);
    layer0_outputs(10931) <= a;
    layer0_outputs(10932) <= not b;
    layer0_outputs(10933) <= not a;
    layer0_outputs(10934) <= not b;
    layer0_outputs(10935) <= not b;
    layer0_outputs(10936) <= b and not a;
    layer0_outputs(10937) <= b;
    layer0_outputs(10938) <= a or b;
    layer0_outputs(10939) <= a;
    layer0_outputs(10940) <= a or b;
    layer0_outputs(10941) <= '0';
    layer0_outputs(10942) <= b and not a;
    layer0_outputs(10943) <= a;
    layer0_outputs(10944) <= a or b;
    layer0_outputs(10945) <= not (a or b);
    layer0_outputs(10946) <= '1';
    layer0_outputs(10947) <= not b or a;
    layer0_outputs(10948) <= not a;
    layer0_outputs(10949) <= '1';
    layer0_outputs(10950) <= not b or a;
    layer0_outputs(10951) <= b;
    layer0_outputs(10952) <= not (a and b);
    layer0_outputs(10953) <= not (a or b);
    layer0_outputs(10954) <= b;
    layer0_outputs(10955) <= not (a xor b);
    layer0_outputs(10956) <= not (a or b);
    layer0_outputs(10957) <= not (a xor b);
    layer0_outputs(10958) <= not (a or b);
    layer0_outputs(10959) <= '0';
    layer0_outputs(10960) <= b and not a;
    layer0_outputs(10961) <= a;
    layer0_outputs(10962) <= a or b;
    layer0_outputs(10963) <= a;
    layer0_outputs(10964) <= not a or b;
    layer0_outputs(10965) <= b and not a;
    layer0_outputs(10966) <= not (a xor b);
    layer0_outputs(10967) <= not a;
    layer0_outputs(10968) <= a and b;
    layer0_outputs(10969) <= not (a xor b);
    layer0_outputs(10970) <= '0';
    layer0_outputs(10971) <= not (a xor b);
    layer0_outputs(10972) <= not b;
    layer0_outputs(10973) <= a or b;
    layer0_outputs(10974) <= not b or a;
    layer0_outputs(10975) <= a or b;
    layer0_outputs(10976) <= '1';
    layer0_outputs(10977) <= not a or b;
    layer0_outputs(10978) <= a or b;
    layer0_outputs(10979) <= '1';
    layer0_outputs(10980) <= b and not a;
    layer0_outputs(10981) <= b and not a;
    layer0_outputs(10982) <= not (a xor b);
    layer0_outputs(10983) <= not (a xor b);
    layer0_outputs(10984) <= a xor b;
    layer0_outputs(10985) <= not b or a;
    layer0_outputs(10986) <= a;
    layer0_outputs(10987) <= '1';
    layer0_outputs(10988) <= not a;
    layer0_outputs(10989) <= not a;
    layer0_outputs(10990) <= not a or b;
    layer0_outputs(10991) <= not a or b;
    layer0_outputs(10992) <= a xor b;
    layer0_outputs(10993) <= not (a xor b);
    layer0_outputs(10994) <= not a;
    layer0_outputs(10995) <= not (a or b);
    layer0_outputs(10996) <= a xor b;
    layer0_outputs(10997) <= '0';
    layer0_outputs(10998) <= a and not b;
    layer0_outputs(10999) <= a and not b;
    layer0_outputs(11000) <= a and not b;
    layer0_outputs(11001) <= a xor b;
    layer0_outputs(11002) <= b;
    layer0_outputs(11003) <= a or b;
    layer0_outputs(11004) <= '1';
    layer0_outputs(11005) <= not a or b;
    layer0_outputs(11006) <= a or b;
    layer0_outputs(11007) <= not a or b;
    layer0_outputs(11008) <= b and not a;
    layer0_outputs(11009) <= b;
    layer0_outputs(11010) <= not a;
    layer0_outputs(11011) <= not (a and b);
    layer0_outputs(11012) <= a and not b;
    layer0_outputs(11013) <= not a;
    layer0_outputs(11014) <= a and b;
    layer0_outputs(11015) <= not (a or b);
    layer0_outputs(11016) <= not b;
    layer0_outputs(11017) <= a and not b;
    layer0_outputs(11018) <= not (a and b);
    layer0_outputs(11019) <= '0';
    layer0_outputs(11020) <= '1';
    layer0_outputs(11021) <= a and not b;
    layer0_outputs(11022) <= not (a or b);
    layer0_outputs(11023) <= a xor b;
    layer0_outputs(11024) <= a and b;
    layer0_outputs(11025) <= not a or b;
    layer0_outputs(11026) <= not (a or b);
    layer0_outputs(11027) <= not a or b;
    layer0_outputs(11028) <= '0';
    layer0_outputs(11029) <= not b or a;
    layer0_outputs(11030) <= not b;
    layer0_outputs(11031) <= not (a and b);
    layer0_outputs(11032) <= not (a xor b);
    layer0_outputs(11033) <= a and not b;
    layer0_outputs(11034) <= b;
    layer0_outputs(11035) <= a xor b;
    layer0_outputs(11036) <= b;
    layer0_outputs(11037) <= not a;
    layer0_outputs(11038) <= b;
    layer0_outputs(11039) <= not (a and b);
    layer0_outputs(11040) <= not b;
    layer0_outputs(11041) <= not (a and b);
    layer0_outputs(11042) <= not (a and b);
    layer0_outputs(11043) <= a;
    layer0_outputs(11044) <= a or b;
    layer0_outputs(11045) <= not a;
    layer0_outputs(11046) <= a and not b;
    layer0_outputs(11047) <= a or b;
    layer0_outputs(11048) <= a or b;
    layer0_outputs(11049) <= a or b;
    layer0_outputs(11050) <= a and not b;
    layer0_outputs(11051) <= a and b;
    layer0_outputs(11052) <= a or b;
    layer0_outputs(11053) <= b and not a;
    layer0_outputs(11054) <= not a or b;
    layer0_outputs(11055) <= b;
    layer0_outputs(11056) <= not (a or b);
    layer0_outputs(11057) <= a xor b;
    layer0_outputs(11058) <= not (a or b);
    layer0_outputs(11059) <= not (a and b);
    layer0_outputs(11060) <= not b or a;
    layer0_outputs(11061) <= a;
    layer0_outputs(11062) <= b;
    layer0_outputs(11063) <= not a;
    layer0_outputs(11064) <= not b or a;
    layer0_outputs(11065) <= not (a xor b);
    layer0_outputs(11066) <= not (a xor b);
    layer0_outputs(11067) <= not a or b;
    layer0_outputs(11068) <= a and b;
    layer0_outputs(11069) <= not (a and b);
    layer0_outputs(11070) <= b and not a;
    layer0_outputs(11071) <= a;
    layer0_outputs(11072) <= '0';
    layer0_outputs(11073) <= not b;
    layer0_outputs(11074) <= a and b;
    layer0_outputs(11075) <= b and not a;
    layer0_outputs(11076) <= a;
    layer0_outputs(11077) <= not a;
    layer0_outputs(11078) <= a or b;
    layer0_outputs(11079) <= not (a and b);
    layer0_outputs(11080) <= a and not b;
    layer0_outputs(11081) <= not b;
    layer0_outputs(11082) <= not a or b;
    layer0_outputs(11083) <= b and not a;
    layer0_outputs(11084) <= a and b;
    layer0_outputs(11085) <= a xor b;
    layer0_outputs(11086) <= '0';
    layer0_outputs(11087) <= not b or a;
    layer0_outputs(11088) <= not (a and b);
    layer0_outputs(11089) <= b and not a;
    layer0_outputs(11090) <= not (a or b);
    layer0_outputs(11091) <= not (a and b);
    layer0_outputs(11092) <= a or b;
    layer0_outputs(11093) <= not b;
    layer0_outputs(11094) <= b and not a;
    layer0_outputs(11095) <= a;
    layer0_outputs(11096) <= a;
    layer0_outputs(11097) <= not (a or b);
    layer0_outputs(11098) <= not b;
    layer0_outputs(11099) <= a;
    layer0_outputs(11100) <= not b or a;
    layer0_outputs(11101) <= not a or b;
    layer0_outputs(11102) <= b;
    layer0_outputs(11103) <= b and not a;
    layer0_outputs(11104) <= not (a or b);
    layer0_outputs(11105) <= not b or a;
    layer0_outputs(11106) <= a;
    layer0_outputs(11107) <= b;
    layer0_outputs(11108) <= not (a xor b);
    layer0_outputs(11109) <= not a;
    layer0_outputs(11110) <= '0';
    layer0_outputs(11111) <= not (a or b);
    layer0_outputs(11112) <= '0';
    layer0_outputs(11113) <= not b;
    layer0_outputs(11114) <= not (a xor b);
    layer0_outputs(11115) <= not (a and b);
    layer0_outputs(11116) <= not b;
    layer0_outputs(11117) <= not (a and b);
    layer0_outputs(11118) <= a or b;
    layer0_outputs(11119) <= not b or a;
    layer0_outputs(11120) <= not a or b;
    layer0_outputs(11121) <= a or b;
    layer0_outputs(11122) <= not b;
    layer0_outputs(11123) <= a or b;
    layer0_outputs(11124) <= '0';
    layer0_outputs(11125) <= not (a and b);
    layer0_outputs(11126) <= not (a or b);
    layer0_outputs(11127) <= b and not a;
    layer0_outputs(11128) <= a;
    layer0_outputs(11129) <= not (a xor b);
    layer0_outputs(11130) <= '0';
    layer0_outputs(11131) <= b;
    layer0_outputs(11132) <= '0';
    layer0_outputs(11133) <= a and not b;
    layer0_outputs(11134) <= not (a or b);
    layer0_outputs(11135) <= not (a and b);
    layer0_outputs(11136) <= not (a or b);
    layer0_outputs(11137) <= not b or a;
    layer0_outputs(11138) <= a;
    layer0_outputs(11139) <= a;
    layer0_outputs(11140) <= a and not b;
    layer0_outputs(11141) <= not (a or b);
    layer0_outputs(11142) <= not a or b;
    layer0_outputs(11143) <= not b;
    layer0_outputs(11144) <= a and b;
    layer0_outputs(11145) <= b and not a;
    layer0_outputs(11146) <= not (a and b);
    layer0_outputs(11147) <= not a;
    layer0_outputs(11148) <= not a or b;
    layer0_outputs(11149) <= a or b;
    layer0_outputs(11150) <= b;
    layer0_outputs(11151) <= a xor b;
    layer0_outputs(11152) <= a or b;
    layer0_outputs(11153) <= not a or b;
    layer0_outputs(11154) <= not b or a;
    layer0_outputs(11155) <= a xor b;
    layer0_outputs(11156) <= a xor b;
    layer0_outputs(11157) <= a xor b;
    layer0_outputs(11158) <= a or b;
    layer0_outputs(11159) <= a and not b;
    layer0_outputs(11160) <= not (a or b);
    layer0_outputs(11161) <= a and not b;
    layer0_outputs(11162) <= a and not b;
    layer0_outputs(11163) <= a xor b;
    layer0_outputs(11164) <= '0';
    layer0_outputs(11165) <= '0';
    layer0_outputs(11166) <= not (a and b);
    layer0_outputs(11167) <= b;
    layer0_outputs(11168) <= not b;
    layer0_outputs(11169) <= b and not a;
    layer0_outputs(11170) <= a and not b;
    layer0_outputs(11171) <= not b or a;
    layer0_outputs(11172) <= '0';
    layer0_outputs(11173) <= b;
    layer0_outputs(11174) <= not (a xor b);
    layer0_outputs(11175) <= b and not a;
    layer0_outputs(11176) <= b and not a;
    layer0_outputs(11177) <= a xor b;
    layer0_outputs(11178) <= a;
    layer0_outputs(11179) <= a or b;
    layer0_outputs(11180) <= not a;
    layer0_outputs(11181) <= a and b;
    layer0_outputs(11182) <= not (a and b);
    layer0_outputs(11183) <= not a;
    layer0_outputs(11184) <= a or b;
    layer0_outputs(11185) <= not b or a;
    layer0_outputs(11186) <= a;
    layer0_outputs(11187) <= not (a xor b);
    layer0_outputs(11188) <= not (a xor b);
    layer0_outputs(11189) <= '1';
    layer0_outputs(11190) <= '1';
    layer0_outputs(11191) <= b;
    layer0_outputs(11192) <= '0';
    layer0_outputs(11193) <= a xor b;
    layer0_outputs(11194) <= b and not a;
    layer0_outputs(11195) <= a and b;
    layer0_outputs(11196) <= a or b;
    layer0_outputs(11197) <= not (a xor b);
    layer0_outputs(11198) <= not (a or b);
    layer0_outputs(11199) <= b;
    layer0_outputs(11200) <= a and b;
    layer0_outputs(11201) <= not b;
    layer0_outputs(11202) <= not a;
    layer0_outputs(11203) <= a;
    layer0_outputs(11204) <= a;
    layer0_outputs(11205) <= not b;
    layer0_outputs(11206) <= not b or a;
    layer0_outputs(11207) <= a xor b;
    layer0_outputs(11208) <= not (a or b);
    layer0_outputs(11209) <= not a or b;
    layer0_outputs(11210) <= not (a or b);
    layer0_outputs(11211) <= not (a or b);
    layer0_outputs(11212) <= not (a xor b);
    layer0_outputs(11213) <= b and not a;
    layer0_outputs(11214) <= a xor b;
    layer0_outputs(11215) <= not b;
    layer0_outputs(11216) <= b;
    layer0_outputs(11217) <= not b or a;
    layer0_outputs(11218) <= not a or b;
    layer0_outputs(11219) <= a and not b;
    layer0_outputs(11220) <= a xor b;
    layer0_outputs(11221) <= a and not b;
    layer0_outputs(11222) <= b;
    layer0_outputs(11223) <= not (a and b);
    layer0_outputs(11224) <= '0';
    layer0_outputs(11225) <= a and b;
    layer0_outputs(11226) <= b and not a;
    layer0_outputs(11227) <= '1';
    layer0_outputs(11228) <= a xor b;
    layer0_outputs(11229) <= not b or a;
    layer0_outputs(11230) <= not b;
    layer0_outputs(11231) <= b and not a;
    layer0_outputs(11232) <= a xor b;
    layer0_outputs(11233) <= not (a or b);
    layer0_outputs(11234) <= a and b;
    layer0_outputs(11235) <= a;
    layer0_outputs(11236) <= not b or a;
    layer0_outputs(11237) <= a or b;
    layer0_outputs(11238) <= not a;
    layer0_outputs(11239) <= not (a xor b);
    layer0_outputs(11240) <= a and not b;
    layer0_outputs(11241) <= b;
    layer0_outputs(11242) <= a;
    layer0_outputs(11243) <= a or b;
    layer0_outputs(11244) <= not b or a;
    layer0_outputs(11245) <= a or b;
    layer0_outputs(11246) <= not b;
    layer0_outputs(11247) <= b and not a;
    layer0_outputs(11248) <= a xor b;
    layer0_outputs(11249) <= not (a xor b);
    layer0_outputs(11250) <= not (a and b);
    layer0_outputs(11251) <= not (a xor b);
    layer0_outputs(11252) <= not a or b;
    layer0_outputs(11253) <= a or b;
    layer0_outputs(11254) <= '1';
    layer0_outputs(11255) <= a and b;
    layer0_outputs(11256) <= b;
    layer0_outputs(11257) <= not (a and b);
    layer0_outputs(11258) <= a and b;
    layer0_outputs(11259) <= not b;
    layer0_outputs(11260) <= b and not a;
    layer0_outputs(11261) <= not (a and b);
    layer0_outputs(11262) <= '0';
    layer0_outputs(11263) <= not b;
    layer0_outputs(11264) <= not b or a;
    layer0_outputs(11265) <= not (a or b);
    layer0_outputs(11266) <= a and b;
    layer0_outputs(11267) <= a and b;
    layer0_outputs(11268) <= not b or a;
    layer0_outputs(11269) <= '1';
    layer0_outputs(11270) <= '1';
    layer0_outputs(11271) <= '1';
    layer0_outputs(11272) <= a or b;
    layer0_outputs(11273) <= a and not b;
    layer0_outputs(11274) <= '1';
    layer0_outputs(11275) <= a or b;
    layer0_outputs(11276) <= '0';
    layer0_outputs(11277) <= '1';
    layer0_outputs(11278) <= a xor b;
    layer0_outputs(11279) <= a xor b;
    layer0_outputs(11280) <= not (a xor b);
    layer0_outputs(11281) <= a;
    layer0_outputs(11282) <= not a or b;
    layer0_outputs(11283) <= not a or b;
    layer0_outputs(11284) <= not a;
    layer0_outputs(11285) <= not (a or b);
    layer0_outputs(11286) <= not (a xor b);
    layer0_outputs(11287) <= not (a or b);
    layer0_outputs(11288) <= not b or a;
    layer0_outputs(11289) <= not (a xor b);
    layer0_outputs(11290) <= a;
    layer0_outputs(11291) <= '0';
    layer0_outputs(11292) <= a and not b;
    layer0_outputs(11293) <= a or b;
    layer0_outputs(11294) <= a or b;
    layer0_outputs(11295) <= a and not b;
    layer0_outputs(11296) <= a and not b;
    layer0_outputs(11297) <= a xor b;
    layer0_outputs(11298) <= a or b;
    layer0_outputs(11299) <= a and b;
    layer0_outputs(11300) <= a and b;
    layer0_outputs(11301) <= a or b;
    layer0_outputs(11302) <= a or b;
    layer0_outputs(11303) <= b;
    layer0_outputs(11304) <= a xor b;
    layer0_outputs(11305) <= a and not b;
    layer0_outputs(11306) <= a xor b;
    layer0_outputs(11307) <= not (a and b);
    layer0_outputs(11308) <= b and not a;
    layer0_outputs(11309) <= not (a xor b);
    layer0_outputs(11310) <= '1';
    layer0_outputs(11311) <= a xor b;
    layer0_outputs(11312) <= a and b;
    layer0_outputs(11313) <= '1';
    layer0_outputs(11314) <= a and b;
    layer0_outputs(11315) <= not b or a;
    layer0_outputs(11316) <= not (a or b);
    layer0_outputs(11317) <= not a;
    layer0_outputs(11318) <= not b or a;
    layer0_outputs(11319) <= not b or a;
    layer0_outputs(11320) <= a and b;
    layer0_outputs(11321) <= not (a or b);
    layer0_outputs(11322) <= not a or b;
    layer0_outputs(11323) <= not b or a;
    layer0_outputs(11324) <= b and not a;
    layer0_outputs(11325) <= a or b;
    layer0_outputs(11326) <= a;
    layer0_outputs(11327) <= not b or a;
    layer0_outputs(11328) <= a and not b;
    layer0_outputs(11329) <= a;
    layer0_outputs(11330) <= not a or b;
    layer0_outputs(11331) <= a or b;
    layer0_outputs(11332) <= not b;
    layer0_outputs(11333) <= a or b;
    layer0_outputs(11334) <= not a;
    layer0_outputs(11335) <= a;
    layer0_outputs(11336) <= '1';
    layer0_outputs(11337) <= not b;
    layer0_outputs(11338) <= not (a and b);
    layer0_outputs(11339) <= not (a and b);
    layer0_outputs(11340) <= '0';
    layer0_outputs(11341) <= not b or a;
    layer0_outputs(11342) <= not (a or b);
    layer0_outputs(11343) <= a xor b;
    layer0_outputs(11344) <= '0';
    layer0_outputs(11345) <= not a or b;
    layer0_outputs(11346) <= '1';
    layer0_outputs(11347) <= a;
    layer0_outputs(11348) <= not (a xor b);
    layer0_outputs(11349) <= not a;
    layer0_outputs(11350) <= not b;
    layer0_outputs(11351) <= not b;
    layer0_outputs(11352) <= not b or a;
    layer0_outputs(11353) <= a and b;
    layer0_outputs(11354) <= not (a or b);
    layer0_outputs(11355) <= a and b;
    layer0_outputs(11356) <= a and not b;
    layer0_outputs(11357) <= not b;
    layer0_outputs(11358) <= a and not b;
    layer0_outputs(11359) <= not b;
    layer0_outputs(11360) <= not (a or b);
    layer0_outputs(11361) <= '0';
    layer0_outputs(11362) <= a and not b;
    layer0_outputs(11363) <= a or b;
    layer0_outputs(11364) <= b;
    layer0_outputs(11365) <= a and b;
    layer0_outputs(11366) <= b;
    layer0_outputs(11367) <= b;
    layer0_outputs(11368) <= not (a xor b);
    layer0_outputs(11369) <= '0';
    layer0_outputs(11370) <= a and not b;
    layer0_outputs(11371) <= not (a or b);
    layer0_outputs(11372) <= '0';
    layer0_outputs(11373) <= not b or a;
    layer0_outputs(11374) <= not a or b;
    layer0_outputs(11375) <= not (a or b);
    layer0_outputs(11376) <= not b;
    layer0_outputs(11377) <= not b;
    layer0_outputs(11378) <= a or b;
    layer0_outputs(11379) <= '0';
    layer0_outputs(11380) <= not a or b;
    layer0_outputs(11381) <= not a;
    layer0_outputs(11382) <= not (a or b);
    layer0_outputs(11383) <= '1';
    layer0_outputs(11384) <= a;
    layer0_outputs(11385) <= not (a or b);
    layer0_outputs(11386) <= not b or a;
    layer0_outputs(11387) <= not a or b;
    layer0_outputs(11388) <= a;
    layer0_outputs(11389) <= b;
    layer0_outputs(11390) <= b;
    layer0_outputs(11391) <= not b or a;
    layer0_outputs(11392) <= a and not b;
    layer0_outputs(11393) <= not b or a;
    layer0_outputs(11394) <= a and not b;
    layer0_outputs(11395) <= not (a or b);
    layer0_outputs(11396) <= a xor b;
    layer0_outputs(11397) <= not (a xor b);
    layer0_outputs(11398) <= not a;
    layer0_outputs(11399) <= not (a or b);
    layer0_outputs(11400) <= b;
    layer0_outputs(11401) <= not a or b;
    layer0_outputs(11402) <= not a or b;
    layer0_outputs(11403) <= a or b;
    layer0_outputs(11404) <= not (a and b);
    layer0_outputs(11405) <= not (a xor b);
    layer0_outputs(11406) <= not b or a;
    layer0_outputs(11407) <= b;
    layer0_outputs(11408) <= not (a or b);
    layer0_outputs(11409) <= not b;
    layer0_outputs(11410) <= not (a xor b);
    layer0_outputs(11411) <= not (a xor b);
    layer0_outputs(11412) <= not b;
    layer0_outputs(11413) <= not a;
    layer0_outputs(11414) <= a and not b;
    layer0_outputs(11415) <= not a or b;
    layer0_outputs(11416) <= '0';
    layer0_outputs(11417) <= a or b;
    layer0_outputs(11418) <= not a or b;
    layer0_outputs(11419) <= not b or a;
    layer0_outputs(11420) <= not (a and b);
    layer0_outputs(11421) <= '0';
    layer0_outputs(11422) <= not (a or b);
    layer0_outputs(11423) <= b and not a;
    layer0_outputs(11424) <= not a;
    layer0_outputs(11425) <= not (a or b);
    layer0_outputs(11426) <= a and not b;
    layer0_outputs(11427) <= a;
    layer0_outputs(11428) <= not (a or b);
    layer0_outputs(11429) <= b;
    layer0_outputs(11430) <= a;
    layer0_outputs(11431) <= not (a or b);
    layer0_outputs(11432) <= not (a or b);
    layer0_outputs(11433) <= a xor b;
    layer0_outputs(11434) <= a or b;
    layer0_outputs(11435) <= b;
    layer0_outputs(11436) <= b;
    layer0_outputs(11437) <= b and not a;
    layer0_outputs(11438) <= not b or a;
    layer0_outputs(11439) <= a and b;
    layer0_outputs(11440) <= '0';
    layer0_outputs(11441) <= not (a and b);
    layer0_outputs(11442) <= b;
    layer0_outputs(11443) <= not (a or b);
    layer0_outputs(11444) <= a;
    layer0_outputs(11445) <= not a;
    layer0_outputs(11446) <= not a;
    layer0_outputs(11447) <= a and not b;
    layer0_outputs(11448) <= a or b;
    layer0_outputs(11449) <= not (a or b);
    layer0_outputs(11450) <= '0';
    layer0_outputs(11451) <= a or b;
    layer0_outputs(11452) <= a;
    layer0_outputs(11453) <= b and not a;
    layer0_outputs(11454) <= a and not b;
    layer0_outputs(11455) <= b and not a;
    layer0_outputs(11456) <= a and not b;
    layer0_outputs(11457) <= not (a or b);
    layer0_outputs(11458) <= not (a or b);
    layer0_outputs(11459) <= a or b;
    layer0_outputs(11460) <= a and b;
    layer0_outputs(11461) <= not (a or b);
    layer0_outputs(11462) <= b;
    layer0_outputs(11463) <= not a;
    layer0_outputs(11464) <= a and not b;
    layer0_outputs(11465) <= b;
    layer0_outputs(11466) <= a;
    layer0_outputs(11467) <= not b or a;
    layer0_outputs(11468) <= not b or a;
    layer0_outputs(11469) <= b;
    layer0_outputs(11470) <= b;
    layer0_outputs(11471) <= a;
    layer0_outputs(11472) <= not b;
    layer0_outputs(11473) <= b and not a;
    layer0_outputs(11474) <= a xor b;
    layer0_outputs(11475) <= not (a or b);
    layer0_outputs(11476) <= a and not b;
    layer0_outputs(11477) <= a and not b;
    layer0_outputs(11478) <= a and not b;
    layer0_outputs(11479) <= b and not a;
    layer0_outputs(11480) <= not (a and b);
    layer0_outputs(11481) <= not a;
    layer0_outputs(11482) <= b and not a;
    layer0_outputs(11483) <= not a or b;
    layer0_outputs(11484) <= not a;
    layer0_outputs(11485) <= b;
    layer0_outputs(11486) <= a xor b;
    layer0_outputs(11487) <= a xor b;
    layer0_outputs(11488) <= a xor b;
    layer0_outputs(11489) <= b and not a;
    layer0_outputs(11490) <= not (a and b);
    layer0_outputs(11491) <= a and b;
    layer0_outputs(11492) <= a and b;
    layer0_outputs(11493) <= a xor b;
    layer0_outputs(11494) <= not b or a;
    layer0_outputs(11495) <= a or b;
    layer0_outputs(11496) <= not a or b;
    layer0_outputs(11497) <= not (a or b);
    layer0_outputs(11498) <= not (a or b);
    layer0_outputs(11499) <= '1';
    layer0_outputs(11500) <= not b;
    layer0_outputs(11501) <= not (a or b);
    layer0_outputs(11502) <= a and b;
    layer0_outputs(11503) <= a or b;
    layer0_outputs(11504) <= not (a or b);
    layer0_outputs(11505) <= '1';
    layer0_outputs(11506) <= not b;
    layer0_outputs(11507) <= a and b;
    layer0_outputs(11508) <= '1';
    layer0_outputs(11509) <= b;
    layer0_outputs(11510) <= not (a and b);
    layer0_outputs(11511) <= b;
    layer0_outputs(11512) <= a;
    layer0_outputs(11513) <= not (a xor b);
    layer0_outputs(11514) <= not (a xor b);
    layer0_outputs(11515) <= not (a or b);
    layer0_outputs(11516) <= not a;
    layer0_outputs(11517) <= '0';
    layer0_outputs(11518) <= not a;
    layer0_outputs(11519) <= b;
    layer0_outputs(11520) <= '1';
    layer0_outputs(11521) <= not (a or b);
    layer0_outputs(11522) <= not (a or b);
    layer0_outputs(11523) <= not b or a;
    layer0_outputs(11524) <= not a or b;
    layer0_outputs(11525) <= '1';
    layer0_outputs(11526) <= a and not b;
    layer0_outputs(11527) <= not a;
    layer0_outputs(11528) <= '1';
    layer0_outputs(11529) <= a and not b;
    layer0_outputs(11530) <= not (a xor b);
    layer0_outputs(11531) <= a and not b;
    layer0_outputs(11532) <= a and not b;
    layer0_outputs(11533) <= a and not b;
    layer0_outputs(11534) <= not a or b;
    layer0_outputs(11535) <= a;
    layer0_outputs(11536) <= not a or b;
    layer0_outputs(11537) <= b and not a;
    layer0_outputs(11538) <= not b or a;
    layer0_outputs(11539) <= not a or b;
    layer0_outputs(11540) <= a and b;
    layer0_outputs(11541) <= a or b;
    layer0_outputs(11542) <= a or b;
    layer0_outputs(11543) <= a xor b;
    layer0_outputs(11544) <= not a or b;
    layer0_outputs(11545) <= a and b;
    layer0_outputs(11546) <= a xor b;
    layer0_outputs(11547) <= not a or b;
    layer0_outputs(11548) <= b and not a;
    layer0_outputs(11549) <= b and not a;
    layer0_outputs(11550) <= not a;
    layer0_outputs(11551) <= a;
    layer0_outputs(11552) <= not (a or b);
    layer0_outputs(11553) <= not (a xor b);
    layer0_outputs(11554) <= b;
    layer0_outputs(11555) <= a xor b;
    layer0_outputs(11556) <= a;
    layer0_outputs(11557) <= not a or b;
    layer0_outputs(11558) <= not (a or b);
    layer0_outputs(11559) <= not a;
    layer0_outputs(11560) <= b;
    layer0_outputs(11561) <= not a or b;
    layer0_outputs(11562) <= not a or b;
    layer0_outputs(11563) <= not a;
    layer0_outputs(11564) <= a or b;
    layer0_outputs(11565) <= b;
    layer0_outputs(11566) <= a and not b;
    layer0_outputs(11567) <= b and not a;
    layer0_outputs(11568) <= not b or a;
    layer0_outputs(11569) <= not (a or b);
    layer0_outputs(11570) <= '1';
    layer0_outputs(11571) <= b and not a;
    layer0_outputs(11572) <= b;
    layer0_outputs(11573) <= b;
    layer0_outputs(11574) <= b;
    layer0_outputs(11575) <= not a or b;
    layer0_outputs(11576) <= '1';
    layer0_outputs(11577) <= not (a xor b);
    layer0_outputs(11578) <= a and b;
    layer0_outputs(11579) <= a or b;
    layer0_outputs(11580) <= a;
    layer0_outputs(11581) <= b;
    layer0_outputs(11582) <= a and b;
    layer0_outputs(11583) <= b;
    layer0_outputs(11584) <= a or b;
    layer0_outputs(11585) <= '1';
    layer0_outputs(11586) <= not b or a;
    layer0_outputs(11587) <= a and not b;
    layer0_outputs(11588) <= not (a and b);
    layer0_outputs(11589) <= b;
    layer0_outputs(11590) <= not a;
    layer0_outputs(11591) <= '0';
    layer0_outputs(11592) <= a or b;
    layer0_outputs(11593) <= a and not b;
    layer0_outputs(11594) <= a and not b;
    layer0_outputs(11595) <= not a;
    layer0_outputs(11596) <= '0';
    layer0_outputs(11597) <= not b;
    layer0_outputs(11598) <= not a;
    layer0_outputs(11599) <= not (a and b);
    layer0_outputs(11600) <= '1';
    layer0_outputs(11601) <= not a;
    layer0_outputs(11602) <= not (a and b);
    layer0_outputs(11603) <= '0';
    layer0_outputs(11604) <= not (a or b);
    layer0_outputs(11605) <= not a or b;
    layer0_outputs(11606) <= not b;
    layer0_outputs(11607) <= not b or a;
    layer0_outputs(11608) <= '1';
    layer0_outputs(11609) <= not a;
    layer0_outputs(11610) <= b;
    layer0_outputs(11611) <= b and not a;
    layer0_outputs(11612) <= not a or b;
    layer0_outputs(11613) <= '1';
    layer0_outputs(11614) <= not b or a;
    layer0_outputs(11615) <= a;
    layer0_outputs(11616) <= not (a xor b);
    layer0_outputs(11617) <= not a or b;
    layer0_outputs(11618) <= a and not b;
    layer0_outputs(11619) <= '1';
    layer0_outputs(11620) <= b;
    layer0_outputs(11621) <= a and b;
    layer0_outputs(11622) <= '0';
    layer0_outputs(11623) <= not b;
    layer0_outputs(11624) <= not (a and b);
    layer0_outputs(11625) <= b and not a;
    layer0_outputs(11626) <= not a;
    layer0_outputs(11627) <= not (a xor b);
    layer0_outputs(11628) <= a or b;
    layer0_outputs(11629) <= a;
    layer0_outputs(11630) <= b;
    layer0_outputs(11631) <= a;
    layer0_outputs(11632) <= not b;
    layer0_outputs(11633) <= b and not a;
    layer0_outputs(11634) <= b;
    layer0_outputs(11635) <= not (a and b);
    layer0_outputs(11636) <= not b;
    layer0_outputs(11637) <= not b;
    layer0_outputs(11638) <= not a;
    layer0_outputs(11639) <= not b;
    layer0_outputs(11640) <= not a or b;
    layer0_outputs(11641) <= a xor b;
    layer0_outputs(11642) <= '0';
    layer0_outputs(11643) <= '0';
    layer0_outputs(11644) <= not (a or b);
    layer0_outputs(11645) <= a and not b;
    layer0_outputs(11646) <= a xor b;
    layer0_outputs(11647) <= not a;
    layer0_outputs(11648) <= not b;
    layer0_outputs(11649) <= a and b;
    layer0_outputs(11650) <= a;
    layer0_outputs(11651) <= '0';
    layer0_outputs(11652) <= not b;
    layer0_outputs(11653) <= b;
    layer0_outputs(11654) <= not (a xor b);
    layer0_outputs(11655) <= not b or a;
    layer0_outputs(11656) <= a and not b;
    layer0_outputs(11657) <= a or b;
    layer0_outputs(11658) <= '1';
    layer0_outputs(11659) <= '1';
    layer0_outputs(11660) <= '1';
    layer0_outputs(11661) <= not (a and b);
    layer0_outputs(11662) <= '1';
    layer0_outputs(11663) <= not a;
    layer0_outputs(11664) <= not (a or b);
    layer0_outputs(11665) <= not (a or b);
    layer0_outputs(11666) <= not b or a;
    layer0_outputs(11667) <= '1';
    layer0_outputs(11668) <= not b or a;
    layer0_outputs(11669) <= b and not a;
    layer0_outputs(11670) <= a xor b;
    layer0_outputs(11671) <= '0';
    layer0_outputs(11672) <= '1';
    layer0_outputs(11673) <= a xor b;
    layer0_outputs(11674) <= not a;
    layer0_outputs(11675) <= a;
    layer0_outputs(11676) <= a and b;
    layer0_outputs(11677) <= not (a xor b);
    layer0_outputs(11678) <= '0';
    layer0_outputs(11679) <= b;
    layer0_outputs(11680) <= a;
    layer0_outputs(11681) <= a;
    layer0_outputs(11682) <= '1';
    layer0_outputs(11683) <= not a or b;
    layer0_outputs(11684) <= a xor b;
    layer0_outputs(11685) <= not (a or b);
    layer0_outputs(11686) <= a and b;
    layer0_outputs(11687) <= not b;
    layer0_outputs(11688) <= not a;
    layer0_outputs(11689) <= b;
    layer0_outputs(11690) <= not (a xor b);
    layer0_outputs(11691) <= not (a xor b);
    layer0_outputs(11692) <= not (a or b);
    layer0_outputs(11693) <= '1';
    layer0_outputs(11694) <= a and not b;
    layer0_outputs(11695) <= not a or b;
    layer0_outputs(11696) <= a or b;
    layer0_outputs(11697) <= b and not a;
    layer0_outputs(11698) <= not a or b;
    layer0_outputs(11699) <= not b;
    layer0_outputs(11700) <= not a or b;
    layer0_outputs(11701) <= not a;
    layer0_outputs(11702) <= a or b;
    layer0_outputs(11703) <= not b or a;
    layer0_outputs(11704) <= a and not b;
    layer0_outputs(11705) <= b;
    layer0_outputs(11706) <= not b or a;
    layer0_outputs(11707) <= a and not b;
    layer0_outputs(11708) <= not (a or b);
    layer0_outputs(11709) <= not b;
    layer0_outputs(11710) <= not (a xor b);
    layer0_outputs(11711) <= a or b;
    layer0_outputs(11712) <= not (a xor b);
    layer0_outputs(11713) <= b and not a;
    layer0_outputs(11714) <= not (a xor b);
    layer0_outputs(11715) <= not b or a;
    layer0_outputs(11716) <= b;
    layer0_outputs(11717) <= '1';
    layer0_outputs(11718) <= a or b;
    layer0_outputs(11719) <= not b or a;
    layer0_outputs(11720) <= a;
    layer0_outputs(11721) <= a and not b;
    layer0_outputs(11722) <= a or b;
    layer0_outputs(11723) <= not (a and b);
    layer0_outputs(11724) <= not b;
    layer0_outputs(11725) <= b;
    layer0_outputs(11726) <= not (a or b);
    layer0_outputs(11727) <= not a or b;
    layer0_outputs(11728) <= not (a or b);
    layer0_outputs(11729) <= not b;
    layer0_outputs(11730) <= a;
    layer0_outputs(11731) <= not a or b;
    layer0_outputs(11732) <= a;
    layer0_outputs(11733) <= b;
    layer0_outputs(11734) <= b and not a;
    layer0_outputs(11735) <= not (a and b);
    layer0_outputs(11736) <= not (a and b);
    layer0_outputs(11737) <= a xor b;
    layer0_outputs(11738) <= not a or b;
    layer0_outputs(11739) <= '0';
    layer0_outputs(11740) <= not (a xor b);
    layer0_outputs(11741) <= not (a and b);
    layer0_outputs(11742) <= '1';
    layer0_outputs(11743) <= b;
    layer0_outputs(11744) <= '0';
    layer0_outputs(11745) <= a and not b;
    layer0_outputs(11746) <= b and not a;
    layer0_outputs(11747) <= not (a or b);
    layer0_outputs(11748) <= not a;
    layer0_outputs(11749) <= not a or b;
    layer0_outputs(11750) <= not a;
    layer0_outputs(11751) <= a and b;
    layer0_outputs(11752) <= b and not a;
    layer0_outputs(11753) <= a xor b;
    layer0_outputs(11754) <= not a or b;
    layer0_outputs(11755) <= a xor b;
    layer0_outputs(11756) <= a or b;
    layer0_outputs(11757) <= not b;
    layer0_outputs(11758) <= a and b;
    layer0_outputs(11759) <= a or b;
    layer0_outputs(11760) <= b;
    layer0_outputs(11761) <= a xor b;
    layer0_outputs(11762) <= a xor b;
    layer0_outputs(11763) <= not b;
    layer0_outputs(11764) <= a and not b;
    layer0_outputs(11765) <= b and not a;
    layer0_outputs(11766) <= b;
    layer0_outputs(11767) <= a or b;
    layer0_outputs(11768) <= b;
    layer0_outputs(11769) <= not b or a;
    layer0_outputs(11770) <= not a or b;
    layer0_outputs(11771) <= a and not b;
    layer0_outputs(11772) <= not a or b;
    layer0_outputs(11773) <= not b or a;
    layer0_outputs(11774) <= not a or b;
    layer0_outputs(11775) <= '0';
    layer0_outputs(11776) <= a and not b;
    layer0_outputs(11777) <= not (a xor b);
    layer0_outputs(11778) <= a or b;
    layer0_outputs(11779) <= '1';
    layer0_outputs(11780) <= b;
    layer0_outputs(11781) <= not b or a;
    layer0_outputs(11782) <= b;
    layer0_outputs(11783) <= '0';
    layer0_outputs(11784) <= a and b;
    layer0_outputs(11785) <= b;
    layer0_outputs(11786) <= a;
    layer0_outputs(11787) <= not (a xor b);
    layer0_outputs(11788) <= not (a and b);
    layer0_outputs(11789) <= not (a or b);
    layer0_outputs(11790) <= not a or b;
    layer0_outputs(11791) <= a or b;
    layer0_outputs(11792) <= a;
    layer0_outputs(11793) <= '1';
    layer0_outputs(11794) <= not a or b;
    layer0_outputs(11795) <= a and b;
    layer0_outputs(11796) <= b and not a;
    layer0_outputs(11797) <= not b or a;
    layer0_outputs(11798) <= b and not a;
    layer0_outputs(11799) <= b;
    layer0_outputs(11800) <= a or b;
    layer0_outputs(11801) <= a and b;
    layer0_outputs(11802) <= not a or b;
    layer0_outputs(11803) <= a or b;
    layer0_outputs(11804) <= not (a and b);
    layer0_outputs(11805) <= b and not a;
    layer0_outputs(11806) <= not a or b;
    layer0_outputs(11807) <= a xor b;
    layer0_outputs(11808) <= a or b;
    layer0_outputs(11809) <= not (a and b);
    layer0_outputs(11810) <= not b;
    layer0_outputs(11811) <= a and not b;
    layer0_outputs(11812) <= not a;
    layer0_outputs(11813) <= b and not a;
    layer0_outputs(11814) <= a or b;
    layer0_outputs(11815) <= a and not b;
    layer0_outputs(11816) <= not a;
    layer0_outputs(11817) <= not (a or b);
    layer0_outputs(11818) <= not (a and b);
    layer0_outputs(11819) <= not a or b;
    layer0_outputs(11820) <= not b or a;
    layer0_outputs(11821) <= '1';
    layer0_outputs(11822) <= not (a or b);
    layer0_outputs(11823) <= not (a or b);
    layer0_outputs(11824) <= a and not b;
    layer0_outputs(11825) <= not b;
    layer0_outputs(11826) <= not b;
    layer0_outputs(11827) <= a xor b;
    layer0_outputs(11828) <= not a;
    layer0_outputs(11829) <= '1';
    layer0_outputs(11830) <= not (a and b);
    layer0_outputs(11831) <= b and not a;
    layer0_outputs(11832) <= a and b;
    layer0_outputs(11833) <= not a;
    layer0_outputs(11834) <= b and not a;
    layer0_outputs(11835) <= a and not b;
    layer0_outputs(11836) <= a xor b;
    layer0_outputs(11837) <= not a;
    layer0_outputs(11838) <= not b or a;
    layer0_outputs(11839) <= not b;
    layer0_outputs(11840) <= not (a xor b);
    layer0_outputs(11841) <= not (a or b);
    layer0_outputs(11842) <= b;
    layer0_outputs(11843) <= not (a and b);
    layer0_outputs(11844) <= a or b;
    layer0_outputs(11845) <= not (a and b);
    layer0_outputs(11846) <= not (a xor b);
    layer0_outputs(11847) <= not (a and b);
    layer0_outputs(11848) <= not b or a;
    layer0_outputs(11849) <= not b or a;
    layer0_outputs(11850) <= not (a or b);
    layer0_outputs(11851) <= not b or a;
    layer0_outputs(11852) <= a and b;
    layer0_outputs(11853) <= not (a xor b);
    layer0_outputs(11854) <= '1';
    layer0_outputs(11855) <= a and not b;
    layer0_outputs(11856) <= not b or a;
    layer0_outputs(11857) <= b;
    layer0_outputs(11858) <= not (a or b);
    layer0_outputs(11859) <= a and b;
    layer0_outputs(11860) <= not a or b;
    layer0_outputs(11861) <= a and b;
    layer0_outputs(11862) <= not (a and b);
    layer0_outputs(11863) <= not b or a;
    layer0_outputs(11864) <= not (a xor b);
    layer0_outputs(11865) <= not b or a;
    layer0_outputs(11866) <= a or b;
    layer0_outputs(11867) <= a and not b;
    layer0_outputs(11868) <= not (a xor b);
    layer0_outputs(11869) <= '1';
    layer0_outputs(11870) <= not b or a;
    layer0_outputs(11871) <= b;
    layer0_outputs(11872) <= a and not b;
    layer0_outputs(11873) <= a and b;
    layer0_outputs(11874) <= a or b;
    layer0_outputs(11875) <= not b;
    layer0_outputs(11876) <= a xor b;
    layer0_outputs(11877) <= a xor b;
    layer0_outputs(11878) <= a xor b;
    layer0_outputs(11879) <= not (a xor b);
    layer0_outputs(11880) <= not b;
    layer0_outputs(11881) <= a and b;
    layer0_outputs(11882) <= not b;
    layer0_outputs(11883) <= not a or b;
    layer0_outputs(11884) <= a;
    layer0_outputs(11885) <= a xor b;
    layer0_outputs(11886) <= not b;
    layer0_outputs(11887) <= not a;
    layer0_outputs(11888) <= a;
    layer0_outputs(11889) <= '0';
    layer0_outputs(11890) <= a and b;
    layer0_outputs(11891) <= a and b;
    layer0_outputs(11892) <= '1';
    layer0_outputs(11893) <= a;
    layer0_outputs(11894) <= not (a and b);
    layer0_outputs(11895) <= not a or b;
    layer0_outputs(11896) <= b;
    layer0_outputs(11897) <= not (a xor b);
    layer0_outputs(11898) <= b;
    layer0_outputs(11899) <= a or b;
    layer0_outputs(11900) <= a and b;
    layer0_outputs(11901) <= a and not b;
    layer0_outputs(11902) <= not (a and b);
    layer0_outputs(11903) <= a xor b;
    layer0_outputs(11904) <= a xor b;
    layer0_outputs(11905) <= not a;
    layer0_outputs(11906) <= a and not b;
    layer0_outputs(11907) <= not b or a;
    layer0_outputs(11908) <= not a;
    layer0_outputs(11909) <= not b or a;
    layer0_outputs(11910) <= b and not a;
    layer0_outputs(11911) <= '0';
    layer0_outputs(11912) <= a and b;
    layer0_outputs(11913) <= not b;
    layer0_outputs(11914) <= not a;
    layer0_outputs(11915) <= a and not b;
    layer0_outputs(11916) <= b;
    layer0_outputs(11917) <= '0';
    layer0_outputs(11918) <= not (a or b);
    layer0_outputs(11919) <= not b or a;
    layer0_outputs(11920) <= not a or b;
    layer0_outputs(11921) <= not b;
    layer0_outputs(11922) <= b and not a;
    layer0_outputs(11923) <= b;
    layer0_outputs(11924) <= a;
    layer0_outputs(11925) <= a;
    layer0_outputs(11926) <= not b;
    layer0_outputs(11927) <= b and not a;
    layer0_outputs(11928) <= a and b;
    layer0_outputs(11929) <= b;
    layer0_outputs(11930) <= b and not a;
    layer0_outputs(11931) <= a and not b;
    layer0_outputs(11932) <= a or b;
    layer0_outputs(11933) <= a and not b;
    layer0_outputs(11934) <= a xor b;
    layer0_outputs(11935) <= not a or b;
    layer0_outputs(11936) <= not (a xor b);
    layer0_outputs(11937) <= a and not b;
    layer0_outputs(11938) <= '1';
    layer0_outputs(11939) <= not a or b;
    layer0_outputs(11940) <= not (a or b);
    layer0_outputs(11941) <= a or b;
    layer0_outputs(11942) <= '1';
    layer0_outputs(11943) <= not (a or b);
    layer0_outputs(11944) <= '0';
    layer0_outputs(11945) <= not a;
    layer0_outputs(11946) <= a and not b;
    layer0_outputs(11947) <= b and not a;
    layer0_outputs(11948) <= '1';
    layer0_outputs(11949) <= b and not a;
    layer0_outputs(11950) <= a or b;
    layer0_outputs(11951) <= '0';
    layer0_outputs(11952) <= a xor b;
    layer0_outputs(11953) <= not a or b;
    layer0_outputs(11954) <= '1';
    layer0_outputs(11955) <= b;
    layer0_outputs(11956) <= not (a and b);
    layer0_outputs(11957) <= not a or b;
    layer0_outputs(11958) <= not (a or b);
    layer0_outputs(11959) <= a xor b;
    layer0_outputs(11960) <= a or b;
    layer0_outputs(11961) <= not b or a;
    layer0_outputs(11962) <= b and not a;
    layer0_outputs(11963) <= not (a and b);
    layer0_outputs(11964) <= b;
    layer0_outputs(11965) <= a or b;
    layer0_outputs(11966) <= not b;
    layer0_outputs(11967) <= a and not b;
    layer0_outputs(11968) <= not (a or b);
    layer0_outputs(11969) <= '1';
    layer0_outputs(11970) <= not (a xor b);
    layer0_outputs(11971) <= not (a xor b);
    layer0_outputs(11972) <= not a;
    layer0_outputs(11973) <= a and b;
    layer0_outputs(11974) <= a and not b;
    layer0_outputs(11975) <= not a;
    layer0_outputs(11976) <= not (a or b);
    layer0_outputs(11977) <= a or b;
    layer0_outputs(11978) <= not (a or b);
    layer0_outputs(11979) <= not (a or b);
    layer0_outputs(11980) <= not b or a;
    layer0_outputs(11981) <= a or b;
    layer0_outputs(11982) <= a or b;
    layer0_outputs(11983) <= a or b;
    layer0_outputs(11984) <= a or b;
    layer0_outputs(11985) <= b;
    layer0_outputs(11986) <= a and not b;
    layer0_outputs(11987) <= a and not b;
    layer0_outputs(11988) <= not (a xor b);
    layer0_outputs(11989) <= not b;
    layer0_outputs(11990) <= not (a or b);
    layer0_outputs(11991) <= not (a or b);
    layer0_outputs(11992) <= not a;
    layer0_outputs(11993) <= b;
    layer0_outputs(11994) <= not b or a;
    layer0_outputs(11995) <= a xor b;
    layer0_outputs(11996) <= a;
    layer0_outputs(11997) <= a;
    layer0_outputs(11998) <= '0';
    layer0_outputs(11999) <= not a or b;
    layer0_outputs(12000) <= not (a and b);
    layer0_outputs(12001) <= a or b;
    layer0_outputs(12002) <= not (a or b);
    layer0_outputs(12003) <= a;
    layer0_outputs(12004) <= a and b;
    layer0_outputs(12005) <= a and not b;
    layer0_outputs(12006) <= a;
    layer0_outputs(12007) <= not a or b;
    layer0_outputs(12008) <= '1';
    layer0_outputs(12009) <= b;
    layer0_outputs(12010) <= not a or b;
    layer0_outputs(12011) <= b;
    layer0_outputs(12012) <= not a;
    layer0_outputs(12013) <= not b;
    layer0_outputs(12014) <= a;
    layer0_outputs(12015) <= a xor b;
    layer0_outputs(12016) <= a xor b;
    layer0_outputs(12017) <= not (a or b);
    layer0_outputs(12018) <= not (a xor b);
    layer0_outputs(12019) <= a xor b;
    layer0_outputs(12020) <= b;
    layer0_outputs(12021) <= a and b;
    layer0_outputs(12022) <= not b or a;
    layer0_outputs(12023) <= a;
    layer0_outputs(12024) <= not b;
    layer0_outputs(12025) <= a;
    layer0_outputs(12026) <= not (a xor b);
    layer0_outputs(12027) <= not a;
    layer0_outputs(12028) <= a or b;
    layer0_outputs(12029) <= b and not a;
    layer0_outputs(12030) <= not (a or b);
    layer0_outputs(12031) <= b;
    layer0_outputs(12032) <= not (a or b);
    layer0_outputs(12033) <= a and not b;
    layer0_outputs(12034) <= a;
    layer0_outputs(12035) <= a xor b;
    layer0_outputs(12036) <= a and b;
    layer0_outputs(12037) <= not a or b;
    layer0_outputs(12038) <= not a;
    layer0_outputs(12039) <= a xor b;
    layer0_outputs(12040) <= not a;
    layer0_outputs(12041) <= not (a or b);
    layer0_outputs(12042) <= a;
    layer0_outputs(12043) <= not a or b;
    layer0_outputs(12044) <= not b;
    layer0_outputs(12045) <= not (a xor b);
    layer0_outputs(12046) <= b and not a;
    layer0_outputs(12047) <= a or b;
    layer0_outputs(12048) <= a xor b;
    layer0_outputs(12049) <= not (a xor b);
    layer0_outputs(12050) <= a;
    layer0_outputs(12051) <= not (a or b);
    layer0_outputs(12052) <= not (a or b);
    layer0_outputs(12053) <= a;
    layer0_outputs(12054) <= not (a or b);
    layer0_outputs(12055) <= a or b;
    layer0_outputs(12056) <= a xor b;
    layer0_outputs(12057) <= not a;
    layer0_outputs(12058) <= not a;
    layer0_outputs(12059) <= not a;
    layer0_outputs(12060) <= not (a and b);
    layer0_outputs(12061) <= not a or b;
    layer0_outputs(12062) <= a or b;
    layer0_outputs(12063) <= '0';
    layer0_outputs(12064) <= a;
    layer0_outputs(12065) <= a;
    layer0_outputs(12066) <= a xor b;
    layer0_outputs(12067) <= '0';
    layer0_outputs(12068) <= not (a xor b);
    layer0_outputs(12069) <= not (a or b);
    layer0_outputs(12070) <= not (a xor b);
    layer0_outputs(12071) <= a and not b;
    layer0_outputs(12072) <= '1';
    layer0_outputs(12073) <= a;
    layer0_outputs(12074) <= b and not a;
    layer0_outputs(12075) <= not (a xor b);
    layer0_outputs(12076) <= not b;
    layer0_outputs(12077) <= not (a and b);
    layer0_outputs(12078) <= a;
    layer0_outputs(12079) <= b and not a;
    layer0_outputs(12080) <= b;
    layer0_outputs(12081) <= not b;
    layer0_outputs(12082) <= not b or a;
    layer0_outputs(12083) <= not (a xor b);
    layer0_outputs(12084) <= not b;
    layer0_outputs(12085) <= a xor b;
    layer0_outputs(12086) <= not (a xor b);
    layer0_outputs(12087) <= not a or b;
    layer0_outputs(12088) <= b and not a;
    layer0_outputs(12089) <= not b;
    layer0_outputs(12090) <= a;
    layer0_outputs(12091) <= not b;
    layer0_outputs(12092) <= b and not a;
    layer0_outputs(12093) <= b;
    layer0_outputs(12094) <= not (a and b);
    layer0_outputs(12095) <= not (a or b);
    layer0_outputs(12096) <= '0';
    layer0_outputs(12097) <= b and not a;
    layer0_outputs(12098) <= a and not b;
    layer0_outputs(12099) <= not (a xor b);
    layer0_outputs(12100) <= b;
    layer0_outputs(12101) <= a xor b;
    layer0_outputs(12102) <= a;
    layer0_outputs(12103) <= not (a and b);
    layer0_outputs(12104) <= not b;
    layer0_outputs(12105) <= not b or a;
    layer0_outputs(12106) <= not a or b;
    layer0_outputs(12107) <= not a or b;
    layer0_outputs(12108) <= b and not a;
    layer0_outputs(12109) <= not (a xor b);
    layer0_outputs(12110) <= '1';
    layer0_outputs(12111) <= not b or a;
    layer0_outputs(12112) <= a;
    layer0_outputs(12113) <= a or b;
    layer0_outputs(12114) <= a and not b;
    layer0_outputs(12115) <= not b;
    layer0_outputs(12116) <= not b;
    layer0_outputs(12117) <= not a;
    layer0_outputs(12118) <= b;
    layer0_outputs(12119) <= b and not a;
    layer0_outputs(12120) <= a;
    layer0_outputs(12121) <= a;
    layer0_outputs(12122) <= not a;
    layer0_outputs(12123) <= b;
    layer0_outputs(12124) <= '1';
    layer0_outputs(12125) <= a or b;
    layer0_outputs(12126) <= a or b;
    layer0_outputs(12127) <= '0';
    layer0_outputs(12128) <= not (a or b);
    layer0_outputs(12129) <= a xor b;
    layer0_outputs(12130) <= a xor b;
    layer0_outputs(12131) <= '0';
    layer0_outputs(12132) <= b and not a;
    layer0_outputs(12133) <= not (a or b);
    layer0_outputs(12134) <= not b;
    layer0_outputs(12135) <= a;
    layer0_outputs(12136) <= not (a xor b);
    layer0_outputs(12137) <= not b;
    layer0_outputs(12138) <= '1';
    layer0_outputs(12139) <= not b;
    layer0_outputs(12140) <= not b or a;
    layer0_outputs(12141) <= a xor b;
    layer0_outputs(12142) <= a or b;
    layer0_outputs(12143) <= a;
    layer0_outputs(12144) <= b and not a;
    layer0_outputs(12145) <= not (a xor b);
    layer0_outputs(12146) <= not (a or b);
    layer0_outputs(12147) <= '0';
    layer0_outputs(12148) <= a;
    layer0_outputs(12149) <= not a;
    layer0_outputs(12150) <= '0';
    layer0_outputs(12151) <= not (a and b);
    layer0_outputs(12152) <= not a or b;
    layer0_outputs(12153) <= a xor b;
    layer0_outputs(12154) <= a;
    layer0_outputs(12155) <= not a;
    layer0_outputs(12156) <= not b or a;
    layer0_outputs(12157) <= a or b;
    layer0_outputs(12158) <= not (a xor b);
    layer0_outputs(12159) <= not a or b;
    layer0_outputs(12160) <= '1';
    layer0_outputs(12161) <= not a;
    layer0_outputs(12162) <= not b or a;
    layer0_outputs(12163) <= not b or a;
    layer0_outputs(12164) <= not (a or b);
    layer0_outputs(12165) <= not b;
    layer0_outputs(12166) <= not a or b;
    layer0_outputs(12167) <= a;
    layer0_outputs(12168) <= not (a or b);
    layer0_outputs(12169) <= not (a or b);
    layer0_outputs(12170) <= '0';
    layer0_outputs(12171) <= not (a or b);
    layer0_outputs(12172) <= b;
    layer0_outputs(12173) <= b;
    layer0_outputs(12174) <= a or b;
    layer0_outputs(12175) <= not a or b;
    layer0_outputs(12176) <= '0';
    layer0_outputs(12177) <= not b;
    layer0_outputs(12178) <= not b or a;
    layer0_outputs(12179) <= a and not b;
    layer0_outputs(12180) <= not a or b;
    layer0_outputs(12181) <= a or b;
    layer0_outputs(12182) <= a and b;
    layer0_outputs(12183) <= not b or a;
    layer0_outputs(12184) <= a;
    layer0_outputs(12185) <= not (a or b);
    layer0_outputs(12186) <= '0';
    layer0_outputs(12187) <= a or b;
    layer0_outputs(12188) <= not (a or b);
    layer0_outputs(12189) <= not (a or b);
    layer0_outputs(12190) <= not a;
    layer0_outputs(12191) <= not a or b;
    layer0_outputs(12192) <= not b or a;
    layer0_outputs(12193) <= not a;
    layer0_outputs(12194) <= not a or b;
    layer0_outputs(12195) <= not a or b;
    layer0_outputs(12196) <= not (a or b);
    layer0_outputs(12197) <= '1';
    layer0_outputs(12198) <= a;
    layer0_outputs(12199) <= '1';
    layer0_outputs(12200) <= a or b;
    layer0_outputs(12201) <= a;
    layer0_outputs(12202) <= not b;
    layer0_outputs(12203) <= not b or a;
    layer0_outputs(12204) <= not (a or b);
    layer0_outputs(12205) <= b;
    layer0_outputs(12206) <= not a;
    layer0_outputs(12207) <= not b or a;
    layer0_outputs(12208) <= a and b;
    layer0_outputs(12209) <= a xor b;
    layer0_outputs(12210) <= a;
    layer0_outputs(12211) <= b;
    layer0_outputs(12212) <= not b or a;
    layer0_outputs(12213) <= '1';
    layer0_outputs(12214) <= a or b;
    layer0_outputs(12215) <= a;
    layer0_outputs(12216) <= b and not a;
    layer0_outputs(12217) <= a and not b;
    layer0_outputs(12218) <= a;
    layer0_outputs(12219) <= a and not b;
    layer0_outputs(12220) <= not a;
    layer0_outputs(12221) <= '1';
    layer0_outputs(12222) <= a xor b;
    layer0_outputs(12223) <= '0';
    layer0_outputs(12224) <= a xor b;
    layer0_outputs(12225) <= not a or b;
    layer0_outputs(12226) <= not a or b;
    layer0_outputs(12227) <= not b;
    layer0_outputs(12228) <= '0';
    layer0_outputs(12229) <= not (a and b);
    layer0_outputs(12230) <= '1';
    layer0_outputs(12231) <= '0';
    layer0_outputs(12232) <= not (a or b);
    layer0_outputs(12233) <= a and b;
    layer0_outputs(12234) <= not b or a;
    layer0_outputs(12235) <= b;
    layer0_outputs(12236) <= not a or b;
    layer0_outputs(12237) <= a and not b;
    layer0_outputs(12238) <= not (a xor b);
    layer0_outputs(12239) <= not (a or b);
    layer0_outputs(12240) <= a and not b;
    layer0_outputs(12241) <= not (a xor b);
    layer0_outputs(12242) <= a or b;
    layer0_outputs(12243) <= not (a or b);
    layer0_outputs(12244) <= not (a xor b);
    layer0_outputs(12245) <= a and not b;
    layer0_outputs(12246) <= not b or a;
    layer0_outputs(12247) <= not (a xor b);
    layer0_outputs(12248) <= not b or a;
    layer0_outputs(12249) <= a or b;
    layer0_outputs(12250) <= not (a xor b);
    layer0_outputs(12251) <= b and not a;
    layer0_outputs(12252) <= not (a and b);
    layer0_outputs(12253) <= a and b;
    layer0_outputs(12254) <= a and not b;
    layer0_outputs(12255) <= not a;
    layer0_outputs(12256) <= b and not a;
    layer0_outputs(12257) <= not a;
    layer0_outputs(12258) <= not (a or b);
    layer0_outputs(12259) <= a and not b;
    layer0_outputs(12260) <= a or b;
    layer0_outputs(12261) <= b;
    layer0_outputs(12262) <= a or b;
    layer0_outputs(12263) <= not (a or b);
    layer0_outputs(12264) <= a;
    layer0_outputs(12265) <= not (a xor b);
    layer0_outputs(12266) <= not a;
    layer0_outputs(12267) <= not b;
    layer0_outputs(12268) <= not (a and b);
    layer0_outputs(12269) <= '0';
    layer0_outputs(12270) <= not b;
    layer0_outputs(12271) <= not (a or b);
    layer0_outputs(12272) <= a and not b;
    layer0_outputs(12273) <= not (a and b);
    layer0_outputs(12274) <= a or b;
    layer0_outputs(12275) <= a and b;
    layer0_outputs(12276) <= b;
    layer0_outputs(12277) <= a and b;
    layer0_outputs(12278) <= not b;
    layer0_outputs(12279) <= a;
    layer0_outputs(12280) <= '0';
    layer0_outputs(12281) <= b;
    layer0_outputs(12282) <= not (a and b);
    layer0_outputs(12283) <= not a;
    layer0_outputs(12284) <= a xor b;
    layer0_outputs(12285) <= not (a or b);
    layer0_outputs(12286) <= b;
    layer0_outputs(12287) <= not b or a;
    layer0_outputs(12288) <= not a;
    layer0_outputs(12289) <= not (a and b);
    layer0_outputs(12290) <= b;
    layer0_outputs(12291) <= not b;
    layer0_outputs(12292) <= a or b;
    layer0_outputs(12293) <= not a or b;
    layer0_outputs(12294) <= not a or b;
    layer0_outputs(12295) <= not b or a;
    layer0_outputs(12296) <= b;
    layer0_outputs(12297) <= '1';
    layer0_outputs(12298) <= b;
    layer0_outputs(12299) <= not (a xor b);
    layer0_outputs(12300) <= b;
    layer0_outputs(12301) <= a and b;
    layer0_outputs(12302) <= a xor b;
    layer0_outputs(12303) <= not (a and b);
    layer0_outputs(12304) <= a;
    layer0_outputs(12305) <= a or b;
    layer0_outputs(12306) <= a and not b;
    layer0_outputs(12307) <= not (a xor b);
    layer0_outputs(12308) <= not (a xor b);
    layer0_outputs(12309) <= not b or a;
    layer0_outputs(12310) <= not b or a;
    layer0_outputs(12311) <= a xor b;
    layer0_outputs(12312) <= not (a or b);
    layer0_outputs(12313) <= not (a or b);
    layer0_outputs(12314) <= not (a and b);
    layer0_outputs(12315) <= b;
    layer0_outputs(12316) <= a;
    layer0_outputs(12317) <= not a;
    layer0_outputs(12318) <= not b;
    layer0_outputs(12319) <= '0';
    layer0_outputs(12320) <= not (a and b);
    layer0_outputs(12321) <= not (a xor b);
    layer0_outputs(12322) <= not b or a;
    layer0_outputs(12323) <= a and not b;
    layer0_outputs(12324) <= not (a and b);
    layer0_outputs(12325) <= a and not b;
    layer0_outputs(12326) <= a xor b;
    layer0_outputs(12327) <= '1';
    layer0_outputs(12328) <= a xor b;
    layer0_outputs(12329) <= not (a or b);
    layer0_outputs(12330) <= a xor b;
    layer0_outputs(12331) <= not a;
    layer0_outputs(12332) <= a and not b;
    layer0_outputs(12333) <= not b;
    layer0_outputs(12334) <= not (a xor b);
    layer0_outputs(12335) <= a xor b;
    layer0_outputs(12336) <= '1';
    layer0_outputs(12337) <= a;
    layer0_outputs(12338) <= '0';
    layer0_outputs(12339) <= not a;
    layer0_outputs(12340) <= not b or a;
    layer0_outputs(12341) <= not a;
    layer0_outputs(12342) <= not b;
    layer0_outputs(12343) <= a and not b;
    layer0_outputs(12344) <= a;
    layer0_outputs(12345) <= a xor b;
    layer0_outputs(12346) <= not b or a;
    layer0_outputs(12347) <= a and not b;
    layer0_outputs(12348) <= not a or b;
    layer0_outputs(12349) <= '1';
    layer0_outputs(12350) <= '0';
    layer0_outputs(12351) <= not a;
    layer0_outputs(12352) <= not a;
    layer0_outputs(12353) <= a;
    layer0_outputs(12354) <= a or b;
    layer0_outputs(12355) <= not (a and b);
    layer0_outputs(12356) <= not b or a;
    layer0_outputs(12357) <= not a or b;
    layer0_outputs(12358) <= not b or a;
    layer0_outputs(12359) <= '1';
    layer0_outputs(12360) <= not a;
    layer0_outputs(12361) <= not (a and b);
    layer0_outputs(12362) <= b and not a;
    layer0_outputs(12363) <= a xor b;
    layer0_outputs(12364) <= a or b;
    layer0_outputs(12365) <= not b or a;
    layer0_outputs(12366) <= a and b;
    layer0_outputs(12367) <= a or b;
    layer0_outputs(12368) <= '0';
    layer0_outputs(12369) <= a;
    layer0_outputs(12370) <= not a;
    layer0_outputs(12371) <= not (a or b);
    layer0_outputs(12372) <= not a;
    layer0_outputs(12373) <= b;
    layer0_outputs(12374) <= a or b;
    layer0_outputs(12375) <= not b or a;
    layer0_outputs(12376) <= not (a or b);
    layer0_outputs(12377) <= not a or b;
    layer0_outputs(12378) <= not (a and b);
    layer0_outputs(12379) <= b;
    layer0_outputs(12380) <= not a or b;
    layer0_outputs(12381) <= not b or a;
    layer0_outputs(12382) <= not (a or b);
    layer0_outputs(12383) <= not (a or b);
    layer0_outputs(12384) <= a or b;
    layer0_outputs(12385) <= b;
    layer0_outputs(12386) <= not b;
    layer0_outputs(12387) <= '0';
    layer0_outputs(12388) <= a;
    layer0_outputs(12389) <= a or b;
    layer0_outputs(12390) <= not (a or b);
    layer0_outputs(12391) <= not a;
    layer0_outputs(12392) <= not (a xor b);
    layer0_outputs(12393) <= not (a xor b);
    layer0_outputs(12394) <= not b;
    layer0_outputs(12395) <= b and not a;
    layer0_outputs(12396) <= not b or a;
    layer0_outputs(12397) <= a and not b;
    layer0_outputs(12398) <= a and b;
    layer0_outputs(12399) <= a;
    layer0_outputs(12400) <= a and not b;
    layer0_outputs(12401) <= a and b;
    layer0_outputs(12402) <= not a or b;
    layer0_outputs(12403) <= not a or b;
    layer0_outputs(12404) <= b and not a;
    layer0_outputs(12405) <= a xor b;
    layer0_outputs(12406) <= not b or a;
    layer0_outputs(12407) <= b;
    layer0_outputs(12408) <= '0';
    layer0_outputs(12409) <= not b or a;
    layer0_outputs(12410) <= not a;
    layer0_outputs(12411) <= a and b;
    layer0_outputs(12412) <= not b;
    layer0_outputs(12413) <= a;
    layer0_outputs(12414) <= not a;
    layer0_outputs(12415) <= not (a or b);
    layer0_outputs(12416) <= a;
    layer0_outputs(12417) <= not b or a;
    layer0_outputs(12418) <= b;
    layer0_outputs(12419) <= not b or a;
    layer0_outputs(12420) <= not a or b;
    layer0_outputs(12421) <= b;
    layer0_outputs(12422) <= b and not a;
    layer0_outputs(12423) <= b and not a;
    layer0_outputs(12424) <= not (a xor b);
    layer0_outputs(12425) <= not b;
    layer0_outputs(12426) <= not b;
    layer0_outputs(12427) <= b and not a;
    layer0_outputs(12428) <= not b;
    layer0_outputs(12429) <= not b or a;
    layer0_outputs(12430) <= a or b;
    layer0_outputs(12431) <= a and not b;
    layer0_outputs(12432) <= not a or b;
    layer0_outputs(12433) <= '0';
    layer0_outputs(12434) <= not (a xor b);
    layer0_outputs(12435) <= not a;
    layer0_outputs(12436) <= not (a and b);
    layer0_outputs(12437) <= a or b;
    layer0_outputs(12438) <= not (a xor b);
    layer0_outputs(12439) <= b;
    layer0_outputs(12440) <= a or b;
    layer0_outputs(12441) <= a and b;
    layer0_outputs(12442) <= '1';
    layer0_outputs(12443) <= not a or b;
    layer0_outputs(12444) <= a or b;
    layer0_outputs(12445) <= b and not a;
    layer0_outputs(12446) <= a or b;
    layer0_outputs(12447) <= not a;
    layer0_outputs(12448) <= a and not b;
    layer0_outputs(12449) <= a;
    layer0_outputs(12450) <= b and not a;
    layer0_outputs(12451) <= b and not a;
    layer0_outputs(12452) <= b;
    layer0_outputs(12453) <= a or b;
    layer0_outputs(12454) <= not (a or b);
    layer0_outputs(12455) <= not b;
    layer0_outputs(12456) <= not a;
    layer0_outputs(12457) <= a and b;
    layer0_outputs(12458) <= not b or a;
    layer0_outputs(12459) <= b;
    layer0_outputs(12460) <= '1';
    layer0_outputs(12461) <= a or b;
    layer0_outputs(12462) <= not (a or b);
    layer0_outputs(12463) <= not b;
    layer0_outputs(12464) <= not b;
    layer0_outputs(12465) <= a or b;
    layer0_outputs(12466) <= not b;
    layer0_outputs(12467) <= not (a or b);
    layer0_outputs(12468) <= '1';
    layer0_outputs(12469) <= a or b;
    layer0_outputs(12470) <= b and not a;
    layer0_outputs(12471) <= not b or a;
    layer0_outputs(12472) <= not a or b;
    layer0_outputs(12473) <= '0';
    layer0_outputs(12474) <= not (a and b);
    layer0_outputs(12475) <= not a;
    layer0_outputs(12476) <= not a;
    layer0_outputs(12477) <= a;
    layer0_outputs(12478) <= a or b;
    layer0_outputs(12479) <= a or b;
    layer0_outputs(12480) <= not b or a;
    layer0_outputs(12481) <= a;
    layer0_outputs(12482) <= '1';
    layer0_outputs(12483) <= not (a and b);
    layer0_outputs(12484) <= not a;
    layer0_outputs(12485) <= '1';
    layer0_outputs(12486) <= not a or b;
    layer0_outputs(12487) <= a or b;
    layer0_outputs(12488) <= a;
    layer0_outputs(12489) <= b and not a;
    layer0_outputs(12490) <= not a;
    layer0_outputs(12491) <= not (a or b);
    layer0_outputs(12492) <= a xor b;
    layer0_outputs(12493) <= not a or b;
    layer0_outputs(12494) <= '0';
    layer0_outputs(12495) <= not b or a;
    layer0_outputs(12496) <= not (a and b);
    layer0_outputs(12497) <= a or b;
    layer0_outputs(12498) <= not (a or b);
    layer0_outputs(12499) <= '0';
    layer0_outputs(12500) <= a and not b;
    layer0_outputs(12501) <= a or b;
    layer0_outputs(12502) <= not a or b;
    layer0_outputs(12503) <= a xor b;
    layer0_outputs(12504) <= a or b;
    layer0_outputs(12505) <= b and not a;
    layer0_outputs(12506) <= a or b;
    layer0_outputs(12507) <= '0';
    layer0_outputs(12508) <= a xor b;
    layer0_outputs(12509) <= not (a xor b);
    layer0_outputs(12510) <= a;
    layer0_outputs(12511) <= not (a or b);
    layer0_outputs(12512) <= a or b;
    layer0_outputs(12513) <= a or b;
    layer0_outputs(12514) <= b and not a;
    layer0_outputs(12515) <= a xor b;
    layer0_outputs(12516) <= b;
    layer0_outputs(12517) <= a xor b;
    layer0_outputs(12518) <= a or b;
    layer0_outputs(12519) <= not b;
    layer0_outputs(12520) <= a and not b;
    layer0_outputs(12521) <= not a;
    layer0_outputs(12522) <= '1';
    layer0_outputs(12523) <= b;
    layer0_outputs(12524) <= '0';
    layer0_outputs(12525) <= a or b;
    layer0_outputs(12526) <= not b;
    layer0_outputs(12527) <= not b or a;
    layer0_outputs(12528) <= '1';
    layer0_outputs(12529) <= '0';
    layer0_outputs(12530) <= not (a or b);
    layer0_outputs(12531) <= not b or a;
    layer0_outputs(12532) <= not (a xor b);
    layer0_outputs(12533) <= not (a and b);
    layer0_outputs(12534) <= not (a or b);
    layer0_outputs(12535) <= a or b;
    layer0_outputs(12536) <= '0';
    layer0_outputs(12537) <= not a;
    layer0_outputs(12538) <= '0';
    layer0_outputs(12539) <= not b or a;
    layer0_outputs(12540) <= '1';
    layer0_outputs(12541) <= a or b;
    layer0_outputs(12542) <= a and not b;
    layer0_outputs(12543) <= not a or b;
    layer0_outputs(12544) <= b;
    layer0_outputs(12545) <= a and b;
    layer0_outputs(12546) <= a;
    layer0_outputs(12547) <= not a;
    layer0_outputs(12548) <= b and not a;
    layer0_outputs(12549) <= not b;
    layer0_outputs(12550) <= b and not a;
    layer0_outputs(12551) <= '0';
    layer0_outputs(12552) <= a or b;
    layer0_outputs(12553) <= a;
    layer0_outputs(12554) <= a and not b;
    layer0_outputs(12555) <= a or b;
    layer0_outputs(12556) <= a xor b;
    layer0_outputs(12557) <= not b;
    layer0_outputs(12558) <= not a or b;
    layer0_outputs(12559) <= not (a and b);
    layer0_outputs(12560) <= not (a xor b);
    layer0_outputs(12561) <= b;
    layer0_outputs(12562) <= not (a and b);
    layer0_outputs(12563) <= '1';
    layer0_outputs(12564) <= not (a xor b);
    layer0_outputs(12565) <= a or b;
    layer0_outputs(12566) <= not a;
    layer0_outputs(12567) <= b;
    layer0_outputs(12568) <= a xor b;
    layer0_outputs(12569) <= not (a and b);
    layer0_outputs(12570) <= b;
    layer0_outputs(12571) <= not (a and b);
    layer0_outputs(12572) <= b and not a;
    layer0_outputs(12573) <= a xor b;
    layer0_outputs(12574) <= not (a and b);
    layer0_outputs(12575) <= not (a xor b);
    layer0_outputs(12576) <= not b;
    layer0_outputs(12577) <= a xor b;
    layer0_outputs(12578) <= not b or a;
    layer0_outputs(12579) <= not (a or b);
    layer0_outputs(12580) <= a;
    layer0_outputs(12581) <= not (a xor b);
    layer0_outputs(12582) <= not (a and b);
    layer0_outputs(12583) <= not (a or b);
    layer0_outputs(12584) <= not b or a;
    layer0_outputs(12585) <= not (a or b);
    layer0_outputs(12586) <= a and not b;
    layer0_outputs(12587) <= b and not a;
    layer0_outputs(12588) <= a;
    layer0_outputs(12589) <= a xor b;
    layer0_outputs(12590) <= '1';
    layer0_outputs(12591) <= '1';
    layer0_outputs(12592) <= a and b;
    layer0_outputs(12593) <= not a;
    layer0_outputs(12594) <= not a;
    layer0_outputs(12595) <= a;
    layer0_outputs(12596) <= a xor b;
    layer0_outputs(12597) <= a and not b;
    layer0_outputs(12598) <= a;
    layer0_outputs(12599) <= '1';
    layer0_outputs(12600) <= a xor b;
    layer0_outputs(12601) <= a or b;
    layer0_outputs(12602) <= b and not a;
    layer0_outputs(12603) <= not (a xor b);
    layer0_outputs(12604) <= a xor b;
    layer0_outputs(12605) <= b;
    layer0_outputs(12606) <= not b;
    layer0_outputs(12607) <= a;
    layer0_outputs(12608) <= b;
    layer0_outputs(12609) <= b and not a;
    layer0_outputs(12610) <= not (a xor b);
    layer0_outputs(12611) <= a;
    layer0_outputs(12612) <= a or b;
    layer0_outputs(12613) <= '1';
    layer0_outputs(12614) <= b and not a;
    layer0_outputs(12615) <= b;
    layer0_outputs(12616) <= '1';
    layer0_outputs(12617) <= '0';
    layer0_outputs(12618) <= b;
    layer0_outputs(12619) <= a and not b;
    layer0_outputs(12620) <= not a or b;
    layer0_outputs(12621) <= not (a or b);
    layer0_outputs(12622) <= not a;
    layer0_outputs(12623) <= not (a and b);
    layer0_outputs(12624) <= not a or b;
    layer0_outputs(12625) <= b;
    layer0_outputs(12626) <= '1';
    layer0_outputs(12627) <= a;
    layer0_outputs(12628) <= not a;
    layer0_outputs(12629) <= not a or b;
    layer0_outputs(12630) <= a or b;
    layer0_outputs(12631) <= not b or a;
    layer0_outputs(12632) <= not (a or b);
    layer0_outputs(12633) <= not a;
    layer0_outputs(12634) <= a and not b;
    layer0_outputs(12635) <= '1';
    layer0_outputs(12636) <= b;
    layer0_outputs(12637) <= not (a and b);
    layer0_outputs(12638) <= b;
    layer0_outputs(12639) <= not b;
    layer0_outputs(12640) <= '1';
    layer0_outputs(12641) <= not a;
    layer0_outputs(12642) <= not a;
    layer0_outputs(12643) <= a xor b;
    layer0_outputs(12644) <= a xor b;
    layer0_outputs(12645) <= b and not a;
    layer0_outputs(12646) <= b;
    layer0_outputs(12647) <= not (a and b);
    layer0_outputs(12648) <= not a;
    layer0_outputs(12649) <= '0';
    layer0_outputs(12650) <= a;
    layer0_outputs(12651) <= not a or b;
    layer0_outputs(12652) <= not a;
    layer0_outputs(12653) <= b;
    layer0_outputs(12654) <= not (a xor b);
    layer0_outputs(12655) <= not b or a;
    layer0_outputs(12656) <= b and not a;
    layer0_outputs(12657) <= not (a xor b);
    layer0_outputs(12658) <= a xor b;
    layer0_outputs(12659) <= a;
    layer0_outputs(12660) <= a and not b;
    layer0_outputs(12661) <= '0';
    layer0_outputs(12662) <= a and b;
    layer0_outputs(12663) <= a xor b;
    layer0_outputs(12664) <= not (a and b);
    layer0_outputs(12665) <= a xor b;
    layer0_outputs(12666) <= not (a or b);
    layer0_outputs(12667) <= not b;
    layer0_outputs(12668) <= not (a xor b);
    layer0_outputs(12669) <= a xor b;
    layer0_outputs(12670) <= '1';
    layer0_outputs(12671) <= a;
    layer0_outputs(12672) <= not a;
    layer0_outputs(12673) <= not b or a;
    layer0_outputs(12674) <= a;
    layer0_outputs(12675) <= not b;
    layer0_outputs(12676) <= a xor b;
    layer0_outputs(12677) <= a and not b;
    layer0_outputs(12678) <= a xor b;
    layer0_outputs(12679) <= a xor b;
    layer0_outputs(12680) <= a and not b;
    layer0_outputs(12681) <= not a;
    layer0_outputs(12682) <= a and not b;
    layer0_outputs(12683) <= not a or b;
    layer0_outputs(12684) <= b and not a;
    layer0_outputs(12685) <= not a;
    layer0_outputs(12686) <= not b or a;
    layer0_outputs(12687) <= a and b;
    layer0_outputs(12688) <= b;
    layer0_outputs(12689) <= not a or b;
    layer0_outputs(12690) <= not b;
    layer0_outputs(12691) <= a;
    layer0_outputs(12692) <= not b;
    layer0_outputs(12693) <= not b;
    layer0_outputs(12694) <= a or b;
    layer0_outputs(12695) <= not a;
    layer0_outputs(12696) <= not b or a;
    layer0_outputs(12697) <= not b;
    layer0_outputs(12698) <= a xor b;
    layer0_outputs(12699) <= not b or a;
    layer0_outputs(12700) <= b;
    layer0_outputs(12701) <= not b or a;
    layer0_outputs(12702) <= a or b;
    layer0_outputs(12703) <= a and not b;
    layer0_outputs(12704) <= not (a or b);
    layer0_outputs(12705) <= not b or a;
    layer0_outputs(12706) <= a and not b;
    layer0_outputs(12707) <= b;
    layer0_outputs(12708) <= a xor b;
    layer0_outputs(12709) <= not a;
    layer0_outputs(12710) <= '1';
    layer0_outputs(12711) <= not b;
    layer0_outputs(12712) <= a and not b;
    layer0_outputs(12713) <= not (a xor b);
    layer0_outputs(12714) <= b;
    layer0_outputs(12715) <= a and not b;
    layer0_outputs(12716) <= a and not b;
    layer0_outputs(12717) <= b;
    layer0_outputs(12718) <= a;
    layer0_outputs(12719) <= not a;
    layer0_outputs(12720) <= not (a or b);
    layer0_outputs(12721) <= not b;
    layer0_outputs(12722) <= '1';
    layer0_outputs(12723) <= '0';
    layer0_outputs(12724) <= not b;
    layer0_outputs(12725) <= not (a and b);
    layer0_outputs(12726) <= a;
    layer0_outputs(12727) <= not b or a;
    layer0_outputs(12728) <= not b or a;
    layer0_outputs(12729) <= a or b;
    layer0_outputs(12730) <= a or b;
    layer0_outputs(12731) <= not b;
    layer0_outputs(12732) <= a or b;
    layer0_outputs(12733) <= b;
    layer0_outputs(12734) <= b and not a;
    layer0_outputs(12735) <= not (a xor b);
    layer0_outputs(12736) <= not (a and b);
    layer0_outputs(12737) <= b and not a;
    layer0_outputs(12738) <= not b;
    layer0_outputs(12739) <= not b;
    layer0_outputs(12740) <= not b or a;
    layer0_outputs(12741) <= a xor b;
    layer0_outputs(12742) <= a or b;
    layer0_outputs(12743) <= '0';
    layer0_outputs(12744) <= b and not a;
    layer0_outputs(12745) <= not a or b;
    layer0_outputs(12746) <= not (a xor b);
    layer0_outputs(12747) <= a and b;
    layer0_outputs(12748) <= not (a or b);
    layer0_outputs(12749) <= b and not a;
    layer0_outputs(12750) <= not a or b;
    layer0_outputs(12751) <= not a;
    layer0_outputs(12752) <= not (a and b);
    layer0_outputs(12753) <= a;
    layer0_outputs(12754) <= not b or a;
    layer0_outputs(12755) <= a xor b;
    layer0_outputs(12756) <= a and not b;
    layer0_outputs(12757) <= a or b;
    layer0_outputs(12758) <= not (a and b);
    layer0_outputs(12759) <= not b or a;
    layer0_outputs(12760) <= b;
    layer0_outputs(12761) <= not (a or b);
    layer0_outputs(12762) <= a xor b;
    layer0_outputs(12763) <= not a or b;
    layer0_outputs(12764) <= a and b;
    layer0_outputs(12765) <= a xor b;
    layer0_outputs(12766) <= not a;
    layer0_outputs(12767) <= '0';
    layer0_outputs(12768) <= not a or b;
    layer0_outputs(12769) <= b;
    layer0_outputs(12770) <= not a or b;
    layer0_outputs(12771) <= not b or a;
    layer0_outputs(12772) <= a;
    layer0_outputs(12773) <= not (a xor b);
    layer0_outputs(12774) <= not (a xor b);
    layer0_outputs(12775) <= b and not a;
    layer0_outputs(12776) <= a;
    layer0_outputs(12777) <= a xor b;
    layer0_outputs(12778) <= not b or a;
    layer0_outputs(12779) <= a xor b;
    layer0_outputs(12780) <= not (a and b);
    layer0_outputs(12781) <= a and b;
    layer0_outputs(12782) <= a xor b;
    layer0_outputs(12783) <= not a;
    layer0_outputs(12784) <= a and not b;
    layer0_outputs(12785) <= not (a or b);
    layer0_outputs(12786) <= a;
    layer0_outputs(12787) <= b;
    layer0_outputs(12788) <= not (a or b);
    layer0_outputs(12789) <= not b or a;
    layer0_outputs(12790) <= not b;
    layer0_outputs(12791) <= a xor b;
    layer0_outputs(12792) <= b;
    layer0_outputs(12793) <= not (a and b);
    layer0_outputs(12794) <= not (a xor b);
    layer0_outputs(12795) <= not (a xor b);
    layer0_outputs(12796) <= not a or b;
    layer0_outputs(12797) <= not (a xor b);
    layer0_outputs(12798) <= not a or b;
    layer0_outputs(12799) <= '1';
    layer1_outputs(0) <= a;
    layer1_outputs(1) <= b and not a;
    layer1_outputs(2) <= b;
    layer1_outputs(3) <= b and not a;
    layer1_outputs(4) <= '1';
    layer1_outputs(5) <= a xor b;
    layer1_outputs(6) <= '1';
    layer1_outputs(7) <= not (a xor b);
    layer1_outputs(8) <= not a;
    layer1_outputs(9) <= a or b;
    layer1_outputs(10) <= not (a xor b);
    layer1_outputs(11) <= not a;
    layer1_outputs(12) <= not b;
    layer1_outputs(13) <= not (a and b);
    layer1_outputs(14) <= not (a xor b);
    layer1_outputs(15) <= not a;
    layer1_outputs(16) <= not b;
    layer1_outputs(17) <= b;
    layer1_outputs(18) <= b and not a;
    layer1_outputs(19) <= not b;
    layer1_outputs(20) <= not a or b;
    layer1_outputs(21) <= b;
    layer1_outputs(22) <= b;
    layer1_outputs(23) <= b and not a;
    layer1_outputs(24) <= b and not a;
    layer1_outputs(25) <= not b or a;
    layer1_outputs(26) <= '0';
    layer1_outputs(27) <= not b;
    layer1_outputs(28) <= a and not b;
    layer1_outputs(29) <= not a or b;
    layer1_outputs(30) <= not a or b;
    layer1_outputs(31) <= a xor b;
    layer1_outputs(32) <= a;
    layer1_outputs(33) <= a or b;
    layer1_outputs(34) <= not (a and b);
    layer1_outputs(35) <= not a;
    layer1_outputs(36) <= not (a and b);
    layer1_outputs(37) <= not a;
    layer1_outputs(38) <= '0';
    layer1_outputs(39) <= b;
    layer1_outputs(40) <= a xor b;
    layer1_outputs(41) <= '1';
    layer1_outputs(42) <= not (a or b);
    layer1_outputs(43) <= not a or b;
    layer1_outputs(44) <= '1';
    layer1_outputs(45) <= b and not a;
    layer1_outputs(46) <= b;
    layer1_outputs(47) <= '0';
    layer1_outputs(48) <= b and not a;
    layer1_outputs(49) <= a;
    layer1_outputs(50) <= not a;
    layer1_outputs(51) <= a;
    layer1_outputs(52) <= a and not b;
    layer1_outputs(53) <= b;
    layer1_outputs(54) <= not a or b;
    layer1_outputs(55) <= a and not b;
    layer1_outputs(56) <= not a;
    layer1_outputs(57) <= a and b;
    layer1_outputs(58) <= not (a and b);
    layer1_outputs(59) <= not (a or b);
    layer1_outputs(60) <= a;
    layer1_outputs(61) <= a;
    layer1_outputs(62) <= a;
    layer1_outputs(63) <= a and b;
    layer1_outputs(64) <= not b;
    layer1_outputs(65) <= b and not a;
    layer1_outputs(66) <= a;
    layer1_outputs(67) <= '1';
    layer1_outputs(68) <= not a;
    layer1_outputs(69) <= not b;
    layer1_outputs(70) <= not b;
    layer1_outputs(71) <= a and not b;
    layer1_outputs(72) <= not a;
    layer1_outputs(73) <= a and not b;
    layer1_outputs(74) <= not b or a;
    layer1_outputs(75) <= not (a or b);
    layer1_outputs(76) <= not a;
    layer1_outputs(77) <= not a or b;
    layer1_outputs(78) <= b and not a;
    layer1_outputs(79) <= not b;
    layer1_outputs(80) <= a or b;
    layer1_outputs(81) <= '0';
    layer1_outputs(82) <= not (a or b);
    layer1_outputs(83) <= '0';
    layer1_outputs(84) <= a and b;
    layer1_outputs(85) <= b;
    layer1_outputs(86) <= a;
    layer1_outputs(87) <= b;
    layer1_outputs(88) <= '0';
    layer1_outputs(89) <= not (a or b);
    layer1_outputs(90) <= not b;
    layer1_outputs(91) <= a;
    layer1_outputs(92) <= '1';
    layer1_outputs(93) <= a or b;
    layer1_outputs(94) <= a and not b;
    layer1_outputs(95) <= a;
    layer1_outputs(96) <= not b;
    layer1_outputs(97) <= not (a and b);
    layer1_outputs(98) <= a xor b;
    layer1_outputs(99) <= not b or a;
    layer1_outputs(100) <= not b or a;
    layer1_outputs(101) <= a and not b;
    layer1_outputs(102) <= not b;
    layer1_outputs(103) <= not a;
    layer1_outputs(104) <= not a or b;
    layer1_outputs(105) <= a and not b;
    layer1_outputs(106) <= '0';
    layer1_outputs(107) <= not b;
    layer1_outputs(108) <= a xor b;
    layer1_outputs(109) <= not a;
    layer1_outputs(110) <= a or b;
    layer1_outputs(111) <= a or b;
    layer1_outputs(112) <= a and not b;
    layer1_outputs(113) <= a and b;
    layer1_outputs(114) <= b;
    layer1_outputs(115) <= '1';
    layer1_outputs(116) <= '1';
    layer1_outputs(117) <= not (a xor b);
    layer1_outputs(118) <= a;
    layer1_outputs(119) <= not (a and b);
    layer1_outputs(120) <= not (a and b);
    layer1_outputs(121) <= a;
    layer1_outputs(122) <= not b;
    layer1_outputs(123) <= not a or b;
    layer1_outputs(124) <= not a or b;
    layer1_outputs(125) <= b and not a;
    layer1_outputs(126) <= a xor b;
    layer1_outputs(127) <= b;
    layer1_outputs(128) <= a;
    layer1_outputs(129) <= a;
    layer1_outputs(130) <= not (a or b);
    layer1_outputs(131) <= not (a and b);
    layer1_outputs(132) <= not (a and b);
    layer1_outputs(133) <= '0';
    layer1_outputs(134) <= not (a and b);
    layer1_outputs(135) <= not (a or b);
    layer1_outputs(136) <= not (a xor b);
    layer1_outputs(137) <= a xor b;
    layer1_outputs(138) <= b and not a;
    layer1_outputs(139) <= b;
    layer1_outputs(140) <= not (a and b);
    layer1_outputs(141) <= a or b;
    layer1_outputs(142) <= not (a and b);
    layer1_outputs(143) <= a or b;
    layer1_outputs(144) <= b and not a;
    layer1_outputs(145) <= a or b;
    layer1_outputs(146) <= a and b;
    layer1_outputs(147) <= not a or b;
    layer1_outputs(148) <= a or b;
    layer1_outputs(149) <= a and not b;
    layer1_outputs(150) <= not a;
    layer1_outputs(151) <= a and not b;
    layer1_outputs(152) <= '0';
    layer1_outputs(153) <= '0';
    layer1_outputs(154) <= a and not b;
    layer1_outputs(155) <= b and not a;
    layer1_outputs(156) <= '1';
    layer1_outputs(157) <= not a;
    layer1_outputs(158) <= '1';
    layer1_outputs(159) <= not (a xor b);
    layer1_outputs(160) <= b;
    layer1_outputs(161) <= not (a and b);
    layer1_outputs(162) <= b;
    layer1_outputs(163) <= not (a and b);
    layer1_outputs(164) <= b and not a;
    layer1_outputs(165) <= a or b;
    layer1_outputs(166) <= not a;
    layer1_outputs(167) <= b and not a;
    layer1_outputs(168) <= b;
    layer1_outputs(169) <= a;
    layer1_outputs(170) <= not a;
    layer1_outputs(171) <= a;
    layer1_outputs(172) <= a or b;
    layer1_outputs(173) <= b and not a;
    layer1_outputs(174) <= not (a and b);
    layer1_outputs(175) <= a;
    layer1_outputs(176) <= '1';
    layer1_outputs(177) <= a and b;
    layer1_outputs(178) <= a xor b;
    layer1_outputs(179) <= not a or b;
    layer1_outputs(180) <= not b or a;
    layer1_outputs(181) <= '0';
    layer1_outputs(182) <= not b;
    layer1_outputs(183) <= not a or b;
    layer1_outputs(184) <= '1';
    layer1_outputs(185) <= not b;
    layer1_outputs(186) <= not b or a;
    layer1_outputs(187) <= '1';
    layer1_outputs(188) <= b;
    layer1_outputs(189) <= a and b;
    layer1_outputs(190) <= not a or b;
    layer1_outputs(191) <= not (a and b);
    layer1_outputs(192) <= a;
    layer1_outputs(193) <= not b or a;
    layer1_outputs(194) <= not b;
    layer1_outputs(195) <= a and b;
    layer1_outputs(196) <= a or b;
    layer1_outputs(197) <= a;
    layer1_outputs(198) <= not (a or b);
    layer1_outputs(199) <= a and b;
    layer1_outputs(200) <= not (a or b);
    layer1_outputs(201) <= not b or a;
    layer1_outputs(202) <= not (a or b);
    layer1_outputs(203) <= b;
    layer1_outputs(204) <= not (a or b);
    layer1_outputs(205) <= not (a or b);
    layer1_outputs(206) <= not (a and b);
    layer1_outputs(207) <= b;
    layer1_outputs(208) <= a or b;
    layer1_outputs(209) <= a and b;
    layer1_outputs(210) <= not a;
    layer1_outputs(211) <= not a or b;
    layer1_outputs(212) <= b;
    layer1_outputs(213) <= not b or a;
    layer1_outputs(214) <= not a;
    layer1_outputs(215) <= b and not a;
    layer1_outputs(216) <= not a;
    layer1_outputs(217) <= a xor b;
    layer1_outputs(218) <= a;
    layer1_outputs(219) <= not b or a;
    layer1_outputs(220) <= b;
    layer1_outputs(221) <= a and b;
    layer1_outputs(222) <= a and not b;
    layer1_outputs(223) <= '0';
    layer1_outputs(224) <= not (a and b);
    layer1_outputs(225) <= a and b;
    layer1_outputs(226) <= not b or a;
    layer1_outputs(227) <= not (a xor b);
    layer1_outputs(228) <= '1';
    layer1_outputs(229) <= not a;
    layer1_outputs(230) <= '0';
    layer1_outputs(231) <= '1';
    layer1_outputs(232) <= not a;
    layer1_outputs(233) <= not (a or b);
    layer1_outputs(234) <= not (a and b);
    layer1_outputs(235) <= '0';
    layer1_outputs(236) <= not (a xor b);
    layer1_outputs(237) <= b;
    layer1_outputs(238) <= '0';
    layer1_outputs(239) <= '1';
    layer1_outputs(240) <= b and not a;
    layer1_outputs(241) <= '0';
    layer1_outputs(242) <= '0';
    layer1_outputs(243) <= a or b;
    layer1_outputs(244) <= b;
    layer1_outputs(245) <= not (a xor b);
    layer1_outputs(246) <= b and not a;
    layer1_outputs(247) <= not b or a;
    layer1_outputs(248) <= b and not a;
    layer1_outputs(249) <= not b or a;
    layer1_outputs(250) <= not a;
    layer1_outputs(251) <= not b or a;
    layer1_outputs(252) <= not b;
    layer1_outputs(253) <= not a or b;
    layer1_outputs(254) <= a xor b;
    layer1_outputs(255) <= not (a xor b);
    layer1_outputs(256) <= not (a and b);
    layer1_outputs(257) <= a and b;
    layer1_outputs(258) <= not a or b;
    layer1_outputs(259) <= '0';
    layer1_outputs(260) <= b;
    layer1_outputs(261) <= a and b;
    layer1_outputs(262) <= not (a or b);
    layer1_outputs(263) <= a and not b;
    layer1_outputs(264) <= not b or a;
    layer1_outputs(265) <= b;
    layer1_outputs(266) <= not (a or b);
    layer1_outputs(267) <= not a or b;
    layer1_outputs(268) <= a and b;
    layer1_outputs(269) <= b and not a;
    layer1_outputs(270) <= a xor b;
    layer1_outputs(271) <= not a;
    layer1_outputs(272) <= a;
    layer1_outputs(273) <= a and not b;
    layer1_outputs(274) <= not (a xor b);
    layer1_outputs(275) <= a and not b;
    layer1_outputs(276) <= not b or a;
    layer1_outputs(277) <= not b;
    layer1_outputs(278) <= b;
    layer1_outputs(279) <= b and not a;
    layer1_outputs(280) <= b;
    layer1_outputs(281) <= b;
    layer1_outputs(282) <= not b;
    layer1_outputs(283) <= not b or a;
    layer1_outputs(284) <= '1';
    layer1_outputs(285) <= not a;
    layer1_outputs(286) <= b;
    layer1_outputs(287) <= '0';
    layer1_outputs(288) <= '1';
    layer1_outputs(289) <= '1';
    layer1_outputs(290) <= not a or b;
    layer1_outputs(291) <= a;
    layer1_outputs(292) <= not (a xor b);
    layer1_outputs(293) <= not a;
    layer1_outputs(294) <= not b;
    layer1_outputs(295) <= a;
    layer1_outputs(296) <= not a or b;
    layer1_outputs(297) <= a or b;
    layer1_outputs(298) <= not (a xor b);
    layer1_outputs(299) <= b;
    layer1_outputs(300) <= not b;
    layer1_outputs(301) <= not (a xor b);
    layer1_outputs(302) <= b;
    layer1_outputs(303) <= a;
    layer1_outputs(304) <= not a or b;
    layer1_outputs(305) <= b;
    layer1_outputs(306) <= b and not a;
    layer1_outputs(307) <= b and not a;
    layer1_outputs(308) <= not b;
    layer1_outputs(309) <= not (a or b);
    layer1_outputs(310) <= '1';
    layer1_outputs(311) <= not (a and b);
    layer1_outputs(312) <= not (a xor b);
    layer1_outputs(313) <= '1';
    layer1_outputs(314) <= b and not a;
    layer1_outputs(315) <= not b or a;
    layer1_outputs(316) <= '0';
    layer1_outputs(317) <= b;
    layer1_outputs(318) <= not b;
    layer1_outputs(319) <= a or b;
    layer1_outputs(320) <= not b or a;
    layer1_outputs(321) <= b;
    layer1_outputs(322) <= a;
    layer1_outputs(323) <= b;
    layer1_outputs(324) <= '1';
    layer1_outputs(325) <= a;
    layer1_outputs(326) <= not b or a;
    layer1_outputs(327) <= b and not a;
    layer1_outputs(328) <= not a or b;
    layer1_outputs(329) <= not b;
    layer1_outputs(330) <= not a;
    layer1_outputs(331) <= not b or a;
    layer1_outputs(332) <= not (a or b);
    layer1_outputs(333) <= b;
    layer1_outputs(334) <= '1';
    layer1_outputs(335) <= not a;
    layer1_outputs(336) <= not (a or b);
    layer1_outputs(337) <= b and not a;
    layer1_outputs(338) <= not (a and b);
    layer1_outputs(339) <= not a;
    layer1_outputs(340) <= not a or b;
    layer1_outputs(341) <= not (a or b);
    layer1_outputs(342) <= '1';
    layer1_outputs(343) <= a or b;
    layer1_outputs(344) <= not b;
    layer1_outputs(345) <= not a;
    layer1_outputs(346) <= a xor b;
    layer1_outputs(347) <= '1';
    layer1_outputs(348) <= a and b;
    layer1_outputs(349) <= not a;
    layer1_outputs(350) <= not (a xor b);
    layer1_outputs(351) <= b;
    layer1_outputs(352) <= not (a and b);
    layer1_outputs(353) <= '1';
    layer1_outputs(354) <= a and b;
    layer1_outputs(355) <= not (a and b);
    layer1_outputs(356) <= a;
    layer1_outputs(357) <= '1';
    layer1_outputs(358) <= a and b;
    layer1_outputs(359) <= not a or b;
    layer1_outputs(360) <= not a or b;
    layer1_outputs(361) <= a and b;
    layer1_outputs(362) <= a;
    layer1_outputs(363) <= '0';
    layer1_outputs(364) <= not a or b;
    layer1_outputs(365) <= b and not a;
    layer1_outputs(366) <= '0';
    layer1_outputs(367) <= a xor b;
    layer1_outputs(368) <= a and not b;
    layer1_outputs(369) <= not (a or b);
    layer1_outputs(370) <= a and not b;
    layer1_outputs(371) <= not a;
    layer1_outputs(372) <= a and not b;
    layer1_outputs(373) <= not a or b;
    layer1_outputs(374) <= a xor b;
    layer1_outputs(375) <= b and not a;
    layer1_outputs(376) <= not (a and b);
    layer1_outputs(377) <= not b;
    layer1_outputs(378) <= a or b;
    layer1_outputs(379) <= a or b;
    layer1_outputs(380) <= not a;
    layer1_outputs(381) <= b and not a;
    layer1_outputs(382) <= a;
    layer1_outputs(383) <= not (a xor b);
    layer1_outputs(384) <= '0';
    layer1_outputs(385) <= not b;
    layer1_outputs(386) <= '1';
    layer1_outputs(387) <= '1';
    layer1_outputs(388) <= '0';
    layer1_outputs(389) <= not (a and b);
    layer1_outputs(390) <= not b;
    layer1_outputs(391) <= a and b;
    layer1_outputs(392) <= not (a and b);
    layer1_outputs(393) <= not b;
    layer1_outputs(394) <= a xor b;
    layer1_outputs(395) <= b;
    layer1_outputs(396) <= a;
    layer1_outputs(397) <= b and not a;
    layer1_outputs(398) <= a and b;
    layer1_outputs(399) <= not a or b;
    layer1_outputs(400) <= not a;
    layer1_outputs(401) <= not a;
    layer1_outputs(402) <= a and b;
    layer1_outputs(403) <= a;
    layer1_outputs(404) <= '1';
    layer1_outputs(405) <= a;
    layer1_outputs(406) <= b and not a;
    layer1_outputs(407) <= not b;
    layer1_outputs(408) <= a and b;
    layer1_outputs(409) <= not b;
    layer1_outputs(410) <= a xor b;
    layer1_outputs(411) <= a or b;
    layer1_outputs(412) <= not (a or b);
    layer1_outputs(413) <= not b or a;
    layer1_outputs(414) <= not (a or b);
    layer1_outputs(415) <= '1';
    layer1_outputs(416) <= '1';
    layer1_outputs(417) <= not b or a;
    layer1_outputs(418) <= a or b;
    layer1_outputs(419) <= a or b;
    layer1_outputs(420) <= a or b;
    layer1_outputs(421) <= '0';
    layer1_outputs(422) <= b and not a;
    layer1_outputs(423) <= a xor b;
    layer1_outputs(424) <= '0';
    layer1_outputs(425) <= '0';
    layer1_outputs(426) <= a xor b;
    layer1_outputs(427) <= b and not a;
    layer1_outputs(428) <= not (a or b);
    layer1_outputs(429) <= b and not a;
    layer1_outputs(430) <= not (a or b);
    layer1_outputs(431) <= a and not b;
    layer1_outputs(432) <= not (a or b);
    layer1_outputs(433) <= not b;
    layer1_outputs(434) <= a xor b;
    layer1_outputs(435) <= a;
    layer1_outputs(436) <= a and b;
    layer1_outputs(437) <= '0';
    layer1_outputs(438) <= not b;
    layer1_outputs(439) <= a or b;
    layer1_outputs(440) <= not b or a;
    layer1_outputs(441) <= b;
    layer1_outputs(442) <= '0';
    layer1_outputs(443) <= '0';
    layer1_outputs(444) <= '1';
    layer1_outputs(445) <= not b;
    layer1_outputs(446) <= not a or b;
    layer1_outputs(447) <= a or b;
    layer1_outputs(448) <= not a;
    layer1_outputs(449) <= b;
    layer1_outputs(450) <= '0';
    layer1_outputs(451) <= '0';
    layer1_outputs(452) <= '0';
    layer1_outputs(453) <= a and b;
    layer1_outputs(454) <= a;
    layer1_outputs(455) <= not (a and b);
    layer1_outputs(456) <= not a or b;
    layer1_outputs(457) <= not a;
    layer1_outputs(458) <= not b or a;
    layer1_outputs(459) <= not a;
    layer1_outputs(460) <= not (a and b);
    layer1_outputs(461) <= a and b;
    layer1_outputs(462) <= a;
    layer1_outputs(463) <= not (a or b);
    layer1_outputs(464) <= not a;
    layer1_outputs(465) <= a;
    layer1_outputs(466) <= not b;
    layer1_outputs(467) <= '0';
    layer1_outputs(468) <= a or b;
    layer1_outputs(469) <= a xor b;
    layer1_outputs(470) <= not (a xor b);
    layer1_outputs(471) <= a;
    layer1_outputs(472) <= not a;
    layer1_outputs(473) <= not (a and b);
    layer1_outputs(474) <= not a or b;
    layer1_outputs(475) <= not b or a;
    layer1_outputs(476) <= not a;
    layer1_outputs(477) <= '0';
    layer1_outputs(478) <= not (a and b);
    layer1_outputs(479) <= '1';
    layer1_outputs(480) <= '0';
    layer1_outputs(481) <= '0';
    layer1_outputs(482) <= a or b;
    layer1_outputs(483) <= not a;
    layer1_outputs(484) <= not a or b;
    layer1_outputs(485) <= not a or b;
    layer1_outputs(486) <= a and b;
    layer1_outputs(487) <= b;
    layer1_outputs(488) <= not (a and b);
    layer1_outputs(489) <= not (a and b);
    layer1_outputs(490) <= b and not a;
    layer1_outputs(491) <= b;
    layer1_outputs(492) <= not a or b;
    layer1_outputs(493) <= a and not b;
    layer1_outputs(494) <= not a;
    layer1_outputs(495) <= a and b;
    layer1_outputs(496) <= a and b;
    layer1_outputs(497) <= a;
    layer1_outputs(498) <= not b;
    layer1_outputs(499) <= not b or a;
    layer1_outputs(500) <= a and not b;
    layer1_outputs(501) <= not (a xor b);
    layer1_outputs(502) <= a xor b;
    layer1_outputs(503) <= not b;
    layer1_outputs(504) <= a and not b;
    layer1_outputs(505) <= not (a and b);
    layer1_outputs(506) <= a;
    layer1_outputs(507) <= '1';
    layer1_outputs(508) <= a;
    layer1_outputs(509) <= '0';
    layer1_outputs(510) <= a and not b;
    layer1_outputs(511) <= not a;
    layer1_outputs(512) <= not b or a;
    layer1_outputs(513) <= not (a and b);
    layer1_outputs(514) <= '1';
    layer1_outputs(515) <= not (a or b);
    layer1_outputs(516) <= b and not a;
    layer1_outputs(517) <= not a;
    layer1_outputs(518) <= b;
    layer1_outputs(519) <= b;
    layer1_outputs(520) <= a and b;
    layer1_outputs(521) <= a or b;
    layer1_outputs(522) <= '1';
    layer1_outputs(523) <= a and b;
    layer1_outputs(524) <= not (a or b);
    layer1_outputs(525) <= not a or b;
    layer1_outputs(526) <= '1';
    layer1_outputs(527) <= not (a or b);
    layer1_outputs(528) <= a and not b;
    layer1_outputs(529) <= '1';
    layer1_outputs(530) <= b;
    layer1_outputs(531) <= a or b;
    layer1_outputs(532) <= not (a and b);
    layer1_outputs(533) <= a;
    layer1_outputs(534) <= '1';
    layer1_outputs(535) <= b;
    layer1_outputs(536) <= not a;
    layer1_outputs(537) <= not b or a;
    layer1_outputs(538) <= not b or a;
    layer1_outputs(539) <= a and not b;
    layer1_outputs(540) <= not a;
    layer1_outputs(541) <= not a or b;
    layer1_outputs(542) <= not (a and b);
    layer1_outputs(543) <= not b or a;
    layer1_outputs(544) <= a or b;
    layer1_outputs(545) <= b and not a;
    layer1_outputs(546) <= not (a or b);
    layer1_outputs(547) <= not a or b;
    layer1_outputs(548) <= not b;
    layer1_outputs(549) <= a and b;
    layer1_outputs(550) <= not a;
    layer1_outputs(551) <= b and not a;
    layer1_outputs(552) <= not b or a;
    layer1_outputs(553) <= a and not b;
    layer1_outputs(554) <= b and not a;
    layer1_outputs(555) <= '0';
    layer1_outputs(556) <= not a;
    layer1_outputs(557) <= not b;
    layer1_outputs(558) <= not a;
    layer1_outputs(559) <= b and not a;
    layer1_outputs(560) <= not a;
    layer1_outputs(561) <= not b;
    layer1_outputs(562) <= not b or a;
    layer1_outputs(563) <= b;
    layer1_outputs(564) <= a and not b;
    layer1_outputs(565) <= not b or a;
    layer1_outputs(566) <= a or b;
    layer1_outputs(567) <= not b or a;
    layer1_outputs(568) <= not (a or b);
    layer1_outputs(569) <= b;
    layer1_outputs(570) <= a or b;
    layer1_outputs(571) <= a or b;
    layer1_outputs(572) <= '0';
    layer1_outputs(573) <= not b or a;
    layer1_outputs(574) <= not (a and b);
    layer1_outputs(575) <= a xor b;
    layer1_outputs(576) <= a;
    layer1_outputs(577) <= a and not b;
    layer1_outputs(578) <= not b or a;
    layer1_outputs(579) <= not b;
    layer1_outputs(580) <= a or b;
    layer1_outputs(581) <= b;
    layer1_outputs(582) <= not (a and b);
    layer1_outputs(583) <= '0';
    layer1_outputs(584) <= not b;
    layer1_outputs(585) <= b and not a;
    layer1_outputs(586) <= not (a and b);
    layer1_outputs(587) <= not a;
    layer1_outputs(588) <= not (a and b);
    layer1_outputs(589) <= a and not b;
    layer1_outputs(590) <= not b or a;
    layer1_outputs(591) <= not (a and b);
    layer1_outputs(592) <= a and b;
    layer1_outputs(593) <= not b;
    layer1_outputs(594) <= not a;
    layer1_outputs(595) <= '0';
    layer1_outputs(596) <= b;
    layer1_outputs(597) <= not a or b;
    layer1_outputs(598) <= '1';
    layer1_outputs(599) <= '1';
    layer1_outputs(600) <= not b;
    layer1_outputs(601) <= not (a xor b);
    layer1_outputs(602) <= a and not b;
    layer1_outputs(603) <= a xor b;
    layer1_outputs(604) <= a xor b;
    layer1_outputs(605) <= b;
    layer1_outputs(606) <= b;
    layer1_outputs(607) <= b;
    layer1_outputs(608) <= '1';
    layer1_outputs(609) <= not (a or b);
    layer1_outputs(610) <= b;
    layer1_outputs(611) <= not (a or b);
    layer1_outputs(612) <= a and b;
    layer1_outputs(613) <= not b;
    layer1_outputs(614) <= a and b;
    layer1_outputs(615) <= a;
    layer1_outputs(616) <= not (a and b);
    layer1_outputs(617) <= a xor b;
    layer1_outputs(618) <= a or b;
    layer1_outputs(619) <= a or b;
    layer1_outputs(620) <= not a;
    layer1_outputs(621) <= b and not a;
    layer1_outputs(622) <= not b;
    layer1_outputs(623) <= '1';
    layer1_outputs(624) <= not a;
    layer1_outputs(625) <= '1';
    layer1_outputs(626) <= not (a or b);
    layer1_outputs(627) <= not a or b;
    layer1_outputs(628) <= not a;
    layer1_outputs(629) <= a and b;
    layer1_outputs(630) <= not b;
    layer1_outputs(631) <= b and not a;
    layer1_outputs(632) <= not (a xor b);
    layer1_outputs(633) <= a and not b;
    layer1_outputs(634) <= a;
    layer1_outputs(635) <= not a or b;
    layer1_outputs(636) <= a or b;
    layer1_outputs(637) <= not b;
    layer1_outputs(638) <= b;
    layer1_outputs(639) <= b;
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= not (a and b);
    layer1_outputs(642) <= not b or a;
    layer1_outputs(643) <= a or b;
    layer1_outputs(644) <= not a;
    layer1_outputs(645) <= not (a or b);
    layer1_outputs(646) <= a and b;
    layer1_outputs(647) <= b;
    layer1_outputs(648) <= b;
    layer1_outputs(649) <= a and not b;
    layer1_outputs(650) <= a and b;
    layer1_outputs(651) <= not b or a;
    layer1_outputs(652) <= b;
    layer1_outputs(653) <= '0';
    layer1_outputs(654) <= '0';
    layer1_outputs(655) <= b;
    layer1_outputs(656) <= b;
    layer1_outputs(657) <= a and b;
    layer1_outputs(658) <= not a or b;
    layer1_outputs(659) <= b;
    layer1_outputs(660) <= not (a and b);
    layer1_outputs(661) <= a and b;
    layer1_outputs(662) <= not (a and b);
    layer1_outputs(663) <= not b or a;
    layer1_outputs(664) <= '0';
    layer1_outputs(665) <= b;
    layer1_outputs(666) <= a and b;
    layer1_outputs(667) <= b and not a;
    layer1_outputs(668) <= '1';
    layer1_outputs(669) <= not b or a;
    layer1_outputs(670) <= not (a and b);
    layer1_outputs(671) <= b;
    layer1_outputs(672) <= not (a or b);
    layer1_outputs(673) <= a;
    layer1_outputs(674) <= a and b;
    layer1_outputs(675) <= b and not a;
    layer1_outputs(676) <= '0';
    layer1_outputs(677) <= a;
    layer1_outputs(678) <= not a or b;
    layer1_outputs(679) <= not a or b;
    layer1_outputs(680) <= not a;
    layer1_outputs(681) <= not (a or b);
    layer1_outputs(682) <= not a or b;
    layer1_outputs(683) <= not b;
    layer1_outputs(684) <= a;
    layer1_outputs(685) <= a and b;
    layer1_outputs(686) <= '0';
    layer1_outputs(687) <= a and not b;
    layer1_outputs(688) <= not b or a;
    layer1_outputs(689) <= '1';
    layer1_outputs(690) <= a and b;
    layer1_outputs(691) <= not b;
    layer1_outputs(692) <= b;
    layer1_outputs(693) <= not a;
    layer1_outputs(694) <= '1';
    layer1_outputs(695) <= not (a or b);
    layer1_outputs(696) <= not (a or b);
    layer1_outputs(697) <= a and not b;
    layer1_outputs(698) <= b and not a;
    layer1_outputs(699) <= b and not a;
    layer1_outputs(700) <= not (a xor b);
    layer1_outputs(701) <= a and not b;
    layer1_outputs(702) <= '1';
    layer1_outputs(703) <= a and not b;
    layer1_outputs(704) <= b;
    layer1_outputs(705) <= not a or b;
    layer1_outputs(706) <= not a or b;
    layer1_outputs(707) <= not b;
    layer1_outputs(708) <= not (a or b);
    layer1_outputs(709) <= a and b;
    layer1_outputs(710) <= not (a and b);
    layer1_outputs(711) <= not (a xor b);
    layer1_outputs(712) <= a xor b;
    layer1_outputs(713) <= not a or b;
    layer1_outputs(714) <= a and not b;
    layer1_outputs(715) <= b and not a;
    layer1_outputs(716) <= a;
    layer1_outputs(717) <= a and b;
    layer1_outputs(718) <= a and b;
    layer1_outputs(719) <= a xor b;
    layer1_outputs(720) <= b;
    layer1_outputs(721) <= not a or b;
    layer1_outputs(722) <= a or b;
    layer1_outputs(723) <= not b;
    layer1_outputs(724) <= not b;
    layer1_outputs(725) <= '1';
    layer1_outputs(726) <= b and not a;
    layer1_outputs(727) <= b;
    layer1_outputs(728) <= '1';
    layer1_outputs(729) <= not (a and b);
    layer1_outputs(730) <= not a or b;
    layer1_outputs(731) <= not (a or b);
    layer1_outputs(732) <= not a;
    layer1_outputs(733) <= not (a xor b);
    layer1_outputs(734) <= not a or b;
    layer1_outputs(735) <= a or b;
    layer1_outputs(736) <= b;
    layer1_outputs(737) <= not b;
    layer1_outputs(738) <= b;
    layer1_outputs(739) <= not b;
    layer1_outputs(740) <= a or b;
    layer1_outputs(741) <= b and not a;
    layer1_outputs(742) <= not a or b;
    layer1_outputs(743) <= a or b;
    layer1_outputs(744) <= a and b;
    layer1_outputs(745) <= not a or b;
    layer1_outputs(746) <= not (a and b);
    layer1_outputs(747) <= not (a or b);
    layer1_outputs(748) <= b and not a;
    layer1_outputs(749) <= a and not b;
    layer1_outputs(750) <= not (a or b);
    layer1_outputs(751) <= not (a or b);
    layer1_outputs(752) <= b;
    layer1_outputs(753) <= a and b;
    layer1_outputs(754) <= b;
    layer1_outputs(755) <= not a;
    layer1_outputs(756) <= a or b;
    layer1_outputs(757) <= not a;
    layer1_outputs(758) <= not (a or b);
    layer1_outputs(759) <= not b;
    layer1_outputs(760) <= not b or a;
    layer1_outputs(761) <= b and not a;
    layer1_outputs(762) <= b;
    layer1_outputs(763) <= not b;
    layer1_outputs(764) <= not b or a;
    layer1_outputs(765) <= not (a or b);
    layer1_outputs(766) <= not a;
    layer1_outputs(767) <= not (a or b);
    layer1_outputs(768) <= not b;
    layer1_outputs(769) <= '0';
    layer1_outputs(770) <= not (a xor b);
    layer1_outputs(771) <= not b;
    layer1_outputs(772) <= b;
    layer1_outputs(773) <= b;
    layer1_outputs(774) <= a and not b;
    layer1_outputs(775) <= b;
    layer1_outputs(776) <= a;
    layer1_outputs(777) <= b and not a;
    layer1_outputs(778) <= not a or b;
    layer1_outputs(779) <= a;
    layer1_outputs(780) <= not a or b;
    layer1_outputs(781) <= a and not b;
    layer1_outputs(782) <= a or b;
    layer1_outputs(783) <= not b;
    layer1_outputs(784) <= a or b;
    layer1_outputs(785) <= a or b;
    layer1_outputs(786) <= not a;
    layer1_outputs(787) <= '0';
    layer1_outputs(788) <= not (a or b);
    layer1_outputs(789) <= a and not b;
    layer1_outputs(790) <= not b;
    layer1_outputs(791) <= '0';
    layer1_outputs(792) <= b and not a;
    layer1_outputs(793) <= a or b;
    layer1_outputs(794) <= not a;
    layer1_outputs(795) <= not a or b;
    layer1_outputs(796) <= a;
    layer1_outputs(797) <= not b;
    layer1_outputs(798) <= not a;
    layer1_outputs(799) <= not (a and b);
    layer1_outputs(800) <= '0';
    layer1_outputs(801) <= b and not a;
    layer1_outputs(802) <= '1';
    layer1_outputs(803) <= a and b;
    layer1_outputs(804) <= not b;
    layer1_outputs(805) <= b;
    layer1_outputs(806) <= '1';
    layer1_outputs(807) <= not (a and b);
    layer1_outputs(808) <= not (a xor b);
    layer1_outputs(809) <= not b;
    layer1_outputs(810) <= b and not a;
    layer1_outputs(811) <= a or b;
    layer1_outputs(812) <= not (a and b);
    layer1_outputs(813) <= not a or b;
    layer1_outputs(814) <= a and not b;
    layer1_outputs(815) <= not (a and b);
    layer1_outputs(816) <= not a or b;
    layer1_outputs(817) <= not a or b;
    layer1_outputs(818) <= a;
    layer1_outputs(819) <= b and not a;
    layer1_outputs(820) <= not a;
    layer1_outputs(821) <= '1';
    layer1_outputs(822) <= not a or b;
    layer1_outputs(823) <= not a;
    layer1_outputs(824) <= '0';
    layer1_outputs(825) <= '1';
    layer1_outputs(826) <= '0';
    layer1_outputs(827) <= not (a and b);
    layer1_outputs(828) <= '0';
    layer1_outputs(829) <= a;
    layer1_outputs(830) <= not b or a;
    layer1_outputs(831) <= '1';
    layer1_outputs(832) <= not b;
    layer1_outputs(833) <= a xor b;
    layer1_outputs(834) <= not (a or b);
    layer1_outputs(835) <= not (a and b);
    layer1_outputs(836) <= not b;
    layer1_outputs(837) <= a xor b;
    layer1_outputs(838) <= not b or a;
    layer1_outputs(839) <= a;
    layer1_outputs(840) <= a;
    layer1_outputs(841) <= not b;
    layer1_outputs(842) <= not b;
    layer1_outputs(843) <= a and b;
    layer1_outputs(844) <= b;
    layer1_outputs(845) <= a and not b;
    layer1_outputs(846) <= '0';
    layer1_outputs(847) <= not a or b;
    layer1_outputs(848) <= not b;
    layer1_outputs(849) <= not a or b;
    layer1_outputs(850) <= b and not a;
    layer1_outputs(851) <= '0';
    layer1_outputs(852) <= not (a xor b);
    layer1_outputs(853) <= not (a and b);
    layer1_outputs(854) <= '0';
    layer1_outputs(855) <= '1';
    layer1_outputs(856) <= a and not b;
    layer1_outputs(857) <= not a;
    layer1_outputs(858) <= not a or b;
    layer1_outputs(859) <= not b or a;
    layer1_outputs(860) <= not (a and b);
    layer1_outputs(861) <= not a;
    layer1_outputs(862) <= a and b;
    layer1_outputs(863) <= not b or a;
    layer1_outputs(864) <= a;
    layer1_outputs(865) <= b;
    layer1_outputs(866) <= not (a xor b);
    layer1_outputs(867) <= a or b;
    layer1_outputs(868) <= not (a and b);
    layer1_outputs(869) <= b;
    layer1_outputs(870) <= not b;
    layer1_outputs(871) <= not (a and b);
    layer1_outputs(872) <= a and not b;
    layer1_outputs(873) <= not b;
    layer1_outputs(874) <= not a or b;
    layer1_outputs(875) <= a and not b;
    layer1_outputs(876) <= not (a or b);
    layer1_outputs(877) <= a or b;
    layer1_outputs(878) <= not a;
    layer1_outputs(879) <= a;
    layer1_outputs(880) <= not (a and b);
    layer1_outputs(881) <= b and not a;
    layer1_outputs(882) <= not b or a;
    layer1_outputs(883) <= not a or b;
    layer1_outputs(884) <= not a;
    layer1_outputs(885) <= not a;
    layer1_outputs(886) <= not (a and b);
    layer1_outputs(887) <= b;
    layer1_outputs(888) <= '0';
    layer1_outputs(889) <= not b;
    layer1_outputs(890) <= a xor b;
    layer1_outputs(891) <= a or b;
    layer1_outputs(892) <= a;
    layer1_outputs(893) <= not a;
    layer1_outputs(894) <= '0';
    layer1_outputs(895) <= not a;
    layer1_outputs(896) <= a and not b;
    layer1_outputs(897) <= '0';
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= not b or a;
    layer1_outputs(900) <= not (a or b);
    layer1_outputs(901) <= not (a or b);
    layer1_outputs(902) <= not a or b;
    layer1_outputs(903) <= not a;
    layer1_outputs(904) <= b and not a;
    layer1_outputs(905) <= not (a xor b);
    layer1_outputs(906) <= not b or a;
    layer1_outputs(907) <= not b or a;
    layer1_outputs(908) <= not b or a;
    layer1_outputs(909) <= b and not a;
    layer1_outputs(910) <= not a;
    layer1_outputs(911) <= not (a or b);
    layer1_outputs(912) <= a xor b;
    layer1_outputs(913) <= not a or b;
    layer1_outputs(914) <= a and not b;
    layer1_outputs(915) <= a or b;
    layer1_outputs(916) <= b and not a;
    layer1_outputs(917) <= b;
    layer1_outputs(918) <= not a or b;
    layer1_outputs(919) <= a and not b;
    layer1_outputs(920) <= not (a or b);
    layer1_outputs(921) <= a;
    layer1_outputs(922) <= a and b;
    layer1_outputs(923) <= not b or a;
    layer1_outputs(924) <= not (a and b);
    layer1_outputs(925) <= a and not b;
    layer1_outputs(926) <= not (a and b);
    layer1_outputs(927) <= not b;
    layer1_outputs(928) <= not (a xor b);
    layer1_outputs(929) <= a and not b;
    layer1_outputs(930) <= a or b;
    layer1_outputs(931) <= not (a and b);
    layer1_outputs(932) <= '0';
    layer1_outputs(933) <= not (a xor b);
    layer1_outputs(934) <= not a or b;
    layer1_outputs(935) <= a;
    layer1_outputs(936) <= '0';
    layer1_outputs(937) <= not (a xor b);
    layer1_outputs(938) <= not b or a;
    layer1_outputs(939) <= not b or a;
    layer1_outputs(940) <= a;
    layer1_outputs(941) <= not (a or b);
    layer1_outputs(942) <= '1';
    layer1_outputs(943) <= '1';
    layer1_outputs(944) <= not b or a;
    layer1_outputs(945) <= b;
    layer1_outputs(946) <= '1';
    layer1_outputs(947) <= not b or a;
    layer1_outputs(948) <= not b;
    layer1_outputs(949) <= a;
    layer1_outputs(950) <= '1';
    layer1_outputs(951) <= b and not a;
    layer1_outputs(952) <= not (a and b);
    layer1_outputs(953) <= b and not a;
    layer1_outputs(954) <= '0';
    layer1_outputs(955) <= a;
    layer1_outputs(956) <= not b;
    layer1_outputs(957) <= b;
    layer1_outputs(958) <= '1';
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= '0';
    layer1_outputs(961) <= not b or a;
    layer1_outputs(962) <= a xor b;
    layer1_outputs(963) <= a;
    layer1_outputs(964) <= not (a or b);
    layer1_outputs(965) <= not b;
    layer1_outputs(966) <= '0';
    layer1_outputs(967) <= a or b;
    layer1_outputs(968) <= not (a or b);
    layer1_outputs(969) <= not a or b;
    layer1_outputs(970) <= not (a or b);
    layer1_outputs(971) <= a or b;
    layer1_outputs(972) <= not b or a;
    layer1_outputs(973) <= not b;
    layer1_outputs(974) <= a xor b;
    layer1_outputs(975) <= '0';
    layer1_outputs(976) <= a and b;
    layer1_outputs(977) <= a or b;
    layer1_outputs(978) <= not b;
    layer1_outputs(979) <= not a;
    layer1_outputs(980) <= '1';
    layer1_outputs(981) <= not b or a;
    layer1_outputs(982) <= '1';
    layer1_outputs(983) <= b and not a;
    layer1_outputs(984) <= not b;
    layer1_outputs(985) <= a or b;
    layer1_outputs(986) <= '1';
    layer1_outputs(987) <= b;
    layer1_outputs(988) <= b;
    layer1_outputs(989) <= not b or a;
    layer1_outputs(990) <= not (a or b);
    layer1_outputs(991) <= not b;
    layer1_outputs(992) <= b;
    layer1_outputs(993) <= not b;
    layer1_outputs(994) <= a;
    layer1_outputs(995) <= not b;
    layer1_outputs(996) <= a or b;
    layer1_outputs(997) <= not (a or b);
    layer1_outputs(998) <= not a or b;
    layer1_outputs(999) <= a or b;
    layer1_outputs(1000) <= a and b;
    layer1_outputs(1001) <= not b;
    layer1_outputs(1002) <= not a;
    layer1_outputs(1003) <= a and b;
    layer1_outputs(1004) <= not (a or b);
    layer1_outputs(1005) <= not b;
    layer1_outputs(1006) <= not a or b;
    layer1_outputs(1007) <= '0';
    layer1_outputs(1008) <= b and not a;
    layer1_outputs(1009) <= b;
    layer1_outputs(1010) <= a xor b;
    layer1_outputs(1011) <= not a;
    layer1_outputs(1012) <= not b or a;
    layer1_outputs(1013) <= a or b;
    layer1_outputs(1014) <= not b;
    layer1_outputs(1015) <= a and b;
    layer1_outputs(1016) <= '0';
    layer1_outputs(1017) <= '1';
    layer1_outputs(1018) <= '0';
    layer1_outputs(1019) <= not a;
    layer1_outputs(1020) <= not (a xor b);
    layer1_outputs(1021) <= not a or b;
    layer1_outputs(1022) <= a xor b;
    layer1_outputs(1023) <= not (a xor b);
    layer1_outputs(1024) <= a and b;
    layer1_outputs(1025) <= a xor b;
    layer1_outputs(1026) <= a and b;
    layer1_outputs(1027) <= a and not b;
    layer1_outputs(1028) <= a;
    layer1_outputs(1029) <= a or b;
    layer1_outputs(1030) <= b and not a;
    layer1_outputs(1031) <= a;
    layer1_outputs(1032) <= a and not b;
    layer1_outputs(1033) <= b;
    layer1_outputs(1034) <= not b or a;
    layer1_outputs(1035) <= a;
    layer1_outputs(1036) <= not b;
    layer1_outputs(1037) <= '1';
    layer1_outputs(1038) <= b;
    layer1_outputs(1039) <= not a or b;
    layer1_outputs(1040) <= not a or b;
    layer1_outputs(1041) <= a and b;
    layer1_outputs(1042) <= a;
    layer1_outputs(1043) <= a or b;
    layer1_outputs(1044) <= not b or a;
    layer1_outputs(1045) <= not (a and b);
    layer1_outputs(1046) <= not (a xor b);
    layer1_outputs(1047) <= not (a and b);
    layer1_outputs(1048) <= a xor b;
    layer1_outputs(1049) <= not a or b;
    layer1_outputs(1050) <= not (a xor b);
    layer1_outputs(1051) <= not a or b;
    layer1_outputs(1052) <= a and b;
    layer1_outputs(1053) <= not b;
    layer1_outputs(1054) <= a or b;
    layer1_outputs(1055) <= b and not a;
    layer1_outputs(1056) <= not a or b;
    layer1_outputs(1057) <= not (a and b);
    layer1_outputs(1058) <= not a;
    layer1_outputs(1059) <= not b or a;
    layer1_outputs(1060) <= not (a and b);
    layer1_outputs(1061) <= a xor b;
    layer1_outputs(1062) <= '1';
    layer1_outputs(1063) <= b and not a;
    layer1_outputs(1064) <= not (a xor b);
    layer1_outputs(1065) <= '0';
    layer1_outputs(1066) <= a or b;
    layer1_outputs(1067) <= not b or a;
    layer1_outputs(1068) <= not a;
    layer1_outputs(1069) <= b and not a;
    layer1_outputs(1070) <= not (a or b);
    layer1_outputs(1071) <= '1';
    layer1_outputs(1072) <= not (a and b);
    layer1_outputs(1073) <= a and b;
    layer1_outputs(1074) <= a or b;
    layer1_outputs(1075) <= b;
    layer1_outputs(1076) <= not (a or b);
    layer1_outputs(1077) <= not a or b;
    layer1_outputs(1078) <= a xor b;
    layer1_outputs(1079) <= not (a or b);
    layer1_outputs(1080) <= not (a or b);
    layer1_outputs(1081) <= not a or b;
    layer1_outputs(1082) <= not (a xor b);
    layer1_outputs(1083) <= not a or b;
    layer1_outputs(1084) <= a or b;
    layer1_outputs(1085) <= not b;
    layer1_outputs(1086) <= not (a or b);
    layer1_outputs(1087) <= a and not b;
    layer1_outputs(1088) <= b and not a;
    layer1_outputs(1089) <= not b;
    layer1_outputs(1090) <= b and not a;
    layer1_outputs(1091) <= a and b;
    layer1_outputs(1092) <= b;
    layer1_outputs(1093) <= '0';
    layer1_outputs(1094) <= a or b;
    layer1_outputs(1095) <= not a;
    layer1_outputs(1096) <= not (a xor b);
    layer1_outputs(1097) <= not b;
    layer1_outputs(1098) <= a and b;
    layer1_outputs(1099) <= not (a and b);
    layer1_outputs(1100) <= b;
    layer1_outputs(1101) <= a or b;
    layer1_outputs(1102) <= a;
    layer1_outputs(1103) <= b and not a;
    layer1_outputs(1104) <= a;
    layer1_outputs(1105) <= a and b;
    layer1_outputs(1106) <= a and not b;
    layer1_outputs(1107) <= not b or a;
    layer1_outputs(1108) <= b;
    layer1_outputs(1109) <= not a;
    layer1_outputs(1110) <= not b;
    layer1_outputs(1111) <= a;
    layer1_outputs(1112) <= a and not b;
    layer1_outputs(1113) <= not (a and b);
    layer1_outputs(1114) <= b;
    layer1_outputs(1115) <= a or b;
    layer1_outputs(1116) <= b;
    layer1_outputs(1117) <= not a or b;
    layer1_outputs(1118) <= not (a or b);
    layer1_outputs(1119) <= a and not b;
    layer1_outputs(1120) <= a or b;
    layer1_outputs(1121) <= a or b;
    layer1_outputs(1122) <= a or b;
    layer1_outputs(1123) <= not b;
    layer1_outputs(1124) <= a and not b;
    layer1_outputs(1125) <= a and not b;
    layer1_outputs(1126) <= not a;
    layer1_outputs(1127) <= a or b;
    layer1_outputs(1128) <= not b or a;
    layer1_outputs(1129) <= not b;
    layer1_outputs(1130) <= not a;
    layer1_outputs(1131) <= not (a and b);
    layer1_outputs(1132) <= '0';
    layer1_outputs(1133) <= b and not a;
    layer1_outputs(1134) <= not (a and b);
    layer1_outputs(1135) <= not (a and b);
    layer1_outputs(1136) <= a and not b;
    layer1_outputs(1137) <= a and b;
    layer1_outputs(1138) <= a and not b;
    layer1_outputs(1139) <= a or b;
    layer1_outputs(1140) <= b;
    layer1_outputs(1141) <= not b;
    layer1_outputs(1142) <= a xor b;
    layer1_outputs(1143) <= not a;
    layer1_outputs(1144) <= a or b;
    layer1_outputs(1145) <= not b;
    layer1_outputs(1146) <= '1';
    layer1_outputs(1147) <= a and b;
    layer1_outputs(1148) <= not b or a;
    layer1_outputs(1149) <= '1';
    layer1_outputs(1150) <= not (a and b);
    layer1_outputs(1151) <= not (a xor b);
    layer1_outputs(1152) <= a and not b;
    layer1_outputs(1153) <= not (a and b);
    layer1_outputs(1154) <= a;
    layer1_outputs(1155) <= a or b;
    layer1_outputs(1156) <= a;
    layer1_outputs(1157) <= a and not b;
    layer1_outputs(1158) <= not a;
    layer1_outputs(1159) <= not b;
    layer1_outputs(1160) <= a;
    layer1_outputs(1161) <= '1';
    layer1_outputs(1162) <= b;
    layer1_outputs(1163) <= '1';
    layer1_outputs(1164) <= b;
    layer1_outputs(1165) <= '1';
    layer1_outputs(1166) <= not (a or b);
    layer1_outputs(1167) <= a or b;
    layer1_outputs(1168) <= '0';
    layer1_outputs(1169) <= a and not b;
    layer1_outputs(1170) <= a and b;
    layer1_outputs(1171) <= a;
    layer1_outputs(1172) <= not b;
    layer1_outputs(1173) <= a or b;
    layer1_outputs(1174) <= not b;
    layer1_outputs(1175) <= not a;
    layer1_outputs(1176) <= b;
    layer1_outputs(1177) <= not b;
    layer1_outputs(1178) <= not (a or b);
    layer1_outputs(1179) <= '0';
    layer1_outputs(1180) <= not (a and b);
    layer1_outputs(1181) <= a and b;
    layer1_outputs(1182) <= a;
    layer1_outputs(1183) <= '0';
    layer1_outputs(1184) <= '0';
    layer1_outputs(1185) <= a or b;
    layer1_outputs(1186) <= a and not b;
    layer1_outputs(1187) <= b and not a;
    layer1_outputs(1188) <= '1';
    layer1_outputs(1189) <= a and b;
    layer1_outputs(1190) <= not (a and b);
    layer1_outputs(1191) <= a and not b;
    layer1_outputs(1192) <= not a or b;
    layer1_outputs(1193) <= not b or a;
    layer1_outputs(1194) <= a;
    layer1_outputs(1195) <= not (a or b);
    layer1_outputs(1196) <= '0';
    layer1_outputs(1197) <= not b;
    layer1_outputs(1198) <= a and not b;
    layer1_outputs(1199) <= not a;
    layer1_outputs(1200) <= not (a and b);
    layer1_outputs(1201) <= not b;
    layer1_outputs(1202) <= not b or a;
    layer1_outputs(1203) <= a and b;
    layer1_outputs(1204) <= a;
    layer1_outputs(1205) <= '1';
    layer1_outputs(1206) <= a;
    layer1_outputs(1207) <= not a or b;
    layer1_outputs(1208) <= not a or b;
    layer1_outputs(1209) <= b and not a;
    layer1_outputs(1210) <= not a or b;
    layer1_outputs(1211) <= a and not b;
    layer1_outputs(1212) <= a and not b;
    layer1_outputs(1213) <= a and b;
    layer1_outputs(1214) <= '1';
    layer1_outputs(1215) <= not (a and b);
    layer1_outputs(1216) <= not a or b;
    layer1_outputs(1217) <= not a or b;
    layer1_outputs(1218) <= '1';
    layer1_outputs(1219) <= not (a and b);
    layer1_outputs(1220) <= not (a or b);
    layer1_outputs(1221) <= '1';
    layer1_outputs(1222) <= a and b;
    layer1_outputs(1223) <= not (a and b);
    layer1_outputs(1224) <= '1';
    layer1_outputs(1225) <= b and not a;
    layer1_outputs(1226) <= b and not a;
    layer1_outputs(1227) <= not (a or b);
    layer1_outputs(1228) <= not a;
    layer1_outputs(1229) <= a and not b;
    layer1_outputs(1230) <= '0';
    layer1_outputs(1231) <= not (a and b);
    layer1_outputs(1232) <= b and not a;
    layer1_outputs(1233) <= not (a or b);
    layer1_outputs(1234) <= not b or a;
    layer1_outputs(1235) <= '0';
    layer1_outputs(1236) <= not (a or b);
    layer1_outputs(1237) <= a and b;
    layer1_outputs(1238) <= not a or b;
    layer1_outputs(1239) <= '0';
    layer1_outputs(1240) <= not (a and b);
    layer1_outputs(1241) <= b and not a;
    layer1_outputs(1242) <= a and not b;
    layer1_outputs(1243) <= a xor b;
    layer1_outputs(1244) <= not a or b;
    layer1_outputs(1245) <= a or b;
    layer1_outputs(1246) <= a and b;
    layer1_outputs(1247) <= not b;
    layer1_outputs(1248) <= not (a and b);
    layer1_outputs(1249) <= b and not a;
    layer1_outputs(1250) <= '0';
    layer1_outputs(1251) <= not b;
    layer1_outputs(1252) <= b;
    layer1_outputs(1253) <= '1';
    layer1_outputs(1254) <= a;
    layer1_outputs(1255) <= '1';
    layer1_outputs(1256) <= b;
    layer1_outputs(1257) <= a xor b;
    layer1_outputs(1258) <= a;
    layer1_outputs(1259) <= a and not b;
    layer1_outputs(1260) <= a;
    layer1_outputs(1261) <= not b or a;
    layer1_outputs(1262) <= b;
    layer1_outputs(1263) <= not a or b;
    layer1_outputs(1264) <= a or b;
    layer1_outputs(1265) <= a and b;
    layer1_outputs(1266) <= b and not a;
    layer1_outputs(1267) <= not b;
    layer1_outputs(1268) <= a;
    layer1_outputs(1269) <= not a;
    layer1_outputs(1270) <= '0';
    layer1_outputs(1271) <= a and b;
    layer1_outputs(1272) <= a or b;
    layer1_outputs(1273) <= '1';
    layer1_outputs(1274) <= b and not a;
    layer1_outputs(1275) <= not a or b;
    layer1_outputs(1276) <= a;
    layer1_outputs(1277) <= a and b;
    layer1_outputs(1278) <= a and b;
    layer1_outputs(1279) <= a and not b;
    layer1_outputs(1280) <= b and not a;
    layer1_outputs(1281) <= not b or a;
    layer1_outputs(1282) <= '0';
    layer1_outputs(1283) <= b;
    layer1_outputs(1284) <= not b or a;
    layer1_outputs(1285) <= b;
    layer1_outputs(1286) <= b;
    layer1_outputs(1287) <= not (a and b);
    layer1_outputs(1288) <= not a;
    layer1_outputs(1289) <= a and b;
    layer1_outputs(1290) <= b and not a;
    layer1_outputs(1291) <= not a or b;
    layer1_outputs(1292) <= not a or b;
    layer1_outputs(1293) <= '0';
    layer1_outputs(1294) <= not b;
    layer1_outputs(1295) <= a or b;
    layer1_outputs(1296) <= not (a or b);
    layer1_outputs(1297) <= not b;
    layer1_outputs(1298) <= b and not a;
    layer1_outputs(1299) <= not b;
    layer1_outputs(1300) <= b;
    layer1_outputs(1301) <= not b;
    layer1_outputs(1302) <= not a or b;
    layer1_outputs(1303) <= not (a and b);
    layer1_outputs(1304) <= not (a or b);
    layer1_outputs(1305) <= a or b;
    layer1_outputs(1306) <= b and not a;
    layer1_outputs(1307) <= not (a and b);
    layer1_outputs(1308) <= a and b;
    layer1_outputs(1309) <= a and b;
    layer1_outputs(1310) <= not b;
    layer1_outputs(1311) <= '0';
    layer1_outputs(1312) <= a and not b;
    layer1_outputs(1313) <= not a or b;
    layer1_outputs(1314) <= a;
    layer1_outputs(1315) <= a and not b;
    layer1_outputs(1316) <= not a;
    layer1_outputs(1317) <= not b or a;
    layer1_outputs(1318) <= b;
    layer1_outputs(1319) <= a;
    layer1_outputs(1320) <= not b or a;
    layer1_outputs(1321) <= not b or a;
    layer1_outputs(1322) <= not a;
    layer1_outputs(1323) <= b and not a;
    layer1_outputs(1324) <= not (a or b);
    layer1_outputs(1325) <= b;
    layer1_outputs(1326) <= b;
    layer1_outputs(1327) <= '1';
    layer1_outputs(1328) <= a and not b;
    layer1_outputs(1329) <= not (a and b);
    layer1_outputs(1330) <= a and b;
    layer1_outputs(1331) <= not a;
    layer1_outputs(1332) <= b and not a;
    layer1_outputs(1333) <= not (a or b);
    layer1_outputs(1334) <= not (a and b);
    layer1_outputs(1335) <= '0';
    layer1_outputs(1336) <= '1';
    layer1_outputs(1337) <= '1';
    layer1_outputs(1338) <= not (a or b);
    layer1_outputs(1339) <= a xor b;
    layer1_outputs(1340) <= not (a xor b);
    layer1_outputs(1341) <= not b;
    layer1_outputs(1342) <= not b;
    layer1_outputs(1343) <= a or b;
    layer1_outputs(1344) <= not (a and b);
    layer1_outputs(1345) <= not (a and b);
    layer1_outputs(1346) <= a xor b;
    layer1_outputs(1347) <= not (a and b);
    layer1_outputs(1348) <= not b;
    layer1_outputs(1349) <= not (a and b);
    layer1_outputs(1350) <= a;
    layer1_outputs(1351) <= '1';
    layer1_outputs(1352) <= b and not a;
    layer1_outputs(1353) <= a and not b;
    layer1_outputs(1354) <= not (a xor b);
    layer1_outputs(1355) <= not b;
    layer1_outputs(1356) <= b;
    layer1_outputs(1357) <= a;
    layer1_outputs(1358) <= not b;
    layer1_outputs(1359) <= not b;
    layer1_outputs(1360) <= a xor b;
    layer1_outputs(1361) <= '0';
    layer1_outputs(1362) <= '1';
    layer1_outputs(1363) <= not (a and b);
    layer1_outputs(1364) <= a;
    layer1_outputs(1365) <= not a;
    layer1_outputs(1366) <= not a or b;
    layer1_outputs(1367) <= a;
    layer1_outputs(1368) <= '1';
    layer1_outputs(1369) <= b;
    layer1_outputs(1370) <= a and b;
    layer1_outputs(1371) <= not a or b;
    layer1_outputs(1372) <= not a;
    layer1_outputs(1373) <= not (a or b);
    layer1_outputs(1374) <= not b;
    layer1_outputs(1375) <= not a;
    layer1_outputs(1376) <= a xor b;
    layer1_outputs(1377) <= b;
    layer1_outputs(1378) <= not (a or b);
    layer1_outputs(1379) <= b and not a;
    layer1_outputs(1380) <= a and not b;
    layer1_outputs(1381) <= a and b;
    layer1_outputs(1382) <= a;
    layer1_outputs(1383) <= not a;
    layer1_outputs(1384) <= a and not b;
    layer1_outputs(1385) <= a and not b;
    layer1_outputs(1386) <= b;
    layer1_outputs(1387) <= not b or a;
    layer1_outputs(1388) <= b and not a;
    layer1_outputs(1389) <= a;
    layer1_outputs(1390) <= a xor b;
    layer1_outputs(1391) <= not (a or b);
    layer1_outputs(1392) <= b and not a;
    layer1_outputs(1393) <= b;
    layer1_outputs(1394) <= not (a and b);
    layer1_outputs(1395) <= not (a or b);
    layer1_outputs(1396) <= '1';
    layer1_outputs(1397) <= '1';
    layer1_outputs(1398) <= a or b;
    layer1_outputs(1399) <= a;
    layer1_outputs(1400) <= not (a xor b);
    layer1_outputs(1401) <= a and b;
    layer1_outputs(1402) <= not (a and b);
    layer1_outputs(1403) <= a and b;
    layer1_outputs(1404) <= not b;
    layer1_outputs(1405) <= a and not b;
    layer1_outputs(1406) <= not b;
    layer1_outputs(1407) <= '0';
    layer1_outputs(1408) <= '0';
    layer1_outputs(1409) <= not a;
    layer1_outputs(1410) <= a;
    layer1_outputs(1411) <= a or b;
    layer1_outputs(1412) <= not a or b;
    layer1_outputs(1413) <= not (a or b);
    layer1_outputs(1414) <= not a or b;
    layer1_outputs(1415) <= a and b;
    layer1_outputs(1416) <= '0';
    layer1_outputs(1417) <= a;
    layer1_outputs(1418) <= not b;
    layer1_outputs(1419) <= a;
    layer1_outputs(1420) <= not b or a;
    layer1_outputs(1421) <= b and not a;
    layer1_outputs(1422) <= a and not b;
    layer1_outputs(1423) <= a xor b;
    layer1_outputs(1424) <= '0';
    layer1_outputs(1425) <= a and b;
    layer1_outputs(1426) <= not (a and b);
    layer1_outputs(1427) <= not (a or b);
    layer1_outputs(1428) <= not (a or b);
    layer1_outputs(1429) <= not (a and b);
    layer1_outputs(1430) <= a or b;
    layer1_outputs(1431) <= a or b;
    layer1_outputs(1432) <= not (a or b);
    layer1_outputs(1433) <= a;
    layer1_outputs(1434) <= b and not a;
    layer1_outputs(1435) <= b;
    layer1_outputs(1436) <= not (a and b);
    layer1_outputs(1437) <= b;
    layer1_outputs(1438) <= b;
    layer1_outputs(1439) <= a and b;
    layer1_outputs(1440) <= a and b;
    layer1_outputs(1441) <= a;
    layer1_outputs(1442) <= not b or a;
    layer1_outputs(1443) <= not a;
    layer1_outputs(1444) <= not (a xor b);
    layer1_outputs(1445) <= not a;
    layer1_outputs(1446) <= not (a or b);
    layer1_outputs(1447) <= a;
    layer1_outputs(1448) <= not a;
    layer1_outputs(1449) <= '1';
    layer1_outputs(1450) <= b and not a;
    layer1_outputs(1451) <= not a or b;
    layer1_outputs(1452) <= not b;
    layer1_outputs(1453) <= not (a xor b);
    layer1_outputs(1454) <= a;
    layer1_outputs(1455) <= not a or b;
    layer1_outputs(1456) <= not a;
    layer1_outputs(1457) <= not a;
    layer1_outputs(1458) <= not b or a;
    layer1_outputs(1459) <= not (a xor b);
    layer1_outputs(1460) <= a or b;
    layer1_outputs(1461) <= not b or a;
    layer1_outputs(1462) <= not b or a;
    layer1_outputs(1463) <= a or b;
    layer1_outputs(1464) <= not (a and b);
    layer1_outputs(1465) <= not (a xor b);
    layer1_outputs(1466) <= '1';
    layer1_outputs(1467) <= not b or a;
    layer1_outputs(1468) <= '1';
    layer1_outputs(1469) <= not b or a;
    layer1_outputs(1470) <= not b;
    layer1_outputs(1471) <= '1';
    layer1_outputs(1472) <= a xor b;
    layer1_outputs(1473) <= not a or b;
    layer1_outputs(1474) <= not (a and b);
    layer1_outputs(1475) <= not (a and b);
    layer1_outputs(1476) <= not a;
    layer1_outputs(1477) <= not (a and b);
    layer1_outputs(1478) <= not (a and b);
    layer1_outputs(1479) <= a;
    layer1_outputs(1480) <= a and b;
    layer1_outputs(1481) <= not b;
    layer1_outputs(1482) <= not a;
    layer1_outputs(1483) <= '1';
    layer1_outputs(1484) <= not a or b;
    layer1_outputs(1485) <= a and not b;
    layer1_outputs(1486) <= b;
    layer1_outputs(1487) <= b and not a;
    layer1_outputs(1488) <= '0';
    layer1_outputs(1489) <= '1';
    layer1_outputs(1490) <= not a;
    layer1_outputs(1491) <= not (a and b);
    layer1_outputs(1492) <= not (a and b);
    layer1_outputs(1493) <= not (a and b);
    layer1_outputs(1494) <= a;
    layer1_outputs(1495) <= not a or b;
    layer1_outputs(1496) <= not (a or b);
    layer1_outputs(1497) <= '1';
    layer1_outputs(1498) <= a;
    layer1_outputs(1499) <= b and not a;
    layer1_outputs(1500) <= not a;
    layer1_outputs(1501) <= a and b;
    layer1_outputs(1502) <= not (a or b);
    layer1_outputs(1503) <= b and not a;
    layer1_outputs(1504) <= not (a and b);
    layer1_outputs(1505) <= not b;
    layer1_outputs(1506) <= b;
    layer1_outputs(1507) <= not b;
    layer1_outputs(1508) <= not (a or b);
    layer1_outputs(1509) <= a and not b;
    layer1_outputs(1510) <= not b;
    layer1_outputs(1511) <= b and not a;
    layer1_outputs(1512) <= '1';
    layer1_outputs(1513) <= not a;
    layer1_outputs(1514) <= not (a and b);
    layer1_outputs(1515) <= b;
    layer1_outputs(1516) <= a;
    layer1_outputs(1517) <= b and not a;
    layer1_outputs(1518) <= a xor b;
    layer1_outputs(1519) <= b;
    layer1_outputs(1520) <= a xor b;
    layer1_outputs(1521) <= '0';
    layer1_outputs(1522) <= '0';
    layer1_outputs(1523) <= not b or a;
    layer1_outputs(1524) <= not (a xor b);
    layer1_outputs(1525) <= a or b;
    layer1_outputs(1526) <= a and not b;
    layer1_outputs(1527) <= a;
    layer1_outputs(1528) <= '1';
    layer1_outputs(1529) <= not a;
    layer1_outputs(1530) <= not a or b;
    layer1_outputs(1531) <= '1';
    layer1_outputs(1532) <= not a;
    layer1_outputs(1533) <= not (a or b);
    layer1_outputs(1534) <= not b or a;
    layer1_outputs(1535) <= a and b;
    layer1_outputs(1536) <= not b or a;
    layer1_outputs(1537) <= a;
    layer1_outputs(1538) <= a or b;
    layer1_outputs(1539) <= b;
    layer1_outputs(1540) <= not (a and b);
    layer1_outputs(1541) <= not (a and b);
    layer1_outputs(1542) <= b;
    layer1_outputs(1543) <= b;
    layer1_outputs(1544) <= not b;
    layer1_outputs(1545) <= not b;
    layer1_outputs(1546) <= a;
    layer1_outputs(1547) <= not (a and b);
    layer1_outputs(1548) <= not (a or b);
    layer1_outputs(1549) <= not a;
    layer1_outputs(1550) <= not a or b;
    layer1_outputs(1551) <= b;
    layer1_outputs(1552) <= not (a or b);
    layer1_outputs(1553) <= a and not b;
    layer1_outputs(1554) <= not (a or b);
    layer1_outputs(1555) <= a and not b;
    layer1_outputs(1556) <= not a or b;
    layer1_outputs(1557) <= not b or a;
    layer1_outputs(1558) <= not (a xor b);
    layer1_outputs(1559) <= b;
    layer1_outputs(1560) <= a or b;
    layer1_outputs(1561) <= b and not a;
    layer1_outputs(1562) <= a and not b;
    layer1_outputs(1563) <= b and not a;
    layer1_outputs(1564) <= b;
    layer1_outputs(1565) <= a xor b;
    layer1_outputs(1566) <= '1';
    layer1_outputs(1567) <= b;
    layer1_outputs(1568) <= a or b;
    layer1_outputs(1569) <= not b or a;
    layer1_outputs(1570) <= a and b;
    layer1_outputs(1571) <= a or b;
    layer1_outputs(1572) <= not b or a;
    layer1_outputs(1573) <= a and not b;
    layer1_outputs(1574) <= '0';
    layer1_outputs(1575) <= a and b;
    layer1_outputs(1576) <= not (a xor b);
    layer1_outputs(1577) <= '0';
    layer1_outputs(1578) <= b;
    layer1_outputs(1579) <= b;
    layer1_outputs(1580) <= not a;
    layer1_outputs(1581) <= '0';
    layer1_outputs(1582) <= not b;
    layer1_outputs(1583) <= a and not b;
    layer1_outputs(1584) <= a or b;
    layer1_outputs(1585) <= not b;
    layer1_outputs(1586) <= not (a and b);
    layer1_outputs(1587) <= a xor b;
    layer1_outputs(1588) <= not b or a;
    layer1_outputs(1589) <= not b;
    layer1_outputs(1590) <= a and not b;
    layer1_outputs(1591) <= not (a or b);
    layer1_outputs(1592) <= a and b;
    layer1_outputs(1593) <= not (a or b);
    layer1_outputs(1594) <= a and not b;
    layer1_outputs(1595) <= a or b;
    layer1_outputs(1596) <= not (a or b);
    layer1_outputs(1597) <= a or b;
    layer1_outputs(1598) <= not (a and b);
    layer1_outputs(1599) <= not a;
    layer1_outputs(1600) <= not (a or b);
    layer1_outputs(1601) <= not b or a;
    layer1_outputs(1602) <= not (a and b);
    layer1_outputs(1603) <= a;
    layer1_outputs(1604) <= not b;
    layer1_outputs(1605) <= '1';
    layer1_outputs(1606) <= not a or b;
    layer1_outputs(1607) <= '0';
    layer1_outputs(1608) <= not (a and b);
    layer1_outputs(1609) <= not (a and b);
    layer1_outputs(1610) <= not (a and b);
    layer1_outputs(1611) <= a and not b;
    layer1_outputs(1612) <= a;
    layer1_outputs(1613) <= not a or b;
    layer1_outputs(1614) <= not a;
    layer1_outputs(1615) <= a and not b;
    layer1_outputs(1616) <= b;
    layer1_outputs(1617) <= not a or b;
    layer1_outputs(1618) <= b and not a;
    layer1_outputs(1619) <= b and not a;
    layer1_outputs(1620) <= not (a and b);
    layer1_outputs(1621) <= b;
    layer1_outputs(1622) <= a and b;
    layer1_outputs(1623) <= b;
    layer1_outputs(1624) <= not b or a;
    layer1_outputs(1625) <= a or b;
    layer1_outputs(1626) <= a xor b;
    layer1_outputs(1627) <= b;
    layer1_outputs(1628) <= b;
    layer1_outputs(1629) <= not a or b;
    layer1_outputs(1630) <= not a or b;
    layer1_outputs(1631) <= not b or a;
    layer1_outputs(1632) <= not (a xor b);
    layer1_outputs(1633) <= a xor b;
    layer1_outputs(1634) <= a xor b;
    layer1_outputs(1635) <= a;
    layer1_outputs(1636) <= not a;
    layer1_outputs(1637) <= not (a and b);
    layer1_outputs(1638) <= a xor b;
    layer1_outputs(1639) <= b;
    layer1_outputs(1640) <= a and b;
    layer1_outputs(1641) <= a or b;
    layer1_outputs(1642) <= not a or b;
    layer1_outputs(1643) <= b;
    layer1_outputs(1644) <= not b;
    layer1_outputs(1645) <= b;
    layer1_outputs(1646) <= a and not b;
    layer1_outputs(1647) <= not b;
    layer1_outputs(1648) <= a and not b;
    layer1_outputs(1649) <= not a;
    layer1_outputs(1650) <= a and not b;
    layer1_outputs(1651) <= not (a and b);
    layer1_outputs(1652) <= not (a or b);
    layer1_outputs(1653) <= not b or a;
    layer1_outputs(1654) <= b and not a;
    layer1_outputs(1655) <= b;
    layer1_outputs(1656) <= '0';
    layer1_outputs(1657) <= a;
    layer1_outputs(1658) <= not a;
    layer1_outputs(1659) <= a or b;
    layer1_outputs(1660) <= not (a and b);
    layer1_outputs(1661) <= not b or a;
    layer1_outputs(1662) <= b;
    layer1_outputs(1663) <= b;
    layer1_outputs(1664) <= b;
    layer1_outputs(1665) <= not a;
    layer1_outputs(1666) <= not b or a;
    layer1_outputs(1667) <= b and not a;
    layer1_outputs(1668) <= not a or b;
    layer1_outputs(1669) <= not (a and b);
    layer1_outputs(1670) <= a;
    layer1_outputs(1671) <= '0';
    layer1_outputs(1672) <= not b;
    layer1_outputs(1673) <= not (a and b);
    layer1_outputs(1674) <= not (a or b);
    layer1_outputs(1675) <= not a;
    layer1_outputs(1676) <= a and not b;
    layer1_outputs(1677) <= not b;
    layer1_outputs(1678) <= a and b;
    layer1_outputs(1679) <= a or b;
    layer1_outputs(1680) <= a;
    layer1_outputs(1681) <= not a;
    layer1_outputs(1682) <= a xor b;
    layer1_outputs(1683) <= not a or b;
    layer1_outputs(1684) <= not b or a;
    layer1_outputs(1685) <= not b or a;
    layer1_outputs(1686) <= a or b;
    layer1_outputs(1687) <= b and not a;
    layer1_outputs(1688) <= b;
    layer1_outputs(1689) <= a;
    layer1_outputs(1690) <= '1';
    layer1_outputs(1691) <= not (a xor b);
    layer1_outputs(1692) <= '1';
    layer1_outputs(1693) <= not (a and b);
    layer1_outputs(1694) <= not (a or b);
    layer1_outputs(1695) <= b and not a;
    layer1_outputs(1696) <= not a;
    layer1_outputs(1697) <= a xor b;
    layer1_outputs(1698) <= not a or b;
    layer1_outputs(1699) <= a;
    layer1_outputs(1700) <= not a;
    layer1_outputs(1701) <= b;
    layer1_outputs(1702) <= not b;
    layer1_outputs(1703) <= not b or a;
    layer1_outputs(1704) <= not a;
    layer1_outputs(1705) <= b;
    layer1_outputs(1706) <= '1';
    layer1_outputs(1707) <= '1';
    layer1_outputs(1708) <= a and b;
    layer1_outputs(1709) <= b;
    layer1_outputs(1710) <= not b;
    layer1_outputs(1711) <= not (a or b);
    layer1_outputs(1712) <= a;
    layer1_outputs(1713) <= not (a xor b);
    layer1_outputs(1714) <= not (a or b);
    layer1_outputs(1715) <= not a;
    layer1_outputs(1716) <= a xor b;
    layer1_outputs(1717) <= '1';
    layer1_outputs(1718) <= a and not b;
    layer1_outputs(1719) <= not a;
    layer1_outputs(1720) <= not b or a;
    layer1_outputs(1721) <= a and b;
    layer1_outputs(1722) <= a;
    layer1_outputs(1723) <= a or b;
    layer1_outputs(1724) <= not (a and b);
    layer1_outputs(1725) <= b and not a;
    layer1_outputs(1726) <= not (a and b);
    layer1_outputs(1727) <= not b;
    layer1_outputs(1728) <= a;
    layer1_outputs(1729) <= not b or a;
    layer1_outputs(1730) <= not (a and b);
    layer1_outputs(1731) <= a xor b;
    layer1_outputs(1732) <= a and not b;
    layer1_outputs(1733) <= not (a and b);
    layer1_outputs(1734) <= not a;
    layer1_outputs(1735) <= not (a or b);
    layer1_outputs(1736) <= not a;
    layer1_outputs(1737) <= not b or a;
    layer1_outputs(1738) <= not b or a;
    layer1_outputs(1739) <= a xor b;
    layer1_outputs(1740) <= a and not b;
    layer1_outputs(1741) <= '0';
    layer1_outputs(1742) <= not b or a;
    layer1_outputs(1743) <= a and not b;
    layer1_outputs(1744) <= not b;
    layer1_outputs(1745) <= '0';
    layer1_outputs(1746) <= not a;
    layer1_outputs(1747) <= a and b;
    layer1_outputs(1748) <= '0';
    layer1_outputs(1749) <= b and not a;
    layer1_outputs(1750) <= '1';
    layer1_outputs(1751) <= not b;
    layer1_outputs(1752) <= a or b;
    layer1_outputs(1753) <= not a;
    layer1_outputs(1754) <= not (a or b);
    layer1_outputs(1755) <= b;
    layer1_outputs(1756) <= a and b;
    layer1_outputs(1757) <= b and not a;
    layer1_outputs(1758) <= b;
    layer1_outputs(1759) <= not a;
    layer1_outputs(1760) <= '1';
    layer1_outputs(1761) <= a or b;
    layer1_outputs(1762) <= b and not a;
    layer1_outputs(1763) <= b;
    layer1_outputs(1764) <= not a or b;
    layer1_outputs(1765) <= not a;
    layer1_outputs(1766) <= not b;
    layer1_outputs(1767) <= '0';
    layer1_outputs(1768) <= b and not a;
    layer1_outputs(1769) <= a and not b;
    layer1_outputs(1770) <= a and not b;
    layer1_outputs(1771) <= not (a or b);
    layer1_outputs(1772) <= a and b;
    layer1_outputs(1773) <= not b or a;
    layer1_outputs(1774) <= not (a and b);
    layer1_outputs(1775) <= not a;
    layer1_outputs(1776) <= a and not b;
    layer1_outputs(1777) <= '1';
    layer1_outputs(1778) <= '0';
    layer1_outputs(1779) <= not (a or b);
    layer1_outputs(1780) <= a and b;
    layer1_outputs(1781) <= b and not a;
    layer1_outputs(1782) <= '1';
    layer1_outputs(1783) <= b;
    layer1_outputs(1784) <= a and b;
    layer1_outputs(1785) <= not b;
    layer1_outputs(1786) <= b;
    layer1_outputs(1787) <= not (a xor b);
    layer1_outputs(1788) <= not (a or b);
    layer1_outputs(1789) <= not a;
    layer1_outputs(1790) <= not (a xor b);
    layer1_outputs(1791) <= b;
    layer1_outputs(1792) <= a xor b;
    layer1_outputs(1793) <= not b or a;
    layer1_outputs(1794) <= not b or a;
    layer1_outputs(1795) <= '0';
    layer1_outputs(1796) <= '1';
    layer1_outputs(1797) <= not a;
    layer1_outputs(1798) <= b;
    layer1_outputs(1799) <= not (a and b);
    layer1_outputs(1800) <= not a;
    layer1_outputs(1801) <= not b;
    layer1_outputs(1802) <= b and not a;
    layer1_outputs(1803) <= '0';
    layer1_outputs(1804) <= not a;
    layer1_outputs(1805) <= not a or b;
    layer1_outputs(1806) <= a;
    layer1_outputs(1807) <= a or b;
    layer1_outputs(1808) <= not a;
    layer1_outputs(1809) <= a and not b;
    layer1_outputs(1810) <= a and b;
    layer1_outputs(1811) <= b and not a;
    layer1_outputs(1812) <= b and not a;
    layer1_outputs(1813) <= not (a and b);
    layer1_outputs(1814) <= not (a and b);
    layer1_outputs(1815) <= not a;
    layer1_outputs(1816) <= b;
    layer1_outputs(1817) <= a and not b;
    layer1_outputs(1818) <= '0';
    layer1_outputs(1819) <= not a or b;
    layer1_outputs(1820) <= not a or b;
    layer1_outputs(1821) <= not (a xor b);
    layer1_outputs(1822) <= not b or a;
    layer1_outputs(1823) <= b;
    layer1_outputs(1824) <= a or b;
    layer1_outputs(1825) <= a and b;
    layer1_outputs(1826) <= a or b;
    layer1_outputs(1827) <= a;
    layer1_outputs(1828) <= not (a and b);
    layer1_outputs(1829) <= not b;
    layer1_outputs(1830) <= not (a or b);
    layer1_outputs(1831) <= not b or a;
    layer1_outputs(1832) <= a and not b;
    layer1_outputs(1833) <= b;
    layer1_outputs(1834) <= a and b;
    layer1_outputs(1835) <= a xor b;
    layer1_outputs(1836) <= not (a or b);
    layer1_outputs(1837) <= '0';
    layer1_outputs(1838) <= a and b;
    layer1_outputs(1839) <= '0';
    layer1_outputs(1840) <= not a;
    layer1_outputs(1841) <= b;
    layer1_outputs(1842) <= '1';
    layer1_outputs(1843) <= a or b;
    layer1_outputs(1844) <= not b or a;
    layer1_outputs(1845) <= not (a and b);
    layer1_outputs(1846) <= not (a and b);
    layer1_outputs(1847) <= b;
    layer1_outputs(1848) <= not (a and b);
    layer1_outputs(1849) <= not (a and b);
    layer1_outputs(1850) <= not b or a;
    layer1_outputs(1851) <= a or b;
    layer1_outputs(1852) <= not a;
    layer1_outputs(1853) <= a or b;
    layer1_outputs(1854) <= '0';
    layer1_outputs(1855) <= not b or a;
    layer1_outputs(1856) <= a;
    layer1_outputs(1857) <= not b or a;
    layer1_outputs(1858) <= not b;
    layer1_outputs(1859) <= not a;
    layer1_outputs(1860) <= '1';
    layer1_outputs(1861) <= a xor b;
    layer1_outputs(1862) <= not a or b;
    layer1_outputs(1863) <= a;
    layer1_outputs(1864) <= b;
    layer1_outputs(1865) <= a or b;
    layer1_outputs(1866) <= a or b;
    layer1_outputs(1867) <= not (a and b);
    layer1_outputs(1868) <= b and not a;
    layer1_outputs(1869) <= a;
    layer1_outputs(1870) <= '0';
    layer1_outputs(1871) <= not (a and b);
    layer1_outputs(1872) <= b and not a;
    layer1_outputs(1873) <= b;
    layer1_outputs(1874) <= a and not b;
    layer1_outputs(1875) <= not a;
    layer1_outputs(1876) <= not (a and b);
    layer1_outputs(1877) <= not (a xor b);
    layer1_outputs(1878) <= a and b;
    layer1_outputs(1879) <= not b;
    layer1_outputs(1880) <= not (a or b);
    layer1_outputs(1881) <= a;
    layer1_outputs(1882) <= not a or b;
    layer1_outputs(1883) <= not a;
    layer1_outputs(1884) <= not (a or b);
    layer1_outputs(1885) <= a and b;
    layer1_outputs(1886) <= '1';
    layer1_outputs(1887) <= not b;
    layer1_outputs(1888) <= not (a and b);
    layer1_outputs(1889) <= not b or a;
    layer1_outputs(1890) <= a;
    layer1_outputs(1891) <= a or b;
    layer1_outputs(1892) <= b;
    layer1_outputs(1893) <= not (a and b);
    layer1_outputs(1894) <= b;
    layer1_outputs(1895) <= not (a and b);
    layer1_outputs(1896) <= not (a and b);
    layer1_outputs(1897) <= a;
    layer1_outputs(1898) <= b and not a;
    layer1_outputs(1899) <= not a;
    layer1_outputs(1900) <= not (a xor b);
    layer1_outputs(1901) <= not (a or b);
    layer1_outputs(1902) <= '1';
    layer1_outputs(1903) <= '1';
    layer1_outputs(1904) <= not a or b;
    layer1_outputs(1905) <= not (a and b);
    layer1_outputs(1906) <= not a;
    layer1_outputs(1907) <= not (a and b);
    layer1_outputs(1908) <= b;
    layer1_outputs(1909) <= b;
    layer1_outputs(1910) <= not (a and b);
    layer1_outputs(1911) <= b;
    layer1_outputs(1912) <= '1';
    layer1_outputs(1913) <= '1';
    layer1_outputs(1914) <= '0';
    layer1_outputs(1915) <= not (a or b);
    layer1_outputs(1916) <= not a;
    layer1_outputs(1917) <= not b;
    layer1_outputs(1918) <= not (a xor b);
    layer1_outputs(1919) <= not (a and b);
    layer1_outputs(1920) <= not a or b;
    layer1_outputs(1921) <= not b;
    layer1_outputs(1922) <= a and not b;
    layer1_outputs(1923) <= b;
    layer1_outputs(1924) <= not (a xor b);
    layer1_outputs(1925) <= '0';
    layer1_outputs(1926) <= a xor b;
    layer1_outputs(1927) <= not b;
    layer1_outputs(1928) <= a and b;
    layer1_outputs(1929) <= not a;
    layer1_outputs(1930) <= '1';
    layer1_outputs(1931) <= a;
    layer1_outputs(1932) <= not (a or b);
    layer1_outputs(1933) <= b and not a;
    layer1_outputs(1934) <= a;
    layer1_outputs(1935) <= '0';
    layer1_outputs(1936) <= not a;
    layer1_outputs(1937) <= not a or b;
    layer1_outputs(1938) <= b;
    layer1_outputs(1939) <= a xor b;
    layer1_outputs(1940) <= a and b;
    layer1_outputs(1941) <= a and b;
    layer1_outputs(1942) <= not (a xor b);
    layer1_outputs(1943) <= a and b;
    layer1_outputs(1944) <= not b or a;
    layer1_outputs(1945) <= not (a and b);
    layer1_outputs(1946) <= b;
    layer1_outputs(1947) <= not a;
    layer1_outputs(1948) <= a xor b;
    layer1_outputs(1949) <= a;
    layer1_outputs(1950) <= not a;
    layer1_outputs(1951) <= a;
    layer1_outputs(1952) <= a;
    layer1_outputs(1953) <= a and not b;
    layer1_outputs(1954) <= not a;
    layer1_outputs(1955) <= not (a and b);
    layer1_outputs(1956) <= not (a and b);
    layer1_outputs(1957) <= not (a or b);
    layer1_outputs(1958) <= b;
    layer1_outputs(1959) <= not a;
    layer1_outputs(1960) <= a or b;
    layer1_outputs(1961) <= a or b;
    layer1_outputs(1962) <= not b or a;
    layer1_outputs(1963) <= a and b;
    layer1_outputs(1964) <= a and not b;
    layer1_outputs(1965) <= not b or a;
    layer1_outputs(1966) <= a xor b;
    layer1_outputs(1967) <= not (a or b);
    layer1_outputs(1968) <= not (a and b);
    layer1_outputs(1969) <= b and not a;
    layer1_outputs(1970) <= a and b;
    layer1_outputs(1971) <= a or b;
    layer1_outputs(1972) <= a xor b;
    layer1_outputs(1973) <= '0';
    layer1_outputs(1974) <= b;
    layer1_outputs(1975) <= not a;
    layer1_outputs(1976) <= not b or a;
    layer1_outputs(1977) <= a or b;
    layer1_outputs(1978) <= a or b;
    layer1_outputs(1979) <= a and b;
    layer1_outputs(1980) <= b;
    layer1_outputs(1981) <= not (a or b);
    layer1_outputs(1982) <= not (a xor b);
    layer1_outputs(1983) <= a and b;
    layer1_outputs(1984) <= a and b;
    layer1_outputs(1985) <= not (a or b);
    layer1_outputs(1986) <= a and b;
    layer1_outputs(1987) <= not (a or b);
    layer1_outputs(1988) <= not b;
    layer1_outputs(1989) <= b;
    layer1_outputs(1990) <= a or b;
    layer1_outputs(1991) <= a;
    layer1_outputs(1992) <= not b or a;
    layer1_outputs(1993) <= '0';
    layer1_outputs(1994) <= '1';
    layer1_outputs(1995) <= not a;
    layer1_outputs(1996) <= not b;
    layer1_outputs(1997) <= a and not b;
    layer1_outputs(1998) <= a and b;
    layer1_outputs(1999) <= a and b;
    layer1_outputs(2000) <= a and not b;
    layer1_outputs(2001) <= a and not b;
    layer1_outputs(2002) <= b;
    layer1_outputs(2003) <= not a or b;
    layer1_outputs(2004) <= a or b;
    layer1_outputs(2005) <= a;
    layer1_outputs(2006) <= not a;
    layer1_outputs(2007) <= not a;
    layer1_outputs(2008) <= '0';
    layer1_outputs(2009) <= '0';
    layer1_outputs(2010) <= not a or b;
    layer1_outputs(2011) <= a and not b;
    layer1_outputs(2012) <= '1';
    layer1_outputs(2013) <= a or b;
    layer1_outputs(2014) <= not b or a;
    layer1_outputs(2015) <= a and not b;
    layer1_outputs(2016) <= a xor b;
    layer1_outputs(2017) <= not (a and b);
    layer1_outputs(2018) <= a and b;
    layer1_outputs(2019) <= not (a xor b);
    layer1_outputs(2020) <= b and not a;
    layer1_outputs(2021) <= a and b;
    layer1_outputs(2022) <= not a or b;
    layer1_outputs(2023) <= not b or a;
    layer1_outputs(2024) <= not (a and b);
    layer1_outputs(2025) <= not (a or b);
    layer1_outputs(2026) <= not (a or b);
    layer1_outputs(2027) <= b and not a;
    layer1_outputs(2028) <= '0';
    layer1_outputs(2029) <= not b;
    layer1_outputs(2030) <= not a;
    layer1_outputs(2031) <= a or b;
    layer1_outputs(2032) <= a or b;
    layer1_outputs(2033) <= '0';
    layer1_outputs(2034) <= not a or b;
    layer1_outputs(2035) <= a and not b;
    layer1_outputs(2036) <= '0';
    layer1_outputs(2037) <= '0';
    layer1_outputs(2038) <= a and not b;
    layer1_outputs(2039) <= a;
    layer1_outputs(2040) <= '1';
    layer1_outputs(2041) <= '1';
    layer1_outputs(2042) <= not a or b;
    layer1_outputs(2043) <= b;
    layer1_outputs(2044) <= not (a or b);
    layer1_outputs(2045) <= not a;
    layer1_outputs(2046) <= not b or a;
    layer1_outputs(2047) <= '0';
    layer1_outputs(2048) <= a or b;
    layer1_outputs(2049) <= a or b;
    layer1_outputs(2050) <= '1';
    layer1_outputs(2051) <= a or b;
    layer1_outputs(2052) <= a and b;
    layer1_outputs(2053) <= not a;
    layer1_outputs(2054) <= b and not a;
    layer1_outputs(2055) <= not b or a;
    layer1_outputs(2056) <= not (a or b);
    layer1_outputs(2057) <= not a or b;
    layer1_outputs(2058) <= b and not a;
    layer1_outputs(2059) <= b;
    layer1_outputs(2060) <= '0';
    layer1_outputs(2061) <= not (a or b);
    layer1_outputs(2062) <= not (a or b);
    layer1_outputs(2063) <= not b or a;
    layer1_outputs(2064) <= '1';
    layer1_outputs(2065) <= a and b;
    layer1_outputs(2066) <= not b or a;
    layer1_outputs(2067) <= '0';
    layer1_outputs(2068) <= a or b;
    layer1_outputs(2069) <= a;
    layer1_outputs(2070) <= '0';
    layer1_outputs(2071) <= not (a or b);
    layer1_outputs(2072) <= '0';
    layer1_outputs(2073) <= '0';
    layer1_outputs(2074) <= a and b;
    layer1_outputs(2075) <= b;
    layer1_outputs(2076) <= not b;
    layer1_outputs(2077) <= a or b;
    layer1_outputs(2078) <= a and not b;
    layer1_outputs(2079) <= '1';
    layer1_outputs(2080) <= a;
    layer1_outputs(2081) <= '0';
    layer1_outputs(2082) <= a or b;
    layer1_outputs(2083) <= a or b;
    layer1_outputs(2084) <= not b;
    layer1_outputs(2085) <= a and not b;
    layer1_outputs(2086) <= b and not a;
    layer1_outputs(2087) <= a;
    layer1_outputs(2088) <= a and b;
    layer1_outputs(2089) <= not b or a;
    layer1_outputs(2090) <= not (a xor b);
    layer1_outputs(2091) <= not b or a;
    layer1_outputs(2092) <= a and not b;
    layer1_outputs(2093) <= a;
    layer1_outputs(2094) <= not b;
    layer1_outputs(2095) <= not b;
    layer1_outputs(2096) <= not b or a;
    layer1_outputs(2097) <= b;
    layer1_outputs(2098) <= not b;
    layer1_outputs(2099) <= a or b;
    layer1_outputs(2100) <= not (a and b);
    layer1_outputs(2101) <= a and b;
    layer1_outputs(2102) <= '0';
    layer1_outputs(2103) <= a or b;
    layer1_outputs(2104) <= not b;
    layer1_outputs(2105) <= a and not b;
    layer1_outputs(2106) <= b;
    layer1_outputs(2107) <= not b;
    layer1_outputs(2108) <= a and b;
    layer1_outputs(2109) <= a xor b;
    layer1_outputs(2110) <= b;
    layer1_outputs(2111) <= '1';
    layer1_outputs(2112) <= b;
    layer1_outputs(2113) <= not b;
    layer1_outputs(2114) <= not (a or b);
    layer1_outputs(2115) <= a or b;
    layer1_outputs(2116) <= not (a or b);
    layer1_outputs(2117) <= a and b;
    layer1_outputs(2118) <= not (a xor b);
    layer1_outputs(2119) <= a and not b;
    layer1_outputs(2120) <= a;
    layer1_outputs(2121) <= not a or b;
    layer1_outputs(2122) <= b;
    layer1_outputs(2123) <= '0';
    layer1_outputs(2124) <= not a or b;
    layer1_outputs(2125) <= '1';
    layer1_outputs(2126) <= not (a and b);
    layer1_outputs(2127) <= '1';
    layer1_outputs(2128) <= '0';
    layer1_outputs(2129) <= b;
    layer1_outputs(2130) <= a and b;
    layer1_outputs(2131) <= not (a xor b);
    layer1_outputs(2132) <= a and b;
    layer1_outputs(2133) <= not b;
    layer1_outputs(2134) <= a;
    layer1_outputs(2135) <= b;
    layer1_outputs(2136) <= '0';
    layer1_outputs(2137) <= '1';
    layer1_outputs(2138) <= a and not b;
    layer1_outputs(2139) <= not b;
    layer1_outputs(2140) <= not b or a;
    layer1_outputs(2141) <= not a or b;
    layer1_outputs(2142) <= not a or b;
    layer1_outputs(2143) <= not b or a;
    layer1_outputs(2144) <= '1';
    layer1_outputs(2145) <= '0';
    layer1_outputs(2146) <= b;
    layer1_outputs(2147) <= a xor b;
    layer1_outputs(2148) <= not b;
    layer1_outputs(2149) <= b and not a;
    layer1_outputs(2150) <= b;
    layer1_outputs(2151) <= not (a or b);
    layer1_outputs(2152) <= a and b;
    layer1_outputs(2153) <= not b;
    layer1_outputs(2154) <= not b;
    layer1_outputs(2155) <= not a;
    layer1_outputs(2156) <= a and b;
    layer1_outputs(2157) <= not (a xor b);
    layer1_outputs(2158) <= not (a xor b);
    layer1_outputs(2159) <= a or b;
    layer1_outputs(2160) <= b;
    layer1_outputs(2161) <= a and b;
    layer1_outputs(2162) <= b;
    layer1_outputs(2163) <= not b;
    layer1_outputs(2164) <= not (a xor b);
    layer1_outputs(2165) <= a and not b;
    layer1_outputs(2166) <= a;
    layer1_outputs(2167) <= '0';
    layer1_outputs(2168) <= not b;
    layer1_outputs(2169) <= a and b;
    layer1_outputs(2170) <= not (a and b);
    layer1_outputs(2171) <= '1';
    layer1_outputs(2172) <= '0';
    layer1_outputs(2173) <= b and not a;
    layer1_outputs(2174) <= '0';
    layer1_outputs(2175) <= '0';
    layer1_outputs(2176) <= not (a or b);
    layer1_outputs(2177) <= not (a or b);
    layer1_outputs(2178) <= a and not b;
    layer1_outputs(2179) <= not a or b;
    layer1_outputs(2180) <= not (a and b);
    layer1_outputs(2181) <= not (a or b);
    layer1_outputs(2182) <= not (a or b);
    layer1_outputs(2183) <= not (a or b);
    layer1_outputs(2184) <= not (a or b);
    layer1_outputs(2185) <= b;
    layer1_outputs(2186) <= not (a and b);
    layer1_outputs(2187) <= not b;
    layer1_outputs(2188) <= b;
    layer1_outputs(2189) <= a xor b;
    layer1_outputs(2190) <= not a or b;
    layer1_outputs(2191) <= not a;
    layer1_outputs(2192) <= not (a and b);
    layer1_outputs(2193) <= not a or b;
    layer1_outputs(2194) <= a;
    layer1_outputs(2195) <= not a;
    layer1_outputs(2196) <= not (a and b);
    layer1_outputs(2197) <= b and not a;
    layer1_outputs(2198) <= a and b;
    layer1_outputs(2199) <= a and b;
    layer1_outputs(2200) <= not b or a;
    layer1_outputs(2201) <= a;
    layer1_outputs(2202) <= a or b;
    layer1_outputs(2203) <= a;
    layer1_outputs(2204) <= a or b;
    layer1_outputs(2205) <= not (a or b);
    layer1_outputs(2206) <= a or b;
    layer1_outputs(2207) <= not a or b;
    layer1_outputs(2208) <= not a;
    layer1_outputs(2209) <= '0';
    layer1_outputs(2210) <= b;
    layer1_outputs(2211) <= '1';
    layer1_outputs(2212) <= a;
    layer1_outputs(2213) <= not b or a;
    layer1_outputs(2214) <= a and not b;
    layer1_outputs(2215) <= '1';
    layer1_outputs(2216) <= a or b;
    layer1_outputs(2217) <= not b;
    layer1_outputs(2218) <= not a or b;
    layer1_outputs(2219) <= '1';
    layer1_outputs(2220) <= '1';
    layer1_outputs(2221) <= a;
    layer1_outputs(2222) <= not b or a;
    layer1_outputs(2223) <= not a or b;
    layer1_outputs(2224) <= not a or b;
    layer1_outputs(2225) <= '0';
    layer1_outputs(2226) <= not (a and b);
    layer1_outputs(2227) <= a xor b;
    layer1_outputs(2228) <= b;
    layer1_outputs(2229) <= '0';
    layer1_outputs(2230) <= b and not a;
    layer1_outputs(2231) <= b and not a;
    layer1_outputs(2232) <= '0';
    layer1_outputs(2233) <= b and not a;
    layer1_outputs(2234) <= a;
    layer1_outputs(2235) <= not a;
    layer1_outputs(2236) <= a;
    layer1_outputs(2237) <= not (a xor b);
    layer1_outputs(2238) <= b;
    layer1_outputs(2239) <= not b;
    layer1_outputs(2240) <= b and not a;
    layer1_outputs(2241) <= not a or b;
    layer1_outputs(2242) <= a or b;
    layer1_outputs(2243) <= a;
    layer1_outputs(2244) <= a and b;
    layer1_outputs(2245) <= a or b;
    layer1_outputs(2246) <= b and not a;
    layer1_outputs(2247) <= a and b;
    layer1_outputs(2248) <= a or b;
    layer1_outputs(2249) <= a and b;
    layer1_outputs(2250) <= a and b;
    layer1_outputs(2251) <= not (a xor b);
    layer1_outputs(2252) <= '0';
    layer1_outputs(2253) <= not a;
    layer1_outputs(2254) <= a xor b;
    layer1_outputs(2255) <= not a or b;
    layer1_outputs(2256) <= a and b;
    layer1_outputs(2257) <= b;
    layer1_outputs(2258) <= a;
    layer1_outputs(2259) <= not (a and b);
    layer1_outputs(2260) <= not b or a;
    layer1_outputs(2261) <= not a;
    layer1_outputs(2262) <= a;
    layer1_outputs(2263) <= not b;
    layer1_outputs(2264) <= a and not b;
    layer1_outputs(2265) <= b and not a;
    layer1_outputs(2266) <= not (a or b);
    layer1_outputs(2267) <= not b or a;
    layer1_outputs(2268) <= not b;
    layer1_outputs(2269) <= not (a xor b);
    layer1_outputs(2270) <= a and b;
    layer1_outputs(2271) <= not a;
    layer1_outputs(2272) <= not a or b;
    layer1_outputs(2273) <= a and b;
    layer1_outputs(2274) <= not a or b;
    layer1_outputs(2275) <= a or b;
    layer1_outputs(2276) <= not (a or b);
    layer1_outputs(2277) <= a;
    layer1_outputs(2278) <= a or b;
    layer1_outputs(2279) <= a and b;
    layer1_outputs(2280) <= a and not b;
    layer1_outputs(2281) <= not a or b;
    layer1_outputs(2282) <= not a;
    layer1_outputs(2283) <= not a;
    layer1_outputs(2284) <= b;
    layer1_outputs(2285) <= a and b;
    layer1_outputs(2286) <= not b;
    layer1_outputs(2287) <= b and not a;
    layer1_outputs(2288) <= a;
    layer1_outputs(2289) <= not a;
    layer1_outputs(2290) <= '0';
    layer1_outputs(2291) <= not (a and b);
    layer1_outputs(2292) <= not a;
    layer1_outputs(2293) <= b;
    layer1_outputs(2294) <= not (a or b);
    layer1_outputs(2295) <= a and not b;
    layer1_outputs(2296) <= not (a or b);
    layer1_outputs(2297) <= not a;
    layer1_outputs(2298) <= not a or b;
    layer1_outputs(2299) <= a;
    layer1_outputs(2300) <= a;
    layer1_outputs(2301) <= '0';
    layer1_outputs(2302) <= not a;
    layer1_outputs(2303) <= not b;
    layer1_outputs(2304) <= a or b;
    layer1_outputs(2305) <= not b;
    layer1_outputs(2306) <= '1';
    layer1_outputs(2307) <= not (a xor b);
    layer1_outputs(2308) <= '1';
    layer1_outputs(2309) <= not b;
    layer1_outputs(2310) <= not b;
    layer1_outputs(2311) <= b;
    layer1_outputs(2312) <= not b;
    layer1_outputs(2313) <= not (a and b);
    layer1_outputs(2314) <= a xor b;
    layer1_outputs(2315) <= '0';
    layer1_outputs(2316) <= a and not b;
    layer1_outputs(2317) <= a or b;
    layer1_outputs(2318) <= '0';
    layer1_outputs(2319) <= a;
    layer1_outputs(2320) <= b and not a;
    layer1_outputs(2321) <= b and not a;
    layer1_outputs(2322) <= not b;
    layer1_outputs(2323) <= a and not b;
    layer1_outputs(2324) <= a or b;
    layer1_outputs(2325) <= not (a or b);
    layer1_outputs(2326) <= b;
    layer1_outputs(2327) <= not b;
    layer1_outputs(2328) <= a and b;
    layer1_outputs(2329) <= '1';
    layer1_outputs(2330) <= not a or b;
    layer1_outputs(2331) <= not a or b;
    layer1_outputs(2332) <= '0';
    layer1_outputs(2333) <= not b;
    layer1_outputs(2334) <= a and not b;
    layer1_outputs(2335) <= not (a and b);
    layer1_outputs(2336) <= not (a and b);
    layer1_outputs(2337) <= not (a xor b);
    layer1_outputs(2338) <= not (a xor b);
    layer1_outputs(2339) <= b and not a;
    layer1_outputs(2340) <= not a or b;
    layer1_outputs(2341) <= not (a xor b);
    layer1_outputs(2342) <= a;
    layer1_outputs(2343) <= not b;
    layer1_outputs(2344) <= a;
    layer1_outputs(2345) <= not b;
    layer1_outputs(2346) <= a;
    layer1_outputs(2347) <= a or b;
    layer1_outputs(2348) <= a or b;
    layer1_outputs(2349) <= not (a or b);
    layer1_outputs(2350) <= '1';
    layer1_outputs(2351) <= a and not b;
    layer1_outputs(2352) <= not b;
    layer1_outputs(2353) <= '0';
    layer1_outputs(2354) <= not (a or b);
    layer1_outputs(2355) <= not b;
    layer1_outputs(2356) <= a and not b;
    layer1_outputs(2357) <= not (a and b);
    layer1_outputs(2358) <= b;
    layer1_outputs(2359) <= b;
    layer1_outputs(2360) <= '1';
    layer1_outputs(2361) <= a xor b;
    layer1_outputs(2362) <= a and b;
    layer1_outputs(2363) <= not (a or b);
    layer1_outputs(2364) <= '0';
    layer1_outputs(2365) <= b and not a;
    layer1_outputs(2366) <= not (a xor b);
    layer1_outputs(2367) <= not (a and b);
    layer1_outputs(2368) <= '0';
    layer1_outputs(2369) <= not b or a;
    layer1_outputs(2370) <= '1';
    layer1_outputs(2371) <= b;
    layer1_outputs(2372) <= not a or b;
    layer1_outputs(2373) <= b;
    layer1_outputs(2374) <= '0';
    layer1_outputs(2375) <= b and not a;
    layer1_outputs(2376) <= not b or a;
    layer1_outputs(2377) <= a or b;
    layer1_outputs(2378) <= '0';
    layer1_outputs(2379) <= not a or b;
    layer1_outputs(2380) <= not b;
    layer1_outputs(2381) <= '0';
    layer1_outputs(2382) <= a;
    layer1_outputs(2383) <= a and b;
    layer1_outputs(2384) <= not a;
    layer1_outputs(2385) <= not b or a;
    layer1_outputs(2386) <= not a or b;
    layer1_outputs(2387) <= not b or a;
    layer1_outputs(2388) <= not a;
    layer1_outputs(2389) <= b;
    layer1_outputs(2390) <= a or b;
    layer1_outputs(2391) <= not a or b;
    layer1_outputs(2392) <= a;
    layer1_outputs(2393) <= '1';
    layer1_outputs(2394) <= not (a and b);
    layer1_outputs(2395) <= not (a or b);
    layer1_outputs(2396) <= b;
    layer1_outputs(2397) <= not a or b;
    layer1_outputs(2398) <= a and b;
    layer1_outputs(2399) <= b;
    layer1_outputs(2400) <= not a;
    layer1_outputs(2401) <= not (a and b);
    layer1_outputs(2402) <= not a;
    layer1_outputs(2403) <= not b;
    layer1_outputs(2404) <= not (a and b);
    layer1_outputs(2405) <= not b or a;
    layer1_outputs(2406) <= not (a and b);
    layer1_outputs(2407) <= b;
    layer1_outputs(2408) <= b and not a;
    layer1_outputs(2409) <= '1';
    layer1_outputs(2410) <= a;
    layer1_outputs(2411) <= not b;
    layer1_outputs(2412) <= not b;
    layer1_outputs(2413) <= not a;
    layer1_outputs(2414) <= a or b;
    layer1_outputs(2415) <= not a;
    layer1_outputs(2416) <= not a or b;
    layer1_outputs(2417) <= '0';
    layer1_outputs(2418) <= a and b;
    layer1_outputs(2419) <= not (a and b);
    layer1_outputs(2420) <= not a;
    layer1_outputs(2421) <= not (a and b);
    layer1_outputs(2422) <= '1';
    layer1_outputs(2423) <= not b or a;
    layer1_outputs(2424) <= not b;
    layer1_outputs(2425) <= not b;
    layer1_outputs(2426) <= not b or a;
    layer1_outputs(2427) <= not (a and b);
    layer1_outputs(2428) <= '1';
    layer1_outputs(2429) <= not a;
    layer1_outputs(2430) <= not b;
    layer1_outputs(2431) <= not (a xor b);
    layer1_outputs(2432) <= a and not b;
    layer1_outputs(2433) <= a or b;
    layer1_outputs(2434) <= b and not a;
    layer1_outputs(2435) <= not a;
    layer1_outputs(2436) <= b and not a;
    layer1_outputs(2437) <= b and not a;
    layer1_outputs(2438) <= not (a and b);
    layer1_outputs(2439) <= not (a and b);
    layer1_outputs(2440) <= a and not b;
    layer1_outputs(2441) <= not b;
    layer1_outputs(2442) <= not a;
    layer1_outputs(2443) <= not (a and b);
    layer1_outputs(2444) <= '1';
    layer1_outputs(2445) <= a and not b;
    layer1_outputs(2446) <= not (a or b);
    layer1_outputs(2447) <= a;
    layer1_outputs(2448) <= b;
    layer1_outputs(2449) <= b;
    layer1_outputs(2450) <= a and b;
    layer1_outputs(2451) <= b;
    layer1_outputs(2452) <= not (a or b);
    layer1_outputs(2453) <= a xor b;
    layer1_outputs(2454) <= not a;
    layer1_outputs(2455) <= not a or b;
    layer1_outputs(2456) <= '0';
    layer1_outputs(2457) <= not a;
    layer1_outputs(2458) <= not b or a;
    layer1_outputs(2459) <= b and not a;
    layer1_outputs(2460) <= not (a or b);
    layer1_outputs(2461) <= '0';
    layer1_outputs(2462) <= a and not b;
    layer1_outputs(2463) <= not (a and b);
    layer1_outputs(2464) <= a and b;
    layer1_outputs(2465) <= not a or b;
    layer1_outputs(2466) <= not a or b;
    layer1_outputs(2467) <= a and b;
    layer1_outputs(2468) <= not b;
    layer1_outputs(2469) <= a and not b;
    layer1_outputs(2470) <= not (a and b);
    layer1_outputs(2471) <= not (a or b);
    layer1_outputs(2472) <= not (a and b);
    layer1_outputs(2473) <= a;
    layer1_outputs(2474) <= not a;
    layer1_outputs(2475) <= a and not b;
    layer1_outputs(2476) <= not b;
    layer1_outputs(2477) <= a;
    layer1_outputs(2478) <= '0';
    layer1_outputs(2479) <= a or b;
    layer1_outputs(2480) <= a or b;
    layer1_outputs(2481) <= a and b;
    layer1_outputs(2482) <= b;
    layer1_outputs(2483) <= a;
    layer1_outputs(2484) <= not b or a;
    layer1_outputs(2485) <= a xor b;
    layer1_outputs(2486) <= b and not a;
    layer1_outputs(2487) <= not a or b;
    layer1_outputs(2488) <= not (a or b);
    layer1_outputs(2489) <= a and b;
    layer1_outputs(2490) <= not b or a;
    layer1_outputs(2491) <= not (a or b);
    layer1_outputs(2492) <= b;
    layer1_outputs(2493) <= not a;
    layer1_outputs(2494) <= not b or a;
    layer1_outputs(2495) <= b and not a;
    layer1_outputs(2496) <= not (a xor b);
    layer1_outputs(2497) <= a or b;
    layer1_outputs(2498) <= not a or b;
    layer1_outputs(2499) <= not b;
    layer1_outputs(2500) <= not (a and b);
    layer1_outputs(2501) <= a and not b;
    layer1_outputs(2502) <= b and not a;
    layer1_outputs(2503) <= not (a xor b);
    layer1_outputs(2504) <= not (a or b);
    layer1_outputs(2505) <= not (a or b);
    layer1_outputs(2506) <= a and not b;
    layer1_outputs(2507) <= a and b;
    layer1_outputs(2508) <= a;
    layer1_outputs(2509) <= b and not a;
    layer1_outputs(2510) <= not (a and b);
    layer1_outputs(2511) <= a and not b;
    layer1_outputs(2512) <= not b;
    layer1_outputs(2513) <= not a or b;
    layer1_outputs(2514) <= '0';
    layer1_outputs(2515) <= '1';
    layer1_outputs(2516) <= not a or b;
    layer1_outputs(2517) <= a;
    layer1_outputs(2518) <= a and b;
    layer1_outputs(2519) <= a and not b;
    layer1_outputs(2520) <= b;
    layer1_outputs(2521) <= a;
    layer1_outputs(2522) <= not a;
    layer1_outputs(2523) <= '0';
    layer1_outputs(2524) <= not (a and b);
    layer1_outputs(2525) <= not b or a;
    layer1_outputs(2526) <= not (a or b);
    layer1_outputs(2527) <= '0';
    layer1_outputs(2528) <= not (a or b);
    layer1_outputs(2529) <= not a;
    layer1_outputs(2530) <= a xor b;
    layer1_outputs(2531) <= a;
    layer1_outputs(2532) <= b;
    layer1_outputs(2533) <= not a or b;
    layer1_outputs(2534) <= '0';
    layer1_outputs(2535) <= '0';
    layer1_outputs(2536) <= not (a or b);
    layer1_outputs(2537) <= not b or a;
    layer1_outputs(2538) <= a xor b;
    layer1_outputs(2539) <= a and not b;
    layer1_outputs(2540) <= '0';
    layer1_outputs(2541) <= a;
    layer1_outputs(2542) <= not a;
    layer1_outputs(2543) <= not b or a;
    layer1_outputs(2544) <= not (a or b);
    layer1_outputs(2545) <= not b or a;
    layer1_outputs(2546) <= not a or b;
    layer1_outputs(2547) <= a and b;
    layer1_outputs(2548) <= b and not a;
    layer1_outputs(2549) <= a and not b;
    layer1_outputs(2550) <= a;
    layer1_outputs(2551) <= b and not a;
    layer1_outputs(2552) <= not a;
    layer1_outputs(2553) <= not a or b;
    layer1_outputs(2554) <= a and b;
    layer1_outputs(2555) <= a;
    layer1_outputs(2556) <= not a or b;
    layer1_outputs(2557) <= b and not a;
    layer1_outputs(2558) <= not b or a;
    layer1_outputs(2559) <= a and not b;
    layer1_outputs(2560) <= a or b;
    layer1_outputs(2561) <= not (a or b);
    layer1_outputs(2562) <= not (a xor b);
    layer1_outputs(2563) <= '0';
    layer1_outputs(2564) <= a and not b;
    layer1_outputs(2565) <= '1';
    layer1_outputs(2566) <= b and not a;
    layer1_outputs(2567) <= not a or b;
    layer1_outputs(2568) <= not (a and b);
    layer1_outputs(2569) <= not b or a;
    layer1_outputs(2570) <= not a or b;
    layer1_outputs(2571) <= not a;
    layer1_outputs(2572) <= not b;
    layer1_outputs(2573) <= a;
    layer1_outputs(2574) <= not a or b;
    layer1_outputs(2575) <= not a;
    layer1_outputs(2576) <= not a;
    layer1_outputs(2577) <= a and b;
    layer1_outputs(2578) <= a and b;
    layer1_outputs(2579) <= not b or a;
    layer1_outputs(2580) <= a xor b;
    layer1_outputs(2581) <= b and not a;
    layer1_outputs(2582) <= a and b;
    layer1_outputs(2583) <= not b;
    layer1_outputs(2584) <= not (a and b);
    layer1_outputs(2585) <= not a or b;
    layer1_outputs(2586) <= a;
    layer1_outputs(2587) <= not (a or b);
    layer1_outputs(2588) <= b;
    layer1_outputs(2589) <= b;
    layer1_outputs(2590) <= '0';
    layer1_outputs(2591) <= '0';
    layer1_outputs(2592) <= not b;
    layer1_outputs(2593) <= a or b;
    layer1_outputs(2594) <= not (a and b);
    layer1_outputs(2595) <= not (a or b);
    layer1_outputs(2596) <= not a or b;
    layer1_outputs(2597) <= not (a xor b);
    layer1_outputs(2598) <= a and b;
    layer1_outputs(2599) <= '1';
    layer1_outputs(2600) <= a and b;
    layer1_outputs(2601) <= a or b;
    layer1_outputs(2602) <= '0';
    layer1_outputs(2603) <= a;
    layer1_outputs(2604) <= not b;
    layer1_outputs(2605) <= not a or b;
    layer1_outputs(2606) <= a or b;
    layer1_outputs(2607) <= b and not a;
    layer1_outputs(2608) <= not a or b;
    layer1_outputs(2609) <= '0';
    layer1_outputs(2610) <= '1';
    layer1_outputs(2611) <= a or b;
    layer1_outputs(2612) <= '0';
    layer1_outputs(2613) <= b and not a;
    layer1_outputs(2614) <= a and b;
    layer1_outputs(2615) <= b and not a;
    layer1_outputs(2616) <= not a;
    layer1_outputs(2617) <= not (a and b);
    layer1_outputs(2618) <= a;
    layer1_outputs(2619) <= '1';
    layer1_outputs(2620) <= not b or a;
    layer1_outputs(2621) <= not (a and b);
    layer1_outputs(2622) <= not (a or b);
    layer1_outputs(2623) <= a or b;
    layer1_outputs(2624) <= a xor b;
    layer1_outputs(2625) <= a;
    layer1_outputs(2626) <= not b or a;
    layer1_outputs(2627) <= b;
    layer1_outputs(2628) <= not a;
    layer1_outputs(2629) <= a and b;
    layer1_outputs(2630) <= not a or b;
    layer1_outputs(2631) <= b and not a;
    layer1_outputs(2632) <= b;
    layer1_outputs(2633) <= not (a and b);
    layer1_outputs(2634) <= not b;
    layer1_outputs(2635) <= not (a or b);
    layer1_outputs(2636) <= '0';
    layer1_outputs(2637) <= not b;
    layer1_outputs(2638) <= '1';
    layer1_outputs(2639) <= not (a or b);
    layer1_outputs(2640) <= a and b;
    layer1_outputs(2641) <= a and not b;
    layer1_outputs(2642) <= a;
    layer1_outputs(2643) <= '1';
    layer1_outputs(2644) <= b and not a;
    layer1_outputs(2645) <= not a or b;
    layer1_outputs(2646) <= '0';
    layer1_outputs(2647) <= a and not b;
    layer1_outputs(2648) <= a and b;
    layer1_outputs(2649) <= b and not a;
    layer1_outputs(2650) <= a xor b;
    layer1_outputs(2651) <= a and not b;
    layer1_outputs(2652) <= b and not a;
    layer1_outputs(2653) <= '1';
    layer1_outputs(2654) <= a xor b;
    layer1_outputs(2655) <= not (a or b);
    layer1_outputs(2656) <= not (a and b);
    layer1_outputs(2657) <= a and not b;
    layer1_outputs(2658) <= not (a and b);
    layer1_outputs(2659) <= not (a or b);
    layer1_outputs(2660) <= a and b;
    layer1_outputs(2661) <= a and not b;
    layer1_outputs(2662) <= not a or b;
    layer1_outputs(2663) <= not a;
    layer1_outputs(2664) <= a or b;
    layer1_outputs(2665) <= not (a xor b);
    layer1_outputs(2666) <= a and b;
    layer1_outputs(2667) <= not b or a;
    layer1_outputs(2668) <= not b or a;
    layer1_outputs(2669) <= not b;
    layer1_outputs(2670) <= not b or a;
    layer1_outputs(2671) <= not a;
    layer1_outputs(2672) <= a;
    layer1_outputs(2673) <= b;
    layer1_outputs(2674) <= not a or b;
    layer1_outputs(2675) <= '0';
    layer1_outputs(2676) <= '0';
    layer1_outputs(2677) <= b;
    layer1_outputs(2678) <= b;
    layer1_outputs(2679) <= not a or b;
    layer1_outputs(2680) <= a xor b;
    layer1_outputs(2681) <= a and b;
    layer1_outputs(2682) <= a or b;
    layer1_outputs(2683) <= not a or b;
    layer1_outputs(2684) <= not a;
    layer1_outputs(2685) <= b and not a;
    layer1_outputs(2686) <= a;
    layer1_outputs(2687) <= '1';
    layer1_outputs(2688) <= not a;
    layer1_outputs(2689) <= not b;
    layer1_outputs(2690) <= not b or a;
    layer1_outputs(2691) <= a and b;
    layer1_outputs(2692) <= not (a xor b);
    layer1_outputs(2693) <= a and b;
    layer1_outputs(2694) <= not a or b;
    layer1_outputs(2695) <= b;
    layer1_outputs(2696) <= b;
    layer1_outputs(2697) <= a;
    layer1_outputs(2698) <= a xor b;
    layer1_outputs(2699) <= not (a or b);
    layer1_outputs(2700) <= a or b;
    layer1_outputs(2701) <= a;
    layer1_outputs(2702) <= not (a or b);
    layer1_outputs(2703) <= not (a or b);
    layer1_outputs(2704) <= not b;
    layer1_outputs(2705) <= '0';
    layer1_outputs(2706) <= not a or b;
    layer1_outputs(2707) <= not a or b;
    layer1_outputs(2708) <= a;
    layer1_outputs(2709) <= not a or b;
    layer1_outputs(2710) <= b;
    layer1_outputs(2711) <= not b or a;
    layer1_outputs(2712) <= a or b;
    layer1_outputs(2713) <= not b or a;
    layer1_outputs(2714) <= not a or b;
    layer1_outputs(2715) <= b;
    layer1_outputs(2716) <= not (a xor b);
    layer1_outputs(2717) <= a;
    layer1_outputs(2718) <= not (a and b);
    layer1_outputs(2719) <= not a;
    layer1_outputs(2720) <= not b or a;
    layer1_outputs(2721) <= a;
    layer1_outputs(2722) <= b and not a;
    layer1_outputs(2723) <= b;
    layer1_outputs(2724) <= a and not b;
    layer1_outputs(2725) <= b and not a;
    layer1_outputs(2726) <= a xor b;
    layer1_outputs(2727) <= a;
    layer1_outputs(2728) <= a or b;
    layer1_outputs(2729) <= a xor b;
    layer1_outputs(2730) <= '1';
    layer1_outputs(2731) <= '1';
    layer1_outputs(2732) <= a xor b;
    layer1_outputs(2733) <= not a or b;
    layer1_outputs(2734) <= not (a and b);
    layer1_outputs(2735) <= not b or a;
    layer1_outputs(2736) <= not b or a;
    layer1_outputs(2737) <= '1';
    layer1_outputs(2738) <= a or b;
    layer1_outputs(2739) <= not b or a;
    layer1_outputs(2740) <= not a;
    layer1_outputs(2741) <= '0';
    layer1_outputs(2742) <= not b;
    layer1_outputs(2743) <= not a;
    layer1_outputs(2744) <= b and not a;
    layer1_outputs(2745) <= not (a and b);
    layer1_outputs(2746) <= b;
    layer1_outputs(2747) <= not b or a;
    layer1_outputs(2748) <= a and b;
    layer1_outputs(2749) <= '0';
    layer1_outputs(2750) <= not a;
    layer1_outputs(2751) <= b and not a;
    layer1_outputs(2752) <= '1';
    layer1_outputs(2753) <= not a or b;
    layer1_outputs(2754) <= not (a or b);
    layer1_outputs(2755) <= not b;
    layer1_outputs(2756) <= b;
    layer1_outputs(2757) <= a and not b;
    layer1_outputs(2758) <= '0';
    layer1_outputs(2759) <= a and b;
    layer1_outputs(2760) <= b;
    layer1_outputs(2761) <= a xor b;
    layer1_outputs(2762) <= a;
    layer1_outputs(2763) <= a;
    layer1_outputs(2764) <= not a;
    layer1_outputs(2765) <= a and b;
    layer1_outputs(2766) <= a and b;
    layer1_outputs(2767) <= not a;
    layer1_outputs(2768) <= a or b;
    layer1_outputs(2769) <= a and b;
    layer1_outputs(2770) <= a xor b;
    layer1_outputs(2771) <= b;
    layer1_outputs(2772) <= not a;
    layer1_outputs(2773) <= '0';
    layer1_outputs(2774) <= a or b;
    layer1_outputs(2775) <= not b;
    layer1_outputs(2776) <= a or b;
    layer1_outputs(2777) <= a and b;
    layer1_outputs(2778) <= a xor b;
    layer1_outputs(2779) <= not b or a;
    layer1_outputs(2780) <= a xor b;
    layer1_outputs(2781) <= '0';
    layer1_outputs(2782) <= not a;
    layer1_outputs(2783) <= not b;
    layer1_outputs(2784) <= a or b;
    layer1_outputs(2785) <= a;
    layer1_outputs(2786) <= b and not a;
    layer1_outputs(2787) <= not a or b;
    layer1_outputs(2788) <= a xor b;
    layer1_outputs(2789) <= a xor b;
    layer1_outputs(2790) <= a;
    layer1_outputs(2791) <= a;
    layer1_outputs(2792) <= not a;
    layer1_outputs(2793) <= not (a and b);
    layer1_outputs(2794) <= b;
    layer1_outputs(2795) <= not (a and b);
    layer1_outputs(2796) <= a;
    layer1_outputs(2797) <= not b;
    layer1_outputs(2798) <= not (a and b);
    layer1_outputs(2799) <= not (a or b);
    layer1_outputs(2800) <= '0';
    layer1_outputs(2801) <= b;
    layer1_outputs(2802) <= a or b;
    layer1_outputs(2803) <= not a or b;
    layer1_outputs(2804) <= not a or b;
    layer1_outputs(2805) <= a or b;
    layer1_outputs(2806) <= not (a or b);
    layer1_outputs(2807) <= a or b;
    layer1_outputs(2808) <= a and b;
    layer1_outputs(2809) <= b;
    layer1_outputs(2810) <= a or b;
    layer1_outputs(2811) <= a and b;
    layer1_outputs(2812) <= b;
    layer1_outputs(2813) <= '1';
    layer1_outputs(2814) <= a;
    layer1_outputs(2815) <= a;
    layer1_outputs(2816) <= a;
    layer1_outputs(2817) <= '0';
    layer1_outputs(2818) <= not b or a;
    layer1_outputs(2819) <= a;
    layer1_outputs(2820) <= b and not a;
    layer1_outputs(2821) <= not b or a;
    layer1_outputs(2822) <= a and not b;
    layer1_outputs(2823) <= not (a and b);
    layer1_outputs(2824) <= not a or b;
    layer1_outputs(2825) <= not a or b;
    layer1_outputs(2826) <= b and not a;
    layer1_outputs(2827) <= '1';
    layer1_outputs(2828) <= a or b;
    layer1_outputs(2829) <= a and b;
    layer1_outputs(2830) <= '1';
    layer1_outputs(2831) <= a and not b;
    layer1_outputs(2832) <= a and b;
    layer1_outputs(2833) <= not a or b;
    layer1_outputs(2834) <= a or b;
    layer1_outputs(2835) <= a xor b;
    layer1_outputs(2836) <= a;
    layer1_outputs(2837) <= not (a or b);
    layer1_outputs(2838) <= a and b;
    layer1_outputs(2839) <= not a;
    layer1_outputs(2840) <= not b or a;
    layer1_outputs(2841) <= not b or a;
    layer1_outputs(2842) <= not (a xor b);
    layer1_outputs(2843) <= not a or b;
    layer1_outputs(2844) <= a xor b;
    layer1_outputs(2845) <= not (a xor b);
    layer1_outputs(2846) <= '1';
    layer1_outputs(2847) <= b and not a;
    layer1_outputs(2848) <= a and b;
    layer1_outputs(2849) <= a and not b;
    layer1_outputs(2850) <= '1';
    layer1_outputs(2851) <= not (a or b);
    layer1_outputs(2852) <= not b;
    layer1_outputs(2853) <= not a;
    layer1_outputs(2854) <= not b or a;
    layer1_outputs(2855) <= not b;
    layer1_outputs(2856) <= not (a and b);
    layer1_outputs(2857) <= a;
    layer1_outputs(2858) <= a or b;
    layer1_outputs(2859) <= a or b;
    layer1_outputs(2860) <= not a or b;
    layer1_outputs(2861) <= not a;
    layer1_outputs(2862) <= '1';
    layer1_outputs(2863) <= not b or a;
    layer1_outputs(2864) <= b;
    layer1_outputs(2865) <= not a;
    layer1_outputs(2866) <= a;
    layer1_outputs(2867) <= a or b;
    layer1_outputs(2868) <= not (a and b);
    layer1_outputs(2869) <= not (a and b);
    layer1_outputs(2870) <= a xor b;
    layer1_outputs(2871) <= a and not b;
    layer1_outputs(2872) <= not a;
    layer1_outputs(2873) <= b;
    layer1_outputs(2874) <= '0';
    layer1_outputs(2875) <= not (a or b);
    layer1_outputs(2876) <= a;
    layer1_outputs(2877) <= not (a or b);
    layer1_outputs(2878) <= not a or b;
    layer1_outputs(2879) <= b and not a;
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= a or b;
    layer1_outputs(2882) <= not a;
    layer1_outputs(2883) <= not b;
    layer1_outputs(2884) <= '0';
    layer1_outputs(2885) <= a and not b;
    layer1_outputs(2886) <= not (a or b);
    layer1_outputs(2887) <= a or b;
    layer1_outputs(2888) <= not a;
    layer1_outputs(2889) <= b;
    layer1_outputs(2890) <= '0';
    layer1_outputs(2891) <= not (a or b);
    layer1_outputs(2892) <= not b;
    layer1_outputs(2893) <= '1';
    layer1_outputs(2894) <= b;
    layer1_outputs(2895) <= a and not b;
    layer1_outputs(2896) <= not (a or b);
    layer1_outputs(2897) <= not (a xor b);
    layer1_outputs(2898) <= '0';
    layer1_outputs(2899) <= a xor b;
    layer1_outputs(2900) <= not b;
    layer1_outputs(2901) <= a or b;
    layer1_outputs(2902) <= a;
    layer1_outputs(2903) <= b and not a;
    layer1_outputs(2904) <= b;
    layer1_outputs(2905) <= b and not a;
    layer1_outputs(2906) <= a;
    layer1_outputs(2907) <= not b;
    layer1_outputs(2908) <= not a or b;
    layer1_outputs(2909) <= not b or a;
    layer1_outputs(2910) <= b and not a;
    layer1_outputs(2911) <= b and not a;
    layer1_outputs(2912) <= a and not b;
    layer1_outputs(2913) <= a and b;
    layer1_outputs(2914) <= not b or a;
    layer1_outputs(2915) <= '1';
    layer1_outputs(2916) <= b and not a;
    layer1_outputs(2917) <= a and not b;
    layer1_outputs(2918) <= '1';
    layer1_outputs(2919) <= a;
    layer1_outputs(2920) <= a and b;
    layer1_outputs(2921) <= not (a or b);
    layer1_outputs(2922) <= a or b;
    layer1_outputs(2923) <= a;
    layer1_outputs(2924) <= not (a or b);
    layer1_outputs(2925) <= a;
    layer1_outputs(2926) <= not b;
    layer1_outputs(2927) <= not (a or b);
    layer1_outputs(2928) <= a and b;
    layer1_outputs(2929) <= b and not a;
    layer1_outputs(2930) <= b;
    layer1_outputs(2931) <= not b;
    layer1_outputs(2932) <= a and not b;
    layer1_outputs(2933) <= a and not b;
    layer1_outputs(2934) <= not (a xor b);
    layer1_outputs(2935) <= '0';
    layer1_outputs(2936) <= not a;
    layer1_outputs(2937) <= not a;
    layer1_outputs(2938) <= '1';
    layer1_outputs(2939) <= b and not a;
    layer1_outputs(2940) <= b;
    layer1_outputs(2941) <= not a;
    layer1_outputs(2942) <= b and not a;
    layer1_outputs(2943) <= a;
    layer1_outputs(2944) <= a and b;
    layer1_outputs(2945) <= not a or b;
    layer1_outputs(2946) <= b and not a;
    layer1_outputs(2947) <= a;
    layer1_outputs(2948) <= a;
    layer1_outputs(2949) <= not (a and b);
    layer1_outputs(2950) <= not a or b;
    layer1_outputs(2951) <= b;
    layer1_outputs(2952) <= b;
    layer1_outputs(2953) <= a and b;
    layer1_outputs(2954) <= not (a or b);
    layer1_outputs(2955) <= a and b;
    layer1_outputs(2956) <= b;
    layer1_outputs(2957) <= not b;
    layer1_outputs(2958) <= not a;
    layer1_outputs(2959) <= not b;
    layer1_outputs(2960) <= b;
    layer1_outputs(2961) <= not (a xor b);
    layer1_outputs(2962) <= a;
    layer1_outputs(2963) <= a xor b;
    layer1_outputs(2964) <= not (a and b);
    layer1_outputs(2965) <= not b or a;
    layer1_outputs(2966) <= b;
    layer1_outputs(2967) <= not (a or b);
    layer1_outputs(2968) <= not b or a;
    layer1_outputs(2969) <= a or b;
    layer1_outputs(2970) <= not a or b;
    layer1_outputs(2971) <= not a;
    layer1_outputs(2972) <= not (a and b);
    layer1_outputs(2973) <= '0';
    layer1_outputs(2974) <= a and b;
    layer1_outputs(2975) <= '0';
    layer1_outputs(2976) <= not (a or b);
    layer1_outputs(2977) <= not a;
    layer1_outputs(2978) <= '1';
    layer1_outputs(2979) <= a or b;
    layer1_outputs(2980) <= not a;
    layer1_outputs(2981) <= b;
    layer1_outputs(2982) <= b and not a;
    layer1_outputs(2983) <= not (a and b);
    layer1_outputs(2984) <= a xor b;
    layer1_outputs(2985) <= not (a and b);
    layer1_outputs(2986) <= not a or b;
    layer1_outputs(2987) <= not a or b;
    layer1_outputs(2988) <= b;
    layer1_outputs(2989) <= '0';
    layer1_outputs(2990) <= not b;
    layer1_outputs(2991) <= a xor b;
    layer1_outputs(2992) <= a and not b;
    layer1_outputs(2993) <= b and not a;
    layer1_outputs(2994) <= a and not b;
    layer1_outputs(2995) <= a and b;
    layer1_outputs(2996) <= not (a and b);
    layer1_outputs(2997) <= not a;
    layer1_outputs(2998) <= b and not a;
    layer1_outputs(2999) <= '1';
    layer1_outputs(3000) <= '0';
    layer1_outputs(3001) <= '1';
    layer1_outputs(3002) <= a or b;
    layer1_outputs(3003) <= not (a or b);
    layer1_outputs(3004) <= not (a xor b);
    layer1_outputs(3005) <= a and not b;
    layer1_outputs(3006) <= not b;
    layer1_outputs(3007) <= not (a xor b);
    layer1_outputs(3008) <= not b or a;
    layer1_outputs(3009) <= a;
    layer1_outputs(3010) <= not b;
    layer1_outputs(3011) <= a;
    layer1_outputs(3012) <= not (a xor b);
    layer1_outputs(3013) <= a or b;
    layer1_outputs(3014) <= not b or a;
    layer1_outputs(3015) <= not a or b;
    layer1_outputs(3016) <= b;
    layer1_outputs(3017) <= not b;
    layer1_outputs(3018) <= b and not a;
    layer1_outputs(3019) <= a;
    layer1_outputs(3020) <= not b or a;
    layer1_outputs(3021) <= a or b;
    layer1_outputs(3022) <= b and not a;
    layer1_outputs(3023) <= not b;
    layer1_outputs(3024) <= a;
    layer1_outputs(3025) <= not (a and b);
    layer1_outputs(3026) <= not a;
    layer1_outputs(3027) <= a and not b;
    layer1_outputs(3028) <= not a or b;
    layer1_outputs(3029) <= b and not a;
    layer1_outputs(3030) <= not (a xor b);
    layer1_outputs(3031) <= b;
    layer1_outputs(3032) <= a and b;
    layer1_outputs(3033) <= not b or a;
    layer1_outputs(3034) <= '1';
    layer1_outputs(3035) <= b and not a;
    layer1_outputs(3036) <= a;
    layer1_outputs(3037) <= '0';
    layer1_outputs(3038) <= '0';
    layer1_outputs(3039) <= a;
    layer1_outputs(3040) <= not (a or b);
    layer1_outputs(3041) <= not b or a;
    layer1_outputs(3042) <= a and b;
    layer1_outputs(3043) <= '1';
    layer1_outputs(3044) <= not (a and b);
    layer1_outputs(3045) <= a or b;
    layer1_outputs(3046) <= not (a and b);
    layer1_outputs(3047) <= not b or a;
    layer1_outputs(3048) <= a and b;
    layer1_outputs(3049) <= not a;
    layer1_outputs(3050) <= a and b;
    layer1_outputs(3051) <= '0';
    layer1_outputs(3052) <= b and not a;
    layer1_outputs(3053) <= not (a or b);
    layer1_outputs(3054) <= '0';
    layer1_outputs(3055) <= not a or b;
    layer1_outputs(3056) <= a and b;
    layer1_outputs(3057) <= b;
    layer1_outputs(3058) <= b;
    layer1_outputs(3059) <= not a or b;
    layer1_outputs(3060) <= a;
    layer1_outputs(3061) <= not (a and b);
    layer1_outputs(3062) <= b;
    layer1_outputs(3063) <= not a;
    layer1_outputs(3064) <= not a;
    layer1_outputs(3065) <= '1';
    layer1_outputs(3066) <= not (a and b);
    layer1_outputs(3067) <= not b;
    layer1_outputs(3068) <= '1';
    layer1_outputs(3069) <= a or b;
    layer1_outputs(3070) <= a and b;
    layer1_outputs(3071) <= b;
    layer1_outputs(3072) <= b;
    layer1_outputs(3073) <= not a or b;
    layer1_outputs(3074) <= a and b;
    layer1_outputs(3075) <= '1';
    layer1_outputs(3076) <= not b or a;
    layer1_outputs(3077) <= not b or a;
    layer1_outputs(3078) <= b;
    layer1_outputs(3079) <= not a;
    layer1_outputs(3080) <= a;
    layer1_outputs(3081) <= a;
    layer1_outputs(3082) <= b and not a;
    layer1_outputs(3083) <= a or b;
    layer1_outputs(3084) <= not (a and b);
    layer1_outputs(3085) <= not a;
    layer1_outputs(3086) <= not b;
    layer1_outputs(3087) <= not a;
    layer1_outputs(3088) <= not b;
    layer1_outputs(3089) <= not a or b;
    layer1_outputs(3090) <= '1';
    layer1_outputs(3091) <= b;
    layer1_outputs(3092) <= not a;
    layer1_outputs(3093) <= not (a and b);
    layer1_outputs(3094) <= not (a or b);
    layer1_outputs(3095) <= not b or a;
    layer1_outputs(3096) <= a;
    layer1_outputs(3097) <= not b;
    layer1_outputs(3098) <= not a;
    layer1_outputs(3099) <= a;
    layer1_outputs(3100) <= not b;
    layer1_outputs(3101) <= not (a or b);
    layer1_outputs(3102) <= not b or a;
    layer1_outputs(3103) <= a or b;
    layer1_outputs(3104) <= not (a xor b);
    layer1_outputs(3105) <= not b or a;
    layer1_outputs(3106) <= not a;
    layer1_outputs(3107) <= not b;
    layer1_outputs(3108) <= a;
    layer1_outputs(3109) <= not a;
    layer1_outputs(3110) <= '0';
    layer1_outputs(3111) <= not (a and b);
    layer1_outputs(3112) <= not a or b;
    layer1_outputs(3113) <= not (a and b);
    layer1_outputs(3114) <= not (a xor b);
    layer1_outputs(3115) <= a;
    layer1_outputs(3116) <= '1';
    layer1_outputs(3117) <= '1';
    layer1_outputs(3118) <= b;
    layer1_outputs(3119) <= a;
    layer1_outputs(3120) <= not (a xor b);
    layer1_outputs(3121) <= not b or a;
    layer1_outputs(3122) <= not (a or b);
    layer1_outputs(3123) <= b and not a;
    layer1_outputs(3124) <= a;
    layer1_outputs(3125) <= not (a or b);
    layer1_outputs(3126) <= '0';
    layer1_outputs(3127) <= a and b;
    layer1_outputs(3128) <= b;
    layer1_outputs(3129) <= a and not b;
    layer1_outputs(3130) <= b and not a;
    layer1_outputs(3131) <= not a;
    layer1_outputs(3132) <= not (a and b);
    layer1_outputs(3133) <= not b or a;
    layer1_outputs(3134) <= '0';
    layer1_outputs(3135) <= not (a or b);
    layer1_outputs(3136) <= '0';
    layer1_outputs(3137) <= not (a and b);
    layer1_outputs(3138) <= not (a or b);
    layer1_outputs(3139) <= a and not b;
    layer1_outputs(3140) <= not (a and b);
    layer1_outputs(3141) <= not b;
    layer1_outputs(3142) <= not b;
    layer1_outputs(3143) <= not a or b;
    layer1_outputs(3144) <= a;
    layer1_outputs(3145) <= not (a or b);
    layer1_outputs(3146) <= a;
    layer1_outputs(3147) <= b and not a;
    layer1_outputs(3148) <= not b;
    layer1_outputs(3149) <= '1';
    layer1_outputs(3150) <= a or b;
    layer1_outputs(3151) <= b;
    layer1_outputs(3152) <= a and not b;
    layer1_outputs(3153) <= b and not a;
    layer1_outputs(3154) <= b;
    layer1_outputs(3155) <= a or b;
    layer1_outputs(3156) <= not b;
    layer1_outputs(3157) <= a and b;
    layer1_outputs(3158) <= '0';
    layer1_outputs(3159) <= b;
    layer1_outputs(3160) <= not (a or b);
    layer1_outputs(3161) <= '0';
    layer1_outputs(3162) <= a or b;
    layer1_outputs(3163) <= a;
    layer1_outputs(3164) <= b;
    layer1_outputs(3165) <= a or b;
    layer1_outputs(3166) <= not b or a;
    layer1_outputs(3167) <= '1';
    layer1_outputs(3168) <= a and not b;
    layer1_outputs(3169) <= b;
    layer1_outputs(3170) <= not b;
    layer1_outputs(3171) <= not (a xor b);
    layer1_outputs(3172) <= b and not a;
    layer1_outputs(3173) <= a and not b;
    layer1_outputs(3174) <= '1';
    layer1_outputs(3175) <= '1';
    layer1_outputs(3176) <= '1';
    layer1_outputs(3177) <= '0';
    layer1_outputs(3178) <= b and not a;
    layer1_outputs(3179) <= not a or b;
    layer1_outputs(3180) <= not (a or b);
    layer1_outputs(3181) <= not b or a;
    layer1_outputs(3182) <= '0';
    layer1_outputs(3183) <= b and not a;
    layer1_outputs(3184) <= not b;
    layer1_outputs(3185) <= not (a and b);
    layer1_outputs(3186) <= b and not a;
    layer1_outputs(3187) <= a or b;
    layer1_outputs(3188) <= '1';
    layer1_outputs(3189) <= not a or b;
    layer1_outputs(3190) <= not b or a;
    layer1_outputs(3191) <= b;
    layer1_outputs(3192) <= not (a or b);
    layer1_outputs(3193) <= not (a and b);
    layer1_outputs(3194) <= not a or b;
    layer1_outputs(3195) <= not (a and b);
    layer1_outputs(3196) <= not a;
    layer1_outputs(3197) <= not b or a;
    layer1_outputs(3198) <= a or b;
    layer1_outputs(3199) <= '1';
    layer1_outputs(3200) <= not (a xor b);
    layer1_outputs(3201) <= '0';
    layer1_outputs(3202) <= b and not a;
    layer1_outputs(3203) <= a and b;
    layer1_outputs(3204) <= not a or b;
    layer1_outputs(3205) <= not b or a;
    layer1_outputs(3206) <= not a;
    layer1_outputs(3207) <= b;
    layer1_outputs(3208) <= '1';
    layer1_outputs(3209) <= a or b;
    layer1_outputs(3210) <= '0';
    layer1_outputs(3211) <= a and b;
    layer1_outputs(3212) <= a xor b;
    layer1_outputs(3213) <= not b or a;
    layer1_outputs(3214) <= a;
    layer1_outputs(3215) <= a and b;
    layer1_outputs(3216) <= not (a xor b);
    layer1_outputs(3217) <= a or b;
    layer1_outputs(3218) <= a and b;
    layer1_outputs(3219) <= not (a or b);
    layer1_outputs(3220) <= b;
    layer1_outputs(3221) <= b;
    layer1_outputs(3222) <= not b;
    layer1_outputs(3223) <= a or b;
    layer1_outputs(3224) <= not a;
    layer1_outputs(3225) <= b and not a;
    layer1_outputs(3226) <= not (a or b);
    layer1_outputs(3227) <= b and not a;
    layer1_outputs(3228) <= not (a or b);
    layer1_outputs(3229) <= not b;
    layer1_outputs(3230) <= not b;
    layer1_outputs(3231) <= a and not b;
    layer1_outputs(3232) <= not a;
    layer1_outputs(3233) <= a;
    layer1_outputs(3234) <= not b;
    layer1_outputs(3235) <= not (a or b);
    layer1_outputs(3236) <= b and not a;
    layer1_outputs(3237) <= a and not b;
    layer1_outputs(3238) <= not a or b;
    layer1_outputs(3239) <= not a or b;
    layer1_outputs(3240) <= a;
    layer1_outputs(3241) <= b and not a;
    layer1_outputs(3242) <= not b or a;
    layer1_outputs(3243) <= not (a xor b);
    layer1_outputs(3244) <= not (a or b);
    layer1_outputs(3245) <= a or b;
    layer1_outputs(3246) <= not a;
    layer1_outputs(3247) <= a and not b;
    layer1_outputs(3248) <= b;
    layer1_outputs(3249) <= not a or b;
    layer1_outputs(3250) <= not (a or b);
    layer1_outputs(3251) <= '0';
    layer1_outputs(3252) <= a;
    layer1_outputs(3253) <= '1';
    layer1_outputs(3254) <= a xor b;
    layer1_outputs(3255) <= a and not b;
    layer1_outputs(3256) <= b;
    layer1_outputs(3257) <= '0';
    layer1_outputs(3258) <= not a;
    layer1_outputs(3259) <= not (a or b);
    layer1_outputs(3260) <= a;
    layer1_outputs(3261) <= a or b;
    layer1_outputs(3262) <= not (a or b);
    layer1_outputs(3263) <= b and not a;
    layer1_outputs(3264) <= b and not a;
    layer1_outputs(3265) <= not (a or b);
    layer1_outputs(3266) <= not b;
    layer1_outputs(3267) <= b and not a;
    layer1_outputs(3268) <= '0';
    layer1_outputs(3269) <= a;
    layer1_outputs(3270) <= not (a and b);
    layer1_outputs(3271) <= a and b;
    layer1_outputs(3272) <= not b;
    layer1_outputs(3273) <= b;
    layer1_outputs(3274) <= not a or b;
    layer1_outputs(3275) <= not b or a;
    layer1_outputs(3276) <= a and b;
    layer1_outputs(3277) <= not a;
    layer1_outputs(3278) <= a and not b;
    layer1_outputs(3279) <= a;
    layer1_outputs(3280) <= not (a xor b);
    layer1_outputs(3281) <= not a or b;
    layer1_outputs(3282) <= '0';
    layer1_outputs(3283) <= not (a or b);
    layer1_outputs(3284) <= a and b;
    layer1_outputs(3285) <= a and not b;
    layer1_outputs(3286) <= a;
    layer1_outputs(3287) <= a and b;
    layer1_outputs(3288) <= b and not a;
    layer1_outputs(3289) <= not (a or b);
    layer1_outputs(3290) <= not a;
    layer1_outputs(3291) <= '1';
    layer1_outputs(3292) <= b and not a;
    layer1_outputs(3293) <= b;
    layer1_outputs(3294) <= not b;
    layer1_outputs(3295) <= a and b;
    layer1_outputs(3296) <= not (a and b);
    layer1_outputs(3297) <= not b or a;
    layer1_outputs(3298) <= a and b;
    layer1_outputs(3299) <= '0';
    layer1_outputs(3300) <= b;
    layer1_outputs(3301) <= not (a or b);
    layer1_outputs(3302) <= not a or b;
    layer1_outputs(3303) <= not b or a;
    layer1_outputs(3304) <= '0';
    layer1_outputs(3305) <= '1';
    layer1_outputs(3306) <= a or b;
    layer1_outputs(3307) <= a and b;
    layer1_outputs(3308) <= '0';
    layer1_outputs(3309) <= '1';
    layer1_outputs(3310) <= '0';
    layer1_outputs(3311) <= not b or a;
    layer1_outputs(3312) <= b and not a;
    layer1_outputs(3313) <= not a;
    layer1_outputs(3314) <= b and not a;
    layer1_outputs(3315) <= not b;
    layer1_outputs(3316) <= b;
    layer1_outputs(3317) <= not (a and b);
    layer1_outputs(3318) <= not b;
    layer1_outputs(3319) <= a;
    layer1_outputs(3320) <= not (a and b);
    layer1_outputs(3321) <= a;
    layer1_outputs(3322) <= not a;
    layer1_outputs(3323) <= not (a xor b);
    layer1_outputs(3324) <= not a;
    layer1_outputs(3325) <= b and not a;
    layer1_outputs(3326) <= a;
    layer1_outputs(3327) <= not b;
    layer1_outputs(3328) <= not b;
    layer1_outputs(3329) <= not b;
    layer1_outputs(3330) <= a or b;
    layer1_outputs(3331) <= not (a and b);
    layer1_outputs(3332) <= a and not b;
    layer1_outputs(3333) <= not b;
    layer1_outputs(3334) <= not b;
    layer1_outputs(3335) <= '0';
    layer1_outputs(3336) <= b and not a;
    layer1_outputs(3337) <= not b or a;
    layer1_outputs(3338) <= a or b;
    layer1_outputs(3339) <= a xor b;
    layer1_outputs(3340) <= a and not b;
    layer1_outputs(3341) <= b;
    layer1_outputs(3342) <= b;
    layer1_outputs(3343) <= '0';
    layer1_outputs(3344) <= '0';
    layer1_outputs(3345) <= a and not b;
    layer1_outputs(3346) <= b;
    layer1_outputs(3347) <= a;
    layer1_outputs(3348) <= not a or b;
    layer1_outputs(3349) <= a or b;
    layer1_outputs(3350) <= not (a and b);
    layer1_outputs(3351) <= '1';
    layer1_outputs(3352) <= not a or b;
    layer1_outputs(3353) <= b;
    layer1_outputs(3354) <= '0';
    layer1_outputs(3355) <= not (a or b);
    layer1_outputs(3356) <= a and not b;
    layer1_outputs(3357) <= not a or b;
    layer1_outputs(3358) <= not b or a;
    layer1_outputs(3359) <= not (a xor b);
    layer1_outputs(3360) <= '0';
    layer1_outputs(3361) <= not b or a;
    layer1_outputs(3362) <= b and not a;
    layer1_outputs(3363) <= not b or a;
    layer1_outputs(3364) <= a and b;
    layer1_outputs(3365) <= a;
    layer1_outputs(3366) <= a and b;
    layer1_outputs(3367) <= not b or a;
    layer1_outputs(3368) <= a and b;
    layer1_outputs(3369) <= a or b;
    layer1_outputs(3370) <= b;
    layer1_outputs(3371) <= b and not a;
    layer1_outputs(3372) <= not (a or b);
    layer1_outputs(3373) <= not (a or b);
    layer1_outputs(3374) <= '1';
    layer1_outputs(3375) <= not (a xor b);
    layer1_outputs(3376) <= a and b;
    layer1_outputs(3377) <= not b;
    layer1_outputs(3378) <= not (a and b);
    layer1_outputs(3379) <= a;
    layer1_outputs(3380) <= b;
    layer1_outputs(3381) <= not a or b;
    layer1_outputs(3382) <= not a;
    layer1_outputs(3383) <= not a or b;
    layer1_outputs(3384) <= b and not a;
    layer1_outputs(3385) <= a and not b;
    layer1_outputs(3386) <= not b;
    layer1_outputs(3387) <= a and b;
    layer1_outputs(3388) <= not b;
    layer1_outputs(3389) <= a;
    layer1_outputs(3390) <= not a or b;
    layer1_outputs(3391) <= a and not b;
    layer1_outputs(3392) <= '0';
    layer1_outputs(3393) <= a xor b;
    layer1_outputs(3394) <= not a or b;
    layer1_outputs(3395) <= '1';
    layer1_outputs(3396) <= b and not a;
    layer1_outputs(3397) <= '0';
    layer1_outputs(3398) <= not a;
    layer1_outputs(3399) <= a and not b;
    layer1_outputs(3400) <= a or b;
    layer1_outputs(3401) <= not b or a;
    layer1_outputs(3402) <= b and not a;
    layer1_outputs(3403) <= b and not a;
    layer1_outputs(3404) <= not a;
    layer1_outputs(3405) <= not a or b;
    layer1_outputs(3406) <= '0';
    layer1_outputs(3407) <= '0';
    layer1_outputs(3408) <= not a or b;
    layer1_outputs(3409) <= b and not a;
    layer1_outputs(3410) <= a and b;
    layer1_outputs(3411) <= '0';
    layer1_outputs(3412) <= '0';
    layer1_outputs(3413) <= a or b;
    layer1_outputs(3414) <= b and not a;
    layer1_outputs(3415) <= a and b;
    layer1_outputs(3416) <= b and not a;
    layer1_outputs(3417) <= not (a and b);
    layer1_outputs(3418) <= not (a xor b);
    layer1_outputs(3419) <= not a or b;
    layer1_outputs(3420) <= not a or b;
    layer1_outputs(3421) <= a;
    layer1_outputs(3422) <= not a or b;
    layer1_outputs(3423) <= b;
    layer1_outputs(3424) <= not b or a;
    layer1_outputs(3425) <= b;
    layer1_outputs(3426) <= not (a or b);
    layer1_outputs(3427) <= not a;
    layer1_outputs(3428) <= not b or a;
    layer1_outputs(3429) <= '1';
    layer1_outputs(3430) <= not (a or b);
    layer1_outputs(3431) <= a;
    layer1_outputs(3432) <= a and b;
    layer1_outputs(3433) <= a and b;
    layer1_outputs(3434) <= not (a and b);
    layer1_outputs(3435) <= not (a or b);
    layer1_outputs(3436) <= '1';
    layer1_outputs(3437) <= a and not b;
    layer1_outputs(3438) <= not a;
    layer1_outputs(3439) <= not a or b;
    layer1_outputs(3440) <= a;
    layer1_outputs(3441) <= not a or b;
    layer1_outputs(3442) <= a and b;
    layer1_outputs(3443) <= a;
    layer1_outputs(3444) <= not a;
    layer1_outputs(3445) <= a xor b;
    layer1_outputs(3446) <= '0';
    layer1_outputs(3447) <= a and not b;
    layer1_outputs(3448) <= a;
    layer1_outputs(3449) <= '0';
    layer1_outputs(3450) <= b;
    layer1_outputs(3451) <= not b;
    layer1_outputs(3452) <= not a or b;
    layer1_outputs(3453) <= not b or a;
    layer1_outputs(3454) <= '1';
    layer1_outputs(3455) <= not a;
    layer1_outputs(3456) <= not b;
    layer1_outputs(3457) <= '0';
    layer1_outputs(3458) <= not (a or b);
    layer1_outputs(3459) <= not b;
    layer1_outputs(3460) <= a and b;
    layer1_outputs(3461) <= not (a xor b);
    layer1_outputs(3462) <= not a;
    layer1_outputs(3463) <= not (a or b);
    layer1_outputs(3464) <= not a;
    layer1_outputs(3465) <= not b;
    layer1_outputs(3466) <= b and not a;
    layer1_outputs(3467) <= a or b;
    layer1_outputs(3468) <= '1';
    layer1_outputs(3469) <= a and not b;
    layer1_outputs(3470) <= not b or a;
    layer1_outputs(3471) <= not (a or b);
    layer1_outputs(3472) <= not b;
    layer1_outputs(3473) <= not (a or b);
    layer1_outputs(3474) <= not (a and b);
    layer1_outputs(3475) <= not (a or b);
    layer1_outputs(3476) <= b and not a;
    layer1_outputs(3477) <= not (a xor b);
    layer1_outputs(3478) <= b and not a;
    layer1_outputs(3479) <= not (a and b);
    layer1_outputs(3480) <= b and not a;
    layer1_outputs(3481) <= not a or b;
    layer1_outputs(3482) <= a and not b;
    layer1_outputs(3483) <= not (a or b);
    layer1_outputs(3484) <= b and not a;
    layer1_outputs(3485) <= not a or b;
    layer1_outputs(3486) <= not (a xor b);
    layer1_outputs(3487) <= a or b;
    layer1_outputs(3488) <= not b;
    layer1_outputs(3489) <= a or b;
    layer1_outputs(3490) <= a;
    layer1_outputs(3491) <= a xor b;
    layer1_outputs(3492) <= not b;
    layer1_outputs(3493) <= b and not a;
    layer1_outputs(3494) <= a;
    layer1_outputs(3495) <= b and not a;
    layer1_outputs(3496) <= not b;
    layer1_outputs(3497) <= not a or b;
    layer1_outputs(3498) <= not (a or b);
    layer1_outputs(3499) <= not b or a;
    layer1_outputs(3500) <= not b;
    layer1_outputs(3501) <= b;
    layer1_outputs(3502) <= '1';
    layer1_outputs(3503) <= '0';
    layer1_outputs(3504) <= a or b;
    layer1_outputs(3505) <= not a;
    layer1_outputs(3506) <= b and not a;
    layer1_outputs(3507) <= a xor b;
    layer1_outputs(3508) <= not a;
    layer1_outputs(3509) <= not (a and b);
    layer1_outputs(3510) <= not b or a;
    layer1_outputs(3511) <= b and not a;
    layer1_outputs(3512) <= b and not a;
    layer1_outputs(3513) <= a and b;
    layer1_outputs(3514) <= a and b;
    layer1_outputs(3515) <= '0';
    layer1_outputs(3516) <= b;
    layer1_outputs(3517) <= a and b;
    layer1_outputs(3518) <= a and b;
    layer1_outputs(3519) <= not (a or b);
    layer1_outputs(3520) <= not a;
    layer1_outputs(3521) <= '0';
    layer1_outputs(3522) <= a;
    layer1_outputs(3523) <= '1';
    layer1_outputs(3524) <= not b or a;
    layer1_outputs(3525) <= a;
    layer1_outputs(3526) <= not a;
    layer1_outputs(3527) <= a and b;
    layer1_outputs(3528) <= a;
    layer1_outputs(3529) <= a or b;
    layer1_outputs(3530) <= b and not a;
    layer1_outputs(3531) <= not a;
    layer1_outputs(3532) <= not a;
    layer1_outputs(3533) <= b;
    layer1_outputs(3534) <= not a;
    layer1_outputs(3535) <= b and not a;
    layer1_outputs(3536) <= not (a and b);
    layer1_outputs(3537) <= a;
    layer1_outputs(3538) <= not b or a;
    layer1_outputs(3539) <= not b or a;
    layer1_outputs(3540) <= a or b;
    layer1_outputs(3541) <= not (a and b);
    layer1_outputs(3542) <= b and not a;
    layer1_outputs(3543) <= not (a xor b);
    layer1_outputs(3544) <= not (a and b);
    layer1_outputs(3545) <= not (a and b);
    layer1_outputs(3546) <= a or b;
    layer1_outputs(3547) <= not b or a;
    layer1_outputs(3548) <= b;
    layer1_outputs(3549) <= not (a and b);
    layer1_outputs(3550) <= b;
    layer1_outputs(3551) <= a and not b;
    layer1_outputs(3552) <= b and not a;
    layer1_outputs(3553) <= not a;
    layer1_outputs(3554) <= not (a or b);
    layer1_outputs(3555) <= b and not a;
    layer1_outputs(3556) <= not (a or b);
    layer1_outputs(3557) <= not a or b;
    layer1_outputs(3558) <= not (a xor b);
    layer1_outputs(3559) <= not (a and b);
    layer1_outputs(3560) <= not b;
    layer1_outputs(3561) <= not a or b;
    layer1_outputs(3562) <= '0';
    layer1_outputs(3563) <= not a;
    layer1_outputs(3564) <= not (a or b);
    layer1_outputs(3565) <= a and not b;
    layer1_outputs(3566) <= '0';
    layer1_outputs(3567) <= not (a and b);
    layer1_outputs(3568) <= not (a or b);
    layer1_outputs(3569) <= '1';
    layer1_outputs(3570) <= not (a xor b);
    layer1_outputs(3571) <= a;
    layer1_outputs(3572) <= a and not b;
    layer1_outputs(3573) <= b;
    layer1_outputs(3574) <= a and not b;
    layer1_outputs(3575) <= not a or b;
    layer1_outputs(3576) <= not b;
    layer1_outputs(3577) <= not b or a;
    layer1_outputs(3578) <= a and not b;
    layer1_outputs(3579) <= not a;
    layer1_outputs(3580) <= not b;
    layer1_outputs(3581) <= not b or a;
    layer1_outputs(3582) <= not b or a;
    layer1_outputs(3583) <= not (a xor b);
    layer1_outputs(3584) <= not (a and b);
    layer1_outputs(3585) <= not a;
    layer1_outputs(3586) <= '0';
    layer1_outputs(3587) <= a or b;
    layer1_outputs(3588) <= not (a or b);
    layer1_outputs(3589) <= b and not a;
    layer1_outputs(3590) <= '0';
    layer1_outputs(3591) <= not b;
    layer1_outputs(3592) <= a and b;
    layer1_outputs(3593) <= not b or a;
    layer1_outputs(3594) <= not (a or b);
    layer1_outputs(3595) <= not (a or b);
    layer1_outputs(3596) <= '1';
    layer1_outputs(3597) <= '0';
    layer1_outputs(3598) <= b;
    layer1_outputs(3599) <= not a;
    layer1_outputs(3600) <= a or b;
    layer1_outputs(3601) <= '0';
    layer1_outputs(3602) <= '0';
    layer1_outputs(3603) <= a and b;
    layer1_outputs(3604) <= '1';
    layer1_outputs(3605) <= '1';
    layer1_outputs(3606) <= not (a xor b);
    layer1_outputs(3607) <= a or b;
    layer1_outputs(3608) <= a and not b;
    layer1_outputs(3609) <= not b;
    layer1_outputs(3610) <= b;
    layer1_outputs(3611) <= not a;
    layer1_outputs(3612) <= not (a xor b);
    layer1_outputs(3613) <= not b;
    layer1_outputs(3614) <= not a;
    layer1_outputs(3615) <= a and not b;
    layer1_outputs(3616) <= not b;
    layer1_outputs(3617) <= not (a and b);
    layer1_outputs(3618) <= not a or b;
    layer1_outputs(3619) <= a or b;
    layer1_outputs(3620) <= a;
    layer1_outputs(3621) <= a;
    layer1_outputs(3622) <= not (a or b);
    layer1_outputs(3623) <= b and not a;
    layer1_outputs(3624) <= b;
    layer1_outputs(3625) <= a and not b;
    layer1_outputs(3626) <= not (a and b);
    layer1_outputs(3627) <= not b or a;
    layer1_outputs(3628) <= b and not a;
    layer1_outputs(3629) <= b and not a;
    layer1_outputs(3630) <= a;
    layer1_outputs(3631) <= not b;
    layer1_outputs(3632) <= not a or b;
    layer1_outputs(3633) <= not b or a;
    layer1_outputs(3634) <= not b or a;
    layer1_outputs(3635) <= not a;
    layer1_outputs(3636) <= not a;
    layer1_outputs(3637) <= a and b;
    layer1_outputs(3638) <= '1';
    layer1_outputs(3639) <= '1';
    layer1_outputs(3640) <= b and not a;
    layer1_outputs(3641) <= not a;
    layer1_outputs(3642) <= not b;
    layer1_outputs(3643) <= a;
    layer1_outputs(3644) <= not b or a;
    layer1_outputs(3645) <= '0';
    layer1_outputs(3646) <= '0';
    layer1_outputs(3647) <= not b or a;
    layer1_outputs(3648) <= not (a or b);
    layer1_outputs(3649) <= not (a xor b);
    layer1_outputs(3650) <= a and not b;
    layer1_outputs(3651) <= '0';
    layer1_outputs(3652) <= a and not b;
    layer1_outputs(3653) <= not a;
    layer1_outputs(3654) <= a;
    layer1_outputs(3655) <= a xor b;
    layer1_outputs(3656) <= not b;
    layer1_outputs(3657) <= not (a or b);
    layer1_outputs(3658) <= not b or a;
    layer1_outputs(3659) <= a or b;
    layer1_outputs(3660) <= not a or b;
    layer1_outputs(3661) <= '0';
    layer1_outputs(3662) <= '1';
    layer1_outputs(3663) <= '0';
    layer1_outputs(3664) <= not b or a;
    layer1_outputs(3665) <= a and b;
    layer1_outputs(3666) <= a and b;
    layer1_outputs(3667) <= a and not b;
    layer1_outputs(3668) <= not b;
    layer1_outputs(3669) <= not a;
    layer1_outputs(3670) <= a xor b;
    layer1_outputs(3671) <= not b;
    layer1_outputs(3672) <= not (a xor b);
    layer1_outputs(3673) <= not b or a;
    layer1_outputs(3674) <= b;
    layer1_outputs(3675) <= not b;
    layer1_outputs(3676) <= not (a or b);
    layer1_outputs(3677) <= not (a or b);
    layer1_outputs(3678) <= b and not a;
    layer1_outputs(3679) <= not (a and b);
    layer1_outputs(3680) <= a;
    layer1_outputs(3681) <= a xor b;
    layer1_outputs(3682) <= not a or b;
    layer1_outputs(3683) <= not (a xor b);
    layer1_outputs(3684) <= '1';
    layer1_outputs(3685) <= not (a and b);
    layer1_outputs(3686) <= not b;
    layer1_outputs(3687) <= not (a or b);
    layer1_outputs(3688) <= not b;
    layer1_outputs(3689) <= b and not a;
    layer1_outputs(3690) <= '0';
    layer1_outputs(3691) <= not (a and b);
    layer1_outputs(3692) <= a and not b;
    layer1_outputs(3693) <= not (a and b);
    layer1_outputs(3694) <= a;
    layer1_outputs(3695) <= not (a and b);
    layer1_outputs(3696) <= not (a or b);
    layer1_outputs(3697) <= not a;
    layer1_outputs(3698) <= a and b;
    layer1_outputs(3699) <= not b;
    layer1_outputs(3700) <= not a;
    layer1_outputs(3701) <= not b or a;
    layer1_outputs(3702) <= '0';
    layer1_outputs(3703) <= a xor b;
    layer1_outputs(3704) <= a or b;
    layer1_outputs(3705) <= not a or b;
    layer1_outputs(3706) <= not a;
    layer1_outputs(3707) <= not a or b;
    layer1_outputs(3708) <= not b or a;
    layer1_outputs(3709) <= not (a and b);
    layer1_outputs(3710) <= not (a or b);
    layer1_outputs(3711) <= not b;
    layer1_outputs(3712) <= not (a or b);
    layer1_outputs(3713) <= a or b;
    layer1_outputs(3714) <= not (a and b);
    layer1_outputs(3715) <= '1';
    layer1_outputs(3716) <= a and b;
    layer1_outputs(3717) <= not (a and b);
    layer1_outputs(3718) <= a and not b;
    layer1_outputs(3719) <= b and not a;
    layer1_outputs(3720) <= '1';
    layer1_outputs(3721) <= '1';
    layer1_outputs(3722) <= a xor b;
    layer1_outputs(3723) <= a or b;
    layer1_outputs(3724) <= not (a or b);
    layer1_outputs(3725) <= not (a or b);
    layer1_outputs(3726) <= a;
    layer1_outputs(3727) <= not (a or b);
    layer1_outputs(3728) <= not (a and b);
    layer1_outputs(3729) <= not a or b;
    layer1_outputs(3730) <= '1';
    layer1_outputs(3731) <= '1';
    layer1_outputs(3732) <= a and not b;
    layer1_outputs(3733) <= not b or a;
    layer1_outputs(3734) <= a and b;
    layer1_outputs(3735) <= not (a and b);
    layer1_outputs(3736) <= '1';
    layer1_outputs(3737) <= a;
    layer1_outputs(3738) <= a;
    layer1_outputs(3739) <= a and not b;
    layer1_outputs(3740) <= '0';
    layer1_outputs(3741) <= a xor b;
    layer1_outputs(3742) <= not b or a;
    layer1_outputs(3743) <= a and b;
    layer1_outputs(3744) <= not (a or b);
    layer1_outputs(3745) <= a and not b;
    layer1_outputs(3746) <= not a;
    layer1_outputs(3747) <= a and not b;
    layer1_outputs(3748) <= a xor b;
    layer1_outputs(3749) <= not (a and b);
    layer1_outputs(3750) <= not a;
    layer1_outputs(3751) <= b and not a;
    layer1_outputs(3752) <= not b;
    layer1_outputs(3753) <= a and not b;
    layer1_outputs(3754) <= a;
    layer1_outputs(3755) <= not b;
    layer1_outputs(3756) <= not b;
    layer1_outputs(3757) <= b and not a;
    layer1_outputs(3758) <= a;
    layer1_outputs(3759) <= not (a xor b);
    layer1_outputs(3760) <= a;
    layer1_outputs(3761) <= not a or b;
    layer1_outputs(3762) <= not a or b;
    layer1_outputs(3763) <= not (a and b);
    layer1_outputs(3764) <= not (a and b);
    layer1_outputs(3765) <= a or b;
    layer1_outputs(3766) <= not (a or b);
    layer1_outputs(3767) <= a xor b;
    layer1_outputs(3768) <= a and not b;
    layer1_outputs(3769) <= not (a and b);
    layer1_outputs(3770) <= not a or b;
    layer1_outputs(3771) <= a or b;
    layer1_outputs(3772) <= not b;
    layer1_outputs(3773) <= a;
    layer1_outputs(3774) <= not b;
    layer1_outputs(3775) <= b and not a;
    layer1_outputs(3776) <= not b;
    layer1_outputs(3777) <= a xor b;
    layer1_outputs(3778) <= b and not a;
    layer1_outputs(3779) <= not (a xor b);
    layer1_outputs(3780) <= b and not a;
    layer1_outputs(3781) <= not a;
    layer1_outputs(3782) <= a and not b;
    layer1_outputs(3783) <= not (a or b);
    layer1_outputs(3784) <= '1';
    layer1_outputs(3785) <= not b;
    layer1_outputs(3786) <= a or b;
    layer1_outputs(3787) <= a or b;
    layer1_outputs(3788) <= not (a and b);
    layer1_outputs(3789) <= a or b;
    layer1_outputs(3790) <= a xor b;
    layer1_outputs(3791) <= not b;
    layer1_outputs(3792) <= a and not b;
    layer1_outputs(3793) <= not b;
    layer1_outputs(3794) <= a;
    layer1_outputs(3795) <= not (a and b);
    layer1_outputs(3796) <= not (a and b);
    layer1_outputs(3797) <= '0';
    layer1_outputs(3798) <= not b;
    layer1_outputs(3799) <= a or b;
    layer1_outputs(3800) <= a xor b;
    layer1_outputs(3801) <= a xor b;
    layer1_outputs(3802) <= a or b;
    layer1_outputs(3803) <= a or b;
    layer1_outputs(3804) <= b and not a;
    layer1_outputs(3805) <= b and not a;
    layer1_outputs(3806) <= not b;
    layer1_outputs(3807) <= b;
    layer1_outputs(3808) <= a and not b;
    layer1_outputs(3809) <= '1';
    layer1_outputs(3810) <= b and not a;
    layer1_outputs(3811) <= not b or a;
    layer1_outputs(3812) <= b and not a;
    layer1_outputs(3813) <= a or b;
    layer1_outputs(3814) <= b;
    layer1_outputs(3815) <= a and not b;
    layer1_outputs(3816) <= not a or b;
    layer1_outputs(3817) <= not (a or b);
    layer1_outputs(3818) <= not b;
    layer1_outputs(3819) <= '1';
    layer1_outputs(3820) <= not a;
    layer1_outputs(3821) <= b;
    layer1_outputs(3822) <= not (a or b);
    layer1_outputs(3823) <= not b or a;
    layer1_outputs(3824) <= a and b;
    layer1_outputs(3825) <= not (a or b);
    layer1_outputs(3826) <= '1';
    layer1_outputs(3827) <= a or b;
    layer1_outputs(3828) <= not a;
    layer1_outputs(3829) <= a;
    layer1_outputs(3830) <= '0';
    layer1_outputs(3831) <= not b;
    layer1_outputs(3832) <= a and b;
    layer1_outputs(3833) <= a;
    layer1_outputs(3834) <= not a or b;
    layer1_outputs(3835) <= a or b;
    layer1_outputs(3836) <= a and not b;
    layer1_outputs(3837) <= a and b;
    layer1_outputs(3838) <= b and not a;
    layer1_outputs(3839) <= a or b;
    layer1_outputs(3840) <= not a;
    layer1_outputs(3841) <= b;
    layer1_outputs(3842) <= b;
    layer1_outputs(3843) <= b and not a;
    layer1_outputs(3844) <= a;
    layer1_outputs(3845) <= not (a or b);
    layer1_outputs(3846) <= not (a xor b);
    layer1_outputs(3847) <= a and b;
    layer1_outputs(3848) <= a xor b;
    layer1_outputs(3849) <= a;
    layer1_outputs(3850) <= a and not b;
    layer1_outputs(3851) <= not (a or b);
    layer1_outputs(3852) <= '1';
    layer1_outputs(3853) <= a and b;
    layer1_outputs(3854) <= a and b;
    layer1_outputs(3855) <= a or b;
    layer1_outputs(3856) <= not a or b;
    layer1_outputs(3857) <= b;
    layer1_outputs(3858) <= not a;
    layer1_outputs(3859) <= b;
    layer1_outputs(3860) <= not a;
    layer1_outputs(3861) <= not (a xor b);
    layer1_outputs(3862) <= a;
    layer1_outputs(3863) <= '0';
    layer1_outputs(3864) <= not (a and b);
    layer1_outputs(3865) <= not a or b;
    layer1_outputs(3866) <= not b;
    layer1_outputs(3867) <= '0';
    layer1_outputs(3868) <= a and b;
    layer1_outputs(3869) <= a and b;
    layer1_outputs(3870) <= a;
    layer1_outputs(3871) <= '1';
    layer1_outputs(3872) <= '1';
    layer1_outputs(3873) <= not b or a;
    layer1_outputs(3874) <= a xor b;
    layer1_outputs(3875) <= a;
    layer1_outputs(3876) <= not a;
    layer1_outputs(3877) <= not (a xor b);
    layer1_outputs(3878) <= not a;
    layer1_outputs(3879) <= not (a xor b);
    layer1_outputs(3880) <= not a;
    layer1_outputs(3881) <= a;
    layer1_outputs(3882) <= '1';
    layer1_outputs(3883) <= a and not b;
    layer1_outputs(3884) <= a and b;
    layer1_outputs(3885) <= a;
    layer1_outputs(3886) <= not b;
    layer1_outputs(3887) <= a;
    layer1_outputs(3888) <= a;
    layer1_outputs(3889) <= a;
    layer1_outputs(3890) <= a and b;
    layer1_outputs(3891) <= a and not b;
    layer1_outputs(3892) <= '0';
    layer1_outputs(3893) <= not b or a;
    layer1_outputs(3894) <= not b;
    layer1_outputs(3895) <= '0';
    layer1_outputs(3896) <= not a or b;
    layer1_outputs(3897) <= b;
    layer1_outputs(3898) <= a xor b;
    layer1_outputs(3899) <= not a;
    layer1_outputs(3900) <= a;
    layer1_outputs(3901) <= '1';
    layer1_outputs(3902) <= not (a and b);
    layer1_outputs(3903) <= a or b;
    layer1_outputs(3904) <= b and not a;
    layer1_outputs(3905) <= '1';
    layer1_outputs(3906) <= not (a and b);
    layer1_outputs(3907) <= a and not b;
    layer1_outputs(3908) <= not (a and b);
    layer1_outputs(3909) <= not (a or b);
    layer1_outputs(3910) <= not (a and b);
    layer1_outputs(3911) <= not b or a;
    layer1_outputs(3912) <= a and b;
    layer1_outputs(3913) <= b and not a;
    layer1_outputs(3914) <= not (a xor b);
    layer1_outputs(3915) <= not a;
    layer1_outputs(3916) <= not a;
    layer1_outputs(3917) <= a;
    layer1_outputs(3918) <= '0';
    layer1_outputs(3919) <= b;
    layer1_outputs(3920) <= '1';
    layer1_outputs(3921) <= a;
    layer1_outputs(3922) <= not (a and b);
    layer1_outputs(3923) <= a or b;
    layer1_outputs(3924) <= a and not b;
    layer1_outputs(3925) <= not (a xor b);
    layer1_outputs(3926) <= a and b;
    layer1_outputs(3927) <= b and not a;
    layer1_outputs(3928) <= not (a or b);
    layer1_outputs(3929) <= not b;
    layer1_outputs(3930) <= a;
    layer1_outputs(3931) <= a and not b;
    layer1_outputs(3932) <= not b;
    layer1_outputs(3933) <= a and not b;
    layer1_outputs(3934) <= a or b;
    layer1_outputs(3935) <= not a or b;
    layer1_outputs(3936) <= b;
    layer1_outputs(3937) <= not (a or b);
    layer1_outputs(3938) <= a xor b;
    layer1_outputs(3939) <= not (a and b);
    layer1_outputs(3940) <= a xor b;
    layer1_outputs(3941) <= '1';
    layer1_outputs(3942) <= not (a and b);
    layer1_outputs(3943) <= a and b;
    layer1_outputs(3944) <= not (a and b);
    layer1_outputs(3945) <= '0';
    layer1_outputs(3946) <= not b;
    layer1_outputs(3947) <= '0';
    layer1_outputs(3948) <= '1';
    layer1_outputs(3949) <= not b;
    layer1_outputs(3950) <= b;
    layer1_outputs(3951) <= not b;
    layer1_outputs(3952) <= not b or a;
    layer1_outputs(3953) <= not a;
    layer1_outputs(3954) <= a;
    layer1_outputs(3955) <= a and not b;
    layer1_outputs(3956) <= not a;
    layer1_outputs(3957) <= '0';
    layer1_outputs(3958) <= a and not b;
    layer1_outputs(3959) <= not b;
    layer1_outputs(3960) <= a or b;
    layer1_outputs(3961) <= a or b;
    layer1_outputs(3962) <= b and not a;
    layer1_outputs(3963) <= a and b;
    layer1_outputs(3964) <= a and b;
    layer1_outputs(3965) <= a;
    layer1_outputs(3966) <= a xor b;
    layer1_outputs(3967) <= a or b;
    layer1_outputs(3968) <= not (a and b);
    layer1_outputs(3969) <= not b or a;
    layer1_outputs(3970) <= b and not a;
    layer1_outputs(3971) <= '1';
    layer1_outputs(3972) <= not (a and b);
    layer1_outputs(3973) <= a;
    layer1_outputs(3974) <= a;
    layer1_outputs(3975) <= a or b;
    layer1_outputs(3976) <= a and not b;
    layer1_outputs(3977) <= not (a xor b);
    layer1_outputs(3978) <= a or b;
    layer1_outputs(3979) <= not (a or b);
    layer1_outputs(3980) <= '0';
    layer1_outputs(3981) <= not b;
    layer1_outputs(3982) <= '0';
    layer1_outputs(3983) <= not (a xor b);
    layer1_outputs(3984) <= not a or b;
    layer1_outputs(3985) <= a and b;
    layer1_outputs(3986) <= not b or a;
    layer1_outputs(3987) <= not b;
    layer1_outputs(3988) <= not b or a;
    layer1_outputs(3989) <= not b or a;
    layer1_outputs(3990) <= not (a or b);
    layer1_outputs(3991) <= '0';
    layer1_outputs(3992) <= b;
    layer1_outputs(3993) <= b;
    layer1_outputs(3994) <= not (a or b);
    layer1_outputs(3995) <= b;
    layer1_outputs(3996) <= a xor b;
    layer1_outputs(3997) <= a and not b;
    layer1_outputs(3998) <= '0';
    layer1_outputs(3999) <= not b;
    layer1_outputs(4000) <= a xor b;
    layer1_outputs(4001) <= not b or a;
    layer1_outputs(4002) <= not (a and b);
    layer1_outputs(4003) <= not b or a;
    layer1_outputs(4004) <= not a;
    layer1_outputs(4005) <= not a or b;
    layer1_outputs(4006) <= a and b;
    layer1_outputs(4007) <= a or b;
    layer1_outputs(4008) <= not b;
    layer1_outputs(4009) <= not a;
    layer1_outputs(4010) <= not a;
    layer1_outputs(4011) <= not b or a;
    layer1_outputs(4012) <= a and b;
    layer1_outputs(4013) <= not b;
    layer1_outputs(4014) <= '1';
    layer1_outputs(4015) <= a;
    layer1_outputs(4016) <= a and b;
    layer1_outputs(4017) <= a and b;
    layer1_outputs(4018) <= '1';
    layer1_outputs(4019) <= not (a and b);
    layer1_outputs(4020) <= a and b;
    layer1_outputs(4021) <= '0';
    layer1_outputs(4022) <= '0';
    layer1_outputs(4023) <= not b or a;
    layer1_outputs(4024) <= b;
    layer1_outputs(4025) <= a;
    layer1_outputs(4026) <= not a;
    layer1_outputs(4027) <= '0';
    layer1_outputs(4028) <= not a;
    layer1_outputs(4029) <= not a or b;
    layer1_outputs(4030) <= a and not b;
    layer1_outputs(4031) <= not b or a;
    layer1_outputs(4032) <= not b;
    layer1_outputs(4033) <= '1';
    layer1_outputs(4034) <= not a or b;
    layer1_outputs(4035) <= '0';
    layer1_outputs(4036) <= not (a and b);
    layer1_outputs(4037) <= a and not b;
    layer1_outputs(4038) <= not (a and b);
    layer1_outputs(4039) <= not a;
    layer1_outputs(4040) <= not (a and b);
    layer1_outputs(4041) <= a and b;
    layer1_outputs(4042) <= not (a or b);
    layer1_outputs(4043) <= a and not b;
    layer1_outputs(4044) <= a;
    layer1_outputs(4045) <= a or b;
    layer1_outputs(4046) <= '0';
    layer1_outputs(4047) <= not (a and b);
    layer1_outputs(4048) <= '1';
    layer1_outputs(4049) <= a or b;
    layer1_outputs(4050) <= not (a and b);
    layer1_outputs(4051) <= a;
    layer1_outputs(4052) <= not b or a;
    layer1_outputs(4053) <= not (a or b);
    layer1_outputs(4054) <= '1';
    layer1_outputs(4055) <= b;
    layer1_outputs(4056) <= not (a and b);
    layer1_outputs(4057) <= a and not b;
    layer1_outputs(4058) <= a and not b;
    layer1_outputs(4059) <= a and b;
    layer1_outputs(4060) <= a and not b;
    layer1_outputs(4061) <= a;
    layer1_outputs(4062) <= not a or b;
    layer1_outputs(4063) <= '1';
    layer1_outputs(4064) <= a or b;
    layer1_outputs(4065) <= b and not a;
    layer1_outputs(4066) <= not a or b;
    layer1_outputs(4067) <= b;
    layer1_outputs(4068) <= '1';
    layer1_outputs(4069) <= not b or a;
    layer1_outputs(4070) <= not b;
    layer1_outputs(4071) <= a;
    layer1_outputs(4072) <= a and b;
    layer1_outputs(4073) <= a or b;
    layer1_outputs(4074) <= '0';
    layer1_outputs(4075) <= not (a or b);
    layer1_outputs(4076) <= b and not a;
    layer1_outputs(4077) <= not b or a;
    layer1_outputs(4078) <= b and not a;
    layer1_outputs(4079) <= not b;
    layer1_outputs(4080) <= not (a xor b);
    layer1_outputs(4081) <= '1';
    layer1_outputs(4082) <= not (a or b);
    layer1_outputs(4083) <= a and b;
    layer1_outputs(4084) <= '1';
    layer1_outputs(4085) <= '0';
    layer1_outputs(4086) <= a and b;
    layer1_outputs(4087) <= a;
    layer1_outputs(4088) <= a and not b;
    layer1_outputs(4089) <= a xor b;
    layer1_outputs(4090) <= b and not a;
    layer1_outputs(4091) <= a and not b;
    layer1_outputs(4092) <= a;
    layer1_outputs(4093) <= not a or b;
    layer1_outputs(4094) <= not a;
    layer1_outputs(4095) <= not (a and b);
    layer1_outputs(4096) <= a or b;
    layer1_outputs(4097) <= '1';
    layer1_outputs(4098) <= b;
    layer1_outputs(4099) <= not (a xor b);
    layer1_outputs(4100) <= not b or a;
    layer1_outputs(4101) <= b and not a;
    layer1_outputs(4102) <= a;
    layer1_outputs(4103) <= b and not a;
    layer1_outputs(4104) <= a;
    layer1_outputs(4105) <= not (a or b);
    layer1_outputs(4106) <= not (a or b);
    layer1_outputs(4107) <= a and not b;
    layer1_outputs(4108) <= not (a or b);
    layer1_outputs(4109) <= not (a xor b);
    layer1_outputs(4110) <= not b;
    layer1_outputs(4111) <= not (a and b);
    layer1_outputs(4112) <= b;
    layer1_outputs(4113) <= b and not a;
    layer1_outputs(4114) <= b;
    layer1_outputs(4115) <= a;
    layer1_outputs(4116) <= not b or a;
    layer1_outputs(4117) <= a and b;
    layer1_outputs(4118) <= a;
    layer1_outputs(4119) <= not a or b;
    layer1_outputs(4120) <= not b or a;
    layer1_outputs(4121) <= not b;
    layer1_outputs(4122) <= not (a and b);
    layer1_outputs(4123) <= a;
    layer1_outputs(4124) <= a or b;
    layer1_outputs(4125) <= b and not a;
    layer1_outputs(4126) <= not b;
    layer1_outputs(4127) <= not a;
    layer1_outputs(4128) <= b;
    layer1_outputs(4129) <= a and b;
    layer1_outputs(4130) <= not b;
    layer1_outputs(4131) <= not (a or b);
    layer1_outputs(4132) <= not b or a;
    layer1_outputs(4133) <= '1';
    layer1_outputs(4134) <= not b;
    layer1_outputs(4135) <= a and b;
    layer1_outputs(4136) <= not a or b;
    layer1_outputs(4137) <= not (a xor b);
    layer1_outputs(4138) <= a or b;
    layer1_outputs(4139) <= not (a xor b);
    layer1_outputs(4140) <= not a or b;
    layer1_outputs(4141) <= a and b;
    layer1_outputs(4142) <= a xor b;
    layer1_outputs(4143) <= not b;
    layer1_outputs(4144) <= a xor b;
    layer1_outputs(4145) <= '1';
    layer1_outputs(4146) <= not a;
    layer1_outputs(4147) <= b and not a;
    layer1_outputs(4148) <= not a or b;
    layer1_outputs(4149) <= a or b;
    layer1_outputs(4150) <= not (a or b);
    layer1_outputs(4151) <= not a or b;
    layer1_outputs(4152) <= not (a or b);
    layer1_outputs(4153) <= a and not b;
    layer1_outputs(4154) <= not a or b;
    layer1_outputs(4155) <= a and b;
    layer1_outputs(4156) <= not a or b;
    layer1_outputs(4157) <= not (a or b);
    layer1_outputs(4158) <= a;
    layer1_outputs(4159) <= a or b;
    layer1_outputs(4160) <= a and b;
    layer1_outputs(4161) <= '1';
    layer1_outputs(4162) <= not (a xor b);
    layer1_outputs(4163) <= not b;
    layer1_outputs(4164) <= a;
    layer1_outputs(4165) <= not (a and b);
    layer1_outputs(4166) <= not a or b;
    layer1_outputs(4167) <= a or b;
    layer1_outputs(4168) <= not a;
    layer1_outputs(4169) <= not (a or b);
    layer1_outputs(4170) <= not b;
    layer1_outputs(4171) <= not (a or b);
    layer1_outputs(4172) <= a and not b;
    layer1_outputs(4173) <= not a;
    layer1_outputs(4174) <= a;
    layer1_outputs(4175) <= not (a or b);
    layer1_outputs(4176) <= '1';
    layer1_outputs(4177) <= not b or a;
    layer1_outputs(4178) <= not a;
    layer1_outputs(4179) <= not b or a;
    layer1_outputs(4180) <= a;
    layer1_outputs(4181) <= a and not b;
    layer1_outputs(4182) <= not b or a;
    layer1_outputs(4183) <= a and not b;
    layer1_outputs(4184) <= b;
    layer1_outputs(4185) <= a or b;
    layer1_outputs(4186) <= not a;
    layer1_outputs(4187) <= b;
    layer1_outputs(4188) <= not b or a;
    layer1_outputs(4189) <= not a;
    layer1_outputs(4190) <= a and not b;
    layer1_outputs(4191) <= '1';
    layer1_outputs(4192) <= not (a or b);
    layer1_outputs(4193) <= b;
    layer1_outputs(4194) <= a;
    layer1_outputs(4195) <= not (a or b);
    layer1_outputs(4196) <= b;
    layer1_outputs(4197) <= a and b;
    layer1_outputs(4198) <= not a;
    layer1_outputs(4199) <= not a or b;
    layer1_outputs(4200) <= not (a and b);
    layer1_outputs(4201) <= not b or a;
    layer1_outputs(4202) <= not (a or b);
    layer1_outputs(4203) <= b;
    layer1_outputs(4204) <= '0';
    layer1_outputs(4205) <= not b;
    layer1_outputs(4206) <= a xor b;
    layer1_outputs(4207) <= '0';
    layer1_outputs(4208) <= not b;
    layer1_outputs(4209) <= not a or b;
    layer1_outputs(4210) <= a;
    layer1_outputs(4211) <= not (a or b);
    layer1_outputs(4212) <= a and not b;
    layer1_outputs(4213) <= '0';
    layer1_outputs(4214) <= not a;
    layer1_outputs(4215) <= not a or b;
    layer1_outputs(4216) <= b;
    layer1_outputs(4217) <= '0';
    layer1_outputs(4218) <= not b or a;
    layer1_outputs(4219) <= b;
    layer1_outputs(4220) <= a or b;
    layer1_outputs(4221) <= not a;
    layer1_outputs(4222) <= a and b;
    layer1_outputs(4223) <= b;
    layer1_outputs(4224) <= a and b;
    layer1_outputs(4225) <= a xor b;
    layer1_outputs(4226) <= a and not b;
    layer1_outputs(4227) <= a or b;
    layer1_outputs(4228) <= a and b;
    layer1_outputs(4229) <= not a or b;
    layer1_outputs(4230) <= a and not b;
    layer1_outputs(4231) <= not b or a;
    layer1_outputs(4232) <= not b or a;
    layer1_outputs(4233) <= not (a and b);
    layer1_outputs(4234) <= a or b;
    layer1_outputs(4235) <= not (a xor b);
    layer1_outputs(4236) <= '1';
    layer1_outputs(4237) <= a;
    layer1_outputs(4238) <= not b or a;
    layer1_outputs(4239) <= '1';
    layer1_outputs(4240) <= a or b;
    layer1_outputs(4241) <= b and not a;
    layer1_outputs(4242) <= not b or a;
    layer1_outputs(4243) <= not (a or b);
    layer1_outputs(4244) <= not (a and b);
    layer1_outputs(4245) <= a or b;
    layer1_outputs(4246) <= '0';
    layer1_outputs(4247) <= a and b;
    layer1_outputs(4248) <= not a;
    layer1_outputs(4249) <= a and b;
    layer1_outputs(4250) <= not (a and b);
    layer1_outputs(4251) <= '1';
    layer1_outputs(4252) <= not (a or b);
    layer1_outputs(4253) <= b and not a;
    layer1_outputs(4254) <= not (a and b);
    layer1_outputs(4255) <= b and not a;
    layer1_outputs(4256) <= not a;
    layer1_outputs(4257) <= a;
    layer1_outputs(4258) <= not a;
    layer1_outputs(4259) <= a and not b;
    layer1_outputs(4260) <= b and not a;
    layer1_outputs(4261) <= a and not b;
    layer1_outputs(4262) <= a and not b;
    layer1_outputs(4263) <= a;
    layer1_outputs(4264) <= not (a and b);
    layer1_outputs(4265) <= not b;
    layer1_outputs(4266) <= b and not a;
    layer1_outputs(4267) <= a and not b;
    layer1_outputs(4268) <= a and not b;
    layer1_outputs(4269) <= b and not a;
    layer1_outputs(4270) <= a and b;
    layer1_outputs(4271) <= not a or b;
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= not a;
    layer1_outputs(4274) <= a and not b;
    layer1_outputs(4275) <= not (a and b);
    layer1_outputs(4276) <= not a;
    layer1_outputs(4277) <= a and not b;
    layer1_outputs(4278) <= a;
    layer1_outputs(4279) <= '0';
    layer1_outputs(4280) <= not b;
    layer1_outputs(4281) <= a xor b;
    layer1_outputs(4282) <= not a;
    layer1_outputs(4283) <= not b or a;
    layer1_outputs(4284) <= not b;
    layer1_outputs(4285) <= '1';
    layer1_outputs(4286) <= a and not b;
    layer1_outputs(4287) <= not b;
    layer1_outputs(4288) <= b and not a;
    layer1_outputs(4289) <= a or b;
    layer1_outputs(4290) <= '1';
    layer1_outputs(4291) <= not (a and b);
    layer1_outputs(4292) <= not a;
    layer1_outputs(4293) <= not (a xor b);
    layer1_outputs(4294) <= b;
    layer1_outputs(4295) <= b;
    layer1_outputs(4296) <= '0';
    layer1_outputs(4297) <= b;
    layer1_outputs(4298) <= '1';
    layer1_outputs(4299) <= not b;
    layer1_outputs(4300) <= not a or b;
    layer1_outputs(4301) <= not a or b;
    layer1_outputs(4302) <= not (a and b);
    layer1_outputs(4303) <= b;
    layer1_outputs(4304) <= '0';
    layer1_outputs(4305) <= b and not a;
    layer1_outputs(4306) <= not (a and b);
    layer1_outputs(4307) <= not a;
    layer1_outputs(4308) <= not a;
    layer1_outputs(4309) <= a and not b;
    layer1_outputs(4310) <= a;
    layer1_outputs(4311) <= a and not b;
    layer1_outputs(4312) <= b and not a;
    layer1_outputs(4313) <= a or b;
    layer1_outputs(4314) <= not b or a;
    layer1_outputs(4315) <= not b;
    layer1_outputs(4316) <= a and not b;
    layer1_outputs(4317) <= '0';
    layer1_outputs(4318) <= not b;
    layer1_outputs(4319) <= b and not a;
    layer1_outputs(4320) <= a;
    layer1_outputs(4321) <= not (a and b);
    layer1_outputs(4322) <= not b;
    layer1_outputs(4323) <= not a;
    layer1_outputs(4324) <= not (a and b);
    layer1_outputs(4325) <= a;
    layer1_outputs(4326) <= not b or a;
    layer1_outputs(4327) <= '1';
    layer1_outputs(4328) <= a or b;
    layer1_outputs(4329) <= not a or b;
    layer1_outputs(4330) <= b and not a;
    layer1_outputs(4331) <= '0';
    layer1_outputs(4332) <= b;
    layer1_outputs(4333) <= a and not b;
    layer1_outputs(4334) <= '1';
    layer1_outputs(4335) <= a;
    layer1_outputs(4336) <= b;
    layer1_outputs(4337) <= a xor b;
    layer1_outputs(4338) <= not (a or b);
    layer1_outputs(4339) <= '1';
    layer1_outputs(4340) <= not a;
    layer1_outputs(4341) <= not (a and b);
    layer1_outputs(4342) <= a;
    layer1_outputs(4343) <= '0';
    layer1_outputs(4344) <= not b or a;
    layer1_outputs(4345) <= b;
    layer1_outputs(4346) <= not b;
    layer1_outputs(4347) <= b;
    layer1_outputs(4348) <= not a;
    layer1_outputs(4349) <= not a or b;
    layer1_outputs(4350) <= not (a and b);
    layer1_outputs(4351) <= not (a and b);
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= not b;
    layer1_outputs(4354) <= a or b;
    layer1_outputs(4355) <= a;
    layer1_outputs(4356) <= a;
    layer1_outputs(4357) <= b;
    layer1_outputs(4358) <= a;
    layer1_outputs(4359) <= not a;
    layer1_outputs(4360) <= a;
    layer1_outputs(4361) <= a and not b;
    layer1_outputs(4362) <= a or b;
    layer1_outputs(4363) <= b;
    layer1_outputs(4364) <= not (a xor b);
    layer1_outputs(4365) <= a and b;
    layer1_outputs(4366) <= not a;
    layer1_outputs(4367) <= b;
    layer1_outputs(4368) <= not (a and b);
    layer1_outputs(4369) <= a and b;
    layer1_outputs(4370) <= '1';
    layer1_outputs(4371) <= not b;
    layer1_outputs(4372) <= not b or a;
    layer1_outputs(4373) <= not a or b;
    layer1_outputs(4374) <= not (a and b);
    layer1_outputs(4375) <= not a;
    layer1_outputs(4376) <= a or b;
    layer1_outputs(4377) <= a or b;
    layer1_outputs(4378) <= not (a xor b);
    layer1_outputs(4379) <= b;
    layer1_outputs(4380) <= b;
    layer1_outputs(4381) <= not (a or b);
    layer1_outputs(4382) <= a and b;
    layer1_outputs(4383) <= not b;
    layer1_outputs(4384) <= not b or a;
    layer1_outputs(4385) <= a or b;
    layer1_outputs(4386) <= not b;
    layer1_outputs(4387) <= not (a or b);
    layer1_outputs(4388) <= not a;
    layer1_outputs(4389) <= '0';
    layer1_outputs(4390) <= b and not a;
    layer1_outputs(4391) <= a and not b;
    layer1_outputs(4392) <= a;
    layer1_outputs(4393) <= not (a and b);
    layer1_outputs(4394) <= not (a or b);
    layer1_outputs(4395) <= b and not a;
    layer1_outputs(4396) <= a;
    layer1_outputs(4397) <= not (a or b);
    layer1_outputs(4398) <= not b;
    layer1_outputs(4399) <= not a;
    layer1_outputs(4400) <= b;
    layer1_outputs(4401) <= not a;
    layer1_outputs(4402) <= '0';
    layer1_outputs(4403) <= not b;
    layer1_outputs(4404) <= a and b;
    layer1_outputs(4405) <= not a;
    layer1_outputs(4406) <= a or b;
    layer1_outputs(4407) <= b;
    layer1_outputs(4408) <= '1';
    layer1_outputs(4409) <= not b or a;
    layer1_outputs(4410) <= a and not b;
    layer1_outputs(4411) <= '0';
    layer1_outputs(4412) <= not a or b;
    layer1_outputs(4413) <= not b or a;
    layer1_outputs(4414) <= not a;
    layer1_outputs(4415) <= b and not a;
    layer1_outputs(4416) <= b and not a;
    layer1_outputs(4417) <= b;
    layer1_outputs(4418) <= a or b;
    layer1_outputs(4419) <= b and not a;
    layer1_outputs(4420) <= not b;
    layer1_outputs(4421) <= not b;
    layer1_outputs(4422) <= b;
    layer1_outputs(4423) <= a and b;
    layer1_outputs(4424) <= not b or a;
    layer1_outputs(4425) <= not (a or b);
    layer1_outputs(4426) <= not a;
    layer1_outputs(4427) <= a xor b;
    layer1_outputs(4428) <= '0';
    layer1_outputs(4429) <= not (a and b);
    layer1_outputs(4430) <= b;
    layer1_outputs(4431) <= not a;
    layer1_outputs(4432) <= not b or a;
    layer1_outputs(4433) <= not (a or b);
    layer1_outputs(4434) <= a and not b;
    layer1_outputs(4435) <= a and b;
    layer1_outputs(4436) <= not b;
    layer1_outputs(4437) <= not (a or b);
    layer1_outputs(4438) <= a;
    layer1_outputs(4439) <= b;
    layer1_outputs(4440) <= not b or a;
    layer1_outputs(4441) <= a;
    layer1_outputs(4442) <= b;
    layer1_outputs(4443) <= b and not a;
    layer1_outputs(4444) <= a;
    layer1_outputs(4445) <= a or b;
    layer1_outputs(4446) <= not (a and b);
    layer1_outputs(4447) <= a and b;
    layer1_outputs(4448) <= not a;
    layer1_outputs(4449) <= '0';
    layer1_outputs(4450) <= a or b;
    layer1_outputs(4451) <= not (a xor b);
    layer1_outputs(4452) <= not a;
    layer1_outputs(4453) <= a;
    layer1_outputs(4454) <= a and b;
    layer1_outputs(4455) <= b;
    layer1_outputs(4456) <= '1';
    layer1_outputs(4457) <= not a;
    layer1_outputs(4458) <= a and b;
    layer1_outputs(4459) <= not (a or b);
    layer1_outputs(4460) <= b;
    layer1_outputs(4461) <= b and not a;
    layer1_outputs(4462) <= not b;
    layer1_outputs(4463) <= '0';
    layer1_outputs(4464) <= a or b;
    layer1_outputs(4465) <= not (a or b);
    layer1_outputs(4466) <= not b;
    layer1_outputs(4467) <= not (a and b);
    layer1_outputs(4468) <= b and not a;
    layer1_outputs(4469) <= not a;
    layer1_outputs(4470) <= b;
    layer1_outputs(4471) <= not (a or b);
    layer1_outputs(4472) <= a and not b;
    layer1_outputs(4473) <= not b;
    layer1_outputs(4474) <= '0';
    layer1_outputs(4475) <= not a;
    layer1_outputs(4476) <= a and b;
    layer1_outputs(4477) <= not (a and b);
    layer1_outputs(4478) <= a or b;
    layer1_outputs(4479) <= '0';
    layer1_outputs(4480) <= a and not b;
    layer1_outputs(4481) <= not (a and b);
    layer1_outputs(4482) <= b and not a;
    layer1_outputs(4483) <= '0';
    layer1_outputs(4484) <= a or b;
    layer1_outputs(4485) <= '1';
    layer1_outputs(4486) <= not b or a;
    layer1_outputs(4487) <= not a;
    layer1_outputs(4488) <= a or b;
    layer1_outputs(4489) <= a and not b;
    layer1_outputs(4490) <= a and b;
    layer1_outputs(4491) <= a and b;
    layer1_outputs(4492) <= not b;
    layer1_outputs(4493) <= '1';
    layer1_outputs(4494) <= '1';
    layer1_outputs(4495) <= not b or a;
    layer1_outputs(4496) <= b;
    layer1_outputs(4497) <= '1';
    layer1_outputs(4498) <= a and not b;
    layer1_outputs(4499) <= '0';
    layer1_outputs(4500) <= not (a or b);
    layer1_outputs(4501) <= b;
    layer1_outputs(4502) <= a;
    layer1_outputs(4503) <= not a;
    layer1_outputs(4504) <= '0';
    layer1_outputs(4505) <= not (a or b);
    layer1_outputs(4506) <= a;
    layer1_outputs(4507) <= '0';
    layer1_outputs(4508) <= not b or a;
    layer1_outputs(4509) <= a;
    layer1_outputs(4510) <= a or b;
    layer1_outputs(4511) <= a;
    layer1_outputs(4512) <= a and b;
    layer1_outputs(4513) <= not (a or b);
    layer1_outputs(4514) <= a and not b;
    layer1_outputs(4515) <= '0';
    layer1_outputs(4516) <= not a;
    layer1_outputs(4517) <= a and b;
    layer1_outputs(4518) <= a and not b;
    layer1_outputs(4519) <= a and b;
    layer1_outputs(4520) <= not (a xor b);
    layer1_outputs(4521) <= a;
    layer1_outputs(4522) <= not (a and b);
    layer1_outputs(4523) <= a and b;
    layer1_outputs(4524) <= b and not a;
    layer1_outputs(4525) <= a xor b;
    layer1_outputs(4526) <= a and b;
    layer1_outputs(4527) <= '0';
    layer1_outputs(4528) <= not a;
    layer1_outputs(4529) <= not a or b;
    layer1_outputs(4530) <= '1';
    layer1_outputs(4531) <= not b or a;
    layer1_outputs(4532) <= a xor b;
    layer1_outputs(4533) <= a;
    layer1_outputs(4534) <= not a;
    layer1_outputs(4535) <= not b;
    layer1_outputs(4536) <= a;
    layer1_outputs(4537) <= not (a or b);
    layer1_outputs(4538) <= a xor b;
    layer1_outputs(4539) <= a;
    layer1_outputs(4540) <= b and not a;
    layer1_outputs(4541) <= a xor b;
    layer1_outputs(4542) <= not a;
    layer1_outputs(4543) <= not b;
    layer1_outputs(4544) <= a and b;
    layer1_outputs(4545) <= not (a or b);
    layer1_outputs(4546) <= not (a and b);
    layer1_outputs(4547) <= not (a and b);
    layer1_outputs(4548) <= not b;
    layer1_outputs(4549) <= b;
    layer1_outputs(4550) <= '0';
    layer1_outputs(4551) <= not a or b;
    layer1_outputs(4552) <= a or b;
    layer1_outputs(4553) <= b and not a;
    layer1_outputs(4554) <= a;
    layer1_outputs(4555) <= not a;
    layer1_outputs(4556) <= not b or a;
    layer1_outputs(4557) <= not b or a;
    layer1_outputs(4558) <= a;
    layer1_outputs(4559) <= b;
    layer1_outputs(4560) <= not (a or b);
    layer1_outputs(4561) <= '1';
    layer1_outputs(4562) <= not (a and b);
    layer1_outputs(4563) <= not (a and b);
    layer1_outputs(4564) <= a and b;
    layer1_outputs(4565) <= '1';
    layer1_outputs(4566) <= a xor b;
    layer1_outputs(4567) <= not a or b;
    layer1_outputs(4568) <= not a;
    layer1_outputs(4569) <= not (a xor b);
    layer1_outputs(4570) <= a;
    layer1_outputs(4571) <= a or b;
    layer1_outputs(4572) <= b and not a;
    layer1_outputs(4573) <= b and not a;
    layer1_outputs(4574) <= not (a and b);
    layer1_outputs(4575) <= a and not b;
    layer1_outputs(4576) <= not a;
    layer1_outputs(4577) <= not a or b;
    layer1_outputs(4578) <= a;
    layer1_outputs(4579) <= not a or b;
    layer1_outputs(4580) <= not (a or b);
    layer1_outputs(4581) <= a and b;
    layer1_outputs(4582) <= a and not b;
    layer1_outputs(4583) <= a xor b;
    layer1_outputs(4584) <= '1';
    layer1_outputs(4585) <= b;
    layer1_outputs(4586) <= '1';
    layer1_outputs(4587) <= a xor b;
    layer1_outputs(4588) <= not (a or b);
    layer1_outputs(4589) <= not a;
    layer1_outputs(4590) <= not a or b;
    layer1_outputs(4591) <= '0';
    layer1_outputs(4592) <= not a;
    layer1_outputs(4593) <= a xor b;
    layer1_outputs(4594) <= not a or b;
    layer1_outputs(4595) <= a xor b;
    layer1_outputs(4596) <= not b or a;
    layer1_outputs(4597) <= not (a xor b);
    layer1_outputs(4598) <= not a or b;
    layer1_outputs(4599) <= not (a or b);
    layer1_outputs(4600) <= b and not a;
    layer1_outputs(4601) <= not b;
    layer1_outputs(4602) <= '1';
    layer1_outputs(4603) <= '1';
    layer1_outputs(4604) <= b;
    layer1_outputs(4605) <= a;
    layer1_outputs(4606) <= not a or b;
    layer1_outputs(4607) <= a;
    layer1_outputs(4608) <= a and not b;
    layer1_outputs(4609) <= a or b;
    layer1_outputs(4610) <= a;
    layer1_outputs(4611) <= a or b;
    layer1_outputs(4612) <= not (a and b);
    layer1_outputs(4613) <= a;
    layer1_outputs(4614) <= not a;
    layer1_outputs(4615) <= a and b;
    layer1_outputs(4616) <= not a;
    layer1_outputs(4617) <= not b;
    layer1_outputs(4618) <= a;
    layer1_outputs(4619) <= a;
    layer1_outputs(4620) <= a;
    layer1_outputs(4621) <= a and b;
    layer1_outputs(4622) <= not b;
    layer1_outputs(4623) <= '1';
    layer1_outputs(4624) <= a or b;
    layer1_outputs(4625) <= not a or b;
    layer1_outputs(4626) <= a;
    layer1_outputs(4627) <= not (a or b);
    layer1_outputs(4628) <= not a;
    layer1_outputs(4629) <= a;
    layer1_outputs(4630) <= a;
    layer1_outputs(4631) <= b;
    layer1_outputs(4632) <= '0';
    layer1_outputs(4633) <= a and b;
    layer1_outputs(4634) <= not a;
    layer1_outputs(4635) <= not b;
    layer1_outputs(4636) <= b;
    layer1_outputs(4637) <= not a or b;
    layer1_outputs(4638) <= a;
    layer1_outputs(4639) <= a and not b;
    layer1_outputs(4640) <= b and not a;
    layer1_outputs(4641) <= not (a or b);
    layer1_outputs(4642) <= a and not b;
    layer1_outputs(4643) <= not b;
    layer1_outputs(4644) <= a and b;
    layer1_outputs(4645) <= a and b;
    layer1_outputs(4646) <= not (a and b);
    layer1_outputs(4647) <= '0';
    layer1_outputs(4648) <= not a;
    layer1_outputs(4649) <= not a or b;
    layer1_outputs(4650) <= b;
    layer1_outputs(4651) <= b;
    layer1_outputs(4652) <= '1';
    layer1_outputs(4653) <= a;
    layer1_outputs(4654) <= not b or a;
    layer1_outputs(4655) <= a and not b;
    layer1_outputs(4656) <= not (a and b);
    layer1_outputs(4657) <= b;
    layer1_outputs(4658) <= a;
    layer1_outputs(4659) <= '1';
    layer1_outputs(4660) <= a or b;
    layer1_outputs(4661) <= not a or b;
    layer1_outputs(4662) <= not b or a;
    layer1_outputs(4663) <= a or b;
    layer1_outputs(4664) <= '1';
    layer1_outputs(4665) <= a and not b;
    layer1_outputs(4666) <= not b;
    layer1_outputs(4667) <= a and not b;
    layer1_outputs(4668) <= '0';
    layer1_outputs(4669) <= '1';
    layer1_outputs(4670) <= not a or b;
    layer1_outputs(4671) <= not b;
    layer1_outputs(4672) <= not (a or b);
    layer1_outputs(4673) <= '0';
    layer1_outputs(4674) <= b;
    layer1_outputs(4675) <= not a or b;
    layer1_outputs(4676) <= a;
    layer1_outputs(4677) <= a or b;
    layer1_outputs(4678) <= not b;
    layer1_outputs(4679) <= not b;
    layer1_outputs(4680) <= b;
    layer1_outputs(4681) <= not (a and b);
    layer1_outputs(4682) <= not b or a;
    layer1_outputs(4683) <= not b or a;
    layer1_outputs(4684) <= a and b;
    layer1_outputs(4685) <= '1';
    layer1_outputs(4686) <= not b;
    layer1_outputs(4687) <= '0';
    layer1_outputs(4688) <= a and not b;
    layer1_outputs(4689) <= b;
    layer1_outputs(4690) <= b;
    layer1_outputs(4691) <= '0';
    layer1_outputs(4692) <= not b;
    layer1_outputs(4693) <= a;
    layer1_outputs(4694) <= a and not b;
    layer1_outputs(4695) <= not a or b;
    layer1_outputs(4696) <= not (a and b);
    layer1_outputs(4697) <= not (a and b);
    layer1_outputs(4698) <= not (a or b);
    layer1_outputs(4699) <= not b;
    layer1_outputs(4700) <= not (a or b);
    layer1_outputs(4701) <= a or b;
    layer1_outputs(4702) <= b and not a;
    layer1_outputs(4703) <= not a or b;
    layer1_outputs(4704) <= b and not a;
    layer1_outputs(4705) <= '1';
    layer1_outputs(4706) <= b;
    layer1_outputs(4707) <= a;
    layer1_outputs(4708) <= '0';
    layer1_outputs(4709) <= not (a and b);
    layer1_outputs(4710) <= not b;
    layer1_outputs(4711) <= not a or b;
    layer1_outputs(4712) <= '1';
    layer1_outputs(4713) <= a;
    layer1_outputs(4714) <= not a;
    layer1_outputs(4715) <= not (a or b);
    layer1_outputs(4716) <= '0';
    layer1_outputs(4717) <= a xor b;
    layer1_outputs(4718) <= b and not a;
    layer1_outputs(4719) <= not b;
    layer1_outputs(4720) <= a;
    layer1_outputs(4721) <= a;
    layer1_outputs(4722) <= b;
    layer1_outputs(4723) <= a and not b;
    layer1_outputs(4724) <= not a or b;
    layer1_outputs(4725) <= not (a or b);
    layer1_outputs(4726) <= b;
    layer1_outputs(4727) <= a and not b;
    layer1_outputs(4728) <= a or b;
    layer1_outputs(4729) <= not (a xor b);
    layer1_outputs(4730) <= '1';
    layer1_outputs(4731) <= not (a or b);
    layer1_outputs(4732) <= a and b;
    layer1_outputs(4733) <= not (a or b);
    layer1_outputs(4734) <= b;
    layer1_outputs(4735) <= a and not b;
    layer1_outputs(4736) <= a or b;
    layer1_outputs(4737) <= a and not b;
    layer1_outputs(4738) <= not (a and b);
    layer1_outputs(4739) <= a and not b;
    layer1_outputs(4740) <= b;
    layer1_outputs(4741) <= not b;
    layer1_outputs(4742) <= not (a or b);
    layer1_outputs(4743) <= a or b;
    layer1_outputs(4744) <= not (a or b);
    layer1_outputs(4745) <= a and b;
    layer1_outputs(4746) <= '0';
    layer1_outputs(4747) <= not b;
    layer1_outputs(4748) <= a;
    layer1_outputs(4749) <= not a or b;
    layer1_outputs(4750) <= not a;
    layer1_outputs(4751) <= a and not b;
    layer1_outputs(4752) <= '0';
    layer1_outputs(4753) <= a and b;
    layer1_outputs(4754) <= '0';
    layer1_outputs(4755) <= a or b;
    layer1_outputs(4756) <= not a;
    layer1_outputs(4757) <= not (a or b);
    layer1_outputs(4758) <= a xor b;
    layer1_outputs(4759) <= not a or b;
    layer1_outputs(4760) <= not b or a;
    layer1_outputs(4761) <= not (a xor b);
    layer1_outputs(4762) <= '0';
    layer1_outputs(4763) <= a and not b;
    layer1_outputs(4764) <= not (a and b);
    layer1_outputs(4765) <= not a;
    layer1_outputs(4766) <= not b or a;
    layer1_outputs(4767) <= a and b;
    layer1_outputs(4768) <= not b;
    layer1_outputs(4769) <= not a;
    layer1_outputs(4770) <= '0';
    layer1_outputs(4771) <= not (a and b);
    layer1_outputs(4772) <= not b;
    layer1_outputs(4773) <= not a;
    layer1_outputs(4774) <= not a;
    layer1_outputs(4775) <= a;
    layer1_outputs(4776) <= b and not a;
    layer1_outputs(4777) <= b;
    layer1_outputs(4778) <= not (a and b);
    layer1_outputs(4779) <= not b;
    layer1_outputs(4780) <= not a;
    layer1_outputs(4781) <= a and b;
    layer1_outputs(4782) <= a and not b;
    layer1_outputs(4783) <= a;
    layer1_outputs(4784) <= '1';
    layer1_outputs(4785) <= b and not a;
    layer1_outputs(4786) <= not b;
    layer1_outputs(4787) <= not (a or b);
    layer1_outputs(4788) <= not b or a;
    layer1_outputs(4789) <= a and not b;
    layer1_outputs(4790) <= a and b;
    layer1_outputs(4791) <= not a or b;
    layer1_outputs(4792) <= a;
    layer1_outputs(4793) <= not a;
    layer1_outputs(4794) <= a and b;
    layer1_outputs(4795) <= b;
    layer1_outputs(4796) <= a and b;
    layer1_outputs(4797) <= a or b;
    layer1_outputs(4798) <= not a or b;
    layer1_outputs(4799) <= a xor b;
    layer1_outputs(4800) <= b;
    layer1_outputs(4801) <= a and b;
    layer1_outputs(4802) <= not a;
    layer1_outputs(4803) <= not (a or b);
    layer1_outputs(4804) <= a;
    layer1_outputs(4805) <= '1';
    layer1_outputs(4806) <= not a;
    layer1_outputs(4807) <= b;
    layer1_outputs(4808) <= '1';
    layer1_outputs(4809) <= a or b;
    layer1_outputs(4810) <= a and not b;
    layer1_outputs(4811) <= not a or b;
    layer1_outputs(4812) <= not b;
    layer1_outputs(4813) <= not a or b;
    layer1_outputs(4814) <= b and not a;
    layer1_outputs(4815) <= not b or a;
    layer1_outputs(4816) <= a and b;
    layer1_outputs(4817) <= a;
    layer1_outputs(4818) <= a or b;
    layer1_outputs(4819) <= not a;
    layer1_outputs(4820) <= a or b;
    layer1_outputs(4821) <= not b;
    layer1_outputs(4822) <= a or b;
    layer1_outputs(4823) <= not (a and b);
    layer1_outputs(4824) <= not b;
    layer1_outputs(4825) <= not (a and b);
    layer1_outputs(4826) <= a;
    layer1_outputs(4827) <= b;
    layer1_outputs(4828) <= a and b;
    layer1_outputs(4829) <= not (a xor b);
    layer1_outputs(4830) <= '0';
    layer1_outputs(4831) <= a and b;
    layer1_outputs(4832) <= a xor b;
    layer1_outputs(4833) <= not a;
    layer1_outputs(4834) <= not a or b;
    layer1_outputs(4835) <= not (a and b);
    layer1_outputs(4836) <= not b;
    layer1_outputs(4837) <= a and not b;
    layer1_outputs(4838) <= a;
    layer1_outputs(4839) <= '0';
    layer1_outputs(4840) <= b and not a;
    layer1_outputs(4841) <= a;
    layer1_outputs(4842) <= not (a or b);
    layer1_outputs(4843) <= a and b;
    layer1_outputs(4844) <= not b;
    layer1_outputs(4845) <= b;
    layer1_outputs(4846) <= a;
    layer1_outputs(4847) <= a and b;
    layer1_outputs(4848) <= b and not a;
    layer1_outputs(4849) <= a;
    layer1_outputs(4850) <= a and b;
    layer1_outputs(4851) <= a;
    layer1_outputs(4852) <= a;
    layer1_outputs(4853) <= b and not a;
    layer1_outputs(4854) <= b;
    layer1_outputs(4855) <= not (a or b);
    layer1_outputs(4856) <= not b;
    layer1_outputs(4857) <= not a or b;
    layer1_outputs(4858) <= a xor b;
    layer1_outputs(4859) <= b;
    layer1_outputs(4860) <= not b;
    layer1_outputs(4861) <= not (a or b);
    layer1_outputs(4862) <= not b;
    layer1_outputs(4863) <= not (a and b);
    layer1_outputs(4864) <= '1';
    layer1_outputs(4865) <= '1';
    layer1_outputs(4866) <= a;
    layer1_outputs(4867) <= b and not a;
    layer1_outputs(4868) <= not b;
    layer1_outputs(4869) <= not b or a;
    layer1_outputs(4870) <= a or b;
    layer1_outputs(4871) <= b;
    layer1_outputs(4872) <= not b or a;
    layer1_outputs(4873) <= b;
    layer1_outputs(4874) <= b;
    layer1_outputs(4875) <= b;
    layer1_outputs(4876) <= b;
    layer1_outputs(4877) <= '0';
    layer1_outputs(4878) <= not (a and b);
    layer1_outputs(4879) <= b;
    layer1_outputs(4880) <= not a;
    layer1_outputs(4881) <= not a;
    layer1_outputs(4882) <= a xor b;
    layer1_outputs(4883) <= not a;
    layer1_outputs(4884) <= not (a xor b);
    layer1_outputs(4885) <= a and not b;
    layer1_outputs(4886) <= not (a or b);
    layer1_outputs(4887) <= a or b;
    layer1_outputs(4888) <= '1';
    layer1_outputs(4889) <= not (a or b);
    layer1_outputs(4890) <= a or b;
    layer1_outputs(4891) <= not b or a;
    layer1_outputs(4892) <= not a;
    layer1_outputs(4893) <= b;
    layer1_outputs(4894) <= not a;
    layer1_outputs(4895) <= not a;
    layer1_outputs(4896) <= not b;
    layer1_outputs(4897) <= not (a or b);
    layer1_outputs(4898) <= b and not a;
    layer1_outputs(4899) <= a;
    layer1_outputs(4900) <= '1';
    layer1_outputs(4901) <= not (a or b);
    layer1_outputs(4902) <= not a;
    layer1_outputs(4903) <= a and b;
    layer1_outputs(4904) <= not b or a;
    layer1_outputs(4905) <= a;
    layer1_outputs(4906) <= b and not a;
    layer1_outputs(4907) <= not a or b;
    layer1_outputs(4908) <= not b;
    layer1_outputs(4909) <= b;
    layer1_outputs(4910) <= a;
    layer1_outputs(4911) <= not a;
    layer1_outputs(4912) <= not b;
    layer1_outputs(4913) <= a;
    layer1_outputs(4914) <= b;
    layer1_outputs(4915) <= a or b;
    layer1_outputs(4916) <= not a;
    layer1_outputs(4917) <= not b or a;
    layer1_outputs(4918) <= not a;
    layer1_outputs(4919) <= a;
    layer1_outputs(4920) <= not (a and b);
    layer1_outputs(4921) <= not (a or b);
    layer1_outputs(4922) <= not a or b;
    layer1_outputs(4923) <= b;
    layer1_outputs(4924) <= not b or a;
    layer1_outputs(4925) <= a or b;
    layer1_outputs(4926) <= a and not b;
    layer1_outputs(4927) <= a and b;
    layer1_outputs(4928) <= a;
    layer1_outputs(4929) <= '0';
    layer1_outputs(4930) <= '0';
    layer1_outputs(4931) <= a;
    layer1_outputs(4932) <= not (a or b);
    layer1_outputs(4933) <= b and not a;
    layer1_outputs(4934) <= not (a xor b);
    layer1_outputs(4935) <= b;
    layer1_outputs(4936) <= not b or a;
    layer1_outputs(4937) <= not a or b;
    layer1_outputs(4938) <= not a;
    layer1_outputs(4939) <= not (a and b);
    layer1_outputs(4940) <= not a or b;
    layer1_outputs(4941) <= not a or b;
    layer1_outputs(4942) <= '1';
    layer1_outputs(4943) <= a and not b;
    layer1_outputs(4944) <= not (a or b);
    layer1_outputs(4945) <= a and not b;
    layer1_outputs(4946) <= a xor b;
    layer1_outputs(4947) <= not b;
    layer1_outputs(4948) <= not (a and b);
    layer1_outputs(4949) <= not (a xor b);
    layer1_outputs(4950) <= not (a and b);
    layer1_outputs(4951) <= '1';
    layer1_outputs(4952) <= not (a xor b);
    layer1_outputs(4953) <= not (a xor b);
    layer1_outputs(4954) <= a;
    layer1_outputs(4955) <= not b;
    layer1_outputs(4956) <= '0';
    layer1_outputs(4957) <= a and b;
    layer1_outputs(4958) <= not (a or b);
    layer1_outputs(4959) <= a and not b;
    layer1_outputs(4960) <= b and not a;
    layer1_outputs(4961) <= not a;
    layer1_outputs(4962) <= b;
    layer1_outputs(4963) <= not (a or b);
    layer1_outputs(4964) <= '0';
    layer1_outputs(4965) <= b;
    layer1_outputs(4966) <= not (a xor b);
    layer1_outputs(4967) <= not b or a;
    layer1_outputs(4968) <= a;
    layer1_outputs(4969) <= not b or a;
    layer1_outputs(4970) <= not a;
    layer1_outputs(4971) <= '0';
    layer1_outputs(4972) <= a;
    layer1_outputs(4973) <= not a;
    layer1_outputs(4974) <= not a or b;
    layer1_outputs(4975) <= '1';
    layer1_outputs(4976) <= not (a or b);
    layer1_outputs(4977) <= a and b;
    layer1_outputs(4978) <= not b;
    layer1_outputs(4979) <= '0';
    layer1_outputs(4980) <= not b or a;
    layer1_outputs(4981) <= a and not b;
    layer1_outputs(4982) <= not (a xor b);
    layer1_outputs(4983) <= not (a or b);
    layer1_outputs(4984) <= a and not b;
    layer1_outputs(4985) <= a;
    layer1_outputs(4986) <= not (a xor b);
    layer1_outputs(4987) <= b;
    layer1_outputs(4988) <= not a;
    layer1_outputs(4989) <= b;
    layer1_outputs(4990) <= b;
    layer1_outputs(4991) <= '0';
    layer1_outputs(4992) <= a and not b;
    layer1_outputs(4993) <= not b;
    layer1_outputs(4994) <= not (a xor b);
    layer1_outputs(4995) <= b;
    layer1_outputs(4996) <= a and b;
    layer1_outputs(4997) <= not (a xor b);
    layer1_outputs(4998) <= b;
    layer1_outputs(4999) <= not (a or b);
    layer1_outputs(5000) <= not (a or b);
    layer1_outputs(5001) <= a or b;
    layer1_outputs(5002) <= not a or b;
    layer1_outputs(5003) <= not a;
    layer1_outputs(5004) <= b;
    layer1_outputs(5005) <= a and not b;
    layer1_outputs(5006) <= b and not a;
    layer1_outputs(5007) <= a and not b;
    layer1_outputs(5008) <= not a or b;
    layer1_outputs(5009) <= '1';
    layer1_outputs(5010) <= a xor b;
    layer1_outputs(5011) <= not b or a;
    layer1_outputs(5012) <= not (a or b);
    layer1_outputs(5013) <= a and not b;
    layer1_outputs(5014) <= b;
    layer1_outputs(5015) <= not a;
    layer1_outputs(5016) <= not (a and b);
    layer1_outputs(5017) <= '1';
    layer1_outputs(5018) <= b and not a;
    layer1_outputs(5019) <= not (a and b);
    layer1_outputs(5020) <= a or b;
    layer1_outputs(5021) <= not (a xor b);
    layer1_outputs(5022) <= not a;
    layer1_outputs(5023) <= not (a or b);
    layer1_outputs(5024) <= b;
    layer1_outputs(5025) <= '0';
    layer1_outputs(5026) <= not b or a;
    layer1_outputs(5027) <= not b;
    layer1_outputs(5028) <= b;
    layer1_outputs(5029) <= a and b;
    layer1_outputs(5030) <= a;
    layer1_outputs(5031) <= not b;
    layer1_outputs(5032) <= b;
    layer1_outputs(5033) <= b;
    layer1_outputs(5034) <= b and not a;
    layer1_outputs(5035) <= not b or a;
    layer1_outputs(5036) <= b and not a;
    layer1_outputs(5037) <= not b;
    layer1_outputs(5038) <= a;
    layer1_outputs(5039) <= a or b;
    layer1_outputs(5040) <= a and b;
    layer1_outputs(5041) <= not b;
    layer1_outputs(5042) <= not b;
    layer1_outputs(5043) <= a;
    layer1_outputs(5044) <= not (a xor b);
    layer1_outputs(5045) <= '1';
    layer1_outputs(5046) <= b and not a;
    layer1_outputs(5047) <= not a;
    layer1_outputs(5048) <= not a or b;
    layer1_outputs(5049) <= not a;
    layer1_outputs(5050) <= a;
    layer1_outputs(5051) <= b and not a;
    layer1_outputs(5052) <= not b;
    layer1_outputs(5053) <= b and not a;
    layer1_outputs(5054) <= not a or b;
    layer1_outputs(5055) <= a and b;
    layer1_outputs(5056) <= not a;
    layer1_outputs(5057) <= not b or a;
    layer1_outputs(5058) <= a or b;
    layer1_outputs(5059) <= a and b;
    layer1_outputs(5060) <= a;
    layer1_outputs(5061) <= '1';
    layer1_outputs(5062) <= not (a and b);
    layer1_outputs(5063) <= '1';
    layer1_outputs(5064) <= b;
    layer1_outputs(5065) <= b;
    layer1_outputs(5066) <= a;
    layer1_outputs(5067) <= not a or b;
    layer1_outputs(5068) <= a;
    layer1_outputs(5069) <= a and b;
    layer1_outputs(5070) <= '0';
    layer1_outputs(5071) <= a or b;
    layer1_outputs(5072) <= b and not a;
    layer1_outputs(5073) <= b and not a;
    layer1_outputs(5074) <= not (a or b);
    layer1_outputs(5075) <= '1';
    layer1_outputs(5076) <= a and b;
    layer1_outputs(5077) <= '0';
    layer1_outputs(5078) <= not (a or b);
    layer1_outputs(5079) <= b;
    layer1_outputs(5080) <= not a;
    layer1_outputs(5081) <= a or b;
    layer1_outputs(5082) <= not a;
    layer1_outputs(5083) <= '0';
    layer1_outputs(5084) <= a;
    layer1_outputs(5085) <= '1';
    layer1_outputs(5086) <= a and not b;
    layer1_outputs(5087) <= not b;
    layer1_outputs(5088) <= b and not a;
    layer1_outputs(5089) <= not (a and b);
    layer1_outputs(5090) <= b and not a;
    layer1_outputs(5091) <= a and b;
    layer1_outputs(5092) <= '1';
    layer1_outputs(5093) <= '0';
    layer1_outputs(5094) <= not (a xor b);
    layer1_outputs(5095) <= not a;
    layer1_outputs(5096) <= not (a or b);
    layer1_outputs(5097) <= b;
    layer1_outputs(5098) <= not b;
    layer1_outputs(5099) <= '1';
    layer1_outputs(5100) <= a xor b;
    layer1_outputs(5101) <= a and not b;
    layer1_outputs(5102) <= not a;
    layer1_outputs(5103) <= '0';
    layer1_outputs(5104) <= a;
    layer1_outputs(5105) <= a or b;
    layer1_outputs(5106) <= not (a and b);
    layer1_outputs(5107) <= not b or a;
    layer1_outputs(5108) <= not (a and b);
    layer1_outputs(5109) <= b;
    layer1_outputs(5110) <= '0';
    layer1_outputs(5111) <= not a or b;
    layer1_outputs(5112) <= a xor b;
    layer1_outputs(5113) <= b;
    layer1_outputs(5114) <= not (a or b);
    layer1_outputs(5115) <= a and not b;
    layer1_outputs(5116) <= not (a xor b);
    layer1_outputs(5117) <= not a;
    layer1_outputs(5118) <= b;
    layer1_outputs(5119) <= not b or a;
    layer1_outputs(5120) <= a xor b;
    layer1_outputs(5121) <= not a;
    layer1_outputs(5122) <= '1';
    layer1_outputs(5123) <= a or b;
    layer1_outputs(5124) <= not (a or b);
    layer1_outputs(5125) <= a or b;
    layer1_outputs(5126) <= not (a or b);
    layer1_outputs(5127) <= not a or b;
    layer1_outputs(5128) <= a;
    layer1_outputs(5129) <= not (a xor b);
    layer1_outputs(5130) <= b and not a;
    layer1_outputs(5131) <= '0';
    layer1_outputs(5132) <= not (a or b);
    layer1_outputs(5133) <= b;
    layer1_outputs(5134) <= not b or a;
    layer1_outputs(5135) <= '0';
    layer1_outputs(5136) <= a and not b;
    layer1_outputs(5137) <= not (a and b);
    layer1_outputs(5138) <= not a;
    layer1_outputs(5139) <= b;
    layer1_outputs(5140) <= a xor b;
    layer1_outputs(5141) <= not (a and b);
    layer1_outputs(5142) <= not (a and b);
    layer1_outputs(5143) <= '1';
    layer1_outputs(5144) <= not a or b;
    layer1_outputs(5145) <= a or b;
    layer1_outputs(5146) <= a;
    layer1_outputs(5147) <= not b;
    layer1_outputs(5148) <= '1';
    layer1_outputs(5149) <= '1';
    layer1_outputs(5150) <= not (a xor b);
    layer1_outputs(5151) <= not b;
    layer1_outputs(5152) <= not a;
    layer1_outputs(5153) <= a;
    layer1_outputs(5154) <= not a;
    layer1_outputs(5155) <= a or b;
    layer1_outputs(5156) <= a;
    layer1_outputs(5157) <= a;
    layer1_outputs(5158) <= a;
    layer1_outputs(5159) <= not a;
    layer1_outputs(5160) <= not a;
    layer1_outputs(5161) <= a xor b;
    layer1_outputs(5162) <= '0';
    layer1_outputs(5163) <= a;
    layer1_outputs(5164) <= not a or b;
    layer1_outputs(5165) <= a and b;
    layer1_outputs(5166) <= not (a or b);
    layer1_outputs(5167) <= not (a or b);
    layer1_outputs(5168) <= not a;
    layer1_outputs(5169) <= a;
    layer1_outputs(5170) <= b and not a;
    layer1_outputs(5171) <= not b or a;
    layer1_outputs(5172) <= a;
    layer1_outputs(5173) <= not a or b;
    layer1_outputs(5174) <= a and b;
    layer1_outputs(5175) <= '0';
    layer1_outputs(5176) <= a;
    layer1_outputs(5177) <= b;
    layer1_outputs(5178) <= a;
    layer1_outputs(5179) <= a and b;
    layer1_outputs(5180) <= '1';
    layer1_outputs(5181) <= not b;
    layer1_outputs(5182) <= not (a xor b);
    layer1_outputs(5183) <= not a or b;
    layer1_outputs(5184) <= not (a xor b);
    layer1_outputs(5185) <= not a or b;
    layer1_outputs(5186) <= a and b;
    layer1_outputs(5187) <= not b or a;
    layer1_outputs(5188) <= '1';
    layer1_outputs(5189) <= not b or a;
    layer1_outputs(5190) <= b and not a;
    layer1_outputs(5191) <= a and b;
    layer1_outputs(5192) <= a and not b;
    layer1_outputs(5193) <= not b;
    layer1_outputs(5194) <= not (a and b);
    layer1_outputs(5195) <= a and b;
    layer1_outputs(5196) <= '0';
    layer1_outputs(5197) <= not (a or b);
    layer1_outputs(5198) <= not (a and b);
    layer1_outputs(5199) <= b;
    layer1_outputs(5200) <= '1';
    layer1_outputs(5201) <= not (a and b);
    layer1_outputs(5202) <= not (a or b);
    layer1_outputs(5203) <= a and not b;
    layer1_outputs(5204) <= a;
    layer1_outputs(5205) <= not a or b;
    layer1_outputs(5206) <= a or b;
    layer1_outputs(5207) <= not (a and b);
    layer1_outputs(5208) <= not (a xor b);
    layer1_outputs(5209) <= a and b;
    layer1_outputs(5210) <= '0';
    layer1_outputs(5211) <= not (a xor b);
    layer1_outputs(5212) <= b and not a;
    layer1_outputs(5213) <= a;
    layer1_outputs(5214) <= not a;
    layer1_outputs(5215) <= b;
    layer1_outputs(5216) <= '0';
    layer1_outputs(5217) <= '0';
    layer1_outputs(5218) <= b;
    layer1_outputs(5219) <= b and not a;
    layer1_outputs(5220) <= not a;
    layer1_outputs(5221) <= '1';
    layer1_outputs(5222) <= not (a and b);
    layer1_outputs(5223) <= a;
    layer1_outputs(5224) <= a and not b;
    layer1_outputs(5225) <= '0';
    layer1_outputs(5226) <= '0';
    layer1_outputs(5227) <= not (a and b);
    layer1_outputs(5228) <= not (a and b);
    layer1_outputs(5229) <= b;
    layer1_outputs(5230) <= not (a or b);
    layer1_outputs(5231) <= a or b;
    layer1_outputs(5232) <= b;
    layer1_outputs(5233) <= not (a or b);
    layer1_outputs(5234) <= not b;
    layer1_outputs(5235) <= not a or b;
    layer1_outputs(5236) <= not a;
    layer1_outputs(5237) <= not a;
    layer1_outputs(5238) <= b;
    layer1_outputs(5239) <= '1';
    layer1_outputs(5240) <= not b or a;
    layer1_outputs(5241) <= not a;
    layer1_outputs(5242) <= not a;
    layer1_outputs(5243) <= a and not b;
    layer1_outputs(5244) <= '1';
    layer1_outputs(5245) <= not (a or b);
    layer1_outputs(5246) <= not (a and b);
    layer1_outputs(5247) <= not (a or b);
    layer1_outputs(5248) <= not a;
    layer1_outputs(5249) <= a or b;
    layer1_outputs(5250) <= '0';
    layer1_outputs(5251) <= a;
    layer1_outputs(5252) <= a;
    layer1_outputs(5253) <= a or b;
    layer1_outputs(5254) <= a and b;
    layer1_outputs(5255) <= a or b;
    layer1_outputs(5256) <= not (a or b);
    layer1_outputs(5257) <= a or b;
    layer1_outputs(5258) <= not b or a;
    layer1_outputs(5259) <= not (a or b);
    layer1_outputs(5260) <= not a or b;
    layer1_outputs(5261) <= not (a or b);
    layer1_outputs(5262) <= b and not a;
    layer1_outputs(5263) <= b and not a;
    layer1_outputs(5264) <= b;
    layer1_outputs(5265) <= not (a or b);
    layer1_outputs(5266) <= '1';
    layer1_outputs(5267) <= b and not a;
    layer1_outputs(5268) <= a and not b;
    layer1_outputs(5269) <= a;
    layer1_outputs(5270) <= a;
    layer1_outputs(5271) <= b;
    layer1_outputs(5272) <= '0';
    layer1_outputs(5273) <= a and b;
    layer1_outputs(5274) <= a and not b;
    layer1_outputs(5275) <= not (a and b);
    layer1_outputs(5276) <= not b;
    layer1_outputs(5277) <= '1';
    layer1_outputs(5278) <= not b;
    layer1_outputs(5279) <= not (a xor b);
    layer1_outputs(5280) <= not (a or b);
    layer1_outputs(5281) <= not a or b;
    layer1_outputs(5282) <= not (a or b);
    layer1_outputs(5283) <= not a;
    layer1_outputs(5284) <= not b or a;
    layer1_outputs(5285) <= b and not a;
    layer1_outputs(5286) <= a and not b;
    layer1_outputs(5287) <= not a;
    layer1_outputs(5288) <= not (a or b);
    layer1_outputs(5289) <= not b;
    layer1_outputs(5290) <= a;
    layer1_outputs(5291) <= a xor b;
    layer1_outputs(5292) <= a and b;
    layer1_outputs(5293) <= b and not a;
    layer1_outputs(5294) <= not a;
    layer1_outputs(5295) <= a xor b;
    layer1_outputs(5296) <= '1';
    layer1_outputs(5297) <= a;
    layer1_outputs(5298) <= not a or b;
    layer1_outputs(5299) <= not a;
    layer1_outputs(5300) <= a xor b;
    layer1_outputs(5301) <= b and not a;
    layer1_outputs(5302) <= not a or b;
    layer1_outputs(5303) <= a;
    layer1_outputs(5304) <= a and not b;
    layer1_outputs(5305) <= a or b;
    layer1_outputs(5306) <= a and b;
    layer1_outputs(5307) <= a and not b;
    layer1_outputs(5308) <= not a or b;
    layer1_outputs(5309) <= not b;
    layer1_outputs(5310) <= a xor b;
    layer1_outputs(5311) <= a or b;
    layer1_outputs(5312) <= not b;
    layer1_outputs(5313) <= '0';
    layer1_outputs(5314) <= b;
    layer1_outputs(5315) <= not b;
    layer1_outputs(5316) <= b and not a;
    layer1_outputs(5317) <= not a;
    layer1_outputs(5318) <= a and not b;
    layer1_outputs(5319) <= b;
    layer1_outputs(5320) <= a and not b;
    layer1_outputs(5321) <= b;
    layer1_outputs(5322) <= not b or a;
    layer1_outputs(5323) <= '1';
    layer1_outputs(5324) <= not (a xor b);
    layer1_outputs(5325) <= '0';
    layer1_outputs(5326) <= a and not b;
    layer1_outputs(5327) <= '1';
    layer1_outputs(5328) <= a and b;
    layer1_outputs(5329) <= b;
    layer1_outputs(5330) <= a or b;
    layer1_outputs(5331) <= '0';
    layer1_outputs(5332) <= not a;
    layer1_outputs(5333) <= not (a or b);
    layer1_outputs(5334) <= b and not a;
    layer1_outputs(5335) <= a or b;
    layer1_outputs(5336) <= a or b;
    layer1_outputs(5337) <= not b or a;
    layer1_outputs(5338) <= not a or b;
    layer1_outputs(5339) <= not (a or b);
    layer1_outputs(5340) <= a or b;
    layer1_outputs(5341) <= '0';
    layer1_outputs(5342) <= a;
    layer1_outputs(5343) <= not a or b;
    layer1_outputs(5344) <= not b;
    layer1_outputs(5345) <= '1';
    layer1_outputs(5346) <= a;
    layer1_outputs(5347) <= not a or b;
    layer1_outputs(5348) <= not a;
    layer1_outputs(5349) <= a or b;
    layer1_outputs(5350) <= a;
    layer1_outputs(5351) <= not (a xor b);
    layer1_outputs(5352) <= not b;
    layer1_outputs(5353) <= not (a and b);
    layer1_outputs(5354) <= '0';
    layer1_outputs(5355) <= '1';
    layer1_outputs(5356) <= not b or a;
    layer1_outputs(5357) <= a and b;
    layer1_outputs(5358) <= b and not a;
    layer1_outputs(5359) <= a;
    layer1_outputs(5360) <= not (a and b);
    layer1_outputs(5361) <= not (a or b);
    layer1_outputs(5362) <= a;
    layer1_outputs(5363) <= not (a and b);
    layer1_outputs(5364) <= not a or b;
    layer1_outputs(5365) <= not b or a;
    layer1_outputs(5366) <= b and not a;
    layer1_outputs(5367) <= not b;
    layer1_outputs(5368) <= not (a or b);
    layer1_outputs(5369) <= not a;
    layer1_outputs(5370) <= b;
    layer1_outputs(5371) <= not b or a;
    layer1_outputs(5372) <= not b;
    layer1_outputs(5373) <= not (a xor b);
    layer1_outputs(5374) <= '0';
    layer1_outputs(5375) <= b;
    layer1_outputs(5376) <= b and not a;
    layer1_outputs(5377) <= not a;
    layer1_outputs(5378) <= not (a and b);
    layer1_outputs(5379) <= not a or b;
    layer1_outputs(5380) <= a and not b;
    layer1_outputs(5381) <= a;
    layer1_outputs(5382) <= a xor b;
    layer1_outputs(5383) <= '0';
    layer1_outputs(5384) <= not (a and b);
    layer1_outputs(5385) <= not (a xor b);
    layer1_outputs(5386) <= a or b;
    layer1_outputs(5387) <= not (a xor b);
    layer1_outputs(5388) <= not b or a;
    layer1_outputs(5389) <= not (a and b);
    layer1_outputs(5390) <= b;
    layer1_outputs(5391) <= '0';
    layer1_outputs(5392) <= not (a or b);
    layer1_outputs(5393) <= b;
    layer1_outputs(5394) <= a or b;
    layer1_outputs(5395) <= not b;
    layer1_outputs(5396) <= not a or b;
    layer1_outputs(5397) <= not a or b;
    layer1_outputs(5398) <= '0';
    layer1_outputs(5399) <= b and not a;
    layer1_outputs(5400) <= not b;
    layer1_outputs(5401) <= not a or b;
    layer1_outputs(5402) <= not (a or b);
    layer1_outputs(5403) <= not b;
    layer1_outputs(5404) <= a;
    layer1_outputs(5405) <= not a;
    layer1_outputs(5406) <= '1';
    layer1_outputs(5407) <= not a;
    layer1_outputs(5408) <= b;
    layer1_outputs(5409) <= a xor b;
    layer1_outputs(5410) <= b and not a;
    layer1_outputs(5411) <= '1';
    layer1_outputs(5412) <= not b;
    layer1_outputs(5413) <= a and not b;
    layer1_outputs(5414) <= not (a or b);
    layer1_outputs(5415) <= not b;
    layer1_outputs(5416) <= not a;
    layer1_outputs(5417) <= a;
    layer1_outputs(5418) <= a;
    layer1_outputs(5419) <= '0';
    layer1_outputs(5420) <= a and b;
    layer1_outputs(5421) <= not a or b;
    layer1_outputs(5422) <= not a or b;
    layer1_outputs(5423) <= not b or a;
    layer1_outputs(5424) <= not b or a;
    layer1_outputs(5425) <= a;
    layer1_outputs(5426) <= a and b;
    layer1_outputs(5427) <= b;
    layer1_outputs(5428) <= a;
    layer1_outputs(5429) <= not b or a;
    layer1_outputs(5430) <= not a or b;
    layer1_outputs(5431) <= not b;
    layer1_outputs(5432) <= not a;
    layer1_outputs(5433) <= '0';
    layer1_outputs(5434) <= a and b;
    layer1_outputs(5435) <= a and not b;
    layer1_outputs(5436) <= b;
    layer1_outputs(5437) <= '0';
    layer1_outputs(5438) <= not a;
    layer1_outputs(5439) <= '1';
    layer1_outputs(5440) <= a and b;
    layer1_outputs(5441) <= not a;
    layer1_outputs(5442) <= a;
    layer1_outputs(5443) <= a;
    layer1_outputs(5444) <= not b or a;
    layer1_outputs(5445) <= '1';
    layer1_outputs(5446) <= not b;
    layer1_outputs(5447) <= not (a and b);
    layer1_outputs(5448) <= not b or a;
    layer1_outputs(5449) <= '0';
    layer1_outputs(5450) <= '1';
    layer1_outputs(5451) <= a or b;
    layer1_outputs(5452) <= b;
    layer1_outputs(5453) <= not a;
    layer1_outputs(5454) <= not a or b;
    layer1_outputs(5455) <= b;
    layer1_outputs(5456) <= a and not b;
    layer1_outputs(5457) <= not b or a;
    layer1_outputs(5458) <= not a or b;
    layer1_outputs(5459) <= not b or a;
    layer1_outputs(5460) <= a;
    layer1_outputs(5461) <= not (a or b);
    layer1_outputs(5462) <= a or b;
    layer1_outputs(5463) <= '1';
    layer1_outputs(5464) <= not b;
    layer1_outputs(5465) <= not b;
    layer1_outputs(5466) <= not (a and b);
    layer1_outputs(5467) <= not a;
    layer1_outputs(5468) <= b and not a;
    layer1_outputs(5469) <= not b or a;
    layer1_outputs(5470) <= not (a and b);
    layer1_outputs(5471) <= a;
    layer1_outputs(5472) <= a and b;
    layer1_outputs(5473) <= '1';
    layer1_outputs(5474) <= a or b;
    layer1_outputs(5475) <= b;
    layer1_outputs(5476) <= not a;
    layer1_outputs(5477) <= not (a and b);
    layer1_outputs(5478) <= a or b;
    layer1_outputs(5479) <= '0';
    layer1_outputs(5480) <= not b or a;
    layer1_outputs(5481) <= not (a xor b);
    layer1_outputs(5482) <= a;
    layer1_outputs(5483) <= a or b;
    layer1_outputs(5484) <= not a or b;
    layer1_outputs(5485) <= not a or b;
    layer1_outputs(5486) <= a and b;
    layer1_outputs(5487) <= a and not b;
    layer1_outputs(5488) <= a and b;
    layer1_outputs(5489) <= not b or a;
    layer1_outputs(5490) <= not (a xor b);
    layer1_outputs(5491) <= not a or b;
    layer1_outputs(5492) <= a and b;
    layer1_outputs(5493) <= a and b;
    layer1_outputs(5494) <= '0';
    layer1_outputs(5495) <= not (a or b);
    layer1_outputs(5496) <= not (a or b);
    layer1_outputs(5497) <= a or b;
    layer1_outputs(5498) <= b;
    layer1_outputs(5499) <= not (a xor b);
    layer1_outputs(5500) <= b;
    layer1_outputs(5501) <= not a or b;
    layer1_outputs(5502) <= not b;
    layer1_outputs(5503) <= not (a xor b);
    layer1_outputs(5504) <= '1';
    layer1_outputs(5505) <= '1';
    layer1_outputs(5506) <= not a or b;
    layer1_outputs(5507) <= not b;
    layer1_outputs(5508) <= b;
    layer1_outputs(5509) <= '0';
    layer1_outputs(5510) <= not a or b;
    layer1_outputs(5511) <= '0';
    layer1_outputs(5512) <= not (a and b);
    layer1_outputs(5513) <= '1';
    layer1_outputs(5514) <= not (a or b);
    layer1_outputs(5515) <= not b or a;
    layer1_outputs(5516) <= not b;
    layer1_outputs(5517) <= b;
    layer1_outputs(5518) <= not a;
    layer1_outputs(5519) <= not (a and b);
    layer1_outputs(5520) <= not (a or b);
    layer1_outputs(5521) <= '0';
    layer1_outputs(5522) <= not (a and b);
    layer1_outputs(5523) <= a;
    layer1_outputs(5524) <= b;
    layer1_outputs(5525) <= b and not a;
    layer1_outputs(5526) <= b;
    layer1_outputs(5527) <= a and not b;
    layer1_outputs(5528) <= b and not a;
    layer1_outputs(5529) <= not (a or b);
    layer1_outputs(5530) <= a and b;
    layer1_outputs(5531) <= '1';
    layer1_outputs(5532) <= a;
    layer1_outputs(5533) <= a;
    layer1_outputs(5534) <= a and not b;
    layer1_outputs(5535) <= not b;
    layer1_outputs(5536) <= a or b;
    layer1_outputs(5537) <= not (a or b);
    layer1_outputs(5538) <= a or b;
    layer1_outputs(5539) <= '0';
    layer1_outputs(5540) <= a and b;
    layer1_outputs(5541) <= not a or b;
    layer1_outputs(5542) <= a or b;
    layer1_outputs(5543) <= a and b;
    layer1_outputs(5544) <= '0';
    layer1_outputs(5545) <= not (a or b);
    layer1_outputs(5546) <= a;
    layer1_outputs(5547) <= a or b;
    layer1_outputs(5548) <= a xor b;
    layer1_outputs(5549) <= b and not a;
    layer1_outputs(5550) <= b;
    layer1_outputs(5551) <= not b;
    layer1_outputs(5552) <= not a or b;
    layer1_outputs(5553) <= b;
    layer1_outputs(5554) <= a and b;
    layer1_outputs(5555) <= not b;
    layer1_outputs(5556) <= not b;
    layer1_outputs(5557) <= not (a and b);
    layer1_outputs(5558) <= a or b;
    layer1_outputs(5559) <= b;
    layer1_outputs(5560) <= '0';
    layer1_outputs(5561) <= b and not a;
    layer1_outputs(5562) <= not a or b;
    layer1_outputs(5563) <= not b;
    layer1_outputs(5564) <= a;
    layer1_outputs(5565) <= not a;
    layer1_outputs(5566) <= b and not a;
    layer1_outputs(5567) <= not b;
    layer1_outputs(5568) <= not b;
    layer1_outputs(5569) <= a and b;
    layer1_outputs(5570) <= not a or b;
    layer1_outputs(5571) <= a or b;
    layer1_outputs(5572) <= a or b;
    layer1_outputs(5573) <= a and b;
    layer1_outputs(5574) <= not (a or b);
    layer1_outputs(5575) <= b;
    layer1_outputs(5576) <= not a;
    layer1_outputs(5577) <= not a;
    layer1_outputs(5578) <= '0';
    layer1_outputs(5579) <= b and not a;
    layer1_outputs(5580) <= not (a or b);
    layer1_outputs(5581) <= '1';
    layer1_outputs(5582) <= not a or b;
    layer1_outputs(5583) <= '1';
    layer1_outputs(5584) <= b;
    layer1_outputs(5585) <= not (a xor b);
    layer1_outputs(5586) <= a or b;
    layer1_outputs(5587) <= a;
    layer1_outputs(5588) <= '1';
    layer1_outputs(5589) <= a and b;
    layer1_outputs(5590) <= '0';
    layer1_outputs(5591) <= not a or b;
    layer1_outputs(5592) <= a xor b;
    layer1_outputs(5593) <= not a;
    layer1_outputs(5594) <= not (a or b);
    layer1_outputs(5595) <= a;
    layer1_outputs(5596) <= not (a and b);
    layer1_outputs(5597) <= a xor b;
    layer1_outputs(5598) <= a or b;
    layer1_outputs(5599) <= not a or b;
    layer1_outputs(5600) <= b and not a;
    layer1_outputs(5601) <= '1';
    layer1_outputs(5602) <= a;
    layer1_outputs(5603) <= '0';
    layer1_outputs(5604) <= not (a and b);
    layer1_outputs(5605) <= '1';
    layer1_outputs(5606) <= not b or a;
    layer1_outputs(5607) <= a;
    layer1_outputs(5608) <= not (a and b);
    layer1_outputs(5609) <= '0';
    layer1_outputs(5610) <= b and not a;
    layer1_outputs(5611) <= '0';
    layer1_outputs(5612) <= a or b;
    layer1_outputs(5613) <= not (a or b);
    layer1_outputs(5614) <= '1';
    layer1_outputs(5615) <= a or b;
    layer1_outputs(5616) <= not (a or b);
    layer1_outputs(5617) <= not (a or b);
    layer1_outputs(5618) <= '1';
    layer1_outputs(5619) <= not (a or b);
    layer1_outputs(5620) <= '1';
    layer1_outputs(5621) <= not a or b;
    layer1_outputs(5622) <= a or b;
    layer1_outputs(5623) <= not a or b;
    layer1_outputs(5624) <= not b;
    layer1_outputs(5625) <= a;
    layer1_outputs(5626) <= a xor b;
    layer1_outputs(5627) <= a and not b;
    layer1_outputs(5628) <= not (a and b);
    layer1_outputs(5629) <= a and not b;
    layer1_outputs(5630) <= a or b;
    layer1_outputs(5631) <= a and not b;
    layer1_outputs(5632) <= a and not b;
    layer1_outputs(5633) <= not a or b;
    layer1_outputs(5634) <= not (a xor b);
    layer1_outputs(5635) <= a and b;
    layer1_outputs(5636) <= not (a or b);
    layer1_outputs(5637) <= a or b;
    layer1_outputs(5638) <= b and not a;
    layer1_outputs(5639) <= b;
    layer1_outputs(5640) <= '1';
    layer1_outputs(5641) <= not (a or b);
    layer1_outputs(5642) <= b and not a;
    layer1_outputs(5643) <= '1';
    layer1_outputs(5644) <= b and not a;
    layer1_outputs(5645) <= '1';
    layer1_outputs(5646) <= a;
    layer1_outputs(5647) <= a and not b;
    layer1_outputs(5648) <= a;
    layer1_outputs(5649) <= not b;
    layer1_outputs(5650) <= '0';
    layer1_outputs(5651) <= a and b;
    layer1_outputs(5652) <= not a;
    layer1_outputs(5653) <= not a or b;
    layer1_outputs(5654) <= b and not a;
    layer1_outputs(5655) <= a and b;
    layer1_outputs(5656) <= not a;
    layer1_outputs(5657) <= not (a and b);
    layer1_outputs(5658) <= a;
    layer1_outputs(5659) <= b and not a;
    layer1_outputs(5660) <= b;
    layer1_outputs(5661) <= not a;
    layer1_outputs(5662) <= not a or b;
    layer1_outputs(5663) <= not (a xor b);
    layer1_outputs(5664) <= not b;
    layer1_outputs(5665) <= a;
    layer1_outputs(5666) <= not b or a;
    layer1_outputs(5667) <= not (a xor b);
    layer1_outputs(5668) <= not b;
    layer1_outputs(5669) <= a;
    layer1_outputs(5670) <= '0';
    layer1_outputs(5671) <= a xor b;
    layer1_outputs(5672) <= not b;
    layer1_outputs(5673) <= a and b;
    layer1_outputs(5674) <= not (a xor b);
    layer1_outputs(5675) <= not (a or b);
    layer1_outputs(5676) <= a;
    layer1_outputs(5677) <= '0';
    layer1_outputs(5678) <= a and not b;
    layer1_outputs(5679) <= not (a or b);
    layer1_outputs(5680) <= b and not a;
    layer1_outputs(5681) <= not b;
    layer1_outputs(5682) <= b and not a;
    layer1_outputs(5683) <= '0';
    layer1_outputs(5684) <= '1';
    layer1_outputs(5685) <= b;
    layer1_outputs(5686) <= not a or b;
    layer1_outputs(5687) <= not b or a;
    layer1_outputs(5688) <= a or b;
    layer1_outputs(5689) <= b and not a;
    layer1_outputs(5690) <= a xor b;
    layer1_outputs(5691) <= not a or b;
    layer1_outputs(5692) <= not a or b;
    layer1_outputs(5693) <= a and b;
    layer1_outputs(5694) <= not (a or b);
    layer1_outputs(5695) <= a and b;
    layer1_outputs(5696) <= not a;
    layer1_outputs(5697) <= a;
    layer1_outputs(5698) <= not b;
    layer1_outputs(5699) <= not b;
    layer1_outputs(5700) <= a and b;
    layer1_outputs(5701) <= b and not a;
    layer1_outputs(5702) <= b;
    layer1_outputs(5703) <= a xor b;
    layer1_outputs(5704) <= a;
    layer1_outputs(5705) <= not a or b;
    layer1_outputs(5706) <= '1';
    layer1_outputs(5707) <= a and b;
    layer1_outputs(5708) <= b;
    layer1_outputs(5709) <= a or b;
    layer1_outputs(5710) <= '0';
    layer1_outputs(5711) <= a and b;
    layer1_outputs(5712) <= b;
    layer1_outputs(5713) <= not (a xor b);
    layer1_outputs(5714) <= not b or a;
    layer1_outputs(5715) <= '1';
    layer1_outputs(5716) <= not a or b;
    layer1_outputs(5717) <= a or b;
    layer1_outputs(5718) <= not b or a;
    layer1_outputs(5719) <= b and not a;
    layer1_outputs(5720) <= a and not b;
    layer1_outputs(5721) <= not a or b;
    layer1_outputs(5722) <= a xor b;
    layer1_outputs(5723) <= not (a or b);
    layer1_outputs(5724) <= b;
    layer1_outputs(5725) <= a and b;
    layer1_outputs(5726) <= not b;
    layer1_outputs(5727) <= a;
    layer1_outputs(5728) <= b;
    layer1_outputs(5729) <= not b or a;
    layer1_outputs(5730) <= '1';
    layer1_outputs(5731) <= b;
    layer1_outputs(5732) <= '0';
    layer1_outputs(5733) <= not (a and b);
    layer1_outputs(5734) <= a or b;
    layer1_outputs(5735) <= not b;
    layer1_outputs(5736) <= a;
    layer1_outputs(5737) <= not a;
    layer1_outputs(5738) <= b;
    layer1_outputs(5739) <= a and not b;
    layer1_outputs(5740) <= a or b;
    layer1_outputs(5741) <= a or b;
    layer1_outputs(5742) <= a and not b;
    layer1_outputs(5743) <= b and not a;
    layer1_outputs(5744) <= b;
    layer1_outputs(5745) <= a xor b;
    layer1_outputs(5746) <= not b;
    layer1_outputs(5747) <= a and b;
    layer1_outputs(5748) <= not a;
    layer1_outputs(5749) <= '1';
    layer1_outputs(5750) <= not b or a;
    layer1_outputs(5751) <= a and b;
    layer1_outputs(5752) <= not b or a;
    layer1_outputs(5753) <= a;
    layer1_outputs(5754) <= b and not a;
    layer1_outputs(5755) <= b;
    layer1_outputs(5756) <= b and not a;
    layer1_outputs(5757) <= b;
    layer1_outputs(5758) <= not (a and b);
    layer1_outputs(5759) <= not (a and b);
    layer1_outputs(5760) <= not a;
    layer1_outputs(5761) <= a and b;
    layer1_outputs(5762) <= not a;
    layer1_outputs(5763) <= not b;
    layer1_outputs(5764) <= a and b;
    layer1_outputs(5765) <= '1';
    layer1_outputs(5766) <= a xor b;
    layer1_outputs(5767) <= not (a xor b);
    layer1_outputs(5768) <= not (a and b);
    layer1_outputs(5769) <= a and not b;
    layer1_outputs(5770) <= a and b;
    layer1_outputs(5771) <= not a;
    layer1_outputs(5772) <= '1';
    layer1_outputs(5773) <= a;
    layer1_outputs(5774) <= not b;
    layer1_outputs(5775) <= not (a or b);
    layer1_outputs(5776) <= a and not b;
    layer1_outputs(5777) <= not (a and b);
    layer1_outputs(5778) <= '0';
    layer1_outputs(5779) <= not (a and b);
    layer1_outputs(5780) <= not (a xor b);
    layer1_outputs(5781) <= not a;
    layer1_outputs(5782) <= not b or a;
    layer1_outputs(5783) <= not b or a;
    layer1_outputs(5784) <= not (a xor b);
    layer1_outputs(5785) <= not a;
    layer1_outputs(5786) <= '1';
    layer1_outputs(5787) <= not (a or b);
    layer1_outputs(5788) <= not a;
    layer1_outputs(5789) <= not (a or b);
    layer1_outputs(5790) <= b and not a;
    layer1_outputs(5791) <= '1';
    layer1_outputs(5792) <= a and b;
    layer1_outputs(5793) <= not a;
    layer1_outputs(5794) <= not b or a;
    layer1_outputs(5795) <= a;
    layer1_outputs(5796) <= not a;
    layer1_outputs(5797) <= a or b;
    layer1_outputs(5798) <= '0';
    layer1_outputs(5799) <= not a;
    layer1_outputs(5800) <= a xor b;
    layer1_outputs(5801) <= '0';
    layer1_outputs(5802) <= b and not a;
    layer1_outputs(5803) <= a xor b;
    layer1_outputs(5804) <= not b;
    layer1_outputs(5805) <= not (a and b);
    layer1_outputs(5806) <= not b or a;
    layer1_outputs(5807) <= '1';
    layer1_outputs(5808) <= a or b;
    layer1_outputs(5809) <= not b or a;
    layer1_outputs(5810) <= b and not a;
    layer1_outputs(5811) <= not b or a;
    layer1_outputs(5812) <= a;
    layer1_outputs(5813) <= a or b;
    layer1_outputs(5814) <= a xor b;
    layer1_outputs(5815) <= not (a and b);
    layer1_outputs(5816) <= a xor b;
    layer1_outputs(5817) <= not a;
    layer1_outputs(5818) <= '0';
    layer1_outputs(5819) <= a or b;
    layer1_outputs(5820) <= not (a xor b);
    layer1_outputs(5821) <= a and not b;
    layer1_outputs(5822) <= b;
    layer1_outputs(5823) <= a;
    layer1_outputs(5824) <= b;
    layer1_outputs(5825) <= '1';
    layer1_outputs(5826) <= '0';
    layer1_outputs(5827) <= not a;
    layer1_outputs(5828) <= a or b;
    layer1_outputs(5829) <= b;
    layer1_outputs(5830) <= a or b;
    layer1_outputs(5831) <= not b or a;
    layer1_outputs(5832) <= a and b;
    layer1_outputs(5833) <= not b;
    layer1_outputs(5834) <= not b or a;
    layer1_outputs(5835) <= b;
    layer1_outputs(5836) <= not a;
    layer1_outputs(5837) <= a and b;
    layer1_outputs(5838) <= a;
    layer1_outputs(5839) <= not (a or b);
    layer1_outputs(5840) <= '1';
    layer1_outputs(5841) <= a or b;
    layer1_outputs(5842) <= not a;
    layer1_outputs(5843) <= not b;
    layer1_outputs(5844) <= not a;
    layer1_outputs(5845) <= not a;
    layer1_outputs(5846) <= not (a or b);
    layer1_outputs(5847) <= not (a or b);
    layer1_outputs(5848) <= not (a and b);
    layer1_outputs(5849) <= not (a and b);
    layer1_outputs(5850) <= a xor b;
    layer1_outputs(5851) <= a or b;
    layer1_outputs(5852) <= '0';
    layer1_outputs(5853) <= not (a or b);
    layer1_outputs(5854) <= not (a and b);
    layer1_outputs(5855) <= not (a and b);
    layer1_outputs(5856) <= not (a xor b);
    layer1_outputs(5857) <= not (a and b);
    layer1_outputs(5858) <= not b;
    layer1_outputs(5859) <= a and not b;
    layer1_outputs(5860) <= not (a or b);
    layer1_outputs(5861) <= '0';
    layer1_outputs(5862) <= a xor b;
    layer1_outputs(5863) <= not (a xor b);
    layer1_outputs(5864) <= not b;
    layer1_outputs(5865) <= not (a or b);
    layer1_outputs(5866) <= '1';
    layer1_outputs(5867) <= not b or a;
    layer1_outputs(5868) <= a and not b;
    layer1_outputs(5869) <= not a or b;
    layer1_outputs(5870) <= '1';
    layer1_outputs(5871) <= b and not a;
    layer1_outputs(5872) <= not (a or b);
    layer1_outputs(5873) <= not (a and b);
    layer1_outputs(5874) <= a or b;
    layer1_outputs(5875) <= not a or b;
    layer1_outputs(5876) <= not b;
    layer1_outputs(5877) <= a;
    layer1_outputs(5878) <= a or b;
    layer1_outputs(5879) <= b;
    layer1_outputs(5880) <= not a;
    layer1_outputs(5881) <= b and not a;
    layer1_outputs(5882) <= not (a and b);
    layer1_outputs(5883) <= a;
    layer1_outputs(5884) <= not b or a;
    layer1_outputs(5885) <= '0';
    layer1_outputs(5886) <= a and b;
    layer1_outputs(5887) <= '0';
    layer1_outputs(5888) <= not a or b;
    layer1_outputs(5889) <= '1';
    layer1_outputs(5890) <= not (a or b);
    layer1_outputs(5891) <= not b or a;
    layer1_outputs(5892) <= '1';
    layer1_outputs(5893) <= a and not b;
    layer1_outputs(5894) <= a or b;
    layer1_outputs(5895) <= a or b;
    layer1_outputs(5896) <= a and not b;
    layer1_outputs(5897) <= not (a or b);
    layer1_outputs(5898) <= not b;
    layer1_outputs(5899) <= '0';
    layer1_outputs(5900) <= not (a or b);
    layer1_outputs(5901) <= b;
    layer1_outputs(5902) <= a and b;
    layer1_outputs(5903) <= a xor b;
    layer1_outputs(5904) <= not a or b;
    layer1_outputs(5905) <= a and not b;
    layer1_outputs(5906) <= a or b;
    layer1_outputs(5907) <= a;
    layer1_outputs(5908) <= not (a or b);
    layer1_outputs(5909) <= a and b;
    layer1_outputs(5910) <= not b;
    layer1_outputs(5911) <= not (a and b);
    layer1_outputs(5912) <= b;
    layer1_outputs(5913) <= not a or b;
    layer1_outputs(5914) <= a;
    layer1_outputs(5915) <= a xor b;
    layer1_outputs(5916) <= b;
    layer1_outputs(5917) <= '0';
    layer1_outputs(5918) <= b and not a;
    layer1_outputs(5919) <= not b;
    layer1_outputs(5920) <= not (a and b);
    layer1_outputs(5921) <= not b;
    layer1_outputs(5922) <= '1';
    layer1_outputs(5923) <= '1';
    layer1_outputs(5924) <= not a or b;
    layer1_outputs(5925) <= a or b;
    layer1_outputs(5926) <= not b or a;
    layer1_outputs(5927) <= b and not a;
    layer1_outputs(5928) <= a and b;
    layer1_outputs(5929) <= b and not a;
    layer1_outputs(5930) <= not b;
    layer1_outputs(5931) <= a;
    layer1_outputs(5932) <= a and not b;
    layer1_outputs(5933) <= not b;
    layer1_outputs(5934) <= not b;
    layer1_outputs(5935) <= a;
    layer1_outputs(5936) <= not (a or b);
    layer1_outputs(5937) <= b and not a;
    layer1_outputs(5938) <= '1';
    layer1_outputs(5939) <= not b;
    layer1_outputs(5940) <= a or b;
    layer1_outputs(5941) <= not b or a;
    layer1_outputs(5942) <= '1';
    layer1_outputs(5943) <= not b;
    layer1_outputs(5944) <= not (a or b);
    layer1_outputs(5945) <= not b;
    layer1_outputs(5946) <= not b or a;
    layer1_outputs(5947) <= not (a or b);
    layer1_outputs(5948) <= not a or b;
    layer1_outputs(5949) <= b and not a;
    layer1_outputs(5950) <= not b or a;
    layer1_outputs(5951) <= a and b;
    layer1_outputs(5952) <= b;
    layer1_outputs(5953) <= '1';
    layer1_outputs(5954) <= not b;
    layer1_outputs(5955) <= not (a or b);
    layer1_outputs(5956) <= a or b;
    layer1_outputs(5957) <= a;
    layer1_outputs(5958) <= '0';
    layer1_outputs(5959) <= a or b;
    layer1_outputs(5960) <= not b or a;
    layer1_outputs(5961) <= not b;
    layer1_outputs(5962) <= a and not b;
    layer1_outputs(5963) <= '1';
    layer1_outputs(5964) <= '1';
    layer1_outputs(5965) <= not b;
    layer1_outputs(5966) <= b and not a;
    layer1_outputs(5967) <= a and b;
    layer1_outputs(5968) <= a;
    layer1_outputs(5969) <= a or b;
    layer1_outputs(5970) <= not b or a;
    layer1_outputs(5971) <= not b or a;
    layer1_outputs(5972) <= a or b;
    layer1_outputs(5973) <= b and not a;
    layer1_outputs(5974) <= b;
    layer1_outputs(5975) <= a;
    layer1_outputs(5976) <= not a or b;
    layer1_outputs(5977) <= not (a and b);
    layer1_outputs(5978) <= not a;
    layer1_outputs(5979) <= a and not b;
    layer1_outputs(5980) <= b and not a;
    layer1_outputs(5981) <= not a or b;
    layer1_outputs(5982) <= a and b;
    layer1_outputs(5983) <= a xor b;
    layer1_outputs(5984) <= not (a and b);
    layer1_outputs(5985) <= a and not b;
    layer1_outputs(5986) <= a or b;
    layer1_outputs(5987) <= not b;
    layer1_outputs(5988) <= not b;
    layer1_outputs(5989) <= a xor b;
    layer1_outputs(5990) <= a xor b;
    layer1_outputs(5991) <= a and not b;
    layer1_outputs(5992) <= b;
    layer1_outputs(5993) <= a and not b;
    layer1_outputs(5994) <= not (a xor b);
    layer1_outputs(5995) <= not (a or b);
    layer1_outputs(5996) <= b and not a;
    layer1_outputs(5997) <= not (a or b);
    layer1_outputs(5998) <= a or b;
    layer1_outputs(5999) <= b and not a;
    layer1_outputs(6000) <= '0';
    layer1_outputs(6001) <= a or b;
    layer1_outputs(6002) <= not b or a;
    layer1_outputs(6003) <= a or b;
    layer1_outputs(6004) <= not b;
    layer1_outputs(6005) <= not a;
    layer1_outputs(6006) <= '0';
    layer1_outputs(6007) <= b and not a;
    layer1_outputs(6008) <= a;
    layer1_outputs(6009) <= not (a or b);
    layer1_outputs(6010) <= a or b;
    layer1_outputs(6011) <= not b;
    layer1_outputs(6012) <= not b;
    layer1_outputs(6013) <= '0';
    layer1_outputs(6014) <= not (a or b);
    layer1_outputs(6015) <= '1';
    layer1_outputs(6016) <= a and b;
    layer1_outputs(6017) <= not b;
    layer1_outputs(6018) <= a or b;
    layer1_outputs(6019) <= '0';
    layer1_outputs(6020) <= a and b;
    layer1_outputs(6021) <= not (a xor b);
    layer1_outputs(6022) <= a and not b;
    layer1_outputs(6023) <= not a;
    layer1_outputs(6024) <= not (a and b);
    layer1_outputs(6025) <= a or b;
    layer1_outputs(6026) <= not a;
    layer1_outputs(6027) <= a and not b;
    layer1_outputs(6028) <= a and not b;
    layer1_outputs(6029) <= a;
    layer1_outputs(6030) <= not a;
    layer1_outputs(6031) <= '0';
    layer1_outputs(6032) <= b and not a;
    layer1_outputs(6033) <= a and not b;
    layer1_outputs(6034) <= a;
    layer1_outputs(6035) <= b and not a;
    layer1_outputs(6036) <= a xor b;
    layer1_outputs(6037) <= not (a or b);
    layer1_outputs(6038) <= '0';
    layer1_outputs(6039) <= a and b;
    layer1_outputs(6040) <= '0';
    layer1_outputs(6041) <= b;
    layer1_outputs(6042) <= '1';
    layer1_outputs(6043) <= b;
    layer1_outputs(6044) <= not a;
    layer1_outputs(6045) <= a and b;
    layer1_outputs(6046) <= not b or a;
    layer1_outputs(6047) <= a and not b;
    layer1_outputs(6048) <= b;
    layer1_outputs(6049) <= b;
    layer1_outputs(6050) <= not (a xor b);
    layer1_outputs(6051) <= not a or b;
    layer1_outputs(6052) <= not (a or b);
    layer1_outputs(6053) <= a;
    layer1_outputs(6054) <= not (a xor b);
    layer1_outputs(6055) <= not (a and b);
    layer1_outputs(6056) <= '1';
    layer1_outputs(6057) <= a;
    layer1_outputs(6058) <= a;
    layer1_outputs(6059) <= not (a or b);
    layer1_outputs(6060) <= a or b;
    layer1_outputs(6061) <= not b;
    layer1_outputs(6062) <= not (a xor b);
    layer1_outputs(6063) <= not a;
    layer1_outputs(6064) <= '0';
    layer1_outputs(6065) <= not b;
    layer1_outputs(6066) <= not b or a;
    layer1_outputs(6067) <= a and not b;
    layer1_outputs(6068) <= a;
    layer1_outputs(6069) <= not a or b;
    layer1_outputs(6070) <= a and not b;
    layer1_outputs(6071) <= a;
    layer1_outputs(6072) <= a and not b;
    layer1_outputs(6073) <= a and not b;
    layer1_outputs(6074) <= not a or b;
    layer1_outputs(6075) <= b;
    layer1_outputs(6076) <= not a or b;
    layer1_outputs(6077) <= a or b;
    layer1_outputs(6078) <= a xor b;
    layer1_outputs(6079) <= a and b;
    layer1_outputs(6080) <= a;
    layer1_outputs(6081) <= b and not a;
    layer1_outputs(6082) <= a or b;
    layer1_outputs(6083) <= a and b;
    layer1_outputs(6084) <= not (a or b);
    layer1_outputs(6085) <= '0';
    layer1_outputs(6086) <= not a;
    layer1_outputs(6087) <= b and not a;
    layer1_outputs(6088) <= not a or b;
    layer1_outputs(6089) <= b;
    layer1_outputs(6090) <= not b or a;
    layer1_outputs(6091) <= not b or a;
    layer1_outputs(6092) <= not b;
    layer1_outputs(6093) <= a and not b;
    layer1_outputs(6094) <= '0';
    layer1_outputs(6095) <= b and not a;
    layer1_outputs(6096) <= not a;
    layer1_outputs(6097) <= not b or a;
    layer1_outputs(6098) <= not (a and b);
    layer1_outputs(6099) <= not b;
    layer1_outputs(6100) <= not a;
    layer1_outputs(6101) <= not a or b;
    layer1_outputs(6102) <= not b;
    layer1_outputs(6103) <= b;
    layer1_outputs(6104) <= not (a and b);
    layer1_outputs(6105) <= not (a and b);
    layer1_outputs(6106) <= a and not b;
    layer1_outputs(6107) <= not (a or b);
    layer1_outputs(6108) <= not a or b;
    layer1_outputs(6109) <= a or b;
    layer1_outputs(6110) <= a and b;
    layer1_outputs(6111) <= not a or b;
    layer1_outputs(6112) <= a or b;
    layer1_outputs(6113) <= a;
    layer1_outputs(6114) <= not a or b;
    layer1_outputs(6115) <= b;
    layer1_outputs(6116) <= b and not a;
    layer1_outputs(6117) <= not b;
    layer1_outputs(6118) <= not a;
    layer1_outputs(6119) <= not (a and b);
    layer1_outputs(6120) <= '0';
    layer1_outputs(6121) <= a or b;
    layer1_outputs(6122) <= not b or a;
    layer1_outputs(6123) <= not (a and b);
    layer1_outputs(6124) <= a and not b;
    layer1_outputs(6125) <= a or b;
    layer1_outputs(6126) <= a;
    layer1_outputs(6127) <= b and not a;
    layer1_outputs(6128) <= not (a and b);
    layer1_outputs(6129) <= not a or b;
    layer1_outputs(6130) <= b and not a;
    layer1_outputs(6131) <= not a;
    layer1_outputs(6132) <= b;
    layer1_outputs(6133) <= a;
    layer1_outputs(6134) <= not a;
    layer1_outputs(6135) <= a and not b;
    layer1_outputs(6136) <= not b or a;
    layer1_outputs(6137) <= b;
    layer1_outputs(6138) <= not b;
    layer1_outputs(6139) <= a;
    layer1_outputs(6140) <= a and not b;
    layer1_outputs(6141) <= a;
    layer1_outputs(6142) <= '1';
    layer1_outputs(6143) <= '1';
    layer1_outputs(6144) <= a;
    layer1_outputs(6145) <= not b or a;
    layer1_outputs(6146) <= not a or b;
    layer1_outputs(6147) <= b and not a;
    layer1_outputs(6148) <= a;
    layer1_outputs(6149) <= a;
    layer1_outputs(6150) <= b and not a;
    layer1_outputs(6151) <= a xor b;
    layer1_outputs(6152) <= a xor b;
    layer1_outputs(6153) <= not b or a;
    layer1_outputs(6154) <= b and not a;
    layer1_outputs(6155) <= a and b;
    layer1_outputs(6156) <= '1';
    layer1_outputs(6157) <= not a or b;
    layer1_outputs(6158) <= b and not a;
    layer1_outputs(6159) <= not (a and b);
    layer1_outputs(6160) <= '1';
    layer1_outputs(6161) <= '1';
    layer1_outputs(6162) <= a and b;
    layer1_outputs(6163) <= a and b;
    layer1_outputs(6164) <= not b or a;
    layer1_outputs(6165) <= b and not a;
    layer1_outputs(6166) <= not b or a;
    layer1_outputs(6167) <= not a;
    layer1_outputs(6168) <= b;
    layer1_outputs(6169) <= '1';
    layer1_outputs(6170) <= a or b;
    layer1_outputs(6171) <= b and not a;
    layer1_outputs(6172) <= a;
    layer1_outputs(6173) <= b and not a;
    layer1_outputs(6174) <= a xor b;
    layer1_outputs(6175) <= not b;
    layer1_outputs(6176) <= '1';
    layer1_outputs(6177) <= '0';
    layer1_outputs(6178) <= not b or a;
    layer1_outputs(6179) <= '1';
    layer1_outputs(6180) <= a and not b;
    layer1_outputs(6181) <= not a;
    layer1_outputs(6182) <= a and not b;
    layer1_outputs(6183) <= not (a and b);
    layer1_outputs(6184) <= b and not a;
    layer1_outputs(6185) <= not (a and b);
    layer1_outputs(6186) <= a and b;
    layer1_outputs(6187) <= not (a or b);
    layer1_outputs(6188) <= b;
    layer1_outputs(6189) <= a and b;
    layer1_outputs(6190) <= a and not b;
    layer1_outputs(6191) <= not a or b;
    layer1_outputs(6192) <= not (a and b);
    layer1_outputs(6193) <= a;
    layer1_outputs(6194) <= not a;
    layer1_outputs(6195) <= a xor b;
    layer1_outputs(6196) <= not (a and b);
    layer1_outputs(6197) <= a and b;
    layer1_outputs(6198) <= a and b;
    layer1_outputs(6199) <= not (a or b);
    layer1_outputs(6200) <= not b;
    layer1_outputs(6201) <= not a;
    layer1_outputs(6202) <= a or b;
    layer1_outputs(6203) <= '1';
    layer1_outputs(6204) <= '1';
    layer1_outputs(6205) <= a or b;
    layer1_outputs(6206) <= b;
    layer1_outputs(6207) <= '1';
    layer1_outputs(6208) <= b;
    layer1_outputs(6209) <= a or b;
    layer1_outputs(6210) <= not b;
    layer1_outputs(6211) <= a and b;
    layer1_outputs(6212) <= not a;
    layer1_outputs(6213) <= a;
    layer1_outputs(6214) <= '0';
    layer1_outputs(6215) <= a and not b;
    layer1_outputs(6216) <= not (a and b);
    layer1_outputs(6217) <= a xor b;
    layer1_outputs(6218) <= not b;
    layer1_outputs(6219) <= not b or a;
    layer1_outputs(6220) <= a and not b;
    layer1_outputs(6221) <= '1';
    layer1_outputs(6222) <= not a;
    layer1_outputs(6223) <= not (a xor b);
    layer1_outputs(6224) <= not (a or b);
    layer1_outputs(6225) <= '1';
    layer1_outputs(6226) <= a;
    layer1_outputs(6227) <= not b or a;
    layer1_outputs(6228) <= not (a xor b);
    layer1_outputs(6229) <= '1';
    layer1_outputs(6230) <= not (a xor b);
    layer1_outputs(6231) <= not a;
    layer1_outputs(6232) <= a and not b;
    layer1_outputs(6233) <= not (a or b);
    layer1_outputs(6234) <= a and b;
    layer1_outputs(6235) <= not a;
    layer1_outputs(6236) <= a and b;
    layer1_outputs(6237) <= a or b;
    layer1_outputs(6238) <= not (a or b);
    layer1_outputs(6239) <= not (a and b);
    layer1_outputs(6240) <= a and not b;
    layer1_outputs(6241) <= b and not a;
    layer1_outputs(6242) <= '0';
    layer1_outputs(6243) <= not b;
    layer1_outputs(6244) <= a;
    layer1_outputs(6245) <= not (a or b);
    layer1_outputs(6246) <= not b or a;
    layer1_outputs(6247) <= '0';
    layer1_outputs(6248) <= not b or a;
    layer1_outputs(6249) <= not a;
    layer1_outputs(6250) <= not a or b;
    layer1_outputs(6251) <= not b or a;
    layer1_outputs(6252) <= '1';
    layer1_outputs(6253) <= b;
    layer1_outputs(6254) <= a;
    layer1_outputs(6255) <= '1';
    layer1_outputs(6256) <= a and b;
    layer1_outputs(6257) <= not a or b;
    layer1_outputs(6258) <= a or b;
    layer1_outputs(6259) <= a and not b;
    layer1_outputs(6260) <= b;
    layer1_outputs(6261) <= not a or b;
    layer1_outputs(6262) <= a or b;
    layer1_outputs(6263) <= a;
    layer1_outputs(6264) <= '0';
    layer1_outputs(6265) <= a or b;
    layer1_outputs(6266) <= a and b;
    layer1_outputs(6267) <= b;
    layer1_outputs(6268) <= '1';
    layer1_outputs(6269) <= not (a or b);
    layer1_outputs(6270) <= b and not a;
    layer1_outputs(6271) <= a xor b;
    layer1_outputs(6272) <= b;
    layer1_outputs(6273) <= a;
    layer1_outputs(6274) <= b;
    layer1_outputs(6275) <= not b or a;
    layer1_outputs(6276) <= a;
    layer1_outputs(6277) <= b;
    layer1_outputs(6278) <= not a;
    layer1_outputs(6279) <= a;
    layer1_outputs(6280) <= not (a xor b);
    layer1_outputs(6281) <= b;
    layer1_outputs(6282) <= a or b;
    layer1_outputs(6283) <= b and not a;
    layer1_outputs(6284) <= not a or b;
    layer1_outputs(6285) <= not b or a;
    layer1_outputs(6286) <= not b;
    layer1_outputs(6287) <= '0';
    layer1_outputs(6288) <= b and not a;
    layer1_outputs(6289) <= not a;
    layer1_outputs(6290) <= '1';
    layer1_outputs(6291) <= a or b;
    layer1_outputs(6292) <= a or b;
    layer1_outputs(6293) <= '0';
    layer1_outputs(6294) <= a or b;
    layer1_outputs(6295) <= '0';
    layer1_outputs(6296) <= b and not a;
    layer1_outputs(6297) <= a and not b;
    layer1_outputs(6298) <= b;
    layer1_outputs(6299) <= a and b;
    layer1_outputs(6300) <= '1';
    layer1_outputs(6301) <= not a or b;
    layer1_outputs(6302) <= a and b;
    layer1_outputs(6303) <= not b;
    layer1_outputs(6304) <= a and b;
    layer1_outputs(6305) <= a and b;
    layer1_outputs(6306) <= a and not b;
    layer1_outputs(6307) <= b;
    layer1_outputs(6308) <= a and not b;
    layer1_outputs(6309) <= a and not b;
    layer1_outputs(6310) <= b;
    layer1_outputs(6311) <= a or b;
    layer1_outputs(6312) <= not a;
    layer1_outputs(6313) <= a;
    layer1_outputs(6314) <= not b or a;
    layer1_outputs(6315) <= not a or b;
    layer1_outputs(6316) <= b;
    layer1_outputs(6317) <= not a;
    layer1_outputs(6318) <= not b;
    layer1_outputs(6319) <= not a or b;
    layer1_outputs(6320) <= b;
    layer1_outputs(6321) <= '1';
    layer1_outputs(6322) <= a;
    layer1_outputs(6323) <= a or b;
    layer1_outputs(6324) <= a xor b;
    layer1_outputs(6325) <= a or b;
    layer1_outputs(6326) <= not (a and b);
    layer1_outputs(6327) <= not (a and b);
    layer1_outputs(6328) <= '1';
    layer1_outputs(6329) <= not a;
    layer1_outputs(6330) <= '1';
    layer1_outputs(6331) <= '1';
    layer1_outputs(6332) <= b;
    layer1_outputs(6333) <= b;
    layer1_outputs(6334) <= a and b;
    layer1_outputs(6335) <= not a;
    layer1_outputs(6336) <= '0';
    layer1_outputs(6337) <= a;
    layer1_outputs(6338) <= not b;
    layer1_outputs(6339) <= not a;
    layer1_outputs(6340) <= a xor b;
    layer1_outputs(6341) <= b;
    layer1_outputs(6342) <= not b;
    layer1_outputs(6343) <= a or b;
    layer1_outputs(6344) <= not (a and b);
    layer1_outputs(6345) <= not a;
    layer1_outputs(6346) <= not b;
    layer1_outputs(6347) <= a and not b;
    layer1_outputs(6348) <= a or b;
    layer1_outputs(6349) <= '1';
    layer1_outputs(6350) <= not a or b;
    layer1_outputs(6351) <= a or b;
    layer1_outputs(6352) <= a xor b;
    layer1_outputs(6353) <= not a or b;
    layer1_outputs(6354) <= b;
    layer1_outputs(6355) <= b and not a;
    layer1_outputs(6356) <= a;
    layer1_outputs(6357) <= not (a xor b);
    layer1_outputs(6358) <= not (a or b);
    layer1_outputs(6359) <= '1';
    layer1_outputs(6360) <= not (a xor b);
    layer1_outputs(6361) <= not b;
    layer1_outputs(6362) <= a xor b;
    layer1_outputs(6363) <= a or b;
    layer1_outputs(6364) <= a xor b;
    layer1_outputs(6365) <= not (a or b);
    layer1_outputs(6366) <= not (a or b);
    layer1_outputs(6367) <= a or b;
    layer1_outputs(6368) <= b and not a;
    layer1_outputs(6369) <= '1';
    layer1_outputs(6370) <= not (a or b);
    layer1_outputs(6371) <= a and b;
    layer1_outputs(6372) <= not (a or b);
    layer1_outputs(6373) <= not b or a;
    layer1_outputs(6374) <= a and not b;
    layer1_outputs(6375) <= b and not a;
    layer1_outputs(6376) <= b;
    layer1_outputs(6377) <= a or b;
    layer1_outputs(6378) <= not a;
    layer1_outputs(6379) <= '0';
    layer1_outputs(6380) <= a and not b;
    layer1_outputs(6381) <= '1';
    layer1_outputs(6382) <= '0';
    layer1_outputs(6383) <= a and not b;
    layer1_outputs(6384) <= not b;
    layer1_outputs(6385) <= a or b;
    layer1_outputs(6386) <= not b or a;
    layer1_outputs(6387) <= not b;
    layer1_outputs(6388) <= not a;
    layer1_outputs(6389) <= a xor b;
    layer1_outputs(6390) <= not (a and b);
    layer1_outputs(6391) <= '1';
    layer1_outputs(6392) <= b and not a;
    layer1_outputs(6393) <= not b or a;
    layer1_outputs(6394) <= '1';
    layer1_outputs(6395) <= a and b;
    layer1_outputs(6396) <= not a;
    layer1_outputs(6397) <= b;
    layer1_outputs(6398) <= a and b;
    layer1_outputs(6399) <= not (a or b);
    layer1_outputs(6400) <= a or b;
    layer1_outputs(6401) <= a or b;
    layer1_outputs(6402) <= not a or b;
    layer1_outputs(6403) <= a;
    layer1_outputs(6404) <= a;
    layer1_outputs(6405) <= not b;
    layer1_outputs(6406) <= '0';
    layer1_outputs(6407) <= b;
    layer1_outputs(6408) <= a;
    layer1_outputs(6409) <= a and b;
    layer1_outputs(6410) <= '1';
    layer1_outputs(6411) <= not (a xor b);
    layer1_outputs(6412) <= a and b;
    layer1_outputs(6413) <= not (a and b);
    layer1_outputs(6414) <= not (a or b);
    layer1_outputs(6415) <= a;
    layer1_outputs(6416) <= a or b;
    layer1_outputs(6417) <= not a;
    layer1_outputs(6418) <= not a or b;
    layer1_outputs(6419) <= '1';
    layer1_outputs(6420) <= not a;
    layer1_outputs(6421) <= not (a xor b);
    layer1_outputs(6422) <= b;
    layer1_outputs(6423) <= not a or b;
    layer1_outputs(6424) <= a and b;
    layer1_outputs(6425) <= not b or a;
    layer1_outputs(6426) <= b;
    layer1_outputs(6427) <= not b;
    layer1_outputs(6428) <= not b or a;
    layer1_outputs(6429) <= not b or a;
    layer1_outputs(6430) <= a;
    layer1_outputs(6431) <= a;
    layer1_outputs(6432) <= not (a xor b);
    layer1_outputs(6433) <= a and b;
    layer1_outputs(6434) <= not (a or b);
    layer1_outputs(6435) <= a and b;
    layer1_outputs(6436) <= a;
    layer1_outputs(6437) <= not a;
    layer1_outputs(6438) <= a or b;
    layer1_outputs(6439) <= b;
    layer1_outputs(6440) <= '1';
    layer1_outputs(6441) <= not b;
    layer1_outputs(6442) <= not a;
    layer1_outputs(6443) <= not (a xor b);
    layer1_outputs(6444) <= '1';
    layer1_outputs(6445) <= a or b;
    layer1_outputs(6446) <= not b or a;
    layer1_outputs(6447) <= a and not b;
    layer1_outputs(6448) <= not b or a;
    layer1_outputs(6449) <= a;
    layer1_outputs(6450) <= '0';
    layer1_outputs(6451) <= b and not a;
    layer1_outputs(6452) <= not a;
    layer1_outputs(6453) <= not (a or b);
    layer1_outputs(6454) <= not (a and b);
    layer1_outputs(6455) <= '1';
    layer1_outputs(6456) <= a and not b;
    layer1_outputs(6457) <= not (a and b);
    layer1_outputs(6458) <= not a;
    layer1_outputs(6459) <= b and not a;
    layer1_outputs(6460) <= not a;
    layer1_outputs(6461) <= b;
    layer1_outputs(6462) <= a;
    layer1_outputs(6463) <= not a or b;
    layer1_outputs(6464) <= '1';
    layer1_outputs(6465) <= b;
    layer1_outputs(6466) <= not a;
    layer1_outputs(6467) <= '0';
    layer1_outputs(6468) <= not (a and b);
    layer1_outputs(6469) <= '0';
    layer1_outputs(6470) <= not (a or b);
    layer1_outputs(6471) <= a and b;
    layer1_outputs(6472) <= not a or b;
    layer1_outputs(6473) <= a xor b;
    layer1_outputs(6474) <= b;
    layer1_outputs(6475) <= not b;
    layer1_outputs(6476) <= not (a or b);
    layer1_outputs(6477) <= a or b;
    layer1_outputs(6478) <= not a;
    layer1_outputs(6479) <= not b;
    layer1_outputs(6480) <= a and not b;
    layer1_outputs(6481) <= b and not a;
    layer1_outputs(6482) <= a or b;
    layer1_outputs(6483) <= a;
    layer1_outputs(6484) <= not a;
    layer1_outputs(6485) <= '0';
    layer1_outputs(6486) <= b and not a;
    layer1_outputs(6487) <= not a or b;
    layer1_outputs(6488) <= b and not a;
    layer1_outputs(6489) <= not a or b;
    layer1_outputs(6490) <= not (a and b);
    layer1_outputs(6491) <= b;
    layer1_outputs(6492) <= a and not b;
    layer1_outputs(6493) <= b;
    layer1_outputs(6494) <= a and not b;
    layer1_outputs(6495) <= a or b;
    layer1_outputs(6496) <= not b or a;
    layer1_outputs(6497) <= a and b;
    layer1_outputs(6498) <= b;
    layer1_outputs(6499) <= not (a and b);
    layer1_outputs(6500) <= not (a or b);
    layer1_outputs(6501) <= not b;
    layer1_outputs(6502) <= a xor b;
    layer1_outputs(6503) <= b;
    layer1_outputs(6504) <= not (a or b);
    layer1_outputs(6505) <= '1';
    layer1_outputs(6506) <= a or b;
    layer1_outputs(6507) <= not (a or b);
    layer1_outputs(6508) <= a and not b;
    layer1_outputs(6509) <= not a or b;
    layer1_outputs(6510) <= a;
    layer1_outputs(6511) <= b;
    layer1_outputs(6512) <= b;
    layer1_outputs(6513) <= not a;
    layer1_outputs(6514) <= not (a and b);
    layer1_outputs(6515) <= b and not a;
    layer1_outputs(6516) <= not a;
    layer1_outputs(6517) <= not a or b;
    layer1_outputs(6518) <= a and b;
    layer1_outputs(6519) <= not (a xor b);
    layer1_outputs(6520) <= not a or b;
    layer1_outputs(6521) <= '1';
    layer1_outputs(6522) <= '0';
    layer1_outputs(6523) <= a;
    layer1_outputs(6524) <= not (a and b);
    layer1_outputs(6525) <= not b;
    layer1_outputs(6526) <= a xor b;
    layer1_outputs(6527) <= not (a and b);
    layer1_outputs(6528) <= not b or a;
    layer1_outputs(6529) <= not a;
    layer1_outputs(6530) <= b;
    layer1_outputs(6531) <= b and not a;
    layer1_outputs(6532) <= not a;
    layer1_outputs(6533) <= b and not a;
    layer1_outputs(6534) <= a and not b;
    layer1_outputs(6535) <= not a;
    layer1_outputs(6536) <= a;
    layer1_outputs(6537) <= '0';
    layer1_outputs(6538) <= not (a xor b);
    layer1_outputs(6539) <= a and b;
    layer1_outputs(6540) <= '1';
    layer1_outputs(6541) <= '0';
    layer1_outputs(6542) <= a and b;
    layer1_outputs(6543) <= not (a and b);
    layer1_outputs(6544) <= not a or b;
    layer1_outputs(6545) <= a and b;
    layer1_outputs(6546) <= a or b;
    layer1_outputs(6547) <= not b or a;
    layer1_outputs(6548) <= not a or b;
    layer1_outputs(6549) <= not (a and b);
    layer1_outputs(6550) <= not b or a;
    layer1_outputs(6551) <= a xor b;
    layer1_outputs(6552) <= not b or a;
    layer1_outputs(6553) <= '0';
    layer1_outputs(6554) <= a;
    layer1_outputs(6555) <= a or b;
    layer1_outputs(6556) <= not a;
    layer1_outputs(6557) <= not (a and b);
    layer1_outputs(6558) <= b;
    layer1_outputs(6559) <= a xor b;
    layer1_outputs(6560) <= not b or a;
    layer1_outputs(6561) <= not a or b;
    layer1_outputs(6562) <= a or b;
    layer1_outputs(6563) <= not b;
    layer1_outputs(6564) <= not b or a;
    layer1_outputs(6565) <= a or b;
    layer1_outputs(6566) <= '0';
    layer1_outputs(6567) <= not a;
    layer1_outputs(6568) <= b and not a;
    layer1_outputs(6569) <= not (a and b);
    layer1_outputs(6570) <= not b or a;
    layer1_outputs(6571) <= '0';
    layer1_outputs(6572) <= '0';
    layer1_outputs(6573) <= '1';
    layer1_outputs(6574) <= a and not b;
    layer1_outputs(6575) <= '0';
    layer1_outputs(6576) <= not a;
    layer1_outputs(6577) <= b;
    layer1_outputs(6578) <= a or b;
    layer1_outputs(6579) <= not b or a;
    layer1_outputs(6580) <= a;
    layer1_outputs(6581) <= a and not b;
    layer1_outputs(6582) <= b;
    layer1_outputs(6583) <= b and not a;
    layer1_outputs(6584) <= not b;
    layer1_outputs(6585) <= a and not b;
    layer1_outputs(6586) <= a xor b;
    layer1_outputs(6587) <= not b or a;
    layer1_outputs(6588) <= a;
    layer1_outputs(6589) <= not (a xor b);
    layer1_outputs(6590) <= not a or b;
    layer1_outputs(6591) <= '0';
    layer1_outputs(6592) <= not b or a;
    layer1_outputs(6593) <= a or b;
    layer1_outputs(6594) <= not a or b;
    layer1_outputs(6595) <= b;
    layer1_outputs(6596) <= a or b;
    layer1_outputs(6597) <= not a;
    layer1_outputs(6598) <= a and not b;
    layer1_outputs(6599) <= '1';
    layer1_outputs(6600) <= not a or b;
    layer1_outputs(6601) <= not a;
    layer1_outputs(6602) <= not b;
    layer1_outputs(6603) <= not a;
    layer1_outputs(6604) <= not (a or b);
    layer1_outputs(6605) <= not (a and b);
    layer1_outputs(6606) <= '0';
    layer1_outputs(6607) <= not (a or b);
    layer1_outputs(6608) <= not b;
    layer1_outputs(6609) <= not b;
    layer1_outputs(6610) <= b;
    layer1_outputs(6611) <= a xor b;
    layer1_outputs(6612) <= not (a and b);
    layer1_outputs(6613) <= b and not a;
    layer1_outputs(6614) <= b and not a;
    layer1_outputs(6615) <= not b;
    layer1_outputs(6616) <= a or b;
    layer1_outputs(6617) <= a and not b;
    layer1_outputs(6618) <= not b or a;
    layer1_outputs(6619) <= not b or a;
    layer1_outputs(6620) <= not a;
    layer1_outputs(6621) <= a and b;
    layer1_outputs(6622) <= not b;
    layer1_outputs(6623) <= a and b;
    layer1_outputs(6624) <= a;
    layer1_outputs(6625) <= a and not b;
    layer1_outputs(6626) <= '0';
    layer1_outputs(6627) <= b;
    layer1_outputs(6628) <= b and not a;
    layer1_outputs(6629) <= not (a or b);
    layer1_outputs(6630) <= a or b;
    layer1_outputs(6631) <= not a or b;
    layer1_outputs(6632) <= not a or b;
    layer1_outputs(6633) <= not b;
    layer1_outputs(6634) <= a;
    layer1_outputs(6635) <= not b or a;
    layer1_outputs(6636) <= a or b;
    layer1_outputs(6637) <= a;
    layer1_outputs(6638) <= a and not b;
    layer1_outputs(6639) <= not (a xor b);
    layer1_outputs(6640) <= not a;
    layer1_outputs(6641) <= not b or a;
    layer1_outputs(6642) <= not a;
    layer1_outputs(6643) <= b and not a;
    layer1_outputs(6644) <= not (a and b);
    layer1_outputs(6645) <= not (a or b);
    layer1_outputs(6646) <= a xor b;
    layer1_outputs(6647) <= not b;
    layer1_outputs(6648) <= not (a and b);
    layer1_outputs(6649) <= not b or a;
    layer1_outputs(6650) <= not b;
    layer1_outputs(6651) <= not (a and b);
    layer1_outputs(6652) <= '1';
    layer1_outputs(6653) <= b;
    layer1_outputs(6654) <= not b or a;
    layer1_outputs(6655) <= b;
    layer1_outputs(6656) <= not a or b;
    layer1_outputs(6657) <= b and not a;
    layer1_outputs(6658) <= a xor b;
    layer1_outputs(6659) <= not a;
    layer1_outputs(6660) <= b and not a;
    layer1_outputs(6661) <= a or b;
    layer1_outputs(6662) <= not b or a;
    layer1_outputs(6663) <= not (a or b);
    layer1_outputs(6664) <= not a or b;
    layer1_outputs(6665) <= b and not a;
    layer1_outputs(6666) <= not (a and b);
    layer1_outputs(6667) <= not b;
    layer1_outputs(6668) <= a;
    layer1_outputs(6669) <= a or b;
    layer1_outputs(6670) <= a and not b;
    layer1_outputs(6671) <= a;
    layer1_outputs(6672) <= a;
    layer1_outputs(6673) <= b;
    layer1_outputs(6674) <= a and not b;
    layer1_outputs(6675) <= b;
    layer1_outputs(6676) <= not a or b;
    layer1_outputs(6677) <= not a or b;
    layer1_outputs(6678) <= not b;
    layer1_outputs(6679) <= not (a or b);
    layer1_outputs(6680) <= '0';
    layer1_outputs(6681) <= not b or a;
    layer1_outputs(6682) <= not b or a;
    layer1_outputs(6683) <= b;
    layer1_outputs(6684) <= a;
    layer1_outputs(6685) <= a;
    layer1_outputs(6686) <= '0';
    layer1_outputs(6687) <= not b or a;
    layer1_outputs(6688) <= b and not a;
    layer1_outputs(6689) <= '1';
    layer1_outputs(6690) <= not b;
    layer1_outputs(6691) <= not a or b;
    layer1_outputs(6692) <= not (a or b);
    layer1_outputs(6693) <= a;
    layer1_outputs(6694) <= not a;
    layer1_outputs(6695) <= a and not b;
    layer1_outputs(6696) <= '1';
    layer1_outputs(6697) <= not (a and b);
    layer1_outputs(6698) <= not a;
    layer1_outputs(6699) <= not a;
    layer1_outputs(6700) <= b;
    layer1_outputs(6701) <= not (a and b);
    layer1_outputs(6702) <= not a or b;
    layer1_outputs(6703) <= a xor b;
    layer1_outputs(6704) <= not b;
    layer1_outputs(6705) <= not b;
    layer1_outputs(6706) <= not a;
    layer1_outputs(6707) <= not b;
    layer1_outputs(6708) <= not (a and b);
    layer1_outputs(6709) <= '1';
    layer1_outputs(6710) <= not a;
    layer1_outputs(6711) <= not (a or b);
    layer1_outputs(6712) <= not b;
    layer1_outputs(6713) <= not b or a;
    layer1_outputs(6714) <= not b or a;
    layer1_outputs(6715) <= not (a and b);
    layer1_outputs(6716) <= a or b;
    layer1_outputs(6717) <= '1';
    layer1_outputs(6718) <= a and b;
    layer1_outputs(6719) <= b and not a;
    layer1_outputs(6720) <= not a or b;
    layer1_outputs(6721) <= a and not b;
    layer1_outputs(6722) <= a and not b;
    layer1_outputs(6723) <= a and not b;
    layer1_outputs(6724) <= not a or b;
    layer1_outputs(6725) <= b;
    layer1_outputs(6726) <= '0';
    layer1_outputs(6727) <= not (a xor b);
    layer1_outputs(6728) <= not a or b;
    layer1_outputs(6729) <= a and b;
    layer1_outputs(6730) <= '1';
    layer1_outputs(6731) <= b;
    layer1_outputs(6732) <= b;
    layer1_outputs(6733) <= a;
    layer1_outputs(6734) <= a and b;
    layer1_outputs(6735) <= a and b;
    layer1_outputs(6736) <= not a;
    layer1_outputs(6737) <= b and not a;
    layer1_outputs(6738) <= '1';
    layer1_outputs(6739) <= not b or a;
    layer1_outputs(6740) <= a and not b;
    layer1_outputs(6741) <= a and b;
    layer1_outputs(6742) <= a or b;
    layer1_outputs(6743) <= a or b;
    layer1_outputs(6744) <= not a;
    layer1_outputs(6745) <= b and not a;
    layer1_outputs(6746) <= a xor b;
    layer1_outputs(6747) <= not a;
    layer1_outputs(6748) <= not a;
    layer1_outputs(6749) <= b;
    layer1_outputs(6750) <= not (a and b);
    layer1_outputs(6751) <= a;
    layer1_outputs(6752) <= b;
    layer1_outputs(6753) <= a xor b;
    layer1_outputs(6754) <= '0';
    layer1_outputs(6755) <= not b;
    layer1_outputs(6756) <= not b;
    layer1_outputs(6757) <= b;
    layer1_outputs(6758) <= a and not b;
    layer1_outputs(6759) <= not b or a;
    layer1_outputs(6760) <= b and not a;
    layer1_outputs(6761) <= a or b;
    layer1_outputs(6762) <= '0';
    layer1_outputs(6763) <= not a;
    layer1_outputs(6764) <= not b;
    layer1_outputs(6765) <= b;
    layer1_outputs(6766) <= not (a and b);
    layer1_outputs(6767) <= a and b;
    layer1_outputs(6768) <= not (a and b);
    layer1_outputs(6769) <= b;
    layer1_outputs(6770) <= b;
    layer1_outputs(6771) <= not (a and b);
    layer1_outputs(6772) <= not a or b;
    layer1_outputs(6773) <= '0';
    layer1_outputs(6774) <= a;
    layer1_outputs(6775) <= a;
    layer1_outputs(6776) <= b;
    layer1_outputs(6777) <= a;
    layer1_outputs(6778) <= b;
    layer1_outputs(6779) <= a and b;
    layer1_outputs(6780) <= not (a or b);
    layer1_outputs(6781) <= not a;
    layer1_outputs(6782) <= a and not b;
    layer1_outputs(6783) <= '0';
    layer1_outputs(6784) <= not (a xor b);
    layer1_outputs(6785) <= not (a xor b);
    layer1_outputs(6786) <= '1';
    layer1_outputs(6787) <= not b;
    layer1_outputs(6788) <= a or b;
    layer1_outputs(6789) <= a;
    layer1_outputs(6790) <= a xor b;
    layer1_outputs(6791) <= not a or b;
    layer1_outputs(6792) <= a;
    layer1_outputs(6793) <= '0';
    layer1_outputs(6794) <= b and not a;
    layer1_outputs(6795) <= not (a and b);
    layer1_outputs(6796) <= a;
    layer1_outputs(6797) <= not b;
    layer1_outputs(6798) <= a;
    layer1_outputs(6799) <= a or b;
    layer1_outputs(6800) <= b and not a;
    layer1_outputs(6801) <= not b;
    layer1_outputs(6802) <= b;
    layer1_outputs(6803) <= not b or a;
    layer1_outputs(6804) <= not b or a;
    layer1_outputs(6805) <= not (a xor b);
    layer1_outputs(6806) <= not b;
    layer1_outputs(6807) <= b and not a;
    layer1_outputs(6808) <= b and not a;
    layer1_outputs(6809) <= '1';
    layer1_outputs(6810) <= not (a or b);
    layer1_outputs(6811) <= not b or a;
    layer1_outputs(6812) <= not (a and b);
    layer1_outputs(6813) <= not a;
    layer1_outputs(6814) <= a or b;
    layer1_outputs(6815) <= not b or a;
    layer1_outputs(6816) <= a and not b;
    layer1_outputs(6817) <= not a or b;
    layer1_outputs(6818) <= '0';
    layer1_outputs(6819) <= a and not b;
    layer1_outputs(6820) <= not a or b;
    layer1_outputs(6821) <= b and not a;
    layer1_outputs(6822) <= a and b;
    layer1_outputs(6823) <= not (a or b);
    layer1_outputs(6824) <= a;
    layer1_outputs(6825) <= not b;
    layer1_outputs(6826) <= a and not b;
    layer1_outputs(6827) <= a and b;
    layer1_outputs(6828) <= a and not b;
    layer1_outputs(6829) <= a;
    layer1_outputs(6830) <= not a;
    layer1_outputs(6831) <= a;
    layer1_outputs(6832) <= not b or a;
    layer1_outputs(6833) <= a xor b;
    layer1_outputs(6834) <= '1';
    layer1_outputs(6835) <= not b;
    layer1_outputs(6836) <= not b;
    layer1_outputs(6837) <= a and not b;
    layer1_outputs(6838) <= a and not b;
    layer1_outputs(6839) <= a;
    layer1_outputs(6840) <= b;
    layer1_outputs(6841) <= not (a or b);
    layer1_outputs(6842) <= b and not a;
    layer1_outputs(6843) <= not b or a;
    layer1_outputs(6844) <= b;
    layer1_outputs(6845) <= a and b;
    layer1_outputs(6846) <= not b;
    layer1_outputs(6847) <= not (a xor b);
    layer1_outputs(6848) <= a or b;
    layer1_outputs(6849) <= a;
    layer1_outputs(6850) <= b;
    layer1_outputs(6851) <= '1';
    layer1_outputs(6852) <= not (a and b);
    layer1_outputs(6853) <= '0';
    layer1_outputs(6854) <= not (a and b);
    layer1_outputs(6855) <= a and b;
    layer1_outputs(6856) <= not (a and b);
    layer1_outputs(6857) <= not (a and b);
    layer1_outputs(6858) <= not (a xor b);
    layer1_outputs(6859) <= '0';
    layer1_outputs(6860) <= not b;
    layer1_outputs(6861) <= a or b;
    layer1_outputs(6862) <= not (a xor b);
    layer1_outputs(6863) <= not (a and b);
    layer1_outputs(6864) <= not (a and b);
    layer1_outputs(6865) <= not b;
    layer1_outputs(6866) <= '0';
    layer1_outputs(6867) <= a and b;
    layer1_outputs(6868) <= '1';
    layer1_outputs(6869) <= not b or a;
    layer1_outputs(6870) <= '0';
    layer1_outputs(6871) <= not (a or b);
    layer1_outputs(6872) <= a xor b;
    layer1_outputs(6873) <= a and b;
    layer1_outputs(6874) <= not a or b;
    layer1_outputs(6875) <= '1';
    layer1_outputs(6876) <= a and b;
    layer1_outputs(6877) <= not b;
    layer1_outputs(6878) <= not a;
    layer1_outputs(6879) <= a and not b;
    layer1_outputs(6880) <= not (a or b);
    layer1_outputs(6881) <= not b or a;
    layer1_outputs(6882) <= b and not a;
    layer1_outputs(6883) <= not a;
    layer1_outputs(6884) <= '0';
    layer1_outputs(6885) <= not b or a;
    layer1_outputs(6886) <= '1';
    layer1_outputs(6887) <= not a or b;
    layer1_outputs(6888) <= '0';
    layer1_outputs(6889) <= not a;
    layer1_outputs(6890) <= b;
    layer1_outputs(6891) <= b;
    layer1_outputs(6892) <= '0';
    layer1_outputs(6893) <= a;
    layer1_outputs(6894) <= not b or a;
    layer1_outputs(6895) <= a or b;
    layer1_outputs(6896) <= not (a and b);
    layer1_outputs(6897) <= '0';
    layer1_outputs(6898) <= '1';
    layer1_outputs(6899) <= not (a and b);
    layer1_outputs(6900) <= b;
    layer1_outputs(6901) <= a and b;
    layer1_outputs(6902) <= '1';
    layer1_outputs(6903) <= '0';
    layer1_outputs(6904) <= not (a xor b);
    layer1_outputs(6905) <= not (a or b);
    layer1_outputs(6906) <= '1';
    layer1_outputs(6907) <= b and not a;
    layer1_outputs(6908) <= not (a and b);
    layer1_outputs(6909) <= a or b;
    layer1_outputs(6910) <= not (a and b);
    layer1_outputs(6911) <= a;
    layer1_outputs(6912) <= not b;
    layer1_outputs(6913) <= not a;
    layer1_outputs(6914) <= not b or a;
    layer1_outputs(6915) <= not a or b;
    layer1_outputs(6916) <= not (a or b);
    layer1_outputs(6917) <= not b or a;
    layer1_outputs(6918) <= not (a and b);
    layer1_outputs(6919) <= not a or b;
    layer1_outputs(6920) <= a and b;
    layer1_outputs(6921) <= not (a and b);
    layer1_outputs(6922) <= b and not a;
    layer1_outputs(6923) <= not b;
    layer1_outputs(6924) <= a or b;
    layer1_outputs(6925) <= a and not b;
    layer1_outputs(6926) <= not b;
    layer1_outputs(6927) <= a;
    layer1_outputs(6928) <= not a or b;
    layer1_outputs(6929) <= not a or b;
    layer1_outputs(6930) <= '1';
    layer1_outputs(6931) <= a xor b;
    layer1_outputs(6932) <= not b;
    layer1_outputs(6933) <= a or b;
    layer1_outputs(6934) <= '0';
    layer1_outputs(6935) <= b;
    layer1_outputs(6936) <= a xor b;
    layer1_outputs(6937) <= not a or b;
    layer1_outputs(6938) <= '0';
    layer1_outputs(6939) <= '0';
    layer1_outputs(6940) <= not a or b;
    layer1_outputs(6941) <= b and not a;
    layer1_outputs(6942) <= b;
    layer1_outputs(6943) <= a or b;
    layer1_outputs(6944) <= a or b;
    layer1_outputs(6945) <= not (a xor b);
    layer1_outputs(6946) <= not b or a;
    layer1_outputs(6947) <= not b;
    layer1_outputs(6948) <= b;
    layer1_outputs(6949) <= a and not b;
    layer1_outputs(6950) <= b;
    layer1_outputs(6951) <= not a;
    layer1_outputs(6952) <= '1';
    layer1_outputs(6953) <= not (a or b);
    layer1_outputs(6954) <= a;
    layer1_outputs(6955) <= '0';
    layer1_outputs(6956) <= not b or a;
    layer1_outputs(6957) <= not a;
    layer1_outputs(6958) <= a;
    layer1_outputs(6959) <= a;
    layer1_outputs(6960) <= b and not a;
    layer1_outputs(6961) <= not a;
    layer1_outputs(6962) <= not b;
    layer1_outputs(6963) <= a and not b;
    layer1_outputs(6964) <= a and not b;
    layer1_outputs(6965) <= b;
    layer1_outputs(6966) <= not a;
    layer1_outputs(6967) <= not a or b;
    layer1_outputs(6968) <= not (a xor b);
    layer1_outputs(6969) <= not a;
    layer1_outputs(6970) <= a and b;
    layer1_outputs(6971) <= not a;
    layer1_outputs(6972) <= not (a and b);
    layer1_outputs(6973) <= '1';
    layer1_outputs(6974) <= not a or b;
    layer1_outputs(6975) <= a or b;
    layer1_outputs(6976) <= '0';
    layer1_outputs(6977) <= not a or b;
    layer1_outputs(6978) <= not (a or b);
    layer1_outputs(6979) <= not a or b;
    layer1_outputs(6980) <= a and b;
    layer1_outputs(6981) <= not a or b;
    layer1_outputs(6982) <= a xor b;
    layer1_outputs(6983) <= a or b;
    layer1_outputs(6984) <= a;
    layer1_outputs(6985) <= not a or b;
    layer1_outputs(6986) <= '0';
    layer1_outputs(6987) <= a and not b;
    layer1_outputs(6988) <= not b or a;
    layer1_outputs(6989) <= a and b;
    layer1_outputs(6990) <= a;
    layer1_outputs(6991) <= a and b;
    layer1_outputs(6992) <= a or b;
    layer1_outputs(6993) <= not b or a;
    layer1_outputs(6994) <= not b or a;
    layer1_outputs(6995) <= a and b;
    layer1_outputs(6996) <= not (a or b);
    layer1_outputs(6997) <= a xor b;
    layer1_outputs(6998) <= b;
    layer1_outputs(6999) <= not b;
    layer1_outputs(7000) <= a;
    layer1_outputs(7001) <= not a;
    layer1_outputs(7002) <= not (a xor b);
    layer1_outputs(7003) <= not a or b;
    layer1_outputs(7004) <= a and b;
    layer1_outputs(7005) <= not a;
    layer1_outputs(7006) <= not (a and b);
    layer1_outputs(7007) <= not a;
    layer1_outputs(7008) <= a;
    layer1_outputs(7009) <= a;
    layer1_outputs(7010) <= not (a and b);
    layer1_outputs(7011) <= a or b;
    layer1_outputs(7012) <= '1';
    layer1_outputs(7013) <= a or b;
    layer1_outputs(7014) <= a xor b;
    layer1_outputs(7015) <= not a;
    layer1_outputs(7016) <= '0';
    layer1_outputs(7017) <= not (a and b);
    layer1_outputs(7018) <= a and not b;
    layer1_outputs(7019) <= not b;
    layer1_outputs(7020) <= not (a and b);
    layer1_outputs(7021) <= a or b;
    layer1_outputs(7022) <= b;
    layer1_outputs(7023) <= not (a or b);
    layer1_outputs(7024) <= a;
    layer1_outputs(7025) <= not a;
    layer1_outputs(7026) <= a and b;
    layer1_outputs(7027) <= a or b;
    layer1_outputs(7028) <= not (a or b);
    layer1_outputs(7029) <= a;
    layer1_outputs(7030) <= not (a or b);
    layer1_outputs(7031) <= not a;
    layer1_outputs(7032) <= a;
    layer1_outputs(7033) <= a or b;
    layer1_outputs(7034) <= b;
    layer1_outputs(7035) <= '0';
    layer1_outputs(7036) <= b;
    layer1_outputs(7037) <= b;
    layer1_outputs(7038) <= '1';
    layer1_outputs(7039) <= b and not a;
    layer1_outputs(7040) <= not a or b;
    layer1_outputs(7041) <= a;
    layer1_outputs(7042) <= b;
    layer1_outputs(7043) <= a or b;
    layer1_outputs(7044) <= '0';
    layer1_outputs(7045) <= '0';
    layer1_outputs(7046) <= '0';
    layer1_outputs(7047) <= '0';
    layer1_outputs(7048) <= not b or a;
    layer1_outputs(7049) <= a or b;
    layer1_outputs(7050) <= not b;
    layer1_outputs(7051) <= b;
    layer1_outputs(7052) <= not a or b;
    layer1_outputs(7053) <= '1';
    layer1_outputs(7054) <= not (a or b);
    layer1_outputs(7055) <= not a or b;
    layer1_outputs(7056) <= not a;
    layer1_outputs(7057) <= a and b;
    layer1_outputs(7058) <= not (a or b);
    layer1_outputs(7059) <= not b or a;
    layer1_outputs(7060) <= not a;
    layer1_outputs(7061) <= not a;
    layer1_outputs(7062) <= not b;
    layer1_outputs(7063) <= not (a or b);
    layer1_outputs(7064) <= not b or a;
    layer1_outputs(7065) <= not a or b;
    layer1_outputs(7066) <= not (a and b);
    layer1_outputs(7067) <= a and b;
    layer1_outputs(7068) <= '0';
    layer1_outputs(7069) <= not (a and b);
    layer1_outputs(7070) <= not b or a;
    layer1_outputs(7071) <= not (a or b);
    layer1_outputs(7072) <= not (a or b);
    layer1_outputs(7073) <= b and not a;
    layer1_outputs(7074) <= a;
    layer1_outputs(7075) <= not (a and b);
    layer1_outputs(7076) <= not b;
    layer1_outputs(7077) <= not a;
    layer1_outputs(7078) <= '1';
    layer1_outputs(7079) <= not (a xor b);
    layer1_outputs(7080) <= a;
    layer1_outputs(7081) <= not (a or b);
    layer1_outputs(7082) <= b;
    layer1_outputs(7083) <= not (a or b);
    layer1_outputs(7084) <= b;
    layer1_outputs(7085) <= not b;
    layer1_outputs(7086) <= not b;
    layer1_outputs(7087) <= not b;
    layer1_outputs(7088) <= b;
    layer1_outputs(7089) <= not (a xor b);
    layer1_outputs(7090) <= '0';
    layer1_outputs(7091) <= '1';
    layer1_outputs(7092) <= '0';
    layer1_outputs(7093) <= a and not b;
    layer1_outputs(7094) <= not (a xor b);
    layer1_outputs(7095) <= a xor b;
    layer1_outputs(7096) <= not b;
    layer1_outputs(7097) <= a and not b;
    layer1_outputs(7098) <= a;
    layer1_outputs(7099) <= a or b;
    layer1_outputs(7100) <= not b;
    layer1_outputs(7101) <= '0';
    layer1_outputs(7102) <= b;
    layer1_outputs(7103) <= not b;
    layer1_outputs(7104) <= not a;
    layer1_outputs(7105) <= a or b;
    layer1_outputs(7106) <= a and b;
    layer1_outputs(7107) <= not a;
    layer1_outputs(7108) <= not a;
    layer1_outputs(7109) <= not a;
    layer1_outputs(7110) <= not b or a;
    layer1_outputs(7111) <= a or b;
    layer1_outputs(7112) <= not b;
    layer1_outputs(7113) <= b and not a;
    layer1_outputs(7114) <= not a;
    layer1_outputs(7115) <= not a;
    layer1_outputs(7116) <= not (a or b);
    layer1_outputs(7117) <= not b;
    layer1_outputs(7118) <= a and b;
    layer1_outputs(7119) <= not b;
    layer1_outputs(7120) <= not (a and b);
    layer1_outputs(7121) <= a;
    layer1_outputs(7122) <= not b;
    layer1_outputs(7123) <= not a;
    layer1_outputs(7124) <= '1';
    layer1_outputs(7125) <= a;
    layer1_outputs(7126) <= not b;
    layer1_outputs(7127) <= b and not a;
    layer1_outputs(7128) <= a and not b;
    layer1_outputs(7129) <= not (a or b);
    layer1_outputs(7130) <= b and not a;
    layer1_outputs(7131) <= not a or b;
    layer1_outputs(7132) <= not (a and b);
    layer1_outputs(7133) <= not b;
    layer1_outputs(7134) <= b;
    layer1_outputs(7135) <= not (a or b);
    layer1_outputs(7136) <= b and not a;
    layer1_outputs(7137) <= a xor b;
    layer1_outputs(7138) <= a and not b;
    layer1_outputs(7139) <= a or b;
    layer1_outputs(7140) <= a xor b;
    layer1_outputs(7141) <= '0';
    layer1_outputs(7142) <= not (a and b);
    layer1_outputs(7143) <= not (a or b);
    layer1_outputs(7144) <= not b or a;
    layer1_outputs(7145) <= not (a or b);
    layer1_outputs(7146) <= not a;
    layer1_outputs(7147) <= not b;
    layer1_outputs(7148) <= a and b;
    layer1_outputs(7149) <= not a or b;
    layer1_outputs(7150) <= '1';
    layer1_outputs(7151) <= not a;
    layer1_outputs(7152) <= b and not a;
    layer1_outputs(7153) <= not a or b;
    layer1_outputs(7154) <= a xor b;
    layer1_outputs(7155) <= not a;
    layer1_outputs(7156) <= b;
    layer1_outputs(7157) <= not a or b;
    layer1_outputs(7158) <= not (a xor b);
    layer1_outputs(7159) <= not (a or b);
    layer1_outputs(7160) <= not a or b;
    layer1_outputs(7161) <= a and b;
    layer1_outputs(7162) <= a or b;
    layer1_outputs(7163) <= not a;
    layer1_outputs(7164) <= not a or b;
    layer1_outputs(7165) <= not a;
    layer1_outputs(7166) <= not b or a;
    layer1_outputs(7167) <= b;
    layer1_outputs(7168) <= a;
    layer1_outputs(7169) <= a or b;
    layer1_outputs(7170) <= not b;
    layer1_outputs(7171) <= not (a xor b);
    layer1_outputs(7172) <= not a or b;
    layer1_outputs(7173) <= a;
    layer1_outputs(7174) <= not (a or b);
    layer1_outputs(7175) <= not b;
    layer1_outputs(7176) <= not b;
    layer1_outputs(7177) <= a and b;
    layer1_outputs(7178) <= a and not b;
    layer1_outputs(7179) <= not (a and b);
    layer1_outputs(7180) <= not b;
    layer1_outputs(7181) <= a and b;
    layer1_outputs(7182) <= not b;
    layer1_outputs(7183) <= not (a xor b);
    layer1_outputs(7184) <= not (a or b);
    layer1_outputs(7185) <= b;
    layer1_outputs(7186) <= a and not b;
    layer1_outputs(7187) <= not b or a;
    layer1_outputs(7188) <= a and not b;
    layer1_outputs(7189) <= a or b;
    layer1_outputs(7190) <= b;
    layer1_outputs(7191) <= not a;
    layer1_outputs(7192) <= a or b;
    layer1_outputs(7193) <= not a or b;
    layer1_outputs(7194) <= b;
    layer1_outputs(7195) <= a and not b;
    layer1_outputs(7196) <= a;
    layer1_outputs(7197) <= a or b;
    layer1_outputs(7198) <= a;
    layer1_outputs(7199) <= a or b;
    layer1_outputs(7200) <= a or b;
    layer1_outputs(7201) <= not a or b;
    layer1_outputs(7202) <= a or b;
    layer1_outputs(7203) <= not (a or b);
    layer1_outputs(7204) <= a and b;
    layer1_outputs(7205) <= not b or a;
    layer1_outputs(7206) <= b;
    layer1_outputs(7207) <= a or b;
    layer1_outputs(7208) <= '1';
    layer1_outputs(7209) <= not (a or b);
    layer1_outputs(7210) <= a;
    layer1_outputs(7211) <= not b or a;
    layer1_outputs(7212) <= a or b;
    layer1_outputs(7213) <= b and not a;
    layer1_outputs(7214) <= '0';
    layer1_outputs(7215) <= a and b;
    layer1_outputs(7216) <= not (a xor b);
    layer1_outputs(7217) <= b;
    layer1_outputs(7218) <= b and not a;
    layer1_outputs(7219) <= not a;
    layer1_outputs(7220) <= b and not a;
    layer1_outputs(7221) <= a;
    layer1_outputs(7222) <= b and not a;
    layer1_outputs(7223) <= b;
    layer1_outputs(7224) <= not (a and b);
    layer1_outputs(7225) <= not (a xor b);
    layer1_outputs(7226) <= '1';
    layer1_outputs(7227) <= not (a and b);
    layer1_outputs(7228) <= not (a or b);
    layer1_outputs(7229) <= '0';
    layer1_outputs(7230) <= not b;
    layer1_outputs(7231) <= a or b;
    layer1_outputs(7232) <= a;
    layer1_outputs(7233) <= not a;
    layer1_outputs(7234) <= a or b;
    layer1_outputs(7235) <= a and not b;
    layer1_outputs(7236) <= not a;
    layer1_outputs(7237) <= '0';
    layer1_outputs(7238) <= not a;
    layer1_outputs(7239) <= a and b;
    layer1_outputs(7240) <= not a or b;
    layer1_outputs(7241) <= not (a or b);
    layer1_outputs(7242) <= '1';
    layer1_outputs(7243) <= a or b;
    layer1_outputs(7244) <= b;
    layer1_outputs(7245) <= not (a and b);
    layer1_outputs(7246) <= b and not a;
    layer1_outputs(7247) <= b;
    layer1_outputs(7248) <= a xor b;
    layer1_outputs(7249) <= a and not b;
    layer1_outputs(7250) <= not b or a;
    layer1_outputs(7251) <= a;
    layer1_outputs(7252) <= a xor b;
    layer1_outputs(7253) <= not (a xor b);
    layer1_outputs(7254) <= b;
    layer1_outputs(7255) <= '1';
    layer1_outputs(7256) <= not b;
    layer1_outputs(7257) <= not b;
    layer1_outputs(7258) <= not b;
    layer1_outputs(7259) <= a;
    layer1_outputs(7260) <= '0';
    layer1_outputs(7261) <= b;
    layer1_outputs(7262) <= not b;
    layer1_outputs(7263) <= not (a and b);
    layer1_outputs(7264) <= '0';
    layer1_outputs(7265) <= '1';
    layer1_outputs(7266) <= not a or b;
    layer1_outputs(7267) <= not (a or b);
    layer1_outputs(7268) <= '0';
    layer1_outputs(7269) <= '0';
    layer1_outputs(7270) <= not a;
    layer1_outputs(7271) <= a and b;
    layer1_outputs(7272) <= a xor b;
    layer1_outputs(7273) <= a;
    layer1_outputs(7274) <= not a;
    layer1_outputs(7275) <= not (a or b);
    layer1_outputs(7276) <= a;
    layer1_outputs(7277) <= a and b;
    layer1_outputs(7278) <= a and b;
    layer1_outputs(7279) <= '0';
    layer1_outputs(7280) <= a and not b;
    layer1_outputs(7281) <= not a;
    layer1_outputs(7282) <= b and not a;
    layer1_outputs(7283) <= not b;
    layer1_outputs(7284) <= a and b;
    layer1_outputs(7285) <= '1';
    layer1_outputs(7286) <= b and not a;
    layer1_outputs(7287) <= not b or a;
    layer1_outputs(7288) <= b and not a;
    layer1_outputs(7289) <= not a;
    layer1_outputs(7290) <= a and not b;
    layer1_outputs(7291) <= a;
    layer1_outputs(7292) <= not a;
    layer1_outputs(7293) <= not (a or b);
    layer1_outputs(7294) <= a or b;
    layer1_outputs(7295) <= b and not a;
    layer1_outputs(7296) <= '0';
    layer1_outputs(7297) <= a or b;
    layer1_outputs(7298) <= not b;
    layer1_outputs(7299) <= not (a xor b);
    layer1_outputs(7300) <= '1';
    layer1_outputs(7301) <= a and not b;
    layer1_outputs(7302) <= not b;
    layer1_outputs(7303) <= not (a or b);
    layer1_outputs(7304) <= not b;
    layer1_outputs(7305) <= a;
    layer1_outputs(7306) <= a;
    layer1_outputs(7307) <= '0';
    layer1_outputs(7308) <= b;
    layer1_outputs(7309) <= '1';
    layer1_outputs(7310) <= not a or b;
    layer1_outputs(7311) <= b and not a;
    layer1_outputs(7312) <= not a;
    layer1_outputs(7313) <= a or b;
    layer1_outputs(7314) <= not (a or b);
    layer1_outputs(7315) <= not b;
    layer1_outputs(7316) <= a;
    layer1_outputs(7317) <= a;
    layer1_outputs(7318) <= a and b;
    layer1_outputs(7319) <= not a or b;
    layer1_outputs(7320) <= '0';
    layer1_outputs(7321) <= not a;
    layer1_outputs(7322) <= a or b;
    layer1_outputs(7323) <= a and not b;
    layer1_outputs(7324) <= a xor b;
    layer1_outputs(7325) <= not a or b;
    layer1_outputs(7326) <= a xor b;
    layer1_outputs(7327) <= not a or b;
    layer1_outputs(7328) <= a or b;
    layer1_outputs(7329) <= '1';
    layer1_outputs(7330) <= a and not b;
    layer1_outputs(7331) <= b;
    layer1_outputs(7332) <= not (a and b);
    layer1_outputs(7333) <= a and b;
    layer1_outputs(7334) <= not (a or b);
    layer1_outputs(7335) <= a;
    layer1_outputs(7336) <= not b;
    layer1_outputs(7337) <= b;
    layer1_outputs(7338) <= a and not b;
    layer1_outputs(7339) <= not (a xor b);
    layer1_outputs(7340) <= not (a or b);
    layer1_outputs(7341) <= not a;
    layer1_outputs(7342) <= not (a xor b);
    layer1_outputs(7343) <= not (a xor b);
    layer1_outputs(7344) <= a;
    layer1_outputs(7345) <= a;
    layer1_outputs(7346) <= a;
    layer1_outputs(7347) <= not b;
    layer1_outputs(7348) <= not a or b;
    layer1_outputs(7349) <= a and not b;
    layer1_outputs(7350) <= not b;
    layer1_outputs(7351) <= not (a or b);
    layer1_outputs(7352) <= '0';
    layer1_outputs(7353) <= a or b;
    layer1_outputs(7354) <= not (a and b);
    layer1_outputs(7355) <= '1';
    layer1_outputs(7356) <= not b or a;
    layer1_outputs(7357) <= not a;
    layer1_outputs(7358) <= not (a and b);
    layer1_outputs(7359) <= '0';
    layer1_outputs(7360) <= b;
    layer1_outputs(7361) <= not (a or b);
    layer1_outputs(7362) <= not (a xor b);
    layer1_outputs(7363) <= b;
    layer1_outputs(7364) <= not a;
    layer1_outputs(7365) <= '1';
    layer1_outputs(7366) <= '0';
    layer1_outputs(7367) <= a and b;
    layer1_outputs(7368) <= '0';
    layer1_outputs(7369) <= a and b;
    layer1_outputs(7370) <= not a;
    layer1_outputs(7371) <= a;
    layer1_outputs(7372) <= a and not b;
    layer1_outputs(7373) <= not b or a;
    layer1_outputs(7374) <= not (a or b);
    layer1_outputs(7375) <= not a or b;
    layer1_outputs(7376) <= a and not b;
    layer1_outputs(7377) <= a and not b;
    layer1_outputs(7378) <= a or b;
    layer1_outputs(7379) <= a xor b;
    layer1_outputs(7380) <= b and not a;
    layer1_outputs(7381) <= not b or a;
    layer1_outputs(7382) <= b;
    layer1_outputs(7383) <= not a or b;
    layer1_outputs(7384) <= a;
    layer1_outputs(7385) <= a;
    layer1_outputs(7386) <= not (a or b);
    layer1_outputs(7387) <= '1';
    layer1_outputs(7388) <= not a or b;
    layer1_outputs(7389) <= a and not b;
    layer1_outputs(7390) <= a and not b;
    layer1_outputs(7391) <= a and not b;
    layer1_outputs(7392) <= a or b;
    layer1_outputs(7393) <= a and not b;
    layer1_outputs(7394) <= not (a and b);
    layer1_outputs(7395) <= a and not b;
    layer1_outputs(7396) <= a xor b;
    layer1_outputs(7397) <= a xor b;
    layer1_outputs(7398) <= a or b;
    layer1_outputs(7399) <= '0';
    layer1_outputs(7400) <= b;
    layer1_outputs(7401) <= '1';
    layer1_outputs(7402) <= a and b;
    layer1_outputs(7403) <= '0';
    layer1_outputs(7404) <= a and not b;
    layer1_outputs(7405) <= not (a and b);
    layer1_outputs(7406) <= not (a or b);
    layer1_outputs(7407) <= a and b;
    layer1_outputs(7408) <= a;
    layer1_outputs(7409) <= not a;
    layer1_outputs(7410) <= '0';
    layer1_outputs(7411) <= not (a and b);
    layer1_outputs(7412) <= a or b;
    layer1_outputs(7413) <= not (a or b);
    layer1_outputs(7414) <= not a;
    layer1_outputs(7415) <= not (a and b);
    layer1_outputs(7416) <= not a;
    layer1_outputs(7417) <= not b or a;
    layer1_outputs(7418) <= '0';
    layer1_outputs(7419) <= a;
    layer1_outputs(7420) <= not (a xor b);
    layer1_outputs(7421) <= not a;
    layer1_outputs(7422) <= not (a xor b);
    layer1_outputs(7423) <= '1';
    layer1_outputs(7424) <= not (a xor b);
    layer1_outputs(7425) <= a;
    layer1_outputs(7426) <= not b;
    layer1_outputs(7427) <= '1';
    layer1_outputs(7428) <= a;
    layer1_outputs(7429) <= not b;
    layer1_outputs(7430) <= not (a and b);
    layer1_outputs(7431) <= not (a xor b);
    layer1_outputs(7432) <= '0';
    layer1_outputs(7433) <= b;
    layer1_outputs(7434) <= not b;
    layer1_outputs(7435) <= b and not a;
    layer1_outputs(7436) <= not b or a;
    layer1_outputs(7437) <= a and b;
    layer1_outputs(7438) <= a;
    layer1_outputs(7439) <= b;
    layer1_outputs(7440) <= b and not a;
    layer1_outputs(7441) <= b and not a;
    layer1_outputs(7442) <= not a or b;
    layer1_outputs(7443) <= not a;
    layer1_outputs(7444) <= not a or b;
    layer1_outputs(7445) <= not b;
    layer1_outputs(7446) <= b and not a;
    layer1_outputs(7447) <= b and not a;
    layer1_outputs(7448) <= not b or a;
    layer1_outputs(7449) <= b;
    layer1_outputs(7450) <= not a or b;
    layer1_outputs(7451) <= '1';
    layer1_outputs(7452) <= b and not a;
    layer1_outputs(7453) <= not (a xor b);
    layer1_outputs(7454) <= a and b;
    layer1_outputs(7455) <= a and not b;
    layer1_outputs(7456) <= a;
    layer1_outputs(7457) <= a and not b;
    layer1_outputs(7458) <= not a;
    layer1_outputs(7459) <= not b or a;
    layer1_outputs(7460) <= not (a and b);
    layer1_outputs(7461) <= b and not a;
    layer1_outputs(7462) <= not a;
    layer1_outputs(7463) <= '0';
    layer1_outputs(7464) <= not (a or b);
    layer1_outputs(7465) <= '0';
    layer1_outputs(7466) <= a;
    layer1_outputs(7467) <= not b or a;
    layer1_outputs(7468) <= '1';
    layer1_outputs(7469) <= a;
    layer1_outputs(7470) <= a and b;
    layer1_outputs(7471) <= not b;
    layer1_outputs(7472) <= not b;
    layer1_outputs(7473) <= not b;
    layer1_outputs(7474) <= b and not a;
    layer1_outputs(7475) <= not (a or b);
    layer1_outputs(7476) <= b and not a;
    layer1_outputs(7477) <= not (a or b);
    layer1_outputs(7478) <= '1';
    layer1_outputs(7479) <= b and not a;
    layer1_outputs(7480) <= a;
    layer1_outputs(7481) <= '1';
    layer1_outputs(7482) <= a or b;
    layer1_outputs(7483) <= not a;
    layer1_outputs(7484) <= not (a or b);
    layer1_outputs(7485) <= a or b;
    layer1_outputs(7486) <= b;
    layer1_outputs(7487) <= a and not b;
    layer1_outputs(7488) <= a;
    layer1_outputs(7489) <= not (a xor b);
    layer1_outputs(7490) <= not b;
    layer1_outputs(7491) <= not b or a;
    layer1_outputs(7492) <= not b;
    layer1_outputs(7493) <= b and not a;
    layer1_outputs(7494) <= b;
    layer1_outputs(7495) <= a;
    layer1_outputs(7496) <= not b;
    layer1_outputs(7497) <= '1';
    layer1_outputs(7498) <= '0';
    layer1_outputs(7499) <= not a or b;
    layer1_outputs(7500) <= '1';
    layer1_outputs(7501) <= not b or a;
    layer1_outputs(7502) <= not (a or b);
    layer1_outputs(7503) <= a;
    layer1_outputs(7504) <= not a;
    layer1_outputs(7505) <= a or b;
    layer1_outputs(7506) <= '0';
    layer1_outputs(7507) <= a and b;
    layer1_outputs(7508) <= not (a and b);
    layer1_outputs(7509) <= '1';
    layer1_outputs(7510) <= not a;
    layer1_outputs(7511) <= not (a and b);
    layer1_outputs(7512) <= not (a or b);
    layer1_outputs(7513) <= a and not b;
    layer1_outputs(7514) <= not b or a;
    layer1_outputs(7515) <= '1';
    layer1_outputs(7516) <= b and not a;
    layer1_outputs(7517) <= b;
    layer1_outputs(7518) <= not a or b;
    layer1_outputs(7519) <= not (a xor b);
    layer1_outputs(7520) <= a and b;
    layer1_outputs(7521) <= not b or a;
    layer1_outputs(7522) <= not (a xor b);
    layer1_outputs(7523) <= a xor b;
    layer1_outputs(7524) <= not (a or b);
    layer1_outputs(7525) <= a and b;
    layer1_outputs(7526) <= not a or b;
    layer1_outputs(7527) <= a and not b;
    layer1_outputs(7528) <= '1';
    layer1_outputs(7529) <= not (a and b);
    layer1_outputs(7530) <= not a or b;
    layer1_outputs(7531) <= '0';
    layer1_outputs(7532) <= '0';
    layer1_outputs(7533) <= b and not a;
    layer1_outputs(7534) <= b;
    layer1_outputs(7535) <= a or b;
    layer1_outputs(7536) <= not a or b;
    layer1_outputs(7537) <= a;
    layer1_outputs(7538) <= not a or b;
    layer1_outputs(7539) <= not a;
    layer1_outputs(7540) <= a;
    layer1_outputs(7541) <= not (a and b);
    layer1_outputs(7542) <= a or b;
    layer1_outputs(7543) <= not (a or b);
    layer1_outputs(7544) <= not b or a;
    layer1_outputs(7545) <= b;
    layer1_outputs(7546) <= a or b;
    layer1_outputs(7547) <= '0';
    layer1_outputs(7548) <= a and b;
    layer1_outputs(7549) <= b and not a;
    layer1_outputs(7550) <= not (a or b);
    layer1_outputs(7551) <= a xor b;
    layer1_outputs(7552) <= b;
    layer1_outputs(7553) <= not (a or b);
    layer1_outputs(7554) <= not (a or b);
    layer1_outputs(7555) <= a;
    layer1_outputs(7556) <= a and b;
    layer1_outputs(7557) <= not b or a;
    layer1_outputs(7558) <= not a or b;
    layer1_outputs(7559) <= not a or b;
    layer1_outputs(7560) <= not a;
    layer1_outputs(7561) <= not a;
    layer1_outputs(7562) <= a or b;
    layer1_outputs(7563) <= not (a xor b);
    layer1_outputs(7564) <= not b or a;
    layer1_outputs(7565) <= a;
    layer1_outputs(7566) <= not a or b;
    layer1_outputs(7567) <= not (a and b);
    layer1_outputs(7568) <= a;
    layer1_outputs(7569) <= '0';
    layer1_outputs(7570) <= a;
    layer1_outputs(7571) <= '1';
    layer1_outputs(7572) <= not a;
    layer1_outputs(7573) <= not b;
    layer1_outputs(7574) <= '1';
    layer1_outputs(7575) <= '1';
    layer1_outputs(7576) <= b and not a;
    layer1_outputs(7577) <= not a;
    layer1_outputs(7578) <= not (a or b);
    layer1_outputs(7579) <= a and not b;
    layer1_outputs(7580) <= a and not b;
    layer1_outputs(7581) <= a or b;
    layer1_outputs(7582) <= not (a xor b);
    layer1_outputs(7583) <= not b or a;
    layer1_outputs(7584) <= a;
    layer1_outputs(7585) <= a and not b;
    layer1_outputs(7586) <= not (a or b);
    layer1_outputs(7587) <= not a;
    layer1_outputs(7588) <= not a or b;
    layer1_outputs(7589) <= a or b;
    layer1_outputs(7590) <= b and not a;
    layer1_outputs(7591) <= not b or a;
    layer1_outputs(7592) <= a or b;
    layer1_outputs(7593) <= a xor b;
    layer1_outputs(7594) <= '1';
    layer1_outputs(7595) <= not b;
    layer1_outputs(7596) <= not a;
    layer1_outputs(7597) <= a or b;
    layer1_outputs(7598) <= '0';
    layer1_outputs(7599) <= not a or b;
    layer1_outputs(7600) <= a and not b;
    layer1_outputs(7601) <= a xor b;
    layer1_outputs(7602) <= not (a and b);
    layer1_outputs(7603) <= a and not b;
    layer1_outputs(7604) <= b;
    layer1_outputs(7605) <= a;
    layer1_outputs(7606) <= '0';
    layer1_outputs(7607) <= a;
    layer1_outputs(7608) <= b and not a;
    layer1_outputs(7609) <= not (a and b);
    layer1_outputs(7610) <= a and not b;
    layer1_outputs(7611) <= b;
    layer1_outputs(7612) <= not (a or b);
    layer1_outputs(7613) <= not b;
    layer1_outputs(7614) <= not (a and b);
    layer1_outputs(7615) <= a xor b;
    layer1_outputs(7616) <= b;
    layer1_outputs(7617) <= not b or a;
    layer1_outputs(7618) <= a or b;
    layer1_outputs(7619) <= a;
    layer1_outputs(7620) <= a;
    layer1_outputs(7621) <= not b;
    layer1_outputs(7622) <= a and not b;
    layer1_outputs(7623) <= not (a or b);
    layer1_outputs(7624) <= '1';
    layer1_outputs(7625) <= not (a and b);
    layer1_outputs(7626) <= not (a or b);
    layer1_outputs(7627) <= not (a and b);
    layer1_outputs(7628) <= a;
    layer1_outputs(7629) <= not a or b;
    layer1_outputs(7630) <= a and b;
    layer1_outputs(7631) <= a or b;
    layer1_outputs(7632) <= not (a or b);
    layer1_outputs(7633) <= a;
    layer1_outputs(7634) <= b and not a;
    layer1_outputs(7635) <= b and not a;
    layer1_outputs(7636) <= '0';
    layer1_outputs(7637) <= not b;
    layer1_outputs(7638) <= a and not b;
    layer1_outputs(7639) <= not (a and b);
    layer1_outputs(7640) <= a;
    layer1_outputs(7641) <= a and b;
    layer1_outputs(7642) <= a and not b;
    layer1_outputs(7643) <= a and b;
    layer1_outputs(7644) <= a and not b;
    layer1_outputs(7645) <= a or b;
    layer1_outputs(7646) <= a;
    layer1_outputs(7647) <= not b or a;
    layer1_outputs(7648) <= b and not a;
    layer1_outputs(7649) <= not b;
    layer1_outputs(7650) <= a;
    layer1_outputs(7651) <= a or b;
    layer1_outputs(7652) <= a xor b;
    layer1_outputs(7653) <= a and not b;
    layer1_outputs(7654) <= not a;
    layer1_outputs(7655) <= '1';
    layer1_outputs(7656) <= '1';
    layer1_outputs(7657) <= not a;
    layer1_outputs(7658) <= not a or b;
    layer1_outputs(7659) <= not a or b;
    layer1_outputs(7660) <= a xor b;
    layer1_outputs(7661) <= not (a and b);
    layer1_outputs(7662) <= not b or a;
    layer1_outputs(7663) <= not b or a;
    layer1_outputs(7664) <= b;
    layer1_outputs(7665) <= a;
    layer1_outputs(7666) <= '0';
    layer1_outputs(7667) <= '1';
    layer1_outputs(7668) <= not (a and b);
    layer1_outputs(7669) <= not b or a;
    layer1_outputs(7670) <= a and not b;
    layer1_outputs(7671) <= b;
    layer1_outputs(7672) <= not b;
    layer1_outputs(7673) <= not a or b;
    layer1_outputs(7674) <= '0';
    layer1_outputs(7675) <= not (a xor b);
    layer1_outputs(7676) <= b and not a;
    layer1_outputs(7677) <= b;
    layer1_outputs(7678) <= a or b;
    layer1_outputs(7679) <= not (a or b);
    layer1_outputs(7680) <= '0';
    layer1_outputs(7681) <= a or b;
    layer1_outputs(7682) <= not a;
    layer1_outputs(7683) <= not (a and b);
    layer1_outputs(7684) <= not a or b;
    layer1_outputs(7685) <= not b;
    layer1_outputs(7686) <= '0';
    layer1_outputs(7687) <= not (a and b);
    layer1_outputs(7688) <= a xor b;
    layer1_outputs(7689) <= a and b;
    layer1_outputs(7690) <= not b or a;
    layer1_outputs(7691) <= not (a xor b);
    layer1_outputs(7692) <= '1';
    layer1_outputs(7693) <= a;
    layer1_outputs(7694) <= '0';
    layer1_outputs(7695) <= not a or b;
    layer1_outputs(7696) <= not a;
    layer1_outputs(7697) <= not b;
    layer1_outputs(7698) <= not (a and b);
    layer1_outputs(7699) <= a or b;
    layer1_outputs(7700) <= a and not b;
    layer1_outputs(7701) <= a and b;
    layer1_outputs(7702) <= a and b;
    layer1_outputs(7703) <= a and b;
    layer1_outputs(7704) <= not (a xor b);
    layer1_outputs(7705) <= a and not b;
    layer1_outputs(7706) <= a;
    layer1_outputs(7707) <= '1';
    layer1_outputs(7708) <= b;
    layer1_outputs(7709) <= a or b;
    layer1_outputs(7710) <= a xor b;
    layer1_outputs(7711) <= a and not b;
    layer1_outputs(7712) <= a and not b;
    layer1_outputs(7713) <= '0';
    layer1_outputs(7714) <= not (a and b);
    layer1_outputs(7715) <= a;
    layer1_outputs(7716) <= not (a and b);
    layer1_outputs(7717) <= a and not b;
    layer1_outputs(7718) <= not (a or b);
    layer1_outputs(7719) <= a and b;
    layer1_outputs(7720) <= not a or b;
    layer1_outputs(7721) <= not a or b;
    layer1_outputs(7722) <= '0';
    layer1_outputs(7723) <= '1';
    layer1_outputs(7724) <= '1';
    layer1_outputs(7725) <= '0';
    layer1_outputs(7726) <= not a;
    layer1_outputs(7727) <= not a or b;
    layer1_outputs(7728) <= not (a and b);
    layer1_outputs(7729) <= a and b;
    layer1_outputs(7730) <= b and not a;
    layer1_outputs(7731) <= a xor b;
    layer1_outputs(7732) <= not (a xor b);
    layer1_outputs(7733) <= '0';
    layer1_outputs(7734) <= '0';
    layer1_outputs(7735) <= a xor b;
    layer1_outputs(7736) <= a and not b;
    layer1_outputs(7737) <= not (a or b);
    layer1_outputs(7738) <= not a;
    layer1_outputs(7739) <= a;
    layer1_outputs(7740) <= a and not b;
    layer1_outputs(7741) <= not a or b;
    layer1_outputs(7742) <= not (a and b);
    layer1_outputs(7743) <= not (a or b);
    layer1_outputs(7744) <= not b;
    layer1_outputs(7745) <= not (a or b);
    layer1_outputs(7746) <= a or b;
    layer1_outputs(7747) <= not (a and b);
    layer1_outputs(7748) <= a and not b;
    layer1_outputs(7749) <= not b or a;
    layer1_outputs(7750) <= not a;
    layer1_outputs(7751) <= '1';
    layer1_outputs(7752) <= not (a or b);
    layer1_outputs(7753) <= not a;
    layer1_outputs(7754) <= b;
    layer1_outputs(7755) <= not b;
    layer1_outputs(7756) <= not a;
    layer1_outputs(7757) <= b and not a;
    layer1_outputs(7758) <= not (a or b);
    layer1_outputs(7759) <= not a;
    layer1_outputs(7760) <= a and b;
    layer1_outputs(7761) <= a and not b;
    layer1_outputs(7762) <= a or b;
    layer1_outputs(7763) <= b and not a;
    layer1_outputs(7764) <= '0';
    layer1_outputs(7765) <= a and not b;
    layer1_outputs(7766) <= '0';
    layer1_outputs(7767) <= not a;
    layer1_outputs(7768) <= not (a xor b);
    layer1_outputs(7769) <= not a;
    layer1_outputs(7770) <= not b;
    layer1_outputs(7771) <= b;
    layer1_outputs(7772) <= not b;
    layer1_outputs(7773) <= not a;
    layer1_outputs(7774) <= a xor b;
    layer1_outputs(7775) <= not a or b;
    layer1_outputs(7776) <= not b or a;
    layer1_outputs(7777) <= not b;
    layer1_outputs(7778) <= not b or a;
    layer1_outputs(7779) <= b and not a;
    layer1_outputs(7780) <= a or b;
    layer1_outputs(7781) <= a and b;
    layer1_outputs(7782) <= not a or b;
    layer1_outputs(7783) <= a;
    layer1_outputs(7784) <= a or b;
    layer1_outputs(7785) <= a and not b;
    layer1_outputs(7786) <= a and not b;
    layer1_outputs(7787) <= not (a and b);
    layer1_outputs(7788) <= not a or b;
    layer1_outputs(7789) <= '1';
    layer1_outputs(7790) <= b;
    layer1_outputs(7791) <= not a or b;
    layer1_outputs(7792) <= a or b;
    layer1_outputs(7793) <= b;
    layer1_outputs(7794) <= b and not a;
    layer1_outputs(7795) <= a and not b;
    layer1_outputs(7796) <= not b;
    layer1_outputs(7797) <= '1';
    layer1_outputs(7798) <= not (a and b);
    layer1_outputs(7799) <= b and not a;
    layer1_outputs(7800) <= b and not a;
    layer1_outputs(7801) <= a;
    layer1_outputs(7802) <= not b or a;
    layer1_outputs(7803) <= not b or a;
    layer1_outputs(7804) <= not b;
    layer1_outputs(7805) <= '1';
    layer1_outputs(7806) <= a and b;
    layer1_outputs(7807) <= not b;
    layer1_outputs(7808) <= not b;
    layer1_outputs(7809) <= not a or b;
    layer1_outputs(7810) <= b;
    layer1_outputs(7811) <= not (a or b);
    layer1_outputs(7812) <= a xor b;
    layer1_outputs(7813) <= not a or b;
    layer1_outputs(7814) <= not a or b;
    layer1_outputs(7815) <= '0';
    layer1_outputs(7816) <= not a;
    layer1_outputs(7817) <= not (a and b);
    layer1_outputs(7818) <= a and b;
    layer1_outputs(7819) <= not b;
    layer1_outputs(7820) <= not b;
    layer1_outputs(7821) <= a and b;
    layer1_outputs(7822) <= b and not a;
    layer1_outputs(7823) <= not a;
    layer1_outputs(7824) <= a;
    layer1_outputs(7825) <= not a or b;
    layer1_outputs(7826) <= not (a or b);
    layer1_outputs(7827) <= not (a or b);
    layer1_outputs(7828) <= a and b;
    layer1_outputs(7829) <= a and not b;
    layer1_outputs(7830) <= a and not b;
    layer1_outputs(7831) <= not b;
    layer1_outputs(7832) <= '1';
    layer1_outputs(7833) <= not b or a;
    layer1_outputs(7834) <= not (a and b);
    layer1_outputs(7835) <= a and b;
    layer1_outputs(7836) <= not (a or b);
    layer1_outputs(7837) <= b;
    layer1_outputs(7838) <= a;
    layer1_outputs(7839) <= not b or a;
    layer1_outputs(7840) <= not b;
    layer1_outputs(7841) <= '0';
    layer1_outputs(7842) <= not (a and b);
    layer1_outputs(7843) <= not b or a;
    layer1_outputs(7844) <= a or b;
    layer1_outputs(7845) <= b and not a;
    layer1_outputs(7846) <= b;
    layer1_outputs(7847) <= a xor b;
    layer1_outputs(7848) <= a or b;
    layer1_outputs(7849) <= not b;
    layer1_outputs(7850) <= not b or a;
    layer1_outputs(7851) <= '1';
    layer1_outputs(7852) <= not a;
    layer1_outputs(7853) <= not a or b;
    layer1_outputs(7854) <= not b;
    layer1_outputs(7855) <= a;
    layer1_outputs(7856) <= not (a or b);
    layer1_outputs(7857) <= not a or b;
    layer1_outputs(7858) <= b;
    layer1_outputs(7859) <= not (a or b);
    layer1_outputs(7860) <= not b;
    layer1_outputs(7861) <= b;
    layer1_outputs(7862) <= not b or a;
    layer1_outputs(7863) <= a or b;
    layer1_outputs(7864) <= not (a xor b);
    layer1_outputs(7865) <= a;
    layer1_outputs(7866) <= not a or b;
    layer1_outputs(7867) <= a and not b;
    layer1_outputs(7868) <= not a or b;
    layer1_outputs(7869) <= a or b;
    layer1_outputs(7870) <= a and not b;
    layer1_outputs(7871) <= a and b;
    layer1_outputs(7872) <= '1';
    layer1_outputs(7873) <= not (a and b);
    layer1_outputs(7874) <= a and b;
    layer1_outputs(7875) <= not a;
    layer1_outputs(7876) <= not b or a;
    layer1_outputs(7877) <= b;
    layer1_outputs(7878) <= not b;
    layer1_outputs(7879) <= not a;
    layer1_outputs(7880) <= not b;
    layer1_outputs(7881) <= not b or a;
    layer1_outputs(7882) <= '1';
    layer1_outputs(7883) <= not a;
    layer1_outputs(7884) <= a;
    layer1_outputs(7885) <= not a;
    layer1_outputs(7886) <= '1';
    layer1_outputs(7887) <= a;
    layer1_outputs(7888) <= b;
    layer1_outputs(7889) <= not b or a;
    layer1_outputs(7890) <= '0';
    layer1_outputs(7891) <= '1';
    layer1_outputs(7892) <= not a;
    layer1_outputs(7893) <= a and not b;
    layer1_outputs(7894) <= b and not a;
    layer1_outputs(7895) <= a or b;
    layer1_outputs(7896) <= '1';
    layer1_outputs(7897) <= b;
    layer1_outputs(7898) <= a xor b;
    layer1_outputs(7899) <= not a;
    layer1_outputs(7900) <= not b or a;
    layer1_outputs(7901) <= '0';
    layer1_outputs(7902) <= not b or a;
    layer1_outputs(7903) <= a;
    layer1_outputs(7904) <= not b or a;
    layer1_outputs(7905) <= not b;
    layer1_outputs(7906) <= not (a xor b);
    layer1_outputs(7907) <= not (a and b);
    layer1_outputs(7908) <= '0';
    layer1_outputs(7909) <= not (a and b);
    layer1_outputs(7910) <= not (a xor b);
    layer1_outputs(7911) <= '1';
    layer1_outputs(7912) <= not b or a;
    layer1_outputs(7913) <= '1';
    layer1_outputs(7914) <= not a;
    layer1_outputs(7915) <= not b or a;
    layer1_outputs(7916) <= not a or b;
    layer1_outputs(7917) <= not b or a;
    layer1_outputs(7918) <= not a;
    layer1_outputs(7919) <= not b or a;
    layer1_outputs(7920) <= '1';
    layer1_outputs(7921) <= a;
    layer1_outputs(7922) <= not b;
    layer1_outputs(7923) <= '0';
    layer1_outputs(7924) <= b and not a;
    layer1_outputs(7925) <= a xor b;
    layer1_outputs(7926) <= not (a and b);
    layer1_outputs(7927) <= not b or a;
    layer1_outputs(7928) <= b and not a;
    layer1_outputs(7929) <= not a;
    layer1_outputs(7930) <= not a;
    layer1_outputs(7931) <= '0';
    layer1_outputs(7932) <= '0';
    layer1_outputs(7933) <= a and b;
    layer1_outputs(7934) <= not a or b;
    layer1_outputs(7935) <= b;
    layer1_outputs(7936) <= not b;
    layer1_outputs(7937) <= a xor b;
    layer1_outputs(7938) <= not (a and b);
    layer1_outputs(7939) <= not a;
    layer1_outputs(7940) <= '1';
    layer1_outputs(7941) <= b;
    layer1_outputs(7942) <= not b;
    layer1_outputs(7943) <= not a or b;
    layer1_outputs(7944) <= not (a and b);
    layer1_outputs(7945) <= not a or b;
    layer1_outputs(7946) <= not (a or b);
    layer1_outputs(7947) <= '0';
    layer1_outputs(7948) <= not a;
    layer1_outputs(7949) <= not (a or b);
    layer1_outputs(7950) <= b and not a;
    layer1_outputs(7951) <= a or b;
    layer1_outputs(7952) <= a and not b;
    layer1_outputs(7953) <= not (a xor b);
    layer1_outputs(7954) <= b and not a;
    layer1_outputs(7955) <= not a;
    layer1_outputs(7956) <= a;
    layer1_outputs(7957) <= a;
    layer1_outputs(7958) <= not (a and b);
    layer1_outputs(7959) <= not b or a;
    layer1_outputs(7960) <= not b or a;
    layer1_outputs(7961) <= b and not a;
    layer1_outputs(7962) <= '0';
    layer1_outputs(7963) <= not a;
    layer1_outputs(7964) <= '0';
    layer1_outputs(7965) <= b;
    layer1_outputs(7966) <= a and not b;
    layer1_outputs(7967) <= not b;
    layer1_outputs(7968) <= not b;
    layer1_outputs(7969) <= not a or b;
    layer1_outputs(7970) <= not a;
    layer1_outputs(7971) <= '1';
    layer1_outputs(7972) <= a and not b;
    layer1_outputs(7973) <= a;
    layer1_outputs(7974) <= not b;
    layer1_outputs(7975) <= a xor b;
    layer1_outputs(7976) <= not (a and b);
    layer1_outputs(7977) <= '0';
    layer1_outputs(7978) <= not a or b;
    layer1_outputs(7979) <= not (a and b);
    layer1_outputs(7980) <= not a or b;
    layer1_outputs(7981) <= not b;
    layer1_outputs(7982) <= a xor b;
    layer1_outputs(7983) <= not b;
    layer1_outputs(7984) <= b;
    layer1_outputs(7985) <= not a;
    layer1_outputs(7986) <= a or b;
    layer1_outputs(7987) <= not (a xor b);
    layer1_outputs(7988) <= not (a or b);
    layer1_outputs(7989) <= a and not b;
    layer1_outputs(7990) <= not a or b;
    layer1_outputs(7991) <= not b;
    layer1_outputs(7992) <= not (a or b);
    layer1_outputs(7993) <= a and b;
    layer1_outputs(7994) <= not b;
    layer1_outputs(7995) <= '0';
    layer1_outputs(7996) <= not (a or b);
    layer1_outputs(7997) <= a or b;
    layer1_outputs(7998) <= not b;
    layer1_outputs(7999) <= a;
    layer1_outputs(8000) <= '0';
    layer1_outputs(8001) <= not (a and b);
    layer1_outputs(8002) <= '0';
    layer1_outputs(8003) <= not a;
    layer1_outputs(8004) <= not b or a;
    layer1_outputs(8005) <= a;
    layer1_outputs(8006) <= '1';
    layer1_outputs(8007) <= a;
    layer1_outputs(8008) <= a and b;
    layer1_outputs(8009) <= not (a and b);
    layer1_outputs(8010) <= not a or b;
    layer1_outputs(8011) <= a;
    layer1_outputs(8012) <= not b;
    layer1_outputs(8013) <= not (a or b);
    layer1_outputs(8014) <= not (a and b);
    layer1_outputs(8015) <= '0';
    layer1_outputs(8016) <= not b;
    layer1_outputs(8017) <= '1';
    layer1_outputs(8018) <= '1';
    layer1_outputs(8019) <= not b;
    layer1_outputs(8020) <= not (a and b);
    layer1_outputs(8021) <= b and not a;
    layer1_outputs(8022) <= a and b;
    layer1_outputs(8023) <= a xor b;
    layer1_outputs(8024) <= not a;
    layer1_outputs(8025) <= not (a and b);
    layer1_outputs(8026) <= b and not a;
    layer1_outputs(8027) <= '1';
    layer1_outputs(8028) <= not b or a;
    layer1_outputs(8029) <= a;
    layer1_outputs(8030) <= not (a xor b);
    layer1_outputs(8031) <= a and b;
    layer1_outputs(8032) <= not b or a;
    layer1_outputs(8033) <= a or b;
    layer1_outputs(8034) <= not a or b;
    layer1_outputs(8035) <= not (a xor b);
    layer1_outputs(8036) <= b and not a;
    layer1_outputs(8037) <= not b or a;
    layer1_outputs(8038) <= not a or b;
    layer1_outputs(8039) <= not a or b;
    layer1_outputs(8040) <= a and not b;
    layer1_outputs(8041) <= a or b;
    layer1_outputs(8042) <= not (a xor b);
    layer1_outputs(8043) <= a xor b;
    layer1_outputs(8044) <= '1';
    layer1_outputs(8045) <= not (a or b);
    layer1_outputs(8046) <= a and b;
    layer1_outputs(8047) <= not a;
    layer1_outputs(8048) <= a and not b;
    layer1_outputs(8049) <= b;
    layer1_outputs(8050) <= '0';
    layer1_outputs(8051) <= '1';
    layer1_outputs(8052) <= a;
    layer1_outputs(8053) <= a and b;
    layer1_outputs(8054) <= b and not a;
    layer1_outputs(8055) <= not (a or b);
    layer1_outputs(8056) <= b and not a;
    layer1_outputs(8057) <= not b or a;
    layer1_outputs(8058) <= '1';
    layer1_outputs(8059) <= not a or b;
    layer1_outputs(8060) <= not b or a;
    layer1_outputs(8061) <= not b;
    layer1_outputs(8062) <= not b;
    layer1_outputs(8063) <= a and b;
    layer1_outputs(8064) <= not (a or b);
    layer1_outputs(8065) <= a and not b;
    layer1_outputs(8066) <= not (a and b);
    layer1_outputs(8067) <= not a or b;
    layer1_outputs(8068) <= not a or b;
    layer1_outputs(8069) <= not b;
    layer1_outputs(8070) <= a and not b;
    layer1_outputs(8071) <= '0';
    layer1_outputs(8072) <= a xor b;
    layer1_outputs(8073) <= a and not b;
    layer1_outputs(8074) <= not a or b;
    layer1_outputs(8075) <= a;
    layer1_outputs(8076) <= '1';
    layer1_outputs(8077) <= b and not a;
    layer1_outputs(8078) <= not b or a;
    layer1_outputs(8079) <= '0';
    layer1_outputs(8080) <= '0';
    layer1_outputs(8081) <= a or b;
    layer1_outputs(8082) <= not (a and b);
    layer1_outputs(8083) <= not (a or b);
    layer1_outputs(8084) <= not a or b;
    layer1_outputs(8085) <= not b or a;
    layer1_outputs(8086) <= a or b;
    layer1_outputs(8087) <= '1';
    layer1_outputs(8088) <= a and not b;
    layer1_outputs(8089) <= not (a xor b);
    layer1_outputs(8090) <= not (a and b);
    layer1_outputs(8091) <= b;
    layer1_outputs(8092) <= not a or b;
    layer1_outputs(8093) <= a or b;
    layer1_outputs(8094) <= not (a or b);
    layer1_outputs(8095) <= not (a and b);
    layer1_outputs(8096) <= a and not b;
    layer1_outputs(8097) <= a xor b;
    layer1_outputs(8098) <= not b;
    layer1_outputs(8099) <= a and b;
    layer1_outputs(8100) <= not (a or b);
    layer1_outputs(8101) <= a;
    layer1_outputs(8102) <= '1';
    layer1_outputs(8103) <= not b or a;
    layer1_outputs(8104) <= b and not a;
    layer1_outputs(8105) <= not (a or b);
    layer1_outputs(8106) <= not b;
    layer1_outputs(8107) <= not a;
    layer1_outputs(8108) <= b;
    layer1_outputs(8109) <= not b or a;
    layer1_outputs(8110) <= not b;
    layer1_outputs(8111) <= not (a and b);
    layer1_outputs(8112) <= a and b;
    layer1_outputs(8113) <= not b;
    layer1_outputs(8114) <= '0';
    layer1_outputs(8115) <= a and not b;
    layer1_outputs(8116) <= a xor b;
    layer1_outputs(8117) <= not a;
    layer1_outputs(8118) <= not (a and b);
    layer1_outputs(8119) <= '0';
    layer1_outputs(8120) <= a and b;
    layer1_outputs(8121) <= not b;
    layer1_outputs(8122) <= a xor b;
    layer1_outputs(8123) <= '1';
    layer1_outputs(8124) <= b;
    layer1_outputs(8125) <= a and b;
    layer1_outputs(8126) <= not a;
    layer1_outputs(8127) <= not a;
    layer1_outputs(8128) <= b;
    layer1_outputs(8129) <= b and not a;
    layer1_outputs(8130) <= a or b;
    layer1_outputs(8131) <= a and b;
    layer1_outputs(8132) <= not a or b;
    layer1_outputs(8133) <= a or b;
    layer1_outputs(8134) <= not a;
    layer1_outputs(8135) <= not b or a;
    layer1_outputs(8136) <= not a;
    layer1_outputs(8137) <= not (a xor b);
    layer1_outputs(8138) <= b;
    layer1_outputs(8139) <= a or b;
    layer1_outputs(8140) <= not a or b;
    layer1_outputs(8141) <= b;
    layer1_outputs(8142) <= a and b;
    layer1_outputs(8143) <= not b;
    layer1_outputs(8144) <= not a;
    layer1_outputs(8145) <= not b or a;
    layer1_outputs(8146) <= b;
    layer1_outputs(8147) <= '0';
    layer1_outputs(8148) <= not a or b;
    layer1_outputs(8149) <= a;
    layer1_outputs(8150) <= not a;
    layer1_outputs(8151) <= not (a and b);
    layer1_outputs(8152) <= '0';
    layer1_outputs(8153) <= '1';
    layer1_outputs(8154) <= not (a and b);
    layer1_outputs(8155) <= b and not a;
    layer1_outputs(8156) <= not (a and b);
    layer1_outputs(8157) <= b;
    layer1_outputs(8158) <= b and not a;
    layer1_outputs(8159) <= a and not b;
    layer1_outputs(8160) <= b;
    layer1_outputs(8161) <= not (a and b);
    layer1_outputs(8162) <= a and not b;
    layer1_outputs(8163) <= a and not b;
    layer1_outputs(8164) <= not (a or b);
    layer1_outputs(8165) <= a;
    layer1_outputs(8166) <= not a or b;
    layer1_outputs(8167) <= a and b;
    layer1_outputs(8168) <= a;
    layer1_outputs(8169) <= not b;
    layer1_outputs(8170) <= a and not b;
    layer1_outputs(8171) <= b and not a;
    layer1_outputs(8172) <= a or b;
    layer1_outputs(8173) <= '0';
    layer1_outputs(8174) <= '0';
    layer1_outputs(8175) <= not a or b;
    layer1_outputs(8176) <= a;
    layer1_outputs(8177) <= not b or a;
    layer1_outputs(8178) <= not (a and b);
    layer1_outputs(8179) <= '1';
    layer1_outputs(8180) <= b and not a;
    layer1_outputs(8181) <= a or b;
    layer1_outputs(8182) <= b;
    layer1_outputs(8183) <= b and not a;
    layer1_outputs(8184) <= '0';
    layer1_outputs(8185) <= not b or a;
    layer1_outputs(8186) <= not (a or b);
    layer1_outputs(8187) <= not (a and b);
    layer1_outputs(8188) <= a;
    layer1_outputs(8189) <= b and not a;
    layer1_outputs(8190) <= '0';
    layer1_outputs(8191) <= not a or b;
    layer1_outputs(8192) <= b and not a;
    layer1_outputs(8193) <= not b or a;
    layer1_outputs(8194) <= a and b;
    layer1_outputs(8195) <= b and not a;
    layer1_outputs(8196) <= a and b;
    layer1_outputs(8197) <= not (a or b);
    layer1_outputs(8198) <= b;
    layer1_outputs(8199) <= not (a xor b);
    layer1_outputs(8200) <= not b;
    layer1_outputs(8201) <= not (a or b);
    layer1_outputs(8202) <= a and b;
    layer1_outputs(8203) <= b and not a;
    layer1_outputs(8204) <= not (a and b);
    layer1_outputs(8205) <= a;
    layer1_outputs(8206) <= a;
    layer1_outputs(8207) <= not a or b;
    layer1_outputs(8208) <= not (a and b);
    layer1_outputs(8209) <= not b;
    layer1_outputs(8210) <= not (a and b);
    layer1_outputs(8211) <= a xor b;
    layer1_outputs(8212) <= a and not b;
    layer1_outputs(8213) <= a xor b;
    layer1_outputs(8214) <= not (a and b);
    layer1_outputs(8215) <= a;
    layer1_outputs(8216) <= b;
    layer1_outputs(8217) <= not a;
    layer1_outputs(8218) <= b;
    layer1_outputs(8219) <= a xor b;
    layer1_outputs(8220) <= not (a and b);
    layer1_outputs(8221) <= a or b;
    layer1_outputs(8222) <= not (a or b);
    layer1_outputs(8223) <= a;
    layer1_outputs(8224) <= not (a and b);
    layer1_outputs(8225) <= a and not b;
    layer1_outputs(8226) <= not b;
    layer1_outputs(8227) <= not (a and b);
    layer1_outputs(8228) <= not b;
    layer1_outputs(8229) <= not b or a;
    layer1_outputs(8230) <= not a;
    layer1_outputs(8231) <= not b or a;
    layer1_outputs(8232) <= a;
    layer1_outputs(8233) <= a and not b;
    layer1_outputs(8234) <= a xor b;
    layer1_outputs(8235) <= '1';
    layer1_outputs(8236) <= not b;
    layer1_outputs(8237) <= not (a or b);
    layer1_outputs(8238) <= not (a and b);
    layer1_outputs(8239) <= not (a or b);
    layer1_outputs(8240) <= not a or b;
    layer1_outputs(8241) <= a and b;
    layer1_outputs(8242) <= a;
    layer1_outputs(8243) <= not (a or b);
    layer1_outputs(8244) <= '0';
    layer1_outputs(8245) <= '1';
    layer1_outputs(8246) <= not b;
    layer1_outputs(8247) <= a;
    layer1_outputs(8248) <= '1';
    layer1_outputs(8249) <= not b or a;
    layer1_outputs(8250) <= a or b;
    layer1_outputs(8251) <= not a or b;
    layer1_outputs(8252) <= a and b;
    layer1_outputs(8253) <= not (a and b);
    layer1_outputs(8254) <= not a or b;
    layer1_outputs(8255) <= not (a xor b);
    layer1_outputs(8256) <= '1';
    layer1_outputs(8257) <= not (a and b);
    layer1_outputs(8258) <= a and b;
    layer1_outputs(8259) <= '1';
    layer1_outputs(8260) <= b and not a;
    layer1_outputs(8261) <= '0';
    layer1_outputs(8262) <= not a or b;
    layer1_outputs(8263) <= a or b;
    layer1_outputs(8264) <= not b;
    layer1_outputs(8265) <= not b or a;
    layer1_outputs(8266) <= not a;
    layer1_outputs(8267) <= a and not b;
    layer1_outputs(8268) <= not a or b;
    layer1_outputs(8269) <= '0';
    layer1_outputs(8270) <= '0';
    layer1_outputs(8271) <= a or b;
    layer1_outputs(8272) <= '1';
    layer1_outputs(8273) <= b;
    layer1_outputs(8274) <= not a or b;
    layer1_outputs(8275) <= not a;
    layer1_outputs(8276) <= not b;
    layer1_outputs(8277) <= b and not a;
    layer1_outputs(8278) <= a;
    layer1_outputs(8279) <= b;
    layer1_outputs(8280) <= not (a and b);
    layer1_outputs(8281) <= b and not a;
    layer1_outputs(8282) <= a;
    layer1_outputs(8283) <= not b;
    layer1_outputs(8284) <= a and b;
    layer1_outputs(8285) <= not a or b;
    layer1_outputs(8286) <= a;
    layer1_outputs(8287) <= b and not a;
    layer1_outputs(8288) <= '1';
    layer1_outputs(8289) <= a or b;
    layer1_outputs(8290) <= a;
    layer1_outputs(8291) <= not (a or b);
    layer1_outputs(8292) <= not a or b;
    layer1_outputs(8293) <= not (a and b);
    layer1_outputs(8294) <= not b;
    layer1_outputs(8295) <= a and not b;
    layer1_outputs(8296) <= b;
    layer1_outputs(8297) <= a or b;
    layer1_outputs(8298) <= a;
    layer1_outputs(8299) <= b and not a;
    layer1_outputs(8300) <= not (a or b);
    layer1_outputs(8301) <= not a;
    layer1_outputs(8302) <= not a;
    layer1_outputs(8303) <= '1';
    layer1_outputs(8304) <= not (a and b);
    layer1_outputs(8305) <= not a or b;
    layer1_outputs(8306) <= not (a xor b);
    layer1_outputs(8307) <= '0';
    layer1_outputs(8308) <= b and not a;
    layer1_outputs(8309) <= a and not b;
    layer1_outputs(8310) <= not (a or b);
    layer1_outputs(8311) <= not b;
    layer1_outputs(8312) <= a or b;
    layer1_outputs(8313) <= not a;
    layer1_outputs(8314) <= a xor b;
    layer1_outputs(8315) <= not a or b;
    layer1_outputs(8316) <= not a;
    layer1_outputs(8317) <= b and not a;
    layer1_outputs(8318) <= not a;
    layer1_outputs(8319) <= not (a and b);
    layer1_outputs(8320) <= not (a or b);
    layer1_outputs(8321) <= b;
    layer1_outputs(8322) <= not a;
    layer1_outputs(8323) <= not a;
    layer1_outputs(8324) <= not b or a;
    layer1_outputs(8325) <= b and not a;
    layer1_outputs(8326) <= a and not b;
    layer1_outputs(8327) <= b;
    layer1_outputs(8328) <= a and b;
    layer1_outputs(8329) <= a or b;
    layer1_outputs(8330) <= a;
    layer1_outputs(8331) <= b;
    layer1_outputs(8332) <= not (a and b);
    layer1_outputs(8333) <= b and not a;
    layer1_outputs(8334) <= a or b;
    layer1_outputs(8335) <= not (a and b);
    layer1_outputs(8336) <= not (a and b);
    layer1_outputs(8337) <= a;
    layer1_outputs(8338) <= a;
    layer1_outputs(8339) <= a or b;
    layer1_outputs(8340) <= a or b;
    layer1_outputs(8341) <= not (a and b);
    layer1_outputs(8342) <= a;
    layer1_outputs(8343) <= not b or a;
    layer1_outputs(8344) <= not (a and b);
    layer1_outputs(8345) <= a or b;
    layer1_outputs(8346) <= not b;
    layer1_outputs(8347) <= a;
    layer1_outputs(8348) <= a and b;
    layer1_outputs(8349) <= a;
    layer1_outputs(8350) <= a;
    layer1_outputs(8351) <= not a;
    layer1_outputs(8352) <= not b;
    layer1_outputs(8353) <= '1';
    layer1_outputs(8354) <= not (a and b);
    layer1_outputs(8355) <= not (a or b);
    layer1_outputs(8356) <= a and b;
    layer1_outputs(8357) <= b;
    layer1_outputs(8358) <= a or b;
    layer1_outputs(8359) <= '1';
    layer1_outputs(8360) <= a and b;
    layer1_outputs(8361) <= '0';
    layer1_outputs(8362) <= not (a or b);
    layer1_outputs(8363) <= b;
    layer1_outputs(8364) <= not a or b;
    layer1_outputs(8365) <= b;
    layer1_outputs(8366) <= b;
    layer1_outputs(8367) <= b;
    layer1_outputs(8368) <= not (a xor b);
    layer1_outputs(8369) <= a;
    layer1_outputs(8370) <= b and not a;
    layer1_outputs(8371) <= not b or a;
    layer1_outputs(8372) <= not a or b;
    layer1_outputs(8373) <= not (a or b);
    layer1_outputs(8374) <= not a;
    layer1_outputs(8375) <= not b or a;
    layer1_outputs(8376) <= not a;
    layer1_outputs(8377) <= not b or a;
    layer1_outputs(8378) <= a and not b;
    layer1_outputs(8379) <= not (a or b);
    layer1_outputs(8380) <= not b;
    layer1_outputs(8381) <= a xor b;
    layer1_outputs(8382) <= not (a and b);
    layer1_outputs(8383) <= b and not a;
    layer1_outputs(8384) <= a xor b;
    layer1_outputs(8385) <= b;
    layer1_outputs(8386) <= not (a or b);
    layer1_outputs(8387) <= not (a and b);
    layer1_outputs(8388) <= '0';
    layer1_outputs(8389) <= a and not b;
    layer1_outputs(8390) <= a and not b;
    layer1_outputs(8391) <= not b;
    layer1_outputs(8392) <= a;
    layer1_outputs(8393) <= not (a or b);
    layer1_outputs(8394) <= not (a or b);
    layer1_outputs(8395) <= not b;
    layer1_outputs(8396) <= '1';
    layer1_outputs(8397) <= a and not b;
    layer1_outputs(8398) <= not (a and b);
    layer1_outputs(8399) <= not b or a;
    layer1_outputs(8400) <= not a;
    layer1_outputs(8401) <= '1';
    layer1_outputs(8402) <= b and not a;
    layer1_outputs(8403) <= not (a xor b);
    layer1_outputs(8404) <= a xor b;
    layer1_outputs(8405) <= a and b;
    layer1_outputs(8406) <= '1';
    layer1_outputs(8407) <= a xor b;
    layer1_outputs(8408) <= a or b;
    layer1_outputs(8409) <= not (a or b);
    layer1_outputs(8410) <= a xor b;
    layer1_outputs(8411) <= a;
    layer1_outputs(8412) <= '0';
    layer1_outputs(8413) <= b and not a;
    layer1_outputs(8414) <= not a or b;
    layer1_outputs(8415) <= not a;
    layer1_outputs(8416) <= not a;
    layer1_outputs(8417) <= a and not b;
    layer1_outputs(8418) <= b and not a;
    layer1_outputs(8419) <= not b or a;
    layer1_outputs(8420) <= not a or b;
    layer1_outputs(8421) <= a and not b;
    layer1_outputs(8422) <= a and b;
    layer1_outputs(8423) <= not (a and b);
    layer1_outputs(8424) <= a or b;
    layer1_outputs(8425) <= not b or a;
    layer1_outputs(8426) <= a;
    layer1_outputs(8427) <= a;
    layer1_outputs(8428) <= a and not b;
    layer1_outputs(8429) <= not (a or b);
    layer1_outputs(8430) <= a;
    layer1_outputs(8431) <= a;
    layer1_outputs(8432) <= a and not b;
    layer1_outputs(8433) <= a;
    layer1_outputs(8434) <= a and b;
    layer1_outputs(8435) <= b and not a;
    layer1_outputs(8436) <= not (a or b);
    layer1_outputs(8437) <= a;
    layer1_outputs(8438) <= '1';
    layer1_outputs(8439) <= not b or a;
    layer1_outputs(8440) <= '1';
    layer1_outputs(8441) <= '0';
    layer1_outputs(8442) <= b and not a;
    layer1_outputs(8443) <= a and not b;
    layer1_outputs(8444) <= not (a and b);
    layer1_outputs(8445) <= a or b;
    layer1_outputs(8446) <= not (a or b);
    layer1_outputs(8447) <= not b or a;
    layer1_outputs(8448) <= not b or a;
    layer1_outputs(8449) <= '0';
    layer1_outputs(8450) <= a xor b;
    layer1_outputs(8451) <= '1';
    layer1_outputs(8452) <= a;
    layer1_outputs(8453) <= a and b;
    layer1_outputs(8454) <= not b;
    layer1_outputs(8455) <= b;
    layer1_outputs(8456) <= b;
    layer1_outputs(8457) <= '0';
    layer1_outputs(8458) <= '0';
    layer1_outputs(8459) <= not a;
    layer1_outputs(8460) <= not (a or b);
    layer1_outputs(8461) <= not (a and b);
    layer1_outputs(8462) <= '0';
    layer1_outputs(8463) <= a or b;
    layer1_outputs(8464) <= not (a or b);
    layer1_outputs(8465) <= b;
    layer1_outputs(8466) <= b and not a;
    layer1_outputs(8467) <= not (a or b);
    layer1_outputs(8468) <= '0';
    layer1_outputs(8469) <= b;
    layer1_outputs(8470) <= a or b;
    layer1_outputs(8471) <= a and not b;
    layer1_outputs(8472) <= '0';
    layer1_outputs(8473) <= a and not b;
    layer1_outputs(8474) <= not a;
    layer1_outputs(8475) <= a xor b;
    layer1_outputs(8476) <= not b;
    layer1_outputs(8477) <= b;
    layer1_outputs(8478) <= not a;
    layer1_outputs(8479) <= not (a or b);
    layer1_outputs(8480) <= a or b;
    layer1_outputs(8481) <= not (a or b);
    layer1_outputs(8482) <= not (a xor b);
    layer1_outputs(8483) <= not (a or b);
    layer1_outputs(8484) <= not (a xor b);
    layer1_outputs(8485) <= a;
    layer1_outputs(8486) <= not b or a;
    layer1_outputs(8487) <= not b;
    layer1_outputs(8488) <= b;
    layer1_outputs(8489) <= a and not b;
    layer1_outputs(8490) <= not b or a;
    layer1_outputs(8491) <= not (a xor b);
    layer1_outputs(8492) <= not b or a;
    layer1_outputs(8493) <= not b or a;
    layer1_outputs(8494) <= a or b;
    layer1_outputs(8495) <= not (a and b);
    layer1_outputs(8496) <= '1';
    layer1_outputs(8497) <= '1';
    layer1_outputs(8498) <= b and not a;
    layer1_outputs(8499) <= not a or b;
    layer1_outputs(8500) <= a;
    layer1_outputs(8501) <= b;
    layer1_outputs(8502) <= not (a xor b);
    layer1_outputs(8503) <= not a;
    layer1_outputs(8504) <= a and not b;
    layer1_outputs(8505) <= not b;
    layer1_outputs(8506) <= b;
    layer1_outputs(8507) <= '0';
    layer1_outputs(8508) <= not a or b;
    layer1_outputs(8509) <= not (a and b);
    layer1_outputs(8510) <= a;
    layer1_outputs(8511) <= '0';
    layer1_outputs(8512) <= b and not a;
    layer1_outputs(8513) <= a and not b;
    layer1_outputs(8514) <= not a or b;
    layer1_outputs(8515) <= '0';
    layer1_outputs(8516) <= not a;
    layer1_outputs(8517) <= not b;
    layer1_outputs(8518) <= a or b;
    layer1_outputs(8519) <= not b or a;
    layer1_outputs(8520) <= a xor b;
    layer1_outputs(8521) <= a and not b;
    layer1_outputs(8522) <= not (a or b);
    layer1_outputs(8523) <= not a;
    layer1_outputs(8524) <= not b or a;
    layer1_outputs(8525) <= a xor b;
    layer1_outputs(8526) <= not b;
    layer1_outputs(8527) <= not a;
    layer1_outputs(8528) <= not b;
    layer1_outputs(8529) <= not a or b;
    layer1_outputs(8530) <= '1';
    layer1_outputs(8531) <= not a or b;
    layer1_outputs(8532) <= a;
    layer1_outputs(8533) <= b and not a;
    layer1_outputs(8534) <= a;
    layer1_outputs(8535) <= a and not b;
    layer1_outputs(8536) <= not b or a;
    layer1_outputs(8537) <= not (a or b);
    layer1_outputs(8538) <= not (a and b);
    layer1_outputs(8539) <= not b or a;
    layer1_outputs(8540) <= '0';
    layer1_outputs(8541) <= b;
    layer1_outputs(8542) <= a xor b;
    layer1_outputs(8543) <= not a;
    layer1_outputs(8544) <= b;
    layer1_outputs(8545) <= b;
    layer1_outputs(8546) <= b;
    layer1_outputs(8547) <= '1';
    layer1_outputs(8548) <= not a;
    layer1_outputs(8549) <= not b or a;
    layer1_outputs(8550) <= '0';
    layer1_outputs(8551) <= not a;
    layer1_outputs(8552) <= '0';
    layer1_outputs(8553) <= b;
    layer1_outputs(8554) <= not (a and b);
    layer1_outputs(8555) <= not (a and b);
    layer1_outputs(8556) <= a;
    layer1_outputs(8557) <= '0';
    layer1_outputs(8558) <= not (a or b);
    layer1_outputs(8559) <= not b or a;
    layer1_outputs(8560) <= '0';
    layer1_outputs(8561) <= a or b;
    layer1_outputs(8562) <= a xor b;
    layer1_outputs(8563) <= b and not a;
    layer1_outputs(8564) <= '0';
    layer1_outputs(8565) <= a or b;
    layer1_outputs(8566) <= '0';
    layer1_outputs(8567) <= '1';
    layer1_outputs(8568) <= not (a or b);
    layer1_outputs(8569) <= not b;
    layer1_outputs(8570) <= a or b;
    layer1_outputs(8571) <= not (a and b);
    layer1_outputs(8572) <= b;
    layer1_outputs(8573) <= a;
    layer1_outputs(8574) <= a and not b;
    layer1_outputs(8575) <= '1';
    layer1_outputs(8576) <= b;
    layer1_outputs(8577) <= not b or a;
    layer1_outputs(8578) <= a xor b;
    layer1_outputs(8579) <= a and not b;
    layer1_outputs(8580) <= '0';
    layer1_outputs(8581) <= a;
    layer1_outputs(8582) <= not (a or b);
    layer1_outputs(8583) <= '0';
    layer1_outputs(8584) <= not a or b;
    layer1_outputs(8585) <= a;
    layer1_outputs(8586) <= b;
    layer1_outputs(8587) <= not a;
    layer1_outputs(8588) <= not (a or b);
    layer1_outputs(8589) <= not a;
    layer1_outputs(8590) <= a xor b;
    layer1_outputs(8591) <= a or b;
    layer1_outputs(8592) <= '1';
    layer1_outputs(8593) <= '0';
    layer1_outputs(8594) <= not a or b;
    layer1_outputs(8595) <= b and not a;
    layer1_outputs(8596) <= not a or b;
    layer1_outputs(8597) <= not (a xor b);
    layer1_outputs(8598) <= '0';
    layer1_outputs(8599) <= not b;
    layer1_outputs(8600) <= '1';
    layer1_outputs(8601) <= a and b;
    layer1_outputs(8602) <= a and not b;
    layer1_outputs(8603) <= not a or b;
    layer1_outputs(8604) <= b and not a;
    layer1_outputs(8605) <= a and b;
    layer1_outputs(8606) <= not (a or b);
    layer1_outputs(8607) <= not (a xor b);
    layer1_outputs(8608) <= a and b;
    layer1_outputs(8609) <= not (a or b);
    layer1_outputs(8610) <= not b;
    layer1_outputs(8611) <= not a;
    layer1_outputs(8612) <= a;
    layer1_outputs(8613) <= b and not a;
    layer1_outputs(8614) <= not (a and b);
    layer1_outputs(8615) <= not b or a;
    layer1_outputs(8616) <= not (a or b);
    layer1_outputs(8617) <= not (a or b);
    layer1_outputs(8618) <= a or b;
    layer1_outputs(8619) <= a and not b;
    layer1_outputs(8620) <= a and not b;
    layer1_outputs(8621) <= a and not b;
    layer1_outputs(8622) <= not a;
    layer1_outputs(8623) <= not (a or b);
    layer1_outputs(8624) <= a or b;
    layer1_outputs(8625) <= a and not b;
    layer1_outputs(8626) <= not (a or b);
    layer1_outputs(8627) <= a and not b;
    layer1_outputs(8628) <= not a or b;
    layer1_outputs(8629) <= a xor b;
    layer1_outputs(8630) <= b;
    layer1_outputs(8631) <= b;
    layer1_outputs(8632) <= a and b;
    layer1_outputs(8633) <= not b;
    layer1_outputs(8634) <= '0';
    layer1_outputs(8635) <= a;
    layer1_outputs(8636) <= b and not a;
    layer1_outputs(8637) <= not b;
    layer1_outputs(8638) <= not (a xor b);
    layer1_outputs(8639) <= not (a or b);
    layer1_outputs(8640) <= not b;
    layer1_outputs(8641) <= a and not b;
    layer1_outputs(8642) <= '1';
    layer1_outputs(8643) <= a or b;
    layer1_outputs(8644) <= a;
    layer1_outputs(8645) <= a xor b;
    layer1_outputs(8646) <= b and not a;
    layer1_outputs(8647) <= not (a xor b);
    layer1_outputs(8648) <= a;
    layer1_outputs(8649) <= '1';
    layer1_outputs(8650) <= a and not b;
    layer1_outputs(8651) <= a or b;
    layer1_outputs(8652) <= '0';
    layer1_outputs(8653) <= a;
    layer1_outputs(8654) <= not a or b;
    layer1_outputs(8655) <= a;
    layer1_outputs(8656) <= not a;
    layer1_outputs(8657) <= not a;
    layer1_outputs(8658) <= a or b;
    layer1_outputs(8659) <= not b;
    layer1_outputs(8660) <= not (a xor b);
    layer1_outputs(8661) <= not (a or b);
    layer1_outputs(8662) <= not (a and b);
    layer1_outputs(8663) <= not (a xor b);
    layer1_outputs(8664) <= '0';
    layer1_outputs(8665) <= not a;
    layer1_outputs(8666) <= a and b;
    layer1_outputs(8667) <= '0';
    layer1_outputs(8668) <= a;
    layer1_outputs(8669) <= not (a or b);
    layer1_outputs(8670) <= a or b;
    layer1_outputs(8671) <= a;
    layer1_outputs(8672) <= b and not a;
    layer1_outputs(8673) <= a and b;
    layer1_outputs(8674) <= a or b;
    layer1_outputs(8675) <= a xor b;
    layer1_outputs(8676) <= b and not a;
    layer1_outputs(8677) <= not a or b;
    layer1_outputs(8678) <= b and not a;
    layer1_outputs(8679) <= not b or a;
    layer1_outputs(8680) <= not a or b;
    layer1_outputs(8681) <= not b or a;
    layer1_outputs(8682) <= not (a or b);
    layer1_outputs(8683) <= not (a xor b);
    layer1_outputs(8684) <= not (a and b);
    layer1_outputs(8685) <= a;
    layer1_outputs(8686) <= not b or a;
    layer1_outputs(8687) <= not b or a;
    layer1_outputs(8688) <= '0';
    layer1_outputs(8689) <= a;
    layer1_outputs(8690) <= b and not a;
    layer1_outputs(8691) <= not (a or b);
    layer1_outputs(8692) <= b;
    layer1_outputs(8693) <= not (a and b);
    layer1_outputs(8694) <= a or b;
    layer1_outputs(8695) <= a or b;
    layer1_outputs(8696) <= not b;
    layer1_outputs(8697) <= a xor b;
    layer1_outputs(8698) <= '0';
    layer1_outputs(8699) <= not (a or b);
    layer1_outputs(8700) <= not a or b;
    layer1_outputs(8701) <= not (a xor b);
    layer1_outputs(8702) <= b and not a;
    layer1_outputs(8703) <= '1';
    layer1_outputs(8704) <= a;
    layer1_outputs(8705) <= b and not a;
    layer1_outputs(8706) <= a and b;
    layer1_outputs(8707) <= b and not a;
    layer1_outputs(8708) <= not b;
    layer1_outputs(8709) <= '0';
    layer1_outputs(8710) <= not (a xor b);
    layer1_outputs(8711) <= not (a and b);
    layer1_outputs(8712) <= not b or a;
    layer1_outputs(8713) <= not b;
    layer1_outputs(8714) <= a and not b;
    layer1_outputs(8715) <= a and b;
    layer1_outputs(8716) <= not (a and b);
    layer1_outputs(8717) <= b;
    layer1_outputs(8718) <= a xor b;
    layer1_outputs(8719) <= not b or a;
    layer1_outputs(8720) <= not a or b;
    layer1_outputs(8721) <= a and b;
    layer1_outputs(8722) <= not b or a;
    layer1_outputs(8723) <= b and not a;
    layer1_outputs(8724) <= a xor b;
    layer1_outputs(8725) <= b and not a;
    layer1_outputs(8726) <= a;
    layer1_outputs(8727) <= not a or b;
    layer1_outputs(8728) <= a;
    layer1_outputs(8729) <= not b or a;
    layer1_outputs(8730) <= a;
    layer1_outputs(8731) <= not a or b;
    layer1_outputs(8732) <= not a;
    layer1_outputs(8733) <= not (a and b);
    layer1_outputs(8734) <= a and not b;
    layer1_outputs(8735) <= not b;
    layer1_outputs(8736) <= not a;
    layer1_outputs(8737) <= not a;
    layer1_outputs(8738) <= a xor b;
    layer1_outputs(8739) <= not a or b;
    layer1_outputs(8740) <= not a or b;
    layer1_outputs(8741) <= a;
    layer1_outputs(8742) <= b;
    layer1_outputs(8743) <= not (a xor b);
    layer1_outputs(8744) <= a and b;
    layer1_outputs(8745) <= a;
    layer1_outputs(8746) <= not a;
    layer1_outputs(8747) <= not a or b;
    layer1_outputs(8748) <= not (a xor b);
    layer1_outputs(8749) <= b;
    layer1_outputs(8750) <= not b;
    layer1_outputs(8751) <= not (a xor b);
    layer1_outputs(8752) <= not (a or b);
    layer1_outputs(8753) <= not a;
    layer1_outputs(8754) <= not b or a;
    layer1_outputs(8755) <= a xor b;
    layer1_outputs(8756) <= not a or b;
    layer1_outputs(8757) <= a and b;
    layer1_outputs(8758) <= a;
    layer1_outputs(8759) <= not b or a;
    layer1_outputs(8760) <= '0';
    layer1_outputs(8761) <= not (a and b);
    layer1_outputs(8762) <= not b or a;
    layer1_outputs(8763) <= a or b;
    layer1_outputs(8764) <= not (a xor b);
    layer1_outputs(8765) <= b;
    layer1_outputs(8766) <= not (a and b);
    layer1_outputs(8767) <= not b or a;
    layer1_outputs(8768) <= not b;
    layer1_outputs(8769) <= not (a or b);
    layer1_outputs(8770) <= b and not a;
    layer1_outputs(8771) <= not b;
    layer1_outputs(8772) <= not (a and b);
    layer1_outputs(8773) <= a and b;
    layer1_outputs(8774) <= a and not b;
    layer1_outputs(8775) <= not b or a;
    layer1_outputs(8776) <= a and b;
    layer1_outputs(8777) <= a and b;
    layer1_outputs(8778) <= '0';
    layer1_outputs(8779) <= not b;
    layer1_outputs(8780) <= '1';
    layer1_outputs(8781) <= a or b;
    layer1_outputs(8782) <= b;
    layer1_outputs(8783) <= a and not b;
    layer1_outputs(8784) <= a and not b;
    layer1_outputs(8785) <= not a or b;
    layer1_outputs(8786) <= a;
    layer1_outputs(8787) <= not a;
    layer1_outputs(8788) <= a;
    layer1_outputs(8789) <= b;
    layer1_outputs(8790) <= not b;
    layer1_outputs(8791) <= a or b;
    layer1_outputs(8792) <= a and not b;
    layer1_outputs(8793) <= not a or b;
    layer1_outputs(8794) <= a and b;
    layer1_outputs(8795) <= '1';
    layer1_outputs(8796) <= not a or b;
    layer1_outputs(8797) <= not a or b;
    layer1_outputs(8798) <= not a;
    layer1_outputs(8799) <= a;
    layer1_outputs(8800) <= not b or a;
    layer1_outputs(8801) <= not (a or b);
    layer1_outputs(8802) <= a and b;
    layer1_outputs(8803) <= not a;
    layer1_outputs(8804) <= not (a xor b);
    layer1_outputs(8805) <= not a or b;
    layer1_outputs(8806) <= a or b;
    layer1_outputs(8807) <= a or b;
    layer1_outputs(8808) <= b;
    layer1_outputs(8809) <= not a;
    layer1_outputs(8810) <= not (a xor b);
    layer1_outputs(8811) <= a xor b;
    layer1_outputs(8812) <= a and not b;
    layer1_outputs(8813) <= not a;
    layer1_outputs(8814) <= not (a and b);
    layer1_outputs(8815) <= not (a or b);
    layer1_outputs(8816) <= not a or b;
    layer1_outputs(8817) <= a or b;
    layer1_outputs(8818) <= not a;
    layer1_outputs(8819) <= a xor b;
    layer1_outputs(8820) <= b;
    layer1_outputs(8821) <= not a or b;
    layer1_outputs(8822) <= a or b;
    layer1_outputs(8823) <= not a;
    layer1_outputs(8824) <= a;
    layer1_outputs(8825) <= not b or a;
    layer1_outputs(8826) <= b;
    layer1_outputs(8827) <= a and not b;
    layer1_outputs(8828) <= not (a and b);
    layer1_outputs(8829) <= b;
    layer1_outputs(8830) <= a;
    layer1_outputs(8831) <= not a or b;
    layer1_outputs(8832) <= a and not b;
    layer1_outputs(8833) <= not b;
    layer1_outputs(8834) <= not a or b;
    layer1_outputs(8835) <= b;
    layer1_outputs(8836) <= a xor b;
    layer1_outputs(8837) <= '0';
    layer1_outputs(8838) <= not (a or b);
    layer1_outputs(8839) <= a and b;
    layer1_outputs(8840) <= b and not a;
    layer1_outputs(8841) <= a;
    layer1_outputs(8842) <= a or b;
    layer1_outputs(8843) <= not a;
    layer1_outputs(8844) <= not a;
    layer1_outputs(8845) <= a and not b;
    layer1_outputs(8846) <= a and not b;
    layer1_outputs(8847) <= a and not b;
    layer1_outputs(8848) <= a or b;
    layer1_outputs(8849) <= '1';
    layer1_outputs(8850) <= not a;
    layer1_outputs(8851) <= not (a xor b);
    layer1_outputs(8852) <= not b or a;
    layer1_outputs(8853) <= not (a and b);
    layer1_outputs(8854) <= b and not a;
    layer1_outputs(8855) <= not b or a;
    layer1_outputs(8856) <= '1';
    layer1_outputs(8857) <= a or b;
    layer1_outputs(8858) <= not a;
    layer1_outputs(8859) <= not b;
    layer1_outputs(8860) <= '1';
    layer1_outputs(8861) <= b and not a;
    layer1_outputs(8862) <= not a;
    layer1_outputs(8863) <= '0';
    layer1_outputs(8864) <= a and not b;
    layer1_outputs(8865) <= a and not b;
    layer1_outputs(8866) <= not (a or b);
    layer1_outputs(8867) <= not b or a;
    layer1_outputs(8868) <= a and not b;
    layer1_outputs(8869) <= not a;
    layer1_outputs(8870) <= b;
    layer1_outputs(8871) <= not a;
    layer1_outputs(8872) <= not (a and b);
    layer1_outputs(8873) <= b and not a;
    layer1_outputs(8874) <= a;
    layer1_outputs(8875) <= a or b;
    layer1_outputs(8876) <= not (a and b);
    layer1_outputs(8877) <= not a;
    layer1_outputs(8878) <= not a;
    layer1_outputs(8879) <= a or b;
    layer1_outputs(8880) <= a and not b;
    layer1_outputs(8881) <= not (a or b);
    layer1_outputs(8882) <= a and b;
    layer1_outputs(8883) <= not b;
    layer1_outputs(8884) <= b;
    layer1_outputs(8885) <= not a;
    layer1_outputs(8886) <= not (a or b);
    layer1_outputs(8887) <= a or b;
    layer1_outputs(8888) <= a and b;
    layer1_outputs(8889) <= a;
    layer1_outputs(8890) <= not b;
    layer1_outputs(8891) <= not (a and b);
    layer1_outputs(8892) <= b;
    layer1_outputs(8893) <= b;
    layer1_outputs(8894) <= not b;
    layer1_outputs(8895) <= not b;
    layer1_outputs(8896) <= a and not b;
    layer1_outputs(8897) <= not (a and b);
    layer1_outputs(8898) <= not (a or b);
    layer1_outputs(8899) <= not (a or b);
    layer1_outputs(8900) <= not a or b;
    layer1_outputs(8901) <= not a or b;
    layer1_outputs(8902) <= '1';
    layer1_outputs(8903) <= b and not a;
    layer1_outputs(8904) <= a;
    layer1_outputs(8905) <= a or b;
    layer1_outputs(8906) <= not b;
    layer1_outputs(8907) <= a;
    layer1_outputs(8908) <= a and not b;
    layer1_outputs(8909) <= not (a and b);
    layer1_outputs(8910) <= b and not a;
    layer1_outputs(8911) <= b and not a;
    layer1_outputs(8912) <= a or b;
    layer1_outputs(8913) <= b;
    layer1_outputs(8914) <= not a or b;
    layer1_outputs(8915) <= not (a or b);
    layer1_outputs(8916) <= a;
    layer1_outputs(8917) <= not (a and b);
    layer1_outputs(8918) <= a and b;
    layer1_outputs(8919) <= not a or b;
    layer1_outputs(8920) <= not (a or b);
    layer1_outputs(8921) <= a and b;
    layer1_outputs(8922) <= b and not a;
    layer1_outputs(8923) <= not (a and b);
    layer1_outputs(8924) <= not (a or b);
    layer1_outputs(8925) <= a and b;
    layer1_outputs(8926) <= not a;
    layer1_outputs(8927) <= not b;
    layer1_outputs(8928) <= b;
    layer1_outputs(8929) <= b and not a;
    layer1_outputs(8930) <= b;
    layer1_outputs(8931) <= not (a and b);
    layer1_outputs(8932) <= a and b;
    layer1_outputs(8933) <= not b or a;
    layer1_outputs(8934) <= a;
    layer1_outputs(8935) <= a and not b;
    layer1_outputs(8936) <= not (a or b);
    layer1_outputs(8937) <= not (a and b);
    layer1_outputs(8938) <= '1';
    layer1_outputs(8939) <= not b;
    layer1_outputs(8940) <= b and not a;
    layer1_outputs(8941) <= not (a or b);
    layer1_outputs(8942) <= a;
    layer1_outputs(8943) <= not (a and b);
    layer1_outputs(8944) <= '1';
    layer1_outputs(8945) <= not b;
    layer1_outputs(8946) <= a;
    layer1_outputs(8947) <= a and b;
    layer1_outputs(8948) <= not b;
    layer1_outputs(8949) <= '1';
    layer1_outputs(8950) <= a and b;
    layer1_outputs(8951) <= not (a or b);
    layer1_outputs(8952) <= b;
    layer1_outputs(8953) <= not (a and b);
    layer1_outputs(8954) <= not b;
    layer1_outputs(8955) <= not (a or b);
    layer1_outputs(8956) <= a and b;
    layer1_outputs(8957) <= not a;
    layer1_outputs(8958) <= '1';
    layer1_outputs(8959) <= a and not b;
    layer1_outputs(8960) <= '1';
    layer1_outputs(8961) <= a and not b;
    layer1_outputs(8962) <= b and not a;
    layer1_outputs(8963) <= b;
    layer1_outputs(8964) <= b and not a;
    layer1_outputs(8965) <= '1';
    layer1_outputs(8966) <= not (a xor b);
    layer1_outputs(8967) <= a xor b;
    layer1_outputs(8968) <= not a;
    layer1_outputs(8969) <= not a;
    layer1_outputs(8970) <= not a or b;
    layer1_outputs(8971) <= b;
    layer1_outputs(8972) <= a xor b;
    layer1_outputs(8973) <= not (a xor b);
    layer1_outputs(8974) <= not a or b;
    layer1_outputs(8975) <= not (a and b);
    layer1_outputs(8976) <= b and not a;
    layer1_outputs(8977) <= not a or b;
    layer1_outputs(8978) <= '0';
    layer1_outputs(8979) <= a xor b;
    layer1_outputs(8980) <= '1';
    layer1_outputs(8981) <= b;
    layer1_outputs(8982) <= not b or a;
    layer1_outputs(8983) <= not a or b;
    layer1_outputs(8984) <= '0';
    layer1_outputs(8985) <= a or b;
    layer1_outputs(8986) <= a;
    layer1_outputs(8987) <= not a;
    layer1_outputs(8988) <= '1';
    layer1_outputs(8989) <= a xor b;
    layer1_outputs(8990) <= b;
    layer1_outputs(8991) <= b;
    layer1_outputs(8992) <= a and not b;
    layer1_outputs(8993) <= a and b;
    layer1_outputs(8994) <= not b or a;
    layer1_outputs(8995) <= not b;
    layer1_outputs(8996) <= b;
    layer1_outputs(8997) <= not a or b;
    layer1_outputs(8998) <= not a;
    layer1_outputs(8999) <= b;
    layer1_outputs(9000) <= '1';
    layer1_outputs(9001) <= not (a and b);
    layer1_outputs(9002) <= a xor b;
    layer1_outputs(9003) <= a xor b;
    layer1_outputs(9004) <= not a or b;
    layer1_outputs(9005) <= not a or b;
    layer1_outputs(9006) <= not b or a;
    layer1_outputs(9007) <= not a;
    layer1_outputs(9008) <= not (a or b);
    layer1_outputs(9009) <= not a;
    layer1_outputs(9010) <= not (a xor b);
    layer1_outputs(9011) <= b;
    layer1_outputs(9012) <= '1';
    layer1_outputs(9013) <= a or b;
    layer1_outputs(9014) <= a and not b;
    layer1_outputs(9015) <= '0';
    layer1_outputs(9016) <= '0';
    layer1_outputs(9017) <= not a;
    layer1_outputs(9018) <= a and b;
    layer1_outputs(9019) <= b and not a;
    layer1_outputs(9020) <= a or b;
    layer1_outputs(9021) <= '1';
    layer1_outputs(9022) <= a;
    layer1_outputs(9023) <= not b;
    layer1_outputs(9024) <= not a;
    layer1_outputs(9025) <= not (a xor b);
    layer1_outputs(9026) <= b;
    layer1_outputs(9027) <= b;
    layer1_outputs(9028) <= '0';
    layer1_outputs(9029) <= not (a xor b);
    layer1_outputs(9030) <= '0';
    layer1_outputs(9031) <= a and b;
    layer1_outputs(9032) <= a;
    layer1_outputs(9033) <= a and b;
    layer1_outputs(9034) <= not (a or b);
    layer1_outputs(9035) <= a;
    layer1_outputs(9036) <= not (a and b);
    layer1_outputs(9037) <= not (a or b);
    layer1_outputs(9038) <= '0';
    layer1_outputs(9039) <= not a;
    layer1_outputs(9040) <= not a or b;
    layer1_outputs(9041) <= not (a xor b);
    layer1_outputs(9042) <= not a;
    layer1_outputs(9043) <= not a or b;
    layer1_outputs(9044) <= not (a xor b);
    layer1_outputs(9045) <= not b;
    layer1_outputs(9046) <= a and not b;
    layer1_outputs(9047) <= a;
    layer1_outputs(9048) <= a and not b;
    layer1_outputs(9049) <= not (a and b);
    layer1_outputs(9050) <= a;
    layer1_outputs(9051) <= not b;
    layer1_outputs(9052) <= a;
    layer1_outputs(9053) <= not (a and b);
    layer1_outputs(9054) <= a and b;
    layer1_outputs(9055) <= not (a xor b);
    layer1_outputs(9056) <= '1';
    layer1_outputs(9057) <= not b or a;
    layer1_outputs(9058) <= '0';
    layer1_outputs(9059) <= '1';
    layer1_outputs(9060) <= b;
    layer1_outputs(9061) <= not a or b;
    layer1_outputs(9062) <= '0';
    layer1_outputs(9063) <= not (a or b);
    layer1_outputs(9064) <= a and not b;
    layer1_outputs(9065) <= not a;
    layer1_outputs(9066) <= a and b;
    layer1_outputs(9067) <= a or b;
    layer1_outputs(9068) <= not (a or b);
    layer1_outputs(9069) <= '0';
    layer1_outputs(9070) <= not a or b;
    layer1_outputs(9071) <= not b;
    layer1_outputs(9072) <= b;
    layer1_outputs(9073) <= not (a and b);
    layer1_outputs(9074) <= '1';
    layer1_outputs(9075) <= not a;
    layer1_outputs(9076) <= a or b;
    layer1_outputs(9077) <= b and not a;
    layer1_outputs(9078) <= a;
    layer1_outputs(9079) <= a and b;
    layer1_outputs(9080) <= not a;
    layer1_outputs(9081) <= not b or a;
    layer1_outputs(9082) <= b;
    layer1_outputs(9083) <= a or b;
    layer1_outputs(9084) <= b;
    layer1_outputs(9085) <= a and b;
    layer1_outputs(9086) <= not (a or b);
    layer1_outputs(9087) <= not a or b;
    layer1_outputs(9088) <= not a;
    layer1_outputs(9089) <= not b;
    layer1_outputs(9090) <= a or b;
    layer1_outputs(9091) <= not a or b;
    layer1_outputs(9092) <= a or b;
    layer1_outputs(9093) <= b;
    layer1_outputs(9094) <= a;
    layer1_outputs(9095) <= not b or a;
    layer1_outputs(9096) <= b and not a;
    layer1_outputs(9097) <= a and b;
    layer1_outputs(9098) <= not b or a;
    layer1_outputs(9099) <= not a or b;
    layer1_outputs(9100) <= a and b;
    layer1_outputs(9101) <= a or b;
    layer1_outputs(9102) <= b and not a;
    layer1_outputs(9103) <= not a;
    layer1_outputs(9104) <= not (a or b);
    layer1_outputs(9105) <= a xor b;
    layer1_outputs(9106) <= a or b;
    layer1_outputs(9107) <= not a;
    layer1_outputs(9108) <= a or b;
    layer1_outputs(9109) <= a xor b;
    layer1_outputs(9110) <= '1';
    layer1_outputs(9111) <= '0';
    layer1_outputs(9112) <= a;
    layer1_outputs(9113) <= not a or b;
    layer1_outputs(9114) <= not a or b;
    layer1_outputs(9115) <= not (a xor b);
    layer1_outputs(9116) <= not a or b;
    layer1_outputs(9117) <= not (a xor b);
    layer1_outputs(9118) <= not (a and b);
    layer1_outputs(9119) <= not (a or b);
    layer1_outputs(9120) <= b and not a;
    layer1_outputs(9121) <= b;
    layer1_outputs(9122) <= a xor b;
    layer1_outputs(9123) <= not b or a;
    layer1_outputs(9124) <= not a or b;
    layer1_outputs(9125) <= a or b;
    layer1_outputs(9126) <= not (a or b);
    layer1_outputs(9127) <= b and not a;
    layer1_outputs(9128) <= b;
    layer1_outputs(9129) <= a or b;
    layer1_outputs(9130) <= not a;
    layer1_outputs(9131) <= not a or b;
    layer1_outputs(9132) <= b;
    layer1_outputs(9133) <= not a or b;
    layer1_outputs(9134) <= a and not b;
    layer1_outputs(9135) <= not (a and b);
    layer1_outputs(9136) <= b;
    layer1_outputs(9137) <= a;
    layer1_outputs(9138) <= not a;
    layer1_outputs(9139) <= a;
    layer1_outputs(9140) <= '0';
    layer1_outputs(9141) <= a and b;
    layer1_outputs(9142) <= not (a and b);
    layer1_outputs(9143) <= a or b;
    layer1_outputs(9144) <= not a;
    layer1_outputs(9145) <= a;
    layer1_outputs(9146) <= a xor b;
    layer1_outputs(9147) <= a;
    layer1_outputs(9148) <= not a or b;
    layer1_outputs(9149) <= a and b;
    layer1_outputs(9150) <= not (a xor b);
    layer1_outputs(9151) <= a or b;
    layer1_outputs(9152) <= '0';
    layer1_outputs(9153) <= not b or a;
    layer1_outputs(9154) <= '0';
    layer1_outputs(9155) <= not (a or b);
    layer1_outputs(9156) <= b;
    layer1_outputs(9157) <= not a or b;
    layer1_outputs(9158) <= not b or a;
    layer1_outputs(9159) <= not (a and b);
    layer1_outputs(9160) <= a and b;
    layer1_outputs(9161) <= b;
    layer1_outputs(9162) <= a;
    layer1_outputs(9163) <= not b;
    layer1_outputs(9164) <= not b;
    layer1_outputs(9165) <= '1';
    layer1_outputs(9166) <= '0';
    layer1_outputs(9167) <= not (a and b);
    layer1_outputs(9168) <= not (a or b);
    layer1_outputs(9169) <= b and not a;
    layer1_outputs(9170) <= b and not a;
    layer1_outputs(9171) <= '0';
    layer1_outputs(9172) <= '1';
    layer1_outputs(9173) <= b and not a;
    layer1_outputs(9174) <= a or b;
    layer1_outputs(9175) <= a xor b;
    layer1_outputs(9176) <= b and not a;
    layer1_outputs(9177) <= '1';
    layer1_outputs(9178) <= a or b;
    layer1_outputs(9179) <= not (a or b);
    layer1_outputs(9180) <= a and not b;
    layer1_outputs(9181) <= '1';
    layer1_outputs(9182) <= '0';
    layer1_outputs(9183) <= not a or b;
    layer1_outputs(9184) <= not b;
    layer1_outputs(9185) <= not (a and b);
    layer1_outputs(9186) <= a and b;
    layer1_outputs(9187) <= not b;
    layer1_outputs(9188) <= b and not a;
    layer1_outputs(9189) <= not b;
    layer1_outputs(9190) <= not b or a;
    layer1_outputs(9191) <= '1';
    layer1_outputs(9192) <= a or b;
    layer1_outputs(9193) <= b;
    layer1_outputs(9194) <= a;
    layer1_outputs(9195) <= not b;
    layer1_outputs(9196) <= b and not a;
    layer1_outputs(9197) <= not b;
    layer1_outputs(9198) <= '0';
    layer1_outputs(9199) <= a;
    layer1_outputs(9200) <= not (a or b);
    layer1_outputs(9201) <= a and not b;
    layer1_outputs(9202) <= not (a xor b);
    layer1_outputs(9203) <= b;
    layer1_outputs(9204) <= a xor b;
    layer1_outputs(9205) <= a xor b;
    layer1_outputs(9206) <= not a or b;
    layer1_outputs(9207) <= a;
    layer1_outputs(9208) <= b and not a;
    layer1_outputs(9209) <= b and not a;
    layer1_outputs(9210) <= not (a or b);
    layer1_outputs(9211) <= not b;
    layer1_outputs(9212) <= b and not a;
    layer1_outputs(9213) <= a;
    layer1_outputs(9214) <= a or b;
    layer1_outputs(9215) <= a xor b;
    layer1_outputs(9216) <= not a or b;
    layer1_outputs(9217) <= not a;
    layer1_outputs(9218) <= b;
    layer1_outputs(9219) <= b;
    layer1_outputs(9220) <= not b or a;
    layer1_outputs(9221) <= not a;
    layer1_outputs(9222) <= b;
    layer1_outputs(9223) <= not (a and b);
    layer1_outputs(9224) <= '0';
    layer1_outputs(9225) <= not a;
    layer1_outputs(9226) <= not b or a;
    layer1_outputs(9227) <= not a;
    layer1_outputs(9228) <= a;
    layer1_outputs(9229) <= not (a and b);
    layer1_outputs(9230) <= not a;
    layer1_outputs(9231) <= a or b;
    layer1_outputs(9232) <= not a;
    layer1_outputs(9233) <= not a;
    layer1_outputs(9234) <= a and b;
    layer1_outputs(9235) <= not b or a;
    layer1_outputs(9236) <= a or b;
    layer1_outputs(9237) <= not b;
    layer1_outputs(9238) <= not a or b;
    layer1_outputs(9239) <= '1';
    layer1_outputs(9240) <= not (a or b);
    layer1_outputs(9241) <= a xor b;
    layer1_outputs(9242) <= a xor b;
    layer1_outputs(9243) <= a;
    layer1_outputs(9244) <= not a;
    layer1_outputs(9245) <= not a;
    layer1_outputs(9246) <= a and b;
    layer1_outputs(9247) <= not b or a;
    layer1_outputs(9248) <= not b or a;
    layer1_outputs(9249) <= not a or b;
    layer1_outputs(9250) <= b and not a;
    layer1_outputs(9251) <= a or b;
    layer1_outputs(9252) <= not (a and b);
    layer1_outputs(9253) <= a xor b;
    layer1_outputs(9254) <= a and b;
    layer1_outputs(9255) <= b;
    layer1_outputs(9256) <= not b;
    layer1_outputs(9257) <= not (a or b);
    layer1_outputs(9258) <= not a or b;
    layer1_outputs(9259) <= not a or b;
    layer1_outputs(9260) <= a;
    layer1_outputs(9261) <= not (a xor b);
    layer1_outputs(9262) <= '1';
    layer1_outputs(9263) <= not (a xor b);
    layer1_outputs(9264) <= not (a or b);
    layer1_outputs(9265) <= a xor b;
    layer1_outputs(9266) <= not b;
    layer1_outputs(9267) <= '1';
    layer1_outputs(9268) <= not a;
    layer1_outputs(9269) <= b and not a;
    layer1_outputs(9270) <= not b;
    layer1_outputs(9271) <= '0';
    layer1_outputs(9272) <= not b or a;
    layer1_outputs(9273) <= not b;
    layer1_outputs(9274) <= not b or a;
    layer1_outputs(9275) <= not (a and b);
    layer1_outputs(9276) <= a or b;
    layer1_outputs(9277) <= not (a xor b);
    layer1_outputs(9278) <= a or b;
    layer1_outputs(9279) <= not a or b;
    layer1_outputs(9280) <= not (a or b);
    layer1_outputs(9281) <= a;
    layer1_outputs(9282) <= not (a and b);
    layer1_outputs(9283) <= not (a and b);
    layer1_outputs(9284) <= not (a xor b);
    layer1_outputs(9285) <= not (a or b);
    layer1_outputs(9286) <= a and not b;
    layer1_outputs(9287) <= not b;
    layer1_outputs(9288) <= b;
    layer1_outputs(9289) <= a;
    layer1_outputs(9290) <= not (a and b);
    layer1_outputs(9291) <= '1';
    layer1_outputs(9292) <= '1';
    layer1_outputs(9293) <= not b;
    layer1_outputs(9294) <= not a or b;
    layer1_outputs(9295) <= not a;
    layer1_outputs(9296) <= not b or a;
    layer1_outputs(9297) <= a and not b;
    layer1_outputs(9298) <= a xor b;
    layer1_outputs(9299) <= '1';
    layer1_outputs(9300) <= not (a and b);
    layer1_outputs(9301) <= a or b;
    layer1_outputs(9302) <= a or b;
    layer1_outputs(9303) <= a and not b;
    layer1_outputs(9304) <= not a;
    layer1_outputs(9305) <= a xor b;
    layer1_outputs(9306) <= not b or a;
    layer1_outputs(9307) <= a;
    layer1_outputs(9308) <= a or b;
    layer1_outputs(9309) <= '0';
    layer1_outputs(9310) <= b;
    layer1_outputs(9311) <= not b or a;
    layer1_outputs(9312) <= a;
    layer1_outputs(9313) <= not (a or b);
    layer1_outputs(9314) <= not b or a;
    layer1_outputs(9315) <= not b;
    layer1_outputs(9316) <= a;
    layer1_outputs(9317) <= not b;
    layer1_outputs(9318) <= not a;
    layer1_outputs(9319) <= a and b;
    layer1_outputs(9320) <= not a;
    layer1_outputs(9321) <= not a;
    layer1_outputs(9322) <= a and b;
    layer1_outputs(9323) <= a and b;
    layer1_outputs(9324) <= b and not a;
    layer1_outputs(9325) <= '1';
    layer1_outputs(9326) <= a;
    layer1_outputs(9327) <= not b or a;
    layer1_outputs(9328) <= '0';
    layer1_outputs(9329) <= not b;
    layer1_outputs(9330) <= not (a and b);
    layer1_outputs(9331) <= b;
    layer1_outputs(9332) <= not a;
    layer1_outputs(9333) <= b and not a;
    layer1_outputs(9334) <= a and b;
    layer1_outputs(9335) <= '0';
    layer1_outputs(9336) <= not (a xor b);
    layer1_outputs(9337) <= a or b;
    layer1_outputs(9338) <= a and b;
    layer1_outputs(9339) <= a and b;
    layer1_outputs(9340) <= b and not a;
    layer1_outputs(9341) <= not (a or b);
    layer1_outputs(9342) <= not b;
    layer1_outputs(9343) <= not a or b;
    layer1_outputs(9344) <= not (a and b);
    layer1_outputs(9345) <= a or b;
    layer1_outputs(9346) <= not b;
    layer1_outputs(9347) <= a;
    layer1_outputs(9348) <= not a;
    layer1_outputs(9349) <= not b;
    layer1_outputs(9350) <= not (a or b);
    layer1_outputs(9351) <= not b;
    layer1_outputs(9352) <= a and not b;
    layer1_outputs(9353) <= a;
    layer1_outputs(9354) <= a xor b;
    layer1_outputs(9355) <= not (a or b);
    layer1_outputs(9356) <= not b;
    layer1_outputs(9357) <= not (a and b);
    layer1_outputs(9358) <= '0';
    layer1_outputs(9359) <= not a;
    layer1_outputs(9360) <= a and not b;
    layer1_outputs(9361) <= not a or b;
    layer1_outputs(9362) <= not b;
    layer1_outputs(9363) <= not (a and b);
    layer1_outputs(9364) <= not b or a;
    layer1_outputs(9365) <= '1';
    layer1_outputs(9366) <= a and b;
    layer1_outputs(9367) <= not a;
    layer1_outputs(9368) <= not a or b;
    layer1_outputs(9369) <= not (a and b);
    layer1_outputs(9370) <= '0';
    layer1_outputs(9371) <= a;
    layer1_outputs(9372) <= a and not b;
    layer1_outputs(9373) <= not a;
    layer1_outputs(9374) <= a;
    layer1_outputs(9375) <= not b or a;
    layer1_outputs(9376) <= not b or a;
    layer1_outputs(9377) <= a and b;
    layer1_outputs(9378) <= not (a or b);
    layer1_outputs(9379) <= a;
    layer1_outputs(9380) <= a xor b;
    layer1_outputs(9381) <= a;
    layer1_outputs(9382) <= a or b;
    layer1_outputs(9383) <= a and not b;
    layer1_outputs(9384) <= not b;
    layer1_outputs(9385) <= '0';
    layer1_outputs(9386) <= not (a or b);
    layer1_outputs(9387) <= b and not a;
    layer1_outputs(9388) <= a and b;
    layer1_outputs(9389) <= b;
    layer1_outputs(9390) <= a or b;
    layer1_outputs(9391) <= not (a xor b);
    layer1_outputs(9392) <= b and not a;
    layer1_outputs(9393) <= not a or b;
    layer1_outputs(9394) <= a or b;
    layer1_outputs(9395) <= a or b;
    layer1_outputs(9396) <= a or b;
    layer1_outputs(9397) <= a and b;
    layer1_outputs(9398) <= '0';
    layer1_outputs(9399) <= a or b;
    layer1_outputs(9400) <= a;
    layer1_outputs(9401) <= not b or a;
    layer1_outputs(9402) <= not a or b;
    layer1_outputs(9403) <= not b;
    layer1_outputs(9404) <= b and not a;
    layer1_outputs(9405) <= a and not b;
    layer1_outputs(9406) <= b and not a;
    layer1_outputs(9407) <= not a or b;
    layer1_outputs(9408) <= '1';
    layer1_outputs(9409) <= not b;
    layer1_outputs(9410) <= a or b;
    layer1_outputs(9411) <= '1';
    layer1_outputs(9412) <= not b or a;
    layer1_outputs(9413) <= '0';
    layer1_outputs(9414) <= not (a and b);
    layer1_outputs(9415) <= not b or a;
    layer1_outputs(9416) <= '1';
    layer1_outputs(9417) <= b;
    layer1_outputs(9418) <= a or b;
    layer1_outputs(9419) <= a or b;
    layer1_outputs(9420) <= not b or a;
    layer1_outputs(9421) <= a and not b;
    layer1_outputs(9422) <= not a;
    layer1_outputs(9423) <= not (a or b);
    layer1_outputs(9424) <= a xor b;
    layer1_outputs(9425) <= not (a and b);
    layer1_outputs(9426) <= not (a or b);
    layer1_outputs(9427) <= not (a or b);
    layer1_outputs(9428) <= a;
    layer1_outputs(9429) <= '0';
    layer1_outputs(9430) <= a or b;
    layer1_outputs(9431) <= not a or b;
    layer1_outputs(9432) <= not a or b;
    layer1_outputs(9433) <= not a or b;
    layer1_outputs(9434) <= '0';
    layer1_outputs(9435) <= not (a or b);
    layer1_outputs(9436) <= not a or b;
    layer1_outputs(9437) <= b;
    layer1_outputs(9438) <= not (a or b);
    layer1_outputs(9439) <= not a;
    layer1_outputs(9440) <= not (a and b);
    layer1_outputs(9441) <= not (a xor b);
    layer1_outputs(9442) <= a and not b;
    layer1_outputs(9443) <= b and not a;
    layer1_outputs(9444) <= not b or a;
    layer1_outputs(9445) <= b and not a;
    layer1_outputs(9446) <= not (a and b);
    layer1_outputs(9447) <= a xor b;
    layer1_outputs(9448) <= a and not b;
    layer1_outputs(9449) <= not b;
    layer1_outputs(9450) <= '0';
    layer1_outputs(9451) <= b and not a;
    layer1_outputs(9452) <= a and b;
    layer1_outputs(9453) <= '1';
    layer1_outputs(9454) <= not a;
    layer1_outputs(9455) <= not (a or b);
    layer1_outputs(9456) <= a and not b;
    layer1_outputs(9457) <= not a or b;
    layer1_outputs(9458) <= not (a xor b);
    layer1_outputs(9459) <= not a;
    layer1_outputs(9460) <= not (a and b);
    layer1_outputs(9461) <= not b;
    layer1_outputs(9462) <= '0';
    layer1_outputs(9463) <= not (a and b);
    layer1_outputs(9464) <= b;
    layer1_outputs(9465) <= a and b;
    layer1_outputs(9466) <= b;
    layer1_outputs(9467) <= a and b;
    layer1_outputs(9468) <= not (a or b);
    layer1_outputs(9469) <= not a or b;
    layer1_outputs(9470) <= '1';
    layer1_outputs(9471) <= not b;
    layer1_outputs(9472) <= not a or b;
    layer1_outputs(9473) <= a and b;
    layer1_outputs(9474) <= a and b;
    layer1_outputs(9475) <= not (a and b);
    layer1_outputs(9476) <= not b;
    layer1_outputs(9477) <= '1';
    layer1_outputs(9478) <= a or b;
    layer1_outputs(9479) <= not a;
    layer1_outputs(9480) <= b and not a;
    layer1_outputs(9481) <= a and not b;
    layer1_outputs(9482) <= not (a xor b);
    layer1_outputs(9483) <= b;
    layer1_outputs(9484) <= not b;
    layer1_outputs(9485) <= b and not a;
    layer1_outputs(9486) <= '0';
    layer1_outputs(9487) <= '0';
    layer1_outputs(9488) <= a or b;
    layer1_outputs(9489) <= not b;
    layer1_outputs(9490) <= a or b;
    layer1_outputs(9491) <= not b;
    layer1_outputs(9492) <= '1';
    layer1_outputs(9493) <= '0';
    layer1_outputs(9494) <= not b;
    layer1_outputs(9495) <= not (a and b);
    layer1_outputs(9496) <= a and b;
    layer1_outputs(9497) <= not (a and b);
    layer1_outputs(9498) <= '1';
    layer1_outputs(9499) <= a or b;
    layer1_outputs(9500) <= a and not b;
    layer1_outputs(9501) <= b and not a;
    layer1_outputs(9502) <= not b;
    layer1_outputs(9503) <= not (a and b);
    layer1_outputs(9504) <= b and not a;
    layer1_outputs(9505) <= a;
    layer1_outputs(9506) <= not (a and b);
    layer1_outputs(9507) <= not b;
    layer1_outputs(9508) <= a;
    layer1_outputs(9509) <= a and b;
    layer1_outputs(9510) <= not (a and b);
    layer1_outputs(9511) <= a and b;
    layer1_outputs(9512) <= b;
    layer1_outputs(9513) <= not b or a;
    layer1_outputs(9514) <= not a or b;
    layer1_outputs(9515) <= a;
    layer1_outputs(9516) <= a and not b;
    layer1_outputs(9517) <= '0';
    layer1_outputs(9518) <= a and not b;
    layer1_outputs(9519) <= a xor b;
    layer1_outputs(9520) <= a and not b;
    layer1_outputs(9521) <= a;
    layer1_outputs(9522) <= '1';
    layer1_outputs(9523) <= '0';
    layer1_outputs(9524) <= a and b;
    layer1_outputs(9525) <= '0';
    layer1_outputs(9526) <= a xor b;
    layer1_outputs(9527) <= b and not a;
    layer1_outputs(9528) <= not a or b;
    layer1_outputs(9529) <= a;
    layer1_outputs(9530) <= not (a and b);
    layer1_outputs(9531) <= not b;
    layer1_outputs(9532) <= not a or b;
    layer1_outputs(9533) <= a xor b;
    layer1_outputs(9534) <= a and b;
    layer1_outputs(9535) <= not a or b;
    layer1_outputs(9536) <= not a or b;
    layer1_outputs(9537) <= a xor b;
    layer1_outputs(9538) <= a or b;
    layer1_outputs(9539) <= not (a xor b);
    layer1_outputs(9540) <= '0';
    layer1_outputs(9541) <= not (a or b);
    layer1_outputs(9542) <= '0';
    layer1_outputs(9543) <= '1';
    layer1_outputs(9544) <= a;
    layer1_outputs(9545) <= not (a or b);
    layer1_outputs(9546) <= b;
    layer1_outputs(9547) <= not (a or b);
    layer1_outputs(9548) <= not a;
    layer1_outputs(9549) <= a and not b;
    layer1_outputs(9550) <= '1';
    layer1_outputs(9551) <= a;
    layer1_outputs(9552) <= not (a and b);
    layer1_outputs(9553) <= a and b;
    layer1_outputs(9554) <= not (a xor b);
    layer1_outputs(9555) <= not a;
    layer1_outputs(9556) <= b and not a;
    layer1_outputs(9557) <= a and b;
    layer1_outputs(9558) <= a xor b;
    layer1_outputs(9559) <= a or b;
    layer1_outputs(9560) <= not a or b;
    layer1_outputs(9561) <= not a;
    layer1_outputs(9562) <= not b;
    layer1_outputs(9563) <= not a or b;
    layer1_outputs(9564) <= not a or b;
    layer1_outputs(9565) <= not b or a;
    layer1_outputs(9566) <= not b;
    layer1_outputs(9567) <= a;
    layer1_outputs(9568) <= not b;
    layer1_outputs(9569) <= not b;
    layer1_outputs(9570) <= not (a xor b);
    layer1_outputs(9571) <= a or b;
    layer1_outputs(9572) <= '1';
    layer1_outputs(9573) <= not b;
    layer1_outputs(9574) <= a and not b;
    layer1_outputs(9575) <= not (a or b);
    layer1_outputs(9576) <= '0';
    layer1_outputs(9577) <= '0';
    layer1_outputs(9578) <= a or b;
    layer1_outputs(9579) <= '0';
    layer1_outputs(9580) <= a and not b;
    layer1_outputs(9581) <= not b;
    layer1_outputs(9582) <= not b or a;
    layer1_outputs(9583) <= a or b;
    layer1_outputs(9584) <= '1';
    layer1_outputs(9585) <= not b;
    layer1_outputs(9586) <= b;
    layer1_outputs(9587) <= not (a and b);
    layer1_outputs(9588) <= not (a and b);
    layer1_outputs(9589) <= b;
    layer1_outputs(9590) <= a or b;
    layer1_outputs(9591) <= not b;
    layer1_outputs(9592) <= a and not b;
    layer1_outputs(9593) <= a or b;
    layer1_outputs(9594) <= a and not b;
    layer1_outputs(9595) <= a;
    layer1_outputs(9596) <= a;
    layer1_outputs(9597) <= '0';
    layer1_outputs(9598) <= not (a xor b);
    layer1_outputs(9599) <= not a or b;
    layer1_outputs(9600) <= not b;
    layer1_outputs(9601) <= not (a and b);
    layer1_outputs(9602) <= a and not b;
    layer1_outputs(9603) <= not b;
    layer1_outputs(9604) <= a;
    layer1_outputs(9605) <= b and not a;
    layer1_outputs(9606) <= '1';
    layer1_outputs(9607) <= a;
    layer1_outputs(9608) <= b and not a;
    layer1_outputs(9609) <= not a;
    layer1_outputs(9610) <= a and b;
    layer1_outputs(9611) <= a;
    layer1_outputs(9612) <= '0';
    layer1_outputs(9613) <= a;
    layer1_outputs(9614) <= a or b;
    layer1_outputs(9615) <= not (a and b);
    layer1_outputs(9616) <= not b;
    layer1_outputs(9617) <= not a;
    layer1_outputs(9618) <= a and not b;
    layer1_outputs(9619) <= not a or b;
    layer1_outputs(9620) <= not a or b;
    layer1_outputs(9621) <= a or b;
    layer1_outputs(9622) <= b and not a;
    layer1_outputs(9623) <= a xor b;
    layer1_outputs(9624) <= not (a or b);
    layer1_outputs(9625) <= '1';
    layer1_outputs(9626) <= a;
    layer1_outputs(9627) <= b;
    layer1_outputs(9628) <= not (a and b);
    layer1_outputs(9629) <= b;
    layer1_outputs(9630) <= b and not a;
    layer1_outputs(9631) <= a and b;
    layer1_outputs(9632) <= a and b;
    layer1_outputs(9633) <= a;
    layer1_outputs(9634) <= b;
    layer1_outputs(9635) <= b and not a;
    layer1_outputs(9636) <= a and b;
    layer1_outputs(9637) <= not (a or b);
    layer1_outputs(9638) <= a or b;
    layer1_outputs(9639) <= a and not b;
    layer1_outputs(9640) <= not a or b;
    layer1_outputs(9641) <= '1';
    layer1_outputs(9642) <= a xor b;
    layer1_outputs(9643) <= not a;
    layer1_outputs(9644) <= a or b;
    layer1_outputs(9645) <= a xor b;
    layer1_outputs(9646) <= '1';
    layer1_outputs(9647) <= a and not b;
    layer1_outputs(9648) <= not b;
    layer1_outputs(9649) <= not b;
    layer1_outputs(9650) <= '1';
    layer1_outputs(9651) <= a or b;
    layer1_outputs(9652) <= '0';
    layer1_outputs(9653) <= a;
    layer1_outputs(9654) <= a or b;
    layer1_outputs(9655) <= not b or a;
    layer1_outputs(9656) <= not b;
    layer1_outputs(9657) <= not a or b;
    layer1_outputs(9658) <= b;
    layer1_outputs(9659) <= not (a and b);
    layer1_outputs(9660) <= not b or a;
    layer1_outputs(9661) <= not b;
    layer1_outputs(9662) <= not (a or b);
    layer1_outputs(9663) <= not b;
    layer1_outputs(9664) <= not (a or b);
    layer1_outputs(9665) <= b and not a;
    layer1_outputs(9666) <= not a;
    layer1_outputs(9667) <= a and not b;
    layer1_outputs(9668) <= not a;
    layer1_outputs(9669) <= not b or a;
    layer1_outputs(9670) <= a xor b;
    layer1_outputs(9671) <= not a;
    layer1_outputs(9672) <= a and b;
    layer1_outputs(9673) <= not (a or b);
    layer1_outputs(9674) <= b and not a;
    layer1_outputs(9675) <= not b;
    layer1_outputs(9676) <= not (a or b);
    layer1_outputs(9677) <= a;
    layer1_outputs(9678) <= b and not a;
    layer1_outputs(9679) <= '0';
    layer1_outputs(9680) <= a or b;
    layer1_outputs(9681) <= a xor b;
    layer1_outputs(9682) <= not (a and b);
    layer1_outputs(9683) <= b;
    layer1_outputs(9684) <= b and not a;
    layer1_outputs(9685) <= a and not b;
    layer1_outputs(9686) <= a or b;
    layer1_outputs(9687) <= a;
    layer1_outputs(9688) <= not (a xor b);
    layer1_outputs(9689) <= not (a and b);
    layer1_outputs(9690) <= a or b;
    layer1_outputs(9691) <= not (a or b);
    layer1_outputs(9692) <= '1';
    layer1_outputs(9693) <= b;
    layer1_outputs(9694) <= b;
    layer1_outputs(9695) <= '1';
    layer1_outputs(9696) <= a or b;
    layer1_outputs(9697) <= '0';
    layer1_outputs(9698) <= not a;
    layer1_outputs(9699) <= '1';
    layer1_outputs(9700) <= not a;
    layer1_outputs(9701) <= not (a and b);
    layer1_outputs(9702) <= not b or a;
    layer1_outputs(9703) <= not a;
    layer1_outputs(9704) <= a or b;
    layer1_outputs(9705) <= a and b;
    layer1_outputs(9706) <= not a;
    layer1_outputs(9707) <= '0';
    layer1_outputs(9708) <= not (a or b);
    layer1_outputs(9709) <= not b;
    layer1_outputs(9710) <= not a;
    layer1_outputs(9711) <= not a;
    layer1_outputs(9712) <= not (a and b);
    layer1_outputs(9713) <= not a or b;
    layer1_outputs(9714) <= not b;
    layer1_outputs(9715) <= a;
    layer1_outputs(9716) <= a;
    layer1_outputs(9717) <= a and not b;
    layer1_outputs(9718) <= b;
    layer1_outputs(9719) <= not b;
    layer1_outputs(9720) <= '1';
    layer1_outputs(9721) <= not (a and b);
    layer1_outputs(9722) <= a or b;
    layer1_outputs(9723) <= a and b;
    layer1_outputs(9724) <= a or b;
    layer1_outputs(9725) <= not a or b;
    layer1_outputs(9726) <= not (a xor b);
    layer1_outputs(9727) <= '0';
    layer1_outputs(9728) <= not a;
    layer1_outputs(9729) <= not a or b;
    layer1_outputs(9730) <= not a or b;
    layer1_outputs(9731) <= a and b;
    layer1_outputs(9732) <= a and b;
    layer1_outputs(9733) <= not b or a;
    layer1_outputs(9734) <= b and not a;
    layer1_outputs(9735) <= not a or b;
    layer1_outputs(9736) <= not b;
    layer1_outputs(9737) <= a and b;
    layer1_outputs(9738) <= '0';
    layer1_outputs(9739) <= '0';
    layer1_outputs(9740) <= a and b;
    layer1_outputs(9741) <= '0';
    layer1_outputs(9742) <= a and not b;
    layer1_outputs(9743) <= b and not a;
    layer1_outputs(9744) <= not a;
    layer1_outputs(9745) <= b and not a;
    layer1_outputs(9746) <= b;
    layer1_outputs(9747) <= not (a and b);
    layer1_outputs(9748) <= not (a or b);
    layer1_outputs(9749) <= not (a and b);
    layer1_outputs(9750) <= not b;
    layer1_outputs(9751) <= not (a and b);
    layer1_outputs(9752) <= b and not a;
    layer1_outputs(9753) <= '1';
    layer1_outputs(9754) <= not a;
    layer1_outputs(9755) <= b and not a;
    layer1_outputs(9756) <= not b or a;
    layer1_outputs(9757) <= not (a or b);
    layer1_outputs(9758) <= a;
    layer1_outputs(9759) <= not b;
    layer1_outputs(9760) <= not b or a;
    layer1_outputs(9761) <= not (a or b);
    layer1_outputs(9762) <= '0';
    layer1_outputs(9763) <= not (a and b);
    layer1_outputs(9764) <= a;
    layer1_outputs(9765) <= not (a or b);
    layer1_outputs(9766) <= not (a and b);
    layer1_outputs(9767) <= not a;
    layer1_outputs(9768) <= b;
    layer1_outputs(9769) <= b;
    layer1_outputs(9770) <= '0';
    layer1_outputs(9771) <= not b or a;
    layer1_outputs(9772) <= b;
    layer1_outputs(9773) <= not a;
    layer1_outputs(9774) <= not a;
    layer1_outputs(9775) <= not (a xor b);
    layer1_outputs(9776) <= not b;
    layer1_outputs(9777) <= not b;
    layer1_outputs(9778) <= not (a or b);
    layer1_outputs(9779) <= not a or b;
    layer1_outputs(9780) <= not (a or b);
    layer1_outputs(9781) <= '1';
    layer1_outputs(9782) <= not a or b;
    layer1_outputs(9783) <= a and b;
    layer1_outputs(9784) <= not (a or b);
    layer1_outputs(9785) <= not a;
    layer1_outputs(9786) <= a and b;
    layer1_outputs(9787) <= not a;
    layer1_outputs(9788) <= b and not a;
    layer1_outputs(9789) <= '1';
    layer1_outputs(9790) <= '0';
    layer1_outputs(9791) <= not a;
    layer1_outputs(9792) <= a and b;
    layer1_outputs(9793) <= a and b;
    layer1_outputs(9794) <= a;
    layer1_outputs(9795) <= not (a and b);
    layer1_outputs(9796) <= a or b;
    layer1_outputs(9797) <= not b or a;
    layer1_outputs(9798) <= not b or a;
    layer1_outputs(9799) <= '1';
    layer1_outputs(9800) <= not (a xor b);
    layer1_outputs(9801) <= not a;
    layer1_outputs(9802) <= b and not a;
    layer1_outputs(9803) <= a xor b;
    layer1_outputs(9804) <= not a or b;
    layer1_outputs(9805) <= a and not b;
    layer1_outputs(9806) <= not (a and b);
    layer1_outputs(9807) <= not a;
    layer1_outputs(9808) <= b and not a;
    layer1_outputs(9809) <= not a;
    layer1_outputs(9810) <= b and not a;
    layer1_outputs(9811) <= b;
    layer1_outputs(9812) <= b and not a;
    layer1_outputs(9813) <= not (a or b);
    layer1_outputs(9814) <= a or b;
    layer1_outputs(9815) <= b and not a;
    layer1_outputs(9816) <= not a;
    layer1_outputs(9817) <= b and not a;
    layer1_outputs(9818) <= not (a and b);
    layer1_outputs(9819) <= a or b;
    layer1_outputs(9820) <= '0';
    layer1_outputs(9821) <= not b;
    layer1_outputs(9822) <= not (a and b);
    layer1_outputs(9823) <= not a or b;
    layer1_outputs(9824) <= a and not b;
    layer1_outputs(9825) <= '0';
    layer1_outputs(9826) <= '1';
    layer1_outputs(9827) <= not (a and b);
    layer1_outputs(9828) <= a or b;
    layer1_outputs(9829) <= not a or b;
    layer1_outputs(9830) <= not (a xor b);
    layer1_outputs(9831) <= not a;
    layer1_outputs(9832) <= not (a and b);
    layer1_outputs(9833) <= a;
    layer1_outputs(9834) <= not b;
    layer1_outputs(9835) <= not b or a;
    layer1_outputs(9836) <= not b;
    layer1_outputs(9837) <= not (a and b);
    layer1_outputs(9838) <= a or b;
    layer1_outputs(9839) <= not (a xor b);
    layer1_outputs(9840) <= '0';
    layer1_outputs(9841) <= not a or b;
    layer1_outputs(9842) <= not (a and b);
    layer1_outputs(9843) <= not a or b;
    layer1_outputs(9844) <= b and not a;
    layer1_outputs(9845) <= '0';
    layer1_outputs(9846) <= not (a and b);
    layer1_outputs(9847) <= not (a xor b);
    layer1_outputs(9848) <= a and not b;
    layer1_outputs(9849) <= not b;
    layer1_outputs(9850) <= a and b;
    layer1_outputs(9851) <= a xor b;
    layer1_outputs(9852) <= a and not b;
    layer1_outputs(9853) <= '1';
    layer1_outputs(9854) <= a;
    layer1_outputs(9855) <= not (a or b);
    layer1_outputs(9856) <= not (a xor b);
    layer1_outputs(9857) <= a xor b;
    layer1_outputs(9858) <= not b;
    layer1_outputs(9859) <= not a or b;
    layer1_outputs(9860) <= not b;
    layer1_outputs(9861) <= a;
    layer1_outputs(9862) <= a and b;
    layer1_outputs(9863) <= not b;
    layer1_outputs(9864) <= not b or a;
    layer1_outputs(9865) <= a;
    layer1_outputs(9866) <= a and b;
    layer1_outputs(9867) <= a and b;
    layer1_outputs(9868) <= a and not b;
    layer1_outputs(9869) <= not b or a;
    layer1_outputs(9870) <= b;
    layer1_outputs(9871) <= b;
    layer1_outputs(9872) <= '1';
    layer1_outputs(9873) <= not a or b;
    layer1_outputs(9874) <= '1';
    layer1_outputs(9875) <= b;
    layer1_outputs(9876) <= a and not b;
    layer1_outputs(9877) <= not (a or b);
    layer1_outputs(9878) <= not a or b;
    layer1_outputs(9879) <= not b or a;
    layer1_outputs(9880) <= not (a xor b);
    layer1_outputs(9881) <= a;
    layer1_outputs(9882) <= not (a or b);
    layer1_outputs(9883) <= not a;
    layer1_outputs(9884) <= a and not b;
    layer1_outputs(9885) <= not (a or b);
    layer1_outputs(9886) <= not a or b;
    layer1_outputs(9887) <= a;
    layer1_outputs(9888) <= not b or a;
    layer1_outputs(9889) <= a and b;
    layer1_outputs(9890) <= not b;
    layer1_outputs(9891) <= not a;
    layer1_outputs(9892) <= not b or a;
    layer1_outputs(9893) <= a or b;
    layer1_outputs(9894) <= not b or a;
    layer1_outputs(9895) <= a and b;
    layer1_outputs(9896) <= a;
    layer1_outputs(9897) <= not (a xor b);
    layer1_outputs(9898) <= not (a and b);
    layer1_outputs(9899) <= a and b;
    layer1_outputs(9900) <= a;
    layer1_outputs(9901) <= not a or b;
    layer1_outputs(9902) <= b and not a;
    layer1_outputs(9903) <= '1';
    layer1_outputs(9904) <= '1';
    layer1_outputs(9905) <= a xor b;
    layer1_outputs(9906) <= not (a or b);
    layer1_outputs(9907) <= a;
    layer1_outputs(9908) <= a xor b;
    layer1_outputs(9909) <= not b;
    layer1_outputs(9910) <= a and not b;
    layer1_outputs(9911) <= not a;
    layer1_outputs(9912) <= not (a xor b);
    layer1_outputs(9913) <= not b;
    layer1_outputs(9914) <= not b or a;
    layer1_outputs(9915) <= b and not a;
    layer1_outputs(9916) <= not a;
    layer1_outputs(9917) <= a xor b;
    layer1_outputs(9918) <= not a or b;
    layer1_outputs(9919) <= '1';
    layer1_outputs(9920) <= not a;
    layer1_outputs(9921) <= a and not b;
    layer1_outputs(9922) <= a and b;
    layer1_outputs(9923) <= not b or a;
    layer1_outputs(9924) <= a or b;
    layer1_outputs(9925) <= a xor b;
    layer1_outputs(9926) <= '0';
    layer1_outputs(9927) <= not (a or b);
    layer1_outputs(9928) <= a xor b;
    layer1_outputs(9929) <= not a;
    layer1_outputs(9930) <= '0';
    layer1_outputs(9931) <= b and not a;
    layer1_outputs(9932) <= '0';
    layer1_outputs(9933) <= b and not a;
    layer1_outputs(9934) <= a and not b;
    layer1_outputs(9935) <= a and b;
    layer1_outputs(9936) <= b;
    layer1_outputs(9937) <= b and not a;
    layer1_outputs(9938) <= not (a xor b);
    layer1_outputs(9939) <= not b;
    layer1_outputs(9940) <= not b;
    layer1_outputs(9941) <= not (a or b);
    layer1_outputs(9942) <= '0';
    layer1_outputs(9943) <= not b;
    layer1_outputs(9944) <= '0';
    layer1_outputs(9945) <= not (a or b);
    layer1_outputs(9946) <= '0';
    layer1_outputs(9947) <= not a;
    layer1_outputs(9948) <= '0';
    layer1_outputs(9949) <= not a or b;
    layer1_outputs(9950) <= b and not a;
    layer1_outputs(9951) <= a and b;
    layer1_outputs(9952) <= a;
    layer1_outputs(9953) <= a and b;
    layer1_outputs(9954) <= not (a and b);
    layer1_outputs(9955) <= not b or a;
    layer1_outputs(9956) <= a and not b;
    layer1_outputs(9957) <= b;
    layer1_outputs(9958) <= not (a and b);
    layer1_outputs(9959) <= a or b;
    layer1_outputs(9960) <= '0';
    layer1_outputs(9961) <= not b;
    layer1_outputs(9962) <= a and b;
    layer1_outputs(9963) <= a xor b;
    layer1_outputs(9964) <= a or b;
    layer1_outputs(9965) <= not b;
    layer1_outputs(9966) <= not b;
    layer1_outputs(9967) <= b and not a;
    layer1_outputs(9968) <= b and not a;
    layer1_outputs(9969) <= a and b;
    layer1_outputs(9970) <= a;
    layer1_outputs(9971) <= not (a xor b);
    layer1_outputs(9972) <= '1';
    layer1_outputs(9973) <= a and b;
    layer1_outputs(9974) <= a or b;
    layer1_outputs(9975) <= a or b;
    layer1_outputs(9976) <= '0';
    layer1_outputs(9977) <= b;
    layer1_outputs(9978) <= b and not a;
    layer1_outputs(9979) <= not (a or b);
    layer1_outputs(9980) <= not b;
    layer1_outputs(9981) <= a or b;
    layer1_outputs(9982) <= not a;
    layer1_outputs(9983) <= '0';
    layer1_outputs(9984) <= '1';
    layer1_outputs(9985) <= '0';
    layer1_outputs(9986) <= not b;
    layer1_outputs(9987) <= a or b;
    layer1_outputs(9988) <= b and not a;
    layer1_outputs(9989) <= a or b;
    layer1_outputs(9990) <= a;
    layer1_outputs(9991) <= a or b;
    layer1_outputs(9992) <= not b or a;
    layer1_outputs(9993) <= a and b;
    layer1_outputs(9994) <= not (a or b);
    layer1_outputs(9995) <= a xor b;
    layer1_outputs(9996) <= a;
    layer1_outputs(9997) <= not a or b;
    layer1_outputs(9998) <= a and not b;
    layer1_outputs(9999) <= not a;
    layer1_outputs(10000) <= not a;
    layer1_outputs(10001) <= a;
    layer1_outputs(10002) <= a;
    layer1_outputs(10003) <= a and not b;
    layer1_outputs(10004) <= not b;
    layer1_outputs(10005) <= b;
    layer1_outputs(10006) <= a or b;
    layer1_outputs(10007) <= a;
    layer1_outputs(10008) <= '1';
    layer1_outputs(10009) <= not a;
    layer1_outputs(10010) <= '1';
    layer1_outputs(10011) <= a and not b;
    layer1_outputs(10012) <= not b or a;
    layer1_outputs(10013) <= not b or a;
    layer1_outputs(10014) <= not b;
    layer1_outputs(10015) <= a;
    layer1_outputs(10016) <= not (a and b);
    layer1_outputs(10017) <= not a or b;
    layer1_outputs(10018) <= '1';
    layer1_outputs(10019) <= a or b;
    layer1_outputs(10020) <= a;
    layer1_outputs(10021) <= a and b;
    layer1_outputs(10022) <= a or b;
    layer1_outputs(10023) <= a or b;
    layer1_outputs(10024) <= '0';
    layer1_outputs(10025) <= not b or a;
    layer1_outputs(10026) <= '0';
    layer1_outputs(10027) <= '0';
    layer1_outputs(10028) <= not b;
    layer1_outputs(10029) <= a or b;
    layer1_outputs(10030) <= a and not b;
    layer1_outputs(10031) <= not a;
    layer1_outputs(10032) <= not b or a;
    layer1_outputs(10033) <= a and not b;
    layer1_outputs(10034) <= a xor b;
    layer1_outputs(10035) <= not (a and b);
    layer1_outputs(10036) <= a or b;
    layer1_outputs(10037) <= not (a and b);
    layer1_outputs(10038) <= b;
    layer1_outputs(10039) <= a or b;
    layer1_outputs(10040) <= not a;
    layer1_outputs(10041) <= a and not b;
    layer1_outputs(10042) <= a and not b;
    layer1_outputs(10043) <= not (a or b);
    layer1_outputs(10044) <= not a;
    layer1_outputs(10045) <= '0';
    layer1_outputs(10046) <= not b;
    layer1_outputs(10047) <= a and not b;
    layer1_outputs(10048) <= b and not a;
    layer1_outputs(10049) <= not a or b;
    layer1_outputs(10050) <= a xor b;
    layer1_outputs(10051) <= a;
    layer1_outputs(10052) <= b and not a;
    layer1_outputs(10053) <= '1';
    layer1_outputs(10054) <= not a;
    layer1_outputs(10055) <= not a;
    layer1_outputs(10056) <= '0';
    layer1_outputs(10057) <= not a;
    layer1_outputs(10058) <= not b or a;
    layer1_outputs(10059) <= a xor b;
    layer1_outputs(10060) <= '1';
    layer1_outputs(10061) <= '0';
    layer1_outputs(10062) <= '1';
    layer1_outputs(10063) <= '1';
    layer1_outputs(10064) <= a xor b;
    layer1_outputs(10065) <= a;
    layer1_outputs(10066) <= a xor b;
    layer1_outputs(10067) <= not b;
    layer1_outputs(10068) <= not b or a;
    layer1_outputs(10069) <= a and b;
    layer1_outputs(10070) <= a and not b;
    layer1_outputs(10071) <= b;
    layer1_outputs(10072) <= '1';
    layer1_outputs(10073) <= not a;
    layer1_outputs(10074) <= '0';
    layer1_outputs(10075) <= not a or b;
    layer1_outputs(10076) <= b;
    layer1_outputs(10077) <= b;
    layer1_outputs(10078) <= '0';
    layer1_outputs(10079) <= '1';
    layer1_outputs(10080) <= not (a xor b);
    layer1_outputs(10081) <= '0';
    layer1_outputs(10082) <= not (a and b);
    layer1_outputs(10083) <= a or b;
    layer1_outputs(10084) <= b;
    layer1_outputs(10085) <= a;
    layer1_outputs(10086) <= '1';
    layer1_outputs(10087) <= a and b;
    layer1_outputs(10088) <= not a;
    layer1_outputs(10089) <= not (a xor b);
    layer1_outputs(10090) <= a;
    layer1_outputs(10091) <= '0';
    layer1_outputs(10092) <= a;
    layer1_outputs(10093) <= a and b;
    layer1_outputs(10094) <= a;
    layer1_outputs(10095) <= b;
    layer1_outputs(10096) <= not a or b;
    layer1_outputs(10097) <= not b or a;
    layer1_outputs(10098) <= a and b;
    layer1_outputs(10099) <= a and b;
    layer1_outputs(10100) <= a and not b;
    layer1_outputs(10101) <= '0';
    layer1_outputs(10102) <= a;
    layer1_outputs(10103) <= not b or a;
    layer1_outputs(10104) <= not a;
    layer1_outputs(10105) <= a and not b;
    layer1_outputs(10106) <= not (a or b);
    layer1_outputs(10107) <= '0';
    layer1_outputs(10108) <= '0';
    layer1_outputs(10109) <= a or b;
    layer1_outputs(10110) <= '0';
    layer1_outputs(10111) <= not a or b;
    layer1_outputs(10112) <= a or b;
    layer1_outputs(10113) <= not a;
    layer1_outputs(10114) <= a xor b;
    layer1_outputs(10115) <= a and b;
    layer1_outputs(10116) <= b;
    layer1_outputs(10117) <= not b;
    layer1_outputs(10118) <= b;
    layer1_outputs(10119) <= not (a and b);
    layer1_outputs(10120) <= not b;
    layer1_outputs(10121) <= not b;
    layer1_outputs(10122) <= not (a and b);
    layer1_outputs(10123) <= not (a or b);
    layer1_outputs(10124) <= '1';
    layer1_outputs(10125) <= not a;
    layer1_outputs(10126) <= a and b;
    layer1_outputs(10127) <= not b or a;
    layer1_outputs(10128) <= a or b;
    layer1_outputs(10129) <= b and not a;
    layer1_outputs(10130) <= not a or b;
    layer1_outputs(10131) <= a;
    layer1_outputs(10132) <= not a;
    layer1_outputs(10133) <= '0';
    layer1_outputs(10134) <= not b or a;
    layer1_outputs(10135) <= b and not a;
    layer1_outputs(10136) <= not b;
    layer1_outputs(10137) <= not b;
    layer1_outputs(10138) <= not a;
    layer1_outputs(10139) <= a;
    layer1_outputs(10140) <= not b;
    layer1_outputs(10141) <= a and b;
    layer1_outputs(10142) <= a;
    layer1_outputs(10143) <= not (a or b);
    layer1_outputs(10144) <= '0';
    layer1_outputs(10145) <= a or b;
    layer1_outputs(10146) <= b and not a;
    layer1_outputs(10147) <= a xor b;
    layer1_outputs(10148) <= not a or b;
    layer1_outputs(10149) <= '1';
    layer1_outputs(10150) <= not a or b;
    layer1_outputs(10151) <= b;
    layer1_outputs(10152) <= not (a xor b);
    layer1_outputs(10153) <= not b;
    layer1_outputs(10154) <= not a;
    layer1_outputs(10155) <= b and not a;
    layer1_outputs(10156) <= a;
    layer1_outputs(10157) <= not (a and b);
    layer1_outputs(10158) <= '1';
    layer1_outputs(10159) <= not a or b;
    layer1_outputs(10160) <= not b or a;
    layer1_outputs(10161) <= a or b;
    layer1_outputs(10162) <= a or b;
    layer1_outputs(10163) <= a or b;
    layer1_outputs(10164) <= not b or a;
    layer1_outputs(10165) <= not (a or b);
    layer1_outputs(10166) <= not a or b;
    layer1_outputs(10167) <= a and not b;
    layer1_outputs(10168) <= a;
    layer1_outputs(10169) <= a;
    layer1_outputs(10170) <= not a;
    layer1_outputs(10171) <= a or b;
    layer1_outputs(10172) <= not b or a;
    layer1_outputs(10173) <= a and b;
    layer1_outputs(10174) <= not a;
    layer1_outputs(10175) <= '0';
    layer1_outputs(10176) <= not (a and b);
    layer1_outputs(10177) <= a or b;
    layer1_outputs(10178) <= not (a xor b);
    layer1_outputs(10179) <= not a;
    layer1_outputs(10180) <= b;
    layer1_outputs(10181) <= not b or a;
    layer1_outputs(10182) <= not a or b;
    layer1_outputs(10183) <= not a or b;
    layer1_outputs(10184) <= not (a xor b);
    layer1_outputs(10185) <= a;
    layer1_outputs(10186) <= not a or b;
    layer1_outputs(10187) <= '1';
    layer1_outputs(10188) <= a or b;
    layer1_outputs(10189) <= not (a or b);
    layer1_outputs(10190) <= not b;
    layer1_outputs(10191) <= not b;
    layer1_outputs(10192) <= '0';
    layer1_outputs(10193) <= b and not a;
    layer1_outputs(10194) <= b;
    layer1_outputs(10195) <= a;
    layer1_outputs(10196) <= not a or b;
    layer1_outputs(10197) <= a;
    layer1_outputs(10198) <= b;
    layer1_outputs(10199) <= b and not a;
    layer1_outputs(10200) <= a and b;
    layer1_outputs(10201) <= not a or b;
    layer1_outputs(10202) <= not (a and b);
    layer1_outputs(10203) <= a;
    layer1_outputs(10204) <= not (a or b);
    layer1_outputs(10205) <= not (a or b);
    layer1_outputs(10206) <= a and b;
    layer1_outputs(10207) <= '0';
    layer1_outputs(10208) <= a or b;
    layer1_outputs(10209) <= b and not a;
    layer1_outputs(10210) <= not (a and b);
    layer1_outputs(10211) <= not a;
    layer1_outputs(10212) <= b;
    layer1_outputs(10213) <= not a;
    layer1_outputs(10214) <= not b;
    layer1_outputs(10215) <= '1';
    layer1_outputs(10216) <= b and not a;
    layer1_outputs(10217) <= not a;
    layer1_outputs(10218) <= a and not b;
    layer1_outputs(10219) <= '1';
    layer1_outputs(10220) <= a and not b;
    layer1_outputs(10221) <= b and not a;
    layer1_outputs(10222) <= b;
    layer1_outputs(10223) <= not b or a;
    layer1_outputs(10224) <= a and b;
    layer1_outputs(10225) <= not (a and b);
    layer1_outputs(10226) <= a and not b;
    layer1_outputs(10227) <= not a;
    layer1_outputs(10228) <= a xor b;
    layer1_outputs(10229) <= not b;
    layer1_outputs(10230) <= not a;
    layer1_outputs(10231) <= a and not b;
    layer1_outputs(10232) <= not a or b;
    layer1_outputs(10233) <= not (a xor b);
    layer1_outputs(10234) <= a and not b;
    layer1_outputs(10235) <= '0';
    layer1_outputs(10236) <= '1';
    layer1_outputs(10237) <= a and not b;
    layer1_outputs(10238) <= a or b;
    layer1_outputs(10239) <= not a or b;
    layer1_outputs(10240) <= not (a or b);
    layer1_outputs(10241) <= a or b;
    layer1_outputs(10242) <= a and b;
    layer1_outputs(10243) <= a and not b;
    layer1_outputs(10244) <= a;
    layer1_outputs(10245) <= '0';
    layer1_outputs(10246) <= not (a or b);
    layer1_outputs(10247) <= b;
    layer1_outputs(10248) <= not a;
    layer1_outputs(10249) <= a xor b;
    layer1_outputs(10250) <= not a or b;
    layer1_outputs(10251) <= not a or b;
    layer1_outputs(10252) <= a;
    layer1_outputs(10253) <= b;
    layer1_outputs(10254) <= '0';
    layer1_outputs(10255) <= b and not a;
    layer1_outputs(10256) <= a;
    layer1_outputs(10257) <= a and b;
    layer1_outputs(10258) <= not (a and b);
    layer1_outputs(10259) <= a;
    layer1_outputs(10260) <= not (a and b);
    layer1_outputs(10261) <= not (a and b);
    layer1_outputs(10262) <= a xor b;
    layer1_outputs(10263) <= a and not b;
    layer1_outputs(10264) <= not a;
    layer1_outputs(10265) <= a;
    layer1_outputs(10266) <= '0';
    layer1_outputs(10267) <= a and b;
    layer1_outputs(10268) <= b;
    layer1_outputs(10269) <= '0';
    layer1_outputs(10270) <= a or b;
    layer1_outputs(10271) <= '1';
    layer1_outputs(10272) <= a;
    layer1_outputs(10273) <= not b;
    layer1_outputs(10274) <= a or b;
    layer1_outputs(10275) <= '1';
    layer1_outputs(10276) <= b and not a;
    layer1_outputs(10277) <= not a;
    layer1_outputs(10278) <= not (a or b);
    layer1_outputs(10279) <= a and b;
    layer1_outputs(10280) <= not a or b;
    layer1_outputs(10281) <= not a or b;
    layer1_outputs(10282) <= a or b;
    layer1_outputs(10283) <= not a or b;
    layer1_outputs(10284) <= not a or b;
    layer1_outputs(10285) <= '1';
    layer1_outputs(10286) <= not (a and b);
    layer1_outputs(10287) <= b and not a;
    layer1_outputs(10288) <= b;
    layer1_outputs(10289) <= a or b;
    layer1_outputs(10290) <= a and not b;
    layer1_outputs(10291) <= a and b;
    layer1_outputs(10292) <= b;
    layer1_outputs(10293) <= a xor b;
    layer1_outputs(10294) <= a;
    layer1_outputs(10295) <= a or b;
    layer1_outputs(10296) <= a and not b;
    layer1_outputs(10297) <= not (a and b);
    layer1_outputs(10298) <= not a or b;
    layer1_outputs(10299) <= not (a or b);
    layer1_outputs(10300) <= b;
    layer1_outputs(10301) <= not b;
    layer1_outputs(10302) <= not a;
    layer1_outputs(10303) <= '1';
    layer1_outputs(10304) <= '0';
    layer1_outputs(10305) <= a;
    layer1_outputs(10306) <= not a;
    layer1_outputs(10307) <= not a;
    layer1_outputs(10308) <= a and b;
    layer1_outputs(10309) <= '0';
    layer1_outputs(10310) <= a;
    layer1_outputs(10311) <= not a;
    layer1_outputs(10312) <= a and b;
    layer1_outputs(10313) <= not b;
    layer1_outputs(10314) <= a;
    layer1_outputs(10315) <= '1';
    layer1_outputs(10316) <= not b or a;
    layer1_outputs(10317) <= '1';
    layer1_outputs(10318) <= a xor b;
    layer1_outputs(10319) <= a;
    layer1_outputs(10320) <= not a;
    layer1_outputs(10321) <= b;
    layer1_outputs(10322) <= not (a and b);
    layer1_outputs(10323) <= not b;
    layer1_outputs(10324) <= a or b;
    layer1_outputs(10325) <= not (a and b);
    layer1_outputs(10326) <= not a;
    layer1_outputs(10327) <= a xor b;
    layer1_outputs(10328) <= not (a or b);
    layer1_outputs(10329) <= a and b;
    layer1_outputs(10330) <= not (a xor b);
    layer1_outputs(10331) <= a and b;
    layer1_outputs(10332) <= a and not b;
    layer1_outputs(10333) <= not (a or b);
    layer1_outputs(10334) <= not b or a;
    layer1_outputs(10335) <= b and not a;
    layer1_outputs(10336) <= a;
    layer1_outputs(10337) <= '0';
    layer1_outputs(10338) <= '1';
    layer1_outputs(10339) <= a and b;
    layer1_outputs(10340) <= not b;
    layer1_outputs(10341) <= a and not b;
    layer1_outputs(10342) <= a;
    layer1_outputs(10343) <= not b or a;
    layer1_outputs(10344) <= not a or b;
    layer1_outputs(10345) <= a xor b;
    layer1_outputs(10346) <= not b;
    layer1_outputs(10347) <= a and not b;
    layer1_outputs(10348) <= b;
    layer1_outputs(10349) <= a and b;
    layer1_outputs(10350) <= not a or b;
    layer1_outputs(10351) <= '1';
    layer1_outputs(10352) <= a xor b;
    layer1_outputs(10353) <= a xor b;
    layer1_outputs(10354) <= not a or b;
    layer1_outputs(10355) <= not b;
    layer1_outputs(10356) <= b;
    layer1_outputs(10357) <= not (a and b);
    layer1_outputs(10358) <= a or b;
    layer1_outputs(10359) <= not b or a;
    layer1_outputs(10360) <= not b or a;
    layer1_outputs(10361) <= not b or a;
    layer1_outputs(10362) <= a and b;
    layer1_outputs(10363) <= not a;
    layer1_outputs(10364) <= a and b;
    layer1_outputs(10365) <= a or b;
    layer1_outputs(10366) <= b;
    layer1_outputs(10367) <= not (a and b);
    layer1_outputs(10368) <= not (a or b);
    layer1_outputs(10369) <= not b or a;
    layer1_outputs(10370) <= not (a and b);
    layer1_outputs(10371) <= '1';
    layer1_outputs(10372) <= not (a xor b);
    layer1_outputs(10373) <= not b;
    layer1_outputs(10374) <= b and not a;
    layer1_outputs(10375) <= a and b;
    layer1_outputs(10376) <= '1';
    layer1_outputs(10377) <= not (a or b);
    layer1_outputs(10378) <= not (a xor b);
    layer1_outputs(10379) <= a;
    layer1_outputs(10380) <= a xor b;
    layer1_outputs(10381) <= not (a and b);
    layer1_outputs(10382) <= a or b;
    layer1_outputs(10383) <= not a or b;
    layer1_outputs(10384) <= '0';
    layer1_outputs(10385) <= a;
    layer1_outputs(10386) <= not b;
    layer1_outputs(10387) <= b and not a;
    layer1_outputs(10388) <= not a or b;
    layer1_outputs(10389) <= not a;
    layer1_outputs(10390) <= a;
    layer1_outputs(10391) <= not a;
    layer1_outputs(10392) <= a or b;
    layer1_outputs(10393) <= b and not a;
    layer1_outputs(10394) <= not b;
    layer1_outputs(10395) <= a and b;
    layer1_outputs(10396) <= not b;
    layer1_outputs(10397) <= not b;
    layer1_outputs(10398) <= not (a and b);
    layer1_outputs(10399) <= a and b;
    layer1_outputs(10400) <= not b;
    layer1_outputs(10401) <= not b;
    layer1_outputs(10402) <= not a or b;
    layer1_outputs(10403) <= a and not b;
    layer1_outputs(10404) <= not a or b;
    layer1_outputs(10405) <= not (a or b);
    layer1_outputs(10406) <= not (a or b);
    layer1_outputs(10407) <= b;
    layer1_outputs(10408) <= a and b;
    layer1_outputs(10409) <= a or b;
    layer1_outputs(10410) <= b and not a;
    layer1_outputs(10411) <= '0';
    layer1_outputs(10412) <= '0';
    layer1_outputs(10413) <= a and not b;
    layer1_outputs(10414) <= a or b;
    layer1_outputs(10415) <= not (a xor b);
    layer1_outputs(10416) <= b and not a;
    layer1_outputs(10417) <= not a;
    layer1_outputs(10418) <= a and b;
    layer1_outputs(10419) <= not (a and b);
    layer1_outputs(10420) <= a or b;
    layer1_outputs(10421) <= a or b;
    layer1_outputs(10422) <= not a or b;
    layer1_outputs(10423) <= b;
    layer1_outputs(10424) <= b and not a;
    layer1_outputs(10425) <= '0';
    layer1_outputs(10426) <= not a;
    layer1_outputs(10427) <= not (a and b);
    layer1_outputs(10428) <= '1';
    layer1_outputs(10429) <= not (a or b);
    layer1_outputs(10430) <= b and not a;
    layer1_outputs(10431) <= a or b;
    layer1_outputs(10432) <= not b;
    layer1_outputs(10433) <= b and not a;
    layer1_outputs(10434) <= a and b;
    layer1_outputs(10435) <= '0';
    layer1_outputs(10436) <= a or b;
    layer1_outputs(10437) <= not a;
    layer1_outputs(10438) <= not a;
    layer1_outputs(10439) <= not b or a;
    layer1_outputs(10440) <= '1';
    layer1_outputs(10441) <= a;
    layer1_outputs(10442) <= a xor b;
    layer1_outputs(10443) <= not a;
    layer1_outputs(10444) <= a and b;
    layer1_outputs(10445) <= not b or a;
    layer1_outputs(10446) <= b;
    layer1_outputs(10447) <= not (a and b);
    layer1_outputs(10448) <= a and not b;
    layer1_outputs(10449) <= not (a and b);
    layer1_outputs(10450) <= '0';
    layer1_outputs(10451) <= a and b;
    layer1_outputs(10452) <= b and not a;
    layer1_outputs(10453) <= not (a and b);
    layer1_outputs(10454) <= not a or b;
    layer1_outputs(10455) <= '0';
    layer1_outputs(10456) <= b;
    layer1_outputs(10457) <= a;
    layer1_outputs(10458) <= a and b;
    layer1_outputs(10459) <= a;
    layer1_outputs(10460) <= not (a xor b);
    layer1_outputs(10461) <= not a;
    layer1_outputs(10462) <= b and not a;
    layer1_outputs(10463) <= not b;
    layer1_outputs(10464) <= a;
    layer1_outputs(10465) <= a and not b;
    layer1_outputs(10466) <= b;
    layer1_outputs(10467) <= b;
    layer1_outputs(10468) <= not a or b;
    layer1_outputs(10469) <= a xor b;
    layer1_outputs(10470) <= not (a or b);
    layer1_outputs(10471) <= a;
    layer1_outputs(10472) <= a and b;
    layer1_outputs(10473) <= a and b;
    layer1_outputs(10474) <= a and b;
    layer1_outputs(10475) <= '1';
    layer1_outputs(10476) <= not (a xor b);
    layer1_outputs(10477) <= b and not a;
    layer1_outputs(10478) <= a and b;
    layer1_outputs(10479) <= not (a and b);
    layer1_outputs(10480) <= b and not a;
    layer1_outputs(10481) <= not a;
    layer1_outputs(10482) <= b;
    layer1_outputs(10483) <= not (a xor b);
    layer1_outputs(10484) <= not a or b;
    layer1_outputs(10485) <= '0';
    layer1_outputs(10486) <= b and not a;
    layer1_outputs(10487) <= not b or a;
    layer1_outputs(10488) <= '0';
    layer1_outputs(10489) <= not b;
    layer1_outputs(10490) <= a xor b;
    layer1_outputs(10491) <= a and not b;
    layer1_outputs(10492) <= b and not a;
    layer1_outputs(10493) <= not a;
    layer1_outputs(10494) <= not (a and b);
    layer1_outputs(10495) <= not b or a;
    layer1_outputs(10496) <= not b or a;
    layer1_outputs(10497) <= b and not a;
    layer1_outputs(10498) <= b;
    layer1_outputs(10499) <= a or b;
    layer1_outputs(10500) <= not (a or b);
    layer1_outputs(10501) <= not a or b;
    layer1_outputs(10502) <= b and not a;
    layer1_outputs(10503) <= a or b;
    layer1_outputs(10504) <= b;
    layer1_outputs(10505) <= a and b;
    layer1_outputs(10506) <= not (a xor b);
    layer1_outputs(10507) <= a and not b;
    layer1_outputs(10508) <= not (a or b);
    layer1_outputs(10509) <= not (a and b);
    layer1_outputs(10510) <= not b;
    layer1_outputs(10511) <= b and not a;
    layer1_outputs(10512) <= '0';
    layer1_outputs(10513) <= '1';
    layer1_outputs(10514) <= not (a or b);
    layer1_outputs(10515) <= a and b;
    layer1_outputs(10516) <= a;
    layer1_outputs(10517) <= '1';
    layer1_outputs(10518) <= a;
    layer1_outputs(10519) <= not b or a;
    layer1_outputs(10520) <= not b or a;
    layer1_outputs(10521) <= not (a or b);
    layer1_outputs(10522) <= a and b;
    layer1_outputs(10523) <= not (a and b);
    layer1_outputs(10524) <= not b;
    layer1_outputs(10525) <= a;
    layer1_outputs(10526) <= not b;
    layer1_outputs(10527) <= a and not b;
    layer1_outputs(10528) <= not a or b;
    layer1_outputs(10529) <= not (a or b);
    layer1_outputs(10530) <= a and b;
    layer1_outputs(10531) <= b and not a;
    layer1_outputs(10532) <= a;
    layer1_outputs(10533) <= a and not b;
    layer1_outputs(10534) <= '0';
    layer1_outputs(10535) <= not a or b;
    layer1_outputs(10536) <= not (a xor b);
    layer1_outputs(10537) <= not b;
    layer1_outputs(10538) <= b and not a;
    layer1_outputs(10539) <= not a or b;
    layer1_outputs(10540) <= b and not a;
    layer1_outputs(10541) <= b;
    layer1_outputs(10542) <= b;
    layer1_outputs(10543) <= b;
    layer1_outputs(10544) <= not a;
    layer1_outputs(10545) <= not a;
    layer1_outputs(10546) <= a and not b;
    layer1_outputs(10547) <= not a;
    layer1_outputs(10548) <= '0';
    layer1_outputs(10549) <= not a or b;
    layer1_outputs(10550) <= not b;
    layer1_outputs(10551) <= a and b;
    layer1_outputs(10552) <= not a;
    layer1_outputs(10553) <= not b or a;
    layer1_outputs(10554) <= '0';
    layer1_outputs(10555) <= b;
    layer1_outputs(10556) <= not a or b;
    layer1_outputs(10557) <= '1';
    layer1_outputs(10558) <= not (a or b);
    layer1_outputs(10559) <= a and not b;
    layer1_outputs(10560) <= not (a xor b);
    layer1_outputs(10561) <= a and b;
    layer1_outputs(10562) <= a or b;
    layer1_outputs(10563) <= not (a or b);
    layer1_outputs(10564) <= '1';
    layer1_outputs(10565) <= b and not a;
    layer1_outputs(10566) <= a;
    layer1_outputs(10567) <= not (a xor b);
    layer1_outputs(10568) <= not (a or b);
    layer1_outputs(10569) <= b and not a;
    layer1_outputs(10570) <= not (a xor b);
    layer1_outputs(10571) <= not (a xor b);
    layer1_outputs(10572) <= b;
    layer1_outputs(10573) <= not a;
    layer1_outputs(10574) <= a or b;
    layer1_outputs(10575) <= b;
    layer1_outputs(10576) <= not b;
    layer1_outputs(10577) <= a and not b;
    layer1_outputs(10578) <= a;
    layer1_outputs(10579) <= b;
    layer1_outputs(10580) <= not a or b;
    layer1_outputs(10581) <= a and b;
    layer1_outputs(10582) <= a and b;
    layer1_outputs(10583) <= not a;
    layer1_outputs(10584) <= '0';
    layer1_outputs(10585) <= a and not b;
    layer1_outputs(10586) <= b;
    layer1_outputs(10587) <= not b or a;
    layer1_outputs(10588) <= not a or b;
    layer1_outputs(10589) <= a;
    layer1_outputs(10590) <= not b;
    layer1_outputs(10591) <= not (a xor b);
    layer1_outputs(10592) <= not a or b;
    layer1_outputs(10593) <= not (a or b);
    layer1_outputs(10594) <= not (a xor b);
    layer1_outputs(10595) <= b;
    layer1_outputs(10596) <= a;
    layer1_outputs(10597) <= b;
    layer1_outputs(10598) <= not b or a;
    layer1_outputs(10599) <= '1';
    layer1_outputs(10600) <= a and not b;
    layer1_outputs(10601) <= a xor b;
    layer1_outputs(10602) <= not b or a;
    layer1_outputs(10603) <= not a;
    layer1_outputs(10604) <= b;
    layer1_outputs(10605) <= '1';
    layer1_outputs(10606) <= b;
    layer1_outputs(10607) <= '0';
    layer1_outputs(10608) <= a;
    layer1_outputs(10609) <= not (a or b);
    layer1_outputs(10610) <= a and b;
    layer1_outputs(10611) <= a and b;
    layer1_outputs(10612) <= b and not a;
    layer1_outputs(10613) <= '0';
    layer1_outputs(10614) <= b;
    layer1_outputs(10615) <= a or b;
    layer1_outputs(10616) <= not b;
    layer1_outputs(10617) <= not a or b;
    layer1_outputs(10618) <= '1';
    layer1_outputs(10619) <= not b or a;
    layer1_outputs(10620) <= a;
    layer1_outputs(10621) <= not a;
    layer1_outputs(10622) <= not a or b;
    layer1_outputs(10623) <= a and b;
    layer1_outputs(10624) <= not (a xor b);
    layer1_outputs(10625) <= b and not a;
    layer1_outputs(10626) <= not (a xor b);
    layer1_outputs(10627) <= a or b;
    layer1_outputs(10628) <= not a;
    layer1_outputs(10629) <= b;
    layer1_outputs(10630) <= not (a or b);
    layer1_outputs(10631) <= b and not a;
    layer1_outputs(10632) <= not (a and b);
    layer1_outputs(10633) <= not a or b;
    layer1_outputs(10634) <= not a;
    layer1_outputs(10635) <= not a;
    layer1_outputs(10636) <= not (a and b);
    layer1_outputs(10637) <= not b;
    layer1_outputs(10638) <= b;
    layer1_outputs(10639) <= '1';
    layer1_outputs(10640) <= not a;
    layer1_outputs(10641) <= '0';
    layer1_outputs(10642) <= '1';
    layer1_outputs(10643) <= a;
    layer1_outputs(10644) <= not a;
    layer1_outputs(10645) <= b and not a;
    layer1_outputs(10646) <= a xor b;
    layer1_outputs(10647) <= not a;
    layer1_outputs(10648) <= not (a and b);
    layer1_outputs(10649) <= a and not b;
    layer1_outputs(10650) <= not (a or b);
    layer1_outputs(10651) <= not b;
    layer1_outputs(10652) <= a;
    layer1_outputs(10653) <= b and not a;
    layer1_outputs(10654) <= a xor b;
    layer1_outputs(10655) <= '1';
    layer1_outputs(10656) <= a or b;
    layer1_outputs(10657) <= '0';
    layer1_outputs(10658) <= a and not b;
    layer1_outputs(10659) <= not b;
    layer1_outputs(10660) <= not b or a;
    layer1_outputs(10661) <= a or b;
    layer1_outputs(10662) <= '0';
    layer1_outputs(10663) <= not (a xor b);
    layer1_outputs(10664) <= a;
    layer1_outputs(10665) <= not a or b;
    layer1_outputs(10666) <= a and not b;
    layer1_outputs(10667) <= not a or b;
    layer1_outputs(10668) <= not a or b;
    layer1_outputs(10669) <= b;
    layer1_outputs(10670) <= '1';
    layer1_outputs(10671) <= a and not b;
    layer1_outputs(10672) <= not (a and b);
    layer1_outputs(10673) <= a and not b;
    layer1_outputs(10674) <= not b;
    layer1_outputs(10675) <= a;
    layer1_outputs(10676) <= b and not a;
    layer1_outputs(10677) <= not (a or b);
    layer1_outputs(10678) <= '1';
    layer1_outputs(10679) <= not (a or b);
    layer1_outputs(10680) <= not b or a;
    layer1_outputs(10681) <= not a;
    layer1_outputs(10682) <= '0';
    layer1_outputs(10683) <= a and not b;
    layer1_outputs(10684) <= not (a or b);
    layer1_outputs(10685) <= '1';
    layer1_outputs(10686) <= not b;
    layer1_outputs(10687) <= b and not a;
    layer1_outputs(10688) <= a xor b;
    layer1_outputs(10689) <= not b;
    layer1_outputs(10690) <= a and b;
    layer1_outputs(10691) <= a;
    layer1_outputs(10692) <= a or b;
    layer1_outputs(10693) <= a xor b;
    layer1_outputs(10694) <= a or b;
    layer1_outputs(10695) <= not b or a;
    layer1_outputs(10696) <= not a or b;
    layer1_outputs(10697) <= a or b;
    layer1_outputs(10698) <= '0';
    layer1_outputs(10699) <= not a;
    layer1_outputs(10700) <= b;
    layer1_outputs(10701) <= not a;
    layer1_outputs(10702) <= not (a and b);
    layer1_outputs(10703) <= b and not a;
    layer1_outputs(10704) <= not (a or b);
    layer1_outputs(10705) <= '0';
    layer1_outputs(10706) <= a;
    layer1_outputs(10707) <= a;
    layer1_outputs(10708) <= '1';
    layer1_outputs(10709) <= a and b;
    layer1_outputs(10710) <= a or b;
    layer1_outputs(10711) <= b;
    layer1_outputs(10712) <= not a or b;
    layer1_outputs(10713) <= a xor b;
    layer1_outputs(10714) <= not b;
    layer1_outputs(10715) <= a xor b;
    layer1_outputs(10716) <= '0';
    layer1_outputs(10717) <= b and not a;
    layer1_outputs(10718) <= '0';
    layer1_outputs(10719) <= b and not a;
    layer1_outputs(10720) <= not b or a;
    layer1_outputs(10721) <= not (a and b);
    layer1_outputs(10722) <= b;
    layer1_outputs(10723) <= not a or b;
    layer1_outputs(10724) <= b and not a;
    layer1_outputs(10725) <= not (a and b);
    layer1_outputs(10726) <= a;
    layer1_outputs(10727) <= not b;
    layer1_outputs(10728) <= not (a and b);
    layer1_outputs(10729) <= not (a and b);
    layer1_outputs(10730) <= b;
    layer1_outputs(10731) <= b and not a;
    layer1_outputs(10732) <= not b or a;
    layer1_outputs(10733) <= b and not a;
    layer1_outputs(10734) <= a and not b;
    layer1_outputs(10735) <= b;
    layer1_outputs(10736) <= b;
    layer1_outputs(10737) <= a and not b;
    layer1_outputs(10738) <= a or b;
    layer1_outputs(10739) <= a xor b;
    layer1_outputs(10740) <= not (a and b);
    layer1_outputs(10741) <= a and b;
    layer1_outputs(10742) <= a;
    layer1_outputs(10743) <= not (a and b);
    layer1_outputs(10744) <= '1';
    layer1_outputs(10745) <= not b;
    layer1_outputs(10746) <= b;
    layer1_outputs(10747) <= not (a and b);
    layer1_outputs(10748) <= b and not a;
    layer1_outputs(10749) <= a;
    layer1_outputs(10750) <= b;
    layer1_outputs(10751) <= not (a or b);
    layer1_outputs(10752) <= not a or b;
    layer1_outputs(10753) <= not a;
    layer1_outputs(10754) <= not b;
    layer1_outputs(10755) <= a and not b;
    layer1_outputs(10756) <= not a;
    layer1_outputs(10757) <= a or b;
    layer1_outputs(10758) <= b;
    layer1_outputs(10759) <= a and b;
    layer1_outputs(10760) <= not a;
    layer1_outputs(10761) <= '1';
    layer1_outputs(10762) <= a and not b;
    layer1_outputs(10763) <= a;
    layer1_outputs(10764) <= '0';
    layer1_outputs(10765) <= a or b;
    layer1_outputs(10766) <= not (a or b);
    layer1_outputs(10767) <= b and not a;
    layer1_outputs(10768) <= not (a and b);
    layer1_outputs(10769) <= not a or b;
    layer1_outputs(10770) <= a or b;
    layer1_outputs(10771) <= a xor b;
    layer1_outputs(10772) <= '1';
    layer1_outputs(10773) <= not (a and b);
    layer1_outputs(10774) <= not (a and b);
    layer1_outputs(10775) <= a;
    layer1_outputs(10776) <= not b or a;
    layer1_outputs(10777) <= a and not b;
    layer1_outputs(10778) <= '0';
    layer1_outputs(10779) <= not (a xor b);
    layer1_outputs(10780) <= a and b;
    layer1_outputs(10781) <= '1';
    layer1_outputs(10782) <= b;
    layer1_outputs(10783) <= '1';
    layer1_outputs(10784) <= not (a or b);
    layer1_outputs(10785) <= not (a or b);
    layer1_outputs(10786) <= not b;
    layer1_outputs(10787) <= '0';
    layer1_outputs(10788) <= a and b;
    layer1_outputs(10789) <= a and not b;
    layer1_outputs(10790) <= '0';
    layer1_outputs(10791) <= '0';
    layer1_outputs(10792) <= not (a and b);
    layer1_outputs(10793) <= not a or b;
    layer1_outputs(10794) <= not b or a;
    layer1_outputs(10795) <= not b or a;
    layer1_outputs(10796) <= '0';
    layer1_outputs(10797) <= not a or b;
    layer1_outputs(10798) <= a;
    layer1_outputs(10799) <= a and not b;
    layer1_outputs(10800) <= b and not a;
    layer1_outputs(10801) <= b and not a;
    layer1_outputs(10802) <= not b or a;
    layer1_outputs(10803) <= not b or a;
    layer1_outputs(10804) <= a xor b;
    layer1_outputs(10805) <= a and not b;
    layer1_outputs(10806) <= a;
    layer1_outputs(10807) <= '0';
    layer1_outputs(10808) <= a or b;
    layer1_outputs(10809) <= not b or a;
    layer1_outputs(10810) <= '1';
    layer1_outputs(10811) <= not (a and b);
    layer1_outputs(10812) <= b;
    layer1_outputs(10813) <= '1';
    layer1_outputs(10814) <= not (a or b);
    layer1_outputs(10815) <= a and b;
    layer1_outputs(10816) <= not b or a;
    layer1_outputs(10817) <= not b;
    layer1_outputs(10818) <= not b or a;
    layer1_outputs(10819) <= a and b;
    layer1_outputs(10820) <= a and not b;
    layer1_outputs(10821) <= a and not b;
    layer1_outputs(10822) <= not (a or b);
    layer1_outputs(10823) <= a and not b;
    layer1_outputs(10824) <= b;
    layer1_outputs(10825) <= not (a or b);
    layer1_outputs(10826) <= not b;
    layer1_outputs(10827) <= not b or a;
    layer1_outputs(10828) <= a and not b;
    layer1_outputs(10829) <= a and b;
    layer1_outputs(10830) <= '0';
    layer1_outputs(10831) <= a or b;
    layer1_outputs(10832) <= a and b;
    layer1_outputs(10833) <= not a or b;
    layer1_outputs(10834) <= not (a or b);
    layer1_outputs(10835) <= a and b;
    layer1_outputs(10836) <= not a;
    layer1_outputs(10837) <= a xor b;
    layer1_outputs(10838) <= '1';
    layer1_outputs(10839) <= '0';
    layer1_outputs(10840) <= b and not a;
    layer1_outputs(10841) <= not (a and b);
    layer1_outputs(10842) <= '0';
    layer1_outputs(10843) <= a and not b;
    layer1_outputs(10844) <= b and not a;
    layer1_outputs(10845) <= a and not b;
    layer1_outputs(10846) <= a and not b;
    layer1_outputs(10847) <= a and b;
    layer1_outputs(10848) <= '0';
    layer1_outputs(10849) <= not b;
    layer1_outputs(10850) <= not b or a;
    layer1_outputs(10851) <= not b or a;
    layer1_outputs(10852) <= b and not a;
    layer1_outputs(10853) <= a and not b;
    layer1_outputs(10854) <= '0';
    layer1_outputs(10855) <= not a or b;
    layer1_outputs(10856) <= b;
    layer1_outputs(10857) <= a and not b;
    layer1_outputs(10858) <= not b;
    layer1_outputs(10859) <= not b;
    layer1_outputs(10860) <= '1';
    layer1_outputs(10861) <= not b;
    layer1_outputs(10862) <= a and not b;
    layer1_outputs(10863) <= not b or a;
    layer1_outputs(10864) <= a and b;
    layer1_outputs(10865) <= b;
    layer1_outputs(10866) <= not b;
    layer1_outputs(10867) <= not (a or b);
    layer1_outputs(10868) <= b;
    layer1_outputs(10869) <= not b or a;
    layer1_outputs(10870) <= not b or a;
    layer1_outputs(10871) <= a;
    layer1_outputs(10872) <= not (a xor b);
    layer1_outputs(10873) <= a xor b;
    layer1_outputs(10874) <= a;
    layer1_outputs(10875) <= not b or a;
    layer1_outputs(10876) <= b and not a;
    layer1_outputs(10877) <= not (a or b);
    layer1_outputs(10878) <= a and b;
    layer1_outputs(10879) <= b and not a;
    layer1_outputs(10880) <= b and not a;
    layer1_outputs(10881) <= not (a and b);
    layer1_outputs(10882) <= a or b;
    layer1_outputs(10883) <= '0';
    layer1_outputs(10884) <= '1';
    layer1_outputs(10885) <= a;
    layer1_outputs(10886) <= not b;
    layer1_outputs(10887) <= a;
    layer1_outputs(10888) <= not (a or b);
    layer1_outputs(10889) <= not (a xor b);
    layer1_outputs(10890) <= not b or a;
    layer1_outputs(10891) <= b and not a;
    layer1_outputs(10892) <= not b or a;
    layer1_outputs(10893) <= a;
    layer1_outputs(10894) <= '1';
    layer1_outputs(10895) <= not a or b;
    layer1_outputs(10896) <= a and b;
    layer1_outputs(10897) <= not (a and b);
    layer1_outputs(10898) <= '1';
    layer1_outputs(10899) <= not a or b;
    layer1_outputs(10900) <= b;
    layer1_outputs(10901) <= not b or a;
    layer1_outputs(10902) <= a and not b;
    layer1_outputs(10903) <= a or b;
    layer1_outputs(10904) <= a;
    layer1_outputs(10905) <= '1';
    layer1_outputs(10906) <= a or b;
    layer1_outputs(10907) <= not (a or b);
    layer1_outputs(10908) <= not b or a;
    layer1_outputs(10909) <= a and not b;
    layer1_outputs(10910) <= not b or a;
    layer1_outputs(10911) <= a or b;
    layer1_outputs(10912) <= not a or b;
    layer1_outputs(10913) <= '1';
    layer1_outputs(10914) <= a or b;
    layer1_outputs(10915) <= a and b;
    layer1_outputs(10916) <= not b or a;
    layer1_outputs(10917) <= a or b;
    layer1_outputs(10918) <= not b;
    layer1_outputs(10919) <= b and not a;
    layer1_outputs(10920) <= not b or a;
    layer1_outputs(10921) <= a or b;
    layer1_outputs(10922) <= '1';
    layer1_outputs(10923) <= a and not b;
    layer1_outputs(10924) <= b;
    layer1_outputs(10925) <= b;
    layer1_outputs(10926) <= '1';
    layer1_outputs(10927) <= not b;
    layer1_outputs(10928) <= a;
    layer1_outputs(10929) <= not a;
    layer1_outputs(10930) <= a or b;
    layer1_outputs(10931) <= a xor b;
    layer1_outputs(10932) <= not b or a;
    layer1_outputs(10933) <= b and not a;
    layer1_outputs(10934) <= not b;
    layer1_outputs(10935) <= a;
    layer1_outputs(10936) <= '0';
    layer1_outputs(10937) <= b and not a;
    layer1_outputs(10938) <= a and not b;
    layer1_outputs(10939) <= '0';
    layer1_outputs(10940) <= not a;
    layer1_outputs(10941) <= not b;
    layer1_outputs(10942) <= not (a or b);
    layer1_outputs(10943) <= not a or b;
    layer1_outputs(10944) <= not (a xor b);
    layer1_outputs(10945) <= not b;
    layer1_outputs(10946) <= a;
    layer1_outputs(10947) <= not a or b;
    layer1_outputs(10948) <= '0';
    layer1_outputs(10949) <= not a or b;
    layer1_outputs(10950) <= not b or a;
    layer1_outputs(10951) <= a xor b;
    layer1_outputs(10952) <= not (a and b);
    layer1_outputs(10953) <= b;
    layer1_outputs(10954) <= not a;
    layer1_outputs(10955) <= a or b;
    layer1_outputs(10956) <= a or b;
    layer1_outputs(10957) <= a or b;
    layer1_outputs(10958) <= not a;
    layer1_outputs(10959) <= not (a and b);
    layer1_outputs(10960) <= not b;
    layer1_outputs(10961) <= '0';
    layer1_outputs(10962) <= a or b;
    layer1_outputs(10963) <= not a or b;
    layer1_outputs(10964) <= not b;
    layer1_outputs(10965) <= not (a xor b);
    layer1_outputs(10966) <= not b;
    layer1_outputs(10967) <= not b or a;
    layer1_outputs(10968) <= a and not b;
    layer1_outputs(10969) <= not (a or b);
    layer1_outputs(10970) <= a or b;
    layer1_outputs(10971) <= '0';
    layer1_outputs(10972) <= not (a xor b);
    layer1_outputs(10973) <= '0';
    layer1_outputs(10974) <= a and b;
    layer1_outputs(10975) <= not (a xor b);
    layer1_outputs(10976) <= a and b;
    layer1_outputs(10977) <= not (a or b);
    layer1_outputs(10978) <= b;
    layer1_outputs(10979) <= b and not a;
    layer1_outputs(10980) <= a and not b;
    layer1_outputs(10981) <= not (a and b);
    layer1_outputs(10982) <= a;
    layer1_outputs(10983) <= not b or a;
    layer1_outputs(10984) <= not b;
    layer1_outputs(10985) <= a or b;
    layer1_outputs(10986) <= not a;
    layer1_outputs(10987) <= a and b;
    layer1_outputs(10988) <= not a or b;
    layer1_outputs(10989) <= b and not a;
    layer1_outputs(10990) <= a;
    layer1_outputs(10991) <= '0';
    layer1_outputs(10992) <= not b;
    layer1_outputs(10993) <= not b or a;
    layer1_outputs(10994) <= a and b;
    layer1_outputs(10995) <= not b or a;
    layer1_outputs(10996) <= a and not b;
    layer1_outputs(10997) <= not (a and b);
    layer1_outputs(10998) <= not b or a;
    layer1_outputs(10999) <= a;
    layer1_outputs(11000) <= a;
    layer1_outputs(11001) <= not (a and b);
    layer1_outputs(11002) <= '0';
    layer1_outputs(11003) <= a and b;
    layer1_outputs(11004) <= not (a xor b);
    layer1_outputs(11005) <= b and not a;
    layer1_outputs(11006) <= a and b;
    layer1_outputs(11007) <= '1';
    layer1_outputs(11008) <= not b or a;
    layer1_outputs(11009) <= b and not a;
    layer1_outputs(11010) <= not a or b;
    layer1_outputs(11011) <= a and b;
    layer1_outputs(11012) <= '0';
    layer1_outputs(11013) <= '0';
    layer1_outputs(11014) <= not b;
    layer1_outputs(11015) <= not (a xor b);
    layer1_outputs(11016) <= b and not a;
    layer1_outputs(11017) <= not (a or b);
    layer1_outputs(11018) <= '1';
    layer1_outputs(11019) <= a;
    layer1_outputs(11020) <= a;
    layer1_outputs(11021) <= a and b;
    layer1_outputs(11022) <= a or b;
    layer1_outputs(11023) <= a and b;
    layer1_outputs(11024) <= a;
    layer1_outputs(11025) <= a;
    layer1_outputs(11026) <= not (a or b);
    layer1_outputs(11027) <= not b or a;
    layer1_outputs(11028) <= not a;
    layer1_outputs(11029) <= a or b;
    layer1_outputs(11030) <= '0';
    layer1_outputs(11031) <= not (a or b);
    layer1_outputs(11032) <= '1';
    layer1_outputs(11033) <= '1';
    layer1_outputs(11034) <= '1';
    layer1_outputs(11035) <= not a or b;
    layer1_outputs(11036) <= not a or b;
    layer1_outputs(11037) <= b;
    layer1_outputs(11038) <= '0';
    layer1_outputs(11039) <= b and not a;
    layer1_outputs(11040) <= not b;
    layer1_outputs(11041) <= '1';
    layer1_outputs(11042) <= not a or b;
    layer1_outputs(11043) <= a and not b;
    layer1_outputs(11044) <= b;
    layer1_outputs(11045) <= not a or b;
    layer1_outputs(11046) <= a and b;
    layer1_outputs(11047) <= '0';
    layer1_outputs(11048) <= a;
    layer1_outputs(11049) <= a and not b;
    layer1_outputs(11050) <= b and not a;
    layer1_outputs(11051) <= not (a or b);
    layer1_outputs(11052) <= a and not b;
    layer1_outputs(11053) <= not a or b;
    layer1_outputs(11054) <= not b;
    layer1_outputs(11055) <= a and not b;
    layer1_outputs(11056) <= not a or b;
    layer1_outputs(11057) <= not (a xor b);
    layer1_outputs(11058) <= '0';
    layer1_outputs(11059) <= a and b;
    layer1_outputs(11060) <= '1';
    layer1_outputs(11061) <= a xor b;
    layer1_outputs(11062) <= a;
    layer1_outputs(11063) <= not (a xor b);
    layer1_outputs(11064) <= b;
    layer1_outputs(11065) <= a and b;
    layer1_outputs(11066) <= '1';
    layer1_outputs(11067) <= not b;
    layer1_outputs(11068) <= a;
    layer1_outputs(11069) <= a and b;
    layer1_outputs(11070) <= not b or a;
    layer1_outputs(11071) <= b and not a;
    layer1_outputs(11072) <= a or b;
    layer1_outputs(11073) <= b;
    layer1_outputs(11074) <= not b;
    layer1_outputs(11075) <= a xor b;
    layer1_outputs(11076) <= b;
    layer1_outputs(11077) <= a;
    layer1_outputs(11078) <= not (a and b);
    layer1_outputs(11079) <= not (a or b);
    layer1_outputs(11080) <= '1';
    layer1_outputs(11081) <= not (a xor b);
    layer1_outputs(11082) <= not b or a;
    layer1_outputs(11083) <= a and not b;
    layer1_outputs(11084) <= '1';
    layer1_outputs(11085) <= b and not a;
    layer1_outputs(11086) <= not b;
    layer1_outputs(11087) <= '0';
    layer1_outputs(11088) <= '1';
    layer1_outputs(11089) <= a xor b;
    layer1_outputs(11090) <= not (a or b);
    layer1_outputs(11091) <= not a or b;
    layer1_outputs(11092) <= a xor b;
    layer1_outputs(11093) <= not b or a;
    layer1_outputs(11094) <= a or b;
    layer1_outputs(11095) <= a and not b;
    layer1_outputs(11096) <= a and not b;
    layer1_outputs(11097) <= not (a or b);
    layer1_outputs(11098) <= not a;
    layer1_outputs(11099) <= a and b;
    layer1_outputs(11100) <= a or b;
    layer1_outputs(11101) <= not (a and b);
    layer1_outputs(11102) <= not a;
    layer1_outputs(11103) <= a;
    layer1_outputs(11104) <= not b;
    layer1_outputs(11105) <= b;
    layer1_outputs(11106) <= not (a and b);
    layer1_outputs(11107) <= not a or b;
    layer1_outputs(11108) <= '0';
    layer1_outputs(11109) <= b and not a;
    layer1_outputs(11110) <= not b or a;
    layer1_outputs(11111) <= b;
    layer1_outputs(11112) <= not (a xor b);
    layer1_outputs(11113) <= a;
    layer1_outputs(11114) <= not (a xor b);
    layer1_outputs(11115) <= not b or a;
    layer1_outputs(11116) <= '0';
    layer1_outputs(11117) <= not b;
    layer1_outputs(11118) <= a and b;
    layer1_outputs(11119) <= not a or b;
    layer1_outputs(11120) <= not b or a;
    layer1_outputs(11121) <= not (a or b);
    layer1_outputs(11122) <= not (a and b);
    layer1_outputs(11123) <= b;
    layer1_outputs(11124) <= a or b;
    layer1_outputs(11125) <= b and not a;
    layer1_outputs(11126) <= not b;
    layer1_outputs(11127) <= '0';
    layer1_outputs(11128) <= not (a xor b);
    layer1_outputs(11129) <= a and not b;
    layer1_outputs(11130) <= not b;
    layer1_outputs(11131) <= a xor b;
    layer1_outputs(11132) <= a and b;
    layer1_outputs(11133) <= a and not b;
    layer1_outputs(11134) <= a and b;
    layer1_outputs(11135) <= a or b;
    layer1_outputs(11136) <= not b;
    layer1_outputs(11137) <= b;
    layer1_outputs(11138) <= b and not a;
    layer1_outputs(11139) <= a;
    layer1_outputs(11140) <= a;
    layer1_outputs(11141) <= a and not b;
    layer1_outputs(11142) <= a and b;
    layer1_outputs(11143) <= a or b;
    layer1_outputs(11144) <= not b;
    layer1_outputs(11145) <= not (a xor b);
    layer1_outputs(11146) <= a and not b;
    layer1_outputs(11147) <= a xor b;
    layer1_outputs(11148) <= not (a or b);
    layer1_outputs(11149) <= b;
    layer1_outputs(11150) <= not a or b;
    layer1_outputs(11151) <= not (a or b);
    layer1_outputs(11152) <= a and not b;
    layer1_outputs(11153) <= not b or a;
    layer1_outputs(11154) <= a and b;
    layer1_outputs(11155) <= not (a or b);
    layer1_outputs(11156) <= not a;
    layer1_outputs(11157) <= '0';
    layer1_outputs(11158) <= not b or a;
    layer1_outputs(11159) <= a and not b;
    layer1_outputs(11160) <= b;
    layer1_outputs(11161) <= a or b;
    layer1_outputs(11162) <= a or b;
    layer1_outputs(11163) <= a and not b;
    layer1_outputs(11164) <= a or b;
    layer1_outputs(11165) <= a and not b;
    layer1_outputs(11166) <= a;
    layer1_outputs(11167) <= b;
    layer1_outputs(11168) <= not (a and b);
    layer1_outputs(11169) <= a and b;
    layer1_outputs(11170) <= a and b;
    layer1_outputs(11171) <= a and not b;
    layer1_outputs(11172) <= b;
    layer1_outputs(11173) <= not (a and b);
    layer1_outputs(11174) <= a and not b;
    layer1_outputs(11175) <= not (a or b);
    layer1_outputs(11176) <= a and b;
    layer1_outputs(11177) <= a or b;
    layer1_outputs(11178) <= not (a and b);
    layer1_outputs(11179) <= '0';
    layer1_outputs(11180) <= not (a or b);
    layer1_outputs(11181) <= a and b;
    layer1_outputs(11182) <= a xor b;
    layer1_outputs(11183) <= a and b;
    layer1_outputs(11184) <= b;
    layer1_outputs(11185) <= not b;
    layer1_outputs(11186) <= not b or a;
    layer1_outputs(11187) <= a;
    layer1_outputs(11188) <= a and b;
    layer1_outputs(11189) <= a or b;
    layer1_outputs(11190) <= a;
    layer1_outputs(11191) <= not (a or b);
    layer1_outputs(11192) <= '0';
    layer1_outputs(11193) <= not a;
    layer1_outputs(11194) <= not a;
    layer1_outputs(11195) <= not (a and b);
    layer1_outputs(11196) <= a or b;
    layer1_outputs(11197) <= not a;
    layer1_outputs(11198) <= a and b;
    layer1_outputs(11199) <= b;
    layer1_outputs(11200) <= not (a and b);
    layer1_outputs(11201) <= a;
    layer1_outputs(11202) <= not (a xor b);
    layer1_outputs(11203) <= '1';
    layer1_outputs(11204) <= a and not b;
    layer1_outputs(11205) <= b;
    layer1_outputs(11206) <= not b or a;
    layer1_outputs(11207) <= not (a xor b);
    layer1_outputs(11208) <= not (a or b);
    layer1_outputs(11209) <= not (a and b);
    layer1_outputs(11210) <= a and not b;
    layer1_outputs(11211) <= not (a xor b);
    layer1_outputs(11212) <= not a;
    layer1_outputs(11213) <= '0';
    layer1_outputs(11214) <= not b;
    layer1_outputs(11215) <= a and b;
    layer1_outputs(11216) <= a;
    layer1_outputs(11217) <= a and b;
    layer1_outputs(11218) <= b and not a;
    layer1_outputs(11219) <= a and b;
    layer1_outputs(11220) <= a and not b;
    layer1_outputs(11221) <= a and b;
    layer1_outputs(11222) <= not (a or b);
    layer1_outputs(11223) <= not b or a;
    layer1_outputs(11224) <= not (a xor b);
    layer1_outputs(11225) <= not a or b;
    layer1_outputs(11226) <= a and not b;
    layer1_outputs(11227) <= a or b;
    layer1_outputs(11228) <= not a or b;
    layer1_outputs(11229) <= a;
    layer1_outputs(11230) <= not b;
    layer1_outputs(11231) <= b and not a;
    layer1_outputs(11232) <= b and not a;
    layer1_outputs(11233) <= '1';
    layer1_outputs(11234) <= not (a and b);
    layer1_outputs(11235) <= '1';
    layer1_outputs(11236) <= not b;
    layer1_outputs(11237) <= not a;
    layer1_outputs(11238) <= not a;
    layer1_outputs(11239) <= a and not b;
    layer1_outputs(11240) <= a and b;
    layer1_outputs(11241) <= not a or b;
    layer1_outputs(11242) <= b and not a;
    layer1_outputs(11243) <= not (a xor b);
    layer1_outputs(11244) <= b;
    layer1_outputs(11245) <= not a;
    layer1_outputs(11246) <= not (a and b);
    layer1_outputs(11247) <= a xor b;
    layer1_outputs(11248) <= a or b;
    layer1_outputs(11249) <= not (a and b);
    layer1_outputs(11250) <= not b or a;
    layer1_outputs(11251) <= not b;
    layer1_outputs(11252) <= b;
    layer1_outputs(11253) <= a and b;
    layer1_outputs(11254) <= not b;
    layer1_outputs(11255) <= not b;
    layer1_outputs(11256) <= a xor b;
    layer1_outputs(11257) <= not (a and b);
    layer1_outputs(11258) <= a;
    layer1_outputs(11259) <= b and not a;
    layer1_outputs(11260) <= not (a xor b);
    layer1_outputs(11261) <= not a or b;
    layer1_outputs(11262) <= '1';
    layer1_outputs(11263) <= '0';
    layer1_outputs(11264) <= '0';
    layer1_outputs(11265) <= a xor b;
    layer1_outputs(11266) <= not b or a;
    layer1_outputs(11267) <= a xor b;
    layer1_outputs(11268) <= a or b;
    layer1_outputs(11269) <= a xor b;
    layer1_outputs(11270) <= not a;
    layer1_outputs(11271) <= not b;
    layer1_outputs(11272) <= '1';
    layer1_outputs(11273) <= a xor b;
    layer1_outputs(11274) <= not b or a;
    layer1_outputs(11275) <= not b;
    layer1_outputs(11276) <= b and not a;
    layer1_outputs(11277) <= a and b;
    layer1_outputs(11278) <= a or b;
    layer1_outputs(11279) <= a and not b;
    layer1_outputs(11280) <= not a or b;
    layer1_outputs(11281) <= a or b;
    layer1_outputs(11282) <= not a or b;
    layer1_outputs(11283) <= a and b;
    layer1_outputs(11284) <= a or b;
    layer1_outputs(11285) <= b;
    layer1_outputs(11286) <= not b;
    layer1_outputs(11287) <= not (a xor b);
    layer1_outputs(11288) <= a;
    layer1_outputs(11289) <= not (a xor b);
    layer1_outputs(11290) <= b and not a;
    layer1_outputs(11291) <= a and b;
    layer1_outputs(11292) <= not (a and b);
    layer1_outputs(11293) <= a or b;
    layer1_outputs(11294) <= not a;
    layer1_outputs(11295) <= '0';
    layer1_outputs(11296) <= '0';
    layer1_outputs(11297) <= b;
    layer1_outputs(11298) <= not b or a;
    layer1_outputs(11299) <= a xor b;
    layer1_outputs(11300) <= not a;
    layer1_outputs(11301) <= not a;
    layer1_outputs(11302) <= not b;
    layer1_outputs(11303) <= b;
    layer1_outputs(11304) <= b;
    layer1_outputs(11305) <= a and not b;
    layer1_outputs(11306) <= not a;
    layer1_outputs(11307) <= not a or b;
    layer1_outputs(11308) <= b;
    layer1_outputs(11309) <= b and not a;
    layer1_outputs(11310) <= not (a xor b);
    layer1_outputs(11311) <= b and not a;
    layer1_outputs(11312) <= not b or a;
    layer1_outputs(11313) <= a and not b;
    layer1_outputs(11314) <= a;
    layer1_outputs(11315) <= a and b;
    layer1_outputs(11316) <= a or b;
    layer1_outputs(11317) <= a and not b;
    layer1_outputs(11318) <= a;
    layer1_outputs(11319) <= a and not b;
    layer1_outputs(11320) <= a xor b;
    layer1_outputs(11321) <= b and not a;
    layer1_outputs(11322) <= a;
    layer1_outputs(11323) <= a;
    layer1_outputs(11324) <= a and b;
    layer1_outputs(11325) <= a and b;
    layer1_outputs(11326) <= not a;
    layer1_outputs(11327) <= not (a xor b);
    layer1_outputs(11328) <= a;
    layer1_outputs(11329) <= a and not b;
    layer1_outputs(11330) <= not a or b;
    layer1_outputs(11331) <= '1';
    layer1_outputs(11332) <= not a or b;
    layer1_outputs(11333) <= a;
    layer1_outputs(11334) <= a and b;
    layer1_outputs(11335) <= not a;
    layer1_outputs(11336) <= not a or b;
    layer1_outputs(11337) <= '1';
    layer1_outputs(11338) <= not (a xor b);
    layer1_outputs(11339) <= not (a or b);
    layer1_outputs(11340) <= b;
    layer1_outputs(11341) <= not b or a;
    layer1_outputs(11342) <= not a or b;
    layer1_outputs(11343) <= a and b;
    layer1_outputs(11344) <= a and not b;
    layer1_outputs(11345) <= not (a and b);
    layer1_outputs(11346) <= not (a xor b);
    layer1_outputs(11347) <= '0';
    layer1_outputs(11348) <= not (a and b);
    layer1_outputs(11349) <= b and not a;
    layer1_outputs(11350) <= b and not a;
    layer1_outputs(11351) <= a xor b;
    layer1_outputs(11352) <= not a;
    layer1_outputs(11353) <= a or b;
    layer1_outputs(11354) <= not (a xor b);
    layer1_outputs(11355) <= not (a and b);
    layer1_outputs(11356) <= b and not a;
    layer1_outputs(11357) <= '0';
    layer1_outputs(11358) <= a or b;
    layer1_outputs(11359) <= not (a and b);
    layer1_outputs(11360) <= a and b;
    layer1_outputs(11361) <= not (a or b);
    layer1_outputs(11362) <= not b or a;
    layer1_outputs(11363) <= a;
    layer1_outputs(11364) <= not (a xor b);
    layer1_outputs(11365) <= '0';
    layer1_outputs(11366) <= a and b;
    layer1_outputs(11367) <= not a;
    layer1_outputs(11368) <= not (a or b);
    layer1_outputs(11369) <= not a or b;
    layer1_outputs(11370) <= not (a and b);
    layer1_outputs(11371) <= '0';
    layer1_outputs(11372) <= a and b;
    layer1_outputs(11373) <= not (a and b);
    layer1_outputs(11374) <= not a or b;
    layer1_outputs(11375) <= a and not b;
    layer1_outputs(11376) <= '1';
    layer1_outputs(11377) <= '0';
    layer1_outputs(11378) <= not a;
    layer1_outputs(11379) <= a and b;
    layer1_outputs(11380) <= not b or a;
    layer1_outputs(11381) <= not b or a;
    layer1_outputs(11382) <= not a or b;
    layer1_outputs(11383) <= a and not b;
    layer1_outputs(11384) <= '1';
    layer1_outputs(11385) <= not (a and b);
    layer1_outputs(11386) <= not (a xor b);
    layer1_outputs(11387) <= b;
    layer1_outputs(11388) <= a and b;
    layer1_outputs(11389) <= not a or b;
    layer1_outputs(11390) <= not a;
    layer1_outputs(11391) <= '1';
    layer1_outputs(11392) <= a xor b;
    layer1_outputs(11393) <= not (a xor b);
    layer1_outputs(11394) <= not a or b;
    layer1_outputs(11395) <= not b or a;
    layer1_outputs(11396) <= not (a xor b);
    layer1_outputs(11397) <= '1';
    layer1_outputs(11398) <= not a;
    layer1_outputs(11399) <= a and b;
    layer1_outputs(11400) <= a xor b;
    layer1_outputs(11401) <= not b or a;
    layer1_outputs(11402) <= not (a or b);
    layer1_outputs(11403) <= b;
    layer1_outputs(11404) <= not a or b;
    layer1_outputs(11405) <= a and not b;
    layer1_outputs(11406) <= not b or a;
    layer1_outputs(11407) <= a and not b;
    layer1_outputs(11408) <= '1';
    layer1_outputs(11409) <= a xor b;
    layer1_outputs(11410) <= a and not b;
    layer1_outputs(11411) <= b and not a;
    layer1_outputs(11412) <= '1';
    layer1_outputs(11413) <= a or b;
    layer1_outputs(11414) <= not b or a;
    layer1_outputs(11415) <= a;
    layer1_outputs(11416) <= b and not a;
    layer1_outputs(11417) <= a and b;
    layer1_outputs(11418) <= a xor b;
    layer1_outputs(11419) <= not b;
    layer1_outputs(11420) <= a and b;
    layer1_outputs(11421) <= a and not b;
    layer1_outputs(11422) <= a and b;
    layer1_outputs(11423) <= not b;
    layer1_outputs(11424) <= not (a and b);
    layer1_outputs(11425) <= b;
    layer1_outputs(11426) <= '0';
    layer1_outputs(11427) <= a or b;
    layer1_outputs(11428) <= a and b;
    layer1_outputs(11429) <= a;
    layer1_outputs(11430) <= a and not b;
    layer1_outputs(11431) <= not a or b;
    layer1_outputs(11432) <= a;
    layer1_outputs(11433) <= not a;
    layer1_outputs(11434) <= a or b;
    layer1_outputs(11435) <= b and not a;
    layer1_outputs(11436) <= not b;
    layer1_outputs(11437) <= '0';
    layer1_outputs(11438) <= not a;
    layer1_outputs(11439) <= a;
    layer1_outputs(11440) <= not (a or b);
    layer1_outputs(11441) <= not b;
    layer1_outputs(11442) <= a and not b;
    layer1_outputs(11443) <= a and b;
    layer1_outputs(11444) <= not a or b;
    layer1_outputs(11445) <= not a;
    layer1_outputs(11446) <= a;
    layer1_outputs(11447) <= a and not b;
    layer1_outputs(11448) <= not (a xor b);
    layer1_outputs(11449) <= a or b;
    layer1_outputs(11450) <= a and not b;
    layer1_outputs(11451) <= a and b;
    layer1_outputs(11452) <= a;
    layer1_outputs(11453) <= a;
    layer1_outputs(11454) <= not (a xor b);
    layer1_outputs(11455) <= a;
    layer1_outputs(11456) <= '1';
    layer1_outputs(11457) <= a;
    layer1_outputs(11458) <= a xor b;
    layer1_outputs(11459) <= b;
    layer1_outputs(11460) <= '1';
    layer1_outputs(11461) <= b and not a;
    layer1_outputs(11462) <= not (a or b);
    layer1_outputs(11463) <= b;
    layer1_outputs(11464) <= '1';
    layer1_outputs(11465) <= not (a or b);
    layer1_outputs(11466) <= '1';
    layer1_outputs(11467) <= a and not b;
    layer1_outputs(11468) <= not b or a;
    layer1_outputs(11469) <= '0';
    layer1_outputs(11470) <= a and not b;
    layer1_outputs(11471) <= b;
    layer1_outputs(11472) <= not b or a;
    layer1_outputs(11473) <= a and not b;
    layer1_outputs(11474) <= a and not b;
    layer1_outputs(11475) <= a and b;
    layer1_outputs(11476) <= a xor b;
    layer1_outputs(11477) <= not a;
    layer1_outputs(11478) <= not a;
    layer1_outputs(11479) <= b;
    layer1_outputs(11480) <= '1';
    layer1_outputs(11481) <= not (a and b);
    layer1_outputs(11482) <= not (a xor b);
    layer1_outputs(11483) <= b;
    layer1_outputs(11484) <= not a or b;
    layer1_outputs(11485) <= b and not a;
    layer1_outputs(11486) <= not a or b;
    layer1_outputs(11487) <= not b;
    layer1_outputs(11488) <= a and not b;
    layer1_outputs(11489) <= not b;
    layer1_outputs(11490) <= a;
    layer1_outputs(11491) <= not b or a;
    layer1_outputs(11492) <= not (a and b);
    layer1_outputs(11493) <= a and not b;
    layer1_outputs(11494) <= a;
    layer1_outputs(11495) <= b;
    layer1_outputs(11496) <= not (a and b);
    layer1_outputs(11497) <= a and not b;
    layer1_outputs(11498) <= a xor b;
    layer1_outputs(11499) <= a xor b;
    layer1_outputs(11500) <= b;
    layer1_outputs(11501) <= not a;
    layer1_outputs(11502) <= not a;
    layer1_outputs(11503) <= not a;
    layer1_outputs(11504) <= not (a and b);
    layer1_outputs(11505) <= not (a or b);
    layer1_outputs(11506) <= a or b;
    layer1_outputs(11507) <= a;
    layer1_outputs(11508) <= not b;
    layer1_outputs(11509) <= not (a or b);
    layer1_outputs(11510) <= not (a or b);
    layer1_outputs(11511) <= not (a xor b);
    layer1_outputs(11512) <= b;
    layer1_outputs(11513) <= b;
    layer1_outputs(11514) <= b and not a;
    layer1_outputs(11515) <= a and b;
    layer1_outputs(11516) <= not a;
    layer1_outputs(11517) <= not b or a;
    layer1_outputs(11518) <= b;
    layer1_outputs(11519) <= a or b;
    layer1_outputs(11520) <= '0';
    layer1_outputs(11521) <= a or b;
    layer1_outputs(11522) <= a and not b;
    layer1_outputs(11523) <= b and not a;
    layer1_outputs(11524) <= not b;
    layer1_outputs(11525) <= a and not b;
    layer1_outputs(11526) <= a and b;
    layer1_outputs(11527) <= not (a and b);
    layer1_outputs(11528) <= not (a and b);
    layer1_outputs(11529) <= a or b;
    layer1_outputs(11530) <= not b;
    layer1_outputs(11531) <= not a;
    layer1_outputs(11532) <= not a;
    layer1_outputs(11533) <= '1';
    layer1_outputs(11534) <= not (a and b);
    layer1_outputs(11535) <= not b or a;
    layer1_outputs(11536) <= not (a and b);
    layer1_outputs(11537) <= b and not a;
    layer1_outputs(11538) <= '1';
    layer1_outputs(11539) <= '1';
    layer1_outputs(11540) <= a and b;
    layer1_outputs(11541) <= b;
    layer1_outputs(11542) <= not a;
    layer1_outputs(11543) <= not b;
    layer1_outputs(11544) <= a and not b;
    layer1_outputs(11545) <= '1';
    layer1_outputs(11546) <= b and not a;
    layer1_outputs(11547) <= a and not b;
    layer1_outputs(11548) <= not a;
    layer1_outputs(11549) <= not (a or b);
    layer1_outputs(11550) <= not a;
    layer1_outputs(11551) <= not b or a;
    layer1_outputs(11552) <= '0';
    layer1_outputs(11553) <= not b;
    layer1_outputs(11554) <= not (a and b);
    layer1_outputs(11555) <= b and not a;
    layer1_outputs(11556) <= a;
    layer1_outputs(11557) <= '1';
    layer1_outputs(11558) <= '1';
    layer1_outputs(11559) <= a xor b;
    layer1_outputs(11560) <= a and not b;
    layer1_outputs(11561) <= a and b;
    layer1_outputs(11562) <= not (a xor b);
    layer1_outputs(11563) <= a and not b;
    layer1_outputs(11564) <= b;
    layer1_outputs(11565) <= a or b;
    layer1_outputs(11566) <= not a;
    layer1_outputs(11567) <= '1';
    layer1_outputs(11568) <= not b;
    layer1_outputs(11569) <= b and not a;
    layer1_outputs(11570) <= not a or b;
    layer1_outputs(11571) <= b and not a;
    layer1_outputs(11572) <= '1';
    layer1_outputs(11573) <= not b;
    layer1_outputs(11574) <= not b or a;
    layer1_outputs(11575) <= b and not a;
    layer1_outputs(11576) <= not a or b;
    layer1_outputs(11577) <= not a or b;
    layer1_outputs(11578) <= not (a and b);
    layer1_outputs(11579) <= not a;
    layer1_outputs(11580) <= not a;
    layer1_outputs(11581) <= not a;
    layer1_outputs(11582) <= not (a or b);
    layer1_outputs(11583) <= '1';
    layer1_outputs(11584) <= a;
    layer1_outputs(11585) <= b;
    layer1_outputs(11586) <= not (a or b);
    layer1_outputs(11587) <= a and not b;
    layer1_outputs(11588) <= b;
    layer1_outputs(11589) <= b and not a;
    layer1_outputs(11590) <= a;
    layer1_outputs(11591) <= '1';
    layer1_outputs(11592) <= a;
    layer1_outputs(11593) <= not b;
    layer1_outputs(11594) <= not a or b;
    layer1_outputs(11595) <= not b;
    layer1_outputs(11596) <= not a or b;
    layer1_outputs(11597) <= a or b;
    layer1_outputs(11598) <= not a or b;
    layer1_outputs(11599) <= not (a and b);
    layer1_outputs(11600) <= b and not a;
    layer1_outputs(11601) <= not (a or b);
    layer1_outputs(11602) <= b and not a;
    layer1_outputs(11603) <= a and not b;
    layer1_outputs(11604) <= a or b;
    layer1_outputs(11605) <= not b;
    layer1_outputs(11606) <= not (a or b);
    layer1_outputs(11607) <= a xor b;
    layer1_outputs(11608) <= not b;
    layer1_outputs(11609) <= a or b;
    layer1_outputs(11610) <= b and not a;
    layer1_outputs(11611) <= not a or b;
    layer1_outputs(11612) <= not b;
    layer1_outputs(11613) <= not b;
    layer1_outputs(11614) <= a;
    layer1_outputs(11615) <= a or b;
    layer1_outputs(11616) <= a and not b;
    layer1_outputs(11617) <= not (a and b);
    layer1_outputs(11618) <= a;
    layer1_outputs(11619) <= not a or b;
    layer1_outputs(11620) <= not a;
    layer1_outputs(11621) <= not (a or b);
    layer1_outputs(11622) <= a;
    layer1_outputs(11623) <= not a or b;
    layer1_outputs(11624) <= not (a or b);
    layer1_outputs(11625) <= not (a and b);
    layer1_outputs(11626) <= not b or a;
    layer1_outputs(11627) <= a;
    layer1_outputs(11628) <= a or b;
    layer1_outputs(11629) <= not (a or b);
    layer1_outputs(11630) <= not (a xor b);
    layer1_outputs(11631) <= not a or b;
    layer1_outputs(11632) <= '0';
    layer1_outputs(11633) <= a or b;
    layer1_outputs(11634) <= not b;
    layer1_outputs(11635) <= '1';
    layer1_outputs(11636) <= a;
    layer1_outputs(11637) <= a;
    layer1_outputs(11638) <= not (a and b);
    layer1_outputs(11639) <= not b or a;
    layer1_outputs(11640) <= b;
    layer1_outputs(11641) <= not (a xor b);
    layer1_outputs(11642) <= b;
    layer1_outputs(11643) <= b and not a;
    layer1_outputs(11644) <= not (a or b);
    layer1_outputs(11645) <= a;
    layer1_outputs(11646) <= not a or b;
    layer1_outputs(11647) <= not b or a;
    layer1_outputs(11648) <= not (a or b);
    layer1_outputs(11649) <= a and b;
    layer1_outputs(11650) <= not a;
    layer1_outputs(11651) <= not (a and b);
    layer1_outputs(11652) <= a xor b;
    layer1_outputs(11653) <= '0';
    layer1_outputs(11654) <= b;
    layer1_outputs(11655) <= '1';
    layer1_outputs(11656) <= not (a or b);
    layer1_outputs(11657) <= a xor b;
    layer1_outputs(11658) <= not b;
    layer1_outputs(11659) <= not b;
    layer1_outputs(11660) <= '0';
    layer1_outputs(11661) <= not (a or b);
    layer1_outputs(11662) <= a or b;
    layer1_outputs(11663) <= '0';
    layer1_outputs(11664) <= not a;
    layer1_outputs(11665) <= a and b;
    layer1_outputs(11666) <= a or b;
    layer1_outputs(11667) <= not a or b;
    layer1_outputs(11668) <= b and not a;
    layer1_outputs(11669) <= not a;
    layer1_outputs(11670) <= b and not a;
    layer1_outputs(11671) <= '0';
    layer1_outputs(11672) <= a;
    layer1_outputs(11673) <= '0';
    layer1_outputs(11674) <= not a;
    layer1_outputs(11675) <= b;
    layer1_outputs(11676) <= not b or a;
    layer1_outputs(11677) <= not (a and b);
    layer1_outputs(11678) <= not b or a;
    layer1_outputs(11679) <= not b or a;
    layer1_outputs(11680) <= not b;
    layer1_outputs(11681) <= not (a or b);
    layer1_outputs(11682) <= not (a or b);
    layer1_outputs(11683) <= not a or b;
    layer1_outputs(11684) <= a and b;
    layer1_outputs(11685) <= b and not a;
    layer1_outputs(11686) <= '0';
    layer1_outputs(11687) <= '0';
    layer1_outputs(11688) <= b;
    layer1_outputs(11689) <= not (a or b);
    layer1_outputs(11690) <= '1';
    layer1_outputs(11691) <= not (a xor b);
    layer1_outputs(11692) <= not a or b;
    layer1_outputs(11693) <= not b;
    layer1_outputs(11694) <= not a or b;
    layer1_outputs(11695) <= not (a and b);
    layer1_outputs(11696) <= not (a xor b);
    layer1_outputs(11697) <= '1';
    layer1_outputs(11698) <= a;
    layer1_outputs(11699) <= not a;
    layer1_outputs(11700) <= b and not a;
    layer1_outputs(11701) <= b and not a;
    layer1_outputs(11702) <= not (a or b);
    layer1_outputs(11703) <= b;
    layer1_outputs(11704) <= a and not b;
    layer1_outputs(11705) <= not a or b;
    layer1_outputs(11706) <= a xor b;
    layer1_outputs(11707) <= b and not a;
    layer1_outputs(11708) <= not b or a;
    layer1_outputs(11709) <= b;
    layer1_outputs(11710) <= not (a or b);
    layer1_outputs(11711) <= not (a or b);
    layer1_outputs(11712) <= a and not b;
    layer1_outputs(11713) <= not b;
    layer1_outputs(11714) <= b;
    layer1_outputs(11715) <= not b or a;
    layer1_outputs(11716) <= a and not b;
    layer1_outputs(11717) <= a and b;
    layer1_outputs(11718) <= a or b;
    layer1_outputs(11719) <= a or b;
    layer1_outputs(11720) <= not a or b;
    layer1_outputs(11721) <= '1';
    layer1_outputs(11722) <= a and b;
    layer1_outputs(11723) <= b and not a;
    layer1_outputs(11724) <= b;
    layer1_outputs(11725) <= a and b;
    layer1_outputs(11726) <= a or b;
    layer1_outputs(11727) <= not b;
    layer1_outputs(11728) <= b;
    layer1_outputs(11729) <= a;
    layer1_outputs(11730) <= not a;
    layer1_outputs(11731) <= not b or a;
    layer1_outputs(11732) <= '0';
    layer1_outputs(11733) <= not a;
    layer1_outputs(11734) <= not a or b;
    layer1_outputs(11735) <= '1';
    layer1_outputs(11736) <= not (a and b);
    layer1_outputs(11737) <= '0';
    layer1_outputs(11738) <= a;
    layer1_outputs(11739) <= not b or a;
    layer1_outputs(11740) <= b;
    layer1_outputs(11741) <= not b or a;
    layer1_outputs(11742) <= not b;
    layer1_outputs(11743) <= not b;
    layer1_outputs(11744) <= '0';
    layer1_outputs(11745) <= not a or b;
    layer1_outputs(11746) <= a and not b;
    layer1_outputs(11747) <= not (a or b);
    layer1_outputs(11748) <= a and b;
    layer1_outputs(11749) <= b;
    layer1_outputs(11750) <= not (a or b);
    layer1_outputs(11751) <= not (a or b);
    layer1_outputs(11752) <= a or b;
    layer1_outputs(11753) <= b;
    layer1_outputs(11754) <= not (a or b);
    layer1_outputs(11755) <= '0';
    layer1_outputs(11756) <= not b or a;
    layer1_outputs(11757) <= b;
    layer1_outputs(11758) <= not a;
    layer1_outputs(11759) <= '0';
    layer1_outputs(11760) <= a;
    layer1_outputs(11761) <= a and not b;
    layer1_outputs(11762) <= not b or a;
    layer1_outputs(11763) <= not b;
    layer1_outputs(11764) <= not b or a;
    layer1_outputs(11765) <= b;
    layer1_outputs(11766) <= not a;
    layer1_outputs(11767) <= '1';
    layer1_outputs(11768) <= '0';
    layer1_outputs(11769) <= not b;
    layer1_outputs(11770) <= '1';
    layer1_outputs(11771) <= not b;
    layer1_outputs(11772) <= not (a xor b);
    layer1_outputs(11773) <= a or b;
    layer1_outputs(11774) <= '0';
    layer1_outputs(11775) <= a or b;
    layer1_outputs(11776) <= a;
    layer1_outputs(11777) <= a and not b;
    layer1_outputs(11778) <= a and b;
    layer1_outputs(11779) <= a and b;
    layer1_outputs(11780) <= not a or b;
    layer1_outputs(11781) <= a xor b;
    layer1_outputs(11782) <= b;
    layer1_outputs(11783) <= not (a xor b);
    layer1_outputs(11784) <= not (a and b);
    layer1_outputs(11785) <= b and not a;
    layer1_outputs(11786) <= '1';
    layer1_outputs(11787) <= b and not a;
    layer1_outputs(11788) <= a or b;
    layer1_outputs(11789) <= b and not a;
    layer1_outputs(11790) <= a and b;
    layer1_outputs(11791) <= b and not a;
    layer1_outputs(11792) <= not (a and b);
    layer1_outputs(11793) <= not (a and b);
    layer1_outputs(11794) <= '0';
    layer1_outputs(11795) <= '1';
    layer1_outputs(11796) <= a and not b;
    layer1_outputs(11797) <= b;
    layer1_outputs(11798) <= not (a xor b);
    layer1_outputs(11799) <= not (a xor b);
    layer1_outputs(11800) <= a and b;
    layer1_outputs(11801) <= not a;
    layer1_outputs(11802) <= a and b;
    layer1_outputs(11803) <= b;
    layer1_outputs(11804) <= b;
    layer1_outputs(11805) <= a and not b;
    layer1_outputs(11806) <= b and not a;
    layer1_outputs(11807) <= b;
    layer1_outputs(11808) <= not (a xor b);
    layer1_outputs(11809) <= a and not b;
    layer1_outputs(11810) <= '0';
    layer1_outputs(11811) <= not a;
    layer1_outputs(11812) <= a or b;
    layer1_outputs(11813) <= '1';
    layer1_outputs(11814) <= b and not a;
    layer1_outputs(11815) <= b;
    layer1_outputs(11816) <= not (a xor b);
    layer1_outputs(11817) <= b and not a;
    layer1_outputs(11818) <= b and not a;
    layer1_outputs(11819) <= not b or a;
    layer1_outputs(11820) <= a and not b;
    layer1_outputs(11821) <= a and not b;
    layer1_outputs(11822) <= a;
    layer1_outputs(11823) <= b;
    layer1_outputs(11824) <= not a;
    layer1_outputs(11825) <= b;
    layer1_outputs(11826) <= a and b;
    layer1_outputs(11827) <= a;
    layer1_outputs(11828) <= '1';
    layer1_outputs(11829) <= not (a or b);
    layer1_outputs(11830) <= not (a and b);
    layer1_outputs(11831) <= not a;
    layer1_outputs(11832) <= b;
    layer1_outputs(11833) <= '0';
    layer1_outputs(11834) <= '1';
    layer1_outputs(11835) <= not (a or b);
    layer1_outputs(11836) <= not (a xor b);
    layer1_outputs(11837) <= a or b;
    layer1_outputs(11838) <= a;
    layer1_outputs(11839) <= not b or a;
    layer1_outputs(11840) <= a and b;
    layer1_outputs(11841) <= not a or b;
    layer1_outputs(11842) <= a xor b;
    layer1_outputs(11843) <= not a;
    layer1_outputs(11844) <= not (a and b);
    layer1_outputs(11845) <= not a;
    layer1_outputs(11846) <= '1';
    layer1_outputs(11847) <= b;
    layer1_outputs(11848) <= b and not a;
    layer1_outputs(11849) <= a and not b;
    layer1_outputs(11850) <= '0';
    layer1_outputs(11851) <= a;
    layer1_outputs(11852) <= not b;
    layer1_outputs(11853) <= not a;
    layer1_outputs(11854) <= a;
    layer1_outputs(11855) <= not a or b;
    layer1_outputs(11856) <= not b or a;
    layer1_outputs(11857) <= b and not a;
    layer1_outputs(11858) <= not b or a;
    layer1_outputs(11859) <= a or b;
    layer1_outputs(11860) <= not (a or b);
    layer1_outputs(11861) <= a;
    layer1_outputs(11862) <= not b or a;
    layer1_outputs(11863) <= not (a or b);
    layer1_outputs(11864) <= not a or b;
    layer1_outputs(11865) <= not (a and b);
    layer1_outputs(11866) <= not a;
    layer1_outputs(11867) <= a;
    layer1_outputs(11868) <= not a;
    layer1_outputs(11869) <= not b;
    layer1_outputs(11870) <= b;
    layer1_outputs(11871) <= a and not b;
    layer1_outputs(11872) <= not (a or b);
    layer1_outputs(11873) <= '0';
    layer1_outputs(11874) <= '1';
    layer1_outputs(11875) <= b and not a;
    layer1_outputs(11876) <= not b or a;
    layer1_outputs(11877) <= b;
    layer1_outputs(11878) <= b and not a;
    layer1_outputs(11879) <= not b;
    layer1_outputs(11880) <= '1';
    layer1_outputs(11881) <= not a;
    layer1_outputs(11882) <= not b;
    layer1_outputs(11883) <= not b or a;
    layer1_outputs(11884) <= b;
    layer1_outputs(11885) <= a xor b;
    layer1_outputs(11886) <= '1';
    layer1_outputs(11887) <= '1';
    layer1_outputs(11888) <= not b;
    layer1_outputs(11889) <= a xor b;
    layer1_outputs(11890) <= a;
    layer1_outputs(11891) <= a or b;
    layer1_outputs(11892) <= not (a xor b);
    layer1_outputs(11893) <= '1';
    layer1_outputs(11894) <= not b;
    layer1_outputs(11895) <= '0';
    layer1_outputs(11896) <= not b;
    layer1_outputs(11897) <= not b;
    layer1_outputs(11898) <= '1';
    layer1_outputs(11899) <= not a;
    layer1_outputs(11900) <= a and not b;
    layer1_outputs(11901) <= not a;
    layer1_outputs(11902) <= not a or b;
    layer1_outputs(11903) <= not a;
    layer1_outputs(11904) <= not (a or b);
    layer1_outputs(11905) <= not (a or b);
    layer1_outputs(11906) <= a;
    layer1_outputs(11907) <= a or b;
    layer1_outputs(11908) <= not b or a;
    layer1_outputs(11909) <= not b or a;
    layer1_outputs(11910) <= not (a or b);
    layer1_outputs(11911) <= not (a or b);
    layer1_outputs(11912) <= b;
    layer1_outputs(11913) <= not b;
    layer1_outputs(11914) <= not b;
    layer1_outputs(11915) <= b;
    layer1_outputs(11916) <= a or b;
    layer1_outputs(11917) <= not b;
    layer1_outputs(11918) <= not a;
    layer1_outputs(11919) <= b and not a;
    layer1_outputs(11920) <= not a;
    layer1_outputs(11921) <= a;
    layer1_outputs(11922) <= a and b;
    layer1_outputs(11923) <= not (a xor b);
    layer1_outputs(11924) <= a or b;
    layer1_outputs(11925) <= a and b;
    layer1_outputs(11926) <= not (a or b);
    layer1_outputs(11927) <= not a or b;
    layer1_outputs(11928) <= not b or a;
    layer1_outputs(11929) <= a;
    layer1_outputs(11930) <= not a;
    layer1_outputs(11931) <= not (a xor b);
    layer1_outputs(11932) <= b and not a;
    layer1_outputs(11933) <= not (a and b);
    layer1_outputs(11934) <= '1';
    layer1_outputs(11935) <= b;
    layer1_outputs(11936) <= a and b;
    layer1_outputs(11937) <= b;
    layer1_outputs(11938) <= a;
    layer1_outputs(11939) <= a and not b;
    layer1_outputs(11940) <= a;
    layer1_outputs(11941) <= a or b;
    layer1_outputs(11942) <= a and b;
    layer1_outputs(11943) <= b and not a;
    layer1_outputs(11944) <= not b or a;
    layer1_outputs(11945) <= b and not a;
    layer1_outputs(11946) <= b and not a;
    layer1_outputs(11947) <= not a;
    layer1_outputs(11948) <= not b;
    layer1_outputs(11949) <= a and not b;
    layer1_outputs(11950) <= not a;
    layer1_outputs(11951) <= a xor b;
    layer1_outputs(11952) <= b and not a;
    layer1_outputs(11953) <= '1';
    layer1_outputs(11954) <= not a or b;
    layer1_outputs(11955) <= a and not b;
    layer1_outputs(11956) <= not (a and b);
    layer1_outputs(11957) <= a and b;
    layer1_outputs(11958) <= b;
    layer1_outputs(11959) <= not b or a;
    layer1_outputs(11960) <= a and b;
    layer1_outputs(11961) <= not b or a;
    layer1_outputs(11962) <= a;
    layer1_outputs(11963) <= not (a xor b);
    layer1_outputs(11964) <= a and not b;
    layer1_outputs(11965) <= not (a and b);
    layer1_outputs(11966) <= a and b;
    layer1_outputs(11967) <= '1';
    layer1_outputs(11968) <= a or b;
    layer1_outputs(11969) <= a;
    layer1_outputs(11970) <= not a;
    layer1_outputs(11971) <= not a;
    layer1_outputs(11972) <= '1';
    layer1_outputs(11973) <= not b or a;
    layer1_outputs(11974) <= a xor b;
    layer1_outputs(11975) <= a;
    layer1_outputs(11976) <= b;
    layer1_outputs(11977) <= b;
    layer1_outputs(11978) <= a;
    layer1_outputs(11979) <= a;
    layer1_outputs(11980) <= not (a or b);
    layer1_outputs(11981) <= not a;
    layer1_outputs(11982) <= '1';
    layer1_outputs(11983) <= not b or a;
    layer1_outputs(11984) <= not a or b;
    layer1_outputs(11985) <= not a or b;
    layer1_outputs(11986) <= a or b;
    layer1_outputs(11987) <= '0';
    layer1_outputs(11988) <= b and not a;
    layer1_outputs(11989) <= b;
    layer1_outputs(11990) <= a;
    layer1_outputs(11991) <= '1';
    layer1_outputs(11992) <= '1';
    layer1_outputs(11993) <= not b;
    layer1_outputs(11994) <= not (a or b);
    layer1_outputs(11995) <= a xor b;
    layer1_outputs(11996) <= a;
    layer1_outputs(11997) <= not a or b;
    layer1_outputs(11998) <= not (a xor b);
    layer1_outputs(11999) <= a xor b;
    layer1_outputs(12000) <= '1';
    layer1_outputs(12001) <= a and not b;
    layer1_outputs(12002) <= not b or a;
    layer1_outputs(12003) <= not a;
    layer1_outputs(12004) <= not (a or b);
    layer1_outputs(12005) <= b;
    layer1_outputs(12006) <= not (a xor b);
    layer1_outputs(12007) <= not a or b;
    layer1_outputs(12008) <= not b;
    layer1_outputs(12009) <= not (a xor b);
    layer1_outputs(12010) <= '1';
    layer1_outputs(12011) <= a and b;
    layer1_outputs(12012) <= a or b;
    layer1_outputs(12013) <= b;
    layer1_outputs(12014) <= not (a and b);
    layer1_outputs(12015) <= b and not a;
    layer1_outputs(12016) <= '1';
    layer1_outputs(12017) <= a;
    layer1_outputs(12018) <= not a;
    layer1_outputs(12019) <= a and b;
    layer1_outputs(12020) <= not b;
    layer1_outputs(12021) <= not b or a;
    layer1_outputs(12022) <= b and not a;
    layer1_outputs(12023) <= not (a and b);
    layer1_outputs(12024) <= '1';
    layer1_outputs(12025) <= not (a or b);
    layer1_outputs(12026) <= a xor b;
    layer1_outputs(12027) <= b;
    layer1_outputs(12028) <= b;
    layer1_outputs(12029) <= '0';
    layer1_outputs(12030) <= not (a or b);
    layer1_outputs(12031) <= '1';
    layer1_outputs(12032) <= a or b;
    layer1_outputs(12033) <= not (a xor b);
    layer1_outputs(12034) <= a and b;
    layer1_outputs(12035) <= a;
    layer1_outputs(12036) <= not b or a;
    layer1_outputs(12037) <= '1';
    layer1_outputs(12038) <= a xor b;
    layer1_outputs(12039) <= '1';
    layer1_outputs(12040) <= '1';
    layer1_outputs(12041) <= not a or b;
    layer1_outputs(12042) <= a and b;
    layer1_outputs(12043) <= b;
    layer1_outputs(12044) <= b;
    layer1_outputs(12045) <= a and b;
    layer1_outputs(12046) <= b;
    layer1_outputs(12047) <= not b or a;
    layer1_outputs(12048) <= '0';
    layer1_outputs(12049) <= b;
    layer1_outputs(12050) <= a and b;
    layer1_outputs(12051) <= a or b;
    layer1_outputs(12052) <= not b or a;
    layer1_outputs(12053) <= not b;
    layer1_outputs(12054) <= '1';
    layer1_outputs(12055) <= a;
    layer1_outputs(12056) <= a and not b;
    layer1_outputs(12057) <= b;
    layer1_outputs(12058) <= a and not b;
    layer1_outputs(12059) <= b and not a;
    layer1_outputs(12060) <= not (a xor b);
    layer1_outputs(12061) <= not (a and b);
    layer1_outputs(12062) <= '1';
    layer1_outputs(12063) <= not a;
    layer1_outputs(12064) <= b and not a;
    layer1_outputs(12065) <= not (a xor b);
    layer1_outputs(12066) <= not a;
    layer1_outputs(12067) <= not (a and b);
    layer1_outputs(12068) <= a or b;
    layer1_outputs(12069) <= not a;
    layer1_outputs(12070) <= not (a and b);
    layer1_outputs(12071) <= a and not b;
    layer1_outputs(12072) <= '0';
    layer1_outputs(12073) <= not b or a;
    layer1_outputs(12074) <= a;
    layer1_outputs(12075) <= not a or b;
    layer1_outputs(12076) <= not (a and b);
    layer1_outputs(12077) <= not b;
    layer1_outputs(12078) <= not (a or b);
    layer1_outputs(12079) <= '0';
    layer1_outputs(12080) <= b and not a;
    layer1_outputs(12081) <= a xor b;
    layer1_outputs(12082) <= b;
    layer1_outputs(12083) <= a and not b;
    layer1_outputs(12084) <= not b;
    layer1_outputs(12085) <= a or b;
    layer1_outputs(12086) <= '1';
    layer1_outputs(12087) <= not b;
    layer1_outputs(12088) <= not a;
    layer1_outputs(12089) <= not b;
    layer1_outputs(12090) <= a;
    layer1_outputs(12091) <= not b;
    layer1_outputs(12092) <= not a or b;
    layer1_outputs(12093) <= not b;
    layer1_outputs(12094) <= a or b;
    layer1_outputs(12095) <= a;
    layer1_outputs(12096) <= not b;
    layer1_outputs(12097) <= not (a or b);
    layer1_outputs(12098) <= not (a or b);
    layer1_outputs(12099) <= not a;
    layer1_outputs(12100) <= a and not b;
    layer1_outputs(12101) <= a and not b;
    layer1_outputs(12102) <= a xor b;
    layer1_outputs(12103) <= a and not b;
    layer1_outputs(12104) <= a;
    layer1_outputs(12105) <= not a;
    layer1_outputs(12106) <= not (a and b);
    layer1_outputs(12107) <= a and not b;
    layer1_outputs(12108) <= a;
    layer1_outputs(12109) <= a and not b;
    layer1_outputs(12110) <= not a or b;
    layer1_outputs(12111) <= a and not b;
    layer1_outputs(12112) <= '0';
    layer1_outputs(12113) <= a and b;
    layer1_outputs(12114) <= a or b;
    layer1_outputs(12115) <= b and not a;
    layer1_outputs(12116) <= '0';
    layer1_outputs(12117) <= b;
    layer1_outputs(12118) <= not b;
    layer1_outputs(12119) <= a or b;
    layer1_outputs(12120) <= not (a or b);
    layer1_outputs(12121) <= a and b;
    layer1_outputs(12122) <= '1';
    layer1_outputs(12123) <= not a;
    layer1_outputs(12124) <= a;
    layer1_outputs(12125) <= a;
    layer1_outputs(12126) <= a;
    layer1_outputs(12127) <= not (a and b);
    layer1_outputs(12128) <= not a;
    layer1_outputs(12129) <= a or b;
    layer1_outputs(12130) <= not a;
    layer1_outputs(12131) <= not b;
    layer1_outputs(12132) <= '1';
    layer1_outputs(12133) <= not a or b;
    layer1_outputs(12134) <= not b;
    layer1_outputs(12135) <= not (a or b);
    layer1_outputs(12136) <= a;
    layer1_outputs(12137) <= not a;
    layer1_outputs(12138) <= a or b;
    layer1_outputs(12139) <= b;
    layer1_outputs(12140) <= a or b;
    layer1_outputs(12141) <= b;
    layer1_outputs(12142) <= not a;
    layer1_outputs(12143) <= a xor b;
    layer1_outputs(12144) <= a;
    layer1_outputs(12145) <= not b;
    layer1_outputs(12146) <= not (a xor b);
    layer1_outputs(12147) <= a;
    layer1_outputs(12148) <= not b or a;
    layer1_outputs(12149) <= b;
    layer1_outputs(12150) <= not b or a;
    layer1_outputs(12151) <= '1';
    layer1_outputs(12152) <= not (a and b);
    layer1_outputs(12153) <= b and not a;
    layer1_outputs(12154) <= a and not b;
    layer1_outputs(12155) <= not a or b;
    layer1_outputs(12156) <= not (a or b);
    layer1_outputs(12157) <= not (a xor b);
    layer1_outputs(12158) <= b;
    layer1_outputs(12159) <= '1';
    layer1_outputs(12160) <= '1';
    layer1_outputs(12161) <= b and not a;
    layer1_outputs(12162) <= a and not b;
    layer1_outputs(12163) <= '1';
    layer1_outputs(12164) <= not a;
    layer1_outputs(12165) <= not b or a;
    layer1_outputs(12166) <= not (a or b);
    layer1_outputs(12167) <= '1';
    layer1_outputs(12168) <= not a;
    layer1_outputs(12169) <= a and not b;
    layer1_outputs(12170) <= a;
    layer1_outputs(12171) <= b;
    layer1_outputs(12172) <= b;
    layer1_outputs(12173) <= '0';
    layer1_outputs(12174) <= '0';
    layer1_outputs(12175) <= '1';
    layer1_outputs(12176) <= not a or b;
    layer1_outputs(12177) <= not (a or b);
    layer1_outputs(12178) <= a;
    layer1_outputs(12179) <= a and not b;
    layer1_outputs(12180) <= a and not b;
    layer1_outputs(12181) <= not (a xor b);
    layer1_outputs(12182) <= a;
    layer1_outputs(12183) <= not b;
    layer1_outputs(12184) <= a or b;
    layer1_outputs(12185) <= a and b;
    layer1_outputs(12186) <= b;
    layer1_outputs(12187) <= a xor b;
    layer1_outputs(12188) <= not b;
    layer1_outputs(12189) <= a;
    layer1_outputs(12190) <= a or b;
    layer1_outputs(12191) <= b;
    layer1_outputs(12192) <= a or b;
    layer1_outputs(12193) <= a or b;
    layer1_outputs(12194) <= a and not b;
    layer1_outputs(12195) <= b;
    layer1_outputs(12196) <= '0';
    layer1_outputs(12197) <= b and not a;
    layer1_outputs(12198) <= a xor b;
    layer1_outputs(12199) <= a and b;
    layer1_outputs(12200) <= '0';
    layer1_outputs(12201) <= '0';
    layer1_outputs(12202) <= b and not a;
    layer1_outputs(12203) <= not (a xor b);
    layer1_outputs(12204) <= a and b;
    layer1_outputs(12205) <= a;
    layer1_outputs(12206) <= a xor b;
    layer1_outputs(12207) <= a;
    layer1_outputs(12208) <= not a or b;
    layer1_outputs(12209) <= '1';
    layer1_outputs(12210) <= a and not b;
    layer1_outputs(12211) <= b and not a;
    layer1_outputs(12212) <= not b;
    layer1_outputs(12213) <= b and not a;
    layer1_outputs(12214) <= not (a or b);
    layer1_outputs(12215) <= not b;
    layer1_outputs(12216) <= '1';
    layer1_outputs(12217) <= a and b;
    layer1_outputs(12218) <= a and not b;
    layer1_outputs(12219) <= not (a or b);
    layer1_outputs(12220) <= not (a and b);
    layer1_outputs(12221) <= '0';
    layer1_outputs(12222) <= '0';
    layer1_outputs(12223) <= a;
    layer1_outputs(12224) <= not a or b;
    layer1_outputs(12225) <= not b;
    layer1_outputs(12226) <= not (a or b);
    layer1_outputs(12227) <= not (a and b);
    layer1_outputs(12228) <= not b;
    layer1_outputs(12229) <= '1';
    layer1_outputs(12230) <= b and not a;
    layer1_outputs(12231) <= b;
    layer1_outputs(12232) <= b;
    layer1_outputs(12233) <= a and not b;
    layer1_outputs(12234) <= not (a and b);
    layer1_outputs(12235) <= a or b;
    layer1_outputs(12236) <= b;
    layer1_outputs(12237) <= b;
    layer1_outputs(12238) <= not a;
    layer1_outputs(12239) <= a or b;
    layer1_outputs(12240) <= not (a xor b);
    layer1_outputs(12241) <= not (a xor b);
    layer1_outputs(12242) <= a and b;
    layer1_outputs(12243) <= not (a and b);
    layer1_outputs(12244) <= a xor b;
    layer1_outputs(12245) <= a xor b;
    layer1_outputs(12246) <= '1';
    layer1_outputs(12247) <= not a;
    layer1_outputs(12248) <= a;
    layer1_outputs(12249) <= not (a or b);
    layer1_outputs(12250) <= b and not a;
    layer1_outputs(12251) <= a;
    layer1_outputs(12252) <= a;
    layer1_outputs(12253) <= not a;
    layer1_outputs(12254) <= a;
    layer1_outputs(12255) <= not (a xor b);
    layer1_outputs(12256) <= b and not a;
    layer1_outputs(12257) <= not a;
    layer1_outputs(12258) <= b and not a;
    layer1_outputs(12259) <= not b;
    layer1_outputs(12260) <= a or b;
    layer1_outputs(12261) <= a;
    layer1_outputs(12262) <= not (a and b);
    layer1_outputs(12263) <= a;
    layer1_outputs(12264) <= a and not b;
    layer1_outputs(12265) <= a xor b;
    layer1_outputs(12266) <= a and b;
    layer1_outputs(12267) <= '1';
    layer1_outputs(12268) <= not a;
    layer1_outputs(12269) <= not b;
    layer1_outputs(12270) <= a and not b;
    layer1_outputs(12271) <= not a or b;
    layer1_outputs(12272) <= b;
    layer1_outputs(12273) <= not b or a;
    layer1_outputs(12274) <= not b;
    layer1_outputs(12275) <= b;
    layer1_outputs(12276) <= not (a and b);
    layer1_outputs(12277) <= a;
    layer1_outputs(12278) <= not (a and b);
    layer1_outputs(12279) <= not (a or b);
    layer1_outputs(12280) <= a;
    layer1_outputs(12281) <= not (a or b);
    layer1_outputs(12282) <= not b;
    layer1_outputs(12283) <= '0';
    layer1_outputs(12284) <= not b;
    layer1_outputs(12285) <= a and b;
    layer1_outputs(12286) <= not a;
    layer1_outputs(12287) <= a xor b;
    layer1_outputs(12288) <= not (a and b);
    layer1_outputs(12289) <= a and b;
    layer1_outputs(12290) <= a xor b;
    layer1_outputs(12291) <= a xor b;
    layer1_outputs(12292) <= not b;
    layer1_outputs(12293) <= not b;
    layer1_outputs(12294) <= not (a or b);
    layer1_outputs(12295) <= not (a and b);
    layer1_outputs(12296) <= b;
    layer1_outputs(12297) <= not a or b;
    layer1_outputs(12298) <= b;
    layer1_outputs(12299) <= a and b;
    layer1_outputs(12300) <= not a or b;
    layer1_outputs(12301) <= a or b;
    layer1_outputs(12302) <= a xor b;
    layer1_outputs(12303) <= not b or a;
    layer1_outputs(12304) <= not b or a;
    layer1_outputs(12305) <= a and b;
    layer1_outputs(12306) <= a;
    layer1_outputs(12307) <= not b or a;
    layer1_outputs(12308) <= '1';
    layer1_outputs(12309) <= b;
    layer1_outputs(12310) <= a;
    layer1_outputs(12311) <= '0';
    layer1_outputs(12312) <= '0';
    layer1_outputs(12313) <= a;
    layer1_outputs(12314) <= '1';
    layer1_outputs(12315) <= a or b;
    layer1_outputs(12316) <= a or b;
    layer1_outputs(12317) <= a and b;
    layer1_outputs(12318) <= a or b;
    layer1_outputs(12319) <= b;
    layer1_outputs(12320) <= not b;
    layer1_outputs(12321) <= a or b;
    layer1_outputs(12322) <= not b;
    layer1_outputs(12323) <= a;
    layer1_outputs(12324) <= b and not a;
    layer1_outputs(12325) <= a and b;
    layer1_outputs(12326) <= not a;
    layer1_outputs(12327) <= b and not a;
    layer1_outputs(12328) <= b;
    layer1_outputs(12329) <= not (a and b);
    layer1_outputs(12330) <= b;
    layer1_outputs(12331) <= not b or a;
    layer1_outputs(12332) <= a or b;
    layer1_outputs(12333) <= not a;
    layer1_outputs(12334) <= not a;
    layer1_outputs(12335) <= a or b;
    layer1_outputs(12336) <= '0';
    layer1_outputs(12337) <= '0';
    layer1_outputs(12338) <= not b or a;
    layer1_outputs(12339) <= b;
    layer1_outputs(12340) <= not a or b;
    layer1_outputs(12341) <= a and b;
    layer1_outputs(12342) <= a and not b;
    layer1_outputs(12343) <= b;
    layer1_outputs(12344) <= not a;
    layer1_outputs(12345) <= not a;
    layer1_outputs(12346) <= a or b;
    layer1_outputs(12347) <= not a;
    layer1_outputs(12348) <= not (a and b);
    layer1_outputs(12349) <= b;
    layer1_outputs(12350) <= not (a and b);
    layer1_outputs(12351) <= '0';
    layer1_outputs(12352) <= a or b;
    layer1_outputs(12353) <= not b or a;
    layer1_outputs(12354) <= a and b;
    layer1_outputs(12355) <= not a or b;
    layer1_outputs(12356) <= b;
    layer1_outputs(12357) <= not a;
    layer1_outputs(12358) <= b;
    layer1_outputs(12359) <= b;
    layer1_outputs(12360) <= not a or b;
    layer1_outputs(12361) <= b;
    layer1_outputs(12362) <= a xor b;
    layer1_outputs(12363) <= a and b;
    layer1_outputs(12364) <= not b;
    layer1_outputs(12365) <= a and not b;
    layer1_outputs(12366) <= '1';
    layer1_outputs(12367) <= not b;
    layer1_outputs(12368) <= a and not b;
    layer1_outputs(12369) <= not a or b;
    layer1_outputs(12370) <= not b;
    layer1_outputs(12371) <= not (a and b);
    layer1_outputs(12372) <= not (a or b);
    layer1_outputs(12373) <= a xor b;
    layer1_outputs(12374) <= a and b;
    layer1_outputs(12375) <= a;
    layer1_outputs(12376) <= a and b;
    layer1_outputs(12377) <= a and not b;
    layer1_outputs(12378) <= not a;
    layer1_outputs(12379) <= '0';
    layer1_outputs(12380) <= a xor b;
    layer1_outputs(12381) <= a xor b;
    layer1_outputs(12382) <= not b or a;
    layer1_outputs(12383) <= '0';
    layer1_outputs(12384) <= '0';
    layer1_outputs(12385) <= a or b;
    layer1_outputs(12386) <= a and not b;
    layer1_outputs(12387) <= a;
    layer1_outputs(12388) <= a and not b;
    layer1_outputs(12389) <= not (a or b);
    layer1_outputs(12390) <= a;
    layer1_outputs(12391) <= not (a and b);
    layer1_outputs(12392) <= not a;
    layer1_outputs(12393) <= b and not a;
    layer1_outputs(12394) <= not b or a;
    layer1_outputs(12395) <= a;
    layer1_outputs(12396) <= b and not a;
    layer1_outputs(12397) <= a xor b;
    layer1_outputs(12398) <= not b;
    layer1_outputs(12399) <= not a or b;
    layer1_outputs(12400) <= not (a and b);
    layer1_outputs(12401) <= not b;
    layer1_outputs(12402) <= not (a or b);
    layer1_outputs(12403) <= '1';
    layer1_outputs(12404) <= a or b;
    layer1_outputs(12405) <= b;
    layer1_outputs(12406) <= a xor b;
    layer1_outputs(12407) <= not a;
    layer1_outputs(12408) <= not a;
    layer1_outputs(12409) <= not a or b;
    layer1_outputs(12410) <= not (a or b);
    layer1_outputs(12411) <= not a;
    layer1_outputs(12412) <= b and not a;
    layer1_outputs(12413) <= a or b;
    layer1_outputs(12414) <= a;
    layer1_outputs(12415) <= b;
    layer1_outputs(12416) <= '1';
    layer1_outputs(12417) <= not a or b;
    layer1_outputs(12418) <= not b;
    layer1_outputs(12419) <= '0';
    layer1_outputs(12420) <= '0';
    layer1_outputs(12421) <= a and not b;
    layer1_outputs(12422) <= a;
    layer1_outputs(12423) <= a;
    layer1_outputs(12424) <= a xor b;
    layer1_outputs(12425) <= not b;
    layer1_outputs(12426) <= not b;
    layer1_outputs(12427) <= b and not a;
    layer1_outputs(12428) <= '1';
    layer1_outputs(12429) <= '1';
    layer1_outputs(12430) <= not a or b;
    layer1_outputs(12431) <= b and not a;
    layer1_outputs(12432) <= a and not b;
    layer1_outputs(12433) <= a and b;
    layer1_outputs(12434) <= a and b;
    layer1_outputs(12435) <= not (a xor b);
    layer1_outputs(12436) <= b;
    layer1_outputs(12437) <= a or b;
    layer1_outputs(12438) <= not a or b;
    layer1_outputs(12439) <= a and b;
    layer1_outputs(12440) <= not b or a;
    layer1_outputs(12441) <= not (a and b);
    layer1_outputs(12442) <= not a;
    layer1_outputs(12443) <= b;
    layer1_outputs(12444) <= a and b;
    layer1_outputs(12445) <= a and b;
    layer1_outputs(12446) <= '1';
    layer1_outputs(12447) <= not b or a;
    layer1_outputs(12448) <= not (a or b);
    layer1_outputs(12449) <= a;
    layer1_outputs(12450) <= b and not a;
    layer1_outputs(12451) <= not b;
    layer1_outputs(12452) <= b and not a;
    layer1_outputs(12453) <= a and not b;
    layer1_outputs(12454) <= not (a and b);
    layer1_outputs(12455) <= b;
    layer1_outputs(12456) <= a xor b;
    layer1_outputs(12457) <= b and not a;
    layer1_outputs(12458) <= not a;
    layer1_outputs(12459) <= a or b;
    layer1_outputs(12460) <= not (a and b);
    layer1_outputs(12461) <= b;
    layer1_outputs(12462) <= a and b;
    layer1_outputs(12463) <= a and not b;
    layer1_outputs(12464) <= b;
    layer1_outputs(12465) <= not b or a;
    layer1_outputs(12466) <= not a or b;
    layer1_outputs(12467) <= not b or a;
    layer1_outputs(12468) <= not (a or b);
    layer1_outputs(12469) <= a;
    layer1_outputs(12470) <= not (a and b);
    layer1_outputs(12471) <= not b;
    layer1_outputs(12472) <= a and b;
    layer1_outputs(12473) <= not (a and b);
    layer1_outputs(12474) <= a and not b;
    layer1_outputs(12475) <= not a;
    layer1_outputs(12476) <= a;
    layer1_outputs(12477) <= not b;
    layer1_outputs(12478) <= a and not b;
    layer1_outputs(12479) <= not (a or b);
    layer1_outputs(12480) <= a or b;
    layer1_outputs(12481) <= a and b;
    layer1_outputs(12482) <= not a or b;
    layer1_outputs(12483) <= b and not a;
    layer1_outputs(12484) <= a;
    layer1_outputs(12485) <= not a or b;
    layer1_outputs(12486) <= a;
    layer1_outputs(12487) <= not b;
    layer1_outputs(12488) <= not a or b;
    layer1_outputs(12489) <= not (a and b);
    layer1_outputs(12490) <= a;
    layer1_outputs(12491) <= not b;
    layer1_outputs(12492) <= not (a and b);
    layer1_outputs(12493) <= not a;
    layer1_outputs(12494) <= a;
    layer1_outputs(12495) <= not b;
    layer1_outputs(12496) <= '1';
    layer1_outputs(12497) <= not (a xor b);
    layer1_outputs(12498) <= a or b;
    layer1_outputs(12499) <= b;
    layer1_outputs(12500) <= a;
    layer1_outputs(12501) <= b and not a;
    layer1_outputs(12502) <= a or b;
    layer1_outputs(12503) <= a and b;
    layer1_outputs(12504) <= not (a xor b);
    layer1_outputs(12505) <= not b or a;
    layer1_outputs(12506) <= '0';
    layer1_outputs(12507) <= a and b;
    layer1_outputs(12508) <= not b or a;
    layer1_outputs(12509) <= '1';
    layer1_outputs(12510) <= a and b;
    layer1_outputs(12511) <= '0';
    layer1_outputs(12512) <= a and not b;
    layer1_outputs(12513) <= not (a or b);
    layer1_outputs(12514) <= not (a or b);
    layer1_outputs(12515) <= a and b;
    layer1_outputs(12516) <= a or b;
    layer1_outputs(12517) <= b;
    layer1_outputs(12518) <= not b;
    layer1_outputs(12519) <= not (a xor b);
    layer1_outputs(12520) <= a or b;
    layer1_outputs(12521) <= not (a xor b);
    layer1_outputs(12522) <= a and not b;
    layer1_outputs(12523) <= not b;
    layer1_outputs(12524) <= not (a or b);
    layer1_outputs(12525) <= a;
    layer1_outputs(12526) <= a;
    layer1_outputs(12527) <= not a or b;
    layer1_outputs(12528) <= a;
    layer1_outputs(12529) <= not a or b;
    layer1_outputs(12530) <= a xor b;
    layer1_outputs(12531) <= b and not a;
    layer1_outputs(12532) <= '1';
    layer1_outputs(12533) <= '0';
    layer1_outputs(12534) <= b and not a;
    layer1_outputs(12535) <= a;
    layer1_outputs(12536) <= a xor b;
    layer1_outputs(12537) <= a;
    layer1_outputs(12538) <= b;
    layer1_outputs(12539) <= b;
    layer1_outputs(12540) <= not a;
    layer1_outputs(12541) <= not a;
    layer1_outputs(12542) <= a;
    layer1_outputs(12543) <= not a or b;
    layer1_outputs(12544) <= not (a and b);
    layer1_outputs(12545) <= not a or b;
    layer1_outputs(12546) <= not b or a;
    layer1_outputs(12547) <= not (a or b);
    layer1_outputs(12548) <= a;
    layer1_outputs(12549) <= not b or a;
    layer1_outputs(12550) <= not b;
    layer1_outputs(12551) <= a;
    layer1_outputs(12552) <= not b;
    layer1_outputs(12553) <= '1';
    layer1_outputs(12554) <= not a;
    layer1_outputs(12555) <= a and not b;
    layer1_outputs(12556) <= a or b;
    layer1_outputs(12557) <= a xor b;
    layer1_outputs(12558) <= '0';
    layer1_outputs(12559) <= not a or b;
    layer1_outputs(12560) <= '1';
    layer1_outputs(12561) <= a and not b;
    layer1_outputs(12562) <= not (a and b);
    layer1_outputs(12563) <= not a or b;
    layer1_outputs(12564) <= a;
    layer1_outputs(12565) <= '1';
    layer1_outputs(12566) <= '0';
    layer1_outputs(12567) <= a xor b;
    layer1_outputs(12568) <= not (a and b);
    layer1_outputs(12569) <= not a or b;
    layer1_outputs(12570) <= not (a or b);
    layer1_outputs(12571) <= not b or a;
    layer1_outputs(12572) <= b and not a;
    layer1_outputs(12573) <= a or b;
    layer1_outputs(12574) <= not (a or b);
    layer1_outputs(12575) <= a and b;
    layer1_outputs(12576) <= a xor b;
    layer1_outputs(12577) <= a and b;
    layer1_outputs(12578) <= not a or b;
    layer1_outputs(12579) <= a and b;
    layer1_outputs(12580) <= '1';
    layer1_outputs(12581) <= a and not b;
    layer1_outputs(12582) <= '0';
    layer1_outputs(12583) <= b;
    layer1_outputs(12584) <= not (a and b);
    layer1_outputs(12585) <= not a or b;
    layer1_outputs(12586) <= a and not b;
    layer1_outputs(12587) <= a and not b;
    layer1_outputs(12588) <= not (a or b);
    layer1_outputs(12589) <= '1';
    layer1_outputs(12590) <= not a;
    layer1_outputs(12591) <= not b or a;
    layer1_outputs(12592) <= '1';
    layer1_outputs(12593) <= not b or a;
    layer1_outputs(12594) <= a or b;
    layer1_outputs(12595) <= a and not b;
    layer1_outputs(12596) <= '0';
    layer1_outputs(12597) <= not a;
    layer1_outputs(12598) <= not a or b;
    layer1_outputs(12599) <= a and b;
    layer1_outputs(12600) <= not b;
    layer1_outputs(12601) <= a and not b;
    layer1_outputs(12602) <= '0';
    layer1_outputs(12603) <= not b or a;
    layer1_outputs(12604) <= a or b;
    layer1_outputs(12605) <= '0';
    layer1_outputs(12606) <= not b or a;
    layer1_outputs(12607) <= not b;
    layer1_outputs(12608) <= b and not a;
    layer1_outputs(12609) <= a or b;
    layer1_outputs(12610) <= b;
    layer1_outputs(12611) <= not (a or b);
    layer1_outputs(12612) <= not a or b;
    layer1_outputs(12613) <= not b or a;
    layer1_outputs(12614) <= '0';
    layer1_outputs(12615) <= '0';
    layer1_outputs(12616) <= a or b;
    layer1_outputs(12617) <= not a or b;
    layer1_outputs(12618) <= not a or b;
    layer1_outputs(12619) <= '1';
    layer1_outputs(12620) <= a and not b;
    layer1_outputs(12621) <= b;
    layer1_outputs(12622) <= not (a or b);
    layer1_outputs(12623) <= b and not a;
    layer1_outputs(12624) <= not a;
    layer1_outputs(12625) <= not a or b;
    layer1_outputs(12626) <= not a;
    layer1_outputs(12627) <= b and not a;
    layer1_outputs(12628) <= a;
    layer1_outputs(12629) <= a xor b;
    layer1_outputs(12630) <= not (a or b);
    layer1_outputs(12631) <= '0';
    layer1_outputs(12632) <= '0';
    layer1_outputs(12633) <= a or b;
    layer1_outputs(12634) <= a or b;
    layer1_outputs(12635) <= '1';
    layer1_outputs(12636) <= '0';
    layer1_outputs(12637) <= not (a or b);
    layer1_outputs(12638) <= b;
    layer1_outputs(12639) <= a xor b;
    layer1_outputs(12640) <= '1';
    layer1_outputs(12641) <= not (a or b);
    layer1_outputs(12642) <= a;
    layer1_outputs(12643) <= a xor b;
    layer1_outputs(12644) <= not a or b;
    layer1_outputs(12645) <= a xor b;
    layer1_outputs(12646) <= not a;
    layer1_outputs(12647) <= '0';
    layer1_outputs(12648) <= b and not a;
    layer1_outputs(12649) <= not (a or b);
    layer1_outputs(12650) <= not b or a;
    layer1_outputs(12651) <= a and b;
    layer1_outputs(12652) <= not a;
    layer1_outputs(12653) <= '1';
    layer1_outputs(12654) <= b and not a;
    layer1_outputs(12655) <= a and not b;
    layer1_outputs(12656) <= not b or a;
    layer1_outputs(12657) <= not a or b;
    layer1_outputs(12658) <= not (a and b);
    layer1_outputs(12659) <= not a or b;
    layer1_outputs(12660) <= not (a and b);
    layer1_outputs(12661) <= a or b;
    layer1_outputs(12662) <= not b or a;
    layer1_outputs(12663) <= not a or b;
    layer1_outputs(12664) <= not (a xor b);
    layer1_outputs(12665) <= b;
    layer1_outputs(12666) <= not (a xor b);
    layer1_outputs(12667) <= '1';
    layer1_outputs(12668) <= a;
    layer1_outputs(12669) <= '0';
    layer1_outputs(12670) <= not a or b;
    layer1_outputs(12671) <= not (a and b);
    layer1_outputs(12672) <= not b;
    layer1_outputs(12673) <= not (a and b);
    layer1_outputs(12674) <= a and b;
    layer1_outputs(12675) <= not a or b;
    layer1_outputs(12676) <= '1';
    layer1_outputs(12677) <= b and not a;
    layer1_outputs(12678) <= a;
    layer1_outputs(12679) <= not (a or b);
    layer1_outputs(12680) <= a and not b;
    layer1_outputs(12681) <= not a;
    layer1_outputs(12682) <= not (a or b);
    layer1_outputs(12683) <= a and not b;
    layer1_outputs(12684) <= not (a xor b);
    layer1_outputs(12685) <= a xor b;
    layer1_outputs(12686) <= not a;
    layer1_outputs(12687) <= not a;
    layer1_outputs(12688) <= '0';
    layer1_outputs(12689) <= not (a or b);
    layer1_outputs(12690) <= a and not b;
    layer1_outputs(12691) <= a and not b;
    layer1_outputs(12692) <= not b;
    layer1_outputs(12693) <= a and b;
    layer1_outputs(12694) <= not b or a;
    layer1_outputs(12695) <= a or b;
    layer1_outputs(12696) <= b;
    layer1_outputs(12697) <= not b;
    layer1_outputs(12698) <= not a;
    layer1_outputs(12699) <= b;
    layer1_outputs(12700) <= not b or a;
    layer1_outputs(12701) <= not b;
    layer1_outputs(12702) <= not b or a;
    layer1_outputs(12703) <= not b or a;
    layer1_outputs(12704) <= b;
    layer1_outputs(12705) <= a xor b;
    layer1_outputs(12706) <= not (a and b);
    layer1_outputs(12707) <= not (a xor b);
    layer1_outputs(12708) <= b;
    layer1_outputs(12709) <= a or b;
    layer1_outputs(12710) <= a and not b;
    layer1_outputs(12711) <= '0';
    layer1_outputs(12712) <= not (a and b);
    layer1_outputs(12713) <= a xor b;
    layer1_outputs(12714) <= a or b;
    layer1_outputs(12715) <= a or b;
    layer1_outputs(12716) <= not b or a;
    layer1_outputs(12717) <= b;
    layer1_outputs(12718) <= not a;
    layer1_outputs(12719) <= not b or a;
    layer1_outputs(12720) <= a xor b;
    layer1_outputs(12721) <= b;
    layer1_outputs(12722) <= b;
    layer1_outputs(12723) <= a xor b;
    layer1_outputs(12724) <= not a or b;
    layer1_outputs(12725) <= b;
    layer1_outputs(12726) <= b;
    layer1_outputs(12727) <= not b;
    layer1_outputs(12728) <= a;
    layer1_outputs(12729) <= not a or b;
    layer1_outputs(12730) <= not a;
    layer1_outputs(12731) <= a and b;
    layer1_outputs(12732) <= not b or a;
    layer1_outputs(12733) <= a or b;
    layer1_outputs(12734) <= '0';
    layer1_outputs(12735) <= '1';
    layer1_outputs(12736) <= a xor b;
    layer1_outputs(12737) <= not (a and b);
    layer1_outputs(12738) <= not a or b;
    layer1_outputs(12739) <= a and not b;
    layer1_outputs(12740) <= b;
    layer1_outputs(12741) <= not b;
    layer1_outputs(12742) <= a or b;
    layer1_outputs(12743) <= a;
    layer1_outputs(12744) <= not a or b;
    layer1_outputs(12745) <= b and not a;
    layer1_outputs(12746) <= b;
    layer1_outputs(12747) <= not b;
    layer1_outputs(12748) <= not a or b;
    layer1_outputs(12749) <= not a;
    layer1_outputs(12750) <= not b;
    layer1_outputs(12751) <= not b;
    layer1_outputs(12752) <= a and not b;
    layer1_outputs(12753) <= not b;
    layer1_outputs(12754) <= a and b;
    layer1_outputs(12755) <= a and not b;
    layer1_outputs(12756) <= not a;
    layer1_outputs(12757) <= not (a and b);
    layer1_outputs(12758) <= not b or a;
    layer1_outputs(12759) <= not b;
    layer1_outputs(12760) <= not a;
    layer1_outputs(12761) <= not a or b;
    layer1_outputs(12762) <= a xor b;
    layer1_outputs(12763) <= not b or a;
    layer1_outputs(12764) <= not (a and b);
    layer1_outputs(12765) <= b;
    layer1_outputs(12766) <= a and b;
    layer1_outputs(12767) <= a and not b;
    layer1_outputs(12768) <= not (a and b);
    layer1_outputs(12769) <= not (a or b);
    layer1_outputs(12770) <= a or b;
    layer1_outputs(12771) <= a or b;
    layer1_outputs(12772) <= not (a xor b);
    layer1_outputs(12773) <= '0';
    layer1_outputs(12774) <= '0';
    layer1_outputs(12775) <= b and not a;
    layer1_outputs(12776) <= b;
    layer1_outputs(12777) <= b and not a;
    layer1_outputs(12778) <= not (a and b);
    layer1_outputs(12779) <= b;
    layer1_outputs(12780) <= a xor b;
    layer1_outputs(12781) <= not (a and b);
    layer1_outputs(12782) <= '0';
    layer1_outputs(12783) <= '1';
    layer1_outputs(12784) <= not b or a;
    layer1_outputs(12785) <= not b;
    layer1_outputs(12786) <= a;
    layer1_outputs(12787) <= not b or a;
    layer1_outputs(12788) <= not b;
    layer1_outputs(12789) <= not a;
    layer1_outputs(12790) <= not b;
    layer1_outputs(12791) <= b;
    layer1_outputs(12792) <= not b;
    layer1_outputs(12793) <= a xor b;
    layer1_outputs(12794) <= not (a and b);
    layer1_outputs(12795) <= b and not a;
    layer1_outputs(12796) <= '1';
    layer1_outputs(12797) <= not a or b;
    layer1_outputs(12798) <= a and b;
    layer1_outputs(12799) <= not a or b;
    layer2_outputs(0) <= not a;
    layer2_outputs(1) <= a xor b;
    layer2_outputs(2) <= '1';
    layer2_outputs(3) <= not a or b;
    layer2_outputs(4) <= a xor b;
    layer2_outputs(5) <= a and b;
    layer2_outputs(6) <= a and not b;
    layer2_outputs(7) <= '0';
    layer2_outputs(8) <= a or b;
    layer2_outputs(9) <= a or b;
    layer2_outputs(10) <= a or b;
    layer2_outputs(11) <= not (a xor b);
    layer2_outputs(12) <= a;
    layer2_outputs(13) <= '1';
    layer2_outputs(14) <= '0';
    layer2_outputs(15) <= not b;
    layer2_outputs(16) <= '0';
    layer2_outputs(17) <= '0';
    layer2_outputs(18) <= a or b;
    layer2_outputs(19) <= not a;
    layer2_outputs(20) <= a or b;
    layer2_outputs(21) <= b and not a;
    layer2_outputs(22) <= not a;
    layer2_outputs(23) <= not b;
    layer2_outputs(24) <= a and not b;
    layer2_outputs(25) <= a xor b;
    layer2_outputs(26) <= b and not a;
    layer2_outputs(27) <= a xor b;
    layer2_outputs(28) <= a and b;
    layer2_outputs(29) <= a and not b;
    layer2_outputs(30) <= not (a or b);
    layer2_outputs(31) <= a and not b;
    layer2_outputs(32) <= not a;
    layer2_outputs(33) <= a and not b;
    layer2_outputs(34) <= not a or b;
    layer2_outputs(35) <= a and b;
    layer2_outputs(36) <= a and b;
    layer2_outputs(37) <= b and not a;
    layer2_outputs(38) <= a or b;
    layer2_outputs(39) <= b;
    layer2_outputs(40) <= b;
    layer2_outputs(41) <= not a;
    layer2_outputs(42) <= '0';
    layer2_outputs(43) <= '1';
    layer2_outputs(44) <= '1';
    layer2_outputs(45) <= b;
    layer2_outputs(46) <= a xor b;
    layer2_outputs(47) <= a;
    layer2_outputs(48) <= b and not a;
    layer2_outputs(49) <= not a or b;
    layer2_outputs(50) <= a xor b;
    layer2_outputs(51) <= not b;
    layer2_outputs(52) <= a and not b;
    layer2_outputs(53) <= a or b;
    layer2_outputs(54) <= not b;
    layer2_outputs(55) <= not (a or b);
    layer2_outputs(56) <= a;
    layer2_outputs(57) <= not b;
    layer2_outputs(58) <= a or b;
    layer2_outputs(59) <= not a or b;
    layer2_outputs(60) <= not (a xor b);
    layer2_outputs(61) <= not b;
    layer2_outputs(62) <= not (a and b);
    layer2_outputs(63) <= not (a and b);
    layer2_outputs(64) <= not b;
    layer2_outputs(65) <= b;
    layer2_outputs(66) <= not a;
    layer2_outputs(67) <= not (a or b);
    layer2_outputs(68) <= not (a or b);
    layer2_outputs(69) <= a xor b;
    layer2_outputs(70) <= b and not a;
    layer2_outputs(71) <= a xor b;
    layer2_outputs(72) <= not a;
    layer2_outputs(73) <= not a;
    layer2_outputs(74) <= not a;
    layer2_outputs(75) <= a;
    layer2_outputs(76) <= not (a or b);
    layer2_outputs(77) <= not b;
    layer2_outputs(78) <= b and not a;
    layer2_outputs(79) <= not (a or b);
    layer2_outputs(80) <= not b or a;
    layer2_outputs(81) <= not (a and b);
    layer2_outputs(82) <= '0';
    layer2_outputs(83) <= a xor b;
    layer2_outputs(84) <= not a or b;
    layer2_outputs(85) <= not (a and b);
    layer2_outputs(86) <= b and not a;
    layer2_outputs(87) <= b;
    layer2_outputs(88) <= '0';
    layer2_outputs(89) <= a;
    layer2_outputs(90) <= not b;
    layer2_outputs(91) <= b;
    layer2_outputs(92) <= not b;
    layer2_outputs(93) <= not (a and b);
    layer2_outputs(94) <= not a;
    layer2_outputs(95) <= '0';
    layer2_outputs(96) <= a and not b;
    layer2_outputs(97) <= a and not b;
    layer2_outputs(98) <= a and not b;
    layer2_outputs(99) <= a and not b;
    layer2_outputs(100) <= not a;
    layer2_outputs(101) <= '1';
    layer2_outputs(102) <= a;
    layer2_outputs(103) <= not (a and b);
    layer2_outputs(104) <= a and b;
    layer2_outputs(105) <= not b;
    layer2_outputs(106) <= not b;
    layer2_outputs(107) <= a or b;
    layer2_outputs(108) <= not b or a;
    layer2_outputs(109) <= not (a or b);
    layer2_outputs(110) <= '1';
    layer2_outputs(111) <= '1';
    layer2_outputs(112) <= not a or b;
    layer2_outputs(113) <= b;
    layer2_outputs(114) <= b and not a;
    layer2_outputs(115) <= not b or a;
    layer2_outputs(116) <= a or b;
    layer2_outputs(117) <= not b or a;
    layer2_outputs(118) <= a and b;
    layer2_outputs(119) <= a xor b;
    layer2_outputs(120) <= '0';
    layer2_outputs(121) <= '1';
    layer2_outputs(122) <= not a;
    layer2_outputs(123) <= '0';
    layer2_outputs(124) <= '1';
    layer2_outputs(125) <= not (a or b);
    layer2_outputs(126) <= not a or b;
    layer2_outputs(127) <= not b;
    layer2_outputs(128) <= '1';
    layer2_outputs(129) <= a or b;
    layer2_outputs(130) <= a or b;
    layer2_outputs(131) <= '1';
    layer2_outputs(132) <= a or b;
    layer2_outputs(133) <= not b;
    layer2_outputs(134) <= b;
    layer2_outputs(135) <= not (a xor b);
    layer2_outputs(136) <= not b or a;
    layer2_outputs(137) <= a or b;
    layer2_outputs(138) <= not a;
    layer2_outputs(139) <= not (a or b);
    layer2_outputs(140) <= not a;
    layer2_outputs(141) <= b and not a;
    layer2_outputs(142) <= not (a and b);
    layer2_outputs(143) <= not (a and b);
    layer2_outputs(144) <= not (a or b);
    layer2_outputs(145) <= not (a xor b);
    layer2_outputs(146) <= not (a and b);
    layer2_outputs(147) <= '1';
    layer2_outputs(148) <= not (a or b);
    layer2_outputs(149) <= not a;
    layer2_outputs(150) <= a xor b;
    layer2_outputs(151) <= b and not a;
    layer2_outputs(152) <= not b;
    layer2_outputs(153) <= a xor b;
    layer2_outputs(154) <= not (a xor b);
    layer2_outputs(155) <= not b;
    layer2_outputs(156) <= a or b;
    layer2_outputs(157) <= not a;
    layer2_outputs(158) <= not (a or b);
    layer2_outputs(159) <= b and not a;
    layer2_outputs(160) <= not (a or b);
    layer2_outputs(161) <= b and not a;
    layer2_outputs(162) <= not a;
    layer2_outputs(163) <= not (a and b);
    layer2_outputs(164) <= not b;
    layer2_outputs(165) <= b;
    layer2_outputs(166) <= '1';
    layer2_outputs(167) <= a or b;
    layer2_outputs(168) <= b and not a;
    layer2_outputs(169) <= not b or a;
    layer2_outputs(170) <= not b or a;
    layer2_outputs(171) <= '0';
    layer2_outputs(172) <= not (a and b);
    layer2_outputs(173) <= not b or a;
    layer2_outputs(174) <= not (a or b);
    layer2_outputs(175) <= not b or a;
    layer2_outputs(176) <= not b or a;
    layer2_outputs(177) <= not b;
    layer2_outputs(178) <= a or b;
    layer2_outputs(179) <= a and not b;
    layer2_outputs(180) <= a and not b;
    layer2_outputs(181) <= not b;
    layer2_outputs(182) <= not (a or b);
    layer2_outputs(183) <= not b;
    layer2_outputs(184) <= not (a or b);
    layer2_outputs(185) <= not b;
    layer2_outputs(186) <= a;
    layer2_outputs(187) <= not (a and b);
    layer2_outputs(188) <= a and not b;
    layer2_outputs(189) <= '0';
    layer2_outputs(190) <= not b;
    layer2_outputs(191) <= a or b;
    layer2_outputs(192) <= '0';
    layer2_outputs(193) <= '1';
    layer2_outputs(194) <= a or b;
    layer2_outputs(195) <= b and not a;
    layer2_outputs(196) <= b;
    layer2_outputs(197) <= not a or b;
    layer2_outputs(198) <= a and b;
    layer2_outputs(199) <= a and not b;
    layer2_outputs(200) <= not (a or b);
    layer2_outputs(201) <= not (a and b);
    layer2_outputs(202) <= a;
    layer2_outputs(203) <= a or b;
    layer2_outputs(204) <= not b;
    layer2_outputs(205) <= not b;
    layer2_outputs(206) <= not b;
    layer2_outputs(207) <= not a;
    layer2_outputs(208) <= a;
    layer2_outputs(209) <= a;
    layer2_outputs(210) <= b;
    layer2_outputs(211) <= b and not a;
    layer2_outputs(212) <= not a;
    layer2_outputs(213) <= b;
    layer2_outputs(214) <= not (a xor b);
    layer2_outputs(215) <= b;
    layer2_outputs(216) <= not a;
    layer2_outputs(217) <= not a or b;
    layer2_outputs(218) <= a;
    layer2_outputs(219) <= b and not a;
    layer2_outputs(220) <= not a or b;
    layer2_outputs(221) <= '1';
    layer2_outputs(222) <= b;
    layer2_outputs(223) <= not b;
    layer2_outputs(224) <= not b;
    layer2_outputs(225) <= b;
    layer2_outputs(226) <= not (a and b);
    layer2_outputs(227) <= '0';
    layer2_outputs(228) <= not a;
    layer2_outputs(229) <= '1';
    layer2_outputs(230) <= not (a or b);
    layer2_outputs(231) <= not (a xor b);
    layer2_outputs(232) <= '0';
    layer2_outputs(233) <= not a;
    layer2_outputs(234) <= '1';
    layer2_outputs(235) <= not b or a;
    layer2_outputs(236) <= b;
    layer2_outputs(237) <= b;
    layer2_outputs(238) <= a;
    layer2_outputs(239) <= a and not b;
    layer2_outputs(240) <= a and not b;
    layer2_outputs(241) <= not a;
    layer2_outputs(242) <= b;
    layer2_outputs(243) <= a;
    layer2_outputs(244) <= b and not a;
    layer2_outputs(245) <= a or b;
    layer2_outputs(246) <= not b or a;
    layer2_outputs(247) <= a and not b;
    layer2_outputs(248) <= '0';
    layer2_outputs(249) <= a;
    layer2_outputs(250) <= a and not b;
    layer2_outputs(251) <= b and not a;
    layer2_outputs(252) <= a or b;
    layer2_outputs(253) <= '0';
    layer2_outputs(254) <= not (a xor b);
    layer2_outputs(255) <= b;
    layer2_outputs(256) <= not (a and b);
    layer2_outputs(257) <= a or b;
    layer2_outputs(258) <= a;
    layer2_outputs(259) <= not b;
    layer2_outputs(260) <= not (a and b);
    layer2_outputs(261) <= a and not b;
    layer2_outputs(262) <= not b;
    layer2_outputs(263) <= b and not a;
    layer2_outputs(264) <= a xor b;
    layer2_outputs(265) <= a and b;
    layer2_outputs(266) <= not (a xor b);
    layer2_outputs(267) <= a or b;
    layer2_outputs(268) <= a and not b;
    layer2_outputs(269) <= not (a or b);
    layer2_outputs(270) <= not a or b;
    layer2_outputs(271) <= b and not a;
    layer2_outputs(272) <= not b;
    layer2_outputs(273) <= a and not b;
    layer2_outputs(274) <= not b;
    layer2_outputs(275) <= b and not a;
    layer2_outputs(276) <= not (a and b);
    layer2_outputs(277) <= a;
    layer2_outputs(278) <= a;
    layer2_outputs(279) <= not b;
    layer2_outputs(280) <= not b;
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= not a;
    layer2_outputs(283) <= not (a and b);
    layer2_outputs(284) <= not a;
    layer2_outputs(285) <= a xor b;
    layer2_outputs(286) <= a;
    layer2_outputs(287) <= a and not b;
    layer2_outputs(288) <= not b or a;
    layer2_outputs(289) <= a;
    layer2_outputs(290) <= not b;
    layer2_outputs(291) <= not b or a;
    layer2_outputs(292) <= not a;
    layer2_outputs(293) <= not (a and b);
    layer2_outputs(294) <= not (a and b);
    layer2_outputs(295) <= b;
    layer2_outputs(296) <= '1';
    layer2_outputs(297) <= a and not b;
    layer2_outputs(298) <= a or b;
    layer2_outputs(299) <= not (a and b);
    layer2_outputs(300) <= b and not a;
    layer2_outputs(301) <= '1';
    layer2_outputs(302) <= not (a or b);
    layer2_outputs(303) <= not (a and b);
    layer2_outputs(304) <= a and not b;
    layer2_outputs(305) <= b and not a;
    layer2_outputs(306) <= '1';
    layer2_outputs(307) <= a xor b;
    layer2_outputs(308) <= a and not b;
    layer2_outputs(309) <= '1';
    layer2_outputs(310) <= not (a or b);
    layer2_outputs(311) <= a and b;
    layer2_outputs(312) <= not (a and b);
    layer2_outputs(313) <= b and not a;
    layer2_outputs(314) <= a and b;
    layer2_outputs(315) <= not a;
    layer2_outputs(316) <= not (a xor b);
    layer2_outputs(317) <= a;
    layer2_outputs(318) <= not (a or b);
    layer2_outputs(319) <= not (a xor b);
    layer2_outputs(320) <= b and not a;
    layer2_outputs(321) <= a;
    layer2_outputs(322) <= not a or b;
    layer2_outputs(323) <= not b or a;
    layer2_outputs(324) <= b;
    layer2_outputs(325) <= '0';
    layer2_outputs(326) <= a xor b;
    layer2_outputs(327) <= b and not a;
    layer2_outputs(328) <= '0';
    layer2_outputs(329) <= not (a or b);
    layer2_outputs(330) <= not a;
    layer2_outputs(331) <= not b;
    layer2_outputs(332) <= a and b;
    layer2_outputs(333) <= not (a and b);
    layer2_outputs(334) <= not (a or b);
    layer2_outputs(335) <= a and b;
    layer2_outputs(336) <= not (a and b);
    layer2_outputs(337) <= '1';
    layer2_outputs(338) <= not a or b;
    layer2_outputs(339) <= a and not b;
    layer2_outputs(340) <= not (a or b);
    layer2_outputs(341) <= '0';
    layer2_outputs(342) <= '1';
    layer2_outputs(343) <= b and not a;
    layer2_outputs(344) <= not b or a;
    layer2_outputs(345) <= not (a and b);
    layer2_outputs(346) <= not a or b;
    layer2_outputs(347) <= a and b;
    layer2_outputs(348) <= not a or b;
    layer2_outputs(349) <= a or b;
    layer2_outputs(350) <= a or b;
    layer2_outputs(351) <= b;
    layer2_outputs(352) <= a and b;
    layer2_outputs(353) <= not a or b;
    layer2_outputs(354) <= not b;
    layer2_outputs(355) <= not a;
    layer2_outputs(356) <= b and not a;
    layer2_outputs(357) <= not a;
    layer2_outputs(358) <= not a;
    layer2_outputs(359) <= b;
    layer2_outputs(360) <= a or b;
    layer2_outputs(361) <= not (a xor b);
    layer2_outputs(362) <= a and b;
    layer2_outputs(363) <= not b or a;
    layer2_outputs(364) <= a or b;
    layer2_outputs(365) <= not b;
    layer2_outputs(366) <= b and not a;
    layer2_outputs(367) <= not (a or b);
    layer2_outputs(368) <= not a or b;
    layer2_outputs(369) <= not b;
    layer2_outputs(370) <= not (a and b);
    layer2_outputs(371) <= not a;
    layer2_outputs(372) <= a and not b;
    layer2_outputs(373) <= a and not b;
    layer2_outputs(374) <= a xor b;
    layer2_outputs(375) <= not b;
    layer2_outputs(376) <= a and b;
    layer2_outputs(377) <= b;
    layer2_outputs(378) <= b;
    layer2_outputs(379) <= not (a and b);
    layer2_outputs(380) <= not a;
    layer2_outputs(381) <= not (a and b);
    layer2_outputs(382) <= '0';
    layer2_outputs(383) <= a and b;
    layer2_outputs(384) <= '1';
    layer2_outputs(385) <= not a or b;
    layer2_outputs(386) <= a and not b;
    layer2_outputs(387) <= '1';
    layer2_outputs(388) <= '0';
    layer2_outputs(389) <= not a or b;
    layer2_outputs(390) <= a and b;
    layer2_outputs(391) <= a or b;
    layer2_outputs(392) <= not (a or b);
    layer2_outputs(393) <= not (a xor b);
    layer2_outputs(394) <= not b;
    layer2_outputs(395) <= not (a and b);
    layer2_outputs(396) <= '0';
    layer2_outputs(397) <= '0';
    layer2_outputs(398) <= a or b;
    layer2_outputs(399) <= b;
    layer2_outputs(400) <= not b or a;
    layer2_outputs(401) <= not b or a;
    layer2_outputs(402) <= b and not a;
    layer2_outputs(403) <= a xor b;
    layer2_outputs(404) <= not b or a;
    layer2_outputs(405) <= not (a and b);
    layer2_outputs(406) <= not a;
    layer2_outputs(407) <= not (a xor b);
    layer2_outputs(408) <= a xor b;
    layer2_outputs(409) <= a or b;
    layer2_outputs(410) <= '0';
    layer2_outputs(411) <= a and not b;
    layer2_outputs(412) <= not a;
    layer2_outputs(413) <= not b;
    layer2_outputs(414) <= a or b;
    layer2_outputs(415) <= a or b;
    layer2_outputs(416) <= a and not b;
    layer2_outputs(417) <= not a;
    layer2_outputs(418) <= a;
    layer2_outputs(419) <= not a or b;
    layer2_outputs(420) <= not a;
    layer2_outputs(421) <= not a;
    layer2_outputs(422) <= not a or b;
    layer2_outputs(423) <= not (a or b);
    layer2_outputs(424) <= '0';
    layer2_outputs(425) <= '1';
    layer2_outputs(426) <= not b;
    layer2_outputs(427) <= '0';
    layer2_outputs(428) <= a and not b;
    layer2_outputs(429) <= not a;
    layer2_outputs(430) <= a;
    layer2_outputs(431) <= not b;
    layer2_outputs(432) <= a or b;
    layer2_outputs(433) <= '0';
    layer2_outputs(434) <= a;
    layer2_outputs(435) <= a or b;
    layer2_outputs(436) <= '1';
    layer2_outputs(437) <= not b or a;
    layer2_outputs(438) <= b and not a;
    layer2_outputs(439) <= b;
    layer2_outputs(440) <= not b;
    layer2_outputs(441) <= a;
    layer2_outputs(442) <= '0';
    layer2_outputs(443) <= a and b;
    layer2_outputs(444) <= not b;
    layer2_outputs(445) <= not (a xor b);
    layer2_outputs(446) <= not b;
    layer2_outputs(447) <= '1';
    layer2_outputs(448) <= a;
    layer2_outputs(449) <= '1';
    layer2_outputs(450) <= a and not b;
    layer2_outputs(451) <= '0';
    layer2_outputs(452) <= '0';
    layer2_outputs(453) <= b;
    layer2_outputs(454) <= not b or a;
    layer2_outputs(455) <= not a;
    layer2_outputs(456) <= not a;
    layer2_outputs(457) <= '0';
    layer2_outputs(458) <= not (a or b);
    layer2_outputs(459) <= a and not b;
    layer2_outputs(460) <= a;
    layer2_outputs(461) <= a and not b;
    layer2_outputs(462) <= a or b;
    layer2_outputs(463) <= b and not a;
    layer2_outputs(464) <= not (a or b);
    layer2_outputs(465) <= not b;
    layer2_outputs(466) <= not a;
    layer2_outputs(467) <= a and b;
    layer2_outputs(468) <= not (a and b);
    layer2_outputs(469) <= a or b;
    layer2_outputs(470) <= not (a xor b);
    layer2_outputs(471) <= a or b;
    layer2_outputs(472) <= b;
    layer2_outputs(473) <= a and not b;
    layer2_outputs(474) <= b and not a;
    layer2_outputs(475) <= b and not a;
    layer2_outputs(476) <= a and b;
    layer2_outputs(477) <= not a;
    layer2_outputs(478) <= a and b;
    layer2_outputs(479) <= not a;
    layer2_outputs(480) <= '0';
    layer2_outputs(481) <= '1';
    layer2_outputs(482) <= b and not a;
    layer2_outputs(483) <= not b or a;
    layer2_outputs(484) <= not (a or b);
    layer2_outputs(485) <= a;
    layer2_outputs(486) <= a or b;
    layer2_outputs(487) <= not a or b;
    layer2_outputs(488) <= not a or b;
    layer2_outputs(489) <= not b;
    layer2_outputs(490) <= a;
    layer2_outputs(491) <= a;
    layer2_outputs(492) <= a or b;
    layer2_outputs(493) <= not a;
    layer2_outputs(494) <= not b;
    layer2_outputs(495) <= a and not b;
    layer2_outputs(496) <= not a;
    layer2_outputs(497) <= not b;
    layer2_outputs(498) <= '0';
    layer2_outputs(499) <= b and not a;
    layer2_outputs(500) <= a;
    layer2_outputs(501) <= not (a or b);
    layer2_outputs(502) <= b and not a;
    layer2_outputs(503) <= a and b;
    layer2_outputs(504) <= '1';
    layer2_outputs(505) <= a;
    layer2_outputs(506) <= b;
    layer2_outputs(507) <= a or b;
    layer2_outputs(508) <= a and b;
    layer2_outputs(509) <= a and b;
    layer2_outputs(510) <= not (a and b);
    layer2_outputs(511) <= '0';
    layer2_outputs(512) <= b;
    layer2_outputs(513) <= a;
    layer2_outputs(514) <= not a;
    layer2_outputs(515) <= b;
    layer2_outputs(516) <= '1';
    layer2_outputs(517) <= b;
    layer2_outputs(518) <= not b or a;
    layer2_outputs(519) <= a or b;
    layer2_outputs(520) <= not a or b;
    layer2_outputs(521) <= a or b;
    layer2_outputs(522) <= not (a xor b);
    layer2_outputs(523) <= b;
    layer2_outputs(524) <= not (a xor b);
    layer2_outputs(525) <= a xor b;
    layer2_outputs(526) <= '0';
    layer2_outputs(527) <= a;
    layer2_outputs(528) <= not a or b;
    layer2_outputs(529) <= a xor b;
    layer2_outputs(530) <= not (a and b);
    layer2_outputs(531) <= a and not b;
    layer2_outputs(532) <= '1';
    layer2_outputs(533) <= a and not b;
    layer2_outputs(534) <= a or b;
    layer2_outputs(535) <= a or b;
    layer2_outputs(536) <= not (a and b);
    layer2_outputs(537) <= a and not b;
    layer2_outputs(538) <= not b or a;
    layer2_outputs(539) <= not (a or b);
    layer2_outputs(540) <= not (a or b);
    layer2_outputs(541) <= not (a or b);
    layer2_outputs(542) <= a and b;
    layer2_outputs(543) <= not (a xor b);
    layer2_outputs(544) <= not a;
    layer2_outputs(545) <= a and b;
    layer2_outputs(546) <= not a or b;
    layer2_outputs(547) <= '1';
    layer2_outputs(548) <= a or b;
    layer2_outputs(549) <= not b;
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= a;
    layer2_outputs(552) <= not b or a;
    layer2_outputs(553) <= not (a or b);
    layer2_outputs(554) <= b and not a;
    layer2_outputs(555) <= a;
    layer2_outputs(556) <= not (a or b);
    layer2_outputs(557) <= b and not a;
    layer2_outputs(558) <= not (a or b);
    layer2_outputs(559) <= not b or a;
    layer2_outputs(560) <= not (a and b);
    layer2_outputs(561) <= a;
    layer2_outputs(562) <= a or b;
    layer2_outputs(563) <= not (a and b);
    layer2_outputs(564) <= not a or b;
    layer2_outputs(565) <= a and not b;
    layer2_outputs(566) <= not (a xor b);
    layer2_outputs(567) <= not a or b;
    layer2_outputs(568) <= not (a or b);
    layer2_outputs(569) <= not b or a;
    layer2_outputs(570) <= not (a xor b);
    layer2_outputs(571) <= b;
    layer2_outputs(572) <= a xor b;
    layer2_outputs(573) <= not b;
    layer2_outputs(574) <= not (a or b);
    layer2_outputs(575) <= a;
    layer2_outputs(576) <= a and not b;
    layer2_outputs(577) <= not b;
    layer2_outputs(578) <= not (a or b);
    layer2_outputs(579) <= b;
    layer2_outputs(580) <= not (a or b);
    layer2_outputs(581) <= a or b;
    layer2_outputs(582) <= a or b;
    layer2_outputs(583) <= '1';
    layer2_outputs(584) <= not (a and b);
    layer2_outputs(585) <= not a or b;
    layer2_outputs(586) <= not b;
    layer2_outputs(587) <= '1';
    layer2_outputs(588) <= not b or a;
    layer2_outputs(589) <= not a;
    layer2_outputs(590) <= a;
    layer2_outputs(591) <= not b;
    layer2_outputs(592) <= not b or a;
    layer2_outputs(593) <= '1';
    layer2_outputs(594) <= b and not a;
    layer2_outputs(595) <= '1';
    layer2_outputs(596) <= '0';
    layer2_outputs(597) <= not a or b;
    layer2_outputs(598) <= not b or a;
    layer2_outputs(599) <= not (a or b);
    layer2_outputs(600) <= '0';
    layer2_outputs(601) <= a;
    layer2_outputs(602) <= not a;
    layer2_outputs(603) <= not a or b;
    layer2_outputs(604) <= a or b;
    layer2_outputs(605) <= a and b;
    layer2_outputs(606) <= not b;
    layer2_outputs(607) <= a or b;
    layer2_outputs(608) <= not a or b;
    layer2_outputs(609) <= b;
    layer2_outputs(610) <= a xor b;
    layer2_outputs(611) <= a;
    layer2_outputs(612) <= not (a xor b);
    layer2_outputs(613) <= not b or a;
    layer2_outputs(614) <= a and b;
    layer2_outputs(615) <= a or b;
    layer2_outputs(616) <= not a;
    layer2_outputs(617) <= a or b;
    layer2_outputs(618) <= '1';
    layer2_outputs(619) <= not (a and b);
    layer2_outputs(620) <= a or b;
    layer2_outputs(621) <= b and not a;
    layer2_outputs(622) <= '1';
    layer2_outputs(623) <= not a;
    layer2_outputs(624) <= a and not b;
    layer2_outputs(625) <= not b or a;
    layer2_outputs(626) <= a;
    layer2_outputs(627) <= not b or a;
    layer2_outputs(628) <= not (a xor b);
    layer2_outputs(629) <= not a or b;
    layer2_outputs(630) <= not b;
    layer2_outputs(631) <= a and not b;
    layer2_outputs(632) <= not b;
    layer2_outputs(633) <= not b;
    layer2_outputs(634) <= '1';
    layer2_outputs(635) <= not (a and b);
    layer2_outputs(636) <= not b;
    layer2_outputs(637) <= not b;
    layer2_outputs(638) <= a;
    layer2_outputs(639) <= '0';
    layer2_outputs(640) <= a and not b;
    layer2_outputs(641) <= b and not a;
    layer2_outputs(642) <= a xor b;
    layer2_outputs(643) <= not b or a;
    layer2_outputs(644) <= a xor b;
    layer2_outputs(645) <= not b;
    layer2_outputs(646) <= '0';
    layer2_outputs(647) <= not b or a;
    layer2_outputs(648) <= not (a and b);
    layer2_outputs(649) <= not a;
    layer2_outputs(650) <= a and b;
    layer2_outputs(651) <= not (a xor b);
    layer2_outputs(652) <= not a or b;
    layer2_outputs(653) <= not (a or b);
    layer2_outputs(654) <= b;
    layer2_outputs(655) <= '1';
    layer2_outputs(656) <= not a;
    layer2_outputs(657) <= b;
    layer2_outputs(658) <= a and not b;
    layer2_outputs(659) <= b;
    layer2_outputs(660) <= b and not a;
    layer2_outputs(661) <= b and not a;
    layer2_outputs(662) <= b;
    layer2_outputs(663) <= not a;
    layer2_outputs(664) <= not (a xor b);
    layer2_outputs(665) <= not b or a;
    layer2_outputs(666) <= not (a or b);
    layer2_outputs(667) <= '1';
    layer2_outputs(668) <= not b;
    layer2_outputs(669) <= '1';
    layer2_outputs(670) <= a xor b;
    layer2_outputs(671) <= '1';
    layer2_outputs(672) <= not (a and b);
    layer2_outputs(673) <= not b or a;
    layer2_outputs(674) <= not a;
    layer2_outputs(675) <= a;
    layer2_outputs(676) <= a and not b;
    layer2_outputs(677) <= not a or b;
    layer2_outputs(678) <= a and not b;
    layer2_outputs(679) <= a xor b;
    layer2_outputs(680) <= not a or b;
    layer2_outputs(681) <= not (a and b);
    layer2_outputs(682) <= not b or a;
    layer2_outputs(683) <= a and b;
    layer2_outputs(684) <= not a or b;
    layer2_outputs(685) <= not (a and b);
    layer2_outputs(686) <= not (a xor b);
    layer2_outputs(687) <= not b;
    layer2_outputs(688) <= a and not b;
    layer2_outputs(689) <= not (a and b);
    layer2_outputs(690) <= not (a or b);
    layer2_outputs(691) <= not a or b;
    layer2_outputs(692) <= not a or b;
    layer2_outputs(693) <= not a;
    layer2_outputs(694) <= '1';
    layer2_outputs(695) <= a xor b;
    layer2_outputs(696) <= a and not b;
    layer2_outputs(697) <= not a;
    layer2_outputs(698) <= a or b;
    layer2_outputs(699) <= not a;
    layer2_outputs(700) <= a or b;
    layer2_outputs(701) <= not a or b;
    layer2_outputs(702) <= b and not a;
    layer2_outputs(703) <= not b or a;
    layer2_outputs(704) <= a and b;
    layer2_outputs(705) <= not (a or b);
    layer2_outputs(706) <= not (a and b);
    layer2_outputs(707) <= a and not b;
    layer2_outputs(708) <= '1';
    layer2_outputs(709) <= a and not b;
    layer2_outputs(710) <= not (a or b);
    layer2_outputs(711) <= not a;
    layer2_outputs(712) <= not a or b;
    layer2_outputs(713) <= not (a and b);
    layer2_outputs(714) <= not (a and b);
    layer2_outputs(715) <= '1';
    layer2_outputs(716) <= not a;
    layer2_outputs(717) <= a or b;
    layer2_outputs(718) <= a;
    layer2_outputs(719) <= '0';
    layer2_outputs(720) <= a and not b;
    layer2_outputs(721) <= not (a and b);
    layer2_outputs(722) <= b;
    layer2_outputs(723) <= '0';
    layer2_outputs(724) <= a xor b;
    layer2_outputs(725) <= not (a and b);
    layer2_outputs(726) <= a and b;
    layer2_outputs(727) <= not b;
    layer2_outputs(728) <= b;
    layer2_outputs(729) <= not (a xor b);
    layer2_outputs(730) <= '0';
    layer2_outputs(731) <= '1';
    layer2_outputs(732) <= not b or a;
    layer2_outputs(733) <= '0';
    layer2_outputs(734) <= a or b;
    layer2_outputs(735) <= not a;
    layer2_outputs(736) <= a and not b;
    layer2_outputs(737) <= not b;
    layer2_outputs(738) <= not (a xor b);
    layer2_outputs(739) <= not b;
    layer2_outputs(740) <= not a;
    layer2_outputs(741) <= '0';
    layer2_outputs(742) <= not a;
    layer2_outputs(743) <= not a;
    layer2_outputs(744) <= b;
    layer2_outputs(745) <= not a or b;
    layer2_outputs(746) <= not b;
    layer2_outputs(747) <= not a or b;
    layer2_outputs(748) <= a xor b;
    layer2_outputs(749) <= b and not a;
    layer2_outputs(750) <= not b or a;
    layer2_outputs(751) <= a or b;
    layer2_outputs(752) <= not a;
    layer2_outputs(753) <= not b or a;
    layer2_outputs(754) <= a;
    layer2_outputs(755) <= not (a and b);
    layer2_outputs(756) <= not (a or b);
    layer2_outputs(757) <= not b;
    layer2_outputs(758) <= b;
    layer2_outputs(759) <= not (a or b);
    layer2_outputs(760) <= b;
    layer2_outputs(761) <= not a;
    layer2_outputs(762) <= '0';
    layer2_outputs(763) <= not a;
    layer2_outputs(764) <= b and not a;
    layer2_outputs(765) <= a and not b;
    layer2_outputs(766) <= not (a or b);
    layer2_outputs(767) <= b and not a;
    layer2_outputs(768) <= not b;
    layer2_outputs(769) <= b and not a;
    layer2_outputs(770) <= b and not a;
    layer2_outputs(771) <= b and not a;
    layer2_outputs(772) <= '0';
    layer2_outputs(773) <= a and not b;
    layer2_outputs(774) <= '0';
    layer2_outputs(775) <= not b;
    layer2_outputs(776) <= not b or a;
    layer2_outputs(777) <= a and not b;
    layer2_outputs(778) <= a and not b;
    layer2_outputs(779) <= not (a or b);
    layer2_outputs(780) <= '0';
    layer2_outputs(781) <= not b;
    layer2_outputs(782) <= '1';
    layer2_outputs(783) <= b and not a;
    layer2_outputs(784) <= a and b;
    layer2_outputs(785) <= b;
    layer2_outputs(786) <= not b;
    layer2_outputs(787) <= '0';
    layer2_outputs(788) <= not (a and b);
    layer2_outputs(789) <= not b;
    layer2_outputs(790) <= not a;
    layer2_outputs(791) <= not a or b;
    layer2_outputs(792) <= not a;
    layer2_outputs(793) <= b and not a;
    layer2_outputs(794) <= '0';
    layer2_outputs(795) <= a;
    layer2_outputs(796) <= a xor b;
    layer2_outputs(797) <= a and not b;
    layer2_outputs(798) <= a xor b;
    layer2_outputs(799) <= not b or a;
    layer2_outputs(800) <= not b or a;
    layer2_outputs(801) <= a;
    layer2_outputs(802) <= b;
    layer2_outputs(803) <= not a;
    layer2_outputs(804) <= a or b;
    layer2_outputs(805) <= not b or a;
    layer2_outputs(806) <= not b;
    layer2_outputs(807) <= b;
    layer2_outputs(808) <= '1';
    layer2_outputs(809) <= a or b;
    layer2_outputs(810) <= not b or a;
    layer2_outputs(811) <= a;
    layer2_outputs(812) <= not b or a;
    layer2_outputs(813) <= b;
    layer2_outputs(814) <= b;
    layer2_outputs(815) <= not (a and b);
    layer2_outputs(816) <= a xor b;
    layer2_outputs(817) <= not b;
    layer2_outputs(818) <= not b;
    layer2_outputs(819) <= '1';
    layer2_outputs(820) <= b and not a;
    layer2_outputs(821) <= not (a or b);
    layer2_outputs(822) <= '0';
    layer2_outputs(823) <= a and not b;
    layer2_outputs(824) <= '0';
    layer2_outputs(825) <= a or b;
    layer2_outputs(826) <= not a;
    layer2_outputs(827) <= b and not a;
    layer2_outputs(828) <= not b;
    layer2_outputs(829) <= a and not b;
    layer2_outputs(830) <= a;
    layer2_outputs(831) <= a;
    layer2_outputs(832) <= b;
    layer2_outputs(833) <= not (a xor b);
    layer2_outputs(834) <= not (a xor b);
    layer2_outputs(835) <= b;
    layer2_outputs(836) <= b;
    layer2_outputs(837) <= not a;
    layer2_outputs(838) <= b;
    layer2_outputs(839) <= '1';
    layer2_outputs(840) <= not a;
    layer2_outputs(841) <= not a or b;
    layer2_outputs(842) <= not (a and b);
    layer2_outputs(843) <= a or b;
    layer2_outputs(844) <= not b or a;
    layer2_outputs(845) <= a and not b;
    layer2_outputs(846) <= not b or a;
    layer2_outputs(847) <= not (a or b);
    layer2_outputs(848) <= not b;
    layer2_outputs(849) <= a and not b;
    layer2_outputs(850) <= not (a xor b);
    layer2_outputs(851) <= '0';
    layer2_outputs(852) <= '1';
    layer2_outputs(853) <= not b or a;
    layer2_outputs(854) <= b;
    layer2_outputs(855) <= a or b;
    layer2_outputs(856) <= not b;
    layer2_outputs(857) <= a or b;
    layer2_outputs(858) <= not b;
    layer2_outputs(859) <= not b;
    layer2_outputs(860) <= not (a and b);
    layer2_outputs(861) <= '0';
    layer2_outputs(862) <= a xor b;
    layer2_outputs(863) <= not b or a;
    layer2_outputs(864) <= not (a and b);
    layer2_outputs(865) <= '1';
    layer2_outputs(866) <= '1';
    layer2_outputs(867) <= b;
    layer2_outputs(868) <= a and not b;
    layer2_outputs(869) <= not a or b;
    layer2_outputs(870) <= a or b;
    layer2_outputs(871) <= not a;
    layer2_outputs(872) <= a xor b;
    layer2_outputs(873) <= '0';
    layer2_outputs(874) <= not b;
    layer2_outputs(875) <= a or b;
    layer2_outputs(876) <= not a;
    layer2_outputs(877) <= a or b;
    layer2_outputs(878) <= b and not a;
    layer2_outputs(879) <= a xor b;
    layer2_outputs(880) <= a or b;
    layer2_outputs(881) <= '0';
    layer2_outputs(882) <= not (a and b);
    layer2_outputs(883) <= a and b;
    layer2_outputs(884) <= a;
    layer2_outputs(885) <= '0';
    layer2_outputs(886) <= b and not a;
    layer2_outputs(887) <= not a or b;
    layer2_outputs(888) <= b;
    layer2_outputs(889) <= not (a or b);
    layer2_outputs(890) <= not b;
    layer2_outputs(891) <= '0';
    layer2_outputs(892) <= not (a and b);
    layer2_outputs(893) <= not b;
    layer2_outputs(894) <= a xor b;
    layer2_outputs(895) <= a;
    layer2_outputs(896) <= not (a and b);
    layer2_outputs(897) <= a and b;
    layer2_outputs(898) <= a;
    layer2_outputs(899) <= not a;
    layer2_outputs(900) <= not (a or b);
    layer2_outputs(901) <= not b;
    layer2_outputs(902) <= not b or a;
    layer2_outputs(903) <= a;
    layer2_outputs(904) <= a or b;
    layer2_outputs(905) <= b and not a;
    layer2_outputs(906) <= not b;
    layer2_outputs(907) <= b;
    layer2_outputs(908) <= b and not a;
    layer2_outputs(909) <= '0';
    layer2_outputs(910) <= not a;
    layer2_outputs(911) <= not (a and b);
    layer2_outputs(912) <= not (a and b);
    layer2_outputs(913) <= not (a or b);
    layer2_outputs(914) <= not (a xor b);
    layer2_outputs(915) <= a or b;
    layer2_outputs(916) <= not a;
    layer2_outputs(917) <= not b;
    layer2_outputs(918) <= a and not b;
    layer2_outputs(919) <= b;
    layer2_outputs(920) <= a and b;
    layer2_outputs(921) <= '0';
    layer2_outputs(922) <= not b;
    layer2_outputs(923) <= a or b;
    layer2_outputs(924) <= '1';
    layer2_outputs(925) <= '0';
    layer2_outputs(926) <= not (a or b);
    layer2_outputs(927) <= a and not b;
    layer2_outputs(928) <= a and b;
    layer2_outputs(929) <= not (a xor b);
    layer2_outputs(930) <= not (a or b);
    layer2_outputs(931) <= a and not b;
    layer2_outputs(932) <= a and not b;
    layer2_outputs(933) <= a or b;
    layer2_outputs(934) <= a;
    layer2_outputs(935) <= not a or b;
    layer2_outputs(936) <= a and not b;
    layer2_outputs(937) <= a and not b;
    layer2_outputs(938) <= not a or b;
    layer2_outputs(939) <= not a;
    layer2_outputs(940) <= not b or a;
    layer2_outputs(941) <= a and not b;
    layer2_outputs(942) <= not b;
    layer2_outputs(943) <= '1';
    layer2_outputs(944) <= not b;
    layer2_outputs(945) <= not a;
    layer2_outputs(946) <= not a;
    layer2_outputs(947) <= not b;
    layer2_outputs(948) <= a or b;
    layer2_outputs(949) <= not b;
    layer2_outputs(950) <= b and not a;
    layer2_outputs(951) <= a or b;
    layer2_outputs(952) <= '0';
    layer2_outputs(953) <= a and not b;
    layer2_outputs(954) <= a xor b;
    layer2_outputs(955) <= not (a and b);
    layer2_outputs(956) <= b;
    layer2_outputs(957) <= '0';
    layer2_outputs(958) <= not (a and b);
    layer2_outputs(959) <= not b;
    layer2_outputs(960) <= not (a and b);
    layer2_outputs(961) <= a and not b;
    layer2_outputs(962) <= b;
    layer2_outputs(963) <= not a;
    layer2_outputs(964) <= not a or b;
    layer2_outputs(965) <= not b;
    layer2_outputs(966) <= not b;
    layer2_outputs(967) <= '0';
    layer2_outputs(968) <= not b;
    layer2_outputs(969) <= not (a or b);
    layer2_outputs(970) <= a or b;
    layer2_outputs(971) <= a and not b;
    layer2_outputs(972) <= not a;
    layer2_outputs(973) <= not (a and b);
    layer2_outputs(974) <= not a;
    layer2_outputs(975) <= a;
    layer2_outputs(976) <= not (a and b);
    layer2_outputs(977) <= not (a and b);
    layer2_outputs(978) <= a and not b;
    layer2_outputs(979) <= not (a and b);
    layer2_outputs(980) <= '0';
    layer2_outputs(981) <= not b;
    layer2_outputs(982) <= b;
    layer2_outputs(983) <= not b or a;
    layer2_outputs(984) <= not b or a;
    layer2_outputs(985) <= '0';
    layer2_outputs(986) <= not a;
    layer2_outputs(987) <= not b;
    layer2_outputs(988) <= a or b;
    layer2_outputs(989) <= not b;
    layer2_outputs(990) <= '0';
    layer2_outputs(991) <= not (a or b);
    layer2_outputs(992) <= not (a xor b);
    layer2_outputs(993) <= b;
    layer2_outputs(994) <= not a;
    layer2_outputs(995) <= a;
    layer2_outputs(996) <= not b;
    layer2_outputs(997) <= not (a or b);
    layer2_outputs(998) <= not a;
    layer2_outputs(999) <= a or b;
    layer2_outputs(1000) <= not b;
    layer2_outputs(1001) <= '1';
    layer2_outputs(1002) <= b;
    layer2_outputs(1003) <= a or b;
    layer2_outputs(1004) <= not a;
    layer2_outputs(1005) <= not (a and b);
    layer2_outputs(1006) <= not b;
    layer2_outputs(1007) <= a;
    layer2_outputs(1008) <= a xor b;
    layer2_outputs(1009) <= not b;
    layer2_outputs(1010) <= not b or a;
    layer2_outputs(1011) <= '0';
    layer2_outputs(1012) <= not a;
    layer2_outputs(1013) <= not (a or b);
    layer2_outputs(1014) <= '0';
    layer2_outputs(1015) <= not b or a;
    layer2_outputs(1016) <= not b;
    layer2_outputs(1017) <= not b or a;
    layer2_outputs(1018) <= '1';
    layer2_outputs(1019) <= a or b;
    layer2_outputs(1020) <= not (a and b);
    layer2_outputs(1021) <= not (a or b);
    layer2_outputs(1022) <= not (a and b);
    layer2_outputs(1023) <= b and not a;
    layer2_outputs(1024) <= not a;
    layer2_outputs(1025) <= not a or b;
    layer2_outputs(1026) <= a or b;
    layer2_outputs(1027) <= not b or a;
    layer2_outputs(1028) <= b and not a;
    layer2_outputs(1029) <= not (a and b);
    layer2_outputs(1030) <= '1';
    layer2_outputs(1031) <= '1';
    layer2_outputs(1032) <= a and b;
    layer2_outputs(1033) <= a and b;
    layer2_outputs(1034) <= a;
    layer2_outputs(1035) <= not b or a;
    layer2_outputs(1036) <= '0';
    layer2_outputs(1037) <= not a or b;
    layer2_outputs(1038) <= not a;
    layer2_outputs(1039) <= a xor b;
    layer2_outputs(1040) <= a and b;
    layer2_outputs(1041) <= not (a or b);
    layer2_outputs(1042) <= not b;
    layer2_outputs(1043) <= '1';
    layer2_outputs(1044) <= not (a xor b);
    layer2_outputs(1045) <= b;
    layer2_outputs(1046) <= not (a or b);
    layer2_outputs(1047) <= b;
    layer2_outputs(1048) <= a xor b;
    layer2_outputs(1049) <= not (a or b);
    layer2_outputs(1050) <= '0';
    layer2_outputs(1051) <= '1';
    layer2_outputs(1052) <= b and not a;
    layer2_outputs(1053) <= a or b;
    layer2_outputs(1054) <= b;
    layer2_outputs(1055) <= not b or a;
    layer2_outputs(1056) <= a and not b;
    layer2_outputs(1057) <= not b or a;
    layer2_outputs(1058) <= a or b;
    layer2_outputs(1059) <= not (a and b);
    layer2_outputs(1060) <= not (a and b);
    layer2_outputs(1061) <= not b;
    layer2_outputs(1062) <= b and not a;
    layer2_outputs(1063) <= not b;
    layer2_outputs(1064) <= b;
    layer2_outputs(1065) <= a or b;
    layer2_outputs(1066) <= not b;
    layer2_outputs(1067) <= '0';
    layer2_outputs(1068) <= b and not a;
    layer2_outputs(1069) <= not (a xor b);
    layer2_outputs(1070) <= not (a and b);
    layer2_outputs(1071) <= not b or a;
    layer2_outputs(1072) <= not a or b;
    layer2_outputs(1073) <= not (a and b);
    layer2_outputs(1074) <= '0';
    layer2_outputs(1075) <= '1';
    layer2_outputs(1076) <= not b or a;
    layer2_outputs(1077) <= a and b;
    layer2_outputs(1078) <= not a;
    layer2_outputs(1079) <= a and b;
    layer2_outputs(1080) <= not (a or b);
    layer2_outputs(1081) <= not b;
    layer2_outputs(1082) <= not (a or b);
    layer2_outputs(1083) <= b;
    layer2_outputs(1084) <= not (a or b);
    layer2_outputs(1085) <= a and not b;
    layer2_outputs(1086) <= a and b;
    layer2_outputs(1087) <= not (a or b);
    layer2_outputs(1088) <= not a;
    layer2_outputs(1089) <= a;
    layer2_outputs(1090) <= b and not a;
    layer2_outputs(1091) <= not b or a;
    layer2_outputs(1092) <= not (a xor b);
    layer2_outputs(1093) <= not b or a;
    layer2_outputs(1094) <= not b or a;
    layer2_outputs(1095) <= not a or b;
    layer2_outputs(1096) <= not a;
    layer2_outputs(1097) <= a;
    layer2_outputs(1098) <= not (a and b);
    layer2_outputs(1099) <= b;
    layer2_outputs(1100) <= not b or a;
    layer2_outputs(1101) <= not (a or b);
    layer2_outputs(1102) <= not (a xor b);
    layer2_outputs(1103) <= a;
    layer2_outputs(1104) <= a or b;
    layer2_outputs(1105) <= not a;
    layer2_outputs(1106) <= a or b;
    layer2_outputs(1107) <= a and not b;
    layer2_outputs(1108) <= a;
    layer2_outputs(1109) <= not a;
    layer2_outputs(1110) <= not a or b;
    layer2_outputs(1111) <= a and b;
    layer2_outputs(1112) <= a and not b;
    layer2_outputs(1113) <= b;
    layer2_outputs(1114) <= a or b;
    layer2_outputs(1115) <= a;
    layer2_outputs(1116) <= '1';
    layer2_outputs(1117) <= a and not b;
    layer2_outputs(1118) <= not b or a;
    layer2_outputs(1119) <= a and b;
    layer2_outputs(1120) <= a and not b;
    layer2_outputs(1121) <= a;
    layer2_outputs(1122) <= a and b;
    layer2_outputs(1123) <= a;
    layer2_outputs(1124) <= a and not b;
    layer2_outputs(1125) <= not (a and b);
    layer2_outputs(1126) <= not b;
    layer2_outputs(1127) <= a;
    layer2_outputs(1128) <= b and not a;
    layer2_outputs(1129) <= not (a or b);
    layer2_outputs(1130) <= not (a xor b);
    layer2_outputs(1131) <= not (a and b);
    layer2_outputs(1132) <= b and not a;
    layer2_outputs(1133) <= not (a and b);
    layer2_outputs(1134) <= not (a xor b);
    layer2_outputs(1135) <= not (a or b);
    layer2_outputs(1136) <= b and not a;
    layer2_outputs(1137) <= not a or b;
    layer2_outputs(1138) <= a and not b;
    layer2_outputs(1139) <= a xor b;
    layer2_outputs(1140) <= a and not b;
    layer2_outputs(1141) <= a and not b;
    layer2_outputs(1142) <= '0';
    layer2_outputs(1143) <= '0';
    layer2_outputs(1144) <= b;
    layer2_outputs(1145) <= not a or b;
    layer2_outputs(1146) <= a xor b;
    layer2_outputs(1147) <= b and not a;
    layer2_outputs(1148) <= not (a or b);
    layer2_outputs(1149) <= not (a and b);
    layer2_outputs(1150) <= not a or b;
    layer2_outputs(1151) <= not b or a;
    layer2_outputs(1152) <= not b;
    layer2_outputs(1153) <= not a;
    layer2_outputs(1154) <= not b;
    layer2_outputs(1155) <= not (a or b);
    layer2_outputs(1156) <= not a;
    layer2_outputs(1157) <= b and not a;
    layer2_outputs(1158) <= b;
    layer2_outputs(1159) <= '0';
    layer2_outputs(1160) <= '1';
    layer2_outputs(1161) <= b;
    layer2_outputs(1162) <= not b;
    layer2_outputs(1163) <= not (a and b);
    layer2_outputs(1164) <= not (a xor b);
    layer2_outputs(1165) <= b and not a;
    layer2_outputs(1166) <= b and not a;
    layer2_outputs(1167) <= not a;
    layer2_outputs(1168) <= '0';
    layer2_outputs(1169) <= a and not b;
    layer2_outputs(1170) <= not a;
    layer2_outputs(1171) <= not a or b;
    layer2_outputs(1172) <= a or b;
    layer2_outputs(1173) <= not a or b;
    layer2_outputs(1174) <= b;
    layer2_outputs(1175) <= not a or b;
    layer2_outputs(1176) <= b;
    layer2_outputs(1177) <= not b;
    layer2_outputs(1178) <= b and not a;
    layer2_outputs(1179) <= a;
    layer2_outputs(1180) <= not (a and b);
    layer2_outputs(1181) <= b;
    layer2_outputs(1182) <= not b or a;
    layer2_outputs(1183) <= not a or b;
    layer2_outputs(1184) <= '0';
    layer2_outputs(1185) <= a;
    layer2_outputs(1186) <= a or b;
    layer2_outputs(1187) <= not a;
    layer2_outputs(1188) <= a and b;
    layer2_outputs(1189) <= b;
    layer2_outputs(1190) <= not (a and b);
    layer2_outputs(1191) <= not b or a;
    layer2_outputs(1192) <= b;
    layer2_outputs(1193) <= not b;
    layer2_outputs(1194) <= a and b;
    layer2_outputs(1195) <= not b;
    layer2_outputs(1196) <= '1';
    layer2_outputs(1197) <= a or b;
    layer2_outputs(1198) <= '1';
    layer2_outputs(1199) <= not b or a;
    layer2_outputs(1200) <= not (a and b);
    layer2_outputs(1201) <= a;
    layer2_outputs(1202) <= a or b;
    layer2_outputs(1203) <= '0';
    layer2_outputs(1204) <= not (a and b);
    layer2_outputs(1205) <= not b;
    layer2_outputs(1206) <= '1';
    layer2_outputs(1207) <= not a or b;
    layer2_outputs(1208) <= '0';
    layer2_outputs(1209) <= '0';
    layer2_outputs(1210) <= a and b;
    layer2_outputs(1211) <= a or b;
    layer2_outputs(1212) <= b;
    layer2_outputs(1213) <= a and not b;
    layer2_outputs(1214) <= not a;
    layer2_outputs(1215) <= a or b;
    layer2_outputs(1216) <= a;
    layer2_outputs(1217) <= not a;
    layer2_outputs(1218) <= a and b;
    layer2_outputs(1219) <= b and not a;
    layer2_outputs(1220) <= b;
    layer2_outputs(1221) <= not a or b;
    layer2_outputs(1222) <= not (a or b);
    layer2_outputs(1223) <= a and b;
    layer2_outputs(1224) <= '0';
    layer2_outputs(1225) <= not a or b;
    layer2_outputs(1226) <= not b or a;
    layer2_outputs(1227) <= a;
    layer2_outputs(1228) <= '1';
    layer2_outputs(1229) <= not a or b;
    layer2_outputs(1230) <= not (a and b);
    layer2_outputs(1231) <= not a;
    layer2_outputs(1232) <= a;
    layer2_outputs(1233) <= b;
    layer2_outputs(1234) <= a and not b;
    layer2_outputs(1235) <= not (a and b);
    layer2_outputs(1236) <= b and not a;
    layer2_outputs(1237) <= not (a xor b);
    layer2_outputs(1238) <= '0';
    layer2_outputs(1239) <= not a;
    layer2_outputs(1240) <= b and not a;
    layer2_outputs(1241) <= '1';
    layer2_outputs(1242) <= '1';
    layer2_outputs(1243) <= a and b;
    layer2_outputs(1244) <= not a or b;
    layer2_outputs(1245) <= b and not a;
    layer2_outputs(1246) <= not (a xor b);
    layer2_outputs(1247) <= '0';
    layer2_outputs(1248) <= a xor b;
    layer2_outputs(1249) <= a and b;
    layer2_outputs(1250) <= not (a or b);
    layer2_outputs(1251) <= not b or a;
    layer2_outputs(1252) <= not a;
    layer2_outputs(1253) <= not a or b;
    layer2_outputs(1254) <= not b or a;
    layer2_outputs(1255) <= a and b;
    layer2_outputs(1256) <= not b or a;
    layer2_outputs(1257) <= not a or b;
    layer2_outputs(1258) <= not b or a;
    layer2_outputs(1259) <= a;
    layer2_outputs(1260) <= a and b;
    layer2_outputs(1261) <= a;
    layer2_outputs(1262) <= not a;
    layer2_outputs(1263) <= '1';
    layer2_outputs(1264) <= not b;
    layer2_outputs(1265) <= not (a and b);
    layer2_outputs(1266) <= a xor b;
    layer2_outputs(1267) <= not a;
    layer2_outputs(1268) <= not (a or b);
    layer2_outputs(1269) <= not (a and b);
    layer2_outputs(1270) <= a;
    layer2_outputs(1271) <= b;
    layer2_outputs(1272) <= not b or a;
    layer2_outputs(1273) <= not a;
    layer2_outputs(1274) <= not a;
    layer2_outputs(1275) <= not b;
    layer2_outputs(1276) <= not (a xor b);
    layer2_outputs(1277) <= b;
    layer2_outputs(1278) <= not (a or b);
    layer2_outputs(1279) <= '0';
    layer2_outputs(1280) <= a;
    layer2_outputs(1281) <= '0';
    layer2_outputs(1282) <= b and not a;
    layer2_outputs(1283) <= b;
    layer2_outputs(1284) <= not a;
    layer2_outputs(1285) <= not (a and b);
    layer2_outputs(1286) <= a or b;
    layer2_outputs(1287) <= a or b;
    layer2_outputs(1288) <= a and b;
    layer2_outputs(1289) <= a or b;
    layer2_outputs(1290) <= a;
    layer2_outputs(1291) <= b;
    layer2_outputs(1292) <= a and b;
    layer2_outputs(1293) <= '1';
    layer2_outputs(1294) <= b;
    layer2_outputs(1295) <= a;
    layer2_outputs(1296) <= not (a xor b);
    layer2_outputs(1297) <= a or b;
    layer2_outputs(1298) <= '1';
    layer2_outputs(1299) <= a;
    layer2_outputs(1300) <= not (a or b);
    layer2_outputs(1301) <= a;
    layer2_outputs(1302) <= not (a and b);
    layer2_outputs(1303) <= b;
    layer2_outputs(1304) <= not a or b;
    layer2_outputs(1305) <= a;
    layer2_outputs(1306) <= not a;
    layer2_outputs(1307) <= b;
    layer2_outputs(1308) <= a or b;
    layer2_outputs(1309) <= '0';
    layer2_outputs(1310) <= a and b;
    layer2_outputs(1311) <= b and not a;
    layer2_outputs(1312) <= not b or a;
    layer2_outputs(1313) <= not (a xor b);
    layer2_outputs(1314) <= not b or a;
    layer2_outputs(1315) <= a and b;
    layer2_outputs(1316) <= a and not b;
    layer2_outputs(1317) <= not a or b;
    layer2_outputs(1318) <= a xor b;
    layer2_outputs(1319) <= not b;
    layer2_outputs(1320) <= a and b;
    layer2_outputs(1321) <= not (a and b);
    layer2_outputs(1322) <= not a;
    layer2_outputs(1323) <= not b;
    layer2_outputs(1324) <= not (a or b);
    layer2_outputs(1325) <= not b;
    layer2_outputs(1326) <= not (a and b);
    layer2_outputs(1327) <= not a;
    layer2_outputs(1328) <= b;
    layer2_outputs(1329) <= a;
    layer2_outputs(1330) <= b and not a;
    layer2_outputs(1331) <= b;
    layer2_outputs(1332) <= not a;
    layer2_outputs(1333) <= a and b;
    layer2_outputs(1334) <= a;
    layer2_outputs(1335) <= not a or b;
    layer2_outputs(1336) <= '0';
    layer2_outputs(1337) <= a or b;
    layer2_outputs(1338) <= not a or b;
    layer2_outputs(1339) <= a;
    layer2_outputs(1340) <= a and not b;
    layer2_outputs(1341) <= a and b;
    layer2_outputs(1342) <= a and b;
    layer2_outputs(1343) <= '0';
    layer2_outputs(1344) <= b;
    layer2_outputs(1345) <= b and not a;
    layer2_outputs(1346) <= b and not a;
    layer2_outputs(1347) <= a or b;
    layer2_outputs(1348) <= not (a and b);
    layer2_outputs(1349) <= not b or a;
    layer2_outputs(1350) <= b;
    layer2_outputs(1351) <= not b or a;
    layer2_outputs(1352) <= not b;
    layer2_outputs(1353) <= a;
    layer2_outputs(1354) <= not a;
    layer2_outputs(1355) <= not b or a;
    layer2_outputs(1356) <= b;
    layer2_outputs(1357) <= b;
    layer2_outputs(1358) <= not (a or b);
    layer2_outputs(1359) <= not (a or b);
    layer2_outputs(1360) <= not (a or b);
    layer2_outputs(1361) <= a;
    layer2_outputs(1362) <= '0';
    layer2_outputs(1363) <= not b or a;
    layer2_outputs(1364) <= b;
    layer2_outputs(1365) <= not a or b;
    layer2_outputs(1366) <= not (a or b);
    layer2_outputs(1367) <= '0';
    layer2_outputs(1368) <= '1';
    layer2_outputs(1369) <= a and not b;
    layer2_outputs(1370) <= not b or a;
    layer2_outputs(1371) <= not (a or b);
    layer2_outputs(1372) <= a;
    layer2_outputs(1373) <= '0';
    layer2_outputs(1374) <= not (a or b);
    layer2_outputs(1375) <= not b or a;
    layer2_outputs(1376) <= a;
    layer2_outputs(1377) <= '0';
    layer2_outputs(1378) <= b;
    layer2_outputs(1379) <= a;
    layer2_outputs(1380) <= a xor b;
    layer2_outputs(1381) <= not a or b;
    layer2_outputs(1382) <= not a;
    layer2_outputs(1383) <= b and not a;
    layer2_outputs(1384) <= not b or a;
    layer2_outputs(1385) <= b and not a;
    layer2_outputs(1386) <= '0';
    layer2_outputs(1387) <= not a;
    layer2_outputs(1388) <= a and not b;
    layer2_outputs(1389) <= not b or a;
    layer2_outputs(1390) <= not (a and b);
    layer2_outputs(1391) <= a;
    layer2_outputs(1392) <= not b;
    layer2_outputs(1393) <= not (a or b);
    layer2_outputs(1394) <= not a or b;
    layer2_outputs(1395) <= a and b;
    layer2_outputs(1396) <= '1';
    layer2_outputs(1397) <= not b;
    layer2_outputs(1398) <= not (a xor b);
    layer2_outputs(1399) <= b;
    layer2_outputs(1400) <= not b;
    layer2_outputs(1401) <= a and b;
    layer2_outputs(1402) <= a and not b;
    layer2_outputs(1403) <= not b or a;
    layer2_outputs(1404) <= b;
    layer2_outputs(1405) <= not a;
    layer2_outputs(1406) <= a;
    layer2_outputs(1407) <= a and b;
    layer2_outputs(1408) <= not b or a;
    layer2_outputs(1409) <= not a;
    layer2_outputs(1410) <= not b or a;
    layer2_outputs(1411) <= a;
    layer2_outputs(1412) <= not a or b;
    layer2_outputs(1413) <= not (a xor b);
    layer2_outputs(1414) <= a or b;
    layer2_outputs(1415) <= a or b;
    layer2_outputs(1416) <= a;
    layer2_outputs(1417) <= not a or b;
    layer2_outputs(1418) <= b and not a;
    layer2_outputs(1419) <= not a;
    layer2_outputs(1420) <= not a;
    layer2_outputs(1421) <= not a or b;
    layer2_outputs(1422) <= a;
    layer2_outputs(1423) <= a;
    layer2_outputs(1424) <= b and not a;
    layer2_outputs(1425) <= b and not a;
    layer2_outputs(1426) <= b;
    layer2_outputs(1427) <= '0';
    layer2_outputs(1428) <= a and not b;
    layer2_outputs(1429) <= not b or a;
    layer2_outputs(1430) <= b and not a;
    layer2_outputs(1431) <= a or b;
    layer2_outputs(1432) <= not (a and b);
    layer2_outputs(1433) <= b and not a;
    layer2_outputs(1434) <= not (a and b);
    layer2_outputs(1435) <= not b or a;
    layer2_outputs(1436) <= a or b;
    layer2_outputs(1437) <= '1';
    layer2_outputs(1438) <= b and not a;
    layer2_outputs(1439) <= a and not b;
    layer2_outputs(1440) <= b;
    layer2_outputs(1441) <= not (a xor b);
    layer2_outputs(1442) <= not (a and b);
    layer2_outputs(1443) <= a and not b;
    layer2_outputs(1444) <= not (a and b);
    layer2_outputs(1445) <= b;
    layer2_outputs(1446) <= not a;
    layer2_outputs(1447) <= a and b;
    layer2_outputs(1448) <= '1';
    layer2_outputs(1449) <= not a;
    layer2_outputs(1450) <= a xor b;
    layer2_outputs(1451) <= not (a and b);
    layer2_outputs(1452) <= b;
    layer2_outputs(1453) <= b and not a;
    layer2_outputs(1454) <= b and not a;
    layer2_outputs(1455) <= b;
    layer2_outputs(1456) <= a and not b;
    layer2_outputs(1457) <= not (a and b);
    layer2_outputs(1458) <= not a or b;
    layer2_outputs(1459) <= a and not b;
    layer2_outputs(1460) <= b and not a;
    layer2_outputs(1461) <= a or b;
    layer2_outputs(1462) <= not a;
    layer2_outputs(1463) <= a or b;
    layer2_outputs(1464) <= b and not a;
    layer2_outputs(1465) <= b;
    layer2_outputs(1466) <= a or b;
    layer2_outputs(1467) <= a;
    layer2_outputs(1468) <= b;
    layer2_outputs(1469) <= b;
    layer2_outputs(1470) <= not (a xor b);
    layer2_outputs(1471) <= b and not a;
    layer2_outputs(1472) <= not a;
    layer2_outputs(1473) <= '1';
    layer2_outputs(1474) <= not (a or b);
    layer2_outputs(1475) <= not b or a;
    layer2_outputs(1476) <= b and not a;
    layer2_outputs(1477) <= b;
    layer2_outputs(1478) <= not (a and b);
    layer2_outputs(1479) <= not (a and b);
    layer2_outputs(1480) <= not a or b;
    layer2_outputs(1481) <= b;
    layer2_outputs(1482) <= not b;
    layer2_outputs(1483) <= '1';
    layer2_outputs(1484) <= b and not a;
    layer2_outputs(1485) <= not b or a;
    layer2_outputs(1486) <= b;
    layer2_outputs(1487) <= not (a and b);
    layer2_outputs(1488) <= a and b;
    layer2_outputs(1489) <= '0';
    layer2_outputs(1490) <= not a;
    layer2_outputs(1491) <= a and b;
    layer2_outputs(1492) <= a and b;
    layer2_outputs(1493) <= not a or b;
    layer2_outputs(1494) <= not (a or b);
    layer2_outputs(1495) <= not (a xor b);
    layer2_outputs(1496) <= not b;
    layer2_outputs(1497) <= '0';
    layer2_outputs(1498) <= a;
    layer2_outputs(1499) <= not a or b;
    layer2_outputs(1500) <= a and not b;
    layer2_outputs(1501) <= a or b;
    layer2_outputs(1502) <= not (a or b);
    layer2_outputs(1503) <= not (a xor b);
    layer2_outputs(1504) <= a xor b;
    layer2_outputs(1505) <= not (a or b);
    layer2_outputs(1506) <= a and not b;
    layer2_outputs(1507) <= not a;
    layer2_outputs(1508) <= b;
    layer2_outputs(1509) <= not (a and b);
    layer2_outputs(1510) <= b and not a;
    layer2_outputs(1511) <= '1';
    layer2_outputs(1512) <= not b or a;
    layer2_outputs(1513) <= a or b;
    layer2_outputs(1514) <= not (a and b);
    layer2_outputs(1515) <= not a or b;
    layer2_outputs(1516) <= '0';
    layer2_outputs(1517) <= b;
    layer2_outputs(1518) <= not (a and b);
    layer2_outputs(1519) <= not a;
    layer2_outputs(1520) <= not (a or b);
    layer2_outputs(1521) <= not (a and b);
    layer2_outputs(1522) <= not (a and b);
    layer2_outputs(1523) <= b and not a;
    layer2_outputs(1524) <= a and b;
    layer2_outputs(1525) <= b;
    layer2_outputs(1526) <= a;
    layer2_outputs(1527) <= a or b;
    layer2_outputs(1528) <= '1';
    layer2_outputs(1529) <= a xor b;
    layer2_outputs(1530) <= '1';
    layer2_outputs(1531) <= '1';
    layer2_outputs(1532) <= not a;
    layer2_outputs(1533) <= not a or b;
    layer2_outputs(1534) <= b;
    layer2_outputs(1535) <= not b or a;
    layer2_outputs(1536) <= '0';
    layer2_outputs(1537) <= a or b;
    layer2_outputs(1538) <= a and b;
    layer2_outputs(1539) <= a;
    layer2_outputs(1540) <= b;
    layer2_outputs(1541) <= not a or b;
    layer2_outputs(1542) <= not b or a;
    layer2_outputs(1543) <= a;
    layer2_outputs(1544) <= b;
    layer2_outputs(1545) <= not (a and b);
    layer2_outputs(1546) <= not b or a;
    layer2_outputs(1547) <= b;
    layer2_outputs(1548) <= a or b;
    layer2_outputs(1549) <= b;
    layer2_outputs(1550) <= a and b;
    layer2_outputs(1551) <= b;
    layer2_outputs(1552) <= a or b;
    layer2_outputs(1553) <= b and not a;
    layer2_outputs(1554) <= not b;
    layer2_outputs(1555) <= '1';
    layer2_outputs(1556) <= not (a and b);
    layer2_outputs(1557) <= not a or b;
    layer2_outputs(1558) <= not a or b;
    layer2_outputs(1559) <= b and not a;
    layer2_outputs(1560) <= not a;
    layer2_outputs(1561) <= a and not b;
    layer2_outputs(1562) <= a and b;
    layer2_outputs(1563) <= a;
    layer2_outputs(1564) <= a or b;
    layer2_outputs(1565) <= b;
    layer2_outputs(1566) <= a;
    layer2_outputs(1567) <= b and not a;
    layer2_outputs(1568) <= not (a or b);
    layer2_outputs(1569) <= not (a and b);
    layer2_outputs(1570) <= a and b;
    layer2_outputs(1571) <= not (a or b);
    layer2_outputs(1572) <= not (a and b);
    layer2_outputs(1573) <= not b or a;
    layer2_outputs(1574) <= not b;
    layer2_outputs(1575) <= '1';
    layer2_outputs(1576) <= '1';
    layer2_outputs(1577) <= b;
    layer2_outputs(1578) <= a or b;
    layer2_outputs(1579) <= not a or b;
    layer2_outputs(1580) <= not a;
    layer2_outputs(1581) <= not b;
    layer2_outputs(1582) <= a;
    layer2_outputs(1583) <= not a or b;
    layer2_outputs(1584) <= not (a and b);
    layer2_outputs(1585) <= not b;
    layer2_outputs(1586) <= not a or b;
    layer2_outputs(1587) <= not (a or b);
    layer2_outputs(1588) <= a;
    layer2_outputs(1589) <= a xor b;
    layer2_outputs(1590) <= a or b;
    layer2_outputs(1591) <= b and not a;
    layer2_outputs(1592) <= b and not a;
    layer2_outputs(1593) <= not a;
    layer2_outputs(1594) <= not b;
    layer2_outputs(1595) <= a or b;
    layer2_outputs(1596) <= a and not b;
    layer2_outputs(1597) <= b;
    layer2_outputs(1598) <= not a;
    layer2_outputs(1599) <= b;
    layer2_outputs(1600) <= not a;
    layer2_outputs(1601) <= b and not a;
    layer2_outputs(1602) <= b and not a;
    layer2_outputs(1603) <= a or b;
    layer2_outputs(1604) <= not (a and b);
    layer2_outputs(1605) <= b;
    layer2_outputs(1606) <= a xor b;
    layer2_outputs(1607) <= b;
    layer2_outputs(1608) <= not a or b;
    layer2_outputs(1609) <= '0';
    layer2_outputs(1610) <= '1';
    layer2_outputs(1611) <= not b;
    layer2_outputs(1612) <= a and not b;
    layer2_outputs(1613) <= a or b;
    layer2_outputs(1614) <= a and not b;
    layer2_outputs(1615) <= a;
    layer2_outputs(1616) <= b;
    layer2_outputs(1617) <= b and not a;
    layer2_outputs(1618) <= not a or b;
    layer2_outputs(1619) <= not a or b;
    layer2_outputs(1620) <= a or b;
    layer2_outputs(1621) <= b and not a;
    layer2_outputs(1622) <= '1';
    layer2_outputs(1623) <= not a;
    layer2_outputs(1624) <= b;
    layer2_outputs(1625) <= '1';
    layer2_outputs(1626) <= not a;
    layer2_outputs(1627) <= not a or b;
    layer2_outputs(1628) <= a xor b;
    layer2_outputs(1629) <= not (a and b);
    layer2_outputs(1630) <= a or b;
    layer2_outputs(1631) <= b and not a;
    layer2_outputs(1632) <= not b or a;
    layer2_outputs(1633) <= a and b;
    layer2_outputs(1634) <= not b;
    layer2_outputs(1635) <= not b or a;
    layer2_outputs(1636) <= a and not b;
    layer2_outputs(1637) <= a and not b;
    layer2_outputs(1638) <= b;
    layer2_outputs(1639) <= a or b;
    layer2_outputs(1640) <= not a;
    layer2_outputs(1641) <= b;
    layer2_outputs(1642) <= not (a or b);
    layer2_outputs(1643) <= a;
    layer2_outputs(1644) <= '0';
    layer2_outputs(1645) <= a or b;
    layer2_outputs(1646) <= not (a xor b);
    layer2_outputs(1647) <= a;
    layer2_outputs(1648) <= b;
    layer2_outputs(1649) <= a;
    layer2_outputs(1650) <= b;
    layer2_outputs(1651) <= a;
    layer2_outputs(1652) <= a;
    layer2_outputs(1653) <= a or b;
    layer2_outputs(1654) <= not a;
    layer2_outputs(1655) <= not b;
    layer2_outputs(1656) <= b;
    layer2_outputs(1657) <= a and b;
    layer2_outputs(1658) <= not (a and b);
    layer2_outputs(1659) <= a;
    layer2_outputs(1660) <= not b;
    layer2_outputs(1661) <= not a;
    layer2_outputs(1662) <= b;
    layer2_outputs(1663) <= not a;
    layer2_outputs(1664) <= not (a xor b);
    layer2_outputs(1665) <= not b;
    layer2_outputs(1666) <= b and not a;
    layer2_outputs(1667) <= not b;
    layer2_outputs(1668) <= not b or a;
    layer2_outputs(1669) <= a and b;
    layer2_outputs(1670) <= not (a or b);
    layer2_outputs(1671) <= a;
    layer2_outputs(1672) <= not a;
    layer2_outputs(1673) <= not b or a;
    layer2_outputs(1674) <= not b or a;
    layer2_outputs(1675) <= not a or b;
    layer2_outputs(1676) <= b and not a;
    layer2_outputs(1677) <= not a;
    layer2_outputs(1678) <= a xor b;
    layer2_outputs(1679) <= a;
    layer2_outputs(1680) <= a xor b;
    layer2_outputs(1681) <= not (a and b);
    layer2_outputs(1682) <= not a or b;
    layer2_outputs(1683) <= a;
    layer2_outputs(1684) <= a;
    layer2_outputs(1685) <= a or b;
    layer2_outputs(1686) <= not b;
    layer2_outputs(1687) <= not a;
    layer2_outputs(1688) <= a and b;
    layer2_outputs(1689) <= '0';
    layer2_outputs(1690) <= a xor b;
    layer2_outputs(1691) <= not b or a;
    layer2_outputs(1692) <= not b;
    layer2_outputs(1693) <= a;
    layer2_outputs(1694) <= a and b;
    layer2_outputs(1695) <= a;
    layer2_outputs(1696) <= not b;
    layer2_outputs(1697) <= not (a and b);
    layer2_outputs(1698) <= not (a and b);
    layer2_outputs(1699) <= a;
    layer2_outputs(1700) <= b and not a;
    layer2_outputs(1701) <= a and b;
    layer2_outputs(1702) <= not a;
    layer2_outputs(1703) <= b and not a;
    layer2_outputs(1704) <= a and b;
    layer2_outputs(1705) <= not b or a;
    layer2_outputs(1706) <= not b;
    layer2_outputs(1707) <= not (a and b);
    layer2_outputs(1708) <= a xor b;
    layer2_outputs(1709) <= not a;
    layer2_outputs(1710) <= a and b;
    layer2_outputs(1711) <= b and not a;
    layer2_outputs(1712) <= not a;
    layer2_outputs(1713) <= not a or b;
    layer2_outputs(1714) <= '0';
    layer2_outputs(1715) <= not b;
    layer2_outputs(1716) <= not b;
    layer2_outputs(1717) <= not (a xor b);
    layer2_outputs(1718) <= not b or a;
    layer2_outputs(1719) <= a or b;
    layer2_outputs(1720) <= not (a or b);
    layer2_outputs(1721) <= not b or a;
    layer2_outputs(1722) <= not (a or b);
    layer2_outputs(1723) <= not a or b;
    layer2_outputs(1724) <= not (a xor b);
    layer2_outputs(1725) <= a and b;
    layer2_outputs(1726) <= not (a xor b);
    layer2_outputs(1727) <= a and not b;
    layer2_outputs(1728) <= a;
    layer2_outputs(1729) <= not b;
    layer2_outputs(1730) <= not (a xor b);
    layer2_outputs(1731) <= not b;
    layer2_outputs(1732) <= not b;
    layer2_outputs(1733) <= not a;
    layer2_outputs(1734) <= not b;
    layer2_outputs(1735) <= a and not b;
    layer2_outputs(1736) <= not (a or b);
    layer2_outputs(1737) <= b;
    layer2_outputs(1738) <= '1';
    layer2_outputs(1739) <= not a or b;
    layer2_outputs(1740) <= '0';
    layer2_outputs(1741) <= a;
    layer2_outputs(1742) <= not (a or b);
    layer2_outputs(1743) <= a and b;
    layer2_outputs(1744) <= '1';
    layer2_outputs(1745) <= a xor b;
    layer2_outputs(1746) <= a;
    layer2_outputs(1747) <= not (a or b);
    layer2_outputs(1748) <= not (a or b);
    layer2_outputs(1749) <= a or b;
    layer2_outputs(1750) <= not a;
    layer2_outputs(1751) <= not (a and b);
    layer2_outputs(1752) <= a;
    layer2_outputs(1753) <= not b or a;
    layer2_outputs(1754) <= '1';
    layer2_outputs(1755) <= a and not b;
    layer2_outputs(1756) <= not b;
    layer2_outputs(1757) <= b;
    layer2_outputs(1758) <= '0';
    layer2_outputs(1759) <= not a or b;
    layer2_outputs(1760) <= not a;
    layer2_outputs(1761) <= b and not a;
    layer2_outputs(1762) <= not b or a;
    layer2_outputs(1763) <= a or b;
    layer2_outputs(1764) <= not (a and b);
    layer2_outputs(1765) <= not a;
    layer2_outputs(1766) <= a and not b;
    layer2_outputs(1767) <= a and not b;
    layer2_outputs(1768) <= b and not a;
    layer2_outputs(1769) <= not b or a;
    layer2_outputs(1770) <= a;
    layer2_outputs(1771) <= not a or b;
    layer2_outputs(1772) <= not (a or b);
    layer2_outputs(1773) <= a or b;
    layer2_outputs(1774) <= a and b;
    layer2_outputs(1775) <= not a;
    layer2_outputs(1776) <= a or b;
    layer2_outputs(1777) <= a or b;
    layer2_outputs(1778) <= b;
    layer2_outputs(1779) <= b;
    layer2_outputs(1780) <= not b or a;
    layer2_outputs(1781) <= not (a xor b);
    layer2_outputs(1782) <= not b or a;
    layer2_outputs(1783) <= not (a xor b);
    layer2_outputs(1784) <= a;
    layer2_outputs(1785) <= not a or b;
    layer2_outputs(1786) <= '1';
    layer2_outputs(1787) <= b and not a;
    layer2_outputs(1788) <= not (a xor b);
    layer2_outputs(1789) <= not (a and b);
    layer2_outputs(1790) <= b;
    layer2_outputs(1791) <= not b;
    layer2_outputs(1792) <= a and b;
    layer2_outputs(1793) <= '0';
    layer2_outputs(1794) <= b;
    layer2_outputs(1795) <= b and not a;
    layer2_outputs(1796) <= '0';
    layer2_outputs(1797) <= '1';
    layer2_outputs(1798) <= b;
    layer2_outputs(1799) <= b;
    layer2_outputs(1800) <= not (a xor b);
    layer2_outputs(1801) <= not a;
    layer2_outputs(1802) <= '1';
    layer2_outputs(1803) <= a and not b;
    layer2_outputs(1804) <= not a or b;
    layer2_outputs(1805) <= not b;
    layer2_outputs(1806) <= '1';
    layer2_outputs(1807) <= '0';
    layer2_outputs(1808) <= not a or b;
    layer2_outputs(1809) <= not (a and b);
    layer2_outputs(1810) <= '1';
    layer2_outputs(1811) <= a;
    layer2_outputs(1812) <= not a or b;
    layer2_outputs(1813) <= b;
    layer2_outputs(1814) <= a;
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= not a;
    layer2_outputs(1817) <= not (a xor b);
    layer2_outputs(1818) <= not a;
    layer2_outputs(1819) <= not (a or b);
    layer2_outputs(1820) <= not (a or b);
    layer2_outputs(1821) <= a and b;
    layer2_outputs(1822) <= not a or b;
    layer2_outputs(1823) <= not a;
    layer2_outputs(1824) <= not b;
    layer2_outputs(1825) <= not b;
    layer2_outputs(1826) <= a and not b;
    layer2_outputs(1827) <= a or b;
    layer2_outputs(1828) <= not (a or b);
    layer2_outputs(1829) <= not a or b;
    layer2_outputs(1830) <= b;
    layer2_outputs(1831) <= b;
    layer2_outputs(1832) <= a xor b;
    layer2_outputs(1833) <= b and not a;
    layer2_outputs(1834) <= a or b;
    layer2_outputs(1835) <= not (a xor b);
    layer2_outputs(1836) <= a and b;
    layer2_outputs(1837) <= not (a and b);
    layer2_outputs(1838) <= not b;
    layer2_outputs(1839) <= a;
    layer2_outputs(1840) <= not (a xor b);
    layer2_outputs(1841) <= a and not b;
    layer2_outputs(1842) <= a and not b;
    layer2_outputs(1843) <= not (a or b);
    layer2_outputs(1844) <= not a or b;
    layer2_outputs(1845) <= not (a or b);
    layer2_outputs(1846) <= not a or b;
    layer2_outputs(1847) <= not a;
    layer2_outputs(1848) <= not (a and b);
    layer2_outputs(1849) <= '0';
    layer2_outputs(1850) <= a xor b;
    layer2_outputs(1851) <= a and not b;
    layer2_outputs(1852) <= not b or a;
    layer2_outputs(1853) <= a and not b;
    layer2_outputs(1854) <= not a;
    layer2_outputs(1855) <= a and b;
    layer2_outputs(1856) <= not (a and b);
    layer2_outputs(1857) <= '1';
    layer2_outputs(1858) <= not b or a;
    layer2_outputs(1859) <= a and not b;
    layer2_outputs(1860) <= a or b;
    layer2_outputs(1861) <= not a;
    layer2_outputs(1862) <= not b or a;
    layer2_outputs(1863) <= '1';
    layer2_outputs(1864) <= a or b;
    layer2_outputs(1865) <= '0';
    layer2_outputs(1866) <= a;
    layer2_outputs(1867) <= a or b;
    layer2_outputs(1868) <= a and not b;
    layer2_outputs(1869) <= b and not a;
    layer2_outputs(1870) <= not a;
    layer2_outputs(1871) <= a and not b;
    layer2_outputs(1872) <= not a;
    layer2_outputs(1873) <= a xor b;
    layer2_outputs(1874) <= not (a or b);
    layer2_outputs(1875) <= '0';
    layer2_outputs(1876) <= a;
    layer2_outputs(1877) <= not a;
    layer2_outputs(1878) <= a and not b;
    layer2_outputs(1879) <= not b;
    layer2_outputs(1880) <= a;
    layer2_outputs(1881) <= not b;
    layer2_outputs(1882) <= a or b;
    layer2_outputs(1883) <= b;
    layer2_outputs(1884) <= b;
    layer2_outputs(1885) <= a and not b;
    layer2_outputs(1886) <= not a or b;
    layer2_outputs(1887) <= b and not a;
    layer2_outputs(1888) <= not a;
    layer2_outputs(1889) <= not a;
    layer2_outputs(1890) <= not (a and b);
    layer2_outputs(1891) <= a and not b;
    layer2_outputs(1892) <= b and not a;
    layer2_outputs(1893) <= a and b;
    layer2_outputs(1894) <= not (a and b);
    layer2_outputs(1895) <= b;
    layer2_outputs(1896) <= not b or a;
    layer2_outputs(1897) <= not a;
    layer2_outputs(1898) <= not b;
    layer2_outputs(1899) <= '1';
    layer2_outputs(1900) <= a or b;
    layer2_outputs(1901) <= a;
    layer2_outputs(1902) <= a and b;
    layer2_outputs(1903) <= a or b;
    layer2_outputs(1904) <= a and not b;
    layer2_outputs(1905) <= not (a and b);
    layer2_outputs(1906) <= not (a xor b);
    layer2_outputs(1907) <= '1';
    layer2_outputs(1908) <= a or b;
    layer2_outputs(1909) <= not (a or b);
    layer2_outputs(1910) <= not (a xor b);
    layer2_outputs(1911) <= not a or b;
    layer2_outputs(1912) <= a or b;
    layer2_outputs(1913) <= not a;
    layer2_outputs(1914) <= not (a and b);
    layer2_outputs(1915) <= not (a or b);
    layer2_outputs(1916) <= a or b;
    layer2_outputs(1917) <= '0';
    layer2_outputs(1918) <= not (a and b);
    layer2_outputs(1919) <= not b;
    layer2_outputs(1920) <= not a or b;
    layer2_outputs(1921) <= not b;
    layer2_outputs(1922) <= not b or a;
    layer2_outputs(1923) <= not a or b;
    layer2_outputs(1924) <= not b;
    layer2_outputs(1925) <= b and not a;
    layer2_outputs(1926) <= not a;
    layer2_outputs(1927) <= not b;
    layer2_outputs(1928) <= a and not b;
    layer2_outputs(1929) <= not b;
    layer2_outputs(1930) <= a;
    layer2_outputs(1931) <= not (a or b);
    layer2_outputs(1932) <= not (a or b);
    layer2_outputs(1933) <= a and b;
    layer2_outputs(1934) <= b;
    layer2_outputs(1935) <= not (a or b);
    layer2_outputs(1936) <= a and not b;
    layer2_outputs(1937) <= a xor b;
    layer2_outputs(1938) <= not a;
    layer2_outputs(1939) <= b;
    layer2_outputs(1940) <= not b;
    layer2_outputs(1941) <= not b;
    layer2_outputs(1942) <= a and b;
    layer2_outputs(1943) <= not b;
    layer2_outputs(1944) <= not (a or b);
    layer2_outputs(1945) <= not a;
    layer2_outputs(1946) <= a or b;
    layer2_outputs(1947) <= a and b;
    layer2_outputs(1948) <= '1';
    layer2_outputs(1949) <= not (a or b);
    layer2_outputs(1950) <= b and not a;
    layer2_outputs(1951) <= not (a xor b);
    layer2_outputs(1952) <= a and not b;
    layer2_outputs(1953) <= b;
    layer2_outputs(1954) <= a or b;
    layer2_outputs(1955) <= not (a and b);
    layer2_outputs(1956) <= not (a and b);
    layer2_outputs(1957) <= a and b;
    layer2_outputs(1958) <= '0';
    layer2_outputs(1959) <= '1';
    layer2_outputs(1960) <= '1';
    layer2_outputs(1961) <= not b or a;
    layer2_outputs(1962) <= a and not b;
    layer2_outputs(1963) <= a and b;
    layer2_outputs(1964) <= not (a xor b);
    layer2_outputs(1965) <= '1';
    layer2_outputs(1966) <= b and not a;
    layer2_outputs(1967) <= not a or b;
    layer2_outputs(1968) <= not b;
    layer2_outputs(1969) <= not b;
    layer2_outputs(1970) <= not b;
    layer2_outputs(1971) <= '0';
    layer2_outputs(1972) <= a and not b;
    layer2_outputs(1973) <= a;
    layer2_outputs(1974) <= not (a or b);
    layer2_outputs(1975) <= not b;
    layer2_outputs(1976) <= a;
    layer2_outputs(1977) <= a and not b;
    layer2_outputs(1978) <= a or b;
    layer2_outputs(1979) <= a and not b;
    layer2_outputs(1980) <= b;
    layer2_outputs(1981) <= not b;
    layer2_outputs(1982) <= a or b;
    layer2_outputs(1983) <= b;
    layer2_outputs(1984) <= not a or b;
    layer2_outputs(1985) <= not a or b;
    layer2_outputs(1986) <= a xor b;
    layer2_outputs(1987) <= a xor b;
    layer2_outputs(1988) <= a;
    layer2_outputs(1989) <= a;
    layer2_outputs(1990) <= '0';
    layer2_outputs(1991) <= a and not b;
    layer2_outputs(1992) <= not a or b;
    layer2_outputs(1993) <= b and not a;
    layer2_outputs(1994) <= not b or a;
    layer2_outputs(1995) <= not (a or b);
    layer2_outputs(1996) <= not b;
    layer2_outputs(1997) <= a;
    layer2_outputs(1998) <= not (a xor b);
    layer2_outputs(1999) <= not b;
    layer2_outputs(2000) <= not (a or b);
    layer2_outputs(2001) <= not b;
    layer2_outputs(2002) <= b and not a;
    layer2_outputs(2003) <= b and not a;
    layer2_outputs(2004) <= a xor b;
    layer2_outputs(2005) <= not b;
    layer2_outputs(2006) <= not (a or b);
    layer2_outputs(2007) <= b and not a;
    layer2_outputs(2008) <= not (a or b);
    layer2_outputs(2009) <= b;
    layer2_outputs(2010) <= b;
    layer2_outputs(2011) <= b and not a;
    layer2_outputs(2012) <= not (a or b);
    layer2_outputs(2013) <= not b or a;
    layer2_outputs(2014) <= not a;
    layer2_outputs(2015) <= not a;
    layer2_outputs(2016) <= a;
    layer2_outputs(2017) <= not a or b;
    layer2_outputs(2018) <= a and b;
    layer2_outputs(2019) <= '1';
    layer2_outputs(2020) <= a or b;
    layer2_outputs(2021) <= a and not b;
    layer2_outputs(2022) <= b;
    layer2_outputs(2023) <= not (a and b);
    layer2_outputs(2024) <= '1';
    layer2_outputs(2025) <= not a or b;
    layer2_outputs(2026) <= b;
    layer2_outputs(2027) <= a xor b;
    layer2_outputs(2028) <= a;
    layer2_outputs(2029) <= not b;
    layer2_outputs(2030) <= a or b;
    layer2_outputs(2031) <= not b or a;
    layer2_outputs(2032) <= not b or a;
    layer2_outputs(2033) <= a or b;
    layer2_outputs(2034) <= not b;
    layer2_outputs(2035) <= not (a and b);
    layer2_outputs(2036) <= '1';
    layer2_outputs(2037) <= not b;
    layer2_outputs(2038) <= not a or b;
    layer2_outputs(2039) <= not b;
    layer2_outputs(2040) <= '1';
    layer2_outputs(2041) <= a or b;
    layer2_outputs(2042) <= not b or a;
    layer2_outputs(2043) <= a;
    layer2_outputs(2044) <= b and not a;
    layer2_outputs(2045) <= a and not b;
    layer2_outputs(2046) <= a;
    layer2_outputs(2047) <= b and not a;
    layer2_outputs(2048) <= not (a and b);
    layer2_outputs(2049) <= not (a and b);
    layer2_outputs(2050) <= b and not a;
    layer2_outputs(2051) <= '1';
    layer2_outputs(2052) <= b and not a;
    layer2_outputs(2053) <= '0';
    layer2_outputs(2054) <= a or b;
    layer2_outputs(2055) <= not a or b;
    layer2_outputs(2056) <= a and not b;
    layer2_outputs(2057) <= not a;
    layer2_outputs(2058) <= not b;
    layer2_outputs(2059) <= a or b;
    layer2_outputs(2060) <= not b;
    layer2_outputs(2061) <= not b;
    layer2_outputs(2062) <= not a;
    layer2_outputs(2063) <= '1';
    layer2_outputs(2064) <= a and not b;
    layer2_outputs(2065) <= a and not b;
    layer2_outputs(2066) <= not b;
    layer2_outputs(2067) <= a and not b;
    layer2_outputs(2068) <= '0';
    layer2_outputs(2069) <= b;
    layer2_outputs(2070) <= not b;
    layer2_outputs(2071) <= '0';
    layer2_outputs(2072) <= a and not b;
    layer2_outputs(2073) <= b and not a;
    layer2_outputs(2074) <= a;
    layer2_outputs(2075) <= b;
    layer2_outputs(2076) <= not b or a;
    layer2_outputs(2077) <= a and not b;
    layer2_outputs(2078) <= not (a or b);
    layer2_outputs(2079) <= not b;
    layer2_outputs(2080) <= not (a and b);
    layer2_outputs(2081) <= a and not b;
    layer2_outputs(2082) <= '0';
    layer2_outputs(2083) <= not (a and b);
    layer2_outputs(2084) <= not a;
    layer2_outputs(2085) <= not b or a;
    layer2_outputs(2086) <= not b or a;
    layer2_outputs(2087) <= b and not a;
    layer2_outputs(2088) <= a;
    layer2_outputs(2089) <= a and not b;
    layer2_outputs(2090) <= '1';
    layer2_outputs(2091) <= a;
    layer2_outputs(2092) <= b;
    layer2_outputs(2093) <= not (a and b);
    layer2_outputs(2094) <= not b;
    layer2_outputs(2095) <= '0';
    layer2_outputs(2096) <= a;
    layer2_outputs(2097) <= not a or b;
    layer2_outputs(2098) <= b and not a;
    layer2_outputs(2099) <= b and not a;
    layer2_outputs(2100) <= not a;
    layer2_outputs(2101) <= not b or a;
    layer2_outputs(2102) <= b and not a;
    layer2_outputs(2103) <= b;
    layer2_outputs(2104) <= not b or a;
    layer2_outputs(2105) <= a;
    layer2_outputs(2106) <= a;
    layer2_outputs(2107) <= a;
    layer2_outputs(2108) <= a or b;
    layer2_outputs(2109) <= a and not b;
    layer2_outputs(2110) <= not b;
    layer2_outputs(2111) <= not (a or b);
    layer2_outputs(2112) <= a or b;
    layer2_outputs(2113) <= not a;
    layer2_outputs(2114) <= b;
    layer2_outputs(2115) <= b and not a;
    layer2_outputs(2116) <= a and not b;
    layer2_outputs(2117) <= not a or b;
    layer2_outputs(2118) <= not a or b;
    layer2_outputs(2119) <= not b or a;
    layer2_outputs(2120) <= not a or b;
    layer2_outputs(2121) <= not b or a;
    layer2_outputs(2122) <= not b;
    layer2_outputs(2123) <= b;
    layer2_outputs(2124) <= a and b;
    layer2_outputs(2125) <= a and b;
    layer2_outputs(2126) <= not b or a;
    layer2_outputs(2127) <= not (a xor b);
    layer2_outputs(2128) <= a;
    layer2_outputs(2129) <= a or b;
    layer2_outputs(2130) <= b and not a;
    layer2_outputs(2131) <= a;
    layer2_outputs(2132) <= b;
    layer2_outputs(2133) <= a;
    layer2_outputs(2134) <= not a or b;
    layer2_outputs(2135) <= not a;
    layer2_outputs(2136) <= a and not b;
    layer2_outputs(2137) <= not a or b;
    layer2_outputs(2138) <= not (a xor b);
    layer2_outputs(2139) <= b;
    layer2_outputs(2140) <= not a;
    layer2_outputs(2141) <= not b;
    layer2_outputs(2142) <= a;
    layer2_outputs(2143) <= not (a xor b);
    layer2_outputs(2144) <= not a or b;
    layer2_outputs(2145) <= not (a xor b);
    layer2_outputs(2146) <= not (a or b);
    layer2_outputs(2147) <= not (a or b);
    layer2_outputs(2148) <= a and b;
    layer2_outputs(2149) <= not a;
    layer2_outputs(2150) <= '0';
    layer2_outputs(2151) <= not a;
    layer2_outputs(2152) <= not (a and b);
    layer2_outputs(2153) <= not b;
    layer2_outputs(2154) <= '1';
    layer2_outputs(2155) <= not (a and b);
    layer2_outputs(2156) <= b;
    layer2_outputs(2157) <= a and not b;
    layer2_outputs(2158) <= b and not a;
    layer2_outputs(2159) <= not (a and b);
    layer2_outputs(2160) <= '0';
    layer2_outputs(2161) <= not b or a;
    layer2_outputs(2162) <= not (a xor b);
    layer2_outputs(2163) <= not b or a;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= a or b;
    layer2_outputs(2166) <= a;
    layer2_outputs(2167) <= not b;
    layer2_outputs(2168) <= a xor b;
    layer2_outputs(2169) <= a and not b;
    layer2_outputs(2170) <= b;
    layer2_outputs(2171) <= a and not b;
    layer2_outputs(2172) <= b;
    layer2_outputs(2173) <= not (a and b);
    layer2_outputs(2174) <= a and b;
    layer2_outputs(2175) <= a;
    layer2_outputs(2176) <= '0';
    layer2_outputs(2177) <= not (a and b);
    layer2_outputs(2178) <= a and b;
    layer2_outputs(2179) <= '1';
    layer2_outputs(2180) <= b and not a;
    layer2_outputs(2181) <= a and b;
    layer2_outputs(2182) <= a or b;
    layer2_outputs(2183) <= not a or b;
    layer2_outputs(2184) <= not (a xor b);
    layer2_outputs(2185) <= not (a and b);
    layer2_outputs(2186) <= b and not a;
    layer2_outputs(2187) <= '1';
    layer2_outputs(2188) <= not a or b;
    layer2_outputs(2189) <= a;
    layer2_outputs(2190) <= not b;
    layer2_outputs(2191) <= not (a or b);
    layer2_outputs(2192) <= not (a and b);
    layer2_outputs(2193) <= '1';
    layer2_outputs(2194) <= not (a and b);
    layer2_outputs(2195) <= a and not b;
    layer2_outputs(2196) <= '0';
    layer2_outputs(2197) <= not a;
    layer2_outputs(2198) <= a or b;
    layer2_outputs(2199) <= not a or b;
    layer2_outputs(2200) <= '0';
    layer2_outputs(2201) <= b;
    layer2_outputs(2202) <= not (a and b);
    layer2_outputs(2203) <= not b;
    layer2_outputs(2204) <= a or b;
    layer2_outputs(2205) <= not a or b;
    layer2_outputs(2206) <= not (a or b);
    layer2_outputs(2207) <= not b;
    layer2_outputs(2208) <= '0';
    layer2_outputs(2209) <= b and not a;
    layer2_outputs(2210) <= not a;
    layer2_outputs(2211) <= b;
    layer2_outputs(2212) <= not (a and b);
    layer2_outputs(2213) <= not b or a;
    layer2_outputs(2214) <= not b or a;
    layer2_outputs(2215) <= not a;
    layer2_outputs(2216) <= not a;
    layer2_outputs(2217) <= a xor b;
    layer2_outputs(2218) <= not b;
    layer2_outputs(2219) <= a;
    layer2_outputs(2220) <= not (a or b);
    layer2_outputs(2221) <= '1';
    layer2_outputs(2222) <= not a;
    layer2_outputs(2223) <= '0';
    layer2_outputs(2224) <= b;
    layer2_outputs(2225) <= '1';
    layer2_outputs(2226) <= '0';
    layer2_outputs(2227) <= not a;
    layer2_outputs(2228) <= b and not a;
    layer2_outputs(2229) <= not (a xor b);
    layer2_outputs(2230) <= not b;
    layer2_outputs(2231) <= not a;
    layer2_outputs(2232) <= not (a and b);
    layer2_outputs(2233) <= not a or b;
    layer2_outputs(2234) <= not (a or b);
    layer2_outputs(2235) <= a and not b;
    layer2_outputs(2236) <= not b or a;
    layer2_outputs(2237) <= b and not a;
    layer2_outputs(2238) <= '1';
    layer2_outputs(2239) <= a and not b;
    layer2_outputs(2240) <= b and not a;
    layer2_outputs(2241) <= '1';
    layer2_outputs(2242) <= not (a or b);
    layer2_outputs(2243) <= a and not b;
    layer2_outputs(2244) <= b and not a;
    layer2_outputs(2245) <= not (a or b);
    layer2_outputs(2246) <= a xor b;
    layer2_outputs(2247) <= not (a and b);
    layer2_outputs(2248) <= b and not a;
    layer2_outputs(2249) <= not (a and b);
    layer2_outputs(2250) <= b and not a;
    layer2_outputs(2251) <= '1';
    layer2_outputs(2252) <= not (a and b);
    layer2_outputs(2253) <= not (a and b);
    layer2_outputs(2254) <= '0';
    layer2_outputs(2255) <= not (a or b);
    layer2_outputs(2256) <= a;
    layer2_outputs(2257) <= a and not b;
    layer2_outputs(2258) <= a and b;
    layer2_outputs(2259) <= not (a and b);
    layer2_outputs(2260) <= a or b;
    layer2_outputs(2261) <= not a;
    layer2_outputs(2262) <= not (a and b);
    layer2_outputs(2263) <= not b or a;
    layer2_outputs(2264) <= a and b;
    layer2_outputs(2265) <= not a;
    layer2_outputs(2266) <= a and b;
    layer2_outputs(2267) <= '0';
    layer2_outputs(2268) <= a or b;
    layer2_outputs(2269) <= '0';
    layer2_outputs(2270) <= not a or b;
    layer2_outputs(2271) <= not a or b;
    layer2_outputs(2272) <= not a;
    layer2_outputs(2273) <= a xor b;
    layer2_outputs(2274) <= b;
    layer2_outputs(2275) <= a and b;
    layer2_outputs(2276) <= a;
    layer2_outputs(2277) <= a;
    layer2_outputs(2278) <= '1';
    layer2_outputs(2279) <= not (a xor b);
    layer2_outputs(2280) <= not b;
    layer2_outputs(2281) <= b;
    layer2_outputs(2282) <= '1';
    layer2_outputs(2283) <= not b;
    layer2_outputs(2284) <= not a;
    layer2_outputs(2285) <= b and not a;
    layer2_outputs(2286) <= '1';
    layer2_outputs(2287) <= a or b;
    layer2_outputs(2288) <= not (a and b);
    layer2_outputs(2289) <= not a;
    layer2_outputs(2290) <= not (a or b);
    layer2_outputs(2291) <= a and b;
    layer2_outputs(2292) <= b and not a;
    layer2_outputs(2293) <= '0';
    layer2_outputs(2294) <= a;
    layer2_outputs(2295) <= not (a xor b);
    layer2_outputs(2296) <= '0';
    layer2_outputs(2297) <= not (a or b);
    layer2_outputs(2298) <= not (a xor b);
    layer2_outputs(2299) <= a and b;
    layer2_outputs(2300) <= a and not b;
    layer2_outputs(2301) <= not (a and b);
    layer2_outputs(2302) <= a xor b;
    layer2_outputs(2303) <= b;
    layer2_outputs(2304) <= not b;
    layer2_outputs(2305) <= '0';
    layer2_outputs(2306) <= a or b;
    layer2_outputs(2307) <= a or b;
    layer2_outputs(2308) <= not b;
    layer2_outputs(2309) <= not (a or b);
    layer2_outputs(2310) <= a;
    layer2_outputs(2311) <= b;
    layer2_outputs(2312) <= not (a and b);
    layer2_outputs(2313) <= not a or b;
    layer2_outputs(2314) <= not b;
    layer2_outputs(2315) <= a and b;
    layer2_outputs(2316) <= b;
    layer2_outputs(2317) <= a and not b;
    layer2_outputs(2318) <= not a;
    layer2_outputs(2319) <= a and not b;
    layer2_outputs(2320) <= not a;
    layer2_outputs(2321) <= '0';
    layer2_outputs(2322) <= not b;
    layer2_outputs(2323) <= not b;
    layer2_outputs(2324) <= not b;
    layer2_outputs(2325) <= not (a xor b);
    layer2_outputs(2326) <= a xor b;
    layer2_outputs(2327) <= '1';
    layer2_outputs(2328) <= not b or a;
    layer2_outputs(2329) <= not b;
    layer2_outputs(2330) <= '0';
    layer2_outputs(2331) <= not b or a;
    layer2_outputs(2332) <= not (a and b);
    layer2_outputs(2333) <= not a;
    layer2_outputs(2334) <= not b;
    layer2_outputs(2335) <= b and not a;
    layer2_outputs(2336) <= not a or b;
    layer2_outputs(2337) <= a;
    layer2_outputs(2338) <= a or b;
    layer2_outputs(2339) <= not (a or b);
    layer2_outputs(2340) <= a and b;
    layer2_outputs(2341) <= b;
    layer2_outputs(2342) <= not b;
    layer2_outputs(2343) <= '1';
    layer2_outputs(2344) <= not (a and b);
    layer2_outputs(2345) <= not a or b;
    layer2_outputs(2346) <= a and not b;
    layer2_outputs(2347) <= '1';
    layer2_outputs(2348) <= not b or a;
    layer2_outputs(2349) <= '1';
    layer2_outputs(2350) <= b;
    layer2_outputs(2351) <= not a or b;
    layer2_outputs(2352) <= a and not b;
    layer2_outputs(2353) <= not b or a;
    layer2_outputs(2354) <= not a;
    layer2_outputs(2355) <= not (a and b);
    layer2_outputs(2356) <= not (a or b);
    layer2_outputs(2357) <= not a;
    layer2_outputs(2358) <= not b or a;
    layer2_outputs(2359) <= a and not b;
    layer2_outputs(2360) <= '0';
    layer2_outputs(2361) <= not (a or b);
    layer2_outputs(2362) <= '1';
    layer2_outputs(2363) <= b;
    layer2_outputs(2364) <= '1';
    layer2_outputs(2365) <= b and not a;
    layer2_outputs(2366) <= not b or a;
    layer2_outputs(2367) <= not (a xor b);
    layer2_outputs(2368) <= '1';
    layer2_outputs(2369) <= not a;
    layer2_outputs(2370) <= a and not b;
    layer2_outputs(2371) <= not a;
    layer2_outputs(2372) <= a and not b;
    layer2_outputs(2373) <= '0';
    layer2_outputs(2374) <= not a;
    layer2_outputs(2375) <= a and not b;
    layer2_outputs(2376) <= '0';
    layer2_outputs(2377) <= a and not b;
    layer2_outputs(2378) <= a and b;
    layer2_outputs(2379) <= not (a and b);
    layer2_outputs(2380) <= not a or b;
    layer2_outputs(2381) <= not a;
    layer2_outputs(2382) <= a;
    layer2_outputs(2383) <= a;
    layer2_outputs(2384) <= not (a and b);
    layer2_outputs(2385) <= not (a or b);
    layer2_outputs(2386) <= not b;
    layer2_outputs(2387) <= not (a and b);
    layer2_outputs(2388) <= b and not a;
    layer2_outputs(2389) <= not (a or b);
    layer2_outputs(2390) <= a or b;
    layer2_outputs(2391) <= '1';
    layer2_outputs(2392) <= not b;
    layer2_outputs(2393) <= not a;
    layer2_outputs(2394) <= a;
    layer2_outputs(2395) <= not (a xor b);
    layer2_outputs(2396) <= '1';
    layer2_outputs(2397) <= not a;
    layer2_outputs(2398) <= a and not b;
    layer2_outputs(2399) <= a or b;
    layer2_outputs(2400) <= b and not a;
    layer2_outputs(2401) <= not (a or b);
    layer2_outputs(2402) <= not b or a;
    layer2_outputs(2403) <= not a;
    layer2_outputs(2404) <= a and b;
    layer2_outputs(2405) <= a or b;
    layer2_outputs(2406) <= a or b;
    layer2_outputs(2407) <= not b;
    layer2_outputs(2408) <= not a;
    layer2_outputs(2409) <= a or b;
    layer2_outputs(2410) <= a and not b;
    layer2_outputs(2411) <= a xor b;
    layer2_outputs(2412) <= '1';
    layer2_outputs(2413) <= a or b;
    layer2_outputs(2414) <= b and not a;
    layer2_outputs(2415) <= a;
    layer2_outputs(2416) <= not b;
    layer2_outputs(2417) <= not (a or b);
    layer2_outputs(2418) <= b and not a;
    layer2_outputs(2419) <= a and not b;
    layer2_outputs(2420) <= not a;
    layer2_outputs(2421) <= not b or a;
    layer2_outputs(2422) <= '1';
    layer2_outputs(2423) <= a and not b;
    layer2_outputs(2424) <= not b;
    layer2_outputs(2425) <= '0';
    layer2_outputs(2426) <= a and b;
    layer2_outputs(2427) <= a xor b;
    layer2_outputs(2428) <= a and not b;
    layer2_outputs(2429) <= '0';
    layer2_outputs(2430) <= a;
    layer2_outputs(2431) <= a and b;
    layer2_outputs(2432) <= a;
    layer2_outputs(2433) <= a;
    layer2_outputs(2434) <= b and not a;
    layer2_outputs(2435) <= b;
    layer2_outputs(2436) <= not a;
    layer2_outputs(2437) <= b;
    layer2_outputs(2438) <= not b or a;
    layer2_outputs(2439) <= b;
    layer2_outputs(2440) <= not a;
    layer2_outputs(2441) <= not b or a;
    layer2_outputs(2442) <= a and b;
    layer2_outputs(2443) <= not a;
    layer2_outputs(2444) <= not b;
    layer2_outputs(2445) <= not a;
    layer2_outputs(2446) <= b and not a;
    layer2_outputs(2447) <= not a or b;
    layer2_outputs(2448) <= a or b;
    layer2_outputs(2449) <= b;
    layer2_outputs(2450) <= not (a xor b);
    layer2_outputs(2451) <= not (a or b);
    layer2_outputs(2452) <= not a;
    layer2_outputs(2453) <= not b or a;
    layer2_outputs(2454) <= b;
    layer2_outputs(2455) <= a and b;
    layer2_outputs(2456) <= not (a or b);
    layer2_outputs(2457) <= b and not a;
    layer2_outputs(2458) <= b and not a;
    layer2_outputs(2459) <= b;
    layer2_outputs(2460) <= b;
    layer2_outputs(2461) <= not (a and b);
    layer2_outputs(2462) <= b;
    layer2_outputs(2463) <= a and not b;
    layer2_outputs(2464) <= a and not b;
    layer2_outputs(2465) <= a;
    layer2_outputs(2466) <= a and b;
    layer2_outputs(2467) <= not (a and b);
    layer2_outputs(2468) <= a;
    layer2_outputs(2469) <= b and not a;
    layer2_outputs(2470) <= not a or b;
    layer2_outputs(2471) <= a and b;
    layer2_outputs(2472) <= not b;
    layer2_outputs(2473) <= not (a and b);
    layer2_outputs(2474) <= not a or b;
    layer2_outputs(2475) <= b;
    layer2_outputs(2476) <= '1';
    layer2_outputs(2477) <= a and b;
    layer2_outputs(2478) <= a or b;
    layer2_outputs(2479) <= not b or a;
    layer2_outputs(2480) <= not (a and b);
    layer2_outputs(2481) <= '0';
    layer2_outputs(2482) <= a;
    layer2_outputs(2483) <= not b;
    layer2_outputs(2484) <= '0';
    layer2_outputs(2485) <= a and not b;
    layer2_outputs(2486) <= '1';
    layer2_outputs(2487) <= not b;
    layer2_outputs(2488) <= not (a or b);
    layer2_outputs(2489) <= not (a or b);
    layer2_outputs(2490) <= a and b;
    layer2_outputs(2491) <= a;
    layer2_outputs(2492) <= not b or a;
    layer2_outputs(2493) <= not (a and b);
    layer2_outputs(2494) <= a and not b;
    layer2_outputs(2495) <= not a;
    layer2_outputs(2496) <= a;
    layer2_outputs(2497) <= not b or a;
    layer2_outputs(2498) <= not a;
    layer2_outputs(2499) <= not (a and b);
    layer2_outputs(2500) <= a;
    layer2_outputs(2501) <= not (a or b);
    layer2_outputs(2502) <= not b or a;
    layer2_outputs(2503) <= not (a or b);
    layer2_outputs(2504) <= not b or a;
    layer2_outputs(2505) <= a or b;
    layer2_outputs(2506) <= b and not a;
    layer2_outputs(2507) <= not b;
    layer2_outputs(2508) <= '1';
    layer2_outputs(2509) <= a and b;
    layer2_outputs(2510) <= not (a or b);
    layer2_outputs(2511) <= '0';
    layer2_outputs(2512) <= a xor b;
    layer2_outputs(2513) <= a;
    layer2_outputs(2514) <= not b or a;
    layer2_outputs(2515) <= '0';
    layer2_outputs(2516) <= not a or b;
    layer2_outputs(2517) <= b;
    layer2_outputs(2518) <= not (a and b);
    layer2_outputs(2519) <= a;
    layer2_outputs(2520) <= a or b;
    layer2_outputs(2521) <= '1';
    layer2_outputs(2522) <= not a or b;
    layer2_outputs(2523) <= a and not b;
    layer2_outputs(2524) <= not b;
    layer2_outputs(2525) <= not a or b;
    layer2_outputs(2526) <= a xor b;
    layer2_outputs(2527) <= not a;
    layer2_outputs(2528) <= not (a and b);
    layer2_outputs(2529) <= not b or a;
    layer2_outputs(2530) <= not a;
    layer2_outputs(2531) <= not (a and b);
    layer2_outputs(2532) <= a and not b;
    layer2_outputs(2533) <= not a;
    layer2_outputs(2534) <= not a;
    layer2_outputs(2535) <= a;
    layer2_outputs(2536) <= '0';
    layer2_outputs(2537) <= '0';
    layer2_outputs(2538) <= '1';
    layer2_outputs(2539) <= a and b;
    layer2_outputs(2540) <= not b or a;
    layer2_outputs(2541) <= a xor b;
    layer2_outputs(2542) <= not (a or b);
    layer2_outputs(2543) <= a;
    layer2_outputs(2544) <= not (a or b);
    layer2_outputs(2545) <= not a;
    layer2_outputs(2546) <= a and not b;
    layer2_outputs(2547) <= not (a or b);
    layer2_outputs(2548) <= b;
    layer2_outputs(2549) <= not b;
    layer2_outputs(2550) <= b;
    layer2_outputs(2551) <= b and not a;
    layer2_outputs(2552) <= not b;
    layer2_outputs(2553) <= a and b;
    layer2_outputs(2554) <= a and not b;
    layer2_outputs(2555) <= not b;
    layer2_outputs(2556) <= a or b;
    layer2_outputs(2557) <= a and b;
    layer2_outputs(2558) <= '0';
    layer2_outputs(2559) <= b and not a;
    layer2_outputs(2560) <= not b;
    layer2_outputs(2561) <= not b;
    layer2_outputs(2562) <= '1';
    layer2_outputs(2563) <= not b;
    layer2_outputs(2564) <= a;
    layer2_outputs(2565) <= not (a or b);
    layer2_outputs(2566) <= not b or a;
    layer2_outputs(2567) <= a or b;
    layer2_outputs(2568) <= not b or a;
    layer2_outputs(2569) <= not a;
    layer2_outputs(2570) <= '0';
    layer2_outputs(2571) <= b;
    layer2_outputs(2572) <= not a or b;
    layer2_outputs(2573) <= a xor b;
    layer2_outputs(2574) <= not a;
    layer2_outputs(2575) <= b;
    layer2_outputs(2576) <= not a or b;
    layer2_outputs(2577) <= b;
    layer2_outputs(2578) <= not a;
    layer2_outputs(2579) <= not a or b;
    layer2_outputs(2580) <= b;
    layer2_outputs(2581) <= a xor b;
    layer2_outputs(2582) <= not a or b;
    layer2_outputs(2583) <= not b;
    layer2_outputs(2584) <= not b or a;
    layer2_outputs(2585) <= a and b;
    layer2_outputs(2586) <= '0';
    layer2_outputs(2587) <= a xor b;
    layer2_outputs(2588) <= a and b;
    layer2_outputs(2589) <= a or b;
    layer2_outputs(2590) <= a and b;
    layer2_outputs(2591) <= not (a and b);
    layer2_outputs(2592) <= a and not b;
    layer2_outputs(2593) <= not a;
    layer2_outputs(2594) <= not b;
    layer2_outputs(2595) <= not b or a;
    layer2_outputs(2596) <= not a;
    layer2_outputs(2597) <= a xor b;
    layer2_outputs(2598) <= not b or a;
    layer2_outputs(2599) <= not (a and b);
    layer2_outputs(2600) <= not (a or b);
    layer2_outputs(2601) <= a xor b;
    layer2_outputs(2602) <= '0';
    layer2_outputs(2603) <= a xor b;
    layer2_outputs(2604) <= a or b;
    layer2_outputs(2605) <= a;
    layer2_outputs(2606) <= '1';
    layer2_outputs(2607) <= a;
    layer2_outputs(2608) <= not b;
    layer2_outputs(2609) <= not (a or b);
    layer2_outputs(2610) <= b;
    layer2_outputs(2611) <= not b or a;
    layer2_outputs(2612) <= a or b;
    layer2_outputs(2613) <= not a or b;
    layer2_outputs(2614) <= not (a or b);
    layer2_outputs(2615) <= '0';
    layer2_outputs(2616) <= b and not a;
    layer2_outputs(2617) <= not b or a;
    layer2_outputs(2618) <= not b;
    layer2_outputs(2619) <= a and not b;
    layer2_outputs(2620) <= not (a or b);
    layer2_outputs(2621) <= not b or a;
    layer2_outputs(2622) <= a;
    layer2_outputs(2623) <= not b;
    layer2_outputs(2624) <= b;
    layer2_outputs(2625) <= a;
    layer2_outputs(2626) <= not a;
    layer2_outputs(2627) <= a or b;
    layer2_outputs(2628) <= a and b;
    layer2_outputs(2629) <= a and b;
    layer2_outputs(2630) <= a and b;
    layer2_outputs(2631) <= not b or a;
    layer2_outputs(2632) <= not a or b;
    layer2_outputs(2633) <= not a;
    layer2_outputs(2634) <= a xor b;
    layer2_outputs(2635) <= b;
    layer2_outputs(2636) <= b and not a;
    layer2_outputs(2637) <= a or b;
    layer2_outputs(2638) <= not b or a;
    layer2_outputs(2639) <= '0';
    layer2_outputs(2640) <= '1';
    layer2_outputs(2641) <= b;
    layer2_outputs(2642) <= b and not a;
    layer2_outputs(2643) <= b;
    layer2_outputs(2644) <= b and not a;
    layer2_outputs(2645) <= a and b;
    layer2_outputs(2646) <= '0';
    layer2_outputs(2647) <= b;
    layer2_outputs(2648) <= a and b;
    layer2_outputs(2649) <= a;
    layer2_outputs(2650) <= b;
    layer2_outputs(2651) <= not (a or b);
    layer2_outputs(2652) <= a and b;
    layer2_outputs(2653) <= not (a or b);
    layer2_outputs(2654) <= not a;
    layer2_outputs(2655) <= '0';
    layer2_outputs(2656) <= not (a xor b);
    layer2_outputs(2657) <= a and not b;
    layer2_outputs(2658) <= not (a and b);
    layer2_outputs(2659) <= not b;
    layer2_outputs(2660) <= not (a and b);
    layer2_outputs(2661) <= '0';
    layer2_outputs(2662) <= not b or a;
    layer2_outputs(2663) <= a;
    layer2_outputs(2664) <= not a;
    layer2_outputs(2665) <= not b;
    layer2_outputs(2666) <= not a or b;
    layer2_outputs(2667) <= a and b;
    layer2_outputs(2668) <= '1';
    layer2_outputs(2669) <= b;
    layer2_outputs(2670) <= not a;
    layer2_outputs(2671) <= b;
    layer2_outputs(2672) <= '0';
    layer2_outputs(2673) <= not a;
    layer2_outputs(2674) <= not b or a;
    layer2_outputs(2675) <= '0';
    layer2_outputs(2676) <= a and not b;
    layer2_outputs(2677) <= not b;
    layer2_outputs(2678) <= not b;
    layer2_outputs(2679) <= not (a or b);
    layer2_outputs(2680) <= a or b;
    layer2_outputs(2681) <= not b;
    layer2_outputs(2682) <= not (a or b);
    layer2_outputs(2683) <= a;
    layer2_outputs(2684) <= b and not a;
    layer2_outputs(2685) <= '1';
    layer2_outputs(2686) <= b;
    layer2_outputs(2687) <= a and not b;
    layer2_outputs(2688) <= a and b;
    layer2_outputs(2689) <= not a;
    layer2_outputs(2690) <= not (a and b);
    layer2_outputs(2691) <= b;
    layer2_outputs(2692) <= a;
    layer2_outputs(2693) <= a and b;
    layer2_outputs(2694) <= a or b;
    layer2_outputs(2695) <= not (a and b);
    layer2_outputs(2696) <= not a or b;
    layer2_outputs(2697) <= b and not a;
    layer2_outputs(2698) <= '1';
    layer2_outputs(2699) <= b and not a;
    layer2_outputs(2700) <= '0';
    layer2_outputs(2701) <= b;
    layer2_outputs(2702) <= not (a or b);
    layer2_outputs(2703) <= not a or b;
    layer2_outputs(2704) <= b and not a;
    layer2_outputs(2705) <= b;
    layer2_outputs(2706) <= a xor b;
    layer2_outputs(2707) <= '1';
    layer2_outputs(2708) <= not b;
    layer2_outputs(2709) <= a;
    layer2_outputs(2710) <= not a or b;
    layer2_outputs(2711) <= not a or b;
    layer2_outputs(2712) <= '1';
    layer2_outputs(2713) <= not a or b;
    layer2_outputs(2714) <= '0';
    layer2_outputs(2715) <= b;
    layer2_outputs(2716) <= '0';
    layer2_outputs(2717) <= b and not a;
    layer2_outputs(2718) <= b;
    layer2_outputs(2719) <= a and b;
    layer2_outputs(2720) <= not b or a;
    layer2_outputs(2721) <= not a;
    layer2_outputs(2722) <= a and b;
    layer2_outputs(2723) <= a and b;
    layer2_outputs(2724) <= a;
    layer2_outputs(2725) <= a;
    layer2_outputs(2726) <= not b;
    layer2_outputs(2727) <= not b;
    layer2_outputs(2728) <= b and not a;
    layer2_outputs(2729) <= not a or b;
    layer2_outputs(2730) <= b;
    layer2_outputs(2731) <= not b or a;
    layer2_outputs(2732) <= not b;
    layer2_outputs(2733) <= a or b;
    layer2_outputs(2734) <= not a;
    layer2_outputs(2735) <= b and not a;
    layer2_outputs(2736) <= not b;
    layer2_outputs(2737) <= a or b;
    layer2_outputs(2738) <= a or b;
    layer2_outputs(2739) <= not a;
    layer2_outputs(2740) <= b;
    layer2_outputs(2741) <= not (a or b);
    layer2_outputs(2742) <= '0';
    layer2_outputs(2743) <= not a or b;
    layer2_outputs(2744) <= a and b;
    layer2_outputs(2745) <= not b or a;
    layer2_outputs(2746) <= not b;
    layer2_outputs(2747) <= a and b;
    layer2_outputs(2748) <= not (a or b);
    layer2_outputs(2749) <= a;
    layer2_outputs(2750) <= '0';
    layer2_outputs(2751) <= a and b;
    layer2_outputs(2752) <= not a or b;
    layer2_outputs(2753) <= b and not a;
    layer2_outputs(2754) <= a and b;
    layer2_outputs(2755) <= b;
    layer2_outputs(2756) <= not b;
    layer2_outputs(2757) <= not a;
    layer2_outputs(2758) <= not a;
    layer2_outputs(2759) <= b;
    layer2_outputs(2760) <= not b;
    layer2_outputs(2761) <= b;
    layer2_outputs(2762) <= a or b;
    layer2_outputs(2763) <= a or b;
    layer2_outputs(2764) <= a and b;
    layer2_outputs(2765) <= not (a and b);
    layer2_outputs(2766) <= not (a or b);
    layer2_outputs(2767) <= not b or a;
    layer2_outputs(2768) <= '0';
    layer2_outputs(2769) <= not (a and b);
    layer2_outputs(2770) <= not (a and b);
    layer2_outputs(2771) <= not a;
    layer2_outputs(2772) <= a and b;
    layer2_outputs(2773) <= b and not a;
    layer2_outputs(2774) <= a and not b;
    layer2_outputs(2775) <= not b;
    layer2_outputs(2776) <= not a;
    layer2_outputs(2777) <= not a or b;
    layer2_outputs(2778) <= b;
    layer2_outputs(2779) <= not a or b;
    layer2_outputs(2780) <= not (a and b);
    layer2_outputs(2781) <= '0';
    layer2_outputs(2782) <= a and not b;
    layer2_outputs(2783) <= b and not a;
    layer2_outputs(2784) <= a and not b;
    layer2_outputs(2785) <= not (a and b);
    layer2_outputs(2786) <= a or b;
    layer2_outputs(2787) <= b and not a;
    layer2_outputs(2788) <= not (a or b);
    layer2_outputs(2789) <= a and b;
    layer2_outputs(2790) <= b;
    layer2_outputs(2791) <= not (a and b);
    layer2_outputs(2792) <= a;
    layer2_outputs(2793) <= not (a and b);
    layer2_outputs(2794) <= '1';
    layer2_outputs(2795) <= not a;
    layer2_outputs(2796) <= '1';
    layer2_outputs(2797) <= a and b;
    layer2_outputs(2798) <= not a;
    layer2_outputs(2799) <= '0';
    layer2_outputs(2800) <= a and b;
    layer2_outputs(2801) <= not (a and b);
    layer2_outputs(2802) <= a and b;
    layer2_outputs(2803) <= b;
    layer2_outputs(2804) <= not (a xor b);
    layer2_outputs(2805) <= not b;
    layer2_outputs(2806) <= not a or b;
    layer2_outputs(2807) <= not (a xor b);
    layer2_outputs(2808) <= a or b;
    layer2_outputs(2809) <= not (a and b);
    layer2_outputs(2810) <= a xor b;
    layer2_outputs(2811) <= b;
    layer2_outputs(2812) <= not (a and b);
    layer2_outputs(2813) <= b and not a;
    layer2_outputs(2814) <= a;
    layer2_outputs(2815) <= a and b;
    layer2_outputs(2816) <= '1';
    layer2_outputs(2817) <= a xor b;
    layer2_outputs(2818) <= a and not b;
    layer2_outputs(2819) <= not a or b;
    layer2_outputs(2820) <= a;
    layer2_outputs(2821) <= '0';
    layer2_outputs(2822) <= a and not b;
    layer2_outputs(2823) <= not a;
    layer2_outputs(2824) <= a or b;
    layer2_outputs(2825) <= '0';
    layer2_outputs(2826) <= not b;
    layer2_outputs(2827) <= not b;
    layer2_outputs(2828) <= not (a and b);
    layer2_outputs(2829) <= not a;
    layer2_outputs(2830) <= b;
    layer2_outputs(2831) <= '1';
    layer2_outputs(2832) <= not a or b;
    layer2_outputs(2833) <= '1';
    layer2_outputs(2834) <= a and not b;
    layer2_outputs(2835) <= not (a and b);
    layer2_outputs(2836) <= not a;
    layer2_outputs(2837) <= a;
    layer2_outputs(2838) <= not b;
    layer2_outputs(2839) <= not b;
    layer2_outputs(2840) <= not a;
    layer2_outputs(2841) <= not (a or b);
    layer2_outputs(2842) <= not b;
    layer2_outputs(2843) <= a;
    layer2_outputs(2844) <= not a or b;
    layer2_outputs(2845) <= b;
    layer2_outputs(2846) <= not b;
    layer2_outputs(2847) <= b;
    layer2_outputs(2848) <= not a or b;
    layer2_outputs(2849) <= not (a or b);
    layer2_outputs(2850) <= b;
    layer2_outputs(2851) <= not (a and b);
    layer2_outputs(2852) <= not b;
    layer2_outputs(2853) <= '0';
    layer2_outputs(2854) <= not b or a;
    layer2_outputs(2855) <= not b;
    layer2_outputs(2856) <= not a;
    layer2_outputs(2857) <= b;
    layer2_outputs(2858) <= '1';
    layer2_outputs(2859) <= a and not b;
    layer2_outputs(2860) <= not (a xor b);
    layer2_outputs(2861) <= b;
    layer2_outputs(2862) <= a;
    layer2_outputs(2863) <= not a or b;
    layer2_outputs(2864) <= not (a and b);
    layer2_outputs(2865) <= a and b;
    layer2_outputs(2866) <= a;
    layer2_outputs(2867) <= a or b;
    layer2_outputs(2868) <= a and b;
    layer2_outputs(2869) <= not b;
    layer2_outputs(2870) <= '1';
    layer2_outputs(2871) <= not b;
    layer2_outputs(2872) <= not (a and b);
    layer2_outputs(2873) <= not b;
    layer2_outputs(2874) <= not a;
    layer2_outputs(2875) <= b and not a;
    layer2_outputs(2876) <= not b;
    layer2_outputs(2877) <= a;
    layer2_outputs(2878) <= not a;
    layer2_outputs(2879) <= b;
    layer2_outputs(2880) <= not a;
    layer2_outputs(2881) <= a and b;
    layer2_outputs(2882) <= not b;
    layer2_outputs(2883) <= a and b;
    layer2_outputs(2884) <= not (a xor b);
    layer2_outputs(2885) <= a;
    layer2_outputs(2886) <= not (a and b);
    layer2_outputs(2887) <= not b or a;
    layer2_outputs(2888) <= b and not a;
    layer2_outputs(2889) <= b;
    layer2_outputs(2890) <= not b;
    layer2_outputs(2891) <= '0';
    layer2_outputs(2892) <= not b;
    layer2_outputs(2893) <= not (a xor b);
    layer2_outputs(2894) <= not a or b;
    layer2_outputs(2895) <= not (a or b);
    layer2_outputs(2896) <= a or b;
    layer2_outputs(2897) <= '1';
    layer2_outputs(2898) <= b and not a;
    layer2_outputs(2899) <= not (a and b);
    layer2_outputs(2900) <= a;
    layer2_outputs(2901) <= not b;
    layer2_outputs(2902) <= '1';
    layer2_outputs(2903) <= a and not b;
    layer2_outputs(2904) <= '0';
    layer2_outputs(2905) <= a and b;
    layer2_outputs(2906) <= '1';
    layer2_outputs(2907) <= a and not b;
    layer2_outputs(2908) <= not b;
    layer2_outputs(2909) <= a and not b;
    layer2_outputs(2910) <= a and not b;
    layer2_outputs(2911) <= '0';
    layer2_outputs(2912) <= a and b;
    layer2_outputs(2913) <= not a or b;
    layer2_outputs(2914) <= b;
    layer2_outputs(2915) <= b and not a;
    layer2_outputs(2916) <= not (a xor b);
    layer2_outputs(2917) <= '1';
    layer2_outputs(2918) <= not (a or b);
    layer2_outputs(2919) <= b and not a;
    layer2_outputs(2920) <= '1';
    layer2_outputs(2921) <= not (a xor b);
    layer2_outputs(2922) <= not a or b;
    layer2_outputs(2923) <= not (a or b);
    layer2_outputs(2924) <= b and not a;
    layer2_outputs(2925) <= b and not a;
    layer2_outputs(2926) <= '1';
    layer2_outputs(2927) <= not b or a;
    layer2_outputs(2928) <= not (a or b);
    layer2_outputs(2929) <= not b or a;
    layer2_outputs(2930) <= a;
    layer2_outputs(2931) <= a and not b;
    layer2_outputs(2932) <= not (a and b);
    layer2_outputs(2933) <= a and b;
    layer2_outputs(2934) <= a;
    layer2_outputs(2935) <= b;
    layer2_outputs(2936) <= a;
    layer2_outputs(2937) <= b;
    layer2_outputs(2938) <= not (a xor b);
    layer2_outputs(2939) <= a xor b;
    layer2_outputs(2940) <= b and not a;
    layer2_outputs(2941) <= b;
    layer2_outputs(2942) <= a and b;
    layer2_outputs(2943) <= not b;
    layer2_outputs(2944) <= a and not b;
    layer2_outputs(2945) <= not a;
    layer2_outputs(2946) <= '0';
    layer2_outputs(2947) <= not (a xor b);
    layer2_outputs(2948) <= not b or a;
    layer2_outputs(2949) <= not (a and b);
    layer2_outputs(2950) <= b and not a;
    layer2_outputs(2951) <= b and not a;
    layer2_outputs(2952) <= a;
    layer2_outputs(2953) <= not a;
    layer2_outputs(2954) <= b and not a;
    layer2_outputs(2955) <= not a or b;
    layer2_outputs(2956) <= a or b;
    layer2_outputs(2957) <= a and not b;
    layer2_outputs(2958) <= '0';
    layer2_outputs(2959) <= not a;
    layer2_outputs(2960) <= b and not a;
    layer2_outputs(2961) <= not (a xor b);
    layer2_outputs(2962) <= not b or a;
    layer2_outputs(2963) <= a or b;
    layer2_outputs(2964) <= a and not b;
    layer2_outputs(2965) <= not a;
    layer2_outputs(2966) <= b;
    layer2_outputs(2967) <= not (a or b);
    layer2_outputs(2968) <= not (a and b);
    layer2_outputs(2969) <= not a or b;
    layer2_outputs(2970) <= a and not b;
    layer2_outputs(2971) <= not (a xor b);
    layer2_outputs(2972) <= a;
    layer2_outputs(2973) <= a xor b;
    layer2_outputs(2974) <= a;
    layer2_outputs(2975) <= a and not b;
    layer2_outputs(2976) <= '0';
    layer2_outputs(2977) <= a and not b;
    layer2_outputs(2978) <= b;
    layer2_outputs(2979) <= '1';
    layer2_outputs(2980) <= not b;
    layer2_outputs(2981) <= '0';
    layer2_outputs(2982) <= not b;
    layer2_outputs(2983) <= a xor b;
    layer2_outputs(2984) <= a;
    layer2_outputs(2985) <= not a or b;
    layer2_outputs(2986) <= a;
    layer2_outputs(2987) <= a;
    layer2_outputs(2988) <= a and not b;
    layer2_outputs(2989) <= not (a or b);
    layer2_outputs(2990) <= not a or b;
    layer2_outputs(2991) <= not (a and b);
    layer2_outputs(2992) <= a and not b;
    layer2_outputs(2993) <= '0';
    layer2_outputs(2994) <= not a;
    layer2_outputs(2995) <= a and not b;
    layer2_outputs(2996) <= '1';
    layer2_outputs(2997) <= a and not b;
    layer2_outputs(2998) <= not (a and b);
    layer2_outputs(2999) <= not b or a;
    layer2_outputs(3000) <= not a;
    layer2_outputs(3001) <= a and b;
    layer2_outputs(3002) <= a xor b;
    layer2_outputs(3003) <= a;
    layer2_outputs(3004) <= '0';
    layer2_outputs(3005) <= a and not b;
    layer2_outputs(3006) <= not b;
    layer2_outputs(3007) <= not b;
    layer2_outputs(3008) <= a and not b;
    layer2_outputs(3009) <= not a;
    layer2_outputs(3010) <= not a;
    layer2_outputs(3011) <= '0';
    layer2_outputs(3012) <= b;
    layer2_outputs(3013) <= a;
    layer2_outputs(3014) <= b;
    layer2_outputs(3015) <= not (a xor b);
    layer2_outputs(3016) <= not (a xor b);
    layer2_outputs(3017) <= '0';
    layer2_outputs(3018) <= a;
    layer2_outputs(3019) <= a or b;
    layer2_outputs(3020) <= not b or a;
    layer2_outputs(3021) <= not b or a;
    layer2_outputs(3022) <= a and b;
    layer2_outputs(3023) <= a and not b;
    layer2_outputs(3024) <= not b or a;
    layer2_outputs(3025) <= a xor b;
    layer2_outputs(3026) <= not b or a;
    layer2_outputs(3027) <= not a;
    layer2_outputs(3028) <= not a or b;
    layer2_outputs(3029) <= not (a and b);
    layer2_outputs(3030) <= '1';
    layer2_outputs(3031) <= a and not b;
    layer2_outputs(3032) <= b;
    layer2_outputs(3033) <= '1';
    layer2_outputs(3034) <= a or b;
    layer2_outputs(3035) <= '1';
    layer2_outputs(3036) <= a;
    layer2_outputs(3037) <= b;
    layer2_outputs(3038) <= b;
    layer2_outputs(3039) <= not (a or b);
    layer2_outputs(3040) <= not (a or b);
    layer2_outputs(3041) <= not (a and b);
    layer2_outputs(3042) <= not (a and b);
    layer2_outputs(3043) <= a or b;
    layer2_outputs(3044) <= a and b;
    layer2_outputs(3045) <= a;
    layer2_outputs(3046) <= b;
    layer2_outputs(3047) <= not b;
    layer2_outputs(3048) <= not b or a;
    layer2_outputs(3049) <= not (a or b);
    layer2_outputs(3050) <= a and b;
    layer2_outputs(3051) <= a;
    layer2_outputs(3052) <= b;
    layer2_outputs(3053) <= not b;
    layer2_outputs(3054) <= not a or b;
    layer2_outputs(3055) <= b and not a;
    layer2_outputs(3056) <= not a;
    layer2_outputs(3057) <= not a;
    layer2_outputs(3058) <= a and b;
    layer2_outputs(3059) <= not (a xor b);
    layer2_outputs(3060) <= not a or b;
    layer2_outputs(3061) <= not a;
    layer2_outputs(3062) <= a xor b;
    layer2_outputs(3063) <= a and not b;
    layer2_outputs(3064) <= '0';
    layer2_outputs(3065) <= not a;
    layer2_outputs(3066) <= not (a or b);
    layer2_outputs(3067) <= not (a or b);
    layer2_outputs(3068) <= b and not a;
    layer2_outputs(3069) <= not b or a;
    layer2_outputs(3070) <= not b;
    layer2_outputs(3071) <= not (a and b);
    layer2_outputs(3072) <= not (a or b);
    layer2_outputs(3073) <= not (a and b);
    layer2_outputs(3074) <= not b or a;
    layer2_outputs(3075) <= a;
    layer2_outputs(3076) <= not (a and b);
    layer2_outputs(3077) <= not (a or b);
    layer2_outputs(3078) <= not b or a;
    layer2_outputs(3079) <= not a;
    layer2_outputs(3080) <= '0';
    layer2_outputs(3081) <= not a;
    layer2_outputs(3082) <= a;
    layer2_outputs(3083) <= '1';
    layer2_outputs(3084) <= '0';
    layer2_outputs(3085) <= not b or a;
    layer2_outputs(3086) <= a xor b;
    layer2_outputs(3087) <= not (a xor b);
    layer2_outputs(3088) <= not a;
    layer2_outputs(3089) <= not b;
    layer2_outputs(3090) <= a and not b;
    layer2_outputs(3091) <= b and not a;
    layer2_outputs(3092) <= '0';
    layer2_outputs(3093) <= b and not a;
    layer2_outputs(3094) <= b;
    layer2_outputs(3095) <= '0';
    layer2_outputs(3096) <= a or b;
    layer2_outputs(3097) <= not b or a;
    layer2_outputs(3098) <= not (a or b);
    layer2_outputs(3099) <= not a;
    layer2_outputs(3100) <= a or b;
    layer2_outputs(3101) <= not (a or b);
    layer2_outputs(3102) <= a and b;
    layer2_outputs(3103) <= b;
    layer2_outputs(3104) <= not (a and b);
    layer2_outputs(3105) <= b and not a;
    layer2_outputs(3106) <= b;
    layer2_outputs(3107) <= b and not a;
    layer2_outputs(3108) <= not a;
    layer2_outputs(3109) <= a xor b;
    layer2_outputs(3110) <= a;
    layer2_outputs(3111) <= not a;
    layer2_outputs(3112) <= b and not a;
    layer2_outputs(3113) <= not b;
    layer2_outputs(3114) <= not (a or b);
    layer2_outputs(3115) <= a;
    layer2_outputs(3116) <= not (a and b);
    layer2_outputs(3117) <= not a;
    layer2_outputs(3118) <= not a;
    layer2_outputs(3119) <= '0';
    layer2_outputs(3120) <= a and b;
    layer2_outputs(3121) <= not a or b;
    layer2_outputs(3122) <= b and not a;
    layer2_outputs(3123) <= a or b;
    layer2_outputs(3124) <= '0';
    layer2_outputs(3125) <= not (a and b);
    layer2_outputs(3126) <= a;
    layer2_outputs(3127) <= a;
    layer2_outputs(3128) <= a and not b;
    layer2_outputs(3129) <= a or b;
    layer2_outputs(3130) <= a or b;
    layer2_outputs(3131) <= a and not b;
    layer2_outputs(3132) <= a and b;
    layer2_outputs(3133) <= a;
    layer2_outputs(3134) <= not b;
    layer2_outputs(3135) <= a;
    layer2_outputs(3136) <= not a;
    layer2_outputs(3137) <= b;
    layer2_outputs(3138) <= '0';
    layer2_outputs(3139) <= a and not b;
    layer2_outputs(3140) <= not b;
    layer2_outputs(3141) <= not (a or b);
    layer2_outputs(3142) <= a and not b;
    layer2_outputs(3143) <= a and b;
    layer2_outputs(3144) <= not b or a;
    layer2_outputs(3145) <= not a or b;
    layer2_outputs(3146) <= not (a or b);
    layer2_outputs(3147) <= not a or b;
    layer2_outputs(3148) <= not b;
    layer2_outputs(3149) <= a or b;
    layer2_outputs(3150) <= a or b;
    layer2_outputs(3151) <= not (a or b);
    layer2_outputs(3152) <= not (a or b);
    layer2_outputs(3153) <= not b;
    layer2_outputs(3154) <= a;
    layer2_outputs(3155) <= b and not a;
    layer2_outputs(3156) <= not b;
    layer2_outputs(3157) <= b;
    layer2_outputs(3158) <= '1';
    layer2_outputs(3159) <= not (a or b);
    layer2_outputs(3160) <= '0';
    layer2_outputs(3161) <= not b or a;
    layer2_outputs(3162) <= '1';
    layer2_outputs(3163) <= not a;
    layer2_outputs(3164) <= a xor b;
    layer2_outputs(3165) <= not b;
    layer2_outputs(3166) <= a and not b;
    layer2_outputs(3167) <= not b or a;
    layer2_outputs(3168) <= b;
    layer2_outputs(3169) <= b and not a;
    layer2_outputs(3170) <= not (a and b);
    layer2_outputs(3171) <= '0';
    layer2_outputs(3172) <= b;
    layer2_outputs(3173) <= not (a and b);
    layer2_outputs(3174) <= a and not b;
    layer2_outputs(3175) <= not a;
    layer2_outputs(3176) <= b and not a;
    layer2_outputs(3177) <= not a or b;
    layer2_outputs(3178) <= a and not b;
    layer2_outputs(3179) <= not (a and b);
    layer2_outputs(3180) <= not a;
    layer2_outputs(3181) <= a and b;
    layer2_outputs(3182) <= not (a and b);
    layer2_outputs(3183) <= '1';
    layer2_outputs(3184) <= a;
    layer2_outputs(3185) <= not b or a;
    layer2_outputs(3186) <= a or b;
    layer2_outputs(3187) <= a and b;
    layer2_outputs(3188) <= not (a or b);
    layer2_outputs(3189) <= b and not a;
    layer2_outputs(3190) <= a or b;
    layer2_outputs(3191) <= b and not a;
    layer2_outputs(3192) <= '1';
    layer2_outputs(3193) <= a or b;
    layer2_outputs(3194) <= b;
    layer2_outputs(3195) <= a and not b;
    layer2_outputs(3196) <= not (a or b);
    layer2_outputs(3197) <= '0';
    layer2_outputs(3198) <= b;
    layer2_outputs(3199) <= '1';
    layer2_outputs(3200) <= not b or a;
    layer2_outputs(3201) <= a;
    layer2_outputs(3202) <= b and not a;
    layer2_outputs(3203) <= not (a xor b);
    layer2_outputs(3204) <= b and not a;
    layer2_outputs(3205) <= not (a xor b);
    layer2_outputs(3206) <= not b;
    layer2_outputs(3207) <= '0';
    layer2_outputs(3208) <= not b;
    layer2_outputs(3209) <= a and not b;
    layer2_outputs(3210) <= b and not a;
    layer2_outputs(3211) <= not (a and b);
    layer2_outputs(3212) <= not b or a;
    layer2_outputs(3213) <= '1';
    layer2_outputs(3214) <= not b;
    layer2_outputs(3215) <= '0';
    layer2_outputs(3216) <= b;
    layer2_outputs(3217) <= b;
    layer2_outputs(3218) <= a and not b;
    layer2_outputs(3219) <= not b;
    layer2_outputs(3220) <= not (a and b);
    layer2_outputs(3221) <= a and not b;
    layer2_outputs(3222) <= a xor b;
    layer2_outputs(3223) <= '1';
    layer2_outputs(3224) <= not a or b;
    layer2_outputs(3225) <= '0';
    layer2_outputs(3226) <= a or b;
    layer2_outputs(3227) <= a;
    layer2_outputs(3228) <= a;
    layer2_outputs(3229) <= '1';
    layer2_outputs(3230) <= a or b;
    layer2_outputs(3231) <= not (a xor b);
    layer2_outputs(3232) <= not (a or b);
    layer2_outputs(3233) <= a;
    layer2_outputs(3234) <= not (a or b);
    layer2_outputs(3235) <= '0';
    layer2_outputs(3236) <= '1';
    layer2_outputs(3237) <= not a;
    layer2_outputs(3238) <= a and b;
    layer2_outputs(3239) <= '0';
    layer2_outputs(3240) <= not b or a;
    layer2_outputs(3241) <= not (a or b);
    layer2_outputs(3242) <= b;
    layer2_outputs(3243) <= not a;
    layer2_outputs(3244) <= '0';
    layer2_outputs(3245) <= not (a and b);
    layer2_outputs(3246) <= a and b;
    layer2_outputs(3247) <= not (a xor b);
    layer2_outputs(3248) <= not (a or b);
    layer2_outputs(3249) <= b;
    layer2_outputs(3250) <= a xor b;
    layer2_outputs(3251) <= a and b;
    layer2_outputs(3252) <= b and not a;
    layer2_outputs(3253) <= a or b;
    layer2_outputs(3254) <= a xor b;
    layer2_outputs(3255) <= b;
    layer2_outputs(3256) <= b;
    layer2_outputs(3257) <= b;
    layer2_outputs(3258) <= b and not a;
    layer2_outputs(3259) <= a;
    layer2_outputs(3260) <= b;
    layer2_outputs(3261) <= not a or b;
    layer2_outputs(3262) <= not a or b;
    layer2_outputs(3263) <= a or b;
    layer2_outputs(3264) <= not (a and b);
    layer2_outputs(3265) <= a;
    layer2_outputs(3266) <= a or b;
    layer2_outputs(3267) <= a and b;
    layer2_outputs(3268) <= a and b;
    layer2_outputs(3269) <= not (a or b);
    layer2_outputs(3270) <= b and not a;
    layer2_outputs(3271) <= not (a or b);
    layer2_outputs(3272) <= not b;
    layer2_outputs(3273) <= '0';
    layer2_outputs(3274) <= a and b;
    layer2_outputs(3275) <= not b;
    layer2_outputs(3276) <= b;
    layer2_outputs(3277) <= not a;
    layer2_outputs(3278) <= a and b;
    layer2_outputs(3279) <= '0';
    layer2_outputs(3280) <= '1';
    layer2_outputs(3281) <= b;
    layer2_outputs(3282) <= a;
    layer2_outputs(3283) <= not a;
    layer2_outputs(3284) <= not (a and b);
    layer2_outputs(3285) <= not b;
    layer2_outputs(3286) <= a;
    layer2_outputs(3287) <= a xor b;
    layer2_outputs(3288) <= b;
    layer2_outputs(3289) <= not b or a;
    layer2_outputs(3290) <= not (a and b);
    layer2_outputs(3291) <= not b or a;
    layer2_outputs(3292) <= not b;
    layer2_outputs(3293) <= '0';
    layer2_outputs(3294) <= not b;
    layer2_outputs(3295) <= not (a or b);
    layer2_outputs(3296) <= not b;
    layer2_outputs(3297) <= '1';
    layer2_outputs(3298) <= a;
    layer2_outputs(3299) <= a or b;
    layer2_outputs(3300) <= not (a xor b);
    layer2_outputs(3301) <= '1';
    layer2_outputs(3302) <= a;
    layer2_outputs(3303) <= a and not b;
    layer2_outputs(3304) <= not (a xor b);
    layer2_outputs(3305) <= b;
    layer2_outputs(3306) <= not (a and b);
    layer2_outputs(3307) <= not a or b;
    layer2_outputs(3308) <= not b;
    layer2_outputs(3309) <= a xor b;
    layer2_outputs(3310) <= a and not b;
    layer2_outputs(3311) <= not (a and b);
    layer2_outputs(3312) <= not a;
    layer2_outputs(3313) <= b;
    layer2_outputs(3314) <= a or b;
    layer2_outputs(3315) <= not (a and b);
    layer2_outputs(3316) <= not (a and b);
    layer2_outputs(3317) <= not b;
    layer2_outputs(3318) <= not a;
    layer2_outputs(3319) <= not b or a;
    layer2_outputs(3320) <= a;
    layer2_outputs(3321) <= not a or b;
    layer2_outputs(3322) <= '0';
    layer2_outputs(3323) <= not b;
    layer2_outputs(3324) <= a or b;
    layer2_outputs(3325) <= not b or a;
    layer2_outputs(3326) <= not a or b;
    layer2_outputs(3327) <= not (a and b);
    layer2_outputs(3328) <= '1';
    layer2_outputs(3329) <= a and not b;
    layer2_outputs(3330) <= not b or a;
    layer2_outputs(3331) <= b;
    layer2_outputs(3332) <= a xor b;
    layer2_outputs(3333) <= '1';
    layer2_outputs(3334) <= not (a and b);
    layer2_outputs(3335) <= '1';
    layer2_outputs(3336) <= not (a xor b);
    layer2_outputs(3337) <= not (a and b);
    layer2_outputs(3338) <= a;
    layer2_outputs(3339) <= b and not a;
    layer2_outputs(3340) <= '0';
    layer2_outputs(3341) <= not b;
    layer2_outputs(3342) <= not b or a;
    layer2_outputs(3343) <= a or b;
    layer2_outputs(3344) <= not a or b;
    layer2_outputs(3345) <= '0';
    layer2_outputs(3346) <= a or b;
    layer2_outputs(3347) <= b and not a;
    layer2_outputs(3348) <= not (a xor b);
    layer2_outputs(3349) <= '0';
    layer2_outputs(3350) <= a or b;
    layer2_outputs(3351) <= b and not a;
    layer2_outputs(3352) <= a;
    layer2_outputs(3353) <= a and not b;
    layer2_outputs(3354) <= b;
    layer2_outputs(3355) <= a xor b;
    layer2_outputs(3356) <= a xor b;
    layer2_outputs(3357) <= not b;
    layer2_outputs(3358) <= not b or a;
    layer2_outputs(3359) <= not a;
    layer2_outputs(3360) <= not a or b;
    layer2_outputs(3361) <= '0';
    layer2_outputs(3362) <= a;
    layer2_outputs(3363) <= not a or b;
    layer2_outputs(3364) <= b;
    layer2_outputs(3365) <= b and not a;
    layer2_outputs(3366) <= a and not b;
    layer2_outputs(3367) <= '0';
    layer2_outputs(3368) <= b;
    layer2_outputs(3369) <= not a;
    layer2_outputs(3370) <= not (a or b);
    layer2_outputs(3371) <= a;
    layer2_outputs(3372) <= b and not a;
    layer2_outputs(3373) <= a and not b;
    layer2_outputs(3374) <= b and not a;
    layer2_outputs(3375) <= not b;
    layer2_outputs(3376) <= a xor b;
    layer2_outputs(3377) <= not a;
    layer2_outputs(3378) <= a;
    layer2_outputs(3379) <= a and b;
    layer2_outputs(3380) <= a and not b;
    layer2_outputs(3381) <= '1';
    layer2_outputs(3382) <= not b or a;
    layer2_outputs(3383) <= not a;
    layer2_outputs(3384) <= not (a xor b);
    layer2_outputs(3385) <= a xor b;
    layer2_outputs(3386) <= '0';
    layer2_outputs(3387) <= not a or b;
    layer2_outputs(3388) <= not b;
    layer2_outputs(3389) <= not a or b;
    layer2_outputs(3390) <= a and b;
    layer2_outputs(3391) <= not a;
    layer2_outputs(3392) <= a and not b;
    layer2_outputs(3393) <= not b or a;
    layer2_outputs(3394) <= '1';
    layer2_outputs(3395) <= not (a or b);
    layer2_outputs(3396) <= a xor b;
    layer2_outputs(3397) <= a xor b;
    layer2_outputs(3398) <= a xor b;
    layer2_outputs(3399) <= a and not b;
    layer2_outputs(3400) <= b;
    layer2_outputs(3401) <= not b;
    layer2_outputs(3402) <= not (a and b);
    layer2_outputs(3403) <= not (a and b);
    layer2_outputs(3404) <= a xor b;
    layer2_outputs(3405) <= not (a and b);
    layer2_outputs(3406) <= not a or b;
    layer2_outputs(3407) <= b;
    layer2_outputs(3408) <= not b;
    layer2_outputs(3409) <= not b;
    layer2_outputs(3410) <= not a;
    layer2_outputs(3411) <= b and not a;
    layer2_outputs(3412) <= '1';
    layer2_outputs(3413) <= a and b;
    layer2_outputs(3414) <= '0';
    layer2_outputs(3415) <= a and b;
    layer2_outputs(3416) <= not (a or b);
    layer2_outputs(3417) <= b;
    layer2_outputs(3418) <= not (a and b);
    layer2_outputs(3419) <= '1';
    layer2_outputs(3420) <= b;
    layer2_outputs(3421) <= b;
    layer2_outputs(3422) <= a and b;
    layer2_outputs(3423) <= b;
    layer2_outputs(3424) <= not a;
    layer2_outputs(3425) <= not a;
    layer2_outputs(3426) <= b;
    layer2_outputs(3427) <= not b;
    layer2_outputs(3428) <= b and not a;
    layer2_outputs(3429) <= not (a or b);
    layer2_outputs(3430) <= not a;
    layer2_outputs(3431) <= a;
    layer2_outputs(3432) <= not (a and b);
    layer2_outputs(3433) <= not (a xor b);
    layer2_outputs(3434) <= not b or a;
    layer2_outputs(3435) <= a;
    layer2_outputs(3436) <= not (a and b);
    layer2_outputs(3437) <= '1';
    layer2_outputs(3438) <= not a or b;
    layer2_outputs(3439) <= not b;
    layer2_outputs(3440) <= a or b;
    layer2_outputs(3441) <= not b;
    layer2_outputs(3442) <= not (a and b);
    layer2_outputs(3443) <= '0';
    layer2_outputs(3444) <= not (a or b);
    layer2_outputs(3445) <= a and b;
    layer2_outputs(3446) <= '1';
    layer2_outputs(3447) <= a and b;
    layer2_outputs(3448) <= a and not b;
    layer2_outputs(3449) <= not b;
    layer2_outputs(3450) <= a or b;
    layer2_outputs(3451) <= b;
    layer2_outputs(3452) <= not a or b;
    layer2_outputs(3453) <= not a or b;
    layer2_outputs(3454) <= not (a xor b);
    layer2_outputs(3455) <= not b;
    layer2_outputs(3456) <= not (a and b);
    layer2_outputs(3457) <= not a;
    layer2_outputs(3458) <= b;
    layer2_outputs(3459) <= not (a and b);
    layer2_outputs(3460) <= not (a xor b);
    layer2_outputs(3461) <= a and b;
    layer2_outputs(3462) <= not a;
    layer2_outputs(3463) <= a or b;
    layer2_outputs(3464) <= not b;
    layer2_outputs(3465) <= a and not b;
    layer2_outputs(3466) <= '1';
    layer2_outputs(3467) <= a and not b;
    layer2_outputs(3468) <= not a or b;
    layer2_outputs(3469) <= not (a and b);
    layer2_outputs(3470) <= '1';
    layer2_outputs(3471) <= a;
    layer2_outputs(3472) <= not (a and b);
    layer2_outputs(3473) <= a or b;
    layer2_outputs(3474) <= '1';
    layer2_outputs(3475) <= not a;
    layer2_outputs(3476) <= not (a and b);
    layer2_outputs(3477) <= a and not b;
    layer2_outputs(3478) <= a;
    layer2_outputs(3479) <= b and not a;
    layer2_outputs(3480) <= '1';
    layer2_outputs(3481) <= '0';
    layer2_outputs(3482) <= a and b;
    layer2_outputs(3483) <= '1';
    layer2_outputs(3484) <= b and not a;
    layer2_outputs(3485) <= not a;
    layer2_outputs(3486) <= a xor b;
    layer2_outputs(3487) <= a and b;
    layer2_outputs(3488) <= b;
    layer2_outputs(3489) <= not (a or b);
    layer2_outputs(3490) <= not a;
    layer2_outputs(3491) <= '0';
    layer2_outputs(3492) <= not b;
    layer2_outputs(3493) <= not (a or b);
    layer2_outputs(3494) <= '1';
    layer2_outputs(3495) <= a xor b;
    layer2_outputs(3496) <= not b;
    layer2_outputs(3497) <= not b or a;
    layer2_outputs(3498) <= not a;
    layer2_outputs(3499) <= b;
    layer2_outputs(3500) <= a or b;
    layer2_outputs(3501) <= a;
    layer2_outputs(3502) <= b;
    layer2_outputs(3503) <= not b;
    layer2_outputs(3504) <= b and not a;
    layer2_outputs(3505) <= not a;
    layer2_outputs(3506) <= '1';
    layer2_outputs(3507) <= b;
    layer2_outputs(3508) <= a and not b;
    layer2_outputs(3509) <= not a or b;
    layer2_outputs(3510) <= b;
    layer2_outputs(3511) <= a;
    layer2_outputs(3512) <= a or b;
    layer2_outputs(3513) <= not a or b;
    layer2_outputs(3514) <= not a;
    layer2_outputs(3515) <= not a;
    layer2_outputs(3516) <= not b;
    layer2_outputs(3517) <= a and not b;
    layer2_outputs(3518) <= not (a or b);
    layer2_outputs(3519) <= not a;
    layer2_outputs(3520) <= '0';
    layer2_outputs(3521) <= a;
    layer2_outputs(3522) <= not a or b;
    layer2_outputs(3523) <= b and not a;
    layer2_outputs(3524) <= a and not b;
    layer2_outputs(3525) <= a;
    layer2_outputs(3526) <= a and b;
    layer2_outputs(3527) <= not (a or b);
    layer2_outputs(3528) <= not a or b;
    layer2_outputs(3529) <= not (a or b);
    layer2_outputs(3530) <= not a or b;
    layer2_outputs(3531) <= b;
    layer2_outputs(3532) <= not b or a;
    layer2_outputs(3533) <= b;
    layer2_outputs(3534) <= a or b;
    layer2_outputs(3535) <= not b;
    layer2_outputs(3536) <= not b or a;
    layer2_outputs(3537) <= '0';
    layer2_outputs(3538) <= a and not b;
    layer2_outputs(3539) <= a and b;
    layer2_outputs(3540) <= not (a xor b);
    layer2_outputs(3541) <= b and not a;
    layer2_outputs(3542) <= a or b;
    layer2_outputs(3543) <= not b or a;
    layer2_outputs(3544) <= not b;
    layer2_outputs(3545) <= not (a or b);
    layer2_outputs(3546) <= b and not a;
    layer2_outputs(3547) <= not (a and b);
    layer2_outputs(3548) <= a;
    layer2_outputs(3549) <= a and not b;
    layer2_outputs(3550) <= not (a or b);
    layer2_outputs(3551) <= b and not a;
    layer2_outputs(3552) <= not b;
    layer2_outputs(3553) <= a;
    layer2_outputs(3554) <= a;
    layer2_outputs(3555) <= not b;
    layer2_outputs(3556) <= a and not b;
    layer2_outputs(3557) <= b;
    layer2_outputs(3558) <= not b or a;
    layer2_outputs(3559) <= a and b;
    layer2_outputs(3560) <= b and not a;
    layer2_outputs(3561) <= not (a or b);
    layer2_outputs(3562) <= b and not a;
    layer2_outputs(3563) <= a or b;
    layer2_outputs(3564) <= not a or b;
    layer2_outputs(3565) <= not b;
    layer2_outputs(3566) <= a and not b;
    layer2_outputs(3567) <= b and not a;
    layer2_outputs(3568) <= not b;
    layer2_outputs(3569) <= a xor b;
    layer2_outputs(3570) <= a or b;
    layer2_outputs(3571) <= not (a and b);
    layer2_outputs(3572) <= b;
    layer2_outputs(3573) <= a or b;
    layer2_outputs(3574) <= b and not a;
    layer2_outputs(3575) <= a;
    layer2_outputs(3576) <= b;
    layer2_outputs(3577) <= not b or a;
    layer2_outputs(3578) <= a or b;
    layer2_outputs(3579) <= '0';
    layer2_outputs(3580) <= not b;
    layer2_outputs(3581) <= not b or a;
    layer2_outputs(3582) <= not a;
    layer2_outputs(3583) <= not (a and b);
    layer2_outputs(3584) <= a;
    layer2_outputs(3585) <= not (a and b);
    layer2_outputs(3586) <= b;
    layer2_outputs(3587) <= a and b;
    layer2_outputs(3588) <= a and not b;
    layer2_outputs(3589) <= not a or b;
    layer2_outputs(3590) <= not (a and b);
    layer2_outputs(3591) <= not a or b;
    layer2_outputs(3592) <= not a or b;
    layer2_outputs(3593) <= not (a and b);
    layer2_outputs(3594) <= a or b;
    layer2_outputs(3595) <= not b;
    layer2_outputs(3596) <= not (a xor b);
    layer2_outputs(3597) <= not b;
    layer2_outputs(3598) <= not a or b;
    layer2_outputs(3599) <= b;
    layer2_outputs(3600) <= not a or b;
    layer2_outputs(3601) <= '1';
    layer2_outputs(3602) <= not b or a;
    layer2_outputs(3603) <= a and b;
    layer2_outputs(3604) <= not a or b;
    layer2_outputs(3605) <= a and b;
    layer2_outputs(3606) <= not b or a;
    layer2_outputs(3607) <= a and b;
    layer2_outputs(3608) <= not b or a;
    layer2_outputs(3609) <= b and not a;
    layer2_outputs(3610) <= '0';
    layer2_outputs(3611) <= b;
    layer2_outputs(3612) <= '1';
    layer2_outputs(3613) <= b and not a;
    layer2_outputs(3614) <= a or b;
    layer2_outputs(3615) <= not (a or b);
    layer2_outputs(3616) <= not a;
    layer2_outputs(3617) <= a;
    layer2_outputs(3618) <= not a;
    layer2_outputs(3619) <= a;
    layer2_outputs(3620) <= a;
    layer2_outputs(3621) <= b;
    layer2_outputs(3622) <= not (a and b);
    layer2_outputs(3623) <= a and not b;
    layer2_outputs(3624) <= not a;
    layer2_outputs(3625) <= not b;
    layer2_outputs(3626) <= b;
    layer2_outputs(3627) <= '0';
    layer2_outputs(3628) <= not a or b;
    layer2_outputs(3629) <= b and not a;
    layer2_outputs(3630) <= a or b;
    layer2_outputs(3631) <= not (a xor b);
    layer2_outputs(3632) <= not (a or b);
    layer2_outputs(3633) <= a and not b;
    layer2_outputs(3634) <= a and not b;
    layer2_outputs(3635) <= not a;
    layer2_outputs(3636) <= b and not a;
    layer2_outputs(3637) <= '0';
    layer2_outputs(3638) <= a;
    layer2_outputs(3639) <= b and not a;
    layer2_outputs(3640) <= '1';
    layer2_outputs(3641) <= not a or b;
    layer2_outputs(3642) <= not b or a;
    layer2_outputs(3643) <= not (a or b);
    layer2_outputs(3644) <= b;
    layer2_outputs(3645) <= a or b;
    layer2_outputs(3646) <= not b;
    layer2_outputs(3647) <= b;
    layer2_outputs(3648) <= not (a or b);
    layer2_outputs(3649) <= not a or b;
    layer2_outputs(3650) <= a and not b;
    layer2_outputs(3651) <= not b;
    layer2_outputs(3652) <= not (a and b);
    layer2_outputs(3653) <= a and not b;
    layer2_outputs(3654) <= a or b;
    layer2_outputs(3655) <= not b or a;
    layer2_outputs(3656) <= not b;
    layer2_outputs(3657) <= not (a or b);
    layer2_outputs(3658) <= not (a or b);
    layer2_outputs(3659) <= b;
    layer2_outputs(3660) <= not a;
    layer2_outputs(3661) <= '0';
    layer2_outputs(3662) <= not (a or b);
    layer2_outputs(3663) <= a or b;
    layer2_outputs(3664) <= not a or b;
    layer2_outputs(3665) <= not a;
    layer2_outputs(3666) <= a and b;
    layer2_outputs(3667) <= not a or b;
    layer2_outputs(3668) <= not (a and b);
    layer2_outputs(3669) <= b;
    layer2_outputs(3670) <= a and not b;
    layer2_outputs(3671) <= a and b;
    layer2_outputs(3672) <= a xor b;
    layer2_outputs(3673) <= b;
    layer2_outputs(3674) <= not b;
    layer2_outputs(3675) <= a;
    layer2_outputs(3676) <= '1';
    layer2_outputs(3677) <= not a or b;
    layer2_outputs(3678) <= a and not b;
    layer2_outputs(3679) <= b;
    layer2_outputs(3680) <= a and not b;
    layer2_outputs(3681) <= a and not b;
    layer2_outputs(3682) <= not b or a;
    layer2_outputs(3683) <= b and not a;
    layer2_outputs(3684) <= b;
    layer2_outputs(3685) <= b and not a;
    layer2_outputs(3686) <= a and not b;
    layer2_outputs(3687) <= a and not b;
    layer2_outputs(3688) <= a xor b;
    layer2_outputs(3689) <= not (a and b);
    layer2_outputs(3690) <= a and not b;
    layer2_outputs(3691) <= not a or b;
    layer2_outputs(3692) <= a and not b;
    layer2_outputs(3693) <= a xor b;
    layer2_outputs(3694) <= b;
    layer2_outputs(3695) <= a and b;
    layer2_outputs(3696) <= not (a or b);
    layer2_outputs(3697) <= a xor b;
    layer2_outputs(3698) <= a;
    layer2_outputs(3699) <= not b;
    layer2_outputs(3700) <= not a;
    layer2_outputs(3701) <= not (a or b);
    layer2_outputs(3702) <= a or b;
    layer2_outputs(3703) <= a or b;
    layer2_outputs(3704) <= not (a or b);
    layer2_outputs(3705) <= '1';
    layer2_outputs(3706) <= b;
    layer2_outputs(3707) <= a and b;
    layer2_outputs(3708) <= a and not b;
    layer2_outputs(3709) <= '1';
    layer2_outputs(3710) <= not (a and b);
    layer2_outputs(3711) <= a;
    layer2_outputs(3712) <= not b;
    layer2_outputs(3713) <= b;
    layer2_outputs(3714) <= not b;
    layer2_outputs(3715) <= a and not b;
    layer2_outputs(3716) <= b and not a;
    layer2_outputs(3717) <= not a;
    layer2_outputs(3718) <= '0';
    layer2_outputs(3719) <= b;
    layer2_outputs(3720) <= a or b;
    layer2_outputs(3721) <= not (a or b);
    layer2_outputs(3722) <= b and not a;
    layer2_outputs(3723) <= not b or a;
    layer2_outputs(3724) <= a and not b;
    layer2_outputs(3725) <= not (a and b);
    layer2_outputs(3726) <= a and b;
    layer2_outputs(3727) <= not (a or b);
    layer2_outputs(3728) <= not a;
    layer2_outputs(3729) <= not b;
    layer2_outputs(3730) <= a and not b;
    layer2_outputs(3731) <= a;
    layer2_outputs(3732) <= b and not a;
    layer2_outputs(3733) <= not (a and b);
    layer2_outputs(3734) <= not b;
    layer2_outputs(3735) <= not a;
    layer2_outputs(3736) <= b and not a;
    layer2_outputs(3737) <= b;
    layer2_outputs(3738) <= not b;
    layer2_outputs(3739) <= b and not a;
    layer2_outputs(3740) <= a and not b;
    layer2_outputs(3741) <= a or b;
    layer2_outputs(3742) <= not b;
    layer2_outputs(3743) <= not b;
    layer2_outputs(3744) <= not (a and b);
    layer2_outputs(3745) <= not b;
    layer2_outputs(3746) <= not b;
    layer2_outputs(3747) <= a and not b;
    layer2_outputs(3748) <= not a;
    layer2_outputs(3749) <= b and not a;
    layer2_outputs(3750) <= not (a or b);
    layer2_outputs(3751) <= not (a or b);
    layer2_outputs(3752) <= b;
    layer2_outputs(3753) <= b;
    layer2_outputs(3754) <= not a;
    layer2_outputs(3755) <= a;
    layer2_outputs(3756) <= not b;
    layer2_outputs(3757) <= not a or b;
    layer2_outputs(3758) <= not a;
    layer2_outputs(3759) <= '0';
    layer2_outputs(3760) <= b and not a;
    layer2_outputs(3761) <= '1';
    layer2_outputs(3762) <= a and not b;
    layer2_outputs(3763) <= b;
    layer2_outputs(3764) <= b;
    layer2_outputs(3765) <= a and b;
    layer2_outputs(3766) <= not b;
    layer2_outputs(3767) <= a;
    layer2_outputs(3768) <= b and not a;
    layer2_outputs(3769) <= '1';
    layer2_outputs(3770) <= b;
    layer2_outputs(3771) <= b;
    layer2_outputs(3772) <= not a or b;
    layer2_outputs(3773) <= a;
    layer2_outputs(3774) <= not b;
    layer2_outputs(3775) <= not a or b;
    layer2_outputs(3776) <= a and not b;
    layer2_outputs(3777) <= '1';
    layer2_outputs(3778) <= not b;
    layer2_outputs(3779) <= not b;
    layer2_outputs(3780) <= a and b;
    layer2_outputs(3781) <= not (a and b);
    layer2_outputs(3782) <= not (a or b);
    layer2_outputs(3783) <= not a;
    layer2_outputs(3784) <= not b or a;
    layer2_outputs(3785) <= not a;
    layer2_outputs(3786) <= a and b;
    layer2_outputs(3787) <= '1';
    layer2_outputs(3788) <= a and not b;
    layer2_outputs(3789) <= not b or a;
    layer2_outputs(3790) <= '1';
    layer2_outputs(3791) <= a xor b;
    layer2_outputs(3792) <= a;
    layer2_outputs(3793) <= not b;
    layer2_outputs(3794) <= a and b;
    layer2_outputs(3795) <= not (a and b);
    layer2_outputs(3796) <= b and not a;
    layer2_outputs(3797) <= not b;
    layer2_outputs(3798) <= not b;
    layer2_outputs(3799) <= a or b;
    layer2_outputs(3800) <= a;
    layer2_outputs(3801) <= b and not a;
    layer2_outputs(3802) <= a;
    layer2_outputs(3803) <= not b;
    layer2_outputs(3804) <= a and b;
    layer2_outputs(3805) <= not (a and b);
    layer2_outputs(3806) <= '1';
    layer2_outputs(3807) <= not b;
    layer2_outputs(3808) <= b;
    layer2_outputs(3809) <= a and not b;
    layer2_outputs(3810) <= '0';
    layer2_outputs(3811) <= not (a and b);
    layer2_outputs(3812) <= not a;
    layer2_outputs(3813) <= '0';
    layer2_outputs(3814) <= a;
    layer2_outputs(3815) <= not (a and b);
    layer2_outputs(3816) <= a xor b;
    layer2_outputs(3817) <= not b or a;
    layer2_outputs(3818) <= not (a or b);
    layer2_outputs(3819) <= not a;
    layer2_outputs(3820) <= not b;
    layer2_outputs(3821) <= not (a or b);
    layer2_outputs(3822) <= not b or a;
    layer2_outputs(3823) <= a or b;
    layer2_outputs(3824) <= b and not a;
    layer2_outputs(3825) <= not (a or b);
    layer2_outputs(3826) <= b;
    layer2_outputs(3827) <= a and not b;
    layer2_outputs(3828) <= a and not b;
    layer2_outputs(3829) <= a or b;
    layer2_outputs(3830) <= not (a or b);
    layer2_outputs(3831) <= not b or a;
    layer2_outputs(3832) <= b and not a;
    layer2_outputs(3833) <= b;
    layer2_outputs(3834) <= not a;
    layer2_outputs(3835) <= a and not b;
    layer2_outputs(3836) <= not b or a;
    layer2_outputs(3837) <= '1';
    layer2_outputs(3838) <= not (a xor b);
    layer2_outputs(3839) <= b and not a;
    layer2_outputs(3840) <= not b or a;
    layer2_outputs(3841) <= '1';
    layer2_outputs(3842) <= a or b;
    layer2_outputs(3843) <= not (a or b);
    layer2_outputs(3844) <= a xor b;
    layer2_outputs(3845) <= a and not b;
    layer2_outputs(3846) <= not (a and b);
    layer2_outputs(3847) <= a or b;
    layer2_outputs(3848) <= not (a and b);
    layer2_outputs(3849) <= '0';
    layer2_outputs(3850) <= '1';
    layer2_outputs(3851) <= a and not b;
    layer2_outputs(3852) <= a and not b;
    layer2_outputs(3853) <= not a;
    layer2_outputs(3854) <= not (a and b);
    layer2_outputs(3855) <= b and not a;
    layer2_outputs(3856) <= not b;
    layer2_outputs(3857) <= not (a and b);
    layer2_outputs(3858) <= '1';
    layer2_outputs(3859) <= not a;
    layer2_outputs(3860) <= not b;
    layer2_outputs(3861) <= not a;
    layer2_outputs(3862) <= a and not b;
    layer2_outputs(3863) <= a xor b;
    layer2_outputs(3864) <= not a;
    layer2_outputs(3865) <= not a;
    layer2_outputs(3866) <= not (a xor b);
    layer2_outputs(3867) <= not (a and b);
    layer2_outputs(3868) <= not b;
    layer2_outputs(3869) <= not a;
    layer2_outputs(3870) <= a and b;
    layer2_outputs(3871) <= a or b;
    layer2_outputs(3872) <= a;
    layer2_outputs(3873) <= not a or b;
    layer2_outputs(3874) <= not a or b;
    layer2_outputs(3875) <= not a;
    layer2_outputs(3876) <= not b;
    layer2_outputs(3877) <= '1';
    layer2_outputs(3878) <= a and b;
    layer2_outputs(3879) <= a;
    layer2_outputs(3880) <= b;
    layer2_outputs(3881) <= b and not a;
    layer2_outputs(3882) <= not b or a;
    layer2_outputs(3883) <= b;
    layer2_outputs(3884) <= a and not b;
    layer2_outputs(3885) <= not a;
    layer2_outputs(3886) <= not a;
    layer2_outputs(3887) <= a or b;
    layer2_outputs(3888) <= a and not b;
    layer2_outputs(3889) <= '1';
    layer2_outputs(3890) <= b;
    layer2_outputs(3891) <= not (a and b);
    layer2_outputs(3892) <= not b;
    layer2_outputs(3893) <= a or b;
    layer2_outputs(3894) <= a and b;
    layer2_outputs(3895) <= a and not b;
    layer2_outputs(3896) <= a and not b;
    layer2_outputs(3897) <= a;
    layer2_outputs(3898) <= not (a or b);
    layer2_outputs(3899) <= not a;
    layer2_outputs(3900) <= not a or b;
    layer2_outputs(3901) <= b;
    layer2_outputs(3902) <= a and not b;
    layer2_outputs(3903) <= not a;
    layer2_outputs(3904) <= '0';
    layer2_outputs(3905) <= b;
    layer2_outputs(3906) <= b;
    layer2_outputs(3907) <= a and not b;
    layer2_outputs(3908) <= not (a and b);
    layer2_outputs(3909) <= a and not b;
    layer2_outputs(3910) <= a;
    layer2_outputs(3911) <= b;
    layer2_outputs(3912) <= not (a or b);
    layer2_outputs(3913) <= a and b;
    layer2_outputs(3914) <= a;
    layer2_outputs(3915) <= '0';
    layer2_outputs(3916) <= not (a xor b);
    layer2_outputs(3917) <= b and not a;
    layer2_outputs(3918) <= not b or a;
    layer2_outputs(3919) <= a or b;
    layer2_outputs(3920) <= not b or a;
    layer2_outputs(3921) <= not b or a;
    layer2_outputs(3922) <= a;
    layer2_outputs(3923) <= not (a or b);
    layer2_outputs(3924) <= not (a and b);
    layer2_outputs(3925) <= '1';
    layer2_outputs(3926) <= b and not a;
    layer2_outputs(3927) <= a and not b;
    layer2_outputs(3928) <= '0';
    layer2_outputs(3929) <= a;
    layer2_outputs(3930) <= not a;
    layer2_outputs(3931) <= a or b;
    layer2_outputs(3932) <= not a;
    layer2_outputs(3933) <= not b;
    layer2_outputs(3934) <= a and not b;
    layer2_outputs(3935) <= not (a or b);
    layer2_outputs(3936) <= not (a or b);
    layer2_outputs(3937) <= not a;
    layer2_outputs(3938) <= a and not b;
    layer2_outputs(3939) <= b and not a;
    layer2_outputs(3940) <= b;
    layer2_outputs(3941) <= not b;
    layer2_outputs(3942) <= not (a and b);
    layer2_outputs(3943) <= not b;
    layer2_outputs(3944) <= a or b;
    layer2_outputs(3945) <= b and not a;
    layer2_outputs(3946) <= a;
    layer2_outputs(3947) <= a and not b;
    layer2_outputs(3948) <= a;
    layer2_outputs(3949) <= not (a xor b);
    layer2_outputs(3950) <= a and not b;
    layer2_outputs(3951) <= b;
    layer2_outputs(3952) <= a;
    layer2_outputs(3953) <= a;
    layer2_outputs(3954) <= a xor b;
    layer2_outputs(3955) <= a and not b;
    layer2_outputs(3956) <= not b;
    layer2_outputs(3957) <= not a;
    layer2_outputs(3958) <= a;
    layer2_outputs(3959) <= not a;
    layer2_outputs(3960) <= b;
    layer2_outputs(3961) <= a xor b;
    layer2_outputs(3962) <= not a;
    layer2_outputs(3963) <= not b or a;
    layer2_outputs(3964) <= not a or b;
    layer2_outputs(3965) <= not b;
    layer2_outputs(3966) <= a;
    layer2_outputs(3967) <= not (a or b);
    layer2_outputs(3968) <= not b or a;
    layer2_outputs(3969) <= not (a and b);
    layer2_outputs(3970) <= a and not b;
    layer2_outputs(3971) <= a or b;
    layer2_outputs(3972) <= not (a or b);
    layer2_outputs(3973) <= not (a or b);
    layer2_outputs(3974) <= b and not a;
    layer2_outputs(3975) <= a;
    layer2_outputs(3976) <= '0';
    layer2_outputs(3977) <= not (a xor b);
    layer2_outputs(3978) <= a;
    layer2_outputs(3979) <= b and not a;
    layer2_outputs(3980) <= not (a xor b);
    layer2_outputs(3981) <= not (a or b);
    layer2_outputs(3982) <= '1';
    layer2_outputs(3983) <= not a;
    layer2_outputs(3984) <= not a or b;
    layer2_outputs(3985) <= b and not a;
    layer2_outputs(3986) <= a and not b;
    layer2_outputs(3987) <= a xor b;
    layer2_outputs(3988) <= a or b;
    layer2_outputs(3989) <= a and not b;
    layer2_outputs(3990) <= not a or b;
    layer2_outputs(3991) <= '1';
    layer2_outputs(3992) <= b;
    layer2_outputs(3993) <= a xor b;
    layer2_outputs(3994) <= not (a xor b);
    layer2_outputs(3995) <= not b or a;
    layer2_outputs(3996) <= '0';
    layer2_outputs(3997) <= a and not b;
    layer2_outputs(3998) <= not a;
    layer2_outputs(3999) <= not a;
    layer2_outputs(4000) <= not (a and b);
    layer2_outputs(4001) <= b;
    layer2_outputs(4002) <= not a;
    layer2_outputs(4003) <= not b;
    layer2_outputs(4004) <= b;
    layer2_outputs(4005) <= not b or a;
    layer2_outputs(4006) <= a and b;
    layer2_outputs(4007) <= not (a or b);
    layer2_outputs(4008) <= a;
    layer2_outputs(4009) <= not (a or b);
    layer2_outputs(4010) <= a xor b;
    layer2_outputs(4011) <= a;
    layer2_outputs(4012) <= a and not b;
    layer2_outputs(4013) <= a or b;
    layer2_outputs(4014) <= not b;
    layer2_outputs(4015) <= b and not a;
    layer2_outputs(4016) <= not (a or b);
    layer2_outputs(4017) <= not b or a;
    layer2_outputs(4018) <= b;
    layer2_outputs(4019) <= not (a or b);
    layer2_outputs(4020) <= not (a xor b);
    layer2_outputs(4021) <= a and b;
    layer2_outputs(4022) <= not (a and b);
    layer2_outputs(4023) <= not a;
    layer2_outputs(4024) <= b and not a;
    layer2_outputs(4025) <= not (a and b);
    layer2_outputs(4026) <= not (a or b);
    layer2_outputs(4027) <= a and not b;
    layer2_outputs(4028) <= b;
    layer2_outputs(4029) <= not a or b;
    layer2_outputs(4030) <= not a or b;
    layer2_outputs(4031) <= not a;
    layer2_outputs(4032) <= b;
    layer2_outputs(4033) <= a;
    layer2_outputs(4034) <= not a;
    layer2_outputs(4035) <= not b;
    layer2_outputs(4036) <= a or b;
    layer2_outputs(4037) <= a or b;
    layer2_outputs(4038) <= '1';
    layer2_outputs(4039) <= not b or a;
    layer2_outputs(4040) <= b and not a;
    layer2_outputs(4041) <= not a;
    layer2_outputs(4042) <= '0';
    layer2_outputs(4043) <= '0';
    layer2_outputs(4044) <= a xor b;
    layer2_outputs(4045) <= a;
    layer2_outputs(4046) <= b and not a;
    layer2_outputs(4047) <= a and b;
    layer2_outputs(4048) <= not a or b;
    layer2_outputs(4049) <= not a or b;
    layer2_outputs(4050) <= b;
    layer2_outputs(4051) <= a;
    layer2_outputs(4052) <= '1';
    layer2_outputs(4053) <= a or b;
    layer2_outputs(4054) <= not a;
    layer2_outputs(4055) <= a;
    layer2_outputs(4056) <= not a;
    layer2_outputs(4057) <= not a;
    layer2_outputs(4058) <= a and b;
    layer2_outputs(4059) <= not (a and b);
    layer2_outputs(4060) <= a and b;
    layer2_outputs(4061) <= b;
    layer2_outputs(4062) <= not b;
    layer2_outputs(4063) <= a xor b;
    layer2_outputs(4064) <= '1';
    layer2_outputs(4065) <= not (a xor b);
    layer2_outputs(4066) <= not b;
    layer2_outputs(4067) <= a and not b;
    layer2_outputs(4068) <= a xor b;
    layer2_outputs(4069) <= a or b;
    layer2_outputs(4070) <= not (a and b);
    layer2_outputs(4071) <= a;
    layer2_outputs(4072) <= a;
    layer2_outputs(4073) <= b and not a;
    layer2_outputs(4074) <= not (a or b);
    layer2_outputs(4075) <= b and not a;
    layer2_outputs(4076) <= '1';
    layer2_outputs(4077) <= a or b;
    layer2_outputs(4078) <= not (a and b);
    layer2_outputs(4079) <= not (a xor b);
    layer2_outputs(4080) <= not b or a;
    layer2_outputs(4081) <= '1';
    layer2_outputs(4082) <= not b;
    layer2_outputs(4083) <= not a;
    layer2_outputs(4084) <= not (a or b);
    layer2_outputs(4085) <= not a or b;
    layer2_outputs(4086) <= not a;
    layer2_outputs(4087) <= a xor b;
    layer2_outputs(4088) <= not b;
    layer2_outputs(4089) <= not a;
    layer2_outputs(4090) <= not a or b;
    layer2_outputs(4091) <= '0';
    layer2_outputs(4092) <= not (a xor b);
    layer2_outputs(4093) <= not b or a;
    layer2_outputs(4094) <= not b or a;
    layer2_outputs(4095) <= not b or a;
    layer2_outputs(4096) <= not b or a;
    layer2_outputs(4097) <= a and b;
    layer2_outputs(4098) <= b;
    layer2_outputs(4099) <= b;
    layer2_outputs(4100) <= a or b;
    layer2_outputs(4101) <= a;
    layer2_outputs(4102) <= b and not a;
    layer2_outputs(4103) <= not (a or b);
    layer2_outputs(4104) <= not (a or b);
    layer2_outputs(4105) <= a and b;
    layer2_outputs(4106) <= not b;
    layer2_outputs(4107) <= not (a or b);
    layer2_outputs(4108) <= b and not a;
    layer2_outputs(4109) <= '0';
    layer2_outputs(4110) <= not b or a;
    layer2_outputs(4111) <= not b;
    layer2_outputs(4112) <= not a;
    layer2_outputs(4113) <= not a;
    layer2_outputs(4114) <= a and b;
    layer2_outputs(4115) <= a xor b;
    layer2_outputs(4116) <= not (a and b);
    layer2_outputs(4117) <= b;
    layer2_outputs(4118) <= not b;
    layer2_outputs(4119) <= '0';
    layer2_outputs(4120) <= not (a xor b);
    layer2_outputs(4121) <= not b or a;
    layer2_outputs(4122) <= b;
    layer2_outputs(4123) <= b;
    layer2_outputs(4124) <= a and b;
    layer2_outputs(4125) <= a and not b;
    layer2_outputs(4126) <= b;
    layer2_outputs(4127) <= a;
    layer2_outputs(4128) <= not b;
    layer2_outputs(4129) <= a;
    layer2_outputs(4130) <= a and not b;
    layer2_outputs(4131) <= not a;
    layer2_outputs(4132) <= b;
    layer2_outputs(4133) <= a and not b;
    layer2_outputs(4134) <= not (a and b);
    layer2_outputs(4135) <= b;
    layer2_outputs(4136) <= a;
    layer2_outputs(4137) <= not (a or b);
    layer2_outputs(4138) <= b and not a;
    layer2_outputs(4139) <= a and b;
    layer2_outputs(4140) <= '1';
    layer2_outputs(4141) <= b;
    layer2_outputs(4142) <= not (a and b);
    layer2_outputs(4143) <= not a or b;
    layer2_outputs(4144) <= a and b;
    layer2_outputs(4145) <= not b or a;
    layer2_outputs(4146) <= not (a and b);
    layer2_outputs(4147) <= not a;
    layer2_outputs(4148) <= a and not b;
    layer2_outputs(4149) <= not a;
    layer2_outputs(4150) <= not (a xor b);
    layer2_outputs(4151) <= b and not a;
    layer2_outputs(4152) <= not (a and b);
    layer2_outputs(4153) <= not (a or b);
    layer2_outputs(4154) <= not a;
    layer2_outputs(4155) <= not a;
    layer2_outputs(4156) <= '0';
    layer2_outputs(4157) <= '1';
    layer2_outputs(4158) <= not (a and b);
    layer2_outputs(4159) <= a or b;
    layer2_outputs(4160) <= not (a and b);
    layer2_outputs(4161) <= not (a and b);
    layer2_outputs(4162) <= b and not a;
    layer2_outputs(4163) <= b;
    layer2_outputs(4164) <= not b or a;
    layer2_outputs(4165) <= a and not b;
    layer2_outputs(4166) <= not (a and b);
    layer2_outputs(4167) <= a and not b;
    layer2_outputs(4168) <= '1';
    layer2_outputs(4169) <= not (a or b);
    layer2_outputs(4170) <= not a or b;
    layer2_outputs(4171) <= not (a and b);
    layer2_outputs(4172) <= '0';
    layer2_outputs(4173) <= not (a and b);
    layer2_outputs(4174) <= not (a and b);
    layer2_outputs(4175) <= a and b;
    layer2_outputs(4176) <= b and not a;
    layer2_outputs(4177) <= b and not a;
    layer2_outputs(4178) <= a or b;
    layer2_outputs(4179) <= not a or b;
    layer2_outputs(4180) <= '1';
    layer2_outputs(4181) <= not b;
    layer2_outputs(4182) <= not b;
    layer2_outputs(4183) <= not b;
    layer2_outputs(4184) <= not a;
    layer2_outputs(4185) <= not b or a;
    layer2_outputs(4186) <= b;
    layer2_outputs(4187) <= '1';
    layer2_outputs(4188) <= b;
    layer2_outputs(4189) <= '1';
    layer2_outputs(4190) <= not (a or b);
    layer2_outputs(4191) <= a or b;
    layer2_outputs(4192) <= not b or a;
    layer2_outputs(4193) <= not b or a;
    layer2_outputs(4194) <= a or b;
    layer2_outputs(4195) <= '1';
    layer2_outputs(4196) <= a xor b;
    layer2_outputs(4197) <= not a;
    layer2_outputs(4198) <= not (a xor b);
    layer2_outputs(4199) <= a and b;
    layer2_outputs(4200) <= not b or a;
    layer2_outputs(4201) <= a;
    layer2_outputs(4202) <= not (a and b);
    layer2_outputs(4203) <= b;
    layer2_outputs(4204) <= not a;
    layer2_outputs(4205) <= not a;
    layer2_outputs(4206) <= a;
    layer2_outputs(4207) <= a;
    layer2_outputs(4208) <= '0';
    layer2_outputs(4209) <= not b or a;
    layer2_outputs(4210) <= a;
    layer2_outputs(4211) <= a and b;
    layer2_outputs(4212) <= not a;
    layer2_outputs(4213) <= not (a or b);
    layer2_outputs(4214) <= not (a and b);
    layer2_outputs(4215) <= not (a xor b);
    layer2_outputs(4216) <= not (a xor b);
    layer2_outputs(4217) <= '0';
    layer2_outputs(4218) <= a and b;
    layer2_outputs(4219) <= not (a or b);
    layer2_outputs(4220) <= a or b;
    layer2_outputs(4221) <= not b;
    layer2_outputs(4222) <= not a or b;
    layer2_outputs(4223) <= b and not a;
    layer2_outputs(4224) <= a and b;
    layer2_outputs(4225) <= a or b;
    layer2_outputs(4226) <= a and not b;
    layer2_outputs(4227) <= a;
    layer2_outputs(4228) <= not b;
    layer2_outputs(4229) <= b;
    layer2_outputs(4230) <= not b or a;
    layer2_outputs(4231) <= not a or b;
    layer2_outputs(4232) <= not a or b;
    layer2_outputs(4233) <= a and not b;
    layer2_outputs(4234) <= not b or a;
    layer2_outputs(4235) <= a;
    layer2_outputs(4236) <= a;
    layer2_outputs(4237) <= a and not b;
    layer2_outputs(4238) <= not b;
    layer2_outputs(4239) <= not b;
    layer2_outputs(4240) <= not a or b;
    layer2_outputs(4241) <= a or b;
    layer2_outputs(4242) <= not a or b;
    layer2_outputs(4243) <= b and not a;
    layer2_outputs(4244) <= not (a or b);
    layer2_outputs(4245) <= a;
    layer2_outputs(4246) <= a;
    layer2_outputs(4247) <= a and not b;
    layer2_outputs(4248) <= not a or b;
    layer2_outputs(4249) <= b;
    layer2_outputs(4250) <= a and b;
    layer2_outputs(4251) <= not b;
    layer2_outputs(4252) <= not a;
    layer2_outputs(4253) <= a and not b;
    layer2_outputs(4254) <= not a;
    layer2_outputs(4255) <= b;
    layer2_outputs(4256) <= a or b;
    layer2_outputs(4257) <= not b or a;
    layer2_outputs(4258) <= not b;
    layer2_outputs(4259) <= not a;
    layer2_outputs(4260) <= '1';
    layer2_outputs(4261) <= not (a and b);
    layer2_outputs(4262) <= not b;
    layer2_outputs(4263) <= not b;
    layer2_outputs(4264) <= not a or b;
    layer2_outputs(4265) <= a or b;
    layer2_outputs(4266) <= a or b;
    layer2_outputs(4267) <= a xor b;
    layer2_outputs(4268) <= not (a and b);
    layer2_outputs(4269) <= not b;
    layer2_outputs(4270) <= a and not b;
    layer2_outputs(4271) <= a and not b;
    layer2_outputs(4272) <= not (a and b);
    layer2_outputs(4273) <= not a or b;
    layer2_outputs(4274) <= not (a or b);
    layer2_outputs(4275) <= a;
    layer2_outputs(4276) <= not (a or b);
    layer2_outputs(4277) <= '0';
    layer2_outputs(4278) <= a;
    layer2_outputs(4279) <= not b or a;
    layer2_outputs(4280) <= a and b;
    layer2_outputs(4281) <= a and b;
    layer2_outputs(4282) <= b and not a;
    layer2_outputs(4283) <= b;
    layer2_outputs(4284) <= not (a or b);
    layer2_outputs(4285) <= a and not b;
    layer2_outputs(4286) <= b and not a;
    layer2_outputs(4287) <= a or b;
    layer2_outputs(4288) <= a;
    layer2_outputs(4289) <= b and not a;
    layer2_outputs(4290) <= not b;
    layer2_outputs(4291) <= a;
    layer2_outputs(4292) <= b and not a;
    layer2_outputs(4293) <= not (a and b);
    layer2_outputs(4294) <= '0';
    layer2_outputs(4295) <= b and not a;
    layer2_outputs(4296) <= a and not b;
    layer2_outputs(4297) <= a and not b;
    layer2_outputs(4298) <= '1';
    layer2_outputs(4299) <= not (a and b);
    layer2_outputs(4300) <= a;
    layer2_outputs(4301) <= a and not b;
    layer2_outputs(4302) <= b;
    layer2_outputs(4303) <= a and not b;
    layer2_outputs(4304) <= '1';
    layer2_outputs(4305) <= not a or b;
    layer2_outputs(4306) <= '1';
    layer2_outputs(4307) <= b and not a;
    layer2_outputs(4308) <= not (a or b);
    layer2_outputs(4309) <= not b;
    layer2_outputs(4310) <= not b;
    layer2_outputs(4311) <= not b or a;
    layer2_outputs(4312) <= not (a or b);
    layer2_outputs(4313) <= a and not b;
    layer2_outputs(4314) <= not (a and b);
    layer2_outputs(4315) <= a and b;
    layer2_outputs(4316) <= not b or a;
    layer2_outputs(4317) <= a;
    layer2_outputs(4318) <= a;
    layer2_outputs(4319) <= not a;
    layer2_outputs(4320) <= a or b;
    layer2_outputs(4321) <= b;
    layer2_outputs(4322) <= not a or b;
    layer2_outputs(4323) <= a or b;
    layer2_outputs(4324) <= not (a and b);
    layer2_outputs(4325) <= b;
    layer2_outputs(4326) <= b and not a;
    layer2_outputs(4327) <= b;
    layer2_outputs(4328) <= not a;
    layer2_outputs(4329) <= not b or a;
    layer2_outputs(4330) <= a;
    layer2_outputs(4331) <= a and not b;
    layer2_outputs(4332) <= a or b;
    layer2_outputs(4333) <= not (a or b);
    layer2_outputs(4334) <= '0';
    layer2_outputs(4335) <= a;
    layer2_outputs(4336) <= not b;
    layer2_outputs(4337) <= not b or a;
    layer2_outputs(4338) <= not b or a;
    layer2_outputs(4339) <= not (a and b);
    layer2_outputs(4340) <= a or b;
    layer2_outputs(4341) <= a and not b;
    layer2_outputs(4342) <= a;
    layer2_outputs(4343) <= not b or a;
    layer2_outputs(4344) <= a or b;
    layer2_outputs(4345) <= b and not a;
    layer2_outputs(4346) <= '0';
    layer2_outputs(4347) <= not (a or b);
    layer2_outputs(4348) <= not (a and b);
    layer2_outputs(4349) <= a or b;
    layer2_outputs(4350) <= not (a xor b);
    layer2_outputs(4351) <= '1';
    layer2_outputs(4352) <= b and not a;
    layer2_outputs(4353) <= not (a or b);
    layer2_outputs(4354) <= not b or a;
    layer2_outputs(4355) <= not (a and b);
    layer2_outputs(4356) <= not (a and b);
    layer2_outputs(4357) <= '1';
    layer2_outputs(4358) <= not (a or b);
    layer2_outputs(4359) <= a and not b;
    layer2_outputs(4360) <= not b;
    layer2_outputs(4361) <= not a or b;
    layer2_outputs(4362) <= a and b;
    layer2_outputs(4363) <= a and not b;
    layer2_outputs(4364) <= not (a xor b);
    layer2_outputs(4365) <= a;
    layer2_outputs(4366) <= a or b;
    layer2_outputs(4367) <= not (a and b);
    layer2_outputs(4368) <= not b;
    layer2_outputs(4369) <= a;
    layer2_outputs(4370) <= a or b;
    layer2_outputs(4371) <= b;
    layer2_outputs(4372) <= not (a or b);
    layer2_outputs(4373) <= b;
    layer2_outputs(4374) <= not (a and b);
    layer2_outputs(4375) <= not b;
    layer2_outputs(4376) <= not (a or b);
    layer2_outputs(4377) <= b;
    layer2_outputs(4378) <= a or b;
    layer2_outputs(4379) <= not b;
    layer2_outputs(4380) <= '0';
    layer2_outputs(4381) <= b;
    layer2_outputs(4382) <= b and not a;
    layer2_outputs(4383) <= '1';
    layer2_outputs(4384) <= not b or a;
    layer2_outputs(4385) <= '1';
    layer2_outputs(4386) <= a and not b;
    layer2_outputs(4387) <= '1';
    layer2_outputs(4388) <= b and not a;
    layer2_outputs(4389) <= b and not a;
    layer2_outputs(4390) <= a and not b;
    layer2_outputs(4391) <= b;
    layer2_outputs(4392) <= '0';
    layer2_outputs(4393) <= a and not b;
    layer2_outputs(4394) <= not a;
    layer2_outputs(4395) <= '1';
    layer2_outputs(4396) <= a;
    layer2_outputs(4397) <= b;
    layer2_outputs(4398) <= b;
    layer2_outputs(4399) <= a and not b;
    layer2_outputs(4400) <= b;
    layer2_outputs(4401) <= a or b;
    layer2_outputs(4402) <= not (a xor b);
    layer2_outputs(4403) <= a and not b;
    layer2_outputs(4404) <= a and b;
    layer2_outputs(4405) <= b;
    layer2_outputs(4406) <= not (a and b);
    layer2_outputs(4407) <= not b;
    layer2_outputs(4408) <= a xor b;
    layer2_outputs(4409) <= b;
    layer2_outputs(4410) <= '0';
    layer2_outputs(4411) <= b;
    layer2_outputs(4412) <= not a;
    layer2_outputs(4413) <= not a;
    layer2_outputs(4414) <= '0';
    layer2_outputs(4415) <= not (a or b);
    layer2_outputs(4416) <= '1';
    layer2_outputs(4417) <= '1';
    layer2_outputs(4418) <= not (a or b);
    layer2_outputs(4419) <= b;
    layer2_outputs(4420) <= not a;
    layer2_outputs(4421) <= not b;
    layer2_outputs(4422) <= a xor b;
    layer2_outputs(4423) <= not b or a;
    layer2_outputs(4424) <= b;
    layer2_outputs(4425) <= a and not b;
    layer2_outputs(4426) <= not (a and b);
    layer2_outputs(4427) <= not b;
    layer2_outputs(4428) <= not (a and b);
    layer2_outputs(4429) <= not b or a;
    layer2_outputs(4430) <= not a;
    layer2_outputs(4431) <= not b;
    layer2_outputs(4432) <= a and not b;
    layer2_outputs(4433) <= a;
    layer2_outputs(4434) <= not b or a;
    layer2_outputs(4435) <= b and not a;
    layer2_outputs(4436) <= a xor b;
    layer2_outputs(4437) <= a xor b;
    layer2_outputs(4438) <= not b or a;
    layer2_outputs(4439) <= not (a and b);
    layer2_outputs(4440) <= not a;
    layer2_outputs(4441) <= not (a or b);
    layer2_outputs(4442) <= not (a xor b);
    layer2_outputs(4443) <= not b;
    layer2_outputs(4444) <= b and not a;
    layer2_outputs(4445) <= not (a or b);
    layer2_outputs(4446) <= b and not a;
    layer2_outputs(4447) <= not b;
    layer2_outputs(4448) <= '1';
    layer2_outputs(4449) <= a and b;
    layer2_outputs(4450) <= b;
    layer2_outputs(4451) <= a;
    layer2_outputs(4452) <= not (a xor b);
    layer2_outputs(4453) <= not a;
    layer2_outputs(4454) <= not b or a;
    layer2_outputs(4455) <= not (a or b);
    layer2_outputs(4456) <= a;
    layer2_outputs(4457) <= b;
    layer2_outputs(4458) <= a and b;
    layer2_outputs(4459) <= b;
    layer2_outputs(4460) <= not a or b;
    layer2_outputs(4461) <= not b;
    layer2_outputs(4462) <= '1';
    layer2_outputs(4463) <= a xor b;
    layer2_outputs(4464) <= b;
    layer2_outputs(4465) <= a and b;
    layer2_outputs(4466) <= not (a xor b);
    layer2_outputs(4467) <= not a;
    layer2_outputs(4468) <= not a or b;
    layer2_outputs(4469) <= '0';
    layer2_outputs(4470) <= '1';
    layer2_outputs(4471) <= b;
    layer2_outputs(4472) <= not a or b;
    layer2_outputs(4473) <= a or b;
    layer2_outputs(4474) <= b and not a;
    layer2_outputs(4475) <= a;
    layer2_outputs(4476) <= not a;
    layer2_outputs(4477) <= not a;
    layer2_outputs(4478) <= not b or a;
    layer2_outputs(4479) <= not a or b;
    layer2_outputs(4480) <= not (a or b);
    layer2_outputs(4481) <= a and not b;
    layer2_outputs(4482) <= not a;
    layer2_outputs(4483) <= not (a xor b);
    layer2_outputs(4484) <= a xor b;
    layer2_outputs(4485) <= a and b;
    layer2_outputs(4486) <= not a;
    layer2_outputs(4487) <= not a or b;
    layer2_outputs(4488) <= not a;
    layer2_outputs(4489) <= a;
    layer2_outputs(4490) <= not a;
    layer2_outputs(4491) <= not a;
    layer2_outputs(4492) <= not b;
    layer2_outputs(4493) <= '1';
    layer2_outputs(4494) <= b;
    layer2_outputs(4495) <= not a;
    layer2_outputs(4496) <= b;
    layer2_outputs(4497) <= a;
    layer2_outputs(4498) <= not (a and b);
    layer2_outputs(4499) <= a or b;
    layer2_outputs(4500) <= not b or a;
    layer2_outputs(4501) <= not (a or b);
    layer2_outputs(4502) <= b;
    layer2_outputs(4503) <= a;
    layer2_outputs(4504) <= a and b;
    layer2_outputs(4505) <= '1';
    layer2_outputs(4506) <= not a or b;
    layer2_outputs(4507) <= b and not a;
    layer2_outputs(4508) <= not a;
    layer2_outputs(4509) <= b;
    layer2_outputs(4510) <= not (a and b);
    layer2_outputs(4511) <= a and not b;
    layer2_outputs(4512) <= not b or a;
    layer2_outputs(4513) <= a and b;
    layer2_outputs(4514) <= not a or b;
    layer2_outputs(4515) <= a or b;
    layer2_outputs(4516) <= a;
    layer2_outputs(4517) <= a xor b;
    layer2_outputs(4518) <= not (a and b);
    layer2_outputs(4519) <= b;
    layer2_outputs(4520) <= not a;
    layer2_outputs(4521) <= not b or a;
    layer2_outputs(4522) <= a and b;
    layer2_outputs(4523) <= not b or a;
    layer2_outputs(4524) <= a or b;
    layer2_outputs(4525) <= b and not a;
    layer2_outputs(4526) <= b;
    layer2_outputs(4527) <= b;
    layer2_outputs(4528) <= b;
    layer2_outputs(4529) <= not (a and b);
    layer2_outputs(4530) <= a xor b;
    layer2_outputs(4531) <= a;
    layer2_outputs(4532) <= not b;
    layer2_outputs(4533) <= b;
    layer2_outputs(4534) <= not (a xor b);
    layer2_outputs(4535) <= not (a or b);
    layer2_outputs(4536) <= a;
    layer2_outputs(4537) <= not a;
    layer2_outputs(4538) <= not b or a;
    layer2_outputs(4539) <= not b;
    layer2_outputs(4540) <= not a or b;
    layer2_outputs(4541) <= not b;
    layer2_outputs(4542) <= not b or a;
    layer2_outputs(4543) <= b and not a;
    layer2_outputs(4544) <= b;
    layer2_outputs(4545) <= a or b;
    layer2_outputs(4546) <= a or b;
    layer2_outputs(4547) <= not b;
    layer2_outputs(4548) <= '0';
    layer2_outputs(4549) <= b and not a;
    layer2_outputs(4550) <= not b;
    layer2_outputs(4551) <= a;
    layer2_outputs(4552) <= not b;
    layer2_outputs(4553) <= '1';
    layer2_outputs(4554) <= a or b;
    layer2_outputs(4555) <= not a;
    layer2_outputs(4556) <= not a or b;
    layer2_outputs(4557) <= not a;
    layer2_outputs(4558) <= not a;
    layer2_outputs(4559) <= not (a and b);
    layer2_outputs(4560) <= b;
    layer2_outputs(4561) <= a;
    layer2_outputs(4562) <= not a;
    layer2_outputs(4563) <= not b;
    layer2_outputs(4564) <= a or b;
    layer2_outputs(4565) <= a;
    layer2_outputs(4566) <= b;
    layer2_outputs(4567) <= '0';
    layer2_outputs(4568) <= not (a xor b);
    layer2_outputs(4569) <= b;
    layer2_outputs(4570) <= a;
    layer2_outputs(4571) <= not a;
    layer2_outputs(4572) <= a and b;
    layer2_outputs(4573) <= a and not b;
    layer2_outputs(4574) <= a;
    layer2_outputs(4575) <= '1';
    layer2_outputs(4576) <= not a;
    layer2_outputs(4577) <= a;
    layer2_outputs(4578) <= not (a or b);
    layer2_outputs(4579) <= a;
    layer2_outputs(4580) <= not b or a;
    layer2_outputs(4581) <= not b or a;
    layer2_outputs(4582) <= a;
    layer2_outputs(4583) <= not a or b;
    layer2_outputs(4584) <= not b;
    layer2_outputs(4585) <= not (a xor b);
    layer2_outputs(4586) <= a xor b;
    layer2_outputs(4587) <= a;
    layer2_outputs(4588) <= not (a or b);
    layer2_outputs(4589) <= '0';
    layer2_outputs(4590) <= a;
    layer2_outputs(4591) <= '0';
    layer2_outputs(4592) <= not a;
    layer2_outputs(4593) <= a;
    layer2_outputs(4594) <= not (a or b);
    layer2_outputs(4595) <= a or b;
    layer2_outputs(4596) <= not a;
    layer2_outputs(4597) <= not (a or b);
    layer2_outputs(4598) <= a and not b;
    layer2_outputs(4599) <= not b;
    layer2_outputs(4600) <= a;
    layer2_outputs(4601) <= a and not b;
    layer2_outputs(4602) <= '0';
    layer2_outputs(4603) <= not a;
    layer2_outputs(4604) <= a and b;
    layer2_outputs(4605) <= not a or b;
    layer2_outputs(4606) <= not (a or b);
    layer2_outputs(4607) <= a and not b;
    layer2_outputs(4608) <= not b or a;
    layer2_outputs(4609) <= b;
    layer2_outputs(4610) <= '0';
    layer2_outputs(4611) <= b;
    layer2_outputs(4612) <= a and b;
    layer2_outputs(4613) <= not (a and b);
    layer2_outputs(4614) <= b and not a;
    layer2_outputs(4615) <= not b;
    layer2_outputs(4616) <= not b or a;
    layer2_outputs(4617) <= a;
    layer2_outputs(4618) <= b;
    layer2_outputs(4619) <= not a;
    layer2_outputs(4620) <= a and b;
    layer2_outputs(4621) <= a and not b;
    layer2_outputs(4622) <= not (a or b);
    layer2_outputs(4623) <= not a;
    layer2_outputs(4624) <= not (a or b);
    layer2_outputs(4625) <= a;
    layer2_outputs(4626) <= b;
    layer2_outputs(4627) <= not a;
    layer2_outputs(4628) <= not b or a;
    layer2_outputs(4629) <= not b;
    layer2_outputs(4630) <= a and not b;
    layer2_outputs(4631) <= a;
    layer2_outputs(4632) <= '0';
    layer2_outputs(4633) <= not b or a;
    layer2_outputs(4634) <= b;
    layer2_outputs(4635) <= a and not b;
    layer2_outputs(4636) <= not a or b;
    layer2_outputs(4637) <= not (a xor b);
    layer2_outputs(4638) <= a;
    layer2_outputs(4639) <= not a;
    layer2_outputs(4640) <= a;
    layer2_outputs(4641) <= not (a and b);
    layer2_outputs(4642) <= a;
    layer2_outputs(4643) <= not a;
    layer2_outputs(4644) <= not (a or b);
    layer2_outputs(4645) <= b and not a;
    layer2_outputs(4646) <= not a;
    layer2_outputs(4647) <= a and not b;
    layer2_outputs(4648) <= not b;
    layer2_outputs(4649) <= a xor b;
    layer2_outputs(4650) <= not b or a;
    layer2_outputs(4651) <= a or b;
    layer2_outputs(4652) <= b and not a;
    layer2_outputs(4653) <= a;
    layer2_outputs(4654) <= a or b;
    layer2_outputs(4655) <= not (a or b);
    layer2_outputs(4656) <= a or b;
    layer2_outputs(4657) <= a and b;
    layer2_outputs(4658) <= '1';
    layer2_outputs(4659) <= not a;
    layer2_outputs(4660) <= not a or b;
    layer2_outputs(4661) <= a and not b;
    layer2_outputs(4662) <= not a or b;
    layer2_outputs(4663) <= not a or b;
    layer2_outputs(4664) <= not a;
    layer2_outputs(4665) <= not b or a;
    layer2_outputs(4666) <= not b;
    layer2_outputs(4667) <= b and not a;
    layer2_outputs(4668) <= a;
    layer2_outputs(4669) <= not a;
    layer2_outputs(4670) <= a;
    layer2_outputs(4671) <= not a;
    layer2_outputs(4672) <= not a or b;
    layer2_outputs(4673) <= a and not b;
    layer2_outputs(4674) <= b and not a;
    layer2_outputs(4675) <= b;
    layer2_outputs(4676) <= not b or a;
    layer2_outputs(4677) <= not b or a;
    layer2_outputs(4678) <= '1';
    layer2_outputs(4679) <= not b;
    layer2_outputs(4680) <= a or b;
    layer2_outputs(4681) <= not (a or b);
    layer2_outputs(4682) <= not (a and b);
    layer2_outputs(4683) <= not (a and b);
    layer2_outputs(4684) <= not a;
    layer2_outputs(4685) <= a and b;
    layer2_outputs(4686) <= a and not b;
    layer2_outputs(4687) <= a and b;
    layer2_outputs(4688) <= not b or a;
    layer2_outputs(4689) <= not (a or b);
    layer2_outputs(4690) <= a and b;
    layer2_outputs(4691) <= not b or a;
    layer2_outputs(4692) <= not (a xor b);
    layer2_outputs(4693) <= b;
    layer2_outputs(4694) <= a;
    layer2_outputs(4695) <= a and b;
    layer2_outputs(4696) <= b;
    layer2_outputs(4697) <= '0';
    layer2_outputs(4698) <= a xor b;
    layer2_outputs(4699) <= not (a or b);
    layer2_outputs(4700) <= a or b;
    layer2_outputs(4701) <= b;
    layer2_outputs(4702) <= b;
    layer2_outputs(4703) <= a;
    layer2_outputs(4704) <= not b or a;
    layer2_outputs(4705) <= not b or a;
    layer2_outputs(4706) <= a and not b;
    layer2_outputs(4707) <= not (a or b);
    layer2_outputs(4708) <= not b or a;
    layer2_outputs(4709) <= not a;
    layer2_outputs(4710) <= a or b;
    layer2_outputs(4711) <= not b;
    layer2_outputs(4712) <= not (a xor b);
    layer2_outputs(4713) <= not (a or b);
    layer2_outputs(4714) <= not a or b;
    layer2_outputs(4715) <= b and not a;
    layer2_outputs(4716) <= not (a or b);
    layer2_outputs(4717) <= a and not b;
    layer2_outputs(4718) <= not (a xor b);
    layer2_outputs(4719) <= b and not a;
    layer2_outputs(4720) <= a or b;
    layer2_outputs(4721) <= '0';
    layer2_outputs(4722) <= b;
    layer2_outputs(4723) <= a;
    layer2_outputs(4724) <= a or b;
    layer2_outputs(4725) <= a;
    layer2_outputs(4726) <= not a;
    layer2_outputs(4727) <= a or b;
    layer2_outputs(4728) <= not b;
    layer2_outputs(4729) <= a or b;
    layer2_outputs(4730) <= not a;
    layer2_outputs(4731) <= b;
    layer2_outputs(4732) <= not (a and b);
    layer2_outputs(4733) <= a;
    layer2_outputs(4734) <= a or b;
    layer2_outputs(4735) <= a;
    layer2_outputs(4736) <= b;
    layer2_outputs(4737) <= a;
    layer2_outputs(4738) <= not b;
    layer2_outputs(4739) <= '0';
    layer2_outputs(4740) <= a;
    layer2_outputs(4741) <= not (a or b);
    layer2_outputs(4742) <= b and not a;
    layer2_outputs(4743) <= a;
    layer2_outputs(4744) <= not b;
    layer2_outputs(4745) <= not (a xor b);
    layer2_outputs(4746) <= not b;
    layer2_outputs(4747) <= not b;
    layer2_outputs(4748) <= not (a and b);
    layer2_outputs(4749) <= a;
    layer2_outputs(4750) <= not b or a;
    layer2_outputs(4751) <= a;
    layer2_outputs(4752) <= '0';
    layer2_outputs(4753) <= not a or b;
    layer2_outputs(4754) <= not a or b;
    layer2_outputs(4755) <= a and b;
    layer2_outputs(4756) <= not a or b;
    layer2_outputs(4757) <= not b or a;
    layer2_outputs(4758) <= a and not b;
    layer2_outputs(4759) <= not b;
    layer2_outputs(4760) <= a;
    layer2_outputs(4761) <= b and not a;
    layer2_outputs(4762) <= not a or b;
    layer2_outputs(4763) <= b;
    layer2_outputs(4764) <= a;
    layer2_outputs(4765) <= a;
    layer2_outputs(4766) <= a and not b;
    layer2_outputs(4767) <= '1';
    layer2_outputs(4768) <= not b;
    layer2_outputs(4769) <= not (a or b);
    layer2_outputs(4770) <= not (a and b);
    layer2_outputs(4771) <= not (a and b);
    layer2_outputs(4772) <= not b or a;
    layer2_outputs(4773) <= not (a or b);
    layer2_outputs(4774) <= '1';
    layer2_outputs(4775) <= a and b;
    layer2_outputs(4776) <= '0';
    layer2_outputs(4777) <= not a;
    layer2_outputs(4778) <= a and b;
    layer2_outputs(4779) <= not b;
    layer2_outputs(4780) <= a and not b;
    layer2_outputs(4781) <= b;
    layer2_outputs(4782) <= b;
    layer2_outputs(4783) <= a xor b;
    layer2_outputs(4784) <= a and b;
    layer2_outputs(4785) <= a and b;
    layer2_outputs(4786) <= '1';
    layer2_outputs(4787) <= b;
    layer2_outputs(4788) <= a and not b;
    layer2_outputs(4789) <= a and not b;
    layer2_outputs(4790) <= not b;
    layer2_outputs(4791) <= a;
    layer2_outputs(4792) <= not a or b;
    layer2_outputs(4793) <= not b;
    layer2_outputs(4794) <= not (a or b);
    layer2_outputs(4795) <= not b;
    layer2_outputs(4796) <= b;
    layer2_outputs(4797) <= not (a or b);
    layer2_outputs(4798) <= a xor b;
    layer2_outputs(4799) <= a;
    layer2_outputs(4800) <= not a;
    layer2_outputs(4801) <= a;
    layer2_outputs(4802) <= a;
    layer2_outputs(4803) <= not (a xor b);
    layer2_outputs(4804) <= a;
    layer2_outputs(4805) <= '1';
    layer2_outputs(4806) <= a;
    layer2_outputs(4807) <= not a;
    layer2_outputs(4808) <= not (a and b);
    layer2_outputs(4809) <= '0';
    layer2_outputs(4810) <= not b or a;
    layer2_outputs(4811) <= not (a and b);
    layer2_outputs(4812) <= a or b;
    layer2_outputs(4813) <= a and not b;
    layer2_outputs(4814) <= not a;
    layer2_outputs(4815) <= '0';
    layer2_outputs(4816) <= not a;
    layer2_outputs(4817) <= not a or b;
    layer2_outputs(4818) <= b;
    layer2_outputs(4819) <= '0';
    layer2_outputs(4820) <= not (a xor b);
    layer2_outputs(4821) <= b;
    layer2_outputs(4822) <= '1';
    layer2_outputs(4823) <= '1';
    layer2_outputs(4824) <= a;
    layer2_outputs(4825) <= not a;
    layer2_outputs(4826) <= not a or b;
    layer2_outputs(4827) <= not a or b;
    layer2_outputs(4828) <= b;
    layer2_outputs(4829) <= not b;
    layer2_outputs(4830) <= not a or b;
    layer2_outputs(4831) <= not (a or b);
    layer2_outputs(4832) <= not a;
    layer2_outputs(4833) <= not (a or b);
    layer2_outputs(4834) <= not (a and b);
    layer2_outputs(4835) <= a;
    layer2_outputs(4836) <= a xor b;
    layer2_outputs(4837) <= a xor b;
    layer2_outputs(4838) <= not a;
    layer2_outputs(4839) <= '0';
    layer2_outputs(4840) <= a or b;
    layer2_outputs(4841) <= a or b;
    layer2_outputs(4842) <= not a;
    layer2_outputs(4843) <= not b or a;
    layer2_outputs(4844) <= '0';
    layer2_outputs(4845) <= a or b;
    layer2_outputs(4846) <= a;
    layer2_outputs(4847) <= b and not a;
    layer2_outputs(4848) <= a and b;
    layer2_outputs(4849) <= not a or b;
    layer2_outputs(4850) <= b and not a;
    layer2_outputs(4851) <= a or b;
    layer2_outputs(4852) <= a and b;
    layer2_outputs(4853) <= b;
    layer2_outputs(4854) <= not (a or b);
    layer2_outputs(4855) <= not a;
    layer2_outputs(4856) <= not b;
    layer2_outputs(4857) <= not (a or b);
    layer2_outputs(4858) <= not b;
    layer2_outputs(4859) <= '1';
    layer2_outputs(4860) <= not b or a;
    layer2_outputs(4861) <= not b;
    layer2_outputs(4862) <= a;
    layer2_outputs(4863) <= '1';
    layer2_outputs(4864) <= '0';
    layer2_outputs(4865) <= not b;
    layer2_outputs(4866) <= b;
    layer2_outputs(4867) <= a and not b;
    layer2_outputs(4868) <= a;
    layer2_outputs(4869) <= a or b;
    layer2_outputs(4870) <= '0';
    layer2_outputs(4871) <= a;
    layer2_outputs(4872) <= b;
    layer2_outputs(4873) <= not (a and b);
    layer2_outputs(4874) <= not a or b;
    layer2_outputs(4875) <= a;
    layer2_outputs(4876) <= not a or b;
    layer2_outputs(4877) <= a and not b;
    layer2_outputs(4878) <= a and b;
    layer2_outputs(4879) <= not (a or b);
    layer2_outputs(4880) <= '0';
    layer2_outputs(4881) <= a or b;
    layer2_outputs(4882) <= not (a or b);
    layer2_outputs(4883) <= b;
    layer2_outputs(4884) <= a or b;
    layer2_outputs(4885) <= not b;
    layer2_outputs(4886) <= '0';
    layer2_outputs(4887) <= not (a or b);
    layer2_outputs(4888) <= a and not b;
    layer2_outputs(4889) <= not (a and b);
    layer2_outputs(4890) <= a;
    layer2_outputs(4891) <= not (a and b);
    layer2_outputs(4892) <= a and not b;
    layer2_outputs(4893) <= not b or a;
    layer2_outputs(4894) <= not a or b;
    layer2_outputs(4895) <= not (a and b);
    layer2_outputs(4896) <= not b;
    layer2_outputs(4897) <= b;
    layer2_outputs(4898) <= not (a and b);
    layer2_outputs(4899) <= not b;
    layer2_outputs(4900) <= a or b;
    layer2_outputs(4901) <= not b;
    layer2_outputs(4902) <= a and not b;
    layer2_outputs(4903) <= a xor b;
    layer2_outputs(4904) <= not a;
    layer2_outputs(4905) <= not (a xor b);
    layer2_outputs(4906) <= b;
    layer2_outputs(4907) <= a or b;
    layer2_outputs(4908) <= not a;
    layer2_outputs(4909) <= a and not b;
    layer2_outputs(4910) <= a and not b;
    layer2_outputs(4911) <= '0';
    layer2_outputs(4912) <= b;
    layer2_outputs(4913) <= not (a or b);
    layer2_outputs(4914) <= a and b;
    layer2_outputs(4915) <= '0';
    layer2_outputs(4916) <= not (a and b);
    layer2_outputs(4917) <= '0';
    layer2_outputs(4918) <= b and not a;
    layer2_outputs(4919) <= not (a and b);
    layer2_outputs(4920) <= not b;
    layer2_outputs(4921) <= not a or b;
    layer2_outputs(4922) <= not (a or b);
    layer2_outputs(4923) <= not b;
    layer2_outputs(4924) <= not (a and b);
    layer2_outputs(4925) <= not b;
    layer2_outputs(4926) <= not a;
    layer2_outputs(4927) <= a xor b;
    layer2_outputs(4928) <= a and b;
    layer2_outputs(4929) <= not (a or b);
    layer2_outputs(4930) <= not b or a;
    layer2_outputs(4931) <= a or b;
    layer2_outputs(4932) <= a;
    layer2_outputs(4933) <= a or b;
    layer2_outputs(4934) <= a or b;
    layer2_outputs(4935) <= '0';
    layer2_outputs(4936) <= '0';
    layer2_outputs(4937) <= a or b;
    layer2_outputs(4938) <= a;
    layer2_outputs(4939) <= not (a and b);
    layer2_outputs(4940) <= not b or a;
    layer2_outputs(4941) <= not b or a;
    layer2_outputs(4942) <= b;
    layer2_outputs(4943) <= not a;
    layer2_outputs(4944) <= a and b;
    layer2_outputs(4945) <= b;
    layer2_outputs(4946) <= not a;
    layer2_outputs(4947) <= b and not a;
    layer2_outputs(4948) <= not (a or b);
    layer2_outputs(4949) <= not b or a;
    layer2_outputs(4950) <= a and b;
    layer2_outputs(4951) <= '0';
    layer2_outputs(4952) <= a and not b;
    layer2_outputs(4953) <= not (a or b);
    layer2_outputs(4954) <= not b or a;
    layer2_outputs(4955) <= not a;
    layer2_outputs(4956) <= b;
    layer2_outputs(4957) <= b and not a;
    layer2_outputs(4958) <= '0';
    layer2_outputs(4959) <= '0';
    layer2_outputs(4960) <= not b or a;
    layer2_outputs(4961) <= not (a and b);
    layer2_outputs(4962) <= b and not a;
    layer2_outputs(4963) <= not (a or b);
    layer2_outputs(4964) <= b;
    layer2_outputs(4965) <= not b or a;
    layer2_outputs(4966) <= not a or b;
    layer2_outputs(4967) <= b;
    layer2_outputs(4968) <= b;
    layer2_outputs(4969) <= '1';
    layer2_outputs(4970) <= not (a and b);
    layer2_outputs(4971) <= not (a or b);
    layer2_outputs(4972) <= a and not b;
    layer2_outputs(4973) <= not a;
    layer2_outputs(4974) <= a;
    layer2_outputs(4975) <= '1';
    layer2_outputs(4976) <= a and not b;
    layer2_outputs(4977) <= not b or a;
    layer2_outputs(4978) <= a and b;
    layer2_outputs(4979) <= b;
    layer2_outputs(4980) <= not a;
    layer2_outputs(4981) <= a and not b;
    layer2_outputs(4982) <= not (a or b);
    layer2_outputs(4983) <= a or b;
    layer2_outputs(4984) <= not b;
    layer2_outputs(4985) <= a;
    layer2_outputs(4986) <= not a or b;
    layer2_outputs(4987) <= not a;
    layer2_outputs(4988) <= not a;
    layer2_outputs(4989) <= b and not a;
    layer2_outputs(4990) <= not b;
    layer2_outputs(4991) <= '0';
    layer2_outputs(4992) <= a;
    layer2_outputs(4993) <= '0';
    layer2_outputs(4994) <= '0';
    layer2_outputs(4995) <= not b;
    layer2_outputs(4996) <= not (a xor b);
    layer2_outputs(4997) <= not (a xor b);
    layer2_outputs(4998) <= '1';
    layer2_outputs(4999) <= not a;
    layer2_outputs(5000) <= not b;
    layer2_outputs(5001) <= a and not b;
    layer2_outputs(5002) <= b and not a;
    layer2_outputs(5003) <= a or b;
    layer2_outputs(5004) <= b;
    layer2_outputs(5005) <= a;
    layer2_outputs(5006) <= a;
    layer2_outputs(5007) <= '1';
    layer2_outputs(5008) <= not (a xor b);
    layer2_outputs(5009) <= '1';
    layer2_outputs(5010) <= b;
    layer2_outputs(5011) <= a;
    layer2_outputs(5012) <= '1';
    layer2_outputs(5013) <= b and not a;
    layer2_outputs(5014) <= a;
    layer2_outputs(5015) <= not b or a;
    layer2_outputs(5016) <= not b or a;
    layer2_outputs(5017) <= b;
    layer2_outputs(5018) <= not (a or b);
    layer2_outputs(5019) <= a;
    layer2_outputs(5020) <= not (a or b);
    layer2_outputs(5021) <= not a or b;
    layer2_outputs(5022) <= not (a and b);
    layer2_outputs(5023) <= not (a and b);
    layer2_outputs(5024) <= '0';
    layer2_outputs(5025) <= a and b;
    layer2_outputs(5026) <= not b;
    layer2_outputs(5027) <= not a or b;
    layer2_outputs(5028) <= b;
    layer2_outputs(5029) <= a and b;
    layer2_outputs(5030) <= not a;
    layer2_outputs(5031) <= not a;
    layer2_outputs(5032) <= a xor b;
    layer2_outputs(5033) <= a and b;
    layer2_outputs(5034) <= not b;
    layer2_outputs(5035) <= a and b;
    layer2_outputs(5036) <= b;
    layer2_outputs(5037) <= a or b;
    layer2_outputs(5038) <= b;
    layer2_outputs(5039) <= not (a and b);
    layer2_outputs(5040) <= b and not a;
    layer2_outputs(5041) <= not (a or b);
    layer2_outputs(5042) <= a xor b;
    layer2_outputs(5043) <= a and b;
    layer2_outputs(5044) <= b;
    layer2_outputs(5045) <= '1';
    layer2_outputs(5046) <= not (a or b);
    layer2_outputs(5047) <= not (a and b);
    layer2_outputs(5048) <= not b;
    layer2_outputs(5049) <= '1';
    layer2_outputs(5050) <= b;
    layer2_outputs(5051) <= b;
    layer2_outputs(5052) <= a or b;
    layer2_outputs(5053) <= b and not a;
    layer2_outputs(5054) <= b and not a;
    layer2_outputs(5055) <= not (a or b);
    layer2_outputs(5056) <= b;
    layer2_outputs(5057) <= a xor b;
    layer2_outputs(5058) <= not a or b;
    layer2_outputs(5059) <= '1';
    layer2_outputs(5060) <= not a;
    layer2_outputs(5061) <= a xor b;
    layer2_outputs(5062) <= not b;
    layer2_outputs(5063) <= a;
    layer2_outputs(5064) <= a or b;
    layer2_outputs(5065) <= b and not a;
    layer2_outputs(5066) <= b and not a;
    layer2_outputs(5067) <= not a or b;
    layer2_outputs(5068) <= a;
    layer2_outputs(5069) <= a and not b;
    layer2_outputs(5070) <= a and b;
    layer2_outputs(5071) <= b;
    layer2_outputs(5072) <= a and b;
    layer2_outputs(5073) <= a or b;
    layer2_outputs(5074) <= b;
    layer2_outputs(5075) <= a and b;
    layer2_outputs(5076) <= not (a or b);
    layer2_outputs(5077) <= not a or b;
    layer2_outputs(5078) <= '1';
    layer2_outputs(5079) <= not b or a;
    layer2_outputs(5080) <= not a or b;
    layer2_outputs(5081) <= '1';
    layer2_outputs(5082) <= '1';
    layer2_outputs(5083) <= b;
    layer2_outputs(5084) <= not (a or b);
    layer2_outputs(5085) <= b and not a;
    layer2_outputs(5086) <= not (a xor b);
    layer2_outputs(5087) <= not b;
    layer2_outputs(5088) <= not (a or b);
    layer2_outputs(5089) <= a;
    layer2_outputs(5090) <= b and not a;
    layer2_outputs(5091) <= not b;
    layer2_outputs(5092) <= not a or b;
    layer2_outputs(5093) <= b;
    layer2_outputs(5094) <= a;
    layer2_outputs(5095) <= not (a or b);
    layer2_outputs(5096) <= '1';
    layer2_outputs(5097) <= '0';
    layer2_outputs(5098) <= a and not b;
    layer2_outputs(5099) <= not b;
    layer2_outputs(5100) <= not a;
    layer2_outputs(5101) <= not b;
    layer2_outputs(5102) <= a and b;
    layer2_outputs(5103) <= a or b;
    layer2_outputs(5104) <= not (a xor b);
    layer2_outputs(5105) <= a and not b;
    layer2_outputs(5106) <= not (a and b);
    layer2_outputs(5107) <= a or b;
    layer2_outputs(5108) <= not (a or b);
    layer2_outputs(5109) <= b;
    layer2_outputs(5110) <= a or b;
    layer2_outputs(5111) <= not (a and b);
    layer2_outputs(5112) <= not a;
    layer2_outputs(5113) <= a;
    layer2_outputs(5114) <= not b;
    layer2_outputs(5115) <= a and not b;
    layer2_outputs(5116) <= not b;
    layer2_outputs(5117) <= not a;
    layer2_outputs(5118) <= not a;
    layer2_outputs(5119) <= b;
    layer2_outputs(5120) <= not (a or b);
    layer2_outputs(5121) <= a;
    layer2_outputs(5122) <= not (a xor b);
    layer2_outputs(5123) <= b and not a;
    layer2_outputs(5124) <= b and not a;
    layer2_outputs(5125) <= not (a xor b);
    layer2_outputs(5126) <= not (a or b);
    layer2_outputs(5127) <= not a or b;
    layer2_outputs(5128) <= not b;
    layer2_outputs(5129) <= not b or a;
    layer2_outputs(5130) <= '0';
    layer2_outputs(5131) <= not a or b;
    layer2_outputs(5132) <= b;
    layer2_outputs(5133) <= a and b;
    layer2_outputs(5134) <= not (a and b);
    layer2_outputs(5135) <= not a or b;
    layer2_outputs(5136) <= not (a or b);
    layer2_outputs(5137) <= not b;
    layer2_outputs(5138) <= a;
    layer2_outputs(5139) <= a and not b;
    layer2_outputs(5140) <= b;
    layer2_outputs(5141) <= a and b;
    layer2_outputs(5142) <= not b or a;
    layer2_outputs(5143) <= a and b;
    layer2_outputs(5144) <= a and b;
    layer2_outputs(5145) <= a;
    layer2_outputs(5146) <= not (a or b);
    layer2_outputs(5147) <= not b or a;
    layer2_outputs(5148) <= b;
    layer2_outputs(5149) <= a and b;
    layer2_outputs(5150) <= '0';
    layer2_outputs(5151) <= '0';
    layer2_outputs(5152) <= not a;
    layer2_outputs(5153) <= b;
    layer2_outputs(5154) <= b and not a;
    layer2_outputs(5155) <= a;
    layer2_outputs(5156) <= not b or a;
    layer2_outputs(5157) <= b and not a;
    layer2_outputs(5158) <= a xor b;
    layer2_outputs(5159) <= a and not b;
    layer2_outputs(5160) <= b;
    layer2_outputs(5161) <= b;
    layer2_outputs(5162) <= b and not a;
    layer2_outputs(5163) <= '0';
    layer2_outputs(5164) <= not b or a;
    layer2_outputs(5165) <= b;
    layer2_outputs(5166) <= a and not b;
    layer2_outputs(5167) <= not b or a;
    layer2_outputs(5168) <= not a or b;
    layer2_outputs(5169) <= a and b;
    layer2_outputs(5170) <= not b;
    layer2_outputs(5171) <= b;
    layer2_outputs(5172) <= a;
    layer2_outputs(5173) <= b;
    layer2_outputs(5174) <= not a or b;
    layer2_outputs(5175) <= not a;
    layer2_outputs(5176) <= not a or b;
    layer2_outputs(5177) <= a and b;
    layer2_outputs(5178) <= a xor b;
    layer2_outputs(5179) <= a;
    layer2_outputs(5180) <= not a or b;
    layer2_outputs(5181) <= not a;
    layer2_outputs(5182) <= not b or a;
    layer2_outputs(5183) <= not b;
    layer2_outputs(5184) <= b;
    layer2_outputs(5185) <= not b or a;
    layer2_outputs(5186) <= b;
    layer2_outputs(5187) <= a or b;
    layer2_outputs(5188) <= a;
    layer2_outputs(5189) <= not (a and b);
    layer2_outputs(5190) <= not (a or b);
    layer2_outputs(5191) <= b;
    layer2_outputs(5192) <= b and not a;
    layer2_outputs(5193) <= not b;
    layer2_outputs(5194) <= b;
    layer2_outputs(5195) <= a and not b;
    layer2_outputs(5196) <= not b;
    layer2_outputs(5197) <= a and b;
    layer2_outputs(5198) <= not b or a;
    layer2_outputs(5199) <= a xor b;
    layer2_outputs(5200) <= not a or b;
    layer2_outputs(5201) <= b and not a;
    layer2_outputs(5202) <= not a;
    layer2_outputs(5203) <= a xor b;
    layer2_outputs(5204) <= a;
    layer2_outputs(5205) <= a;
    layer2_outputs(5206) <= not a or b;
    layer2_outputs(5207) <= not (a and b);
    layer2_outputs(5208) <= '0';
    layer2_outputs(5209) <= b;
    layer2_outputs(5210) <= not a;
    layer2_outputs(5211) <= b;
    layer2_outputs(5212) <= a;
    layer2_outputs(5213) <= b and not a;
    layer2_outputs(5214) <= not (a and b);
    layer2_outputs(5215) <= not (a or b);
    layer2_outputs(5216) <= a and not b;
    layer2_outputs(5217) <= not a;
    layer2_outputs(5218) <= '1';
    layer2_outputs(5219) <= a and b;
    layer2_outputs(5220) <= a;
    layer2_outputs(5221) <= a or b;
    layer2_outputs(5222) <= '0';
    layer2_outputs(5223) <= a xor b;
    layer2_outputs(5224) <= b and not a;
    layer2_outputs(5225) <= '1';
    layer2_outputs(5226) <= a and b;
    layer2_outputs(5227) <= a;
    layer2_outputs(5228) <= not (a xor b);
    layer2_outputs(5229) <= not b or a;
    layer2_outputs(5230) <= not a;
    layer2_outputs(5231) <= b and not a;
    layer2_outputs(5232) <= a and b;
    layer2_outputs(5233) <= not (a or b);
    layer2_outputs(5234) <= a xor b;
    layer2_outputs(5235) <= '1';
    layer2_outputs(5236) <= not a or b;
    layer2_outputs(5237) <= not a or b;
    layer2_outputs(5238) <= a;
    layer2_outputs(5239) <= not (a and b);
    layer2_outputs(5240) <= a xor b;
    layer2_outputs(5241) <= b;
    layer2_outputs(5242) <= a and b;
    layer2_outputs(5243) <= a and b;
    layer2_outputs(5244) <= not b or a;
    layer2_outputs(5245) <= '1';
    layer2_outputs(5246) <= '1';
    layer2_outputs(5247) <= not b or a;
    layer2_outputs(5248) <= not b;
    layer2_outputs(5249) <= a and not b;
    layer2_outputs(5250) <= not a;
    layer2_outputs(5251) <= a;
    layer2_outputs(5252) <= not a;
    layer2_outputs(5253) <= not (a and b);
    layer2_outputs(5254) <= a;
    layer2_outputs(5255) <= '1';
    layer2_outputs(5256) <= not (a and b);
    layer2_outputs(5257) <= a and b;
    layer2_outputs(5258) <= b;
    layer2_outputs(5259) <= not (a xor b);
    layer2_outputs(5260) <= '0';
    layer2_outputs(5261) <= not (a and b);
    layer2_outputs(5262) <= '0';
    layer2_outputs(5263) <= not b;
    layer2_outputs(5264) <= not (a and b);
    layer2_outputs(5265) <= not (a xor b);
    layer2_outputs(5266) <= not a;
    layer2_outputs(5267) <= not (a and b);
    layer2_outputs(5268) <= a;
    layer2_outputs(5269) <= '1';
    layer2_outputs(5270) <= not (a or b);
    layer2_outputs(5271) <= not a;
    layer2_outputs(5272) <= not b;
    layer2_outputs(5273) <= not a;
    layer2_outputs(5274) <= not (a or b);
    layer2_outputs(5275) <= a;
    layer2_outputs(5276) <= b and not a;
    layer2_outputs(5277) <= not a;
    layer2_outputs(5278) <= a;
    layer2_outputs(5279) <= '0';
    layer2_outputs(5280) <= not b or a;
    layer2_outputs(5281) <= a xor b;
    layer2_outputs(5282) <= not (a xor b);
    layer2_outputs(5283) <= not a;
    layer2_outputs(5284) <= b;
    layer2_outputs(5285) <= a or b;
    layer2_outputs(5286) <= not b;
    layer2_outputs(5287) <= not b or a;
    layer2_outputs(5288) <= not (a and b);
    layer2_outputs(5289) <= not a or b;
    layer2_outputs(5290) <= a;
    layer2_outputs(5291) <= a and b;
    layer2_outputs(5292) <= not b;
    layer2_outputs(5293) <= not (a and b);
    layer2_outputs(5294) <= not (a or b);
    layer2_outputs(5295) <= a;
    layer2_outputs(5296) <= not a or b;
    layer2_outputs(5297) <= a or b;
    layer2_outputs(5298) <= a xor b;
    layer2_outputs(5299) <= b;
    layer2_outputs(5300) <= a;
    layer2_outputs(5301) <= a;
    layer2_outputs(5302) <= b and not a;
    layer2_outputs(5303) <= a xor b;
    layer2_outputs(5304) <= not (a or b);
    layer2_outputs(5305) <= not a or b;
    layer2_outputs(5306) <= b;
    layer2_outputs(5307) <= not a;
    layer2_outputs(5308) <= not a or b;
    layer2_outputs(5309) <= not a;
    layer2_outputs(5310) <= a and b;
    layer2_outputs(5311) <= not (a and b);
    layer2_outputs(5312) <= not b;
    layer2_outputs(5313) <= a;
    layer2_outputs(5314) <= not b;
    layer2_outputs(5315) <= not a;
    layer2_outputs(5316) <= a and b;
    layer2_outputs(5317) <= a and not b;
    layer2_outputs(5318) <= not (a or b);
    layer2_outputs(5319) <= not (a and b);
    layer2_outputs(5320) <= a xor b;
    layer2_outputs(5321) <= '1';
    layer2_outputs(5322) <= b and not a;
    layer2_outputs(5323) <= b;
    layer2_outputs(5324) <= '1';
    layer2_outputs(5325) <= a or b;
    layer2_outputs(5326) <= a and b;
    layer2_outputs(5327) <= a and b;
    layer2_outputs(5328) <= not b or a;
    layer2_outputs(5329) <= a and b;
    layer2_outputs(5330) <= a xor b;
    layer2_outputs(5331) <= b and not a;
    layer2_outputs(5332) <= not a;
    layer2_outputs(5333) <= b;
    layer2_outputs(5334) <= not a;
    layer2_outputs(5335) <= not (a and b);
    layer2_outputs(5336) <= b and not a;
    layer2_outputs(5337) <= '0';
    layer2_outputs(5338) <= not a;
    layer2_outputs(5339) <= a or b;
    layer2_outputs(5340) <= not (a or b);
    layer2_outputs(5341) <= a xor b;
    layer2_outputs(5342) <= not (a and b);
    layer2_outputs(5343) <= a;
    layer2_outputs(5344) <= a and not b;
    layer2_outputs(5345) <= not a;
    layer2_outputs(5346) <= not a;
    layer2_outputs(5347) <= a xor b;
    layer2_outputs(5348) <= a and b;
    layer2_outputs(5349) <= '0';
    layer2_outputs(5350) <= a and not b;
    layer2_outputs(5351) <= not (a or b);
    layer2_outputs(5352) <= a;
    layer2_outputs(5353) <= a xor b;
    layer2_outputs(5354) <= a and not b;
    layer2_outputs(5355) <= not (a xor b);
    layer2_outputs(5356) <= a or b;
    layer2_outputs(5357) <= b and not a;
    layer2_outputs(5358) <= not a or b;
    layer2_outputs(5359) <= not a;
    layer2_outputs(5360) <= a xor b;
    layer2_outputs(5361) <= b and not a;
    layer2_outputs(5362) <= a and b;
    layer2_outputs(5363) <= not b;
    layer2_outputs(5364) <= a;
    layer2_outputs(5365) <= a and not b;
    layer2_outputs(5366) <= not (a and b);
    layer2_outputs(5367) <= not a;
    layer2_outputs(5368) <= a xor b;
    layer2_outputs(5369) <= not a or b;
    layer2_outputs(5370) <= a xor b;
    layer2_outputs(5371) <= a and b;
    layer2_outputs(5372) <= not (a or b);
    layer2_outputs(5373) <= b;
    layer2_outputs(5374) <= a;
    layer2_outputs(5375) <= not (a and b);
    layer2_outputs(5376) <= a or b;
    layer2_outputs(5377) <= not (a and b);
    layer2_outputs(5378) <= not a or b;
    layer2_outputs(5379) <= '0';
    layer2_outputs(5380) <= '1';
    layer2_outputs(5381) <= b and not a;
    layer2_outputs(5382) <= b;
    layer2_outputs(5383) <= not b or a;
    layer2_outputs(5384) <= not b;
    layer2_outputs(5385) <= not a;
    layer2_outputs(5386) <= not b;
    layer2_outputs(5387) <= not (a and b);
    layer2_outputs(5388) <= b;
    layer2_outputs(5389) <= a or b;
    layer2_outputs(5390) <= a;
    layer2_outputs(5391) <= not b;
    layer2_outputs(5392) <= a or b;
    layer2_outputs(5393) <= not (a xor b);
    layer2_outputs(5394) <= a and not b;
    layer2_outputs(5395) <= not (a and b);
    layer2_outputs(5396) <= a and not b;
    layer2_outputs(5397) <= not (a xor b);
    layer2_outputs(5398) <= not b;
    layer2_outputs(5399) <= a and not b;
    layer2_outputs(5400) <= a;
    layer2_outputs(5401) <= a and not b;
    layer2_outputs(5402) <= a;
    layer2_outputs(5403) <= a;
    layer2_outputs(5404) <= '0';
    layer2_outputs(5405) <= a;
    layer2_outputs(5406) <= b;
    layer2_outputs(5407) <= not (a xor b);
    layer2_outputs(5408) <= a and not b;
    layer2_outputs(5409) <= a;
    layer2_outputs(5410) <= a and not b;
    layer2_outputs(5411) <= b;
    layer2_outputs(5412) <= a;
    layer2_outputs(5413) <= not b or a;
    layer2_outputs(5414) <= not (a xor b);
    layer2_outputs(5415) <= '1';
    layer2_outputs(5416) <= a and not b;
    layer2_outputs(5417) <= not b;
    layer2_outputs(5418) <= not b;
    layer2_outputs(5419) <= a and not b;
    layer2_outputs(5420) <= a;
    layer2_outputs(5421) <= not b;
    layer2_outputs(5422) <= a or b;
    layer2_outputs(5423) <= a and not b;
    layer2_outputs(5424) <= not (a xor b);
    layer2_outputs(5425) <= not a;
    layer2_outputs(5426) <= not a;
    layer2_outputs(5427) <= a or b;
    layer2_outputs(5428) <= b;
    layer2_outputs(5429) <= a;
    layer2_outputs(5430) <= a;
    layer2_outputs(5431) <= not a;
    layer2_outputs(5432) <= b;
    layer2_outputs(5433) <= a;
    layer2_outputs(5434) <= a xor b;
    layer2_outputs(5435) <= a xor b;
    layer2_outputs(5436) <= not b;
    layer2_outputs(5437) <= '1';
    layer2_outputs(5438) <= a;
    layer2_outputs(5439) <= not (a or b);
    layer2_outputs(5440) <= '0';
    layer2_outputs(5441) <= not b or a;
    layer2_outputs(5442) <= not b or a;
    layer2_outputs(5443) <= b and not a;
    layer2_outputs(5444) <= not b;
    layer2_outputs(5445) <= b and not a;
    layer2_outputs(5446) <= not (a or b);
    layer2_outputs(5447) <= not a;
    layer2_outputs(5448) <= a and b;
    layer2_outputs(5449) <= not a;
    layer2_outputs(5450) <= not b;
    layer2_outputs(5451) <= b;
    layer2_outputs(5452) <= a and not b;
    layer2_outputs(5453) <= b;
    layer2_outputs(5454) <= a and b;
    layer2_outputs(5455) <= a and not b;
    layer2_outputs(5456) <= not a or b;
    layer2_outputs(5457) <= a or b;
    layer2_outputs(5458) <= not b;
    layer2_outputs(5459) <= a and not b;
    layer2_outputs(5460) <= not b or a;
    layer2_outputs(5461) <= not a;
    layer2_outputs(5462) <= b and not a;
    layer2_outputs(5463) <= '1';
    layer2_outputs(5464) <= not a or b;
    layer2_outputs(5465) <= a and b;
    layer2_outputs(5466) <= '1';
    layer2_outputs(5467) <= not a;
    layer2_outputs(5468) <= b and not a;
    layer2_outputs(5469) <= not (a xor b);
    layer2_outputs(5470) <= a and b;
    layer2_outputs(5471) <= not (a and b);
    layer2_outputs(5472) <= '0';
    layer2_outputs(5473) <= b;
    layer2_outputs(5474) <= b and not a;
    layer2_outputs(5475) <= b and not a;
    layer2_outputs(5476) <= not a;
    layer2_outputs(5477) <= not a;
    layer2_outputs(5478) <= not b or a;
    layer2_outputs(5479) <= a and not b;
    layer2_outputs(5480) <= a or b;
    layer2_outputs(5481) <= '0';
    layer2_outputs(5482) <= not a or b;
    layer2_outputs(5483) <= b and not a;
    layer2_outputs(5484) <= a or b;
    layer2_outputs(5485) <= not (a xor b);
    layer2_outputs(5486) <= a and b;
    layer2_outputs(5487) <= a;
    layer2_outputs(5488) <= b;
    layer2_outputs(5489) <= '0';
    layer2_outputs(5490) <= b;
    layer2_outputs(5491) <= b and not a;
    layer2_outputs(5492) <= a or b;
    layer2_outputs(5493) <= a or b;
    layer2_outputs(5494) <= a or b;
    layer2_outputs(5495) <= not b or a;
    layer2_outputs(5496) <= '1';
    layer2_outputs(5497) <= '1';
    layer2_outputs(5498) <= a and not b;
    layer2_outputs(5499) <= a;
    layer2_outputs(5500) <= a and b;
    layer2_outputs(5501) <= not (a and b);
    layer2_outputs(5502) <= not b or a;
    layer2_outputs(5503) <= b;
    layer2_outputs(5504) <= not (a or b);
    layer2_outputs(5505) <= a and b;
    layer2_outputs(5506) <= not b;
    layer2_outputs(5507) <= b;
    layer2_outputs(5508) <= not (a and b);
    layer2_outputs(5509) <= not b or a;
    layer2_outputs(5510) <= a;
    layer2_outputs(5511) <= '1';
    layer2_outputs(5512) <= not a;
    layer2_outputs(5513) <= not (a or b);
    layer2_outputs(5514) <= not (a or b);
    layer2_outputs(5515) <= a or b;
    layer2_outputs(5516) <= not b;
    layer2_outputs(5517) <= a;
    layer2_outputs(5518) <= a or b;
    layer2_outputs(5519) <= '0';
    layer2_outputs(5520) <= b and not a;
    layer2_outputs(5521) <= not a or b;
    layer2_outputs(5522) <= '0';
    layer2_outputs(5523) <= a and not b;
    layer2_outputs(5524) <= not a or b;
    layer2_outputs(5525) <= not (a or b);
    layer2_outputs(5526) <= not b or a;
    layer2_outputs(5527) <= a;
    layer2_outputs(5528) <= a and not b;
    layer2_outputs(5529) <= b;
    layer2_outputs(5530) <= a or b;
    layer2_outputs(5531) <= not (a or b);
    layer2_outputs(5532) <= a and not b;
    layer2_outputs(5533) <= a and b;
    layer2_outputs(5534) <= not (a xor b);
    layer2_outputs(5535) <= not (a xor b);
    layer2_outputs(5536) <= not b or a;
    layer2_outputs(5537) <= b;
    layer2_outputs(5538) <= not (a xor b);
    layer2_outputs(5539) <= not b;
    layer2_outputs(5540) <= a or b;
    layer2_outputs(5541) <= '1';
    layer2_outputs(5542) <= not (a and b);
    layer2_outputs(5543) <= a or b;
    layer2_outputs(5544) <= not b;
    layer2_outputs(5545) <= a xor b;
    layer2_outputs(5546) <= '0';
    layer2_outputs(5547) <= a or b;
    layer2_outputs(5548) <= not b or a;
    layer2_outputs(5549) <= not a;
    layer2_outputs(5550) <= not b or a;
    layer2_outputs(5551) <= b;
    layer2_outputs(5552) <= not b;
    layer2_outputs(5553) <= b and not a;
    layer2_outputs(5554) <= a and not b;
    layer2_outputs(5555) <= a and b;
    layer2_outputs(5556) <= a and b;
    layer2_outputs(5557) <= not (a xor b);
    layer2_outputs(5558) <= b;
    layer2_outputs(5559) <= a;
    layer2_outputs(5560) <= a and not b;
    layer2_outputs(5561) <= not b;
    layer2_outputs(5562) <= not (a and b);
    layer2_outputs(5563) <= not (a or b);
    layer2_outputs(5564) <= not (a or b);
    layer2_outputs(5565) <= a;
    layer2_outputs(5566) <= a xor b;
    layer2_outputs(5567) <= b and not a;
    layer2_outputs(5568) <= a or b;
    layer2_outputs(5569) <= a and not b;
    layer2_outputs(5570) <= not (a and b);
    layer2_outputs(5571) <= a;
    layer2_outputs(5572) <= not (a and b);
    layer2_outputs(5573) <= b and not a;
    layer2_outputs(5574) <= b;
    layer2_outputs(5575) <= a and not b;
    layer2_outputs(5576) <= a and not b;
    layer2_outputs(5577) <= not b;
    layer2_outputs(5578) <= a and b;
    layer2_outputs(5579) <= not (a xor b);
    layer2_outputs(5580) <= b;
    layer2_outputs(5581) <= a or b;
    layer2_outputs(5582) <= a xor b;
    layer2_outputs(5583) <= a xor b;
    layer2_outputs(5584) <= '1';
    layer2_outputs(5585) <= a;
    layer2_outputs(5586) <= a;
    layer2_outputs(5587) <= not a or b;
    layer2_outputs(5588) <= not b or a;
    layer2_outputs(5589) <= not a or b;
    layer2_outputs(5590) <= not a or b;
    layer2_outputs(5591) <= a;
    layer2_outputs(5592) <= not b or a;
    layer2_outputs(5593) <= not a;
    layer2_outputs(5594) <= not b or a;
    layer2_outputs(5595) <= a or b;
    layer2_outputs(5596) <= a and not b;
    layer2_outputs(5597) <= b;
    layer2_outputs(5598) <= not (a xor b);
    layer2_outputs(5599) <= not a or b;
    layer2_outputs(5600) <= b;
    layer2_outputs(5601) <= not a or b;
    layer2_outputs(5602) <= '0';
    layer2_outputs(5603) <= not (a and b);
    layer2_outputs(5604) <= a or b;
    layer2_outputs(5605) <= '0';
    layer2_outputs(5606) <= not a or b;
    layer2_outputs(5607) <= b;
    layer2_outputs(5608) <= not b;
    layer2_outputs(5609) <= '0';
    layer2_outputs(5610) <= not (a xor b);
    layer2_outputs(5611) <= not b or a;
    layer2_outputs(5612) <= a;
    layer2_outputs(5613) <= '0';
    layer2_outputs(5614) <= a or b;
    layer2_outputs(5615) <= '1';
    layer2_outputs(5616) <= not a or b;
    layer2_outputs(5617) <= b;
    layer2_outputs(5618) <= not b or a;
    layer2_outputs(5619) <= not b or a;
    layer2_outputs(5620) <= a and b;
    layer2_outputs(5621) <= a and b;
    layer2_outputs(5622) <= not b or a;
    layer2_outputs(5623) <= a;
    layer2_outputs(5624) <= b;
    layer2_outputs(5625) <= b;
    layer2_outputs(5626) <= a and not b;
    layer2_outputs(5627) <= b;
    layer2_outputs(5628) <= not b;
    layer2_outputs(5629) <= '1';
    layer2_outputs(5630) <= a xor b;
    layer2_outputs(5631) <= a and not b;
    layer2_outputs(5632) <= b;
    layer2_outputs(5633) <= b;
    layer2_outputs(5634) <= not a;
    layer2_outputs(5635) <= not a;
    layer2_outputs(5636) <= '1';
    layer2_outputs(5637) <= b and not a;
    layer2_outputs(5638) <= not b;
    layer2_outputs(5639) <= a and not b;
    layer2_outputs(5640) <= not a or b;
    layer2_outputs(5641) <= not a or b;
    layer2_outputs(5642) <= b and not a;
    layer2_outputs(5643) <= b;
    layer2_outputs(5644) <= a;
    layer2_outputs(5645) <= b and not a;
    layer2_outputs(5646) <= a;
    layer2_outputs(5647) <= a and b;
    layer2_outputs(5648) <= a and not b;
    layer2_outputs(5649) <= not b;
    layer2_outputs(5650) <= b and not a;
    layer2_outputs(5651) <= not b or a;
    layer2_outputs(5652) <= '1';
    layer2_outputs(5653) <= not a or b;
    layer2_outputs(5654) <= b;
    layer2_outputs(5655) <= a and not b;
    layer2_outputs(5656) <= not a;
    layer2_outputs(5657) <= a xor b;
    layer2_outputs(5658) <= not b or a;
    layer2_outputs(5659) <= not b or a;
    layer2_outputs(5660) <= b and not a;
    layer2_outputs(5661) <= not a;
    layer2_outputs(5662) <= a;
    layer2_outputs(5663) <= b and not a;
    layer2_outputs(5664) <= not (a and b);
    layer2_outputs(5665) <= b;
    layer2_outputs(5666) <= not b;
    layer2_outputs(5667) <= '0';
    layer2_outputs(5668) <= not a;
    layer2_outputs(5669) <= a and not b;
    layer2_outputs(5670) <= not b or a;
    layer2_outputs(5671) <= b;
    layer2_outputs(5672) <= not (a and b);
    layer2_outputs(5673) <= a and not b;
    layer2_outputs(5674) <= '0';
    layer2_outputs(5675) <= b;
    layer2_outputs(5676) <= a and not b;
    layer2_outputs(5677) <= a and b;
    layer2_outputs(5678) <= not a or b;
    layer2_outputs(5679) <= not b;
    layer2_outputs(5680) <= not (a and b);
    layer2_outputs(5681) <= a xor b;
    layer2_outputs(5682) <= '0';
    layer2_outputs(5683) <= not (a and b);
    layer2_outputs(5684) <= not (a xor b);
    layer2_outputs(5685) <= not (a or b);
    layer2_outputs(5686) <= not a;
    layer2_outputs(5687) <= a xor b;
    layer2_outputs(5688) <= not (a or b);
    layer2_outputs(5689) <= '0';
    layer2_outputs(5690) <= not b or a;
    layer2_outputs(5691) <= '1';
    layer2_outputs(5692) <= not b;
    layer2_outputs(5693) <= not a;
    layer2_outputs(5694) <= b and not a;
    layer2_outputs(5695) <= a xor b;
    layer2_outputs(5696) <= a or b;
    layer2_outputs(5697) <= b;
    layer2_outputs(5698) <= '0';
    layer2_outputs(5699) <= not b;
    layer2_outputs(5700) <= not a or b;
    layer2_outputs(5701) <= b and not a;
    layer2_outputs(5702) <= not (a or b);
    layer2_outputs(5703) <= not a or b;
    layer2_outputs(5704) <= b and not a;
    layer2_outputs(5705) <= a;
    layer2_outputs(5706) <= a and b;
    layer2_outputs(5707) <= b;
    layer2_outputs(5708) <= a or b;
    layer2_outputs(5709) <= not a or b;
    layer2_outputs(5710) <= b and not a;
    layer2_outputs(5711) <= not a;
    layer2_outputs(5712) <= b;
    layer2_outputs(5713) <= a and b;
    layer2_outputs(5714) <= not b or a;
    layer2_outputs(5715) <= b;
    layer2_outputs(5716) <= '0';
    layer2_outputs(5717) <= not a;
    layer2_outputs(5718) <= b;
    layer2_outputs(5719) <= not a or b;
    layer2_outputs(5720) <= b and not a;
    layer2_outputs(5721) <= not a;
    layer2_outputs(5722) <= not b or a;
    layer2_outputs(5723) <= not b or a;
    layer2_outputs(5724) <= not a;
    layer2_outputs(5725) <= not a or b;
    layer2_outputs(5726) <= b;
    layer2_outputs(5727) <= a and not b;
    layer2_outputs(5728) <= b;
    layer2_outputs(5729) <= not a or b;
    layer2_outputs(5730) <= b;
    layer2_outputs(5731) <= a and not b;
    layer2_outputs(5732) <= a xor b;
    layer2_outputs(5733) <= a and not b;
    layer2_outputs(5734) <= '1';
    layer2_outputs(5735) <= a;
    layer2_outputs(5736) <= not (a xor b);
    layer2_outputs(5737) <= a and b;
    layer2_outputs(5738) <= b and not a;
    layer2_outputs(5739) <= not a;
    layer2_outputs(5740) <= '0';
    layer2_outputs(5741) <= not a;
    layer2_outputs(5742) <= '0';
    layer2_outputs(5743) <= not b or a;
    layer2_outputs(5744) <= not (a or b);
    layer2_outputs(5745) <= a or b;
    layer2_outputs(5746) <= b;
    layer2_outputs(5747) <= not a;
    layer2_outputs(5748) <= '0';
    layer2_outputs(5749) <= b and not a;
    layer2_outputs(5750) <= b and not a;
    layer2_outputs(5751) <= not (a xor b);
    layer2_outputs(5752) <= a;
    layer2_outputs(5753) <= '0';
    layer2_outputs(5754) <= not (a or b);
    layer2_outputs(5755) <= not b or a;
    layer2_outputs(5756) <= b and not a;
    layer2_outputs(5757) <= a and b;
    layer2_outputs(5758) <= not a;
    layer2_outputs(5759) <= '1';
    layer2_outputs(5760) <= not a or b;
    layer2_outputs(5761) <= b;
    layer2_outputs(5762) <= not a;
    layer2_outputs(5763) <= not b or a;
    layer2_outputs(5764) <= not (a or b);
    layer2_outputs(5765) <= a;
    layer2_outputs(5766) <= not (a xor b);
    layer2_outputs(5767) <= not (a or b);
    layer2_outputs(5768) <= not (a and b);
    layer2_outputs(5769) <= '0';
    layer2_outputs(5770) <= a;
    layer2_outputs(5771) <= not b;
    layer2_outputs(5772) <= a;
    layer2_outputs(5773) <= a or b;
    layer2_outputs(5774) <= not b or a;
    layer2_outputs(5775) <= a;
    layer2_outputs(5776) <= not (a or b);
    layer2_outputs(5777) <= b and not a;
    layer2_outputs(5778) <= b and not a;
    layer2_outputs(5779) <= not a;
    layer2_outputs(5780) <= a and not b;
    layer2_outputs(5781) <= a xor b;
    layer2_outputs(5782) <= '0';
    layer2_outputs(5783) <= a or b;
    layer2_outputs(5784) <= not (a or b);
    layer2_outputs(5785) <= b and not a;
    layer2_outputs(5786) <= not b or a;
    layer2_outputs(5787) <= a and b;
    layer2_outputs(5788) <= a and b;
    layer2_outputs(5789) <= not a;
    layer2_outputs(5790) <= b and not a;
    layer2_outputs(5791) <= not b;
    layer2_outputs(5792) <= not (a and b);
    layer2_outputs(5793) <= not a or b;
    layer2_outputs(5794) <= b and not a;
    layer2_outputs(5795) <= b;
    layer2_outputs(5796) <= a and not b;
    layer2_outputs(5797) <= not b or a;
    layer2_outputs(5798) <= b and not a;
    layer2_outputs(5799) <= b;
    layer2_outputs(5800) <= not (a or b);
    layer2_outputs(5801) <= a and not b;
    layer2_outputs(5802) <= '1';
    layer2_outputs(5803) <= not b or a;
    layer2_outputs(5804) <= a or b;
    layer2_outputs(5805) <= a;
    layer2_outputs(5806) <= '1';
    layer2_outputs(5807) <= a or b;
    layer2_outputs(5808) <= a and b;
    layer2_outputs(5809) <= a;
    layer2_outputs(5810) <= not (a or b);
    layer2_outputs(5811) <= not (a and b);
    layer2_outputs(5812) <= a;
    layer2_outputs(5813) <= not b;
    layer2_outputs(5814) <= not (a and b);
    layer2_outputs(5815) <= not (a or b);
    layer2_outputs(5816) <= '1';
    layer2_outputs(5817) <= a and b;
    layer2_outputs(5818) <= not (a and b);
    layer2_outputs(5819) <= b;
    layer2_outputs(5820) <= '1';
    layer2_outputs(5821) <= not b;
    layer2_outputs(5822) <= not (a xor b);
    layer2_outputs(5823) <= not b or a;
    layer2_outputs(5824) <= b and not a;
    layer2_outputs(5825) <= a and b;
    layer2_outputs(5826) <= not (a or b);
    layer2_outputs(5827) <= b and not a;
    layer2_outputs(5828) <= not b;
    layer2_outputs(5829) <= not (a or b);
    layer2_outputs(5830) <= b;
    layer2_outputs(5831) <= b;
    layer2_outputs(5832) <= not (a xor b);
    layer2_outputs(5833) <= not b;
    layer2_outputs(5834) <= a and b;
    layer2_outputs(5835) <= b;
    layer2_outputs(5836) <= not b;
    layer2_outputs(5837) <= b and not a;
    layer2_outputs(5838) <= a or b;
    layer2_outputs(5839) <= not a;
    layer2_outputs(5840) <= a and b;
    layer2_outputs(5841) <= not b;
    layer2_outputs(5842) <= a and not b;
    layer2_outputs(5843) <= not b or a;
    layer2_outputs(5844) <= a and not b;
    layer2_outputs(5845) <= not a;
    layer2_outputs(5846) <= not (a xor b);
    layer2_outputs(5847) <= not a or b;
    layer2_outputs(5848) <= not a;
    layer2_outputs(5849) <= b and not a;
    layer2_outputs(5850) <= a or b;
    layer2_outputs(5851) <= '1';
    layer2_outputs(5852) <= not a;
    layer2_outputs(5853) <= not (a and b);
    layer2_outputs(5854) <= b;
    layer2_outputs(5855) <= b;
    layer2_outputs(5856) <= not (a and b);
    layer2_outputs(5857) <= a and b;
    layer2_outputs(5858) <= '0';
    layer2_outputs(5859) <= a or b;
    layer2_outputs(5860) <= a;
    layer2_outputs(5861) <= not a or b;
    layer2_outputs(5862) <= not a;
    layer2_outputs(5863) <= not a or b;
    layer2_outputs(5864) <= not b or a;
    layer2_outputs(5865) <= a or b;
    layer2_outputs(5866) <= not a or b;
    layer2_outputs(5867) <= b and not a;
    layer2_outputs(5868) <= a xor b;
    layer2_outputs(5869) <= '0';
    layer2_outputs(5870) <= not a;
    layer2_outputs(5871) <= not a or b;
    layer2_outputs(5872) <= not a or b;
    layer2_outputs(5873) <= b;
    layer2_outputs(5874) <= not a or b;
    layer2_outputs(5875) <= not b or a;
    layer2_outputs(5876) <= not a;
    layer2_outputs(5877) <= '0';
    layer2_outputs(5878) <= a;
    layer2_outputs(5879) <= not (a xor b);
    layer2_outputs(5880) <= '0';
    layer2_outputs(5881) <= b;
    layer2_outputs(5882) <= not (a xor b);
    layer2_outputs(5883) <= a;
    layer2_outputs(5884) <= not a;
    layer2_outputs(5885) <= a and not b;
    layer2_outputs(5886) <= not a or b;
    layer2_outputs(5887) <= not (a or b);
    layer2_outputs(5888) <= a or b;
    layer2_outputs(5889) <= '0';
    layer2_outputs(5890) <= a and not b;
    layer2_outputs(5891) <= a;
    layer2_outputs(5892) <= a and not b;
    layer2_outputs(5893) <= not a or b;
    layer2_outputs(5894) <= '1';
    layer2_outputs(5895) <= '0';
    layer2_outputs(5896) <= not a or b;
    layer2_outputs(5897) <= a;
    layer2_outputs(5898) <= not (a and b);
    layer2_outputs(5899) <= not b;
    layer2_outputs(5900) <= a xor b;
    layer2_outputs(5901) <= not b or a;
    layer2_outputs(5902) <= b and not a;
    layer2_outputs(5903) <= '0';
    layer2_outputs(5904) <= a and not b;
    layer2_outputs(5905) <= not (a xor b);
    layer2_outputs(5906) <= '1';
    layer2_outputs(5907) <= '1';
    layer2_outputs(5908) <= a;
    layer2_outputs(5909) <= b;
    layer2_outputs(5910) <= not (a and b);
    layer2_outputs(5911) <= b;
    layer2_outputs(5912) <= not b or a;
    layer2_outputs(5913) <= not a;
    layer2_outputs(5914) <= not b or a;
    layer2_outputs(5915) <= a and b;
    layer2_outputs(5916) <= a xor b;
    layer2_outputs(5917) <= a;
    layer2_outputs(5918) <= not a;
    layer2_outputs(5919) <= not (a and b);
    layer2_outputs(5920) <= a;
    layer2_outputs(5921) <= not b or a;
    layer2_outputs(5922) <= not a or b;
    layer2_outputs(5923) <= '1';
    layer2_outputs(5924) <= a xor b;
    layer2_outputs(5925) <= a;
    layer2_outputs(5926) <= not a or b;
    layer2_outputs(5927) <= '0';
    layer2_outputs(5928) <= a;
    layer2_outputs(5929) <= '1';
    layer2_outputs(5930) <= '0';
    layer2_outputs(5931) <= not b;
    layer2_outputs(5932) <= '1';
    layer2_outputs(5933) <= not a or b;
    layer2_outputs(5934) <= not (a or b);
    layer2_outputs(5935) <= a xor b;
    layer2_outputs(5936) <= b;
    layer2_outputs(5937) <= a or b;
    layer2_outputs(5938) <= not a;
    layer2_outputs(5939) <= not b;
    layer2_outputs(5940) <= not (a or b);
    layer2_outputs(5941) <= not b;
    layer2_outputs(5942) <= a or b;
    layer2_outputs(5943) <= '1';
    layer2_outputs(5944) <= a xor b;
    layer2_outputs(5945) <= not a or b;
    layer2_outputs(5946) <= a;
    layer2_outputs(5947) <= not a;
    layer2_outputs(5948) <= b;
    layer2_outputs(5949) <= not b;
    layer2_outputs(5950) <= a and b;
    layer2_outputs(5951) <= not b;
    layer2_outputs(5952) <= not b or a;
    layer2_outputs(5953) <= not a;
    layer2_outputs(5954) <= '0';
    layer2_outputs(5955) <= not b or a;
    layer2_outputs(5956) <= b;
    layer2_outputs(5957) <= a and b;
    layer2_outputs(5958) <= not b;
    layer2_outputs(5959) <= '1';
    layer2_outputs(5960) <= not (a and b);
    layer2_outputs(5961) <= a and b;
    layer2_outputs(5962) <= a;
    layer2_outputs(5963) <= not (a and b);
    layer2_outputs(5964) <= a and not b;
    layer2_outputs(5965) <= not a;
    layer2_outputs(5966) <= b;
    layer2_outputs(5967) <= a and not b;
    layer2_outputs(5968) <= not a;
    layer2_outputs(5969) <= '1';
    layer2_outputs(5970) <= not b or a;
    layer2_outputs(5971) <= not (a or b);
    layer2_outputs(5972) <= '0';
    layer2_outputs(5973) <= '0';
    layer2_outputs(5974) <= not b or a;
    layer2_outputs(5975) <= not (a and b);
    layer2_outputs(5976) <= not b;
    layer2_outputs(5977) <= a;
    layer2_outputs(5978) <= not b;
    layer2_outputs(5979) <= not b or a;
    layer2_outputs(5980) <= not (a and b);
    layer2_outputs(5981) <= '0';
    layer2_outputs(5982) <= not a or b;
    layer2_outputs(5983) <= b and not a;
    layer2_outputs(5984) <= not a;
    layer2_outputs(5985) <= '0';
    layer2_outputs(5986) <= not b or a;
    layer2_outputs(5987) <= '0';
    layer2_outputs(5988) <= not b or a;
    layer2_outputs(5989) <= a and not b;
    layer2_outputs(5990) <= not a;
    layer2_outputs(5991) <= not b;
    layer2_outputs(5992) <= not b or a;
    layer2_outputs(5993) <= not b;
    layer2_outputs(5994) <= '1';
    layer2_outputs(5995) <= a;
    layer2_outputs(5996) <= not b or a;
    layer2_outputs(5997) <= a;
    layer2_outputs(5998) <= b and not a;
    layer2_outputs(5999) <= '1';
    layer2_outputs(6000) <= b;
    layer2_outputs(6001) <= not a;
    layer2_outputs(6002) <= not b;
    layer2_outputs(6003) <= b;
    layer2_outputs(6004) <= '1';
    layer2_outputs(6005) <= not b or a;
    layer2_outputs(6006) <= '1';
    layer2_outputs(6007) <= not a;
    layer2_outputs(6008) <= '0';
    layer2_outputs(6009) <= a and not b;
    layer2_outputs(6010) <= '1';
    layer2_outputs(6011) <= not b or a;
    layer2_outputs(6012) <= a and b;
    layer2_outputs(6013) <= not a or b;
    layer2_outputs(6014) <= not b;
    layer2_outputs(6015) <= a;
    layer2_outputs(6016) <= not a or b;
    layer2_outputs(6017) <= not b or a;
    layer2_outputs(6018) <= not (a or b);
    layer2_outputs(6019) <= a;
    layer2_outputs(6020) <= not (a and b);
    layer2_outputs(6021) <= not (a or b);
    layer2_outputs(6022) <= not (a or b);
    layer2_outputs(6023) <= a and b;
    layer2_outputs(6024) <= a;
    layer2_outputs(6025) <= not b;
    layer2_outputs(6026) <= not a or b;
    layer2_outputs(6027) <= not (a and b);
    layer2_outputs(6028) <= a or b;
    layer2_outputs(6029) <= not (a or b);
    layer2_outputs(6030) <= not a;
    layer2_outputs(6031) <= '1';
    layer2_outputs(6032) <= a;
    layer2_outputs(6033) <= '0';
    layer2_outputs(6034) <= b;
    layer2_outputs(6035) <= a;
    layer2_outputs(6036) <= a or b;
    layer2_outputs(6037) <= a and b;
    layer2_outputs(6038) <= a;
    layer2_outputs(6039) <= b;
    layer2_outputs(6040) <= not b;
    layer2_outputs(6041) <= b;
    layer2_outputs(6042) <= b;
    layer2_outputs(6043) <= a and b;
    layer2_outputs(6044) <= not a;
    layer2_outputs(6045) <= not a;
    layer2_outputs(6046) <= not a;
    layer2_outputs(6047) <= a or b;
    layer2_outputs(6048) <= '0';
    layer2_outputs(6049) <= a and not b;
    layer2_outputs(6050) <= not b or a;
    layer2_outputs(6051) <= not a;
    layer2_outputs(6052) <= not (a or b);
    layer2_outputs(6053) <= not b;
    layer2_outputs(6054) <= not a;
    layer2_outputs(6055) <= b;
    layer2_outputs(6056) <= not a;
    layer2_outputs(6057) <= not (a and b);
    layer2_outputs(6058) <= b;
    layer2_outputs(6059) <= '1';
    layer2_outputs(6060) <= not b;
    layer2_outputs(6061) <= not (a and b);
    layer2_outputs(6062) <= not a or b;
    layer2_outputs(6063) <= not (a and b);
    layer2_outputs(6064) <= not b or a;
    layer2_outputs(6065) <= a and b;
    layer2_outputs(6066) <= a or b;
    layer2_outputs(6067) <= a;
    layer2_outputs(6068) <= not (a and b);
    layer2_outputs(6069) <= a;
    layer2_outputs(6070) <= b and not a;
    layer2_outputs(6071) <= a and not b;
    layer2_outputs(6072) <= b;
    layer2_outputs(6073) <= not a;
    layer2_outputs(6074) <= '0';
    layer2_outputs(6075) <= not (a or b);
    layer2_outputs(6076) <= '0';
    layer2_outputs(6077) <= b;
    layer2_outputs(6078) <= not b;
    layer2_outputs(6079) <= b;
    layer2_outputs(6080) <= not a or b;
    layer2_outputs(6081) <= a and not b;
    layer2_outputs(6082) <= a and b;
    layer2_outputs(6083) <= b and not a;
    layer2_outputs(6084) <= not b;
    layer2_outputs(6085) <= not b;
    layer2_outputs(6086) <= not b;
    layer2_outputs(6087) <= not a or b;
    layer2_outputs(6088) <= a and b;
    layer2_outputs(6089) <= b and not a;
    layer2_outputs(6090) <= a xor b;
    layer2_outputs(6091) <= not b;
    layer2_outputs(6092) <= b;
    layer2_outputs(6093) <= not a;
    layer2_outputs(6094) <= a or b;
    layer2_outputs(6095) <= b;
    layer2_outputs(6096) <= not b;
    layer2_outputs(6097) <= not (a and b);
    layer2_outputs(6098) <= a and b;
    layer2_outputs(6099) <= '0';
    layer2_outputs(6100) <= not a;
    layer2_outputs(6101) <= a and b;
    layer2_outputs(6102) <= b;
    layer2_outputs(6103) <= not a or b;
    layer2_outputs(6104) <= not b;
    layer2_outputs(6105) <= '0';
    layer2_outputs(6106) <= '1';
    layer2_outputs(6107) <= b;
    layer2_outputs(6108) <= a and not b;
    layer2_outputs(6109) <= not a;
    layer2_outputs(6110) <= b;
    layer2_outputs(6111) <= a xor b;
    layer2_outputs(6112) <= b;
    layer2_outputs(6113) <= not (a and b);
    layer2_outputs(6114) <= not b;
    layer2_outputs(6115) <= '1';
    layer2_outputs(6116) <= '1';
    layer2_outputs(6117) <= not (a xor b);
    layer2_outputs(6118) <= a or b;
    layer2_outputs(6119) <= not b or a;
    layer2_outputs(6120) <= not b;
    layer2_outputs(6121) <= not b;
    layer2_outputs(6122) <= not (a or b);
    layer2_outputs(6123) <= not a;
    layer2_outputs(6124) <= b;
    layer2_outputs(6125) <= not a or b;
    layer2_outputs(6126) <= a or b;
    layer2_outputs(6127) <= a;
    layer2_outputs(6128) <= '1';
    layer2_outputs(6129) <= not a;
    layer2_outputs(6130) <= not a or b;
    layer2_outputs(6131) <= a;
    layer2_outputs(6132) <= not b;
    layer2_outputs(6133) <= b;
    layer2_outputs(6134) <= not (a xor b);
    layer2_outputs(6135) <= a and b;
    layer2_outputs(6136) <= a or b;
    layer2_outputs(6137) <= not (a and b);
    layer2_outputs(6138) <= not (a and b);
    layer2_outputs(6139) <= not (a and b);
    layer2_outputs(6140) <= b;
    layer2_outputs(6141) <= b and not a;
    layer2_outputs(6142) <= '1';
    layer2_outputs(6143) <= a and b;
    layer2_outputs(6144) <= '1';
    layer2_outputs(6145) <= b and not a;
    layer2_outputs(6146) <= a or b;
    layer2_outputs(6147) <= a;
    layer2_outputs(6148) <= a or b;
    layer2_outputs(6149) <= '0';
    layer2_outputs(6150) <= not (a xor b);
    layer2_outputs(6151) <= a and not b;
    layer2_outputs(6152) <= not (a or b);
    layer2_outputs(6153) <= not a;
    layer2_outputs(6154) <= a;
    layer2_outputs(6155) <= not a or b;
    layer2_outputs(6156) <= not (a and b);
    layer2_outputs(6157) <= b;
    layer2_outputs(6158) <= '0';
    layer2_outputs(6159) <= a and b;
    layer2_outputs(6160) <= b;
    layer2_outputs(6161) <= b;
    layer2_outputs(6162) <= a xor b;
    layer2_outputs(6163) <= not (a or b);
    layer2_outputs(6164) <= not b;
    layer2_outputs(6165) <= not (a or b);
    layer2_outputs(6166) <= not a;
    layer2_outputs(6167) <= a xor b;
    layer2_outputs(6168) <= b;
    layer2_outputs(6169) <= a and b;
    layer2_outputs(6170) <= b;
    layer2_outputs(6171) <= a or b;
    layer2_outputs(6172) <= a and b;
    layer2_outputs(6173) <= not (a and b);
    layer2_outputs(6174) <= a and b;
    layer2_outputs(6175) <= not b or a;
    layer2_outputs(6176) <= not a;
    layer2_outputs(6177) <= '1';
    layer2_outputs(6178) <= not (a or b);
    layer2_outputs(6179) <= not (a or b);
    layer2_outputs(6180) <= not b or a;
    layer2_outputs(6181) <= '0';
    layer2_outputs(6182) <= not (a xor b);
    layer2_outputs(6183) <= not b or a;
    layer2_outputs(6184) <= a;
    layer2_outputs(6185) <= not (a and b);
    layer2_outputs(6186) <= not b;
    layer2_outputs(6187) <= b;
    layer2_outputs(6188) <= not (a or b);
    layer2_outputs(6189) <= a xor b;
    layer2_outputs(6190) <= '0';
    layer2_outputs(6191) <= a;
    layer2_outputs(6192) <= not b or a;
    layer2_outputs(6193) <= not (a and b);
    layer2_outputs(6194) <= a and not b;
    layer2_outputs(6195) <= not b;
    layer2_outputs(6196) <= a;
    layer2_outputs(6197) <= a;
    layer2_outputs(6198) <= not b;
    layer2_outputs(6199) <= a xor b;
    layer2_outputs(6200) <= not (a or b);
    layer2_outputs(6201) <= b;
    layer2_outputs(6202) <= '0';
    layer2_outputs(6203) <= a and b;
    layer2_outputs(6204) <= a and b;
    layer2_outputs(6205) <= b;
    layer2_outputs(6206) <= not b or a;
    layer2_outputs(6207) <= a and b;
    layer2_outputs(6208) <= not a;
    layer2_outputs(6209) <= a and not b;
    layer2_outputs(6210) <= not a;
    layer2_outputs(6211) <= a and b;
    layer2_outputs(6212) <= not (a and b);
    layer2_outputs(6213) <= b;
    layer2_outputs(6214) <= a or b;
    layer2_outputs(6215) <= not b;
    layer2_outputs(6216) <= not a;
    layer2_outputs(6217) <= not (a or b);
    layer2_outputs(6218) <= not (a and b);
    layer2_outputs(6219) <= not b;
    layer2_outputs(6220) <= b and not a;
    layer2_outputs(6221) <= not b;
    layer2_outputs(6222) <= a;
    layer2_outputs(6223) <= not a;
    layer2_outputs(6224) <= not b or a;
    layer2_outputs(6225) <= a and b;
    layer2_outputs(6226) <= not a;
    layer2_outputs(6227) <= not a or b;
    layer2_outputs(6228) <= not a;
    layer2_outputs(6229) <= a;
    layer2_outputs(6230) <= not a or b;
    layer2_outputs(6231) <= a;
    layer2_outputs(6232) <= b;
    layer2_outputs(6233) <= not (a and b);
    layer2_outputs(6234) <= a or b;
    layer2_outputs(6235) <= not a or b;
    layer2_outputs(6236) <= not a;
    layer2_outputs(6237) <= not b or a;
    layer2_outputs(6238) <= a or b;
    layer2_outputs(6239) <= a or b;
    layer2_outputs(6240) <= b and not a;
    layer2_outputs(6241) <= a xor b;
    layer2_outputs(6242) <= b and not a;
    layer2_outputs(6243) <= a and b;
    layer2_outputs(6244) <= not (a xor b);
    layer2_outputs(6245) <= a and not b;
    layer2_outputs(6246) <= a and b;
    layer2_outputs(6247) <= not b or a;
    layer2_outputs(6248) <= a and not b;
    layer2_outputs(6249) <= b and not a;
    layer2_outputs(6250) <= a;
    layer2_outputs(6251) <= a;
    layer2_outputs(6252) <= not b or a;
    layer2_outputs(6253) <= '0';
    layer2_outputs(6254) <= '1';
    layer2_outputs(6255) <= a;
    layer2_outputs(6256) <= a xor b;
    layer2_outputs(6257) <= not b or a;
    layer2_outputs(6258) <= not (a or b);
    layer2_outputs(6259) <= not (a xor b);
    layer2_outputs(6260) <= '1';
    layer2_outputs(6261) <= b;
    layer2_outputs(6262) <= not (a or b);
    layer2_outputs(6263) <= a and b;
    layer2_outputs(6264) <= not a;
    layer2_outputs(6265) <= not (a or b);
    layer2_outputs(6266) <= a and not b;
    layer2_outputs(6267) <= a and not b;
    layer2_outputs(6268) <= not (a or b);
    layer2_outputs(6269) <= not (a and b);
    layer2_outputs(6270) <= a and not b;
    layer2_outputs(6271) <= not (a and b);
    layer2_outputs(6272) <= '0';
    layer2_outputs(6273) <= not a;
    layer2_outputs(6274) <= a and b;
    layer2_outputs(6275) <= b;
    layer2_outputs(6276) <= not (a or b);
    layer2_outputs(6277) <= b and not a;
    layer2_outputs(6278) <= not a;
    layer2_outputs(6279) <= not (a xor b);
    layer2_outputs(6280) <= not (a and b);
    layer2_outputs(6281) <= a;
    layer2_outputs(6282) <= '0';
    layer2_outputs(6283) <= '0';
    layer2_outputs(6284) <= b and not a;
    layer2_outputs(6285) <= not (a and b);
    layer2_outputs(6286) <= not b;
    layer2_outputs(6287) <= a or b;
    layer2_outputs(6288) <= b;
    layer2_outputs(6289) <= not b;
    layer2_outputs(6290) <= a and b;
    layer2_outputs(6291) <= a and b;
    layer2_outputs(6292) <= a or b;
    layer2_outputs(6293) <= b;
    layer2_outputs(6294) <= not a or b;
    layer2_outputs(6295) <= not b or a;
    layer2_outputs(6296) <= not a;
    layer2_outputs(6297) <= a and b;
    layer2_outputs(6298) <= b;
    layer2_outputs(6299) <= not a;
    layer2_outputs(6300) <= not (a and b);
    layer2_outputs(6301) <= a or b;
    layer2_outputs(6302) <= not (a or b);
    layer2_outputs(6303) <= not b;
    layer2_outputs(6304) <= a xor b;
    layer2_outputs(6305) <= not a;
    layer2_outputs(6306) <= a;
    layer2_outputs(6307) <= not (a or b);
    layer2_outputs(6308) <= not a or b;
    layer2_outputs(6309) <= not a or b;
    layer2_outputs(6310) <= a or b;
    layer2_outputs(6311) <= not (a or b);
    layer2_outputs(6312) <= b;
    layer2_outputs(6313) <= not (a and b);
    layer2_outputs(6314) <= not (a or b);
    layer2_outputs(6315) <= a and b;
    layer2_outputs(6316) <= '0';
    layer2_outputs(6317) <= not b or a;
    layer2_outputs(6318) <= a and not b;
    layer2_outputs(6319) <= b and not a;
    layer2_outputs(6320) <= not b;
    layer2_outputs(6321) <= a and b;
    layer2_outputs(6322) <= '0';
    layer2_outputs(6323) <= not (a or b);
    layer2_outputs(6324) <= a or b;
    layer2_outputs(6325) <= not (a and b);
    layer2_outputs(6326) <= not (a and b);
    layer2_outputs(6327) <= a and b;
    layer2_outputs(6328) <= not (a or b);
    layer2_outputs(6329) <= not a;
    layer2_outputs(6330) <= not (a or b);
    layer2_outputs(6331) <= b and not a;
    layer2_outputs(6332) <= not a or b;
    layer2_outputs(6333) <= b;
    layer2_outputs(6334) <= a and b;
    layer2_outputs(6335) <= a;
    layer2_outputs(6336) <= a and b;
    layer2_outputs(6337) <= a xor b;
    layer2_outputs(6338) <= not (a or b);
    layer2_outputs(6339) <= '0';
    layer2_outputs(6340) <= not a or b;
    layer2_outputs(6341) <= not (a and b);
    layer2_outputs(6342) <= a or b;
    layer2_outputs(6343) <= not a or b;
    layer2_outputs(6344) <= not b;
    layer2_outputs(6345) <= b and not a;
    layer2_outputs(6346) <= b;
    layer2_outputs(6347) <= not b;
    layer2_outputs(6348) <= a xor b;
    layer2_outputs(6349) <= a and b;
    layer2_outputs(6350) <= not a;
    layer2_outputs(6351) <= a or b;
    layer2_outputs(6352) <= not (a and b);
    layer2_outputs(6353) <= a and not b;
    layer2_outputs(6354) <= not a or b;
    layer2_outputs(6355) <= not a or b;
    layer2_outputs(6356) <= not b;
    layer2_outputs(6357) <= b;
    layer2_outputs(6358) <= not (a or b);
    layer2_outputs(6359) <= a or b;
    layer2_outputs(6360) <= a or b;
    layer2_outputs(6361) <= not a or b;
    layer2_outputs(6362) <= not a;
    layer2_outputs(6363) <= a or b;
    layer2_outputs(6364) <= a xor b;
    layer2_outputs(6365) <= not b or a;
    layer2_outputs(6366) <= not a or b;
    layer2_outputs(6367) <= a or b;
    layer2_outputs(6368) <= a;
    layer2_outputs(6369) <= not a;
    layer2_outputs(6370) <= not (a xor b);
    layer2_outputs(6371) <= a;
    layer2_outputs(6372) <= not b;
    layer2_outputs(6373) <= not b;
    layer2_outputs(6374) <= a and not b;
    layer2_outputs(6375) <= not b;
    layer2_outputs(6376) <= not a or b;
    layer2_outputs(6377) <= b and not a;
    layer2_outputs(6378) <= not (a or b);
    layer2_outputs(6379) <= '0';
    layer2_outputs(6380) <= not a;
    layer2_outputs(6381) <= not a or b;
    layer2_outputs(6382) <= not (a or b);
    layer2_outputs(6383) <= not (a and b);
    layer2_outputs(6384) <= a and not b;
    layer2_outputs(6385) <= not b or a;
    layer2_outputs(6386) <= not (a and b);
    layer2_outputs(6387) <= a xor b;
    layer2_outputs(6388) <= a and not b;
    layer2_outputs(6389) <= not (a xor b);
    layer2_outputs(6390) <= '1';
    layer2_outputs(6391) <= not b;
    layer2_outputs(6392) <= not (a and b);
    layer2_outputs(6393) <= a or b;
    layer2_outputs(6394) <= '0';
    layer2_outputs(6395) <= a xor b;
    layer2_outputs(6396) <= not (a xor b);
    layer2_outputs(6397) <= b and not a;
    layer2_outputs(6398) <= a or b;
    layer2_outputs(6399) <= a;
    layer2_outputs(6400) <= b;
    layer2_outputs(6401) <= a;
    layer2_outputs(6402) <= b and not a;
    layer2_outputs(6403) <= not a or b;
    layer2_outputs(6404) <= b and not a;
    layer2_outputs(6405) <= not (a xor b);
    layer2_outputs(6406) <= a and b;
    layer2_outputs(6407) <= not b or a;
    layer2_outputs(6408) <= a and not b;
    layer2_outputs(6409) <= not a or b;
    layer2_outputs(6410) <= a xor b;
    layer2_outputs(6411) <= a xor b;
    layer2_outputs(6412) <= not a or b;
    layer2_outputs(6413) <= not b or a;
    layer2_outputs(6414) <= a and b;
    layer2_outputs(6415) <= not b or a;
    layer2_outputs(6416) <= a or b;
    layer2_outputs(6417) <= not a;
    layer2_outputs(6418) <= a and not b;
    layer2_outputs(6419) <= a;
    layer2_outputs(6420) <= '0';
    layer2_outputs(6421) <= not (a or b);
    layer2_outputs(6422) <= not a or b;
    layer2_outputs(6423) <= b and not a;
    layer2_outputs(6424) <= not b or a;
    layer2_outputs(6425) <= a and b;
    layer2_outputs(6426) <= a and b;
    layer2_outputs(6427) <= not b;
    layer2_outputs(6428) <= a and not b;
    layer2_outputs(6429) <= not b;
    layer2_outputs(6430) <= not a or b;
    layer2_outputs(6431) <= a and not b;
    layer2_outputs(6432) <= not b;
    layer2_outputs(6433) <= a;
    layer2_outputs(6434) <= b;
    layer2_outputs(6435) <= not b;
    layer2_outputs(6436) <= b and not a;
    layer2_outputs(6437) <= not (a and b);
    layer2_outputs(6438) <= not a or b;
    layer2_outputs(6439) <= not b;
    layer2_outputs(6440) <= a;
    layer2_outputs(6441) <= a;
    layer2_outputs(6442) <= not a or b;
    layer2_outputs(6443) <= not b;
    layer2_outputs(6444) <= b;
    layer2_outputs(6445) <= '0';
    layer2_outputs(6446) <= not (a xor b);
    layer2_outputs(6447) <= a and not b;
    layer2_outputs(6448) <= not b;
    layer2_outputs(6449) <= '0';
    layer2_outputs(6450) <= '1';
    layer2_outputs(6451) <= not (a and b);
    layer2_outputs(6452) <= a xor b;
    layer2_outputs(6453) <= a and not b;
    layer2_outputs(6454) <= a and not b;
    layer2_outputs(6455) <= a and not b;
    layer2_outputs(6456) <= a xor b;
    layer2_outputs(6457) <= not b or a;
    layer2_outputs(6458) <= not b;
    layer2_outputs(6459) <= a or b;
    layer2_outputs(6460) <= b and not a;
    layer2_outputs(6461) <= not a;
    layer2_outputs(6462) <= not a or b;
    layer2_outputs(6463) <= a and b;
    layer2_outputs(6464) <= '0';
    layer2_outputs(6465) <= a and not b;
    layer2_outputs(6466) <= not b;
    layer2_outputs(6467) <= not b or a;
    layer2_outputs(6468) <= not b;
    layer2_outputs(6469) <= '1';
    layer2_outputs(6470) <= a;
    layer2_outputs(6471) <= not b;
    layer2_outputs(6472) <= not a;
    layer2_outputs(6473) <= b and not a;
    layer2_outputs(6474) <= not a or b;
    layer2_outputs(6475) <= not a;
    layer2_outputs(6476) <= a xor b;
    layer2_outputs(6477) <= '1';
    layer2_outputs(6478) <= a;
    layer2_outputs(6479) <= not (a and b);
    layer2_outputs(6480) <= b;
    layer2_outputs(6481) <= a or b;
    layer2_outputs(6482) <= not a;
    layer2_outputs(6483) <= not (a and b);
    layer2_outputs(6484) <= not b;
    layer2_outputs(6485) <= a and not b;
    layer2_outputs(6486) <= a or b;
    layer2_outputs(6487) <= not b;
    layer2_outputs(6488) <= not (a and b);
    layer2_outputs(6489) <= a xor b;
    layer2_outputs(6490) <= not b;
    layer2_outputs(6491) <= not a;
    layer2_outputs(6492) <= not b;
    layer2_outputs(6493) <= a and not b;
    layer2_outputs(6494) <= b;
    layer2_outputs(6495) <= not (a and b);
    layer2_outputs(6496) <= not b;
    layer2_outputs(6497) <= '1';
    layer2_outputs(6498) <= not b or a;
    layer2_outputs(6499) <= not b;
    layer2_outputs(6500) <= '0';
    layer2_outputs(6501) <= not b;
    layer2_outputs(6502) <= not (a or b);
    layer2_outputs(6503) <= not (a or b);
    layer2_outputs(6504) <= '0';
    layer2_outputs(6505) <= a and b;
    layer2_outputs(6506) <= a or b;
    layer2_outputs(6507) <= '1';
    layer2_outputs(6508) <= not (a or b);
    layer2_outputs(6509) <= not a or b;
    layer2_outputs(6510) <= b;
    layer2_outputs(6511) <= a;
    layer2_outputs(6512) <= b and not a;
    layer2_outputs(6513) <= not (a or b);
    layer2_outputs(6514) <= not (a or b);
    layer2_outputs(6515) <= '0';
    layer2_outputs(6516) <= not a;
    layer2_outputs(6517) <= a and b;
    layer2_outputs(6518) <= not b or a;
    layer2_outputs(6519) <= a and b;
    layer2_outputs(6520) <= not (a or b);
    layer2_outputs(6521) <= not (a or b);
    layer2_outputs(6522) <= not a;
    layer2_outputs(6523) <= not a;
    layer2_outputs(6524) <= '0';
    layer2_outputs(6525) <= a xor b;
    layer2_outputs(6526) <= a and not b;
    layer2_outputs(6527) <= a or b;
    layer2_outputs(6528) <= a or b;
    layer2_outputs(6529) <= not a;
    layer2_outputs(6530) <= not b or a;
    layer2_outputs(6531) <= a;
    layer2_outputs(6532) <= '1';
    layer2_outputs(6533) <= not (a and b);
    layer2_outputs(6534) <= not b or a;
    layer2_outputs(6535) <= a;
    layer2_outputs(6536) <= not a or b;
    layer2_outputs(6537) <= not b;
    layer2_outputs(6538) <= not a or b;
    layer2_outputs(6539) <= not (a and b);
    layer2_outputs(6540) <= a or b;
    layer2_outputs(6541) <= '1';
    layer2_outputs(6542) <= not b or a;
    layer2_outputs(6543) <= not a;
    layer2_outputs(6544) <= a and b;
    layer2_outputs(6545) <= a or b;
    layer2_outputs(6546) <= a;
    layer2_outputs(6547) <= '0';
    layer2_outputs(6548) <= not a or b;
    layer2_outputs(6549) <= not b or a;
    layer2_outputs(6550) <= not a or b;
    layer2_outputs(6551) <= not (a xor b);
    layer2_outputs(6552) <= '1';
    layer2_outputs(6553) <= a and b;
    layer2_outputs(6554) <= a;
    layer2_outputs(6555) <= a;
    layer2_outputs(6556) <= not (a xor b);
    layer2_outputs(6557) <= a or b;
    layer2_outputs(6558) <= b and not a;
    layer2_outputs(6559) <= a or b;
    layer2_outputs(6560) <= not a;
    layer2_outputs(6561) <= '1';
    layer2_outputs(6562) <= a and b;
    layer2_outputs(6563) <= not a or b;
    layer2_outputs(6564) <= a or b;
    layer2_outputs(6565) <= not a;
    layer2_outputs(6566) <= '0';
    layer2_outputs(6567) <= b;
    layer2_outputs(6568) <= not (a xor b);
    layer2_outputs(6569) <= not (a and b);
    layer2_outputs(6570) <= not b or a;
    layer2_outputs(6571) <= b and not a;
    layer2_outputs(6572) <= '1';
    layer2_outputs(6573) <= a;
    layer2_outputs(6574) <= a;
    layer2_outputs(6575) <= a and b;
    layer2_outputs(6576) <= a or b;
    layer2_outputs(6577) <= b and not a;
    layer2_outputs(6578) <= a or b;
    layer2_outputs(6579) <= a;
    layer2_outputs(6580) <= a and b;
    layer2_outputs(6581) <= not a or b;
    layer2_outputs(6582) <= a;
    layer2_outputs(6583) <= b;
    layer2_outputs(6584) <= a or b;
    layer2_outputs(6585) <= not (a and b);
    layer2_outputs(6586) <= not b;
    layer2_outputs(6587) <= a and not b;
    layer2_outputs(6588) <= a and b;
    layer2_outputs(6589) <= not a or b;
    layer2_outputs(6590) <= not (a xor b);
    layer2_outputs(6591) <= a and b;
    layer2_outputs(6592) <= not a;
    layer2_outputs(6593) <= not b;
    layer2_outputs(6594) <= not (a and b);
    layer2_outputs(6595) <= not b;
    layer2_outputs(6596) <= not a or b;
    layer2_outputs(6597) <= a or b;
    layer2_outputs(6598) <= '1';
    layer2_outputs(6599) <= '1';
    layer2_outputs(6600) <= a;
    layer2_outputs(6601) <= not (a or b);
    layer2_outputs(6602) <= a;
    layer2_outputs(6603) <= a;
    layer2_outputs(6604) <= a or b;
    layer2_outputs(6605) <= not (a and b);
    layer2_outputs(6606) <= not a;
    layer2_outputs(6607) <= '1';
    layer2_outputs(6608) <= not a or b;
    layer2_outputs(6609) <= not (a and b);
    layer2_outputs(6610) <= a xor b;
    layer2_outputs(6611) <= a and b;
    layer2_outputs(6612) <= '1';
    layer2_outputs(6613) <= a;
    layer2_outputs(6614) <= b and not a;
    layer2_outputs(6615) <= b;
    layer2_outputs(6616) <= not a or b;
    layer2_outputs(6617) <= not a;
    layer2_outputs(6618) <= not b or a;
    layer2_outputs(6619) <= a and not b;
    layer2_outputs(6620) <= not (a or b);
    layer2_outputs(6621) <= '0';
    layer2_outputs(6622) <= '0';
    layer2_outputs(6623) <= not a;
    layer2_outputs(6624) <= b and not a;
    layer2_outputs(6625) <= a and not b;
    layer2_outputs(6626) <= b and not a;
    layer2_outputs(6627) <= b and not a;
    layer2_outputs(6628) <= b;
    layer2_outputs(6629) <= '1';
    layer2_outputs(6630) <= a or b;
    layer2_outputs(6631) <= a and b;
    layer2_outputs(6632) <= not (a and b);
    layer2_outputs(6633) <= a;
    layer2_outputs(6634) <= not (a or b);
    layer2_outputs(6635) <= not b;
    layer2_outputs(6636) <= a;
    layer2_outputs(6637) <= not a;
    layer2_outputs(6638) <= b and not a;
    layer2_outputs(6639) <= not b or a;
    layer2_outputs(6640) <= not a;
    layer2_outputs(6641) <= a and not b;
    layer2_outputs(6642) <= a and not b;
    layer2_outputs(6643) <= a;
    layer2_outputs(6644) <= not a or b;
    layer2_outputs(6645) <= not b;
    layer2_outputs(6646) <= not a or b;
    layer2_outputs(6647) <= '0';
    layer2_outputs(6648) <= not a or b;
    layer2_outputs(6649) <= a and not b;
    layer2_outputs(6650) <= a;
    layer2_outputs(6651) <= b;
    layer2_outputs(6652) <= not (a and b);
    layer2_outputs(6653) <= not a or b;
    layer2_outputs(6654) <= not a;
    layer2_outputs(6655) <= b and not a;
    layer2_outputs(6656) <= not (a and b);
    layer2_outputs(6657) <= a or b;
    layer2_outputs(6658) <= not b or a;
    layer2_outputs(6659) <= a or b;
    layer2_outputs(6660) <= not a;
    layer2_outputs(6661) <= not b or a;
    layer2_outputs(6662) <= not b;
    layer2_outputs(6663) <= a and b;
    layer2_outputs(6664) <= a;
    layer2_outputs(6665) <= not b;
    layer2_outputs(6666) <= b;
    layer2_outputs(6667) <= not b or a;
    layer2_outputs(6668) <= b and not a;
    layer2_outputs(6669) <= a and b;
    layer2_outputs(6670) <= b and not a;
    layer2_outputs(6671) <= b and not a;
    layer2_outputs(6672) <= not b or a;
    layer2_outputs(6673) <= '1';
    layer2_outputs(6674) <= not a or b;
    layer2_outputs(6675) <= not (a xor b);
    layer2_outputs(6676) <= not (a and b);
    layer2_outputs(6677) <= not a;
    layer2_outputs(6678) <= a and b;
    layer2_outputs(6679) <= b;
    layer2_outputs(6680) <= b and not a;
    layer2_outputs(6681) <= not b or a;
    layer2_outputs(6682) <= not (a and b);
    layer2_outputs(6683) <= '1';
    layer2_outputs(6684) <= not (a or b);
    layer2_outputs(6685) <= a and b;
    layer2_outputs(6686) <= a or b;
    layer2_outputs(6687) <= b and not a;
    layer2_outputs(6688) <= a xor b;
    layer2_outputs(6689) <= b;
    layer2_outputs(6690) <= not a or b;
    layer2_outputs(6691) <= not a or b;
    layer2_outputs(6692) <= a;
    layer2_outputs(6693) <= not b;
    layer2_outputs(6694) <= a and b;
    layer2_outputs(6695) <= not (a or b);
    layer2_outputs(6696) <= not a or b;
    layer2_outputs(6697) <= a;
    layer2_outputs(6698) <= a or b;
    layer2_outputs(6699) <= not b;
    layer2_outputs(6700) <= not a or b;
    layer2_outputs(6701) <= '1';
    layer2_outputs(6702) <= not (a and b);
    layer2_outputs(6703) <= '0';
    layer2_outputs(6704) <= not (a xor b);
    layer2_outputs(6705) <= not (a or b);
    layer2_outputs(6706) <= a;
    layer2_outputs(6707) <= not a or b;
    layer2_outputs(6708) <= not (a and b);
    layer2_outputs(6709) <= not (a or b);
    layer2_outputs(6710) <= a;
    layer2_outputs(6711) <= not a or b;
    layer2_outputs(6712) <= not b;
    layer2_outputs(6713) <= not a or b;
    layer2_outputs(6714) <= not (a or b);
    layer2_outputs(6715) <= not b;
    layer2_outputs(6716) <= '0';
    layer2_outputs(6717) <= '0';
    layer2_outputs(6718) <= not (a and b);
    layer2_outputs(6719) <= '1';
    layer2_outputs(6720) <= '0';
    layer2_outputs(6721) <= a;
    layer2_outputs(6722) <= b and not a;
    layer2_outputs(6723) <= not (a or b);
    layer2_outputs(6724) <= b;
    layer2_outputs(6725) <= not a;
    layer2_outputs(6726) <= b and not a;
    layer2_outputs(6727) <= a;
    layer2_outputs(6728) <= b;
    layer2_outputs(6729) <= not (a xor b);
    layer2_outputs(6730) <= '0';
    layer2_outputs(6731) <= a and b;
    layer2_outputs(6732) <= '0';
    layer2_outputs(6733) <= a and not b;
    layer2_outputs(6734) <= '1';
    layer2_outputs(6735) <= a and not b;
    layer2_outputs(6736) <= b;
    layer2_outputs(6737) <= a and b;
    layer2_outputs(6738) <= not b or a;
    layer2_outputs(6739) <= '1';
    layer2_outputs(6740) <= a or b;
    layer2_outputs(6741) <= not (a xor b);
    layer2_outputs(6742) <= not a or b;
    layer2_outputs(6743) <= a or b;
    layer2_outputs(6744) <= '0';
    layer2_outputs(6745) <= not a;
    layer2_outputs(6746) <= a;
    layer2_outputs(6747) <= a;
    layer2_outputs(6748) <= a and b;
    layer2_outputs(6749) <= a or b;
    layer2_outputs(6750) <= a;
    layer2_outputs(6751) <= a and not b;
    layer2_outputs(6752) <= a and b;
    layer2_outputs(6753) <= not a or b;
    layer2_outputs(6754) <= not a;
    layer2_outputs(6755) <= a;
    layer2_outputs(6756) <= b;
    layer2_outputs(6757) <= b and not a;
    layer2_outputs(6758) <= a and not b;
    layer2_outputs(6759) <= not (a xor b);
    layer2_outputs(6760) <= not (a or b);
    layer2_outputs(6761) <= a and not b;
    layer2_outputs(6762) <= not (a xor b);
    layer2_outputs(6763) <= '1';
    layer2_outputs(6764) <= not (a xor b);
    layer2_outputs(6765) <= not a;
    layer2_outputs(6766) <= a and b;
    layer2_outputs(6767) <= a and b;
    layer2_outputs(6768) <= not b or a;
    layer2_outputs(6769) <= not b or a;
    layer2_outputs(6770) <= not (a and b);
    layer2_outputs(6771) <= not b or a;
    layer2_outputs(6772) <= a and not b;
    layer2_outputs(6773) <= not (a xor b);
    layer2_outputs(6774) <= not b or a;
    layer2_outputs(6775) <= not a;
    layer2_outputs(6776) <= b;
    layer2_outputs(6777) <= not b or a;
    layer2_outputs(6778) <= not (a xor b);
    layer2_outputs(6779) <= not (a and b);
    layer2_outputs(6780) <= '1';
    layer2_outputs(6781) <= not a;
    layer2_outputs(6782) <= not a;
    layer2_outputs(6783) <= a;
    layer2_outputs(6784) <= not (a or b);
    layer2_outputs(6785) <= not (a xor b);
    layer2_outputs(6786) <= a;
    layer2_outputs(6787) <= a;
    layer2_outputs(6788) <= b and not a;
    layer2_outputs(6789) <= a;
    layer2_outputs(6790) <= not (a and b);
    layer2_outputs(6791) <= a;
    layer2_outputs(6792) <= not (a and b);
    layer2_outputs(6793) <= a and not b;
    layer2_outputs(6794) <= '0';
    layer2_outputs(6795) <= not b or a;
    layer2_outputs(6796) <= a;
    layer2_outputs(6797) <= not b;
    layer2_outputs(6798) <= '0';
    layer2_outputs(6799) <= not (a or b);
    layer2_outputs(6800) <= a and b;
    layer2_outputs(6801) <= b;
    layer2_outputs(6802) <= a;
    layer2_outputs(6803) <= a and b;
    layer2_outputs(6804) <= a or b;
    layer2_outputs(6805) <= not b or a;
    layer2_outputs(6806) <= not b;
    layer2_outputs(6807) <= b and not a;
    layer2_outputs(6808) <= not b or a;
    layer2_outputs(6809) <= not b or a;
    layer2_outputs(6810) <= b;
    layer2_outputs(6811) <= a and not b;
    layer2_outputs(6812) <= not a or b;
    layer2_outputs(6813) <= not (a or b);
    layer2_outputs(6814) <= '0';
    layer2_outputs(6815) <= b and not a;
    layer2_outputs(6816) <= not a;
    layer2_outputs(6817) <= not (a and b);
    layer2_outputs(6818) <= a and b;
    layer2_outputs(6819) <= a;
    layer2_outputs(6820) <= not a;
    layer2_outputs(6821) <= not a;
    layer2_outputs(6822) <= not b or a;
    layer2_outputs(6823) <= not b;
    layer2_outputs(6824) <= not a or b;
    layer2_outputs(6825) <= a and not b;
    layer2_outputs(6826) <= not a;
    layer2_outputs(6827) <= not (a and b);
    layer2_outputs(6828) <= not a or b;
    layer2_outputs(6829) <= not b;
    layer2_outputs(6830) <= a;
    layer2_outputs(6831) <= not (a and b);
    layer2_outputs(6832) <= a or b;
    layer2_outputs(6833) <= not a or b;
    layer2_outputs(6834) <= a and b;
    layer2_outputs(6835) <= not a or b;
    layer2_outputs(6836) <= not b or a;
    layer2_outputs(6837) <= not (a xor b);
    layer2_outputs(6838) <= b and not a;
    layer2_outputs(6839) <= '1';
    layer2_outputs(6840) <= not (a or b);
    layer2_outputs(6841) <= b and not a;
    layer2_outputs(6842) <= b;
    layer2_outputs(6843) <= a and b;
    layer2_outputs(6844) <= not a;
    layer2_outputs(6845) <= not b;
    layer2_outputs(6846) <= not b;
    layer2_outputs(6847) <= not (a or b);
    layer2_outputs(6848) <= not b;
    layer2_outputs(6849) <= not b or a;
    layer2_outputs(6850) <= not b or a;
    layer2_outputs(6851) <= '1';
    layer2_outputs(6852) <= not b;
    layer2_outputs(6853) <= not b;
    layer2_outputs(6854) <= not a;
    layer2_outputs(6855) <= a and not b;
    layer2_outputs(6856) <= '0';
    layer2_outputs(6857) <= not b or a;
    layer2_outputs(6858) <= b and not a;
    layer2_outputs(6859) <= a;
    layer2_outputs(6860) <= '0';
    layer2_outputs(6861) <= not b;
    layer2_outputs(6862) <= a and b;
    layer2_outputs(6863) <= b and not a;
    layer2_outputs(6864) <= not a;
    layer2_outputs(6865) <= '0';
    layer2_outputs(6866) <= not (a xor b);
    layer2_outputs(6867) <= '1';
    layer2_outputs(6868) <= a and b;
    layer2_outputs(6869) <= not a;
    layer2_outputs(6870) <= not (a and b);
    layer2_outputs(6871) <= not a;
    layer2_outputs(6872) <= not b or a;
    layer2_outputs(6873) <= not a;
    layer2_outputs(6874) <= not b;
    layer2_outputs(6875) <= not a or b;
    layer2_outputs(6876) <= not b;
    layer2_outputs(6877) <= '1';
    layer2_outputs(6878) <= not (a or b);
    layer2_outputs(6879) <= a;
    layer2_outputs(6880) <= b;
    layer2_outputs(6881) <= a;
    layer2_outputs(6882) <= not (a or b);
    layer2_outputs(6883) <= not (a or b);
    layer2_outputs(6884) <= b and not a;
    layer2_outputs(6885) <= '0';
    layer2_outputs(6886) <= a;
    layer2_outputs(6887) <= not a;
    layer2_outputs(6888) <= a;
    layer2_outputs(6889) <= a;
    layer2_outputs(6890) <= a and b;
    layer2_outputs(6891) <= not (a and b);
    layer2_outputs(6892) <= b and not a;
    layer2_outputs(6893) <= not a;
    layer2_outputs(6894) <= not a;
    layer2_outputs(6895) <= '0';
    layer2_outputs(6896) <= not a or b;
    layer2_outputs(6897) <= not (a xor b);
    layer2_outputs(6898) <= not (a and b);
    layer2_outputs(6899) <= '0';
    layer2_outputs(6900) <= '0';
    layer2_outputs(6901) <= b;
    layer2_outputs(6902) <= not (a or b);
    layer2_outputs(6903) <= '0';
    layer2_outputs(6904) <= '0';
    layer2_outputs(6905) <= not (a xor b);
    layer2_outputs(6906) <= not b;
    layer2_outputs(6907) <= not a;
    layer2_outputs(6908) <= '1';
    layer2_outputs(6909) <= a or b;
    layer2_outputs(6910) <= a and b;
    layer2_outputs(6911) <= b and not a;
    layer2_outputs(6912) <= '0';
    layer2_outputs(6913) <= b;
    layer2_outputs(6914) <= a or b;
    layer2_outputs(6915) <= '0';
    layer2_outputs(6916) <= not a or b;
    layer2_outputs(6917) <= a or b;
    layer2_outputs(6918) <= not (a and b);
    layer2_outputs(6919) <= a or b;
    layer2_outputs(6920) <= a;
    layer2_outputs(6921) <= a and not b;
    layer2_outputs(6922) <= not a or b;
    layer2_outputs(6923) <= a and b;
    layer2_outputs(6924) <= a and b;
    layer2_outputs(6925) <= not a or b;
    layer2_outputs(6926) <= not a;
    layer2_outputs(6927) <= not (a and b);
    layer2_outputs(6928) <= a;
    layer2_outputs(6929) <= not (a and b);
    layer2_outputs(6930) <= not b or a;
    layer2_outputs(6931) <= not b or a;
    layer2_outputs(6932) <= not a;
    layer2_outputs(6933) <= not (a or b);
    layer2_outputs(6934) <= b;
    layer2_outputs(6935) <= a or b;
    layer2_outputs(6936) <= a;
    layer2_outputs(6937) <= not b;
    layer2_outputs(6938) <= a;
    layer2_outputs(6939) <= not (a and b);
    layer2_outputs(6940) <= not a;
    layer2_outputs(6941) <= b and not a;
    layer2_outputs(6942) <= a or b;
    layer2_outputs(6943) <= a;
    layer2_outputs(6944) <= not b or a;
    layer2_outputs(6945) <= not b or a;
    layer2_outputs(6946) <= not (a or b);
    layer2_outputs(6947) <= '1';
    layer2_outputs(6948) <= b;
    layer2_outputs(6949) <= not b;
    layer2_outputs(6950) <= not b;
    layer2_outputs(6951) <= a;
    layer2_outputs(6952) <= not a or b;
    layer2_outputs(6953) <= not a;
    layer2_outputs(6954) <= a and not b;
    layer2_outputs(6955) <= not b or a;
    layer2_outputs(6956) <= a and not b;
    layer2_outputs(6957) <= not a or b;
    layer2_outputs(6958) <= '0';
    layer2_outputs(6959) <= a or b;
    layer2_outputs(6960) <= a or b;
    layer2_outputs(6961) <= '0';
    layer2_outputs(6962) <= not (a or b);
    layer2_outputs(6963) <= not a or b;
    layer2_outputs(6964) <= a and not b;
    layer2_outputs(6965) <= '0';
    layer2_outputs(6966) <= '0';
    layer2_outputs(6967) <= '0';
    layer2_outputs(6968) <= '1';
    layer2_outputs(6969) <= a;
    layer2_outputs(6970) <= '1';
    layer2_outputs(6971) <= a and b;
    layer2_outputs(6972) <= a and b;
    layer2_outputs(6973) <= a;
    layer2_outputs(6974) <= not b or a;
    layer2_outputs(6975) <= not (a or b);
    layer2_outputs(6976) <= '1';
    layer2_outputs(6977) <= '0';
    layer2_outputs(6978) <= b;
    layer2_outputs(6979) <= not b;
    layer2_outputs(6980) <= '1';
    layer2_outputs(6981) <= not (a and b);
    layer2_outputs(6982) <= a;
    layer2_outputs(6983) <= not a;
    layer2_outputs(6984) <= '1';
    layer2_outputs(6985) <= a and b;
    layer2_outputs(6986) <= not a;
    layer2_outputs(6987) <= a and not b;
    layer2_outputs(6988) <= not (a or b);
    layer2_outputs(6989) <= a and not b;
    layer2_outputs(6990) <= not a;
    layer2_outputs(6991) <= '1';
    layer2_outputs(6992) <= '0';
    layer2_outputs(6993) <= b;
    layer2_outputs(6994) <= not (a xor b);
    layer2_outputs(6995) <= not b or a;
    layer2_outputs(6996) <= not b;
    layer2_outputs(6997) <= '0';
    layer2_outputs(6998) <= '0';
    layer2_outputs(6999) <= b;
    layer2_outputs(7000) <= not b;
    layer2_outputs(7001) <= b;
    layer2_outputs(7002) <= not b;
    layer2_outputs(7003) <= a or b;
    layer2_outputs(7004) <= not (a and b);
    layer2_outputs(7005) <= not b;
    layer2_outputs(7006) <= not a;
    layer2_outputs(7007) <= a;
    layer2_outputs(7008) <= a or b;
    layer2_outputs(7009) <= a and not b;
    layer2_outputs(7010) <= not (a or b);
    layer2_outputs(7011) <= '0';
    layer2_outputs(7012) <= not a;
    layer2_outputs(7013) <= '1';
    layer2_outputs(7014) <= a;
    layer2_outputs(7015) <= '0';
    layer2_outputs(7016) <= not a or b;
    layer2_outputs(7017) <= a;
    layer2_outputs(7018) <= a or b;
    layer2_outputs(7019) <= a xor b;
    layer2_outputs(7020) <= a or b;
    layer2_outputs(7021) <= b and not a;
    layer2_outputs(7022) <= not (a xor b);
    layer2_outputs(7023) <= not a;
    layer2_outputs(7024) <= b;
    layer2_outputs(7025) <= '0';
    layer2_outputs(7026) <= not b;
    layer2_outputs(7027) <= a;
    layer2_outputs(7028) <= not (a xor b);
    layer2_outputs(7029) <= a;
    layer2_outputs(7030) <= not (a or b);
    layer2_outputs(7031) <= a or b;
    layer2_outputs(7032) <= '0';
    layer2_outputs(7033) <= not (a and b);
    layer2_outputs(7034) <= not (a or b);
    layer2_outputs(7035) <= a and b;
    layer2_outputs(7036) <= not b or a;
    layer2_outputs(7037) <= a or b;
    layer2_outputs(7038) <= a and b;
    layer2_outputs(7039) <= b;
    layer2_outputs(7040) <= not (a or b);
    layer2_outputs(7041) <= not (a and b);
    layer2_outputs(7042) <= a;
    layer2_outputs(7043) <= b and not a;
    layer2_outputs(7044) <= not a or b;
    layer2_outputs(7045) <= a;
    layer2_outputs(7046) <= b;
    layer2_outputs(7047) <= b and not a;
    layer2_outputs(7048) <= b;
    layer2_outputs(7049) <= not b or a;
    layer2_outputs(7050) <= not a or b;
    layer2_outputs(7051) <= not b;
    layer2_outputs(7052) <= not (a xor b);
    layer2_outputs(7053) <= '0';
    layer2_outputs(7054) <= not a;
    layer2_outputs(7055) <= not a or b;
    layer2_outputs(7056) <= a or b;
    layer2_outputs(7057) <= not (a and b);
    layer2_outputs(7058) <= a or b;
    layer2_outputs(7059) <= '0';
    layer2_outputs(7060) <= not (a or b);
    layer2_outputs(7061) <= a or b;
    layer2_outputs(7062) <= a xor b;
    layer2_outputs(7063) <= a xor b;
    layer2_outputs(7064) <= not (a or b);
    layer2_outputs(7065) <= a;
    layer2_outputs(7066) <= a;
    layer2_outputs(7067) <= not a or b;
    layer2_outputs(7068) <= b;
    layer2_outputs(7069) <= not (a or b);
    layer2_outputs(7070) <= a and b;
    layer2_outputs(7071) <= a or b;
    layer2_outputs(7072) <= b;
    layer2_outputs(7073) <= b and not a;
    layer2_outputs(7074) <= b and not a;
    layer2_outputs(7075) <= not (a or b);
    layer2_outputs(7076) <= not (a and b);
    layer2_outputs(7077) <= not a;
    layer2_outputs(7078) <= a and not b;
    layer2_outputs(7079) <= not a;
    layer2_outputs(7080) <= '0';
    layer2_outputs(7081) <= a and not b;
    layer2_outputs(7082) <= b and not a;
    layer2_outputs(7083) <= a or b;
    layer2_outputs(7084) <= a and not b;
    layer2_outputs(7085) <= not b;
    layer2_outputs(7086) <= not b;
    layer2_outputs(7087) <= a and not b;
    layer2_outputs(7088) <= a xor b;
    layer2_outputs(7089) <= not a or b;
    layer2_outputs(7090) <= a;
    layer2_outputs(7091) <= not b or a;
    layer2_outputs(7092) <= not b;
    layer2_outputs(7093) <= a;
    layer2_outputs(7094) <= b;
    layer2_outputs(7095) <= a;
    layer2_outputs(7096) <= '1';
    layer2_outputs(7097) <= a or b;
    layer2_outputs(7098) <= not b or a;
    layer2_outputs(7099) <= not a;
    layer2_outputs(7100) <= a and b;
    layer2_outputs(7101) <= a and b;
    layer2_outputs(7102) <= b and not a;
    layer2_outputs(7103) <= not (a or b);
    layer2_outputs(7104) <= not b;
    layer2_outputs(7105) <= not a;
    layer2_outputs(7106) <= not a;
    layer2_outputs(7107) <= not b;
    layer2_outputs(7108) <= a and not b;
    layer2_outputs(7109) <= not a;
    layer2_outputs(7110) <= '0';
    layer2_outputs(7111) <= not (a and b);
    layer2_outputs(7112) <= a;
    layer2_outputs(7113) <= a and b;
    layer2_outputs(7114) <= not (a and b);
    layer2_outputs(7115) <= a or b;
    layer2_outputs(7116) <= not a or b;
    layer2_outputs(7117) <= not b or a;
    layer2_outputs(7118) <= not (a xor b);
    layer2_outputs(7119) <= not (a and b);
    layer2_outputs(7120) <= not b;
    layer2_outputs(7121) <= not b or a;
    layer2_outputs(7122) <= not (a xor b);
    layer2_outputs(7123) <= a;
    layer2_outputs(7124) <= not a;
    layer2_outputs(7125) <= not (a xor b);
    layer2_outputs(7126) <= not a;
    layer2_outputs(7127) <= not b or a;
    layer2_outputs(7128) <= '1';
    layer2_outputs(7129) <= b;
    layer2_outputs(7130) <= not a;
    layer2_outputs(7131) <= '0';
    layer2_outputs(7132) <= not (a and b);
    layer2_outputs(7133) <= a xor b;
    layer2_outputs(7134) <= not (a or b);
    layer2_outputs(7135) <= '1';
    layer2_outputs(7136) <= b and not a;
    layer2_outputs(7137) <= b and not a;
    layer2_outputs(7138) <= not b or a;
    layer2_outputs(7139) <= b and not a;
    layer2_outputs(7140) <= not b or a;
    layer2_outputs(7141) <= a xor b;
    layer2_outputs(7142) <= not b or a;
    layer2_outputs(7143) <= not (a and b);
    layer2_outputs(7144) <= not (a or b);
    layer2_outputs(7145) <= b and not a;
    layer2_outputs(7146) <= not a;
    layer2_outputs(7147) <= b;
    layer2_outputs(7148) <= a and not b;
    layer2_outputs(7149) <= a or b;
    layer2_outputs(7150) <= not a or b;
    layer2_outputs(7151) <= not a or b;
    layer2_outputs(7152) <= not b or a;
    layer2_outputs(7153) <= a;
    layer2_outputs(7154) <= not (a xor b);
    layer2_outputs(7155) <= '1';
    layer2_outputs(7156) <= b and not a;
    layer2_outputs(7157) <= not a;
    layer2_outputs(7158) <= b and not a;
    layer2_outputs(7159) <= not b or a;
    layer2_outputs(7160) <= a;
    layer2_outputs(7161) <= a;
    layer2_outputs(7162) <= '1';
    layer2_outputs(7163) <= a or b;
    layer2_outputs(7164) <= a;
    layer2_outputs(7165) <= not a;
    layer2_outputs(7166) <= not b;
    layer2_outputs(7167) <= b;
    layer2_outputs(7168) <= not b or a;
    layer2_outputs(7169) <= a and not b;
    layer2_outputs(7170) <= not (a or b);
    layer2_outputs(7171) <= b and not a;
    layer2_outputs(7172) <= a;
    layer2_outputs(7173) <= not (a or b);
    layer2_outputs(7174) <= '0';
    layer2_outputs(7175) <= not (a and b);
    layer2_outputs(7176) <= not a or b;
    layer2_outputs(7177) <= not (a or b);
    layer2_outputs(7178) <= not (a and b);
    layer2_outputs(7179) <= b and not a;
    layer2_outputs(7180) <= a;
    layer2_outputs(7181) <= not (a or b);
    layer2_outputs(7182) <= a and b;
    layer2_outputs(7183) <= a;
    layer2_outputs(7184) <= a and not b;
    layer2_outputs(7185) <= b;
    layer2_outputs(7186) <= not a;
    layer2_outputs(7187) <= not b;
    layer2_outputs(7188) <= a or b;
    layer2_outputs(7189) <= a and not b;
    layer2_outputs(7190) <= a and not b;
    layer2_outputs(7191) <= a;
    layer2_outputs(7192) <= not a;
    layer2_outputs(7193) <= not b;
    layer2_outputs(7194) <= not (a and b);
    layer2_outputs(7195) <= b and not a;
    layer2_outputs(7196) <= a or b;
    layer2_outputs(7197) <= '0';
    layer2_outputs(7198) <= b;
    layer2_outputs(7199) <= not (a and b);
    layer2_outputs(7200) <= not (a or b);
    layer2_outputs(7201) <= b;
    layer2_outputs(7202) <= a and not b;
    layer2_outputs(7203) <= not a or b;
    layer2_outputs(7204) <= a and b;
    layer2_outputs(7205) <= b;
    layer2_outputs(7206) <= a;
    layer2_outputs(7207) <= b;
    layer2_outputs(7208) <= not a or b;
    layer2_outputs(7209) <= not b;
    layer2_outputs(7210) <= a xor b;
    layer2_outputs(7211) <= a and not b;
    layer2_outputs(7212) <= a and b;
    layer2_outputs(7213) <= a or b;
    layer2_outputs(7214) <= '1';
    layer2_outputs(7215) <= a xor b;
    layer2_outputs(7216) <= not (a or b);
    layer2_outputs(7217) <= b and not a;
    layer2_outputs(7218) <= a or b;
    layer2_outputs(7219) <= a;
    layer2_outputs(7220) <= not (a and b);
    layer2_outputs(7221) <= not (a and b);
    layer2_outputs(7222) <= b;
    layer2_outputs(7223) <= a;
    layer2_outputs(7224) <= not a;
    layer2_outputs(7225) <= a and not b;
    layer2_outputs(7226) <= b;
    layer2_outputs(7227) <= '1';
    layer2_outputs(7228) <= b;
    layer2_outputs(7229) <= not b or a;
    layer2_outputs(7230) <= a or b;
    layer2_outputs(7231) <= not b;
    layer2_outputs(7232) <= '1';
    layer2_outputs(7233) <= not (a or b);
    layer2_outputs(7234) <= a and b;
    layer2_outputs(7235) <= not a;
    layer2_outputs(7236) <= not a;
    layer2_outputs(7237) <= not (a xor b);
    layer2_outputs(7238) <= a;
    layer2_outputs(7239) <= b;
    layer2_outputs(7240) <= not b;
    layer2_outputs(7241) <= '0';
    layer2_outputs(7242) <= not a or b;
    layer2_outputs(7243) <= b;
    layer2_outputs(7244) <= a or b;
    layer2_outputs(7245) <= not b;
    layer2_outputs(7246) <= b and not a;
    layer2_outputs(7247) <= a or b;
    layer2_outputs(7248) <= not a or b;
    layer2_outputs(7249) <= not b;
    layer2_outputs(7250) <= a or b;
    layer2_outputs(7251) <= not (a xor b);
    layer2_outputs(7252) <= a;
    layer2_outputs(7253) <= not (a and b);
    layer2_outputs(7254) <= not (a xor b);
    layer2_outputs(7255) <= not a;
    layer2_outputs(7256) <= a and b;
    layer2_outputs(7257) <= '1';
    layer2_outputs(7258) <= a and not b;
    layer2_outputs(7259) <= a or b;
    layer2_outputs(7260) <= not a or b;
    layer2_outputs(7261) <= '1';
    layer2_outputs(7262) <= b;
    layer2_outputs(7263) <= not (a xor b);
    layer2_outputs(7264) <= not a or b;
    layer2_outputs(7265) <= not a or b;
    layer2_outputs(7266) <= a and b;
    layer2_outputs(7267) <= not b;
    layer2_outputs(7268) <= '1';
    layer2_outputs(7269) <= b and not a;
    layer2_outputs(7270) <= not (a and b);
    layer2_outputs(7271) <= b;
    layer2_outputs(7272) <= '0';
    layer2_outputs(7273) <= a or b;
    layer2_outputs(7274) <= not a;
    layer2_outputs(7275) <= not (a and b);
    layer2_outputs(7276) <= not a or b;
    layer2_outputs(7277) <= not a or b;
    layer2_outputs(7278) <= not (a and b);
    layer2_outputs(7279) <= not (a xor b);
    layer2_outputs(7280) <= not b;
    layer2_outputs(7281) <= not (a xor b);
    layer2_outputs(7282) <= b and not a;
    layer2_outputs(7283) <= not b or a;
    layer2_outputs(7284) <= a;
    layer2_outputs(7285) <= not a;
    layer2_outputs(7286) <= a;
    layer2_outputs(7287) <= not b;
    layer2_outputs(7288) <= not b or a;
    layer2_outputs(7289) <= a;
    layer2_outputs(7290) <= a;
    layer2_outputs(7291) <= not (a or b);
    layer2_outputs(7292) <= b;
    layer2_outputs(7293) <= a;
    layer2_outputs(7294) <= not a;
    layer2_outputs(7295) <= not b;
    layer2_outputs(7296) <= not (a xor b);
    layer2_outputs(7297) <= b;
    layer2_outputs(7298) <= not (a xor b);
    layer2_outputs(7299) <= not (a xor b);
    layer2_outputs(7300) <= not a;
    layer2_outputs(7301) <= not (a and b);
    layer2_outputs(7302) <= b and not a;
    layer2_outputs(7303) <= not a;
    layer2_outputs(7304) <= b;
    layer2_outputs(7305) <= not a;
    layer2_outputs(7306) <= not b;
    layer2_outputs(7307) <= not a;
    layer2_outputs(7308) <= not b;
    layer2_outputs(7309) <= b;
    layer2_outputs(7310) <= not b;
    layer2_outputs(7311) <= '1';
    layer2_outputs(7312) <= '0';
    layer2_outputs(7313) <= '0';
    layer2_outputs(7314) <= a xor b;
    layer2_outputs(7315) <= not b;
    layer2_outputs(7316) <= b;
    layer2_outputs(7317) <= not b;
    layer2_outputs(7318) <= a and b;
    layer2_outputs(7319) <= a and b;
    layer2_outputs(7320) <= not (a and b);
    layer2_outputs(7321) <= not b;
    layer2_outputs(7322) <= not (a and b);
    layer2_outputs(7323) <= not a;
    layer2_outputs(7324) <= not a or b;
    layer2_outputs(7325) <= not a;
    layer2_outputs(7326) <= not (a and b);
    layer2_outputs(7327) <= '0';
    layer2_outputs(7328) <= a or b;
    layer2_outputs(7329) <= a or b;
    layer2_outputs(7330) <= not (a and b);
    layer2_outputs(7331) <= a and b;
    layer2_outputs(7332) <= a;
    layer2_outputs(7333) <= not (a xor b);
    layer2_outputs(7334) <= not b or a;
    layer2_outputs(7335) <= not a or b;
    layer2_outputs(7336) <= a and not b;
    layer2_outputs(7337) <= a or b;
    layer2_outputs(7338) <= '0';
    layer2_outputs(7339) <= a and not b;
    layer2_outputs(7340) <= not b;
    layer2_outputs(7341) <= '0';
    layer2_outputs(7342) <= a;
    layer2_outputs(7343) <= not a or b;
    layer2_outputs(7344) <= a;
    layer2_outputs(7345) <= '0';
    layer2_outputs(7346) <= not a;
    layer2_outputs(7347) <= not b or a;
    layer2_outputs(7348) <= not b;
    layer2_outputs(7349) <= b;
    layer2_outputs(7350) <= b and not a;
    layer2_outputs(7351) <= a and b;
    layer2_outputs(7352) <= '0';
    layer2_outputs(7353) <= a;
    layer2_outputs(7354) <= not a or b;
    layer2_outputs(7355) <= b and not a;
    layer2_outputs(7356) <= not a;
    layer2_outputs(7357) <= a and b;
    layer2_outputs(7358) <= a;
    layer2_outputs(7359) <= not (a or b);
    layer2_outputs(7360) <= a and b;
    layer2_outputs(7361) <= not b;
    layer2_outputs(7362) <= not (a xor b);
    layer2_outputs(7363) <= a;
    layer2_outputs(7364) <= '1';
    layer2_outputs(7365) <= not b or a;
    layer2_outputs(7366) <= a;
    layer2_outputs(7367) <= not (a and b);
    layer2_outputs(7368) <= not (a and b);
    layer2_outputs(7369) <= not b or a;
    layer2_outputs(7370) <= a and b;
    layer2_outputs(7371) <= a or b;
    layer2_outputs(7372) <= '0';
    layer2_outputs(7373) <= not (a and b);
    layer2_outputs(7374) <= not b or a;
    layer2_outputs(7375) <= not (a and b);
    layer2_outputs(7376) <= b;
    layer2_outputs(7377) <= a or b;
    layer2_outputs(7378) <= not b;
    layer2_outputs(7379) <= not a or b;
    layer2_outputs(7380) <= not (a or b);
    layer2_outputs(7381) <= not (a and b);
    layer2_outputs(7382) <= a;
    layer2_outputs(7383) <= b and not a;
    layer2_outputs(7384) <= not a;
    layer2_outputs(7385) <= not b;
    layer2_outputs(7386) <= not (a and b);
    layer2_outputs(7387) <= not b;
    layer2_outputs(7388) <= a;
    layer2_outputs(7389) <= not (a xor b);
    layer2_outputs(7390) <= not a;
    layer2_outputs(7391) <= not (a and b);
    layer2_outputs(7392) <= not (a and b);
    layer2_outputs(7393) <= a and b;
    layer2_outputs(7394) <= not (a xor b);
    layer2_outputs(7395) <= a and not b;
    layer2_outputs(7396) <= '0';
    layer2_outputs(7397) <= a;
    layer2_outputs(7398) <= '0';
    layer2_outputs(7399) <= not b or a;
    layer2_outputs(7400) <= not a;
    layer2_outputs(7401) <= not b;
    layer2_outputs(7402) <= a and not b;
    layer2_outputs(7403) <= not b;
    layer2_outputs(7404) <= a and b;
    layer2_outputs(7405) <= b;
    layer2_outputs(7406) <= not a;
    layer2_outputs(7407) <= '1';
    layer2_outputs(7408) <= not a;
    layer2_outputs(7409) <= a;
    layer2_outputs(7410) <= a or b;
    layer2_outputs(7411) <= a;
    layer2_outputs(7412) <= b and not a;
    layer2_outputs(7413) <= not (a or b);
    layer2_outputs(7414) <= a;
    layer2_outputs(7415) <= a or b;
    layer2_outputs(7416) <= a and b;
    layer2_outputs(7417) <= a or b;
    layer2_outputs(7418) <= '1';
    layer2_outputs(7419) <= not a;
    layer2_outputs(7420) <= not (a and b);
    layer2_outputs(7421) <= '1';
    layer2_outputs(7422) <= not b;
    layer2_outputs(7423) <= b;
    layer2_outputs(7424) <= not a;
    layer2_outputs(7425) <= a and b;
    layer2_outputs(7426) <= a;
    layer2_outputs(7427) <= not (a and b);
    layer2_outputs(7428) <= b and not a;
    layer2_outputs(7429) <= a or b;
    layer2_outputs(7430) <= a and not b;
    layer2_outputs(7431) <= not (a or b);
    layer2_outputs(7432) <= a xor b;
    layer2_outputs(7433) <= not a;
    layer2_outputs(7434) <= not b or a;
    layer2_outputs(7435) <= not (a and b);
    layer2_outputs(7436) <= b;
    layer2_outputs(7437) <= b and not a;
    layer2_outputs(7438) <= not a or b;
    layer2_outputs(7439) <= b and not a;
    layer2_outputs(7440) <= not b;
    layer2_outputs(7441) <= not (a or b);
    layer2_outputs(7442) <= a or b;
    layer2_outputs(7443) <= b;
    layer2_outputs(7444) <= b and not a;
    layer2_outputs(7445) <= not b or a;
    layer2_outputs(7446) <= b;
    layer2_outputs(7447) <= a and b;
    layer2_outputs(7448) <= b and not a;
    layer2_outputs(7449) <= not a;
    layer2_outputs(7450) <= a and not b;
    layer2_outputs(7451) <= not (a xor b);
    layer2_outputs(7452) <= b and not a;
    layer2_outputs(7453) <= b and not a;
    layer2_outputs(7454) <= not b or a;
    layer2_outputs(7455) <= '1';
    layer2_outputs(7456) <= b and not a;
    layer2_outputs(7457) <= not b;
    layer2_outputs(7458) <= b;
    layer2_outputs(7459) <= a;
    layer2_outputs(7460) <= b and not a;
    layer2_outputs(7461) <= a and b;
    layer2_outputs(7462) <= not b;
    layer2_outputs(7463) <= a;
    layer2_outputs(7464) <= a or b;
    layer2_outputs(7465) <= b and not a;
    layer2_outputs(7466) <= a or b;
    layer2_outputs(7467) <= a and not b;
    layer2_outputs(7468) <= not (a and b);
    layer2_outputs(7469) <= b;
    layer2_outputs(7470) <= a;
    layer2_outputs(7471) <= a or b;
    layer2_outputs(7472) <= a and b;
    layer2_outputs(7473) <= b;
    layer2_outputs(7474) <= not b;
    layer2_outputs(7475) <= a;
    layer2_outputs(7476) <= not b or a;
    layer2_outputs(7477) <= a xor b;
    layer2_outputs(7478) <= a;
    layer2_outputs(7479) <= a and not b;
    layer2_outputs(7480) <= not a;
    layer2_outputs(7481) <= not (a xor b);
    layer2_outputs(7482) <= a and b;
    layer2_outputs(7483) <= not b;
    layer2_outputs(7484) <= not (a and b);
    layer2_outputs(7485) <= not a;
    layer2_outputs(7486) <= a or b;
    layer2_outputs(7487) <= not a or b;
    layer2_outputs(7488) <= a and b;
    layer2_outputs(7489) <= not a or b;
    layer2_outputs(7490) <= b and not a;
    layer2_outputs(7491) <= a and not b;
    layer2_outputs(7492) <= not (a and b);
    layer2_outputs(7493) <= '0';
    layer2_outputs(7494) <= a and not b;
    layer2_outputs(7495) <= not (a or b);
    layer2_outputs(7496) <= not a or b;
    layer2_outputs(7497) <= not (a and b);
    layer2_outputs(7498) <= not (a and b);
    layer2_outputs(7499) <= a and not b;
    layer2_outputs(7500) <= not a;
    layer2_outputs(7501) <= not a;
    layer2_outputs(7502) <= '0';
    layer2_outputs(7503) <= a and b;
    layer2_outputs(7504) <= not a;
    layer2_outputs(7505) <= b and not a;
    layer2_outputs(7506) <= '1';
    layer2_outputs(7507) <= a and b;
    layer2_outputs(7508) <= a and b;
    layer2_outputs(7509) <= not (a or b);
    layer2_outputs(7510) <= b;
    layer2_outputs(7511) <= not b or a;
    layer2_outputs(7512) <= not a;
    layer2_outputs(7513) <= a and not b;
    layer2_outputs(7514) <= not a;
    layer2_outputs(7515) <= not a;
    layer2_outputs(7516) <= not (a or b);
    layer2_outputs(7517) <= '1';
    layer2_outputs(7518) <= a and not b;
    layer2_outputs(7519) <= a and not b;
    layer2_outputs(7520) <= not b;
    layer2_outputs(7521) <= a or b;
    layer2_outputs(7522) <= not b or a;
    layer2_outputs(7523) <= a and not b;
    layer2_outputs(7524) <= '1';
    layer2_outputs(7525) <= a;
    layer2_outputs(7526) <= not b;
    layer2_outputs(7527) <= not b;
    layer2_outputs(7528) <= a;
    layer2_outputs(7529) <= not (a and b);
    layer2_outputs(7530) <= a or b;
    layer2_outputs(7531) <= not (a or b);
    layer2_outputs(7532) <= a and b;
    layer2_outputs(7533) <= not (a or b);
    layer2_outputs(7534) <= not b;
    layer2_outputs(7535) <= not (a and b);
    layer2_outputs(7536) <= not (a or b);
    layer2_outputs(7537) <= b and not a;
    layer2_outputs(7538) <= not a or b;
    layer2_outputs(7539) <= a;
    layer2_outputs(7540) <= '0';
    layer2_outputs(7541) <= a and not b;
    layer2_outputs(7542) <= not b;
    layer2_outputs(7543) <= a and b;
    layer2_outputs(7544) <= '0';
    layer2_outputs(7545) <= b;
    layer2_outputs(7546) <= not a or b;
    layer2_outputs(7547) <= not (a or b);
    layer2_outputs(7548) <= a;
    layer2_outputs(7549) <= a;
    layer2_outputs(7550) <= b;
    layer2_outputs(7551) <= '1';
    layer2_outputs(7552) <= not b or a;
    layer2_outputs(7553) <= '0';
    layer2_outputs(7554) <= not b or a;
    layer2_outputs(7555) <= not b;
    layer2_outputs(7556) <= not a or b;
    layer2_outputs(7557) <= not a;
    layer2_outputs(7558) <= b;
    layer2_outputs(7559) <= a and not b;
    layer2_outputs(7560) <= b and not a;
    layer2_outputs(7561) <= a or b;
    layer2_outputs(7562) <= a and not b;
    layer2_outputs(7563) <= b and not a;
    layer2_outputs(7564) <= '1';
    layer2_outputs(7565) <= b;
    layer2_outputs(7566) <= not (a or b);
    layer2_outputs(7567) <= '0';
    layer2_outputs(7568) <= not a;
    layer2_outputs(7569) <= not a;
    layer2_outputs(7570) <= not a;
    layer2_outputs(7571) <= not a;
    layer2_outputs(7572) <= a;
    layer2_outputs(7573) <= not b;
    layer2_outputs(7574) <= not (a or b);
    layer2_outputs(7575) <= not a or b;
    layer2_outputs(7576) <= a or b;
    layer2_outputs(7577) <= a or b;
    layer2_outputs(7578) <= a or b;
    layer2_outputs(7579) <= not b;
    layer2_outputs(7580) <= not b;
    layer2_outputs(7581) <= a and b;
    layer2_outputs(7582) <= b;
    layer2_outputs(7583) <= a;
    layer2_outputs(7584) <= not (a or b);
    layer2_outputs(7585) <= b;
    layer2_outputs(7586) <= not b or a;
    layer2_outputs(7587) <= not (a or b);
    layer2_outputs(7588) <= b and not a;
    layer2_outputs(7589) <= not a;
    layer2_outputs(7590) <= not a or b;
    layer2_outputs(7591) <= '0';
    layer2_outputs(7592) <= not (a and b);
    layer2_outputs(7593) <= '0';
    layer2_outputs(7594) <= not (a or b);
    layer2_outputs(7595) <= not (a and b);
    layer2_outputs(7596) <= a;
    layer2_outputs(7597) <= a and not b;
    layer2_outputs(7598) <= a and b;
    layer2_outputs(7599) <= not b or a;
    layer2_outputs(7600) <= not a;
    layer2_outputs(7601) <= not b;
    layer2_outputs(7602) <= not b;
    layer2_outputs(7603) <= '1';
    layer2_outputs(7604) <= b;
    layer2_outputs(7605) <= not a;
    layer2_outputs(7606) <= a or b;
    layer2_outputs(7607) <= not a;
    layer2_outputs(7608) <= not (a and b);
    layer2_outputs(7609) <= a or b;
    layer2_outputs(7610) <= not a;
    layer2_outputs(7611) <= not b;
    layer2_outputs(7612) <= a and b;
    layer2_outputs(7613) <= not b;
    layer2_outputs(7614) <= b;
    layer2_outputs(7615) <= a and not b;
    layer2_outputs(7616) <= not b;
    layer2_outputs(7617) <= not (a or b);
    layer2_outputs(7618) <= a;
    layer2_outputs(7619) <= b;
    layer2_outputs(7620) <= b;
    layer2_outputs(7621) <= b;
    layer2_outputs(7622) <= b;
    layer2_outputs(7623) <= not b;
    layer2_outputs(7624) <= not (a and b);
    layer2_outputs(7625) <= not (a and b);
    layer2_outputs(7626) <= not (a or b);
    layer2_outputs(7627) <= '0';
    layer2_outputs(7628) <= not a;
    layer2_outputs(7629) <= a and not b;
    layer2_outputs(7630) <= not b or a;
    layer2_outputs(7631) <= b;
    layer2_outputs(7632) <= not b;
    layer2_outputs(7633) <= a or b;
    layer2_outputs(7634) <= not (a xor b);
    layer2_outputs(7635) <= a and b;
    layer2_outputs(7636) <= not (a and b);
    layer2_outputs(7637) <= a and not b;
    layer2_outputs(7638) <= a and b;
    layer2_outputs(7639) <= not b;
    layer2_outputs(7640) <= not a;
    layer2_outputs(7641) <= not (a and b);
    layer2_outputs(7642) <= not b or a;
    layer2_outputs(7643) <= b;
    layer2_outputs(7644) <= not a;
    layer2_outputs(7645) <= not b;
    layer2_outputs(7646) <= not b or a;
    layer2_outputs(7647) <= not b or a;
    layer2_outputs(7648) <= not a or b;
    layer2_outputs(7649) <= a;
    layer2_outputs(7650) <= a or b;
    layer2_outputs(7651) <= not (a or b);
    layer2_outputs(7652) <= not b or a;
    layer2_outputs(7653) <= a and b;
    layer2_outputs(7654) <= '1';
    layer2_outputs(7655) <= b;
    layer2_outputs(7656) <= b;
    layer2_outputs(7657) <= b;
    layer2_outputs(7658) <= a xor b;
    layer2_outputs(7659) <= not (a or b);
    layer2_outputs(7660) <= not (a and b);
    layer2_outputs(7661) <= not (a or b);
    layer2_outputs(7662) <= not (a and b);
    layer2_outputs(7663) <= not (a and b);
    layer2_outputs(7664) <= b;
    layer2_outputs(7665) <= b;
    layer2_outputs(7666) <= not a;
    layer2_outputs(7667) <= b and not a;
    layer2_outputs(7668) <= a and b;
    layer2_outputs(7669) <= not b;
    layer2_outputs(7670) <= not b;
    layer2_outputs(7671) <= a;
    layer2_outputs(7672) <= not (a xor b);
    layer2_outputs(7673) <= a and b;
    layer2_outputs(7674) <= not (a and b);
    layer2_outputs(7675) <= not b;
    layer2_outputs(7676) <= b;
    layer2_outputs(7677) <= not (a and b);
    layer2_outputs(7678) <= not (a or b);
    layer2_outputs(7679) <= not a or b;
    layer2_outputs(7680) <= not b;
    layer2_outputs(7681) <= b;
    layer2_outputs(7682) <= not a;
    layer2_outputs(7683) <= a and b;
    layer2_outputs(7684) <= a xor b;
    layer2_outputs(7685) <= a xor b;
    layer2_outputs(7686) <= a;
    layer2_outputs(7687) <= not b;
    layer2_outputs(7688) <= not (a and b);
    layer2_outputs(7689) <= not b;
    layer2_outputs(7690) <= a or b;
    layer2_outputs(7691) <= a;
    layer2_outputs(7692) <= '1';
    layer2_outputs(7693) <= not (a or b);
    layer2_outputs(7694) <= b and not a;
    layer2_outputs(7695) <= not b or a;
    layer2_outputs(7696) <= not a;
    layer2_outputs(7697) <= not b or a;
    layer2_outputs(7698) <= a or b;
    layer2_outputs(7699) <= a;
    layer2_outputs(7700) <= a or b;
    layer2_outputs(7701) <= b and not a;
    layer2_outputs(7702) <= a and not b;
    layer2_outputs(7703) <= '0';
    layer2_outputs(7704) <= not a;
    layer2_outputs(7705) <= not (a or b);
    layer2_outputs(7706) <= a;
    layer2_outputs(7707) <= not a;
    layer2_outputs(7708) <= a and not b;
    layer2_outputs(7709) <= '1';
    layer2_outputs(7710) <= '0';
    layer2_outputs(7711) <= not b or a;
    layer2_outputs(7712) <= '1';
    layer2_outputs(7713) <= not a or b;
    layer2_outputs(7714) <= '1';
    layer2_outputs(7715) <= not (a and b);
    layer2_outputs(7716) <= a or b;
    layer2_outputs(7717) <= not b;
    layer2_outputs(7718) <= a xor b;
    layer2_outputs(7719) <= '1';
    layer2_outputs(7720) <= not b or a;
    layer2_outputs(7721) <= a;
    layer2_outputs(7722) <= not b or a;
    layer2_outputs(7723) <= not a;
    layer2_outputs(7724) <= a or b;
    layer2_outputs(7725) <= not (a or b);
    layer2_outputs(7726) <= a and not b;
    layer2_outputs(7727) <= b and not a;
    layer2_outputs(7728) <= not b;
    layer2_outputs(7729) <= a xor b;
    layer2_outputs(7730) <= not a;
    layer2_outputs(7731) <= '0';
    layer2_outputs(7732) <= not (a xor b);
    layer2_outputs(7733) <= '1';
    layer2_outputs(7734) <= not a;
    layer2_outputs(7735) <= b;
    layer2_outputs(7736) <= a xor b;
    layer2_outputs(7737) <= not (a or b);
    layer2_outputs(7738) <= a and not b;
    layer2_outputs(7739) <= a;
    layer2_outputs(7740) <= a;
    layer2_outputs(7741) <= not b or a;
    layer2_outputs(7742) <= b and not a;
    layer2_outputs(7743) <= not b;
    layer2_outputs(7744) <= '0';
    layer2_outputs(7745) <= not a;
    layer2_outputs(7746) <= not b;
    layer2_outputs(7747) <= not b;
    layer2_outputs(7748) <= not (a or b);
    layer2_outputs(7749) <= b;
    layer2_outputs(7750) <= a or b;
    layer2_outputs(7751) <= not (a xor b);
    layer2_outputs(7752) <= not b;
    layer2_outputs(7753) <= not (a and b);
    layer2_outputs(7754) <= a and not b;
    layer2_outputs(7755) <= a and not b;
    layer2_outputs(7756) <= not (a or b);
    layer2_outputs(7757) <= not b;
    layer2_outputs(7758) <= a and b;
    layer2_outputs(7759) <= b and not a;
    layer2_outputs(7760) <= not a;
    layer2_outputs(7761) <= not (a xor b);
    layer2_outputs(7762) <= a or b;
    layer2_outputs(7763) <= a or b;
    layer2_outputs(7764) <= not a or b;
    layer2_outputs(7765) <= a;
    layer2_outputs(7766) <= a;
    layer2_outputs(7767) <= not b;
    layer2_outputs(7768) <= a or b;
    layer2_outputs(7769) <= '0';
    layer2_outputs(7770) <= not a;
    layer2_outputs(7771) <= not (a and b);
    layer2_outputs(7772) <= not a or b;
    layer2_outputs(7773) <= not (a and b);
    layer2_outputs(7774) <= not a;
    layer2_outputs(7775) <= not a;
    layer2_outputs(7776) <= '0';
    layer2_outputs(7777) <= '1';
    layer2_outputs(7778) <= a and not b;
    layer2_outputs(7779) <= not (a or b);
    layer2_outputs(7780) <= not a;
    layer2_outputs(7781) <= not a;
    layer2_outputs(7782) <= b;
    layer2_outputs(7783) <= a or b;
    layer2_outputs(7784) <= not a;
    layer2_outputs(7785) <= a and b;
    layer2_outputs(7786) <= a or b;
    layer2_outputs(7787) <= a xor b;
    layer2_outputs(7788) <= not b;
    layer2_outputs(7789) <= a xor b;
    layer2_outputs(7790) <= b and not a;
    layer2_outputs(7791) <= a or b;
    layer2_outputs(7792) <= b and not a;
    layer2_outputs(7793) <= a or b;
    layer2_outputs(7794) <= not a;
    layer2_outputs(7795) <= a;
    layer2_outputs(7796) <= a or b;
    layer2_outputs(7797) <= a and b;
    layer2_outputs(7798) <= a and not b;
    layer2_outputs(7799) <= b and not a;
    layer2_outputs(7800) <= '1';
    layer2_outputs(7801) <= a and b;
    layer2_outputs(7802) <= not b or a;
    layer2_outputs(7803) <= '1';
    layer2_outputs(7804) <= not b or a;
    layer2_outputs(7805) <= not a;
    layer2_outputs(7806) <= not (a or b);
    layer2_outputs(7807) <= not (a or b);
    layer2_outputs(7808) <= a and not b;
    layer2_outputs(7809) <= a;
    layer2_outputs(7810) <= not b or a;
    layer2_outputs(7811) <= not a or b;
    layer2_outputs(7812) <= not (a or b);
    layer2_outputs(7813) <= b and not a;
    layer2_outputs(7814) <= not (a and b);
    layer2_outputs(7815) <= b;
    layer2_outputs(7816) <= b and not a;
    layer2_outputs(7817) <= b and not a;
    layer2_outputs(7818) <= a or b;
    layer2_outputs(7819) <= '0';
    layer2_outputs(7820) <= a and b;
    layer2_outputs(7821) <= a;
    layer2_outputs(7822) <= not (a xor b);
    layer2_outputs(7823) <= b;
    layer2_outputs(7824) <= not a;
    layer2_outputs(7825) <= not a or b;
    layer2_outputs(7826) <= a or b;
    layer2_outputs(7827) <= b and not a;
    layer2_outputs(7828) <= b and not a;
    layer2_outputs(7829) <= not (a and b);
    layer2_outputs(7830) <= not b or a;
    layer2_outputs(7831) <= a;
    layer2_outputs(7832) <= not b or a;
    layer2_outputs(7833) <= '0';
    layer2_outputs(7834) <= not (a or b);
    layer2_outputs(7835) <= not (a and b);
    layer2_outputs(7836) <= a xor b;
    layer2_outputs(7837) <= not (a and b);
    layer2_outputs(7838) <= not a;
    layer2_outputs(7839) <= a;
    layer2_outputs(7840) <= a or b;
    layer2_outputs(7841) <= a and b;
    layer2_outputs(7842) <= b;
    layer2_outputs(7843) <= not a or b;
    layer2_outputs(7844) <= b;
    layer2_outputs(7845) <= not (a or b);
    layer2_outputs(7846) <= a and b;
    layer2_outputs(7847) <= not (a or b);
    layer2_outputs(7848) <= b and not a;
    layer2_outputs(7849) <= not a;
    layer2_outputs(7850) <= not b;
    layer2_outputs(7851) <= not b or a;
    layer2_outputs(7852) <= not a or b;
    layer2_outputs(7853) <= a or b;
    layer2_outputs(7854) <= not (a and b);
    layer2_outputs(7855) <= not (a and b);
    layer2_outputs(7856) <= a and not b;
    layer2_outputs(7857) <= not a or b;
    layer2_outputs(7858) <= not (a or b);
    layer2_outputs(7859) <= not (a xor b);
    layer2_outputs(7860) <= not a;
    layer2_outputs(7861) <= '1';
    layer2_outputs(7862) <= b;
    layer2_outputs(7863) <= not a;
    layer2_outputs(7864) <= b and not a;
    layer2_outputs(7865) <= b and not a;
    layer2_outputs(7866) <= a and b;
    layer2_outputs(7867) <= a and b;
    layer2_outputs(7868) <= '1';
    layer2_outputs(7869) <= a and b;
    layer2_outputs(7870) <= '1';
    layer2_outputs(7871) <= a and not b;
    layer2_outputs(7872) <= not b;
    layer2_outputs(7873) <= a xor b;
    layer2_outputs(7874) <= not a;
    layer2_outputs(7875) <= not b;
    layer2_outputs(7876) <= a;
    layer2_outputs(7877) <= not a;
    layer2_outputs(7878) <= not (a and b);
    layer2_outputs(7879) <= not b or a;
    layer2_outputs(7880) <= b and not a;
    layer2_outputs(7881) <= a;
    layer2_outputs(7882) <= not (a xor b);
    layer2_outputs(7883) <= not a or b;
    layer2_outputs(7884) <= not b or a;
    layer2_outputs(7885) <= a and b;
    layer2_outputs(7886) <= not a or b;
    layer2_outputs(7887) <= not a;
    layer2_outputs(7888) <= b;
    layer2_outputs(7889) <= a or b;
    layer2_outputs(7890) <= not (a or b);
    layer2_outputs(7891) <= b and not a;
    layer2_outputs(7892) <= not a or b;
    layer2_outputs(7893) <= not (a and b);
    layer2_outputs(7894) <= not (a or b);
    layer2_outputs(7895) <= not b;
    layer2_outputs(7896) <= not a;
    layer2_outputs(7897) <= not b or a;
    layer2_outputs(7898) <= not (a or b);
    layer2_outputs(7899) <= '1';
    layer2_outputs(7900) <= a or b;
    layer2_outputs(7901) <= not (a and b);
    layer2_outputs(7902) <= not a;
    layer2_outputs(7903) <= a;
    layer2_outputs(7904) <= b and not a;
    layer2_outputs(7905) <= '0';
    layer2_outputs(7906) <= not (a or b);
    layer2_outputs(7907) <= '1';
    layer2_outputs(7908) <= a and b;
    layer2_outputs(7909) <= a;
    layer2_outputs(7910) <= not b;
    layer2_outputs(7911) <= '0';
    layer2_outputs(7912) <= not a or b;
    layer2_outputs(7913) <= b and not a;
    layer2_outputs(7914) <= a;
    layer2_outputs(7915) <= a or b;
    layer2_outputs(7916) <= not (a and b);
    layer2_outputs(7917) <= a;
    layer2_outputs(7918) <= not b;
    layer2_outputs(7919) <= not a;
    layer2_outputs(7920) <= a and not b;
    layer2_outputs(7921) <= not a;
    layer2_outputs(7922) <= not (a or b);
    layer2_outputs(7923) <= b;
    layer2_outputs(7924) <= a and not b;
    layer2_outputs(7925) <= a and b;
    layer2_outputs(7926) <= not b or a;
    layer2_outputs(7927) <= '0';
    layer2_outputs(7928) <= not b or a;
    layer2_outputs(7929) <= not b;
    layer2_outputs(7930) <= b and not a;
    layer2_outputs(7931) <= a;
    layer2_outputs(7932) <= b;
    layer2_outputs(7933) <= not b;
    layer2_outputs(7934) <= a and b;
    layer2_outputs(7935) <= a;
    layer2_outputs(7936) <= not (a or b);
    layer2_outputs(7937) <= b;
    layer2_outputs(7938) <= '1';
    layer2_outputs(7939) <= not a;
    layer2_outputs(7940) <= '0';
    layer2_outputs(7941) <= not a;
    layer2_outputs(7942) <= a or b;
    layer2_outputs(7943) <= b and not a;
    layer2_outputs(7944) <= not b;
    layer2_outputs(7945) <= not a;
    layer2_outputs(7946) <= not a;
    layer2_outputs(7947) <= not (a and b);
    layer2_outputs(7948) <= not b or a;
    layer2_outputs(7949) <= a;
    layer2_outputs(7950) <= not a or b;
    layer2_outputs(7951) <= not b;
    layer2_outputs(7952) <= not (a or b);
    layer2_outputs(7953) <= b and not a;
    layer2_outputs(7954) <= not b;
    layer2_outputs(7955) <= not a;
    layer2_outputs(7956) <= a or b;
    layer2_outputs(7957) <= b and not a;
    layer2_outputs(7958) <= b;
    layer2_outputs(7959) <= b and not a;
    layer2_outputs(7960) <= not a or b;
    layer2_outputs(7961) <= a and not b;
    layer2_outputs(7962) <= b;
    layer2_outputs(7963) <= not (a and b);
    layer2_outputs(7964) <= not (a and b);
    layer2_outputs(7965) <= not b or a;
    layer2_outputs(7966) <= not b or a;
    layer2_outputs(7967) <= a and b;
    layer2_outputs(7968) <= not b;
    layer2_outputs(7969) <= not (a or b);
    layer2_outputs(7970) <= '1';
    layer2_outputs(7971) <= a;
    layer2_outputs(7972) <= a and not b;
    layer2_outputs(7973) <= a and b;
    layer2_outputs(7974) <= not a;
    layer2_outputs(7975) <= a and b;
    layer2_outputs(7976) <= a;
    layer2_outputs(7977) <= a;
    layer2_outputs(7978) <= not (a and b);
    layer2_outputs(7979) <= not a or b;
    layer2_outputs(7980) <= a and b;
    layer2_outputs(7981) <= not (a xor b);
    layer2_outputs(7982) <= '0';
    layer2_outputs(7983) <= '1';
    layer2_outputs(7984) <= not b;
    layer2_outputs(7985) <= a and b;
    layer2_outputs(7986) <= not (a and b);
    layer2_outputs(7987) <= not a;
    layer2_outputs(7988) <= not (a or b);
    layer2_outputs(7989) <= not b;
    layer2_outputs(7990) <= not b;
    layer2_outputs(7991) <= not b;
    layer2_outputs(7992) <= a;
    layer2_outputs(7993) <= not b;
    layer2_outputs(7994) <= b;
    layer2_outputs(7995) <= a and b;
    layer2_outputs(7996) <= a xor b;
    layer2_outputs(7997) <= not a or b;
    layer2_outputs(7998) <= not b;
    layer2_outputs(7999) <= not b;
    layer2_outputs(8000) <= b and not a;
    layer2_outputs(8001) <= not a;
    layer2_outputs(8002) <= a and b;
    layer2_outputs(8003) <= a or b;
    layer2_outputs(8004) <= not a or b;
    layer2_outputs(8005) <= '1';
    layer2_outputs(8006) <= not b;
    layer2_outputs(8007) <= not (a and b);
    layer2_outputs(8008) <= a and not b;
    layer2_outputs(8009) <= b and not a;
    layer2_outputs(8010) <= a and b;
    layer2_outputs(8011) <= not (a or b);
    layer2_outputs(8012) <= not (a or b);
    layer2_outputs(8013) <= not (a or b);
    layer2_outputs(8014) <= a and b;
    layer2_outputs(8015) <= b;
    layer2_outputs(8016) <= a xor b;
    layer2_outputs(8017) <= not a or b;
    layer2_outputs(8018) <= '0';
    layer2_outputs(8019) <= '0';
    layer2_outputs(8020) <= b;
    layer2_outputs(8021) <= a and b;
    layer2_outputs(8022) <= a and not b;
    layer2_outputs(8023) <= b and not a;
    layer2_outputs(8024) <= '0';
    layer2_outputs(8025) <= not b;
    layer2_outputs(8026) <= b and not a;
    layer2_outputs(8027) <= '1';
    layer2_outputs(8028) <= '0';
    layer2_outputs(8029) <= '1';
    layer2_outputs(8030) <= a;
    layer2_outputs(8031) <= a;
    layer2_outputs(8032) <= b;
    layer2_outputs(8033) <= not (a xor b);
    layer2_outputs(8034) <= a xor b;
    layer2_outputs(8035) <= a and b;
    layer2_outputs(8036) <= not a;
    layer2_outputs(8037) <= not a;
    layer2_outputs(8038) <= not (a or b);
    layer2_outputs(8039) <= '0';
    layer2_outputs(8040) <= '1';
    layer2_outputs(8041) <= not b;
    layer2_outputs(8042) <= a xor b;
    layer2_outputs(8043) <= a and not b;
    layer2_outputs(8044) <= a or b;
    layer2_outputs(8045) <= not a or b;
    layer2_outputs(8046) <= a;
    layer2_outputs(8047) <= not a;
    layer2_outputs(8048) <= '1';
    layer2_outputs(8049) <= b;
    layer2_outputs(8050) <= not (a and b);
    layer2_outputs(8051) <= not a;
    layer2_outputs(8052) <= not a;
    layer2_outputs(8053) <= a and b;
    layer2_outputs(8054) <= b;
    layer2_outputs(8055) <= not (a and b);
    layer2_outputs(8056) <= a;
    layer2_outputs(8057) <= not b;
    layer2_outputs(8058) <= not a;
    layer2_outputs(8059) <= '1';
    layer2_outputs(8060) <= not (a and b);
    layer2_outputs(8061) <= not (a and b);
    layer2_outputs(8062) <= b and not a;
    layer2_outputs(8063) <= a and b;
    layer2_outputs(8064) <= b;
    layer2_outputs(8065) <= not b;
    layer2_outputs(8066) <= a;
    layer2_outputs(8067) <= a;
    layer2_outputs(8068) <= a;
    layer2_outputs(8069) <= a and not b;
    layer2_outputs(8070) <= '1';
    layer2_outputs(8071) <= '1';
    layer2_outputs(8072) <= a and not b;
    layer2_outputs(8073) <= not a;
    layer2_outputs(8074) <= not a;
    layer2_outputs(8075) <= b and not a;
    layer2_outputs(8076) <= not b or a;
    layer2_outputs(8077) <= a;
    layer2_outputs(8078) <= not (a xor b);
    layer2_outputs(8079) <= not (a and b);
    layer2_outputs(8080) <= b;
    layer2_outputs(8081) <= a;
    layer2_outputs(8082) <= '0';
    layer2_outputs(8083) <= '0';
    layer2_outputs(8084) <= a xor b;
    layer2_outputs(8085) <= '0';
    layer2_outputs(8086) <= a and not b;
    layer2_outputs(8087) <= '0';
    layer2_outputs(8088) <= '1';
    layer2_outputs(8089) <= '0';
    layer2_outputs(8090) <= not b or a;
    layer2_outputs(8091) <= not (a and b);
    layer2_outputs(8092) <= not a;
    layer2_outputs(8093) <= not (a or b);
    layer2_outputs(8094) <= not (a and b);
    layer2_outputs(8095) <= b;
    layer2_outputs(8096) <= a or b;
    layer2_outputs(8097) <= a;
    layer2_outputs(8098) <= a and b;
    layer2_outputs(8099) <= not b or a;
    layer2_outputs(8100) <= not b;
    layer2_outputs(8101) <= not b;
    layer2_outputs(8102) <= a and b;
    layer2_outputs(8103) <= b and not a;
    layer2_outputs(8104) <= not (a or b);
    layer2_outputs(8105) <= a;
    layer2_outputs(8106) <= '1';
    layer2_outputs(8107) <= not (a xor b);
    layer2_outputs(8108) <= a or b;
    layer2_outputs(8109) <= a;
    layer2_outputs(8110) <= not b or a;
    layer2_outputs(8111) <= not a or b;
    layer2_outputs(8112) <= not a or b;
    layer2_outputs(8113) <= not (a xor b);
    layer2_outputs(8114) <= a and not b;
    layer2_outputs(8115) <= not (a and b);
    layer2_outputs(8116) <= not a;
    layer2_outputs(8117) <= not a;
    layer2_outputs(8118) <= a and b;
    layer2_outputs(8119) <= not b;
    layer2_outputs(8120) <= not (a xor b);
    layer2_outputs(8121) <= b;
    layer2_outputs(8122) <= a and b;
    layer2_outputs(8123) <= not (a or b);
    layer2_outputs(8124) <= a;
    layer2_outputs(8125) <= a and not b;
    layer2_outputs(8126) <= a;
    layer2_outputs(8127) <= not a;
    layer2_outputs(8128) <= not (a and b);
    layer2_outputs(8129) <= not a;
    layer2_outputs(8130) <= not a;
    layer2_outputs(8131) <= a and not b;
    layer2_outputs(8132) <= not a or b;
    layer2_outputs(8133) <= not b;
    layer2_outputs(8134) <= a xor b;
    layer2_outputs(8135) <= a or b;
    layer2_outputs(8136) <= not b;
    layer2_outputs(8137) <= '0';
    layer2_outputs(8138) <= a or b;
    layer2_outputs(8139) <= a and b;
    layer2_outputs(8140) <= a xor b;
    layer2_outputs(8141) <= not a or b;
    layer2_outputs(8142) <= not a or b;
    layer2_outputs(8143) <= not a or b;
    layer2_outputs(8144) <= b;
    layer2_outputs(8145) <= not a or b;
    layer2_outputs(8146) <= b and not a;
    layer2_outputs(8147) <= '0';
    layer2_outputs(8148) <= b and not a;
    layer2_outputs(8149) <= b and not a;
    layer2_outputs(8150) <= not a;
    layer2_outputs(8151) <= not b or a;
    layer2_outputs(8152) <= not (a and b);
    layer2_outputs(8153) <= a and b;
    layer2_outputs(8154) <= not (a and b);
    layer2_outputs(8155) <= not b;
    layer2_outputs(8156) <= b;
    layer2_outputs(8157) <= not a;
    layer2_outputs(8158) <= not a;
    layer2_outputs(8159) <= not b;
    layer2_outputs(8160) <= not (a xor b);
    layer2_outputs(8161) <= not b;
    layer2_outputs(8162) <= a and not b;
    layer2_outputs(8163) <= not b;
    layer2_outputs(8164) <= a or b;
    layer2_outputs(8165) <= a and not b;
    layer2_outputs(8166) <= b;
    layer2_outputs(8167) <= not (a xor b);
    layer2_outputs(8168) <= not (a or b);
    layer2_outputs(8169) <= '0';
    layer2_outputs(8170) <= b and not a;
    layer2_outputs(8171) <= not b or a;
    layer2_outputs(8172) <= not b or a;
    layer2_outputs(8173) <= not (a or b);
    layer2_outputs(8174) <= '1';
    layer2_outputs(8175) <= not (a or b);
    layer2_outputs(8176) <= not a or b;
    layer2_outputs(8177) <= not b or a;
    layer2_outputs(8178) <= not (a and b);
    layer2_outputs(8179) <= not b or a;
    layer2_outputs(8180) <= not (a or b);
    layer2_outputs(8181) <= a;
    layer2_outputs(8182) <= a and not b;
    layer2_outputs(8183) <= not (a and b);
    layer2_outputs(8184) <= not (a xor b);
    layer2_outputs(8185) <= a and b;
    layer2_outputs(8186) <= a and b;
    layer2_outputs(8187) <= '1';
    layer2_outputs(8188) <= not (a and b);
    layer2_outputs(8189) <= not a;
    layer2_outputs(8190) <= a and b;
    layer2_outputs(8191) <= not a or b;
    layer2_outputs(8192) <= a xor b;
    layer2_outputs(8193) <= a or b;
    layer2_outputs(8194) <= not a;
    layer2_outputs(8195) <= a;
    layer2_outputs(8196) <= not b or a;
    layer2_outputs(8197) <= a and b;
    layer2_outputs(8198) <= a and b;
    layer2_outputs(8199) <= not a;
    layer2_outputs(8200) <= a or b;
    layer2_outputs(8201) <= b and not a;
    layer2_outputs(8202) <= not (a and b);
    layer2_outputs(8203) <= not a;
    layer2_outputs(8204) <= not a;
    layer2_outputs(8205) <= a or b;
    layer2_outputs(8206) <= a;
    layer2_outputs(8207) <= not a or b;
    layer2_outputs(8208) <= not a;
    layer2_outputs(8209) <= a xor b;
    layer2_outputs(8210) <= a;
    layer2_outputs(8211) <= a xor b;
    layer2_outputs(8212) <= not (a and b);
    layer2_outputs(8213) <= a or b;
    layer2_outputs(8214) <= b;
    layer2_outputs(8215) <= a xor b;
    layer2_outputs(8216) <= b;
    layer2_outputs(8217) <= a;
    layer2_outputs(8218) <= a;
    layer2_outputs(8219) <= a;
    layer2_outputs(8220) <= a;
    layer2_outputs(8221) <= a or b;
    layer2_outputs(8222) <= a;
    layer2_outputs(8223) <= a xor b;
    layer2_outputs(8224) <= not b;
    layer2_outputs(8225) <= not b;
    layer2_outputs(8226) <= a or b;
    layer2_outputs(8227) <= not b;
    layer2_outputs(8228) <= '0';
    layer2_outputs(8229) <= b and not a;
    layer2_outputs(8230) <= '0';
    layer2_outputs(8231) <= not a;
    layer2_outputs(8232) <= not (a or b);
    layer2_outputs(8233) <= not b;
    layer2_outputs(8234) <= a and b;
    layer2_outputs(8235) <= not a or b;
    layer2_outputs(8236) <= b and not a;
    layer2_outputs(8237) <= not b or a;
    layer2_outputs(8238) <= not b;
    layer2_outputs(8239) <= not b;
    layer2_outputs(8240) <= not a;
    layer2_outputs(8241) <= '1';
    layer2_outputs(8242) <= not a;
    layer2_outputs(8243) <= a and not b;
    layer2_outputs(8244) <= not b;
    layer2_outputs(8245) <= a and b;
    layer2_outputs(8246) <= '1';
    layer2_outputs(8247) <= not b or a;
    layer2_outputs(8248) <= b;
    layer2_outputs(8249) <= b and not a;
    layer2_outputs(8250) <= b;
    layer2_outputs(8251) <= a or b;
    layer2_outputs(8252) <= '0';
    layer2_outputs(8253) <= a or b;
    layer2_outputs(8254) <= a and not b;
    layer2_outputs(8255) <= not a or b;
    layer2_outputs(8256) <= a and b;
    layer2_outputs(8257) <= a xor b;
    layer2_outputs(8258) <= a and b;
    layer2_outputs(8259) <= not b or a;
    layer2_outputs(8260) <= not b;
    layer2_outputs(8261) <= '1';
    layer2_outputs(8262) <= a and b;
    layer2_outputs(8263) <= not a or b;
    layer2_outputs(8264) <= not b;
    layer2_outputs(8265) <= a and not b;
    layer2_outputs(8266) <= a xor b;
    layer2_outputs(8267) <= not (a xor b);
    layer2_outputs(8268) <= a and b;
    layer2_outputs(8269) <= a or b;
    layer2_outputs(8270) <= b and not a;
    layer2_outputs(8271) <= not (a and b);
    layer2_outputs(8272) <= '1';
    layer2_outputs(8273) <= a;
    layer2_outputs(8274) <= not (a and b);
    layer2_outputs(8275) <= b;
    layer2_outputs(8276) <= not a or b;
    layer2_outputs(8277) <= not a;
    layer2_outputs(8278) <= '0';
    layer2_outputs(8279) <= a xor b;
    layer2_outputs(8280) <= not a or b;
    layer2_outputs(8281) <= b;
    layer2_outputs(8282) <= b;
    layer2_outputs(8283) <= a;
    layer2_outputs(8284) <= a and b;
    layer2_outputs(8285) <= b;
    layer2_outputs(8286) <= '0';
    layer2_outputs(8287) <= a and not b;
    layer2_outputs(8288) <= not a;
    layer2_outputs(8289) <= a and not b;
    layer2_outputs(8290) <= not a;
    layer2_outputs(8291) <= b;
    layer2_outputs(8292) <= a;
    layer2_outputs(8293) <= '1';
    layer2_outputs(8294) <= b and not a;
    layer2_outputs(8295) <= '1';
    layer2_outputs(8296) <= not a;
    layer2_outputs(8297) <= not a or b;
    layer2_outputs(8298) <= a xor b;
    layer2_outputs(8299) <= not b;
    layer2_outputs(8300) <= not b;
    layer2_outputs(8301) <= not b;
    layer2_outputs(8302) <= not (a and b);
    layer2_outputs(8303) <= a and b;
    layer2_outputs(8304) <= not (a xor b);
    layer2_outputs(8305) <= not b or a;
    layer2_outputs(8306) <= a and b;
    layer2_outputs(8307) <= not b;
    layer2_outputs(8308) <= not b or a;
    layer2_outputs(8309) <= not b or a;
    layer2_outputs(8310) <= '1';
    layer2_outputs(8311) <= not a;
    layer2_outputs(8312) <= a;
    layer2_outputs(8313) <= a and b;
    layer2_outputs(8314) <= not b;
    layer2_outputs(8315) <= not (a xor b);
    layer2_outputs(8316) <= '0';
    layer2_outputs(8317) <= not b;
    layer2_outputs(8318) <= not (a or b);
    layer2_outputs(8319) <= '0';
    layer2_outputs(8320) <= not a or b;
    layer2_outputs(8321) <= a and b;
    layer2_outputs(8322) <= not (a and b);
    layer2_outputs(8323) <= '1';
    layer2_outputs(8324) <= not (a or b);
    layer2_outputs(8325) <= a or b;
    layer2_outputs(8326) <= '1';
    layer2_outputs(8327) <= a xor b;
    layer2_outputs(8328) <= a;
    layer2_outputs(8329) <= '1';
    layer2_outputs(8330) <= not a or b;
    layer2_outputs(8331) <= not b or a;
    layer2_outputs(8332) <= b;
    layer2_outputs(8333) <= b;
    layer2_outputs(8334) <= not b or a;
    layer2_outputs(8335) <= a and not b;
    layer2_outputs(8336) <= not b or a;
    layer2_outputs(8337) <= a xor b;
    layer2_outputs(8338) <= a and not b;
    layer2_outputs(8339) <= a xor b;
    layer2_outputs(8340) <= a xor b;
    layer2_outputs(8341) <= not a;
    layer2_outputs(8342) <= not b or a;
    layer2_outputs(8343) <= not (a xor b);
    layer2_outputs(8344) <= a or b;
    layer2_outputs(8345) <= '1';
    layer2_outputs(8346) <= a;
    layer2_outputs(8347) <= not (a xor b);
    layer2_outputs(8348) <= '1';
    layer2_outputs(8349) <= a or b;
    layer2_outputs(8350) <= not a;
    layer2_outputs(8351) <= b and not a;
    layer2_outputs(8352) <= not (a and b);
    layer2_outputs(8353) <= b;
    layer2_outputs(8354) <= '0';
    layer2_outputs(8355) <= not a;
    layer2_outputs(8356) <= '1';
    layer2_outputs(8357) <= a or b;
    layer2_outputs(8358) <= a or b;
    layer2_outputs(8359) <= b and not a;
    layer2_outputs(8360) <= not (a xor b);
    layer2_outputs(8361) <= a or b;
    layer2_outputs(8362) <= a and not b;
    layer2_outputs(8363) <= '0';
    layer2_outputs(8364) <= a;
    layer2_outputs(8365) <= a and not b;
    layer2_outputs(8366) <= a;
    layer2_outputs(8367) <= a and not b;
    layer2_outputs(8368) <= '1';
    layer2_outputs(8369) <= b and not a;
    layer2_outputs(8370) <= '1';
    layer2_outputs(8371) <= a xor b;
    layer2_outputs(8372) <= not a;
    layer2_outputs(8373) <= not b or a;
    layer2_outputs(8374) <= a and b;
    layer2_outputs(8375) <= a;
    layer2_outputs(8376) <= a;
    layer2_outputs(8377) <= a and b;
    layer2_outputs(8378) <= '0';
    layer2_outputs(8379) <= a xor b;
    layer2_outputs(8380) <= not a;
    layer2_outputs(8381) <= '0';
    layer2_outputs(8382) <= b and not a;
    layer2_outputs(8383) <= a and not b;
    layer2_outputs(8384) <= a;
    layer2_outputs(8385) <= not (a or b);
    layer2_outputs(8386) <= not (a and b);
    layer2_outputs(8387) <= not b;
    layer2_outputs(8388) <= b;
    layer2_outputs(8389) <= not b;
    layer2_outputs(8390) <= a and b;
    layer2_outputs(8391) <= a and not b;
    layer2_outputs(8392) <= not (a or b);
    layer2_outputs(8393) <= b;
    layer2_outputs(8394) <= a;
    layer2_outputs(8395) <= a or b;
    layer2_outputs(8396) <= '1';
    layer2_outputs(8397) <= not (a and b);
    layer2_outputs(8398) <= not (a and b);
    layer2_outputs(8399) <= b and not a;
    layer2_outputs(8400) <= b;
    layer2_outputs(8401) <= not b;
    layer2_outputs(8402) <= b;
    layer2_outputs(8403) <= not a or b;
    layer2_outputs(8404) <= not b or a;
    layer2_outputs(8405) <= not b;
    layer2_outputs(8406) <= not (a xor b);
    layer2_outputs(8407) <= a;
    layer2_outputs(8408) <= not (a or b);
    layer2_outputs(8409) <= a and not b;
    layer2_outputs(8410) <= b and not a;
    layer2_outputs(8411) <= a or b;
    layer2_outputs(8412) <= b;
    layer2_outputs(8413) <= a;
    layer2_outputs(8414) <= not a;
    layer2_outputs(8415) <= '0';
    layer2_outputs(8416) <= a and not b;
    layer2_outputs(8417) <= not a or b;
    layer2_outputs(8418) <= not a or b;
    layer2_outputs(8419) <= not a or b;
    layer2_outputs(8420) <= a xor b;
    layer2_outputs(8421) <= a and b;
    layer2_outputs(8422) <= not (a xor b);
    layer2_outputs(8423) <= not a;
    layer2_outputs(8424) <= a;
    layer2_outputs(8425) <= not a;
    layer2_outputs(8426) <= not b or a;
    layer2_outputs(8427) <= not b;
    layer2_outputs(8428) <= not a or b;
    layer2_outputs(8429) <= not b or a;
    layer2_outputs(8430) <= not (a or b);
    layer2_outputs(8431) <= not a or b;
    layer2_outputs(8432) <= not a;
    layer2_outputs(8433) <= not a or b;
    layer2_outputs(8434) <= b;
    layer2_outputs(8435) <= b and not a;
    layer2_outputs(8436) <= a and b;
    layer2_outputs(8437) <= b;
    layer2_outputs(8438) <= not (a and b);
    layer2_outputs(8439) <= a;
    layer2_outputs(8440) <= a;
    layer2_outputs(8441) <= not a or b;
    layer2_outputs(8442) <= '1';
    layer2_outputs(8443) <= '0';
    layer2_outputs(8444) <= not (a and b);
    layer2_outputs(8445) <= not b;
    layer2_outputs(8446) <= a xor b;
    layer2_outputs(8447) <= '1';
    layer2_outputs(8448) <= not b;
    layer2_outputs(8449) <= not b;
    layer2_outputs(8450) <= a;
    layer2_outputs(8451) <= b and not a;
    layer2_outputs(8452) <= b;
    layer2_outputs(8453) <= a and b;
    layer2_outputs(8454) <= a and b;
    layer2_outputs(8455) <= a xor b;
    layer2_outputs(8456) <= not a;
    layer2_outputs(8457) <= a;
    layer2_outputs(8458) <= not b or a;
    layer2_outputs(8459) <= b;
    layer2_outputs(8460) <= a;
    layer2_outputs(8461) <= '1';
    layer2_outputs(8462) <= b and not a;
    layer2_outputs(8463) <= not a;
    layer2_outputs(8464) <= a and b;
    layer2_outputs(8465) <= '1';
    layer2_outputs(8466) <= a;
    layer2_outputs(8467) <= '1';
    layer2_outputs(8468) <= b;
    layer2_outputs(8469) <= not b;
    layer2_outputs(8470) <= a;
    layer2_outputs(8471) <= not a;
    layer2_outputs(8472) <= not b or a;
    layer2_outputs(8473) <= b and not a;
    layer2_outputs(8474) <= not (a and b);
    layer2_outputs(8475) <= not a;
    layer2_outputs(8476) <= not b;
    layer2_outputs(8477) <= b;
    layer2_outputs(8478) <= a and b;
    layer2_outputs(8479) <= a xor b;
    layer2_outputs(8480) <= not b or a;
    layer2_outputs(8481) <= '0';
    layer2_outputs(8482) <= not b or a;
    layer2_outputs(8483) <= not b or a;
    layer2_outputs(8484) <= not (a or b);
    layer2_outputs(8485) <= a or b;
    layer2_outputs(8486) <= not (a or b);
    layer2_outputs(8487) <= a and not b;
    layer2_outputs(8488) <= not (a or b);
    layer2_outputs(8489) <= not a;
    layer2_outputs(8490) <= not a;
    layer2_outputs(8491) <= a;
    layer2_outputs(8492) <= not (a and b);
    layer2_outputs(8493) <= '0';
    layer2_outputs(8494) <= a and not b;
    layer2_outputs(8495) <= not a;
    layer2_outputs(8496) <= not (a and b);
    layer2_outputs(8497) <= b;
    layer2_outputs(8498) <= a or b;
    layer2_outputs(8499) <= a and b;
    layer2_outputs(8500) <= b and not a;
    layer2_outputs(8501) <= not (a or b);
    layer2_outputs(8502) <= b;
    layer2_outputs(8503) <= not a;
    layer2_outputs(8504) <= a and b;
    layer2_outputs(8505) <= b and not a;
    layer2_outputs(8506) <= not a;
    layer2_outputs(8507) <= a and not b;
    layer2_outputs(8508) <= not (a and b);
    layer2_outputs(8509) <= b;
    layer2_outputs(8510) <= a and not b;
    layer2_outputs(8511) <= not a;
    layer2_outputs(8512) <= not (a or b);
    layer2_outputs(8513) <= not b or a;
    layer2_outputs(8514) <= not (a and b);
    layer2_outputs(8515) <= '0';
    layer2_outputs(8516) <= '0';
    layer2_outputs(8517) <= b and not a;
    layer2_outputs(8518) <= not (a and b);
    layer2_outputs(8519) <= a and b;
    layer2_outputs(8520) <= a or b;
    layer2_outputs(8521) <= not a or b;
    layer2_outputs(8522) <= not (a or b);
    layer2_outputs(8523) <= a;
    layer2_outputs(8524) <= not b or a;
    layer2_outputs(8525) <= not b or a;
    layer2_outputs(8526) <= a or b;
    layer2_outputs(8527) <= not a or b;
    layer2_outputs(8528) <= not b or a;
    layer2_outputs(8529) <= b;
    layer2_outputs(8530) <= b;
    layer2_outputs(8531) <= b and not a;
    layer2_outputs(8532) <= '1';
    layer2_outputs(8533) <= not a or b;
    layer2_outputs(8534) <= not a or b;
    layer2_outputs(8535) <= not a or b;
    layer2_outputs(8536) <= a;
    layer2_outputs(8537) <= a or b;
    layer2_outputs(8538) <= not a or b;
    layer2_outputs(8539) <= not a;
    layer2_outputs(8540) <= not b;
    layer2_outputs(8541) <= b;
    layer2_outputs(8542) <= b;
    layer2_outputs(8543) <= not a or b;
    layer2_outputs(8544) <= not b;
    layer2_outputs(8545) <= a xor b;
    layer2_outputs(8546) <= not b;
    layer2_outputs(8547) <= not (a or b);
    layer2_outputs(8548) <= b and not a;
    layer2_outputs(8549) <= a and b;
    layer2_outputs(8550) <= b and not a;
    layer2_outputs(8551) <= a;
    layer2_outputs(8552) <= a;
    layer2_outputs(8553) <= b;
    layer2_outputs(8554) <= not b or a;
    layer2_outputs(8555) <= '0';
    layer2_outputs(8556) <= not a or b;
    layer2_outputs(8557) <= b;
    layer2_outputs(8558) <= a or b;
    layer2_outputs(8559) <= not (a and b);
    layer2_outputs(8560) <= not (a xor b);
    layer2_outputs(8561) <= not (a or b);
    layer2_outputs(8562) <= not b;
    layer2_outputs(8563) <= not (a and b);
    layer2_outputs(8564) <= b and not a;
    layer2_outputs(8565) <= a xor b;
    layer2_outputs(8566) <= a or b;
    layer2_outputs(8567) <= a;
    layer2_outputs(8568) <= a and not b;
    layer2_outputs(8569) <= b and not a;
    layer2_outputs(8570) <= not a or b;
    layer2_outputs(8571) <= not a or b;
    layer2_outputs(8572) <= not b;
    layer2_outputs(8573) <= not b;
    layer2_outputs(8574) <= not a;
    layer2_outputs(8575) <= not a or b;
    layer2_outputs(8576) <= not (a or b);
    layer2_outputs(8577) <= not a or b;
    layer2_outputs(8578) <= '1';
    layer2_outputs(8579) <= b;
    layer2_outputs(8580) <= not b;
    layer2_outputs(8581) <= a;
    layer2_outputs(8582) <= not a;
    layer2_outputs(8583) <= '0';
    layer2_outputs(8584) <= a or b;
    layer2_outputs(8585) <= a;
    layer2_outputs(8586) <= not a or b;
    layer2_outputs(8587) <= not b or a;
    layer2_outputs(8588) <= a and not b;
    layer2_outputs(8589) <= not b or a;
    layer2_outputs(8590) <= a or b;
    layer2_outputs(8591) <= not a;
    layer2_outputs(8592) <= b;
    layer2_outputs(8593) <= a or b;
    layer2_outputs(8594) <= a;
    layer2_outputs(8595) <= not b or a;
    layer2_outputs(8596) <= b and not a;
    layer2_outputs(8597) <= a and b;
    layer2_outputs(8598) <= not (a or b);
    layer2_outputs(8599) <= not a;
    layer2_outputs(8600) <= b;
    layer2_outputs(8601) <= b;
    layer2_outputs(8602) <= a or b;
    layer2_outputs(8603) <= not (a or b);
    layer2_outputs(8604) <= a;
    layer2_outputs(8605) <= b;
    layer2_outputs(8606) <= not (a or b);
    layer2_outputs(8607) <= not b or a;
    layer2_outputs(8608) <= b;
    layer2_outputs(8609) <= '1';
    layer2_outputs(8610) <= not a or b;
    layer2_outputs(8611) <= not a or b;
    layer2_outputs(8612) <= a xor b;
    layer2_outputs(8613) <= not a;
    layer2_outputs(8614) <= a and b;
    layer2_outputs(8615) <= not a;
    layer2_outputs(8616) <= b and not a;
    layer2_outputs(8617) <= not a;
    layer2_outputs(8618) <= b and not a;
    layer2_outputs(8619) <= a and b;
    layer2_outputs(8620) <= not (a xor b);
    layer2_outputs(8621) <= not b or a;
    layer2_outputs(8622) <= not a;
    layer2_outputs(8623) <= not b;
    layer2_outputs(8624) <= not a;
    layer2_outputs(8625) <= not (a or b);
    layer2_outputs(8626) <= not a;
    layer2_outputs(8627) <= not b;
    layer2_outputs(8628) <= a;
    layer2_outputs(8629) <= a;
    layer2_outputs(8630) <= not a;
    layer2_outputs(8631) <= '1';
    layer2_outputs(8632) <= not (a or b);
    layer2_outputs(8633) <= not (a xor b);
    layer2_outputs(8634) <= not (a xor b);
    layer2_outputs(8635) <= a or b;
    layer2_outputs(8636) <= not a or b;
    layer2_outputs(8637) <= b;
    layer2_outputs(8638) <= '0';
    layer2_outputs(8639) <= not b or a;
    layer2_outputs(8640) <= not (a and b);
    layer2_outputs(8641) <= not a;
    layer2_outputs(8642) <= b and not a;
    layer2_outputs(8643) <= b and not a;
    layer2_outputs(8644) <= not (a and b);
    layer2_outputs(8645) <= not b or a;
    layer2_outputs(8646) <= '1';
    layer2_outputs(8647) <= not b or a;
    layer2_outputs(8648) <= not b or a;
    layer2_outputs(8649) <= a and b;
    layer2_outputs(8650) <= not a or b;
    layer2_outputs(8651) <= '1';
    layer2_outputs(8652) <= not b;
    layer2_outputs(8653) <= not a or b;
    layer2_outputs(8654) <= not (a xor b);
    layer2_outputs(8655) <= a and not b;
    layer2_outputs(8656) <= not b;
    layer2_outputs(8657) <= not b or a;
    layer2_outputs(8658) <= '1';
    layer2_outputs(8659) <= b;
    layer2_outputs(8660) <= not a;
    layer2_outputs(8661) <= not a;
    layer2_outputs(8662) <= not b;
    layer2_outputs(8663) <= not b or a;
    layer2_outputs(8664) <= b;
    layer2_outputs(8665) <= a and b;
    layer2_outputs(8666) <= not a;
    layer2_outputs(8667) <= b;
    layer2_outputs(8668) <= not b;
    layer2_outputs(8669) <= b and not a;
    layer2_outputs(8670) <= not (a and b);
    layer2_outputs(8671) <= a and b;
    layer2_outputs(8672) <= not a;
    layer2_outputs(8673) <= a;
    layer2_outputs(8674) <= not b or a;
    layer2_outputs(8675) <= a and not b;
    layer2_outputs(8676) <= a;
    layer2_outputs(8677) <= '1';
    layer2_outputs(8678) <= a;
    layer2_outputs(8679) <= not b or a;
    layer2_outputs(8680) <= a xor b;
    layer2_outputs(8681) <= '1';
    layer2_outputs(8682) <= not (a and b);
    layer2_outputs(8683) <= '0';
    layer2_outputs(8684) <= a;
    layer2_outputs(8685) <= not a;
    layer2_outputs(8686) <= b;
    layer2_outputs(8687) <= a;
    layer2_outputs(8688) <= b;
    layer2_outputs(8689) <= '1';
    layer2_outputs(8690) <= a and b;
    layer2_outputs(8691) <= '0';
    layer2_outputs(8692) <= not b;
    layer2_outputs(8693) <= a;
    layer2_outputs(8694) <= b;
    layer2_outputs(8695) <= not a;
    layer2_outputs(8696) <= not (a or b);
    layer2_outputs(8697) <= not (a and b);
    layer2_outputs(8698) <= a or b;
    layer2_outputs(8699) <= '0';
    layer2_outputs(8700) <= not a or b;
    layer2_outputs(8701) <= a or b;
    layer2_outputs(8702) <= not b;
    layer2_outputs(8703) <= a xor b;
    layer2_outputs(8704) <= b;
    layer2_outputs(8705) <= not a or b;
    layer2_outputs(8706) <= b;
    layer2_outputs(8707) <= not b;
    layer2_outputs(8708) <= b;
    layer2_outputs(8709) <= not b;
    layer2_outputs(8710) <= not a;
    layer2_outputs(8711) <= a;
    layer2_outputs(8712) <= b;
    layer2_outputs(8713) <= not b or a;
    layer2_outputs(8714) <= a and b;
    layer2_outputs(8715) <= a and b;
    layer2_outputs(8716) <= a and not b;
    layer2_outputs(8717) <= a and b;
    layer2_outputs(8718) <= not (a and b);
    layer2_outputs(8719) <= '0';
    layer2_outputs(8720) <= not (a and b);
    layer2_outputs(8721) <= b and not a;
    layer2_outputs(8722) <= a or b;
    layer2_outputs(8723) <= not a or b;
    layer2_outputs(8724) <= not b;
    layer2_outputs(8725) <= '0';
    layer2_outputs(8726) <= not b;
    layer2_outputs(8727) <= a and not b;
    layer2_outputs(8728) <= a;
    layer2_outputs(8729) <= a and not b;
    layer2_outputs(8730) <= '0';
    layer2_outputs(8731) <= b and not a;
    layer2_outputs(8732) <= b;
    layer2_outputs(8733) <= not b;
    layer2_outputs(8734) <= not b or a;
    layer2_outputs(8735) <= a xor b;
    layer2_outputs(8736) <= a;
    layer2_outputs(8737) <= b and not a;
    layer2_outputs(8738) <= not a or b;
    layer2_outputs(8739) <= not b;
    layer2_outputs(8740) <= not a;
    layer2_outputs(8741) <= not (a or b);
    layer2_outputs(8742) <= '1';
    layer2_outputs(8743) <= b;
    layer2_outputs(8744) <= not a or b;
    layer2_outputs(8745) <= '1';
    layer2_outputs(8746) <= a;
    layer2_outputs(8747) <= '0';
    layer2_outputs(8748) <= b;
    layer2_outputs(8749) <= not (a xor b);
    layer2_outputs(8750) <= '1';
    layer2_outputs(8751) <= a and b;
    layer2_outputs(8752) <= '1';
    layer2_outputs(8753) <= not (a xor b);
    layer2_outputs(8754) <= not a or b;
    layer2_outputs(8755) <= not (a and b);
    layer2_outputs(8756) <= not b or a;
    layer2_outputs(8757) <= a and not b;
    layer2_outputs(8758) <= not (a and b);
    layer2_outputs(8759) <= not a or b;
    layer2_outputs(8760) <= not b or a;
    layer2_outputs(8761) <= not b or a;
    layer2_outputs(8762) <= not (a xor b);
    layer2_outputs(8763) <= a xor b;
    layer2_outputs(8764) <= not a or b;
    layer2_outputs(8765) <= not (a or b);
    layer2_outputs(8766) <= b;
    layer2_outputs(8767) <= not b or a;
    layer2_outputs(8768) <= not a or b;
    layer2_outputs(8769) <= not (a or b);
    layer2_outputs(8770) <= a and not b;
    layer2_outputs(8771) <= a and not b;
    layer2_outputs(8772) <= a or b;
    layer2_outputs(8773) <= a and not b;
    layer2_outputs(8774) <= a and b;
    layer2_outputs(8775) <= not a;
    layer2_outputs(8776) <= a;
    layer2_outputs(8777) <= a;
    layer2_outputs(8778) <= a;
    layer2_outputs(8779) <= b;
    layer2_outputs(8780) <= not (a xor b);
    layer2_outputs(8781) <= a and b;
    layer2_outputs(8782) <= not b;
    layer2_outputs(8783) <= a and not b;
    layer2_outputs(8784) <= not b;
    layer2_outputs(8785) <= not (a xor b);
    layer2_outputs(8786) <= a;
    layer2_outputs(8787) <= b and not a;
    layer2_outputs(8788) <= not b;
    layer2_outputs(8789) <= b and not a;
    layer2_outputs(8790) <= not b or a;
    layer2_outputs(8791) <= not (a or b);
    layer2_outputs(8792) <= not b or a;
    layer2_outputs(8793) <= not b;
    layer2_outputs(8794) <= b;
    layer2_outputs(8795) <= a and not b;
    layer2_outputs(8796) <= not b;
    layer2_outputs(8797) <= a and not b;
    layer2_outputs(8798) <= not (a and b);
    layer2_outputs(8799) <= a xor b;
    layer2_outputs(8800) <= not (a xor b);
    layer2_outputs(8801) <= a or b;
    layer2_outputs(8802) <= '0';
    layer2_outputs(8803) <= not b or a;
    layer2_outputs(8804) <= a and b;
    layer2_outputs(8805) <= a and not b;
    layer2_outputs(8806) <= not (a or b);
    layer2_outputs(8807) <= a and not b;
    layer2_outputs(8808) <= a;
    layer2_outputs(8809) <= not a;
    layer2_outputs(8810) <= a or b;
    layer2_outputs(8811) <= not a or b;
    layer2_outputs(8812) <= b;
    layer2_outputs(8813) <= not b;
    layer2_outputs(8814) <= '0';
    layer2_outputs(8815) <= '1';
    layer2_outputs(8816) <= b and not a;
    layer2_outputs(8817) <= b and not a;
    layer2_outputs(8818) <= not (a or b);
    layer2_outputs(8819) <= not a;
    layer2_outputs(8820) <= not (a or b);
    layer2_outputs(8821) <= not b;
    layer2_outputs(8822) <= a or b;
    layer2_outputs(8823) <= not a;
    layer2_outputs(8824) <= a;
    layer2_outputs(8825) <= not a;
    layer2_outputs(8826) <= a or b;
    layer2_outputs(8827) <= '1';
    layer2_outputs(8828) <= '0';
    layer2_outputs(8829) <= a;
    layer2_outputs(8830) <= not a;
    layer2_outputs(8831) <= not b;
    layer2_outputs(8832) <= a xor b;
    layer2_outputs(8833) <= not (a and b);
    layer2_outputs(8834) <= not a;
    layer2_outputs(8835) <= '0';
    layer2_outputs(8836) <= not (a and b);
    layer2_outputs(8837) <= b;
    layer2_outputs(8838) <= '0';
    layer2_outputs(8839) <= '1';
    layer2_outputs(8840) <= not b;
    layer2_outputs(8841) <= not a;
    layer2_outputs(8842) <= not a or b;
    layer2_outputs(8843) <= '0';
    layer2_outputs(8844) <= not (a xor b);
    layer2_outputs(8845) <= not (a or b);
    layer2_outputs(8846) <= not b;
    layer2_outputs(8847) <= not a;
    layer2_outputs(8848) <= '1';
    layer2_outputs(8849) <= a and not b;
    layer2_outputs(8850) <= not a;
    layer2_outputs(8851) <= not b;
    layer2_outputs(8852) <= b;
    layer2_outputs(8853) <= not a;
    layer2_outputs(8854) <= '1';
    layer2_outputs(8855) <= not b or a;
    layer2_outputs(8856) <= not (a or b);
    layer2_outputs(8857) <= not a or b;
    layer2_outputs(8858) <= not b;
    layer2_outputs(8859) <= '1';
    layer2_outputs(8860) <= not b;
    layer2_outputs(8861) <= not a;
    layer2_outputs(8862) <= not b;
    layer2_outputs(8863) <= not (a or b);
    layer2_outputs(8864) <= a or b;
    layer2_outputs(8865) <= a or b;
    layer2_outputs(8866) <= not b or a;
    layer2_outputs(8867) <= a and not b;
    layer2_outputs(8868) <= a or b;
    layer2_outputs(8869) <= a;
    layer2_outputs(8870) <= '0';
    layer2_outputs(8871) <= not b;
    layer2_outputs(8872) <= b and not a;
    layer2_outputs(8873) <= a xor b;
    layer2_outputs(8874) <= not a;
    layer2_outputs(8875) <= not (a xor b);
    layer2_outputs(8876) <= b;
    layer2_outputs(8877) <= not (a xor b);
    layer2_outputs(8878) <= a and not b;
    layer2_outputs(8879) <= a or b;
    layer2_outputs(8880) <= '1';
    layer2_outputs(8881) <= not b;
    layer2_outputs(8882) <= b;
    layer2_outputs(8883) <= '0';
    layer2_outputs(8884) <= not (a or b);
    layer2_outputs(8885) <= a;
    layer2_outputs(8886) <= b;
    layer2_outputs(8887) <= b and not a;
    layer2_outputs(8888) <= a;
    layer2_outputs(8889) <= not (a xor b);
    layer2_outputs(8890) <= b and not a;
    layer2_outputs(8891) <= '0';
    layer2_outputs(8892) <= not b or a;
    layer2_outputs(8893) <= a and not b;
    layer2_outputs(8894) <= not a or b;
    layer2_outputs(8895) <= a or b;
    layer2_outputs(8896) <= not a;
    layer2_outputs(8897) <= a or b;
    layer2_outputs(8898) <= '0';
    layer2_outputs(8899) <= a;
    layer2_outputs(8900) <= not (a and b);
    layer2_outputs(8901) <= a and b;
    layer2_outputs(8902) <= '0';
    layer2_outputs(8903) <= not a;
    layer2_outputs(8904) <= not b or a;
    layer2_outputs(8905) <= a or b;
    layer2_outputs(8906) <= a and b;
    layer2_outputs(8907) <= a and not b;
    layer2_outputs(8908) <= '1';
    layer2_outputs(8909) <= a and not b;
    layer2_outputs(8910) <= a or b;
    layer2_outputs(8911) <= not a;
    layer2_outputs(8912) <= not (a or b);
    layer2_outputs(8913) <= not b or a;
    layer2_outputs(8914) <= b;
    layer2_outputs(8915) <= a;
    layer2_outputs(8916) <= a;
    layer2_outputs(8917) <= not b or a;
    layer2_outputs(8918) <= a or b;
    layer2_outputs(8919) <= '0';
    layer2_outputs(8920) <= not b;
    layer2_outputs(8921) <= a and b;
    layer2_outputs(8922) <= a and not b;
    layer2_outputs(8923) <= not b or a;
    layer2_outputs(8924) <= not a or b;
    layer2_outputs(8925) <= a or b;
    layer2_outputs(8926) <= not b;
    layer2_outputs(8927) <= not (a xor b);
    layer2_outputs(8928) <= not b or a;
    layer2_outputs(8929) <= not a;
    layer2_outputs(8930) <= a and not b;
    layer2_outputs(8931) <= not a;
    layer2_outputs(8932) <= '0';
    layer2_outputs(8933) <= not a;
    layer2_outputs(8934) <= a and not b;
    layer2_outputs(8935) <= a and b;
    layer2_outputs(8936) <= b;
    layer2_outputs(8937) <= a or b;
    layer2_outputs(8938) <= a and not b;
    layer2_outputs(8939) <= not a or b;
    layer2_outputs(8940) <= '0';
    layer2_outputs(8941) <= not b or a;
    layer2_outputs(8942) <= '0';
    layer2_outputs(8943) <= not a;
    layer2_outputs(8944) <= a and not b;
    layer2_outputs(8945) <= a or b;
    layer2_outputs(8946) <= not (a and b);
    layer2_outputs(8947) <= a and not b;
    layer2_outputs(8948) <= a and not b;
    layer2_outputs(8949) <= b;
    layer2_outputs(8950) <= not a or b;
    layer2_outputs(8951) <= not a or b;
    layer2_outputs(8952) <= '1';
    layer2_outputs(8953) <= not b;
    layer2_outputs(8954) <= a and b;
    layer2_outputs(8955) <= not a or b;
    layer2_outputs(8956) <= b and not a;
    layer2_outputs(8957) <= not b or a;
    layer2_outputs(8958) <= not a;
    layer2_outputs(8959) <= not b or a;
    layer2_outputs(8960) <= a;
    layer2_outputs(8961) <= not (a and b);
    layer2_outputs(8962) <= not a;
    layer2_outputs(8963) <= a or b;
    layer2_outputs(8964) <= not (a and b);
    layer2_outputs(8965) <= not b or a;
    layer2_outputs(8966) <= a xor b;
    layer2_outputs(8967) <= a or b;
    layer2_outputs(8968) <= '1';
    layer2_outputs(8969) <= '0';
    layer2_outputs(8970) <= a or b;
    layer2_outputs(8971) <= not b or a;
    layer2_outputs(8972) <= a or b;
    layer2_outputs(8973) <= not (a xor b);
    layer2_outputs(8974) <= '1';
    layer2_outputs(8975) <= not a or b;
    layer2_outputs(8976) <= not a or b;
    layer2_outputs(8977) <= a and b;
    layer2_outputs(8978) <= '0';
    layer2_outputs(8979) <= b and not a;
    layer2_outputs(8980) <= a and b;
    layer2_outputs(8981) <= a;
    layer2_outputs(8982) <= not a;
    layer2_outputs(8983) <= not b or a;
    layer2_outputs(8984) <= a;
    layer2_outputs(8985) <= not a;
    layer2_outputs(8986) <= not b or a;
    layer2_outputs(8987) <= a and not b;
    layer2_outputs(8988) <= not a or b;
    layer2_outputs(8989) <= '1';
    layer2_outputs(8990) <= not (a or b);
    layer2_outputs(8991) <= b and not a;
    layer2_outputs(8992) <= a xor b;
    layer2_outputs(8993) <= not (a and b);
    layer2_outputs(8994) <= b;
    layer2_outputs(8995) <= not a or b;
    layer2_outputs(8996) <= b and not a;
    layer2_outputs(8997) <= a and not b;
    layer2_outputs(8998) <= a or b;
    layer2_outputs(8999) <= a xor b;
    layer2_outputs(9000) <= a and b;
    layer2_outputs(9001) <= a and not b;
    layer2_outputs(9002) <= not (a xor b);
    layer2_outputs(9003) <= not (a xor b);
    layer2_outputs(9004) <= not b;
    layer2_outputs(9005) <= not a or b;
    layer2_outputs(9006) <= a and not b;
    layer2_outputs(9007) <= a and b;
    layer2_outputs(9008) <= not (a or b);
    layer2_outputs(9009) <= not b;
    layer2_outputs(9010) <= not b or a;
    layer2_outputs(9011) <= not (a xor b);
    layer2_outputs(9012) <= a and b;
    layer2_outputs(9013) <= b;
    layer2_outputs(9014) <= a and not b;
    layer2_outputs(9015) <= b;
    layer2_outputs(9016) <= a and b;
    layer2_outputs(9017) <= not (a xor b);
    layer2_outputs(9018) <= not a;
    layer2_outputs(9019) <= a and not b;
    layer2_outputs(9020) <= not (a or b);
    layer2_outputs(9021) <= '0';
    layer2_outputs(9022) <= not (a and b);
    layer2_outputs(9023) <= not a;
    layer2_outputs(9024) <= a;
    layer2_outputs(9025) <= not a or b;
    layer2_outputs(9026) <= not a;
    layer2_outputs(9027) <= not b or a;
    layer2_outputs(9028) <= '1';
    layer2_outputs(9029) <= '0';
    layer2_outputs(9030) <= a;
    layer2_outputs(9031) <= a xor b;
    layer2_outputs(9032) <= a xor b;
    layer2_outputs(9033) <= b and not a;
    layer2_outputs(9034) <= b;
    layer2_outputs(9035) <= not a or b;
    layer2_outputs(9036) <= b and not a;
    layer2_outputs(9037) <= not a;
    layer2_outputs(9038) <= b and not a;
    layer2_outputs(9039) <= a;
    layer2_outputs(9040) <= a xor b;
    layer2_outputs(9041) <= b and not a;
    layer2_outputs(9042) <= not (a and b);
    layer2_outputs(9043) <= not b or a;
    layer2_outputs(9044) <= b;
    layer2_outputs(9045) <= not b or a;
    layer2_outputs(9046) <= '0';
    layer2_outputs(9047) <= not b;
    layer2_outputs(9048) <= a;
    layer2_outputs(9049) <= '0';
    layer2_outputs(9050) <= b and not a;
    layer2_outputs(9051) <= a xor b;
    layer2_outputs(9052) <= not b;
    layer2_outputs(9053) <= b and not a;
    layer2_outputs(9054) <= b and not a;
    layer2_outputs(9055) <= a xor b;
    layer2_outputs(9056) <= not b;
    layer2_outputs(9057) <= a;
    layer2_outputs(9058) <= a xor b;
    layer2_outputs(9059) <= a or b;
    layer2_outputs(9060) <= a or b;
    layer2_outputs(9061) <= a or b;
    layer2_outputs(9062) <= not b or a;
    layer2_outputs(9063) <= '0';
    layer2_outputs(9064) <= not b;
    layer2_outputs(9065) <= not a;
    layer2_outputs(9066) <= not b or a;
    layer2_outputs(9067) <= a and b;
    layer2_outputs(9068) <= '1';
    layer2_outputs(9069) <= '1';
    layer2_outputs(9070) <= not b or a;
    layer2_outputs(9071) <= b;
    layer2_outputs(9072) <= '1';
    layer2_outputs(9073) <= b;
    layer2_outputs(9074) <= not b;
    layer2_outputs(9075) <= a and not b;
    layer2_outputs(9076) <= a and b;
    layer2_outputs(9077) <= not (a xor b);
    layer2_outputs(9078) <= not a;
    layer2_outputs(9079) <= not b;
    layer2_outputs(9080) <= a or b;
    layer2_outputs(9081) <= a or b;
    layer2_outputs(9082) <= b and not a;
    layer2_outputs(9083) <= not (a or b);
    layer2_outputs(9084) <= not b or a;
    layer2_outputs(9085) <= '0';
    layer2_outputs(9086) <= a;
    layer2_outputs(9087) <= not (a or b);
    layer2_outputs(9088) <= not b or a;
    layer2_outputs(9089) <= not (a and b);
    layer2_outputs(9090) <= a or b;
    layer2_outputs(9091) <= a;
    layer2_outputs(9092) <= a and b;
    layer2_outputs(9093) <= b;
    layer2_outputs(9094) <= not b;
    layer2_outputs(9095) <= not a;
    layer2_outputs(9096) <= b;
    layer2_outputs(9097) <= b and not a;
    layer2_outputs(9098) <= a and not b;
    layer2_outputs(9099) <= '0';
    layer2_outputs(9100) <= not b or a;
    layer2_outputs(9101) <= not a or b;
    layer2_outputs(9102) <= '0';
    layer2_outputs(9103) <= not a;
    layer2_outputs(9104) <= a xor b;
    layer2_outputs(9105) <= b and not a;
    layer2_outputs(9106) <= '0';
    layer2_outputs(9107) <= a;
    layer2_outputs(9108) <= not (a or b);
    layer2_outputs(9109) <= a;
    layer2_outputs(9110) <= a xor b;
    layer2_outputs(9111) <= a or b;
    layer2_outputs(9112) <= a;
    layer2_outputs(9113) <= a and b;
    layer2_outputs(9114) <= not a or b;
    layer2_outputs(9115) <= not a or b;
    layer2_outputs(9116) <= a and not b;
    layer2_outputs(9117) <= a xor b;
    layer2_outputs(9118) <= not a;
    layer2_outputs(9119) <= not a;
    layer2_outputs(9120) <= b;
    layer2_outputs(9121) <= b;
    layer2_outputs(9122) <= a and not b;
    layer2_outputs(9123) <= not a;
    layer2_outputs(9124) <= '1';
    layer2_outputs(9125) <= a or b;
    layer2_outputs(9126) <= '1';
    layer2_outputs(9127) <= a and not b;
    layer2_outputs(9128) <= b;
    layer2_outputs(9129) <= a or b;
    layer2_outputs(9130) <= a and not b;
    layer2_outputs(9131) <= '0';
    layer2_outputs(9132) <= not b;
    layer2_outputs(9133) <= a;
    layer2_outputs(9134) <= not a;
    layer2_outputs(9135) <= a or b;
    layer2_outputs(9136) <= b;
    layer2_outputs(9137) <= not a;
    layer2_outputs(9138) <= not (a and b);
    layer2_outputs(9139) <= b and not a;
    layer2_outputs(9140) <= a;
    layer2_outputs(9141) <= a xor b;
    layer2_outputs(9142) <= not a or b;
    layer2_outputs(9143) <= a or b;
    layer2_outputs(9144) <= b;
    layer2_outputs(9145) <= a;
    layer2_outputs(9146) <= b;
    layer2_outputs(9147) <= '0';
    layer2_outputs(9148) <= b;
    layer2_outputs(9149) <= not (a xor b);
    layer2_outputs(9150) <= '1';
    layer2_outputs(9151) <= a or b;
    layer2_outputs(9152) <= not a or b;
    layer2_outputs(9153) <= not b or a;
    layer2_outputs(9154) <= not (a or b);
    layer2_outputs(9155) <= not a;
    layer2_outputs(9156) <= a xor b;
    layer2_outputs(9157) <= b and not a;
    layer2_outputs(9158) <= not b;
    layer2_outputs(9159) <= a and not b;
    layer2_outputs(9160) <= a and not b;
    layer2_outputs(9161) <= not b or a;
    layer2_outputs(9162) <= '1';
    layer2_outputs(9163) <= not a or b;
    layer2_outputs(9164) <= a and not b;
    layer2_outputs(9165) <= not a;
    layer2_outputs(9166) <= not b;
    layer2_outputs(9167) <= not a or b;
    layer2_outputs(9168) <= '0';
    layer2_outputs(9169) <= not a or b;
    layer2_outputs(9170) <= '1';
    layer2_outputs(9171) <= a;
    layer2_outputs(9172) <= '1';
    layer2_outputs(9173) <= b;
    layer2_outputs(9174) <= not a;
    layer2_outputs(9175) <= not (a or b);
    layer2_outputs(9176) <= '1';
    layer2_outputs(9177) <= a and b;
    layer2_outputs(9178) <= a and not b;
    layer2_outputs(9179) <= not b;
    layer2_outputs(9180) <= a xor b;
    layer2_outputs(9181) <= a and not b;
    layer2_outputs(9182) <= not a;
    layer2_outputs(9183) <= not a;
    layer2_outputs(9184) <= a or b;
    layer2_outputs(9185) <= not (a or b);
    layer2_outputs(9186) <= not b or a;
    layer2_outputs(9187) <= a and not b;
    layer2_outputs(9188) <= a;
    layer2_outputs(9189) <= a;
    layer2_outputs(9190) <= b;
    layer2_outputs(9191) <= '0';
    layer2_outputs(9192) <= not b or a;
    layer2_outputs(9193) <= not (a and b);
    layer2_outputs(9194) <= not a;
    layer2_outputs(9195) <= not a;
    layer2_outputs(9196) <= not a or b;
    layer2_outputs(9197) <= a and not b;
    layer2_outputs(9198) <= b and not a;
    layer2_outputs(9199) <= '0';
    layer2_outputs(9200) <= not b;
    layer2_outputs(9201) <= not (a or b);
    layer2_outputs(9202) <= b;
    layer2_outputs(9203) <= b and not a;
    layer2_outputs(9204) <= a or b;
    layer2_outputs(9205) <= not a;
    layer2_outputs(9206) <= not a or b;
    layer2_outputs(9207) <= not b or a;
    layer2_outputs(9208) <= a xor b;
    layer2_outputs(9209) <= not a or b;
    layer2_outputs(9210) <= a or b;
    layer2_outputs(9211) <= '1';
    layer2_outputs(9212) <= a and not b;
    layer2_outputs(9213) <= not (a or b);
    layer2_outputs(9214) <= not b;
    layer2_outputs(9215) <= not b;
    layer2_outputs(9216) <= b and not a;
    layer2_outputs(9217) <= a or b;
    layer2_outputs(9218) <= not b;
    layer2_outputs(9219) <= not (a xor b);
    layer2_outputs(9220) <= not b;
    layer2_outputs(9221) <= not b;
    layer2_outputs(9222) <= a and not b;
    layer2_outputs(9223) <= not (a xor b);
    layer2_outputs(9224) <= not b or a;
    layer2_outputs(9225) <= not b;
    layer2_outputs(9226) <= a or b;
    layer2_outputs(9227) <= not a or b;
    layer2_outputs(9228) <= b;
    layer2_outputs(9229) <= a or b;
    layer2_outputs(9230) <= not b;
    layer2_outputs(9231) <= b and not a;
    layer2_outputs(9232) <= a and not b;
    layer2_outputs(9233) <= b and not a;
    layer2_outputs(9234) <= not a;
    layer2_outputs(9235) <= not (a or b);
    layer2_outputs(9236) <= a;
    layer2_outputs(9237) <= not (a and b);
    layer2_outputs(9238) <= b and not a;
    layer2_outputs(9239) <= a;
    layer2_outputs(9240) <= not a;
    layer2_outputs(9241) <= b;
    layer2_outputs(9242) <= a or b;
    layer2_outputs(9243) <= '0';
    layer2_outputs(9244) <= a and b;
    layer2_outputs(9245) <= not a;
    layer2_outputs(9246) <= '0';
    layer2_outputs(9247) <= a;
    layer2_outputs(9248) <= not (a or b);
    layer2_outputs(9249) <= not b;
    layer2_outputs(9250) <= a and b;
    layer2_outputs(9251) <= not (a or b);
    layer2_outputs(9252) <= not a or b;
    layer2_outputs(9253) <= a and b;
    layer2_outputs(9254) <= a or b;
    layer2_outputs(9255) <= b;
    layer2_outputs(9256) <= b and not a;
    layer2_outputs(9257) <= not a;
    layer2_outputs(9258) <= '1';
    layer2_outputs(9259) <= b and not a;
    layer2_outputs(9260) <= a and not b;
    layer2_outputs(9261) <= b;
    layer2_outputs(9262) <= not (a xor b);
    layer2_outputs(9263) <= not a;
    layer2_outputs(9264) <= not a;
    layer2_outputs(9265) <= '0';
    layer2_outputs(9266) <= a and not b;
    layer2_outputs(9267) <= not a;
    layer2_outputs(9268) <= not (a xor b);
    layer2_outputs(9269) <= not (a or b);
    layer2_outputs(9270) <= a;
    layer2_outputs(9271) <= not (a and b);
    layer2_outputs(9272) <= a and b;
    layer2_outputs(9273) <= a;
    layer2_outputs(9274) <= not b or a;
    layer2_outputs(9275) <= not a;
    layer2_outputs(9276) <= a xor b;
    layer2_outputs(9277) <= not a or b;
    layer2_outputs(9278) <= a;
    layer2_outputs(9279) <= not a or b;
    layer2_outputs(9280) <= not b or a;
    layer2_outputs(9281) <= not b or a;
    layer2_outputs(9282) <= not a;
    layer2_outputs(9283) <= '0';
    layer2_outputs(9284) <= not b;
    layer2_outputs(9285) <= a and b;
    layer2_outputs(9286) <= '0';
    layer2_outputs(9287) <= not (a and b);
    layer2_outputs(9288) <= not b;
    layer2_outputs(9289) <= not (a and b);
    layer2_outputs(9290) <= not b or a;
    layer2_outputs(9291) <= b and not a;
    layer2_outputs(9292) <= not a;
    layer2_outputs(9293) <= not a or b;
    layer2_outputs(9294) <= not a or b;
    layer2_outputs(9295) <= '0';
    layer2_outputs(9296) <= b;
    layer2_outputs(9297) <= not (a or b);
    layer2_outputs(9298) <= '0';
    layer2_outputs(9299) <= not (a or b);
    layer2_outputs(9300) <= not b;
    layer2_outputs(9301) <= a;
    layer2_outputs(9302) <= not b or a;
    layer2_outputs(9303) <= b;
    layer2_outputs(9304) <= a xor b;
    layer2_outputs(9305) <= a or b;
    layer2_outputs(9306) <= '1';
    layer2_outputs(9307) <= not b or a;
    layer2_outputs(9308) <= a and not b;
    layer2_outputs(9309) <= b;
    layer2_outputs(9310) <= not (a or b);
    layer2_outputs(9311) <= '0';
    layer2_outputs(9312) <= a or b;
    layer2_outputs(9313) <= '0';
    layer2_outputs(9314) <= not (a or b);
    layer2_outputs(9315) <= b and not a;
    layer2_outputs(9316) <= not (a xor b);
    layer2_outputs(9317) <= '1';
    layer2_outputs(9318) <= '1';
    layer2_outputs(9319) <= not (a or b);
    layer2_outputs(9320) <= not b or a;
    layer2_outputs(9321) <= not a;
    layer2_outputs(9322) <= not a;
    layer2_outputs(9323) <= a xor b;
    layer2_outputs(9324) <= b and not a;
    layer2_outputs(9325) <= not b or a;
    layer2_outputs(9326) <= b and not a;
    layer2_outputs(9327) <= not a;
    layer2_outputs(9328) <= not a or b;
    layer2_outputs(9329) <= not (a and b);
    layer2_outputs(9330) <= a;
    layer2_outputs(9331) <= not b;
    layer2_outputs(9332) <= b and not a;
    layer2_outputs(9333) <= not (a xor b);
    layer2_outputs(9334) <= not b;
    layer2_outputs(9335) <= not a or b;
    layer2_outputs(9336) <= a xor b;
    layer2_outputs(9337) <= not (a or b);
    layer2_outputs(9338) <= '0';
    layer2_outputs(9339) <= a or b;
    layer2_outputs(9340) <= b and not a;
    layer2_outputs(9341) <= '0';
    layer2_outputs(9342) <= b;
    layer2_outputs(9343) <= b;
    layer2_outputs(9344) <= a and b;
    layer2_outputs(9345) <= not b;
    layer2_outputs(9346) <= not b or a;
    layer2_outputs(9347) <= '1';
    layer2_outputs(9348) <= not (a and b);
    layer2_outputs(9349) <= a;
    layer2_outputs(9350) <= not b;
    layer2_outputs(9351) <= not b;
    layer2_outputs(9352) <= not (a xor b);
    layer2_outputs(9353) <= b and not a;
    layer2_outputs(9354) <= '1';
    layer2_outputs(9355) <= not a;
    layer2_outputs(9356) <= a and not b;
    layer2_outputs(9357) <= b and not a;
    layer2_outputs(9358) <= not a;
    layer2_outputs(9359) <= a;
    layer2_outputs(9360) <= a and not b;
    layer2_outputs(9361) <= b and not a;
    layer2_outputs(9362) <= a and not b;
    layer2_outputs(9363) <= b;
    layer2_outputs(9364) <= not a;
    layer2_outputs(9365) <= b and not a;
    layer2_outputs(9366) <= not b;
    layer2_outputs(9367) <= b;
    layer2_outputs(9368) <= b;
    layer2_outputs(9369) <= a;
    layer2_outputs(9370) <= not (a and b);
    layer2_outputs(9371) <= a and not b;
    layer2_outputs(9372) <= b;
    layer2_outputs(9373) <= a;
    layer2_outputs(9374) <= a and not b;
    layer2_outputs(9375) <= b;
    layer2_outputs(9376) <= not (a and b);
    layer2_outputs(9377) <= not b or a;
    layer2_outputs(9378) <= a or b;
    layer2_outputs(9379) <= not b or a;
    layer2_outputs(9380) <= b and not a;
    layer2_outputs(9381) <= b;
    layer2_outputs(9382) <= a and b;
    layer2_outputs(9383) <= not b;
    layer2_outputs(9384) <= a and b;
    layer2_outputs(9385) <= not a or b;
    layer2_outputs(9386) <= not b;
    layer2_outputs(9387) <= a;
    layer2_outputs(9388) <= a or b;
    layer2_outputs(9389) <= not (a or b);
    layer2_outputs(9390) <= b;
    layer2_outputs(9391) <= not a;
    layer2_outputs(9392) <= a;
    layer2_outputs(9393) <= a and b;
    layer2_outputs(9394) <= not (a or b);
    layer2_outputs(9395) <= b;
    layer2_outputs(9396) <= a or b;
    layer2_outputs(9397) <= not b or a;
    layer2_outputs(9398) <= not a;
    layer2_outputs(9399) <= not a;
    layer2_outputs(9400) <= not (a and b);
    layer2_outputs(9401) <= b;
    layer2_outputs(9402) <= '1';
    layer2_outputs(9403) <= a xor b;
    layer2_outputs(9404) <= a;
    layer2_outputs(9405) <= '0';
    layer2_outputs(9406) <= b;
    layer2_outputs(9407) <= a and not b;
    layer2_outputs(9408) <= a and not b;
    layer2_outputs(9409) <= a or b;
    layer2_outputs(9410) <= a;
    layer2_outputs(9411) <= a or b;
    layer2_outputs(9412) <= not b or a;
    layer2_outputs(9413) <= not (a or b);
    layer2_outputs(9414) <= not (a xor b);
    layer2_outputs(9415) <= not b or a;
    layer2_outputs(9416) <= '0';
    layer2_outputs(9417) <= not b or a;
    layer2_outputs(9418) <= a;
    layer2_outputs(9419) <= not (a and b);
    layer2_outputs(9420) <= a;
    layer2_outputs(9421) <= not a or b;
    layer2_outputs(9422) <= not (a xor b);
    layer2_outputs(9423) <= b;
    layer2_outputs(9424) <= not b;
    layer2_outputs(9425) <= '1';
    layer2_outputs(9426) <= a xor b;
    layer2_outputs(9427) <= a and b;
    layer2_outputs(9428) <= '0';
    layer2_outputs(9429) <= not a or b;
    layer2_outputs(9430) <= not a;
    layer2_outputs(9431) <= b and not a;
    layer2_outputs(9432) <= not (a xor b);
    layer2_outputs(9433) <= b;
    layer2_outputs(9434) <= not b;
    layer2_outputs(9435) <= not (a xor b);
    layer2_outputs(9436) <= '1';
    layer2_outputs(9437) <= not (a or b);
    layer2_outputs(9438) <= a;
    layer2_outputs(9439) <= a xor b;
    layer2_outputs(9440) <= a and not b;
    layer2_outputs(9441) <= not (a xor b);
    layer2_outputs(9442) <= not a;
    layer2_outputs(9443) <= a;
    layer2_outputs(9444) <= b;
    layer2_outputs(9445) <= not a;
    layer2_outputs(9446) <= a and b;
    layer2_outputs(9447) <= a xor b;
    layer2_outputs(9448) <= a xor b;
    layer2_outputs(9449) <= not b or a;
    layer2_outputs(9450) <= not a;
    layer2_outputs(9451) <= b and not a;
    layer2_outputs(9452) <= not (a or b);
    layer2_outputs(9453) <= '0';
    layer2_outputs(9454) <= not b or a;
    layer2_outputs(9455) <= not (a xor b);
    layer2_outputs(9456) <= not (a xor b);
    layer2_outputs(9457) <= a or b;
    layer2_outputs(9458) <= a;
    layer2_outputs(9459) <= not (a or b);
    layer2_outputs(9460) <= a;
    layer2_outputs(9461) <= not b;
    layer2_outputs(9462) <= a;
    layer2_outputs(9463) <= b;
    layer2_outputs(9464) <= a;
    layer2_outputs(9465) <= not b;
    layer2_outputs(9466) <= not b;
    layer2_outputs(9467) <= not b;
    layer2_outputs(9468) <= not a or b;
    layer2_outputs(9469) <= a;
    layer2_outputs(9470) <= b and not a;
    layer2_outputs(9471) <= b;
    layer2_outputs(9472) <= not a;
    layer2_outputs(9473) <= b;
    layer2_outputs(9474) <= b and not a;
    layer2_outputs(9475) <= not b or a;
    layer2_outputs(9476) <= not b;
    layer2_outputs(9477) <= '0';
    layer2_outputs(9478) <= '0';
    layer2_outputs(9479) <= not a or b;
    layer2_outputs(9480) <= a;
    layer2_outputs(9481) <= '1';
    layer2_outputs(9482) <= not a or b;
    layer2_outputs(9483) <= not a;
    layer2_outputs(9484) <= a or b;
    layer2_outputs(9485) <= not b;
    layer2_outputs(9486) <= a and not b;
    layer2_outputs(9487) <= b and not a;
    layer2_outputs(9488) <= not a;
    layer2_outputs(9489) <= '0';
    layer2_outputs(9490) <= a and b;
    layer2_outputs(9491) <= '1';
    layer2_outputs(9492) <= a and not b;
    layer2_outputs(9493) <= not b;
    layer2_outputs(9494) <= not (a and b);
    layer2_outputs(9495) <= a;
    layer2_outputs(9496) <= b;
    layer2_outputs(9497) <= a and b;
    layer2_outputs(9498) <= '1';
    layer2_outputs(9499) <= not (a or b);
    layer2_outputs(9500) <= a or b;
    layer2_outputs(9501) <= a and b;
    layer2_outputs(9502) <= a and not b;
    layer2_outputs(9503) <= '0';
    layer2_outputs(9504) <= b;
    layer2_outputs(9505) <= a and not b;
    layer2_outputs(9506) <= b and not a;
    layer2_outputs(9507) <= not b or a;
    layer2_outputs(9508) <= '1';
    layer2_outputs(9509) <= not a or b;
    layer2_outputs(9510) <= a;
    layer2_outputs(9511) <= a;
    layer2_outputs(9512) <= not (a and b);
    layer2_outputs(9513) <= '1';
    layer2_outputs(9514) <= a;
    layer2_outputs(9515) <= a;
    layer2_outputs(9516) <= not a;
    layer2_outputs(9517) <= not a or b;
    layer2_outputs(9518) <= not b;
    layer2_outputs(9519) <= not b or a;
    layer2_outputs(9520) <= not (a xor b);
    layer2_outputs(9521) <= not (a xor b);
    layer2_outputs(9522) <= not a or b;
    layer2_outputs(9523) <= a or b;
    layer2_outputs(9524) <= a;
    layer2_outputs(9525) <= not b or a;
    layer2_outputs(9526) <= a xor b;
    layer2_outputs(9527) <= not (a and b);
    layer2_outputs(9528) <= b;
    layer2_outputs(9529) <= a and not b;
    layer2_outputs(9530) <= b;
    layer2_outputs(9531) <= b and not a;
    layer2_outputs(9532) <= b and not a;
    layer2_outputs(9533) <= not (a or b);
    layer2_outputs(9534) <= b and not a;
    layer2_outputs(9535) <= not a;
    layer2_outputs(9536) <= a and b;
    layer2_outputs(9537) <= '0';
    layer2_outputs(9538) <= not (a xor b);
    layer2_outputs(9539) <= not (a and b);
    layer2_outputs(9540) <= a;
    layer2_outputs(9541) <= a or b;
    layer2_outputs(9542) <= '1';
    layer2_outputs(9543) <= not (a and b);
    layer2_outputs(9544) <= not (a and b);
    layer2_outputs(9545) <= a;
    layer2_outputs(9546) <= not a or b;
    layer2_outputs(9547) <= b;
    layer2_outputs(9548) <= not a or b;
    layer2_outputs(9549) <= not b;
    layer2_outputs(9550) <= a and not b;
    layer2_outputs(9551) <= a and not b;
    layer2_outputs(9552) <= not (a and b);
    layer2_outputs(9553) <= '1';
    layer2_outputs(9554) <= b;
    layer2_outputs(9555) <= a or b;
    layer2_outputs(9556) <= not a or b;
    layer2_outputs(9557) <= not a or b;
    layer2_outputs(9558) <= not a or b;
    layer2_outputs(9559) <= not b;
    layer2_outputs(9560) <= a xor b;
    layer2_outputs(9561) <= not a;
    layer2_outputs(9562) <= not a or b;
    layer2_outputs(9563) <= b;
    layer2_outputs(9564) <= not a or b;
    layer2_outputs(9565) <= not b or a;
    layer2_outputs(9566) <= a;
    layer2_outputs(9567) <= a and b;
    layer2_outputs(9568) <= not a or b;
    layer2_outputs(9569) <= b;
    layer2_outputs(9570) <= not (a or b);
    layer2_outputs(9571) <= '0';
    layer2_outputs(9572) <= b;
    layer2_outputs(9573) <= not (a xor b);
    layer2_outputs(9574) <= b and not a;
    layer2_outputs(9575) <= b and not a;
    layer2_outputs(9576) <= a and b;
    layer2_outputs(9577) <= '1';
    layer2_outputs(9578) <= a and b;
    layer2_outputs(9579) <= not b;
    layer2_outputs(9580) <= not (a or b);
    layer2_outputs(9581) <= not b;
    layer2_outputs(9582) <= b and not a;
    layer2_outputs(9583) <= not (a xor b);
    layer2_outputs(9584) <= '0';
    layer2_outputs(9585) <= not a or b;
    layer2_outputs(9586) <= b;
    layer2_outputs(9587) <= not (a xor b);
    layer2_outputs(9588) <= a and not b;
    layer2_outputs(9589) <= not (a or b);
    layer2_outputs(9590) <= '0';
    layer2_outputs(9591) <= not b;
    layer2_outputs(9592) <= not a;
    layer2_outputs(9593) <= not a;
    layer2_outputs(9594) <= not b;
    layer2_outputs(9595) <= a and b;
    layer2_outputs(9596) <= '1';
    layer2_outputs(9597) <= a;
    layer2_outputs(9598) <= a and b;
    layer2_outputs(9599) <= a;
    layer2_outputs(9600) <= not (a and b);
    layer2_outputs(9601) <= a or b;
    layer2_outputs(9602) <= not a;
    layer2_outputs(9603) <= not a or b;
    layer2_outputs(9604) <= not a;
    layer2_outputs(9605) <= a xor b;
    layer2_outputs(9606) <= '0';
    layer2_outputs(9607) <= not b;
    layer2_outputs(9608) <= a;
    layer2_outputs(9609) <= b and not a;
    layer2_outputs(9610) <= a and b;
    layer2_outputs(9611) <= not a;
    layer2_outputs(9612) <= not a;
    layer2_outputs(9613) <= a;
    layer2_outputs(9614) <= b;
    layer2_outputs(9615) <= not (a or b);
    layer2_outputs(9616) <= not b or a;
    layer2_outputs(9617) <= not b;
    layer2_outputs(9618) <= a;
    layer2_outputs(9619) <= not (a and b);
    layer2_outputs(9620) <= a;
    layer2_outputs(9621) <= b;
    layer2_outputs(9622) <= a;
    layer2_outputs(9623) <= b;
    layer2_outputs(9624) <= not (a or b);
    layer2_outputs(9625) <= not (a and b);
    layer2_outputs(9626) <= b and not a;
    layer2_outputs(9627) <= not (a or b);
    layer2_outputs(9628) <= not (a and b);
    layer2_outputs(9629) <= '0';
    layer2_outputs(9630) <= not (a or b);
    layer2_outputs(9631) <= not b or a;
    layer2_outputs(9632) <= a;
    layer2_outputs(9633) <= a and not b;
    layer2_outputs(9634) <= not (a or b);
    layer2_outputs(9635) <= b and not a;
    layer2_outputs(9636) <= '1';
    layer2_outputs(9637) <= b;
    layer2_outputs(9638) <= a;
    layer2_outputs(9639) <= a and b;
    layer2_outputs(9640) <= a and b;
    layer2_outputs(9641) <= a;
    layer2_outputs(9642) <= b;
    layer2_outputs(9643) <= '0';
    layer2_outputs(9644) <= not a;
    layer2_outputs(9645) <= b;
    layer2_outputs(9646) <= b and not a;
    layer2_outputs(9647) <= not b or a;
    layer2_outputs(9648) <= a or b;
    layer2_outputs(9649) <= not a;
    layer2_outputs(9650) <= b;
    layer2_outputs(9651) <= not a;
    layer2_outputs(9652) <= not b;
    layer2_outputs(9653) <= not b;
    layer2_outputs(9654) <= '0';
    layer2_outputs(9655) <= not (a or b);
    layer2_outputs(9656) <= b;
    layer2_outputs(9657) <= not (a and b);
    layer2_outputs(9658) <= a;
    layer2_outputs(9659) <= a and not b;
    layer2_outputs(9660) <= b;
    layer2_outputs(9661) <= not a;
    layer2_outputs(9662) <= a or b;
    layer2_outputs(9663) <= a and b;
    layer2_outputs(9664) <= a and not b;
    layer2_outputs(9665) <= not (a and b);
    layer2_outputs(9666) <= b and not a;
    layer2_outputs(9667) <= '0';
    layer2_outputs(9668) <= a xor b;
    layer2_outputs(9669) <= '0';
    layer2_outputs(9670) <= '0';
    layer2_outputs(9671) <= b;
    layer2_outputs(9672) <= a and b;
    layer2_outputs(9673) <= a xor b;
    layer2_outputs(9674) <= not (a or b);
    layer2_outputs(9675) <= b and not a;
    layer2_outputs(9676) <= a and b;
    layer2_outputs(9677) <= not a or b;
    layer2_outputs(9678) <= a;
    layer2_outputs(9679) <= not (a and b);
    layer2_outputs(9680) <= b;
    layer2_outputs(9681) <= not a or b;
    layer2_outputs(9682) <= b;
    layer2_outputs(9683) <= a;
    layer2_outputs(9684) <= not (a and b);
    layer2_outputs(9685) <= b and not a;
    layer2_outputs(9686) <= b and not a;
    layer2_outputs(9687) <= not (a xor b);
    layer2_outputs(9688) <= a and b;
    layer2_outputs(9689) <= not a;
    layer2_outputs(9690) <= not b or a;
    layer2_outputs(9691) <= not a;
    layer2_outputs(9692) <= b;
    layer2_outputs(9693) <= not (a and b);
    layer2_outputs(9694) <= a and b;
    layer2_outputs(9695) <= a;
    layer2_outputs(9696) <= a;
    layer2_outputs(9697) <= '1';
    layer2_outputs(9698) <= a;
    layer2_outputs(9699) <= b;
    layer2_outputs(9700) <= '0';
    layer2_outputs(9701) <= b and not a;
    layer2_outputs(9702) <= a;
    layer2_outputs(9703) <= a and b;
    layer2_outputs(9704) <= not (a xor b);
    layer2_outputs(9705) <= b;
    layer2_outputs(9706) <= not a;
    layer2_outputs(9707) <= '0';
    layer2_outputs(9708) <= '0';
    layer2_outputs(9709) <= a;
    layer2_outputs(9710) <= not b;
    layer2_outputs(9711) <= not b;
    layer2_outputs(9712) <= not b;
    layer2_outputs(9713) <= a;
    layer2_outputs(9714) <= a and not b;
    layer2_outputs(9715) <= not b or a;
    layer2_outputs(9716) <= not b;
    layer2_outputs(9717) <= not a;
    layer2_outputs(9718) <= not (a or b);
    layer2_outputs(9719) <= not (a and b);
    layer2_outputs(9720) <= not a or b;
    layer2_outputs(9721) <= a and b;
    layer2_outputs(9722) <= a or b;
    layer2_outputs(9723) <= b;
    layer2_outputs(9724) <= not a or b;
    layer2_outputs(9725) <= not b;
    layer2_outputs(9726) <= not (a and b);
    layer2_outputs(9727) <= '0';
    layer2_outputs(9728) <= b;
    layer2_outputs(9729) <= not b or a;
    layer2_outputs(9730) <= not b;
    layer2_outputs(9731) <= a;
    layer2_outputs(9732) <= not a;
    layer2_outputs(9733) <= not b;
    layer2_outputs(9734) <= not (a and b);
    layer2_outputs(9735) <= a and not b;
    layer2_outputs(9736) <= not b;
    layer2_outputs(9737) <= b and not a;
    layer2_outputs(9738) <= not (a or b);
    layer2_outputs(9739) <= b and not a;
    layer2_outputs(9740) <= not (a or b);
    layer2_outputs(9741) <= a and b;
    layer2_outputs(9742) <= '1';
    layer2_outputs(9743) <= not a or b;
    layer2_outputs(9744) <= '0';
    layer2_outputs(9745) <= not b or a;
    layer2_outputs(9746) <= b;
    layer2_outputs(9747) <= '1';
    layer2_outputs(9748) <= '0';
    layer2_outputs(9749) <= not b;
    layer2_outputs(9750) <= a and b;
    layer2_outputs(9751) <= a and not b;
    layer2_outputs(9752) <= not (a or b);
    layer2_outputs(9753) <= not a or b;
    layer2_outputs(9754) <= a;
    layer2_outputs(9755) <= a and not b;
    layer2_outputs(9756) <= '1';
    layer2_outputs(9757) <= not a;
    layer2_outputs(9758) <= b and not a;
    layer2_outputs(9759) <= b and not a;
    layer2_outputs(9760) <= a and not b;
    layer2_outputs(9761) <= not b or a;
    layer2_outputs(9762) <= a and b;
    layer2_outputs(9763) <= not a;
    layer2_outputs(9764) <= not a or b;
    layer2_outputs(9765) <= '1';
    layer2_outputs(9766) <= a;
    layer2_outputs(9767) <= not (a and b);
    layer2_outputs(9768) <= not (a and b);
    layer2_outputs(9769) <= a xor b;
    layer2_outputs(9770) <= not (a and b);
    layer2_outputs(9771) <= not b;
    layer2_outputs(9772) <= a and b;
    layer2_outputs(9773) <= not (a and b);
    layer2_outputs(9774) <= a and not b;
    layer2_outputs(9775) <= not b;
    layer2_outputs(9776) <= not b or a;
    layer2_outputs(9777) <= '0';
    layer2_outputs(9778) <= a and not b;
    layer2_outputs(9779) <= not (a or b);
    layer2_outputs(9780) <= b;
    layer2_outputs(9781) <= '1';
    layer2_outputs(9782) <= '1';
    layer2_outputs(9783) <= not (a or b);
    layer2_outputs(9784) <= b;
    layer2_outputs(9785) <= a or b;
    layer2_outputs(9786) <= not a or b;
    layer2_outputs(9787) <= a;
    layer2_outputs(9788) <= b;
    layer2_outputs(9789) <= not (a and b);
    layer2_outputs(9790) <= not (a or b);
    layer2_outputs(9791) <= '0';
    layer2_outputs(9792) <= a or b;
    layer2_outputs(9793) <= not a;
    layer2_outputs(9794) <= '0';
    layer2_outputs(9795) <= a xor b;
    layer2_outputs(9796) <= not a;
    layer2_outputs(9797) <= not (a xor b);
    layer2_outputs(9798) <= not (a xor b);
    layer2_outputs(9799) <= a or b;
    layer2_outputs(9800) <= a and b;
    layer2_outputs(9801) <= not b or a;
    layer2_outputs(9802) <= not a or b;
    layer2_outputs(9803) <= not b;
    layer2_outputs(9804) <= not (a and b);
    layer2_outputs(9805) <= not a or b;
    layer2_outputs(9806) <= not b or a;
    layer2_outputs(9807) <= a and not b;
    layer2_outputs(9808) <= '1';
    layer2_outputs(9809) <= b;
    layer2_outputs(9810) <= not b or a;
    layer2_outputs(9811) <= b and not a;
    layer2_outputs(9812) <= '1';
    layer2_outputs(9813) <= not b or a;
    layer2_outputs(9814) <= not a;
    layer2_outputs(9815) <= a;
    layer2_outputs(9816) <= a and b;
    layer2_outputs(9817) <= not (a and b);
    layer2_outputs(9818) <= not (a or b);
    layer2_outputs(9819) <= b and not a;
    layer2_outputs(9820) <= not b;
    layer2_outputs(9821) <= not (a xor b);
    layer2_outputs(9822) <= a or b;
    layer2_outputs(9823) <= b and not a;
    layer2_outputs(9824) <= b;
    layer2_outputs(9825) <= not b or a;
    layer2_outputs(9826) <= not b;
    layer2_outputs(9827) <= '0';
    layer2_outputs(9828) <= not a or b;
    layer2_outputs(9829) <= '0';
    layer2_outputs(9830) <= b and not a;
    layer2_outputs(9831) <= not b or a;
    layer2_outputs(9832) <= not b;
    layer2_outputs(9833) <= not b or a;
    layer2_outputs(9834) <= a and b;
    layer2_outputs(9835) <= not (a or b);
    layer2_outputs(9836) <= not b or a;
    layer2_outputs(9837) <= not a or b;
    layer2_outputs(9838) <= not b or a;
    layer2_outputs(9839) <= a;
    layer2_outputs(9840) <= a and not b;
    layer2_outputs(9841) <= '0';
    layer2_outputs(9842) <= not b;
    layer2_outputs(9843) <= a and b;
    layer2_outputs(9844) <= '1';
    layer2_outputs(9845) <= not b or a;
    layer2_outputs(9846) <= a and b;
    layer2_outputs(9847) <= a or b;
    layer2_outputs(9848) <= b;
    layer2_outputs(9849) <= b;
    layer2_outputs(9850) <= not b;
    layer2_outputs(9851) <= a and not b;
    layer2_outputs(9852) <= b;
    layer2_outputs(9853) <= not a or b;
    layer2_outputs(9854) <= a and b;
    layer2_outputs(9855) <= not b;
    layer2_outputs(9856) <= not (a or b);
    layer2_outputs(9857) <= '0';
    layer2_outputs(9858) <= not (a and b);
    layer2_outputs(9859) <= not b;
    layer2_outputs(9860) <= not b;
    layer2_outputs(9861) <= b and not a;
    layer2_outputs(9862) <= a and b;
    layer2_outputs(9863) <= not a or b;
    layer2_outputs(9864) <= b;
    layer2_outputs(9865) <= not b;
    layer2_outputs(9866) <= not (a and b);
    layer2_outputs(9867) <= a;
    layer2_outputs(9868) <= not (a and b);
    layer2_outputs(9869) <= a xor b;
    layer2_outputs(9870) <= '1';
    layer2_outputs(9871) <= a xor b;
    layer2_outputs(9872) <= not b;
    layer2_outputs(9873) <= not a;
    layer2_outputs(9874) <= b and not a;
    layer2_outputs(9875) <= not b;
    layer2_outputs(9876) <= b;
    layer2_outputs(9877) <= not b;
    layer2_outputs(9878) <= a xor b;
    layer2_outputs(9879) <= a and b;
    layer2_outputs(9880) <= a or b;
    layer2_outputs(9881) <= not (a xor b);
    layer2_outputs(9882) <= b;
    layer2_outputs(9883) <= a;
    layer2_outputs(9884) <= not b;
    layer2_outputs(9885) <= not (a and b);
    layer2_outputs(9886) <= '1';
    layer2_outputs(9887) <= not a or b;
    layer2_outputs(9888) <= b and not a;
    layer2_outputs(9889) <= not (a and b);
    layer2_outputs(9890) <= a or b;
    layer2_outputs(9891) <= not a or b;
    layer2_outputs(9892) <= a and b;
    layer2_outputs(9893) <= not b;
    layer2_outputs(9894) <= not b;
    layer2_outputs(9895) <= '1';
    layer2_outputs(9896) <= not (a or b);
    layer2_outputs(9897) <= not a or b;
    layer2_outputs(9898) <= a xor b;
    layer2_outputs(9899) <= not (a and b);
    layer2_outputs(9900) <= b and not a;
    layer2_outputs(9901) <= not a or b;
    layer2_outputs(9902) <= not a;
    layer2_outputs(9903) <= b;
    layer2_outputs(9904) <= a and not b;
    layer2_outputs(9905) <= b and not a;
    layer2_outputs(9906) <= not (a xor b);
    layer2_outputs(9907) <= b;
    layer2_outputs(9908) <= a and b;
    layer2_outputs(9909) <= b;
    layer2_outputs(9910) <= '1';
    layer2_outputs(9911) <= not (a and b);
    layer2_outputs(9912) <= not a;
    layer2_outputs(9913) <= not b or a;
    layer2_outputs(9914) <= a and not b;
    layer2_outputs(9915) <= not (a or b);
    layer2_outputs(9916) <= a;
    layer2_outputs(9917) <= not a;
    layer2_outputs(9918) <= not b or a;
    layer2_outputs(9919) <= not b;
    layer2_outputs(9920) <= not b or a;
    layer2_outputs(9921) <= not b or a;
    layer2_outputs(9922) <= b;
    layer2_outputs(9923) <= not b or a;
    layer2_outputs(9924) <= b and not a;
    layer2_outputs(9925) <= not (a or b);
    layer2_outputs(9926) <= not (a and b);
    layer2_outputs(9927) <= not (a and b);
    layer2_outputs(9928) <= b;
    layer2_outputs(9929) <= '0';
    layer2_outputs(9930) <= not (a and b);
    layer2_outputs(9931) <= not a;
    layer2_outputs(9932) <= not a;
    layer2_outputs(9933) <= b and not a;
    layer2_outputs(9934) <= not b;
    layer2_outputs(9935) <= b and not a;
    layer2_outputs(9936) <= not a or b;
    layer2_outputs(9937) <= '1';
    layer2_outputs(9938) <= not b;
    layer2_outputs(9939) <= a;
    layer2_outputs(9940) <= a;
    layer2_outputs(9941) <= not a or b;
    layer2_outputs(9942) <= b and not a;
    layer2_outputs(9943) <= a;
    layer2_outputs(9944) <= a and b;
    layer2_outputs(9945) <= not b or a;
    layer2_outputs(9946) <= '0';
    layer2_outputs(9947) <= b;
    layer2_outputs(9948) <= a or b;
    layer2_outputs(9949) <= b and not a;
    layer2_outputs(9950) <= a;
    layer2_outputs(9951) <= a;
    layer2_outputs(9952) <= not (a or b);
    layer2_outputs(9953) <= a;
    layer2_outputs(9954) <= not (a xor b);
    layer2_outputs(9955) <= '1';
    layer2_outputs(9956) <= not b or a;
    layer2_outputs(9957) <= not (a or b);
    layer2_outputs(9958) <= not (a or b);
    layer2_outputs(9959) <= b and not a;
    layer2_outputs(9960) <= not a or b;
    layer2_outputs(9961) <= b and not a;
    layer2_outputs(9962) <= a;
    layer2_outputs(9963) <= not b;
    layer2_outputs(9964) <= a xor b;
    layer2_outputs(9965) <= '1';
    layer2_outputs(9966) <= '1';
    layer2_outputs(9967) <= a and not b;
    layer2_outputs(9968) <= '1';
    layer2_outputs(9969) <= a;
    layer2_outputs(9970) <= not (a or b);
    layer2_outputs(9971) <= '0';
    layer2_outputs(9972) <= not (a or b);
    layer2_outputs(9973) <= a and not b;
    layer2_outputs(9974) <= a and b;
    layer2_outputs(9975) <= a;
    layer2_outputs(9976) <= not b or a;
    layer2_outputs(9977) <= a and b;
    layer2_outputs(9978) <= b;
    layer2_outputs(9979) <= '0';
    layer2_outputs(9980) <= not b or a;
    layer2_outputs(9981) <= a or b;
    layer2_outputs(9982) <= b and not a;
    layer2_outputs(9983) <= not a or b;
    layer2_outputs(9984) <= a or b;
    layer2_outputs(9985) <= '1';
    layer2_outputs(9986) <= a xor b;
    layer2_outputs(9987) <= b;
    layer2_outputs(9988) <= not b or a;
    layer2_outputs(9989) <= not a;
    layer2_outputs(9990) <= not a;
    layer2_outputs(9991) <= '1';
    layer2_outputs(9992) <= not (a or b);
    layer2_outputs(9993) <= not b;
    layer2_outputs(9994) <= not a or b;
    layer2_outputs(9995) <= '0';
    layer2_outputs(9996) <= not b;
    layer2_outputs(9997) <= not a;
    layer2_outputs(9998) <= b;
    layer2_outputs(9999) <= b;
    layer2_outputs(10000) <= not (a or b);
    layer2_outputs(10001) <= b and not a;
    layer2_outputs(10002) <= a xor b;
    layer2_outputs(10003) <= a;
    layer2_outputs(10004) <= b;
    layer2_outputs(10005) <= '1';
    layer2_outputs(10006) <= b;
    layer2_outputs(10007) <= a;
    layer2_outputs(10008) <= not (a or b);
    layer2_outputs(10009) <= a and not b;
    layer2_outputs(10010) <= not b;
    layer2_outputs(10011) <= b;
    layer2_outputs(10012) <= not (a xor b);
    layer2_outputs(10013) <= a and not b;
    layer2_outputs(10014) <= a;
    layer2_outputs(10015) <= a and b;
    layer2_outputs(10016) <= a or b;
    layer2_outputs(10017) <= not (a or b);
    layer2_outputs(10018) <= not b;
    layer2_outputs(10019) <= not b;
    layer2_outputs(10020) <= not (a and b);
    layer2_outputs(10021) <= a;
    layer2_outputs(10022) <= a and b;
    layer2_outputs(10023) <= a and not b;
    layer2_outputs(10024) <= not a;
    layer2_outputs(10025) <= a and not b;
    layer2_outputs(10026) <= not b;
    layer2_outputs(10027) <= a;
    layer2_outputs(10028) <= not a;
    layer2_outputs(10029) <= b;
    layer2_outputs(10030) <= '1';
    layer2_outputs(10031) <= not (a and b);
    layer2_outputs(10032) <= not a or b;
    layer2_outputs(10033) <= a or b;
    layer2_outputs(10034) <= not b;
    layer2_outputs(10035) <= not b;
    layer2_outputs(10036) <= b;
    layer2_outputs(10037) <= a;
    layer2_outputs(10038) <= not b;
    layer2_outputs(10039) <= not b;
    layer2_outputs(10040) <= b;
    layer2_outputs(10041) <= not b or a;
    layer2_outputs(10042) <= not a;
    layer2_outputs(10043) <= not (a xor b);
    layer2_outputs(10044) <= b and not a;
    layer2_outputs(10045) <= '1';
    layer2_outputs(10046) <= not a;
    layer2_outputs(10047) <= a xor b;
    layer2_outputs(10048) <= a and not b;
    layer2_outputs(10049) <= a or b;
    layer2_outputs(10050) <= not a or b;
    layer2_outputs(10051) <= not a;
    layer2_outputs(10052) <= not a;
    layer2_outputs(10053) <= not b or a;
    layer2_outputs(10054) <= a xor b;
    layer2_outputs(10055) <= not (a or b);
    layer2_outputs(10056) <= not b;
    layer2_outputs(10057) <= '0';
    layer2_outputs(10058) <= a or b;
    layer2_outputs(10059) <= a and b;
    layer2_outputs(10060) <= a and b;
    layer2_outputs(10061) <= a or b;
    layer2_outputs(10062) <= a;
    layer2_outputs(10063) <= a and b;
    layer2_outputs(10064) <= not a;
    layer2_outputs(10065) <= '1';
    layer2_outputs(10066) <= b;
    layer2_outputs(10067) <= b and not a;
    layer2_outputs(10068) <= not (a and b);
    layer2_outputs(10069) <= not a;
    layer2_outputs(10070) <= not b;
    layer2_outputs(10071) <= a or b;
    layer2_outputs(10072) <= not a;
    layer2_outputs(10073) <= not a or b;
    layer2_outputs(10074) <= a and b;
    layer2_outputs(10075) <= a or b;
    layer2_outputs(10076) <= not (a or b);
    layer2_outputs(10077) <= not a;
    layer2_outputs(10078) <= a;
    layer2_outputs(10079) <= b and not a;
    layer2_outputs(10080) <= not b;
    layer2_outputs(10081) <= not b or a;
    layer2_outputs(10082) <= not b;
    layer2_outputs(10083) <= a;
    layer2_outputs(10084) <= not b;
    layer2_outputs(10085) <= a xor b;
    layer2_outputs(10086) <= a or b;
    layer2_outputs(10087) <= a;
    layer2_outputs(10088) <= b and not a;
    layer2_outputs(10089) <= a xor b;
    layer2_outputs(10090) <= not (a or b);
    layer2_outputs(10091) <= b;
    layer2_outputs(10092) <= not (a or b);
    layer2_outputs(10093) <= b;
    layer2_outputs(10094) <= b;
    layer2_outputs(10095) <= not a or b;
    layer2_outputs(10096) <= not a;
    layer2_outputs(10097) <= a and b;
    layer2_outputs(10098) <= not a or b;
    layer2_outputs(10099) <= not (a and b);
    layer2_outputs(10100) <= a xor b;
    layer2_outputs(10101) <= not a or b;
    layer2_outputs(10102) <= a or b;
    layer2_outputs(10103) <= '0';
    layer2_outputs(10104) <= not b;
    layer2_outputs(10105) <= not a or b;
    layer2_outputs(10106) <= a and not b;
    layer2_outputs(10107) <= not a or b;
    layer2_outputs(10108) <= a and not b;
    layer2_outputs(10109) <= not (a or b);
    layer2_outputs(10110) <= b;
    layer2_outputs(10111) <= not (a and b);
    layer2_outputs(10112) <= not (a and b);
    layer2_outputs(10113) <= not b;
    layer2_outputs(10114) <= not b or a;
    layer2_outputs(10115) <= not (a xor b);
    layer2_outputs(10116) <= '1';
    layer2_outputs(10117) <= a or b;
    layer2_outputs(10118) <= not (a or b);
    layer2_outputs(10119) <= not a or b;
    layer2_outputs(10120) <= '1';
    layer2_outputs(10121) <= a xor b;
    layer2_outputs(10122) <= not b;
    layer2_outputs(10123) <= not a;
    layer2_outputs(10124) <= b;
    layer2_outputs(10125) <= not a;
    layer2_outputs(10126) <= not b;
    layer2_outputs(10127) <= b;
    layer2_outputs(10128) <= b;
    layer2_outputs(10129) <= a or b;
    layer2_outputs(10130) <= not b;
    layer2_outputs(10131) <= b;
    layer2_outputs(10132) <= a and b;
    layer2_outputs(10133) <= '1';
    layer2_outputs(10134) <= b;
    layer2_outputs(10135) <= not (a or b);
    layer2_outputs(10136) <= not a;
    layer2_outputs(10137) <= not b or a;
    layer2_outputs(10138) <= a or b;
    layer2_outputs(10139) <= a;
    layer2_outputs(10140) <= not b or a;
    layer2_outputs(10141) <= not (a and b);
    layer2_outputs(10142) <= a and b;
    layer2_outputs(10143) <= not (a or b);
    layer2_outputs(10144) <= not b;
    layer2_outputs(10145) <= b;
    layer2_outputs(10146) <= not (a or b);
    layer2_outputs(10147) <= not b or a;
    layer2_outputs(10148) <= not a;
    layer2_outputs(10149) <= a and not b;
    layer2_outputs(10150) <= not b;
    layer2_outputs(10151) <= b;
    layer2_outputs(10152) <= b;
    layer2_outputs(10153) <= not b;
    layer2_outputs(10154) <= not b;
    layer2_outputs(10155) <= a and b;
    layer2_outputs(10156) <= not b or a;
    layer2_outputs(10157) <= a;
    layer2_outputs(10158) <= a and b;
    layer2_outputs(10159) <= a and not b;
    layer2_outputs(10160) <= not b;
    layer2_outputs(10161) <= a or b;
    layer2_outputs(10162) <= not a;
    layer2_outputs(10163) <= not a or b;
    layer2_outputs(10164) <= a and not b;
    layer2_outputs(10165) <= '0';
    layer2_outputs(10166) <= not b;
    layer2_outputs(10167) <= not b;
    layer2_outputs(10168) <= not a;
    layer2_outputs(10169) <= not (a or b);
    layer2_outputs(10170) <= '0';
    layer2_outputs(10171) <= a;
    layer2_outputs(10172) <= b;
    layer2_outputs(10173) <= b and not a;
    layer2_outputs(10174) <= '0';
    layer2_outputs(10175) <= a;
    layer2_outputs(10176) <= not a or b;
    layer2_outputs(10177) <= a;
    layer2_outputs(10178) <= not (a or b);
    layer2_outputs(10179) <= a and b;
    layer2_outputs(10180) <= not a;
    layer2_outputs(10181) <= not (a or b);
    layer2_outputs(10182) <= not (a or b);
    layer2_outputs(10183) <= a and b;
    layer2_outputs(10184) <= not (a or b);
    layer2_outputs(10185) <= a or b;
    layer2_outputs(10186) <= not b or a;
    layer2_outputs(10187) <= not a or b;
    layer2_outputs(10188) <= not (a and b);
    layer2_outputs(10189) <= a;
    layer2_outputs(10190) <= a and not b;
    layer2_outputs(10191) <= not (a and b);
    layer2_outputs(10192) <= a and b;
    layer2_outputs(10193) <= b;
    layer2_outputs(10194) <= a or b;
    layer2_outputs(10195) <= a or b;
    layer2_outputs(10196) <= a or b;
    layer2_outputs(10197) <= not b;
    layer2_outputs(10198) <= a;
    layer2_outputs(10199) <= a or b;
    layer2_outputs(10200) <= '0';
    layer2_outputs(10201) <= '1';
    layer2_outputs(10202) <= '0';
    layer2_outputs(10203) <= a;
    layer2_outputs(10204) <= not a;
    layer2_outputs(10205) <= not b;
    layer2_outputs(10206) <= not a or b;
    layer2_outputs(10207) <= not (a or b);
    layer2_outputs(10208) <= not (a or b);
    layer2_outputs(10209) <= a;
    layer2_outputs(10210) <= not b;
    layer2_outputs(10211) <= a and b;
    layer2_outputs(10212) <= a;
    layer2_outputs(10213) <= not a or b;
    layer2_outputs(10214) <= a;
    layer2_outputs(10215) <= a and b;
    layer2_outputs(10216) <= not a;
    layer2_outputs(10217) <= not b;
    layer2_outputs(10218) <= not a;
    layer2_outputs(10219) <= not (a or b);
    layer2_outputs(10220) <= b;
    layer2_outputs(10221) <= not a;
    layer2_outputs(10222) <= a;
    layer2_outputs(10223) <= not (a or b);
    layer2_outputs(10224) <= not b or a;
    layer2_outputs(10225) <= not a;
    layer2_outputs(10226) <= b;
    layer2_outputs(10227) <= b;
    layer2_outputs(10228) <= a;
    layer2_outputs(10229) <= b;
    layer2_outputs(10230) <= not a;
    layer2_outputs(10231) <= not a or b;
    layer2_outputs(10232) <= b;
    layer2_outputs(10233) <= not b;
    layer2_outputs(10234) <= b and not a;
    layer2_outputs(10235) <= b and not a;
    layer2_outputs(10236) <= not a;
    layer2_outputs(10237) <= not (a and b);
    layer2_outputs(10238) <= a xor b;
    layer2_outputs(10239) <= a or b;
    layer2_outputs(10240) <= '1';
    layer2_outputs(10241) <= b and not a;
    layer2_outputs(10242) <= a xor b;
    layer2_outputs(10243) <= b;
    layer2_outputs(10244) <= not a;
    layer2_outputs(10245) <= a or b;
    layer2_outputs(10246) <= a;
    layer2_outputs(10247) <= not (a or b);
    layer2_outputs(10248) <= a and not b;
    layer2_outputs(10249) <= not (a xor b);
    layer2_outputs(10250) <= not b or a;
    layer2_outputs(10251) <= not b or a;
    layer2_outputs(10252) <= not a or b;
    layer2_outputs(10253) <= not a;
    layer2_outputs(10254) <= not a;
    layer2_outputs(10255) <= a and not b;
    layer2_outputs(10256) <= not (a or b);
    layer2_outputs(10257) <= not (a xor b);
    layer2_outputs(10258) <= not a;
    layer2_outputs(10259) <= not b or a;
    layer2_outputs(10260) <= not (a or b);
    layer2_outputs(10261) <= not (a xor b);
    layer2_outputs(10262) <= not a or b;
    layer2_outputs(10263) <= not (a and b);
    layer2_outputs(10264) <= not b;
    layer2_outputs(10265) <= not b;
    layer2_outputs(10266) <= b;
    layer2_outputs(10267) <= not a;
    layer2_outputs(10268) <= b;
    layer2_outputs(10269) <= not b or a;
    layer2_outputs(10270) <= a or b;
    layer2_outputs(10271) <= not b;
    layer2_outputs(10272) <= not (a or b);
    layer2_outputs(10273) <= not b;
    layer2_outputs(10274) <= not b;
    layer2_outputs(10275) <= b;
    layer2_outputs(10276) <= b and not a;
    layer2_outputs(10277) <= '0';
    layer2_outputs(10278) <= a xor b;
    layer2_outputs(10279) <= a and b;
    layer2_outputs(10280) <= not a;
    layer2_outputs(10281) <= not a;
    layer2_outputs(10282) <= not a or b;
    layer2_outputs(10283) <= not b;
    layer2_outputs(10284) <= b and not a;
    layer2_outputs(10285) <= '1';
    layer2_outputs(10286) <= '0';
    layer2_outputs(10287) <= a and not b;
    layer2_outputs(10288) <= b;
    layer2_outputs(10289) <= not b or a;
    layer2_outputs(10290) <= '1';
    layer2_outputs(10291) <= not a or b;
    layer2_outputs(10292) <= a and not b;
    layer2_outputs(10293) <= a and b;
    layer2_outputs(10294) <= not b or a;
    layer2_outputs(10295) <= b and not a;
    layer2_outputs(10296) <= not b;
    layer2_outputs(10297) <= b and not a;
    layer2_outputs(10298) <= a or b;
    layer2_outputs(10299) <= a;
    layer2_outputs(10300) <= not a;
    layer2_outputs(10301) <= a;
    layer2_outputs(10302) <= not a or b;
    layer2_outputs(10303) <= a xor b;
    layer2_outputs(10304) <= not a or b;
    layer2_outputs(10305) <= a and not b;
    layer2_outputs(10306) <= a or b;
    layer2_outputs(10307) <= b;
    layer2_outputs(10308) <= not a or b;
    layer2_outputs(10309) <= not (a and b);
    layer2_outputs(10310) <= '0';
    layer2_outputs(10311) <= not b;
    layer2_outputs(10312) <= not a;
    layer2_outputs(10313) <= not (a xor b);
    layer2_outputs(10314) <= not b;
    layer2_outputs(10315) <= not b or a;
    layer2_outputs(10316) <= not a;
    layer2_outputs(10317) <= a and b;
    layer2_outputs(10318) <= b;
    layer2_outputs(10319) <= not a;
    layer2_outputs(10320) <= not (a or b);
    layer2_outputs(10321) <= not b;
    layer2_outputs(10322) <= not (a and b);
    layer2_outputs(10323) <= not a;
    layer2_outputs(10324) <= b;
    layer2_outputs(10325) <= not b;
    layer2_outputs(10326) <= a;
    layer2_outputs(10327) <= not a or b;
    layer2_outputs(10328) <= b and not a;
    layer2_outputs(10329) <= not (a or b);
    layer2_outputs(10330) <= not a;
    layer2_outputs(10331) <= b;
    layer2_outputs(10332) <= a and not b;
    layer2_outputs(10333) <= not b;
    layer2_outputs(10334) <= not b or a;
    layer2_outputs(10335) <= '0';
    layer2_outputs(10336) <= '0';
    layer2_outputs(10337) <= not a;
    layer2_outputs(10338) <= not (a and b);
    layer2_outputs(10339) <= not (a xor b);
    layer2_outputs(10340) <= not b;
    layer2_outputs(10341) <= a and b;
    layer2_outputs(10342) <= a and b;
    layer2_outputs(10343) <= b;
    layer2_outputs(10344) <= b and not a;
    layer2_outputs(10345) <= not (a or b);
    layer2_outputs(10346) <= not b or a;
    layer2_outputs(10347) <= b;
    layer2_outputs(10348) <= not b;
    layer2_outputs(10349) <= a or b;
    layer2_outputs(10350) <= a and b;
    layer2_outputs(10351) <= a;
    layer2_outputs(10352) <= not (a or b);
    layer2_outputs(10353) <= not b;
    layer2_outputs(10354) <= not (a or b);
    layer2_outputs(10355) <= not a;
    layer2_outputs(10356) <= '1';
    layer2_outputs(10357) <= not a;
    layer2_outputs(10358) <= not (a or b);
    layer2_outputs(10359) <= a and b;
    layer2_outputs(10360) <= '0';
    layer2_outputs(10361) <= '1';
    layer2_outputs(10362) <= a;
    layer2_outputs(10363) <= not a;
    layer2_outputs(10364) <= b;
    layer2_outputs(10365) <= b;
    layer2_outputs(10366) <= '0';
    layer2_outputs(10367) <= b and not a;
    layer2_outputs(10368) <= a;
    layer2_outputs(10369) <= not a;
    layer2_outputs(10370) <= not (a and b);
    layer2_outputs(10371) <= a;
    layer2_outputs(10372) <= not b or a;
    layer2_outputs(10373) <= not b;
    layer2_outputs(10374) <= not b;
    layer2_outputs(10375) <= b;
    layer2_outputs(10376) <= b and not a;
    layer2_outputs(10377) <= b and not a;
    layer2_outputs(10378) <= a or b;
    layer2_outputs(10379) <= not b or a;
    layer2_outputs(10380) <= a xor b;
    layer2_outputs(10381) <= b;
    layer2_outputs(10382) <= b;
    layer2_outputs(10383) <= not b;
    layer2_outputs(10384) <= a or b;
    layer2_outputs(10385) <= a and b;
    layer2_outputs(10386) <= a;
    layer2_outputs(10387) <= a and b;
    layer2_outputs(10388) <= not b;
    layer2_outputs(10389) <= b;
    layer2_outputs(10390) <= b and not a;
    layer2_outputs(10391) <= b;
    layer2_outputs(10392) <= not b;
    layer2_outputs(10393) <= a or b;
    layer2_outputs(10394) <= a or b;
    layer2_outputs(10395) <= a;
    layer2_outputs(10396) <= not a;
    layer2_outputs(10397) <= b;
    layer2_outputs(10398) <= not b;
    layer2_outputs(10399) <= not (a and b);
    layer2_outputs(10400) <= not b;
    layer2_outputs(10401) <= b;
    layer2_outputs(10402) <= b and not a;
    layer2_outputs(10403) <= not b;
    layer2_outputs(10404) <= a or b;
    layer2_outputs(10405) <= a;
    layer2_outputs(10406) <= b;
    layer2_outputs(10407) <= not a;
    layer2_outputs(10408) <= a xor b;
    layer2_outputs(10409) <= not a;
    layer2_outputs(10410) <= not a;
    layer2_outputs(10411) <= not (a or b);
    layer2_outputs(10412) <= not (a and b);
    layer2_outputs(10413) <= b;
    layer2_outputs(10414) <= a;
    layer2_outputs(10415) <= not b or a;
    layer2_outputs(10416) <= not (a and b);
    layer2_outputs(10417) <= a xor b;
    layer2_outputs(10418) <= not a;
    layer2_outputs(10419) <= not (a and b);
    layer2_outputs(10420) <= not b or a;
    layer2_outputs(10421) <= not a;
    layer2_outputs(10422) <= b;
    layer2_outputs(10423) <= a;
    layer2_outputs(10424) <= a or b;
    layer2_outputs(10425) <= b;
    layer2_outputs(10426) <= b and not a;
    layer2_outputs(10427) <= b and not a;
    layer2_outputs(10428) <= b and not a;
    layer2_outputs(10429) <= not a;
    layer2_outputs(10430) <= a;
    layer2_outputs(10431) <= b and not a;
    layer2_outputs(10432) <= a;
    layer2_outputs(10433) <= a or b;
    layer2_outputs(10434) <= b;
    layer2_outputs(10435) <= not b;
    layer2_outputs(10436) <= a or b;
    layer2_outputs(10437) <= not (a and b);
    layer2_outputs(10438) <= b;
    layer2_outputs(10439) <= a or b;
    layer2_outputs(10440) <= '0';
    layer2_outputs(10441) <= a or b;
    layer2_outputs(10442) <= '0';
    layer2_outputs(10443) <= not b or a;
    layer2_outputs(10444) <= a;
    layer2_outputs(10445) <= not a;
    layer2_outputs(10446) <= not a;
    layer2_outputs(10447) <= a;
    layer2_outputs(10448) <= a and b;
    layer2_outputs(10449) <= a;
    layer2_outputs(10450) <= not b;
    layer2_outputs(10451) <= a and b;
    layer2_outputs(10452) <= not b or a;
    layer2_outputs(10453) <= not a or b;
    layer2_outputs(10454) <= not b or a;
    layer2_outputs(10455) <= not b or a;
    layer2_outputs(10456) <= '1';
    layer2_outputs(10457) <= not (a or b);
    layer2_outputs(10458) <= not a or b;
    layer2_outputs(10459) <= a;
    layer2_outputs(10460) <= not (a and b);
    layer2_outputs(10461) <= a and not b;
    layer2_outputs(10462) <= b and not a;
    layer2_outputs(10463) <= not (a or b);
    layer2_outputs(10464) <= a and not b;
    layer2_outputs(10465) <= a;
    layer2_outputs(10466) <= not a or b;
    layer2_outputs(10467) <= not a;
    layer2_outputs(10468) <= not (a and b);
    layer2_outputs(10469) <= '1';
    layer2_outputs(10470) <= a and b;
    layer2_outputs(10471) <= a and not b;
    layer2_outputs(10472) <= b;
    layer2_outputs(10473) <= not (a or b);
    layer2_outputs(10474) <= a xor b;
    layer2_outputs(10475) <= a or b;
    layer2_outputs(10476) <= a and not b;
    layer2_outputs(10477) <= '1';
    layer2_outputs(10478) <= a and b;
    layer2_outputs(10479) <= not a or b;
    layer2_outputs(10480) <= not a;
    layer2_outputs(10481) <= '0';
    layer2_outputs(10482) <= b and not a;
    layer2_outputs(10483) <= a and not b;
    layer2_outputs(10484) <= a;
    layer2_outputs(10485) <= a xor b;
    layer2_outputs(10486) <= not (a or b);
    layer2_outputs(10487) <= a and not b;
    layer2_outputs(10488) <= a or b;
    layer2_outputs(10489) <= not a;
    layer2_outputs(10490) <= not b;
    layer2_outputs(10491) <= '1';
    layer2_outputs(10492) <= not b;
    layer2_outputs(10493) <= not (a and b);
    layer2_outputs(10494) <= not a;
    layer2_outputs(10495) <= not a;
    layer2_outputs(10496) <= not a or b;
    layer2_outputs(10497) <= not (a or b);
    layer2_outputs(10498) <= not (a or b);
    layer2_outputs(10499) <= '1';
    layer2_outputs(10500) <= not b;
    layer2_outputs(10501) <= '0';
    layer2_outputs(10502) <= not a or b;
    layer2_outputs(10503) <= not b;
    layer2_outputs(10504) <= b;
    layer2_outputs(10505) <= '0';
    layer2_outputs(10506) <= a;
    layer2_outputs(10507) <= '0';
    layer2_outputs(10508) <= a;
    layer2_outputs(10509) <= a or b;
    layer2_outputs(10510) <= not b or a;
    layer2_outputs(10511) <= not b or a;
    layer2_outputs(10512) <= not b;
    layer2_outputs(10513) <= not (a or b);
    layer2_outputs(10514) <= a and not b;
    layer2_outputs(10515) <= b;
    layer2_outputs(10516) <= not (a and b);
    layer2_outputs(10517) <= not b;
    layer2_outputs(10518) <= a and b;
    layer2_outputs(10519) <= '0';
    layer2_outputs(10520) <= not b or a;
    layer2_outputs(10521) <= a and b;
    layer2_outputs(10522) <= a or b;
    layer2_outputs(10523) <= not (a and b);
    layer2_outputs(10524) <= not (a and b);
    layer2_outputs(10525) <= a;
    layer2_outputs(10526) <= a and b;
    layer2_outputs(10527) <= a xor b;
    layer2_outputs(10528) <= not a or b;
    layer2_outputs(10529) <= not a;
    layer2_outputs(10530) <= b;
    layer2_outputs(10531) <= a xor b;
    layer2_outputs(10532) <= a and not b;
    layer2_outputs(10533) <= not (a or b);
    layer2_outputs(10534) <= a and not b;
    layer2_outputs(10535) <= '0';
    layer2_outputs(10536) <= a and not b;
    layer2_outputs(10537) <= a xor b;
    layer2_outputs(10538) <= not b or a;
    layer2_outputs(10539) <= b;
    layer2_outputs(10540) <= a and b;
    layer2_outputs(10541) <= b;
    layer2_outputs(10542) <= not a;
    layer2_outputs(10543) <= not a or b;
    layer2_outputs(10544) <= a or b;
    layer2_outputs(10545) <= not b or a;
    layer2_outputs(10546) <= not a;
    layer2_outputs(10547) <= a;
    layer2_outputs(10548) <= not (a or b);
    layer2_outputs(10549) <= not (a and b);
    layer2_outputs(10550) <= '1';
    layer2_outputs(10551) <= b;
    layer2_outputs(10552) <= a and not b;
    layer2_outputs(10553) <= '0';
    layer2_outputs(10554) <= not (a or b);
    layer2_outputs(10555) <= b and not a;
    layer2_outputs(10556) <= a;
    layer2_outputs(10557) <= b;
    layer2_outputs(10558) <= b;
    layer2_outputs(10559) <= '0';
    layer2_outputs(10560) <= a and not b;
    layer2_outputs(10561) <= not a or b;
    layer2_outputs(10562) <= a and not b;
    layer2_outputs(10563) <= not a or b;
    layer2_outputs(10564) <= not a or b;
    layer2_outputs(10565) <= not a or b;
    layer2_outputs(10566) <= not b or a;
    layer2_outputs(10567) <= not (a and b);
    layer2_outputs(10568) <= not a or b;
    layer2_outputs(10569) <= a and b;
    layer2_outputs(10570) <= '1';
    layer2_outputs(10571) <= not a;
    layer2_outputs(10572) <= b;
    layer2_outputs(10573) <= not (a and b);
    layer2_outputs(10574) <= a and not b;
    layer2_outputs(10575) <= a and b;
    layer2_outputs(10576) <= a and b;
    layer2_outputs(10577) <= not (a and b);
    layer2_outputs(10578) <= a and not b;
    layer2_outputs(10579) <= a and b;
    layer2_outputs(10580) <= '1';
    layer2_outputs(10581) <= not (a or b);
    layer2_outputs(10582) <= not (a xor b);
    layer2_outputs(10583) <= b;
    layer2_outputs(10584) <= '0';
    layer2_outputs(10585) <= not a;
    layer2_outputs(10586) <= not (a and b);
    layer2_outputs(10587) <= not (a or b);
    layer2_outputs(10588) <= '1';
    layer2_outputs(10589) <= not a or b;
    layer2_outputs(10590) <= a;
    layer2_outputs(10591) <= not a;
    layer2_outputs(10592) <= a xor b;
    layer2_outputs(10593) <= a and b;
    layer2_outputs(10594) <= b;
    layer2_outputs(10595) <= not b;
    layer2_outputs(10596) <= not a;
    layer2_outputs(10597) <= not a;
    layer2_outputs(10598) <= a and b;
    layer2_outputs(10599) <= not a;
    layer2_outputs(10600) <= '0';
    layer2_outputs(10601) <= not b;
    layer2_outputs(10602) <= b;
    layer2_outputs(10603) <= not (a and b);
    layer2_outputs(10604) <= not a or b;
    layer2_outputs(10605) <= b and not a;
    layer2_outputs(10606) <= a and not b;
    layer2_outputs(10607) <= '1';
    layer2_outputs(10608) <= not b;
    layer2_outputs(10609) <= a;
    layer2_outputs(10610) <= not (a xor b);
    layer2_outputs(10611) <= a xor b;
    layer2_outputs(10612) <= a and b;
    layer2_outputs(10613) <= b;
    layer2_outputs(10614) <= not a;
    layer2_outputs(10615) <= b;
    layer2_outputs(10616) <= not b or a;
    layer2_outputs(10617) <= not a;
    layer2_outputs(10618) <= a or b;
    layer2_outputs(10619) <= b and not a;
    layer2_outputs(10620) <= a xor b;
    layer2_outputs(10621) <= not b or a;
    layer2_outputs(10622) <= '1';
    layer2_outputs(10623) <= not b;
    layer2_outputs(10624) <= not b;
    layer2_outputs(10625) <= not b or a;
    layer2_outputs(10626) <= a;
    layer2_outputs(10627) <= not a;
    layer2_outputs(10628) <= a and not b;
    layer2_outputs(10629) <= not a;
    layer2_outputs(10630) <= not b or a;
    layer2_outputs(10631) <= not b;
    layer2_outputs(10632) <= not b;
    layer2_outputs(10633) <= '0';
    layer2_outputs(10634) <= not (a or b);
    layer2_outputs(10635) <= '0';
    layer2_outputs(10636) <= '1';
    layer2_outputs(10637) <= not b;
    layer2_outputs(10638) <= b and not a;
    layer2_outputs(10639) <= a xor b;
    layer2_outputs(10640) <= not a;
    layer2_outputs(10641) <= not b or a;
    layer2_outputs(10642) <= not b;
    layer2_outputs(10643) <= not (a and b);
    layer2_outputs(10644) <= b and not a;
    layer2_outputs(10645) <= not a;
    layer2_outputs(10646) <= b and not a;
    layer2_outputs(10647) <= not (a or b);
    layer2_outputs(10648) <= '1';
    layer2_outputs(10649) <= not b or a;
    layer2_outputs(10650) <= a and not b;
    layer2_outputs(10651) <= a and not b;
    layer2_outputs(10652) <= a xor b;
    layer2_outputs(10653) <= a xor b;
    layer2_outputs(10654) <= a xor b;
    layer2_outputs(10655) <= '1';
    layer2_outputs(10656) <= not a or b;
    layer2_outputs(10657) <= a;
    layer2_outputs(10658) <= a or b;
    layer2_outputs(10659) <= a or b;
    layer2_outputs(10660) <= not b;
    layer2_outputs(10661) <= not a or b;
    layer2_outputs(10662) <= a and not b;
    layer2_outputs(10663) <= a and b;
    layer2_outputs(10664) <= '0';
    layer2_outputs(10665) <= not b or a;
    layer2_outputs(10666) <= not (a or b);
    layer2_outputs(10667) <= '1';
    layer2_outputs(10668) <= a and b;
    layer2_outputs(10669) <= not b or a;
    layer2_outputs(10670) <= not (a or b);
    layer2_outputs(10671) <= not a;
    layer2_outputs(10672) <= not (a xor b);
    layer2_outputs(10673) <= a or b;
    layer2_outputs(10674) <= a or b;
    layer2_outputs(10675) <= not b;
    layer2_outputs(10676) <= a and not b;
    layer2_outputs(10677) <= not b;
    layer2_outputs(10678) <= a and b;
    layer2_outputs(10679) <= not (a or b);
    layer2_outputs(10680) <= not a;
    layer2_outputs(10681) <= a and not b;
    layer2_outputs(10682) <= not b or a;
    layer2_outputs(10683) <= not a;
    layer2_outputs(10684) <= '0';
    layer2_outputs(10685) <= a;
    layer2_outputs(10686) <= '0';
    layer2_outputs(10687) <= a;
    layer2_outputs(10688) <= a and not b;
    layer2_outputs(10689) <= '0';
    layer2_outputs(10690) <= a and not b;
    layer2_outputs(10691) <= not b;
    layer2_outputs(10692) <= not (a and b);
    layer2_outputs(10693) <= '1';
    layer2_outputs(10694) <= a or b;
    layer2_outputs(10695) <= not b;
    layer2_outputs(10696) <= a and not b;
    layer2_outputs(10697) <= not b;
    layer2_outputs(10698) <= '1';
    layer2_outputs(10699) <= not (a and b);
    layer2_outputs(10700) <= b;
    layer2_outputs(10701) <= a or b;
    layer2_outputs(10702) <= '1';
    layer2_outputs(10703) <= b;
    layer2_outputs(10704) <= a and not b;
    layer2_outputs(10705) <= not b or a;
    layer2_outputs(10706) <= not a or b;
    layer2_outputs(10707) <= not a or b;
    layer2_outputs(10708) <= a xor b;
    layer2_outputs(10709) <= not b;
    layer2_outputs(10710) <= '1';
    layer2_outputs(10711) <= not (a and b);
    layer2_outputs(10712) <= a xor b;
    layer2_outputs(10713) <= not b;
    layer2_outputs(10714) <= not b or a;
    layer2_outputs(10715) <= a or b;
    layer2_outputs(10716) <= '1';
    layer2_outputs(10717) <= not a or b;
    layer2_outputs(10718) <= not b or a;
    layer2_outputs(10719) <= a;
    layer2_outputs(10720) <= b;
    layer2_outputs(10721) <= a and not b;
    layer2_outputs(10722) <= a;
    layer2_outputs(10723) <= not a or b;
    layer2_outputs(10724) <= not (a or b);
    layer2_outputs(10725) <= not a;
    layer2_outputs(10726) <= not a;
    layer2_outputs(10727) <= '1';
    layer2_outputs(10728) <= b and not a;
    layer2_outputs(10729) <= '1';
    layer2_outputs(10730) <= not a;
    layer2_outputs(10731) <= a and b;
    layer2_outputs(10732) <= b;
    layer2_outputs(10733) <= '1';
    layer2_outputs(10734) <= b;
    layer2_outputs(10735) <= not b or a;
    layer2_outputs(10736) <= not b;
    layer2_outputs(10737) <= a;
    layer2_outputs(10738) <= a;
    layer2_outputs(10739) <= a and not b;
    layer2_outputs(10740) <= not b;
    layer2_outputs(10741) <= a;
    layer2_outputs(10742) <= a;
    layer2_outputs(10743) <= b;
    layer2_outputs(10744) <= '1';
    layer2_outputs(10745) <= '0';
    layer2_outputs(10746) <= b;
    layer2_outputs(10747) <= not a;
    layer2_outputs(10748) <= a and b;
    layer2_outputs(10749) <= not b or a;
    layer2_outputs(10750) <= not b;
    layer2_outputs(10751) <= not (a and b);
    layer2_outputs(10752) <= a and b;
    layer2_outputs(10753) <= '1';
    layer2_outputs(10754) <= '1';
    layer2_outputs(10755) <= a;
    layer2_outputs(10756) <= not b;
    layer2_outputs(10757) <= a;
    layer2_outputs(10758) <= a xor b;
    layer2_outputs(10759) <= a;
    layer2_outputs(10760) <= not b or a;
    layer2_outputs(10761) <= not a;
    layer2_outputs(10762) <= a and b;
    layer2_outputs(10763) <= a xor b;
    layer2_outputs(10764) <= a;
    layer2_outputs(10765) <= a;
    layer2_outputs(10766) <= a or b;
    layer2_outputs(10767) <= a and b;
    layer2_outputs(10768) <= a;
    layer2_outputs(10769) <= not b;
    layer2_outputs(10770) <= '1';
    layer2_outputs(10771) <= '1';
    layer2_outputs(10772) <= not (a or b);
    layer2_outputs(10773) <= a and b;
    layer2_outputs(10774) <= not a;
    layer2_outputs(10775) <= not b;
    layer2_outputs(10776) <= not (a or b);
    layer2_outputs(10777) <= not a;
    layer2_outputs(10778) <= b and not a;
    layer2_outputs(10779) <= a;
    layer2_outputs(10780) <= a and b;
    layer2_outputs(10781) <= a and not b;
    layer2_outputs(10782) <= not b;
    layer2_outputs(10783) <= a or b;
    layer2_outputs(10784) <= a and b;
    layer2_outputs(10785) <= not (a xor b);
    layer2_outputs(10786) <= not (a or b);
    layer2_outputs(10787) <= not a;
    layer2_outputs(10788) <= not a;
    layer2_outputs(10789) <= a;
    layer2_outputs(10790) <= a and not b;
    layer2_outputs(10791) <= a;
    layer2_outputs(10792) <= a xor b;
    layer2_outputs(10793) <= a and not b;
    layer2_outputs(10794) <= b and not a;
    layer2_outputs(10795) <= b;
    layer2_outputs(10796) <= a;
    layer2_outputs(10797) <= not a or b;
    layer2_outputs(10798) <= not (a and b);
    layer2_outputs(10799) <= not b or a;
    layer2_outputs(10800) <= a and not b;
    layer2_outputs(10801) <= not b or a;
    layer2_outputs(10802) <= '0';
    layer2_outputs(10803) <= '1';
    layer2_outputs(10804) <= b and not a;
    layer2_outputs(10805) <= not b or a;
    layer2_outputs(10806) <= not (a or b);
    layer2_outputs(10807) <= b;
    layer2_outputs(10808) <= b and not a;
    layer2_outputs(10809) <= '1';
    layer2_outputs(10810) <= a and b;
    layer2_outputs(10811) <= a and b;
    layer2_outputs(10812) <= a;
    layer2_outputs(10813) <= a and not b;
    layer2_outputs(10814) <= b;
    layer2_outputs(10815) <= b and not a;
    layer2_outputs(10816) <= a and not b;
    layer2_outputs(10817) <= not b or a;
    layer2_outputs(10818) <= a and not b;
    layer2_outputs(10819) <= a xor b;
    layer2_outputs(10820) <= a;
    layer2_outputs(10821) <= b;
    layer2_outputs(10822) <= a;
    layer2_outputs(10823) <= b;
    layer2_outputs(10824) <= not (a and b);
    layer2_outputs(10825) <= b;
    layer2_outputs(10826) <= not (a xor b);
    layer2_outputs(10827) <= b and not a;
    layer2_outputs(10828) <= a and b;
    layer2_outputs(10829) <= a or b;
    layer2_outputs(10830) <= a or b;
    layer2_outputs(10831) <= not (a or b);
    layer2_outputs(10832) <= not a;
    layer2_outputs(10833) <= b and not a;
    layer2_outputs(10834) <= not a or b;
    layer2_outputs(10835) <= not (a and b);
    layer2_outputs(10836) <= not (a or b);
    layer2_outputs(10837) <= a;
    layer2_outputs(10838) <= not a;
    layer2_outputs(10839) <= not a;
    layer2_outputs(10840) <= a and not b;
    layer2_outputs(10841) <= b;
    layer2_outputs(10842) <= a and b;
    layer2_outputs(10843) <= a;
    layer2_outputs(10844) <= '0';
    layer2_outputs(10845) <= a;
    layer2_outputs(10846) <= '0';
    layer2_outputs(10847) <= not (a and b);
    layer2_outputs(10848) <= b;
    layer2_outputs(10849) <= not b;
    layer2_outputs(10850) <= a or b;
    layer2_outputs(10851) <= b;
    layer2_outputs(10852) <= b and not a;
    layer2_outputs(10853) <= not a;
    layer2_outputs(10854) <= '0';
    layer2_outputs(10855) <= not b or a;
    layer2_outputs(10856) <= not (a and b);
    layer2_outputs(10857) <= '1';
    layer2_outputs(10858) <= a and not b;
    layer2_outputs(10859) <= a or b;
    layer2_outputs(10860) <= '0';
    layer2_outputs(10861) <= a;
    layer2_outputs(10862) <= not b;
    layer2_outputs(10863) <= not (a or b);
    layer2_outputs(10864) <= not (a xor b);
    layer2_outputs(10865) <= not b or a;
    layer2_outputs(10866) <= not b or a;
    layer2_outputs(10867) <= a;
    layer2_outputs(10868) <= not (a or b);
    layer2_outputs(10869) <= '1';
    layer2_outputs(10870) <= '0';
    layer2_outputs(10871) <= '0';
    layer2_outputs(10872) <= not (a xor b);
    layer2_outputs(10873) <= a;
    layer2_outputs(10874) <= a or b;
    layer2_outputs(10875) <= not b;
    layer2_outputs(10876) <= not b;
    layer2_outputs(10877) <= not b;
    layer2_outputs(10878) <= not (a or b);
    layer2_outputs(10879) <= b;
    layer2_outputs(10880) <= a;
    layer2_outputs(10881) <= b and not a;
    layer2_outputs(10882) <= a;
    layer2_outputs(10883) <= '0';
    layer2_outputs(10884) <= not b;
    layer2_outputs(10885) <= b and not a;
    layer2_outputs(10886) <= b;
    layer2_outputs(10887) <= a and b;
    layer2_outputs(10888) <= a;
    layer2_outputs(10889) <= not b;
    layer2_outputs(10890) <= not (a or b);
    layer2_outputs(10891) <= a or b;
    layer2_outputs(10892) <= b and not a;
    layer2_outputs(10893) <= not b or a;
    layer2_outputs(10894) <= b;
    layer2_outputs(10895) <= '0';
    layer2_outputs(10896) <= a and not b;
    layer2_outputs(10897) <= a and not b;
    layer2_outputs(10898) <= a and b;
    layer2_outputs(10899) <= a and b;
    layer2_outputs(10900) <= not a;
    layer2_outputs(10901) <= not b;
    layer2_outputs(10902) <= not b;
    layer2_outputs(10903) <= a;
    layer2_outputs(10904) <= b;
    layer2_outputs(10905) <= a;
    layer2_outputs(10906) <= b and not a;
    layer2_outputs(10907) <= a or b;
    layer2_outputs(10908) <= not (a xor b);
    layer2_outputs(10909) <= a;
    layer2_outputs(10910) <= b and not a;
    layer2_outputs(10911) <= not a or b;
    layer2_outputs(10912) <= b;
    layer2_outputs(10913) <= '1';
    layer2_outputs(10914) <= a;
    layer2_outputs(10915) <= not (a and b);
    layer2_outputs(10916) <= '1';
    layer2_outputs(10917) <= b;
    layer2_outputs(10918) <= not b;
    layer2_outputs(10919) <= not b or a;
    layer2_outputs(10920) <= not (a and b);
    layer2_outputs(10921) <= b;
    layer2_outputs(10922) <= not (a and b);
    layer2_outputs(10923) <= b and not a;
    layer2_outputs(10924) <= a and not b;
    layer2_outputs(10925) <= not b;
    layer2_outputs(10926) <= not (a and b);
    layer2_outputs(10927) <= a;
    layer2_outputs(10928) <= not (a and b);
    layer2_outputs(10929) <= not b;
    layer2_outputs(10930) <= a and not b;
    layer2_outputs(10931) <= not b;
    layer2_outputs(10932) <= b and not a;
    layer2_outputs(10933) <= a and not b;
    layer2_outputs(10934) <= not (a xor b);
    layer2_outputs(10935) <= a;
    layer2_outputs(10936) <= not (a and b);
    layer2_outputs(10937) <= a;
    layer2_outputs(10938) <= a and b;
    layer2_outputs(10939) <= not a or b;
    layer2_outputs(10940) <= not a;
    layer2_outputs(10941) <= a and not b;
    layer2_outputs(10942) <= b;
    layer2_outputs(10943) <= '1';
    layer2_outputs(10944) <= b;
    layer2_outputs(10945) <= a and b;
    layer2_outputs(10946) <= not b;
    layer2_outputs(10947) <= not a;
    layer2_outputs(10948) <= a and b;
    layer2_outputs(10949) <= not a;
    layer2_outputs(10950) <= not a;
    layer2_outputs(10951) <= b;
    layer2_outputs(10952) <= not a;
    layer2_outputs(10953) <= not b;
    layer2_outputs(10954) <= a;
    layer2_outputs(10955) <= not a or b;
    layer2_outputs(10956) <= not a;
    layer2_outputs(10957) <= not (a and b);
    layer2_outputs(10958) <= a or b;
    layer2_outputs(10959) <= not (a or b);
    layer2_outputs(10960) <= not a or b;
    layer2_outputs(10961) <= b and not a;
    layer2_outputs(10962) <= not a or b;
    layer2_outputs(10963) <= not b;
    layer2_outputs(10964) <= not a;
    layer2_outputs(10965) <= '1';
    layer2_outputs(10966) <= not (a xor b);
    layer2_outputs(10967) <= not a;
    layer2_outputs(10968) <= not a;
    layer2_outputs(10969) <= not b or a;
    layer2_outputs(10970) <= a and not b;
    layer2_outputs(10971) <= not b;
    layer2_outputs(10972) <= b;
    layer2_outputs(10973) <= not (a or b);
    layer2_outputs(10974) <= a;
    layer2_outputs(10975) <= '0';
    layer2_outputs(10976) <= b;
    layer2_outputs(10977) <= a and b;
    layer2_outputs(10978) <= a;
    layer2_outputs(10979) <= b;
    layer2_outputs(10980) <= not a;
    layer2_outputs(10981) <= not a or b;
    layer2_outputs(10982) <= a;
    layer2_outputs(10983) <= a or b;
    layer2_outputs(10984) <= not a;
    layer2_outputs(10985) <= a;
    layer2_outputs(10986) <= not b or a;
    layer2_outputs(10987) <= a and b;
    layer2_outputs(10988) <= not (a or b);
    layer2_outputs(10989) <= not a or b;
    layer2_outputs(10990) <= not a or b;
    layer2_outputs(10991) <= a and not b;
    layer2_outputs(10992) <= not b;
    layer2_outputs(10993) <= a;
    layer2_outputs(10994) <= a xor b;
    layer2_outputs(10995) <= b and not a;
    layer2_outputs(10996) <= not (a or b);
    layer2_outputs(10997) <= a;
    layer2_outputs(10998) <= b;
    layer2_outputs(10999) <= a;
    layer2_outputs(11000) <= a or b;
    layer2_outputs(11001) <= not (a xor b);
    layer2_outputs(11002) <= a and not b;
    layer2_outputs(11003) <= not a;
    layer2_outputs(11004) <= not (a and b);
    layer2_outputs(11005) <= b;
    layer2_outputs(11006) <= '0';
    layer2_outputs(11007) <= a;
    layer2_outputs(11008) <= '0';
    layer2_outputs(11009) <= not (a xor b);
    layer2_outputs(11010) <= a;
    layer2_outputs(11011) <= a and not b;
    layer2_outputs(11012) <= '0';
    layer2_outputs(11013) <= not b;
    layer2_outputs(11014) <= b and not a;
    layer2_outputs(11015) <= a and b;
    layer2_outputs(11016) <= a and b;
    layer2_outputs(11017) <= not a;
    layer2_outputs(11018) <= not a or b;
    layer2_outputs(11019) <= a and b;
    layer2_outputs(11020) <= a or b;
    layer2_outputs(11021) <= a xor b;
    layer2_outputs(11022) <= b and not a;
    layer2_outputs(11023) <= not (a xor b);
    layer2_outputs(11024) <= '0';
    layer2_outputs(11025) <= not b;
    layer2_outputs(11026) <= not (a and b);
    layer2_outputs(11027) <= a or b;
    layer2_outputs(11028) <= not b;
    layer2_outputs(11029) <= not (a and b);
    layer2_outputs(11030) <= '1';
    layer2_outputs(11031) <= a;
    layer2_outputs(11032) <= a or b;
    layer2_outputs(11033) <= not b;
    layer2_outputs(11034) <= b;
    layer2_outputs(11035) <= a or b;
    layer2_outputs(11036) <= not (a or b);
    layer2_outputs(11037) <= '0';
    layer2_outputs(11038) <= not b;
    layer2_outputs(11039) <= b;
    layer2_outputs(11040) <= not b;
    layer2_outputs(11041) <= not a;
    layer2_outputs(11042) <= a;
    layer2_outputs(11043) <= b and not a;
    layer2_outputs(11044) <= a or b;
    layer2_outputs(11045) <= not b;
    layer2_outputs(11046) <= not a;
    layer2_outputs(11047) <= not a or b;
    layer2_outputs(11048) <= a and b;
    layer2_outputs(11049) <= '0';
    layer2_outputs(11050) <= not b;
    layer2_outputs(11051) <= b;
    layer2_outputs(11052) <= a and not b;
    layer2_outputs(11053) <= a or b;
    layer2_outputs(11054) <= b;
    layer2_outputs(11055) <= not a;
    layer2_outputs(11056) <= '0';
    layer2_outputs(11057) <= '0';
    layer2_outputs(11058) <= a or b;
    layer2_outputs(11059) <= a;
    layer2_outputs(11060) <= a or b;
    layer2_outputs(11061) <= b and not a;
    layer2_outputs(11062) <= not b or a;
    layer2_outputs(11063) <= a or b;
    layer2_outputs(11064) <= a or b;
    layer2_outputs(11065) <= a;
    layer2_outputs(11066) <= '0';
    layer2_outputs(11067) <= not a;
    layer2_outputs(11068) <= a;
    layer2_outputs(11069) <= a and b;
    layer2_outputs(11070) <= not (a and b);
    layer2_outputs(11071) <= not (a or b);
    layer2_outputs(11072) <= not a;
    layer2_outputs(11073) <= not b or a;
    layer2_outputs(11074) <= a;
    layer2_outputs(11075) <= a xor b;
    layer2_outputs(11076) <= not (a and b);
    layer2_outputs(11077) <= not (a or b);
    layer2_outputs(11078) <= '1';
    layer2_outputs(11079) <= a;
    layer2_outputs(11080) <= not (a and b);
    layer2_outputs(11081) <= not b or a;
    layer2_outputs(11082) <= not a;
    layer2_outputs(11083) <= a;
    layer2_outputs(11084) <= a or b;
    layer2_outputs(11085) <= b;
    layer2_outputs(11086) <= a or b;
    layer2_outputs(11087) <= not a;
    layer2_outputs(11088) <= not a;
    layer2_outputs(11089) <= a;
    layer2_outputs(11090) <= not a;
    layer2_outputs(11091) <= b;
    layer2_outputs(11092) <= not (a and b);
    layer2_outputs(11093) <= b and not a;
    layer2_outputs(11094) <= a and not b;
    layer2_outputs(11095) <= b;
    layer2_outputs(11096) <= not b;
    layer2_outputs(11097) <= b;
    layer2_outputs(11098) <= a or b;
    layer2_outputs(11099) <= not a;
    layer2_outputs(11100) <= a and b;
    layer2_outputs(11101) <= b;
    layer2_outputs(11102) <= a xor b;
    layer2_outputs(11103) <= a and not b;
    layer2_outputs(11104) <= a or b;
    layer2_outputs(11105) <= not a or b;
    layer2_outputs(11106) <= not a;
    layer2_outputs(11107) <= a and not b;
    layer2_outputs(11108) <= '1';
    layer2_outputs(11109) <= not (a and b);
    layer2_outputs(11110) <= not b or a;
    layer2_outputs(11111) <= '1';
    layer2_outputs(11112) <= not a or b;
    layer2_outputs(11113) <= a or b;
    layer2_outputs(11114) <= not a;
    layer2_outputs(11115) <= a and b;
    layer2_outputs(11116) <= not a;
    layer2_outputs(11117) <= b;
    layer2_outputs(11118) <= not (a or b);
    layer2_outputs(11119) <= b;
    layer2_outputs(11120) <= not a;
    layer2_outputs(11121) <= b;
    layer2_outputs(11122) <= a or b;
    layer2_outputs(11123) <= a or b;
    layer2_outputs(11124) <= a xor b;
    layer2_outputs(11125) <= not (a or b);
    layer2_outputs(11126) <= b and not a;
    layer2_outputs(11127) <= not a or b;
    layer2_outputs(11128) <= not a or b;
    layer2_outputs(11129) <= not b or a;
    layer2_outputs(11130) <= a and not b;
    layer2_outputs(11131) <= b and not a;
    layer2_outputs(11132) <= not a;
    layer2_outputs(11133) <= not a or b;
    layer2_outputs(11134) <= not b or a;
    layer2_outputs(11135) <= not a;
    layer2_outputs(11136) <= '0';
    layer2_outputs(11137) <= not b or a;
    layer2_outputs(11138) <= '0';
    layer2_outputs(11139) <= a and b;
    layer2_outputs(11140) <= a;
    layer2_outputs(11141) <= not b;
    layer2_outputs(11142) <= not a or b;
    layer2_outputs(11143) <= b and not a;
    layer2_outputs(11144) <= a and not b;
    layer2_outputs(11145) <= not a;
    layer2_outputs(11146) <= a xor b;
    layer2_outputs(11147) <= not (a or b);
    layer2_outputs(11148) <= a;
    layer2_outputs(11149) <= not b;
    layer2_outputs(11150) <= b;
    layer2_outputs(11151) <= not b or a;
    layer2_outputs(11152) <= a;
    layer2_outputs(11153) <= a xor b;
    layer2_outputs(11154) <= '1';
    layer2_outputs(11155) <= a or b;
    layer2_outputs(11156) <= a and b;
    layer2_outputs(11157) <= b;
    layer2_outputs(11158) <= a;
    layer2_outputs(11159) <= a or b;
    layer2_outputs(11160) <= b and not a;
    layer2_outputs(11161) <= not (a xor b);
    layer2_outputs(11162) <= not (a or b);
    layer2_outputs(11163) <= not (a or b);
    layer2_outputs(11164) <= not a;
    layer2_outputs(11165) <= not b or a;
    layer2_outputs(11166) <= a xor b;
    layer2_outputs(11167) <= not a;
    layer2_outputs(11168) <= not (a and b);
    layer2_outputs(11169) <= not b;
    layer2_outputs(11170) <= not a or b;
    layer2_outputs(11171) <= '1';
    layer2_outputs(11172) <= not a;
    layer2_outputs(11173) <= '1';
    layer2_outputs(11174) <= not a or b;
    layer2_outputs(11175) <= not (a or b);
    layer2_outputs(11176) <= not a;
    layer2_outputs(11177) <= a;
    layer2_outputs(11178) <= not a;
    layer2_outputs(11179) <= '1';
    layer2_outputs(11180) <= not b;
    layer2_outputs(11181) <= '1';
    layer2_outputs(11182) <= not b;
    layer2_outputs(11183) <= '0';
    layer2_outputs(11184) <= a and not b;
    layer2_outputs(11185) <= a;
    layer2_outputs(11186) <= b and not a;
    layer2_outputs(11187) <= not b or a;
    layer2_outputs(11188) <= a;
    layer2_outputs(11189) <= not a or b;
    layer2_outputs(11190) <= a and not b;
    layer2_outputs(11191) <= not b;
    layer2_outputs(11192) <= not a or b;
    layer2_outputs(11193) <= a and not b;
    layer2_outputs(11194) <= not b;
    layer2_outputs(11195) <= a and not b;
    layer2_outputs(11196) <= not b or a;
    layer2_outputs(11197) <= not b;
    layer2_outputs(11198) <= '1';
    layer2_outputs(11199) <= not b;
    layer2_outputs(11200) <= b and not a;
    layer2_outputs(11201) <= b and not a;
    layer2_outputs(11202) <= a or b;
    layer2_outputs(11203) <= a;
    layer2_outputs(11204) <= not a;
    layer2_outputs(11205) <= a or b;
    layer2_outputs(11206) <= '0';
    layer2_outputs(11207) <= not (a and b);
    layer2_outputs(11208) <= a or b;
    layer2_outputs(11209) <= a and b;
    layer2_outputs(11210) <= b;
    layer2_outputs(11211) <= a and b;
    layer2_outputs(11212) <= a or b;
    layer2_outputs(11213) <= a or b;
    layer2_outputs(11214) <= a xor b;
    layer2_outputs(11215) <= b;
    layer2_outputs(11216) <= not a or b;
    layer2_outputs(11217) <= a and b;
    layer2_outputs(11218) <= not a;
    layer2_outputs(11219) <= not (a or b);
    layer2_outputs(11220) <= '0';
    layer2_outputs(11221) <= '0';
    layer2_outputs(11222) <= b;
    layer2_outputs(11223) <= a xor b;
    layer2_outputs(11224) <= a;
    layer2_outputs(11225) <= '1';
    layer2_outputs(11226) <= b;
    layer2_outputs(11227) <= not (a or b);
    layer2_outputs(11228) <= not a;
    layer2_outputs(11229) <= not (a and b);
    layer2_outputs(11230) <= a;
    layer2_outputs(11231) <= not b;
    layer2_outputs(11232) <= a;
    layer2_outputs(11233) <= not a or b;
    layer2_outputs(11234) <= a;
    layer2_outputs(11235) <= not b or a;
    layer2_outputs(11236) <= a and b;
    layer2_outputs(11237) <= a and b;
    layer2_outputs(11238) <= not a or b;
    layer2_outputs(11239) <= a or b;
    layer2_outputs(11240) <= a or b;
    layer2_outputs(11241) <= b and not a;
    layer2_outputs(11242) <= not b;
    layer2_outputs(11243) <= a and not b;
    layer2_outputs(11244) <= b;
    layer2_outputs(11245) <= not b;
    layer2_outputs(11246) <= '1';
    layer2_outputs(11247) <= '0';
    layer2_outputs(11248) <= not a;
    layer2_outputs(11249) <= not b or a;
    layer2_outputs(11250) <= '0';
    layer2_outputs(11251) <= not a or b;
    layer2_outputs(11252) <= a;
    layer2_outputs(11253) <= a and not b;
    layer2_outputs(11254) <= not (a or b);
    layer2_outputs(11255) <= b and not a;
    layer2_outputs(11256) <= b and not a;
    layer2_outputs(11257) <= not (a or b);
    layer2_outputs(11258) <= b and not a;
    layer2_outputs(11259) <= a and not b;
    layer2_outputs(11260) <= a and b;
    layer2_outputs(11261) <= not (a and b);
    layer2_outputs(11262) <= not b or a;
    layer2_outputs(11263) <= a xor b;
    layer2_outputs(11264) <= b;
    layer2_outputs(11265) <= a and b;
    layer2_outputs(11266) <= a or b;
    layer2_outputs(11267) <= a and b;
    layer2_outputs(11268) <= not (a xor b);
    layer2_outputs(11269) <= b;
    layer2_outputs(11270) <= b and not a;
    layer2_outputs(11271) <= b and not a;
    layer2_outputs(11272) <= b;
    layer2_outputs(11273) <= not b or a;
    layer2_outputs(11274) <= not b or a;
    layer2_outputs(11275) <= a;
    layer2_outputs(11276) <= b;
    layer2_outputs(11277) <= not b;
    layer2_outputs(11278) <= b;
    layer2_outputs(11279) <= a or b;
    layer2_outputs(11280) <= a;
    layer2_outputs(11281) <= not (a xor b);
    layer2_outputs(11282) <= not (a or b);
    layer2_outputs(11283) <= '0';
    layer2_outputs(11284) <= a and b;
    layer2_outputs(11285) <= not a or b;
    layer2_outputs(11286) <= not a;
    layer2_outputs(11287) <= not b or a;
    layer2_outputs(11288) <= a or b;
    layer2_outputs(11289) <= b;
    layer2_outputs(11290) <= a and b;
    layer2_outputs(11291) <= not b;
    layer2_outputs(11292) <= a or b;
    layer2_outputs(11293) <= '1';
    layer2_outputs(11294) <= a and not b;
    layer2_outputs(11295) <= not (a or b);
    layer2_outputs(11296) <= not b;
    layer2_outputs(11297) <= b;
    layer2_outputs(11298) <= not (a or b);
    layer2_outputs(11299) <= a;
    layer2_outputs(11300) <= not a or b;
    layer2_outputs(11301) <= '1';
    layer2_outputs(11302) <= not b or a;
    layer2_outputs(11303) <= a;
    layer2_outputs(11304) <= a or b;
    layer2_outputs(11305) <= not (a or b);
    layer2_outputs(11306) <= b;
    layer2_outputs(11307) <= '1';
    layer2_outputs(11308) <= a;
    layer2_outputs(11309) <= not (a xor b);
    layer2_outputs(11310) <= not (a or b);
    layer2_outputs(11311) <= not b;
    layer2_outputs(11312) <= not (a xor b);
    layer2_outputs(11313) <= a and not b;
    layer2_outputs(11314) <= not (a or b);
    layer2_outputs(11315) <= a and not b;
    layer2_outputs(11316) <= '1';
    layer2_outputs(11317) <= not (a or b);
    layer2_outputs(11318) <= not a;
    layer2_outputs(11319) <= not a;
    layer2_outputs(11320) <= not a or b;
    layer2_outputs(11321) <= a;
    layer2_outputs(11322) <= not (a or b);
    layer2_outputs(11323) <= not b;
    layer2_outputs(11324) <= b and not a;
    layer2_outputs(11325) <= '1';
    layer2_outputs(11326) <= '0';
    layer2_outputs(11327) <= not (a xor b);
    layer2_outputs(11328) <= not (a and b);
    layer2_outputs(11329) <= not b;
    layer2_outputs(11330) <= a xor b;
    layer2_outputs(11331) <= b;
    layer2_outputs(11332) <= b;
    layer2_outputs(11333) <= b and not a;
    layer2_outputs(11334) <= not b or a;
    layer2_outputs(11335) <= not a;
    layer2_outputs(11336) <= '1';
    layer2_outputs(11337) <= not a;
    layer2_outputs(11338) <= '1';
    layer2_outputs(11339) <= not (a or b);
    layer2_outputs(11340) <= not (a or b);
    layer2_outputs(11341) <= a;
    layer2_outputs(11342) <= b and not a;
    layer2_outputs(11343) <= b and not a;
    layer2_outputs(11344) <= a and not b;
    layer2_outputs(11345) <= not (a or b);
    layer2_outputs(11346) <= a xor b;
    layer2_outputs(11347) <= not b or a;
    layer2_outputs(11348) <= not (a and b);
    layer2_outputs(11349) <= a;
    layer2_outputs(11350) <= a and not b;
    layer2_outputs(11351) <= not (a and b);
    layer2_outputs(11352) <= not (a and b);
    layer2_outputs(11353) <= '0';
    layer2_outputs(11354) <= not (a or b);
    layer2_outputs(11355) <= not (a or b);
    layer2_outputs(11356) <= not b or a;
    layer2_outputs(11357) <= a and not b;
    layer2_outputs(11358) <= not a;
    layer2_outputs(11359) <= not a;
    layer2_outputs(11360) <= b;
    layer2_outputs(11361) <= not b;
    layer2_outputs(11362) <= b and not a;
    layer2_outputs(11363) <= not (a or b);
    layer2_outputs(11364) <= not a;
    layer2_outputs(11365) <= a or b;
    layer2_outputs(11366) <= a or b;
    layer2_outputs(11367) <= b;
    layer2_outputs(11368) <= a and not b;
    layer2_outputs(11369) <= b;
    layer2_outputs(11370) <= not a;
    layer2_outputs(11371) <= a and not b;
    layer2_outputs(11372) <= '1';
    layer2_outputs(11373) <= b;
    layer2_outputs(11374) <= a or b;
    layer2_outputs(11375) <= a and b;
    layer2_outputs(11376) <= a or b;
    layer2_outputs(11377) <= a;
    layer2_outputs(11378) <= not a or b;
    layer2_outputs(11379) <= a or b;
    layer2_outputs(11380) <= '1';
    layer2_outputs(11381) <= b;
    layer2_outputs(11382) <= not b or a;
    layer2_outputs(11383) <= b;
    layer2_outputs(11384) <= a and not b;
    layer2_outputs(11385) <= '1';
    layer2_outputs(11386) <= not b;
    layer2_outputs(11387) <= not a;
    layer2_outputs(11388) <= not b or a;
    layer2_outputs(11389) <= '1';
    layer2_outputs(11390) <= not b;
    layer2_outputs(11391) <= not (a and b);
    layer2_outputs(11392) <= not a;
    layer2_outputs(11393) <= b and not a;
    layer2_outputs(11394) <= not (a and b);
    layer2_outputs(11395) <= a and not b;
    layer2_outputs(11396) <= a and b;
    layer2_outputs(11397) <= b;
    layer2_outputs(11398) <= not b;
    layer2_outputs(11399) <= not (a or b);
    layer2_outputs(11400) <= not a or b;
    layer2_outputs(11401) <= a xor b;
    layer2_outputs(11402) <= not a;
    layer2_outputs(11403) <= not b;
    layer2_outputs(11404) <= not b;
    layer2_outputs(11405) <= b and not a;
    layer2_outputs(11406) <= '1';
    layer2_outputs(11407) <= a or b;
    layer2_outputs(11408) <= not b;
    layer2_outputs(11409) <= a and b;
    layer2_outputs(11410) <= not (a or b);
    layer2_outputs(11411) <= b and not a;
    layer2_outputs(11412) <= not b;
    layer2_outputs(11413) <= a or b;
    layer2_outputs(11414) <= not b;
    layer2_outputs(11415) <= a and b;
    layer2_outputs(11416) <= a and not b;
    layer2_outputs(11417) <= b and not a;
    layer2_outputs(11418) <= '1';
    layer2_outputs(11419) <= b;
    layer2_outputs(11420) <= b;
    layer2_outputs(11421) <= '0';
    layer2_outputs(11422) <= not a;
    layer2_outputs(11423) <= a or b;
    layer2_outputs(11424) <= a and not b;
    layer2_outputs(11425) <= a;
    layer2_outputs(11426) <= not (a xor b);
    layer2_outputs(11427) <= a or b;
    layer2_outputs(11428) <= a or b;
    layer2_outputs(11429) <= a and b;
    layer2_outputs(11430) <= b and not a;
    layer2_outputs(11431) <= not a;
    layer2_outputs(11432) <= b;
    layer2_outputs(11433) <= a;
    layer2_outputs(11434) <= not (a and b);
    layer2_outputs(11435) <= not b or a;
    layer2_outputs(11436) <= not b;
    layer2_outputs(11437) <= a xor b;
    layer2_outputs(11438) <= not (a and b);
    layer2_outputs(11439) <= not (a and b);
    layer2_outputs(11440) <= a xor b;
    layer2_outputs(11441) <= '0';
    layer2_outputs(11442) <= a xor b;
    layer2_outputs(11443) <= not (a or b);
    layer2_outputs(11444) <= not a;
    layer2_outputs(11445) <= a and not b;
    layer2_outputs(11446) <= not a;
    layer2_outputs(11447) <= '1';
    layer2_outputs(11448) <= not b;
    layer2_outputs(11449) <= not b;
    layer2_outputs(11450) <= not (a or b);
    layer2_outputs(11451) <= a or b;
    layer2_outputs(11452) <= a;
    layer2_outputs(11453) <= not b or a;
    layer2_outputs(11454) <= b;
    layer2_outputs(11455) <= not (a xor b);
    layer2_outputs(11456) <= a;
    layer2_outputs(11457) <= a;
    layer2_outputs(11458) <= not b;
    layer2_outputs(11459) <= not (a or b);
    layer2_outputs(11460) <= not a;
    layer2_outputs(11461) <= b and not a;
    layer2_outputs(11462) <= a and not b;
    layer2_outputs(11463) <= not (a and b);
    layer2_outputs(11464) <= not a;
    layer2_outputs(11465) <= b and not a;
    layer2_outputs(11466) <= not (a and b);
    layer2_outputs(11467) <= a and b;
    layer2_outputs(11468) <= a;
    layer2_outputs(11469) <= '0';
    layer2_outputs(11470) <= not a;
    layer2_outputs(11471) <= a and not b;
    layer2_outputs(11472) <= '0';
    layer2_outputs(11473) <= a and b;
    layer2_outputs(11474) <= not (a or b);
    layer2_outputs(11475) <= b;
    layer2_outputs(11476) <= '1';
    layer2_outputs(11477) <= b;
    layer2_outputs(11478) <= not b or a;
    layer2_outputs(11479) <= a or b;
    layer2_outputs(11480) <= a;
    layer2_outputs(11481) <= not b or a;
    layer2_outputs(11482) <= not a or b;
    layer2_outputs(11483) <= '0';
    layer2_outputs(11484) <= a;
    layer2_outputs(11485) <= not b;
    layer2_outputs(11486) <= '1';
    layer2_outputs(11487) <= a and b;
    layer2_outputs(11488) <= b and not a;
    layer2_outputs(11489) <= not (a or b);
    layer2_outputs(11490) <= b and not a;
    layer2_outputs(11491) <= a and b;
    layer2_outputs(11492) <= b;
    layer2_outputs(11493) <= a or b;
    layer2_outputs(11494) <= a and not b;
    layer2_outputs(11495) <= not a or b;
    layer2_outputs(11496) <= not a;
    layer2_outputs(11497) <= not a;
    layer2_outputs(11498) <= not (a and b);
    layer2_outputs(11499) <= a;
    layer2_outputs(11500) <= a and b;
    layer2_outputs(11501) <= a and not b;
    layer2_outputs(11502) <= not b;
    layer2_outputs(11503) <= not b or a;
    layer2_outputs(11504) <= b and not a;
    layer2_outputs(11505) <= b;
    layer2_outputs(11506) <= a and b;
    layer2_outputs(11507) <= not a;
    layer2_outputs(11508) <= a and b;
    layer2_outputs(11509) <= not (a or b);
    layer2_outputs(11510) <= not b or a;
    layer2_outputs(11511) <= a;
    layer2_outputs(11512) <= a or b;
    layer2_outputs(11513) <= '0';
    layer2_outputs(11514) <= a and b;
    layer2_outputs(11515) <= b;
    layer2_outputs(11516) <= b;
    layer2_outputs(11517) <= a xor b;
    layer2_outputs(11518) <= not b;
    layer2_outputs(11519) <= not (a or b);
    layer2_outputs(11520) <= a and not b;
    layer2_outputs(11521) <= a;
    layer2_outputs(11522) <= a;
    layer2_outputs(11523) <= not (a and b);
    layer2_outputs(11524) <= a;
    layer2_outputs(11525) <= not a;
    layer2_outputs(11526) <= b and not a;
    layer2_outputs(11527) <= not a;
    layer2_outputs(11528) <= a;
    layer2_outputs(11529) <= b and not a;
    layer2_outputs(11530) <= not b;
    layer2_outputs(11531) <= a or b;
    layer2_outputs(11532) <= a and not b;
    layer2_outputs(11533) <= a;
    layer2_outputs(11534) <= not b or a;
    layer2_outputs(11535) <= not b;
    layer2_outputs(11536) <= '1';
    layer2_outputs(11537) <= not a or b;
    layer2_outputs(11538) <= a or b;
    layer2_outputs(11539) <= b;
    layer2_outputs(11540) <= '1';
    layer2_outputs(11541) <= not a or b;
    layer2_outputs(11542) <= not a;
    layer2_outputs(11543) <= a and not b;
    layer2_outputs(11544) <= a and b;
    layer2_outputs(11545) <= not b;
    layer2_outputs(11546) <= '1';
    layer2_outputs(11547) <= a;
    layer2_outputs(11548) <= a and not b;
    layer2_outputs(11549) <= b;
    layer2_outputs(11550) <= a xor b;
    layer2_outputs(11551) <= not a or b;
    layer2_outputs(11552) <= b;
    layer2_outputs(11553) <= a and b;
    layer2_outputs(11554) <= a xor b;
    layer2_outputs(11555) <= not (a xor b);
    layer2_outputs(11556) <= not a;
    layer2_outputs(11557) <= not b or a;
    layer2_outputs(11558) <= a and b;
    layer2_outputs(11559) <= not a;
    layer2_outputs(11560) <= not b or a;
    layer2_outputs(11561) <= not b or a;
    layer2_outputs(11562) <= not a or b;
    layer2_outputs(11563) <= a or b;
    layer2_outputs(11564) <= a and b;
    layer2_outputs(11565) <= not (a and b);
    layer2_outputs(11566) <= not b;
    layer2_outputs(11567) <= b;
    layer2_outputs(11568) <= not a or b;
    layer2_outputs(11569) <= a and not b;
    layer2_outputs(11570) <= b;
    layer2_outputs(11571) <= a and not b;
    layer2_outputs(11572) <= a;
    layer2_outputs(11573) <= not b;
    layer2_outputs(11574) <= not b;
    layer2_outputs(11575) <= a or b;
    layer2_outputs(11576) <= b;
    layer2_outputs(11577) <= not b;
    layer2_outputs(11578) <= not b;
    layer2_outputs(11579) <= b and not a;
    layer2_outputs(11580) <= not b or a;
    layer2_outputs(11581) <= not b;
    layer2_outputs(11582) <= not (a or b);
    layer2_outputs(11583) <= not a;
    layer2_outputs(11584) <= not b;
    layer2_outputs(11585) <= not a;
    layer2_outputs(11586) <= a or b;
    layer2_outputs(11587) <= not a;
    layer2_outputs(11588) <= not b;
    layer2_outputs(11589) <= not a;
    layer2_outputs(11590) <= not a or b;
    layer2_outputs(11591) <= '0';
    layer2_outputs(11592) <= not (a or b);
    layer2_outputs(11593) <= '1';
    layer2_outputs(11594) <= a or b;
    layer2_outputs(11595) <= not (a or b);
    layer2_outputs(11596) <= not (a xor b);
    layer2_outputs(11597) <= not b or a;
    layer2_outputs(11598) <= a;
    layer2_outputs(11599) <= not b;
    layer2_outputs(11600) <= not a or b;
    layer2_outputs(11601) <= not (a and b);
    layer2_outputs(11602) <= not a;
    layer2_outputs(11603) <= a;
    layer2_outputs(11604) <= a;
    layer2_outputs(11605) <= b and not a;
    layer2_outputs(11606) <= '1';
    layer2_outputs(11607) <= a;
    layer2_outputs(11608) <= '0';
    layer2_outputs(11609) <= not a;
    layer2_outputs(11610) <= a or b;
    layer2_outputs(11611) <= '1';
    layer2_outputs(11612) <= b;
    layer2_outputs(11613) <= not a;
    layer2_outputs(11614) <= not a;
    layer2_outputs(11615) <= not (a or b);
    layer2_outputs(11616) <= not a or b;
    layer2_outputs(11617) <= a and b;
    layer2_outputs(11618) <= '0';
    layer2_outputs(11619) <= not a or b;
    layer2_outputs(11620) <= '1';
    layer2_outputs(11621) <= '0';
    layer2_outputs(11622) <= not a;
    layer2_outputs(11623) <= not (a and b);
    layer2_outputs(11624) <= a or b;
    layer2_outputs(11625) <= not a;
    layer2_outputs(11626) <= not a or b;
    layer2_outputs(11627) <= a;
    layer2_outputs(11628) <= a or b;
    layer2_outputs(11629) <= not (a and b);
    layer2_outputs(11630) <= not a;
    layer2_outputs(11631) <= a and b;
    layer2_outputs(11632) <= b;
    layer2_outputs(11633) <= a or b;
    layer2_outputs(11634) <= a and b;
    layer2_outputs(11635) <= a and b;
    layer2_outputs(11636) <= not (a or b);
    layer2_outputs(11637) <= a or b;
    layer2_outputs(11638) <= not b;
    layer2_outputs(11639) <= not b or a;
    layer2_outputs(11640) <= a or b;
    layer2_outputs(11641) <= a;
    layer2_outputs(11642) <= a and not b;
    layer2_outputs(11643) <= not b;
    layer2_outputs(11644) <= a or b;
    layer2_outputs(11645) <= not b;
    layer2_outputs(11646) <= b and not a;
    layer2_outputs(11647) <= not a or b;
    layer2_outputs(11648) <= '1';
    layer2_outputs(11649) <= '1';
    layer2_outputs(11650) <= not (a or b);
    layer2_outputs(11651) <= a;
    layer2_outputs(11652) <= b and not a;
    layer2_outputs(11653) <= '1';
    layer2_outputs(11654) <= not a;
    layer2_outputs(11655) <= a and not b;
    layer2_outputs(11656) <= not a or b;
    layer2_outputs(11657) <= b;
    layer2_outputs(11658) <= not b;
    layer2_outputs(11659) <= not a;
    layer2_outputs(11660) <= not a;
    layer2_outputs(11661) <= a xor b;
    layer2_outputs(11662) <= a and not b;
    layer2_outputs(11663) <= a and b;
    layer2_outputs(11664) <= not b;
    layer2_outputs(11665) <= '0';
    layer2_outputs(11666) <= not (a xor b);
    layer2_outputs(11667) <= a and not b;
    layer2_outputs(11668) <= not (a and b);
    layer2_outputs(11669) <= not (a and b);
    layer2_outputs(11670) <= a and b;
    layer2_outputs(11671) <= not (a and b);
    layer2_outputs(11672) <= b and not a;
    layer2_outputs(11673) <= not b or a;
    layer2_outputs(11674) <= not b or a;
    layer2_outputs(11675) <= b;
    layer2_outputs(11676) <= a;
    layer2_outputs(11677) <= a and b;
    layer2_outputs(11678) <= not (a xor b);
    layer2_outputs(11679) <= not a;
    layer2_outputs(11680) <= not (a xor b);
    layer2_outputs(11681) <= a;
    layer2_outputs(11682) <= not b;
    layer2_outputs(11683) <= a and not b;
    layer2_outputs(11684) <= b;
    layer2_outputs(11685) <= a;
    layer2_outputs(11686) <= not b;
    layer2_outputs(11687) <= not (a or b);
    layer2_outputs(11688) <= '0';
    layer2_outputs(11689) <= a;
    layer2_outputs(11690) <= a;
    layer2_outputs(11691) <= a;
    layer2_outputs(11692) <= not b;
    layer2_outputs(11693) <= '0';
    layer2_outputs(11694) <= not a or b;
    layer2_outputs(11695) <= not a or b;
    layer2_outputs(11696) <= a or b;
    layer2_outputs(11697) <= not a or b;
    layer2_outputs(11698) <= b and not a;
    layer2_outputs(11699) <= a and not b;
    layer2_outputs(11700) <= a and b;
    layer2_outputs(11701) <= '0';
    layer2_outputs(11702) <= not a or b;
    layer2_outputs(11703) <= b;
    layer2_outputs(11704) <= '0';
    layer2_outputs(11705) <= not (a or b);
    layer2_outputs(11706) <= not (a xor b);
    layer2_outputs(11707) <= b;
    layer2_outputs(11708) <= b;
    layer2_outputs(11709) <= not a or b;
    layer2_outputs(11710) <= a;
    layer2_outputs(11711) <= not (a and b);
    layer2_outputs(11712) <= not a or b;
    layer2_outputs(11713) <= a xor b;
    layer2_outputs(11714) <= not a or b;
    layer2_outputs(11715) <= b;
    layer2_outputs(11716) <= '1';
    layer2_outputs(11717) <= a or b;
    layer2_outputs(11718) <= not b or a;
    layer2_outputs(11719) <= not a or b;
    layer2_outputs(11720) <= not (a and b);
    layer2_outputs(11721) <= a and not b;
    layer2_outputs(11722) <= not a;
    layer2_outputs(11723) <= '1';
    layer2_outputs(11724) <= a xor b;
    layer2_outputs(11725) <= a or b;
    layer2_outputs(11726) <= '1';
    layer2_outputs(11727) <= '1';
    layer2_outputs(11728) <= a and b;
    layer2_outputs(11729) <= b and not a;
    layer2_outputs(11730) <= a and b;
    layer2_outputs(11731) <= not b;
    layer2_outputs(11732) <= a xor b;
    layer2_outputs(11733) <= a;
    layer2_outputs(11734) <= not (a and b);
    layer2_outputs(11735) <= not a;
    layer2_outputs(11736) <= not a or b;
    layer2_outputs(11737) <= not (a or b);
    layer2_outputs(11738) <= a or b;
    layer2_outputs(11739) <= '0';
    layer2_outputs(11740) <= not b;
    layer2_outputs(11741) <= not b;
    layer2_outputs(11742) <= a xor b;
    layer2_outputs(11743) <= b and not a;
    layer2_outputs(11744) <= not (a or b);
    layer2_outputs(11745) <= a;
    layer2_outputs(11746) <= a xor b;
    layer2_outputs(11747) <= '0';
    layer2_outputs(11748) <= not b or a;
    layer2_outputs(11749) <= not b;
    layer2_outputs(11750) <= '1';
    layer2_outputs(11751) <= b;
    layer2_outputs(11752) <= a;
    layer2_outputs(11753) <= a and not b;
    layer2_outputs(11754) <= not b;
    layer2_outputs(11755) <= not a or b;
    layer2_outputs(11756) <= a and b;
    layer2_outputs(11757) <= b;
    layer2_outputs(11758) <= not a;
    layer2_outputs(11759) <= not b;
    layer2_outputs(11760) <= a;
    layer2_outputs(11761) <= not a or b;
    layer2_outputs(11762) <= a and b;
    layer2_outputs(11763) <= a and not b;
    layer2_outputs(11764) <= '0';
    layer2_outputs(11765) <= not a or b;
    layer2_outputs(11766) <= b and not a;
    layer2_outputs(11767) <= not a;
    layer2_outputs(11768) <= not a;
    layer2_outputs(11769) <= b and not a;
    layer2_outputs(11770) <= not a;
    layer2_outputs(11771) <= not a;
    layer2_outputs(11772) <= not (a xor b);
    layer2_outputs(11773) <= not b or a;
    layer2_outputs(11774) <= a or b;
    layer2_outputs(11775) <= not b or a;
    layer2_outputs(11776) <= a and not b;
    layer2_outputs(11777) <= a and b;
    layer2_outputs(11778) <= not (a or b);
    layer2_outputs(11779) <= a and not b;
    layer2_outputs(11780) <= '1';
    layer2_outputs(11781) <= b;
    layer2_outputs(11782) <= a xor b;
    layer2_outputs(11783) <= not (a or b);
    layer2_outputs(11784) <= a or b;
    layer2_outputs(11785) <= b;
    layer2_outputs(11786) <= a;
    layer2_outputs(11787) <= not (a or b);
    layer2_outputs(11788) <= a;
    layer2_outputs(11789) <= a;
    layer2_outputs(11790) <= not (a and b);
    layer2_outputs(11791) <= not (a and b);
    layer2_outputs(11792) <= a or b;
    layer2_outputs(11793) <= '1';
    layer2_outputs(11794) <= a;
    layer2_outputs(11795) <= a and not b;
    layer2_outputs(11796) <= not b;
    layer2_outputs(11797) <= a and b;
    layer2_outputs(11798) <= not a;
    layer2_outputs(11799) <= not a or b;
    layer2_outputs(11800) <= not (a or b);
    layer2_outputs(11801) <= b and not a;
    layer2_outputs(11802) <= b;
    layer2_outputs(11803) <= b;
    layer2_outputs(11804) <= not b;
    layer2_outputs(11805) <= b;
    layer2_outputs(11806) <= not b;
    layer2_outputs(11807) <= a and not b;
    layer2_outputs(11808) <= a;
    layer2_outputs(11809) <= b;
    layer2_outputs(11810) <= a and not b;
    layer2_outputs(11811) <= a or b;
    layer2_outputs(11812) <= not a;
    layer2_outputs(11813) <= not (a or b);
    layer2_outputs(11814) <= not (a or b);
    layer2_outputs(11815) <= not a;
    layer2_outputs(11816) <= not (a xor b);
    layer2_outputs(11817) <= a and not b;
    layer2_outputs(11818) <= a xor b;
    layer2_outputs(11819) <= '0';
    layer2_outputs(11820) <= a and b;
    layer2_outputs(11821) <= not a or b;
    layer2_outputs(11822) <= a and not b;
    layer2_outputs(11823) <= '0';
    layer2_outputs(11824) <= not b or a;
    layer2_outputs(11825) <= '1';
    layer2_outputs(11826) <= a xor b;
    layer2_outputs(11827) <= a;
    layer2_outputs(11828) <= not a;
    layer2_outputs(11829) <= b;
    layer2_outputs(11830) <= b;
    layer2_outputs(11831) <= not a or b;
    layer2_outputs(11832) <= a and not b;
    layer2_outputs(11833) <= not b;
    layer2_outputs(11834) <= not b or a;
    layer2_outputs(11835) <= not b;
    layer2_outputs(11836) <= a xor b;
    layer2_outputs(11837) <= not b;
    layer2_outputs(11838) <= not a;
    layer2_outputs(11839) <= b;
    layer2_outputs(11840) <= not (a or b);
    layer2_outputs(11841) <= not (a or b);
    layer2_outputs(11842) <= not a or b;
    layer2_outputs(11843) <= a xor b;
    layer2_outputs(11844) <= not (a or b);
    layer2_outputs(11845) <= a and not b;
    layer2_outputs(11846) <= a and not b;
    layer2_outputs(11847) <= a or b;
    layer2_outputs(11848) <= not b;
    layer2_outputs(11849) <= a or b;
    layer2_outputs(11850) <= a or b;
    layer2_outputs(11851) <= not b;
    layer2_outputs(11852) <= '0';
    layer2_outputs(11853) <= '0';
    layer2_outputs(11854) <= a and b;
    layer2_outputs(11855) <= a or b;
    layer2_outputs(11856) <= a;
    layer2_outputs(11857) <= not b or a;
    layer2_outputs(11858) <= not (a and b);
    layer2_outputs(11859) <= not a;
    layer2_outputs(11860) <= not (a and b);
    layer2_outputs(11861) <= not a;
    layer2_outputs(11862) <= not b;
    layer2_outputs(11863) <= not b;
    layer2_outputs(11864) <= a and not b;
    layer2_outputs(11865) <= '1';
    layer2_outputs(11866) <= not b or a;
    layer2_outputs(11867) <= a and b;
    layer2_outputs(11868) <= a;
    layer2_outputs(11869) <= b and not a;
    layer2_outputs(11870) <= not b;
    layer2_outputs(11871) <= not (a or b);
    layer2_outputs(11872) <= not b or a;
    layer2_outputs(11873) <= a and not b;
    layer2_outputs(11874) <= a and not b;
    layer2_outputs(11875) <= not (a xor b);
    layer2_outputs(11876) <= a;
    layer2_outputs(11877) <= a and not b;
    layer2_outputs(11878) <= a or b;
    layer2_outputs(11879) <= a or b;
    layer2_outputs(11880) <= b;
    layer2_outputs(11881) <= not b;
    layer2_outputs(11882) <= '0';
    layer2_outputs(11883) <= a and not b;
    layer2_outputs(11884) <= not a;
    layer2_outputs(11885) <= not a;
    layer2_outputs(11886) <= not (a or b);
    layer2_outputs(11887) <= not (a and b);
    layer2_outputs(11888) <= a or b;
    layer2_outputs(11889) <= a and b;
    layer2_outputs(11890) <= not (a and b);
    layer2_outputs(11891) <= a xor b;
    layer2_outputs(11892) <= a or b;
    layer2_outputs(11893) <= not (a and b);
    layer2_outputs(11894) <= a and b;
    layer2_outputs(11895) <= a and b;
    layer2_outputs(11896) <= b and not a;
    layer2_outputs(11897) <= '1';
    layer2_outputs(11898) <= not a;
    layer2_outputs(11899) <= a or b;
    layer2_outputs(11900) <= a and b;
    layer2_outputs(11901) <= not a;
    layer2_outputs(11902) <= not (a xor b);
    layer2_outputs(11903) <= not (a xor b);
    layer2_outputs(11904) <= b;
    layer2_outputs(11905) <= not a;
    layer2_outputs(11906) <= not b;
    layer2_outputs(11907) <= b;
    layer2_outputs(11908) <= not a;
    layer2_outputs(11909) <= '0';
    layer2_outputs(11910) <= a or b;
    layer2_outputs(11911) <= a or b;
    layer2_outputs(11912) <= '0';
    layer2_outputs(11913) <= a;
    layer2_outputs(11914) <= a and not b;
    layer2_outputs(11915) <= not b;
    layer2_outputs(11916) <= not (a xor b);
    layer2_outputs(11917) <= a or b;
    layer2_outputs(11918) <= '1';
    layer2_outputs(11919) <= not (a and b);
    layer2_outputs(11920) <= a;
    layer2_outputs(11921) <= not b or a;
    layer2_outputs(11922) <= not a or b;
    layer2_outputs(11923) <= not a or b;
    layer2_outputs(11924) <= not b;
    layer2_outputs(11925) <= '1';
    layer2_outputs(11926) <= a and not b;
    layer2_outputs(11927) <= a;
    layer2_outputs(11928) <= a xor b;
    layer2_outputs(11929) <= not b;
    layer2_outputs(11930) <= a and b;
    layer2_outputs(11931) <= b;
    layer2_outputs(11932) <= not a or b;
    layer2_outputs(11933) <= not (a or b);
    layer2_outputs(11934) <= a and b;
    layer2_outputs(11935) <= not (a and b);
    layer2_outputs(11936) <= not a or b;
    layer2_outputs(11937) <= not b;
    layer2_outputs(11938) <= not b or a;
    layer2_outputs(11939) <= b and not a;
    layer2_outputs(11940) <= b;
    layer2_outputs(11941) <= a and not b;
    layer2_outputs(11942) <= not a or b;
    layer2_outputs(11943) <= not (a or b);
    layer2_outputs(11944) <= a;
    layer2_outputs(11945) <= not a;
    layer2_outputs(11946) <= '1';
    layer2_outputs(11947) <= '1';
    layer2_outputs(11948) <= b;
    layer2_outputs(11949) <= a;
    layer2_outputs(11950) <= a;
    layer2_outputs(11951) <= b and not a;
    layer2_outputs(11952) <= b and not a;
    layer2_outputs(11953) <= '0';
    layer2_outputs(11954) <= a;
    layer2_outputs(11955) <= not b;
    layer2_outputs(11956) <= a or b;
    layer2_outputs(11957) <= not b or a;
    layer2_outputs(11958) <= a or b;
    layer2_outputs(11959) <= a and b;
    layer2_outputs(11960) <= not (a or b);
    layer2_outputs(11961) <= b and not a;
    layer2_outputs(11962) <= not a or b;
    layer2_outputs(11963) <= a xor b;
    layer2_outputs(11964) <= a and not b;
    layer2_outputs(11965) <= not (a or b);
    layer2_outputs(11966) <= not b or a;
    layer2_outputs(11967) <= a or b;
    layer2_outputs(11968) <= not (a and b);
    layer2_outputs(11969) <= not (a and b);
    layer2_outputs(11970) <= a;
    layer2_outputs(11971) <= not b;
    layer2_outputs(11972) <= a xor b;
    layer2_outputs(11973) <= not a;
    layer2_outputs(11974) <= not (a or b);
    layer2_outputs(11975) <= a and not b;
    layer2_outputs(11976) <= a xor b;
    layer2_outputs(11977) <= a or b;
    layer2_outputs(11978) <= '0';
    layer2_outputs(11979) <= a;
    layer2_outputs(11980) <= '0';
    layer2_outputs(11981) <= a xor b;
    layer2_outputs(11982) <= b;
    layer2_outputs(11983) <= not a;
    layer2_outputs(11984) <= not b;
    layer2_outputs(11985) <= not (a or b);
    layer2_outputs(11986) <= not b;
    layer2_outputs(11987) <= not (a or b);
    layer2_outputs(11988) <= a and not b;
    layer2_outputs(11989) <= not (a and b);
    layer2_outputs(11990) <= '1';
    layer2_outputs(11991) <= b;
    layer2_outputs(11992) <= not a or b;
    layer2_outputs(11993) <= not (a or b);
    layer2_outputs(11994) <= not (a and b);
    layer2_outputs(11995) <= not b or a;
    layer2_outputs(11996) <= a;
    layer2_outputs(11997) <= b;
    layer2_outputs(11998) <= not a;
    layer2_outputs(11999) <= a and b;
    layer2_outputs(12000) <= a;
    layer2_outputs(12001) <= a or b;
    layer2_outputs(12002) <= not (a and b);
    layer2_outputs(12003) <= not a;
    layer2_outputs(12004) <= a;
    layer2_outputs(12005) <= not (a or b);
    layer2_outputs(12006) <= a and not b;
    layer2_outputs(12007) <= '0';
    layer2_outputs(12008) <= a;
    layer2_outputs(12009) <= a and not b;
    layer2_outputs(12010) <= not a;
    layer2_outputs(12011) <= '1';
    layer2_outputs(12012) <= b;
    layer2_outputs(12013) <= not (a xor b);
    layer2_outputs(12014) <= not a;
    layer2_outputs(12015) <= not a;
    layer2_outputs(12016) <= a xor b;
    layer2_outputs(12017) <= '0';
    layer2_outputs(12018) <= a xor b;
    layer2_outputs(12019) <= '0';
    layer2_outputs(12020) <= a and not b;
    layer2_outputs(12021) <= not b or a;
    layer2_outputs(12022) <= not a;
    layer2_outputs(12023) <= not b;
    layer2_outputs(12024) <= a;
    layer2_outputs(12025) <= not (a xor b);
    layer2_outputs(12026) <= not a;
    layer2_outputs(12027) <= a and not b;
    layer2_outputs(12028) <= b;
    layer2_outputs(12029) <= not (a xor b);
    layer2_outputs(12030) <= b;
    layer2_outputs(12031) <= not (a and b);
    layer2_outputs(12032) <= not (a and b);
    layer2_outputs(12033) <= not (a and b);
    layer2_outputs(12034) <= a;
    layer2_outputs(12035) <= not b;
    layer2_outputs(12036) <= not b;
    layer2_outputs(12037) <= b and not a;
    layer2_outputs(12038) <= not a or b;
    layer2_outputs(12039) <= not a or b;
    layer2_outputs(12040) <= not a;
    layer2_outputs(12041) <= not b;
    layer2_outputs(12042) <= a or b;
    layer2_outputs(12043) <= b;
    layer2_outputs(12044) <= a and b;
    layer2_outputs(12045) <= not a or b;
    layer2_outputs(12046) <= b;
    layer2_outputs(12047) <= b;
    layer2_outputs(12048) <= a and b;
    layer2_outputs(12049) <= '0';
    layer2_outputs(12050) <= b and not a;
    layer2_outputs(12051) <= not (a xor b);
    layer2_outputs(12052) <= not (a or b);
    layer2_outputs(12053) <= '0';
    layer2_outputs(12054) <= a and not b;
    layer2_outputs(12055) <= a or b;
    layer2_outputs(12056) <= not (a or b);
    layer2_outputs(12057) <= a xor b;
    layer2_outputs(12058) <= not (a xor b);
    layer2_outputs(12059) <= not b;
    layer2_outputs(12060) <= b;
    layer2_outputs(12061) <= a;
    layer2_outputs(12062) <= a xor b;
    layer2_outputs(12063) <= a;
    layer2_outputs(12064) <= '1';
    layer2_outputs(12065) <= not b;
    layer2_outputs(12066) <= not (a or b);
    layer2_outputs(12067) <= not (a and b);
    layer2_outputs(12068) <= not (a or b);
    layer2_outputs(12069) <= not (a or b);
    layer2_outputs(12070) <= '0';
    layer2_outputs(12071) <= a or b;
    layer2_outputs(12072) <= not a;
    layer2_outputs(12073) <= a or b;
    layer2_outputs(12074) <= not (a or b);
    layer2_outputs(12075) <= not (a and b);
    layer2_outputs(12076) <= b;
    layer2_outputs(12077) <= a xor b;
    layer2_outputs(12078) <= not (a or b);
    layer2_outputs(12079) <= b;
    layer2_outputs(12080) <= not (a and b);
    layer2_outputs(12081) <= not (a or b);
    layer2_outputs(12082) <= a and b;
    layer2_outputs(12083) <= not b;
    layer2_outputs(12084) <= '0';
    layer2_outputs(12085) <= not (a and b);
    layer2_outputs(12086) <= not a or b;
    layer2_outputs(12087) <= a;
    layer2_outputs(12088) <= a or b;
    layer2_outputs(12089) <= not (a or b);
    layer2_outputs(12090) <= '1';
    layer2_outputs(12091) <= not (a and b);
    layer2_outputs(12092) <= not a;
    layer2_outputs(12093) <= not b;
    layer2_outputs(12094) <= not a or b;
    layer2_outputs(12095) <= b;
    layer2_outputs(12096) <= not a or b;
    layer2_outputs(12097) <= not (a or b);
    layer2_outputs(12098) <= a;
    layer2_outputs(12099) <= a;
    layer2_outputs(12100) <= a xor b;
    layer2_outputs(12101) <= '1';
    layer2_outputs(12102) <= a and not b;
    layer2_outputs(12103) <= not b;
    layer2_outputs(12104) <= b;
    layer2_outputs(12105) <= not (a and b);
    layer2_outputs(12106) <= '0';
    layer2_outputs(12107) <= not (a xor b);
    layer2_outputs(12108) <= a;
    layer2_outputs(12109) <= '0';
    layer2_outputs(12110) <= a and b;
    layer2_outputs(12111) <= not b;
    layer2_outputs(12112) <= b and not a;
    layer2_outputs(12113) <= a;
    layer2_outputs(12114) <= not b or a;
    layer2_outputs(12115) <= b and not a;
    layer2_outputs(12116) <= a and not b;
    layer2_outputs(12117) <= a;
    layer2_outputs(12118) <= not (a and b);
    layer2_outputs(12119) <= not b;
    layer2_outputs(12120) <= '0';
    layer2_outputs(12121) <= not b or a;
    layer2_outputs(12122) <= not b or a;
    layer2_outputs(12123) <= not (a and b);
    layer2_outputs(12124) <= not (a or b);
    layer2_outputs(12125) <= b and not a;
    layer2_outputs(12126) <= a;
    layer2_outputs(12127) <= b;
    layer2_outputs(12128) <= not (a xor b);
    layer2_outputs(12129) <= not b;
    layer2_outputs(12130) <= not a or b;
    layer2_outputs(12131) <= a and b;
    layer2_outputs(12132) <= a or b;
    layer2_outputs(12133) <= not (a or b);
    layer2_outputs(12134) <= b;
    layer2_outputs(12135) <= '1';
    layer2_outputs(12136) <= not a;
    layer2_outputs(12137) <= a and b;
    layer2_outputs(12138) <= not b;
    layer2_outputs(12139) <= '1';
    layer2_outputs(12140) <= not (a xor b);
    layer2_outputs(12141) <= a or b;
    layer2_outputs(12142) <= not b;
    layer2_outputs(12143) <= a;
    layer2_outputs(12144) <= b;
    layer2_outputs(12145) <= a;
    layer2_outputs(12146) <= b;
    layer2_outputs(12147) <= not b or a;
    layer2_outputs(12148) <= a and b;
    layer2_outputs(12149) <= a and b;
    layer2_outputs(12150) <= not b or a;
    layer2_outputs(12151) <= a;
    layer2_outputs(12152) <= not (a and b);
    layer2_outputs(12153) <= not a;
    layer2_outputs(12154) <= not (a or b);
    layer2_outputs(12155) <= not (a and b);
    layer2_outputs(12156) <= not a or b;
    layer2_outputs(12157) <= a and not b;
    layer2_outputs(12158) <= not a;
    layer2_outputs(12159) <= not a or b;
    layer2_outputs(12160) <= not b or a;
    layer2_outputs(12161) <= a;
    layer2_outputs(12162) <= a and b;
    layer2_outputs(12163) <= a or b;
    layer2_outputs(12164) <= a;
    layer2_outputs(12165) <= not b or a;
    layer2_outputs(12166) <= not b;
    layer2_outputs(12167) <= a;
    layer2_outputs(12168) <= not a or b;
    layer2_outputs(12169) <= not (a xor b);
    layer2_outputs(12170) <= not b or a;
    layer2_outputs(12171) <= not b or a;
    layer2_outputs(12172) <= a and not b;
    layer2_outputs(12173) <= a and not b;
    layer2_outputs(12174) <= not b or a;
    layer2_outputs(12175) <= not a or b;
    layer2_outputs(12176) <= a xor b;
    layer2_outputs(12177) <= not b;
    layer2_outputs(12178) <= a or b;
    layer2_outputs(12179) <= not (a xor b);
    layer2_outputs(12180) <= not b or a;
    layer2_outputs(12181) <= a and not b;
    layer2_outputs(12182) <= not a;
    layer2_outputs(12183) <= a;
    layer2_outputs(12184) <= a;
    layer2_outputs(12185) <= b;
    layer2_outputs(12186) <= a and not b;
    layer2_outputs(12187) <= b;
    layer2_outputs(12188) <= a;
    layer2_outputs(12189) <= not b;
    layer2_outputs(12190) <= '1';
    layer2_outputs(12191) <= not (a and b);
    layer2_outputs(12192) <= not b;
    layer2_outputs(12193) <= a and b;
    layer2_outputs(12194) <= not b or a;
    layer2_outputs(12195) <= not a or b;
    layer2_outputs(12196) <= '0';
    layer2_outputs(12197) <= not (a xor b);
    layer2_outputs(12198) <= '0';
    layer2_outputs(12199) <= b and not a;
    layer2_outputs(12200) <= a xor b;
    layer2_outputs(12201) <= a and b;
    layer2_outputs(12202) <= not b or a;
    layer2_outputs(12203) <= not a;
    layer2_outputs(12204) <= a;
    layer2_outputs(12205) <= not b or a;
    layer2_outputs(12206) <= not a;
    layer2_outputs(12207) <= not (a or b);
    layer2_outputs(12208) <= not (a or b);
    layer2_outputs(12209) <= not (a or b);
    layer2_outputs(12210) <= '1';
    layer2_outputs(12211) <= b and not a;
    layer2_outputs(12212) <= a;
    layer2_outputs(12213) <= a and b;
    layer2_outputs(12214) <= a;
    layer2_outputs(12215) <= a and not b;
    layer2_outputs(12216) <= b;
    layer2_outputs(12217) <= a or b;
    layer2_outputs(12218) <= not (a or b);
    layer2_outputs(12219) <= b and not a;
    layer2_outputs(12220) <= b;
    layer2_outputs(12221) <= not a;
    layer2_outputs(12222) <= b and not a;
    layer2_outputs(12223) <= b;
    layer2_outputs(12224) <= not a;
    layer2_outputs(12225) <= '0';
    layer2_outputs(12226) <= a and b;
    layer2_outputs(12227) <= not b or a;
    layer2_outputs(12228) <= not a or b;
    layer2_outputs(12229) <= not (a or b);
    layer2_outputs(12230) <= not (a or b);
    layer2_outputs(12231) <= not b or a;
    layer2_outputs(12232) <= not a;
    layer2_outputs(12233) <= not b or a;
    layer2_outputs(12234) <= a or b;
    layer2_outputs(12235) <= a or b;
    layer2_outputs(12236) <= '0';
    layer2_outputs(12237) <= not b or a;
    layer2_outputs(12238) <= not b;
    layer2_outputs(12239) <= b and not a;
    layer2_outputs(12240) <= a;
    layer2_outputs(12241) <= a or b;
    layer2_outputs(12242) <= not a;
    layer2_outputs(12243) <= not (a and b);
    layer2_outputs(12244) <= b;
    layer2_outputs(12245) <= a and not b;
    layer2_outputs(12246) <= not (a and b);
    layer2_outputs(12247) <= a;
    layer2_outputs(12248) <= not (a and b);
    layer2_outputs(12249) <= '0';
    layer2_outputs(12250) <= b;
    layer2_outputs(12251) <= not a;
    layer2_outputs(12252) <= b;
    layer2_outputs(12253) <= '0';
    layer2_outputs(12254) <= a;
    layer2_outputs(12255) <= not b or a;
    layer2_outputs(12256) <= b and not a;
    layer2_outputs(12257) <= a or b;
    layer2_outputs(12258) <= not a;
    layer2_outputs(12259) <= '1';
    layer2_outputs(12260) <= a or b;
    layer2_outputs(12261) <= not (a and b);
    layer2_outputs(12262) <= b;
    layer2_outputs(12263) <= '1';
    layer2_outputs(12264) <= not a;
    layer2_outputs(12265) <= a or b;
    layer2_outputs(12266) <= a;
    layer2_outputs(12267) <= '1';
    layer2_outputs(12268) <= not (a xor b);
    layer2_outputs(12269) <= a;
    layer2_outputs(12270) <= a and not b;
    layer2_outputs(12271) <= a and not b;
    layer2_outputs(12272) <= not a or b;
    layer2_outputs(12273) <= not b;
    layer2_outputs(12274) <= not (a xor b);
    layer2_outputs(12275) <= not b;
    layer2_outputs(12276) <= b and not a;
    layer2_outputs(12277) <= not a;
    layer2_outputs(12278) <= not (a xor b);
    layer2_outputs(12279) <= b;
    layer2_outputs(12280) <= not b or a;
    layer2_outputs(12281) <= a or b;
    layer2_outputs(12282) <= not a or b;
    layer2_outputs(12283) <= not b or a;
    layer2_outputs(12284) <= not a or b;
    layer2_outputs(12285) <= '0';
    layer2_outputs(12286) <= not a;
    layer2_outputs(12287) <= not b;
    layer2_outputs(12288) <= not (a or b);
    layer2_outputs(12289) <= a xor b;
    layer2_outputs(12290) <= a or b;
    layer2_outputs(12291) <= '0';
    layer2_outputs(12292) <= '1';
    layer2_outputs(12293) <= b and not a;
    layer2_outputs(12294) <= a or b;
    layer2_outputs(12295) <= b and not a;
    layer2_outputs(12296) <= not (a and b);
    layer2_outputs(12297) <= a;
    layer2_outputs(12298) <= b;
    layer2_outputs(12299) <= a or b;
    layer2_outputs(12300) <= not a;
    layer2_outputs(12301) <= not b or a;
    layer2_outputs(12302) <= b and not a;
    layer2_outputs(12303) <= '0';
    layer2_outputs(12304) <= a;
    layer2_outputs(12305) <= a;
    layer2_outputs(12306) <= b and not a;
    layer2_outputs(12307) <= '0';
    layer2_outputs(12308) <= not (a or b);
    layer2_outputs(12309) <= not (a or b);
    layer2_outputs(12310) <= a xor b;
    layer2_outputs(12311) <= '0';
    layer2_outputs(12312) <= a and b;
    layer2_outputs(12313) <= not (a xor b);
    layer2_outputs(12314) <= a;
    layer2_outputs(12315) <= not b or a;
    layer2_outputs(12316) <= b;
    layer2_outputs(12317) <= not b;
    layer2_outputs(12318) <= not a;
    layer2_outputs(12319) <= b;
    layer2_outputs(12320) <= '1';
    layer2_outputs(12321) <= not b or a;
    layer2_outputs(12322) <= '1';
    layer2_outputs(12323) <= b and not a;
    layer2_outputs(12324) <= not (a or b);
    layer2_outputs(12325) <= b;
    layer2_outputs(12326) <= not b;
    layer2_outputs(12327) <= not (a and b);
    layer2_outputs(12328) <= '0';
    layer2_outputs(12329) <= b;
    layer2_outputs(12330) <= a;
    layer2_outputs(12331) <= not a;
    layer2_outputs(12332) <= not b;
    layer2_outputs(12333) <= not b;
    layer2_outputs(12334) <= b and not a;
    layer2_outputs(12335) <= not a;
    layer2_outputs(12336) <= not a or b;
    layer2_outputs(12337) <= not a;
    layer2_outputs(12338) <= a and b;
    layer2_outputs(12339) <= not b;
    layer2_outputs(12340) <= b and not a;
    layer2_outputs(12341) <= a and not b;
    layer2_outputs(12342) <= not a or b;
    layer2_outputs(12343) <= '0';
    layer2_outputs(12344) <= not a;
    layer2_outputs(12345) <= not b or a;
    layer2_outputs(12346) <= b and not a;
    layer2_outputs(12347) <= a and not b;
    layer2_outputs(12348) <= a;
    layer2_outputs(12349) <= '1';
    layer2_outputs(12350) <= b;
    layer2_outputs(12351) <= not (a or b);
    layer2_outputs(12352) <= not a;
    layer2_outputs(12353) <= b;
    layer2_outputs(12354) <= not (a and b);
    layer2_outputs(12355) <= b;
    layer2_outputs(12356) <= not (a or b);
    layer2_outputs(12357) <= not (a and b);
    layer2_outputs(12358) <= a or b;
    layer2_outputs(12359) <= '0';
    layer2_outputs(12360) <= a;
    layer2_outputs(12361) <= a and b;
    layer2_outputs(12362) <= a and not b;
    layer2_outputs(12363) <= a and b;
    layer2_outputs(12364) <= b and not a;
    layer2_outputs(12365) <= b and not a;
    layer2_outputs(12366) <= not (a or b);
    layer2_outputs(12367) <= b and not a;
    layer2_outputs(12368) <= '1';
    layer2_outputs(12369) <= not (a or b);
    layer2_outputs(12370) <= not a;
    layer2_outputs(12371) <= a;
    layer2_outputs(12372) <= not b;
    layer2_outputs(12373) <= not (a and b);
    layer2_outputs(12374) <= not b or a;
    layer2_outputs(12375) <= a or b;
    layer2_outputs(12376) <= not b;
    layer2_outputs(12377) <= '0';
    layer2_outputs(12378) <= b;
    layer2_outputs(12379) <= not b;
    layer2_outputs(12380) <= a or b;
    layer2_outputs(12381) <= a;
    layer2_outputs(12382) <= not a;
    layer2_outputs(12383) <= not b;
    layer2_outputs(12384) <= not b;
    layer2_outputs(12385) <= a and b;
    layer2_outputs(12386) <= '1';
    layer2_outputs(12387) <= not (a or b);
    layer2_outputs(12388) <= a;
    layer2_outputs(12389) <= not (a xor b);
    layer2_outputs(12390) <= a;
    layer2_outputs(12391) <= a or b;
    layer2_outputs(12392) <= a;
    layer2_outputs(12393) <= a and b;
    layer2_outputs(12394) <= b and not a;
    layer2_outputs(12395) <= not (a and b);
    layer2_outputs(12396) <= not a or b;
    layer2_outputs(12397) <= not (a and b);
    layer2_outputs(12398) <= a or b;
    layer2_outputs(12399) <= not (a and b);
    layer2_outputs(12400) <= not a;
    layer2_outputs(12401) <= not a or b;
    layer2_outputs(12402) <= a;
    layer2_outputs(12403) <= not b;
    layer2_outputs(12404) <= a;
    layer2_outputs(12405) <= b and not a;
    layer2_outputs(12406) <= '1';
    layer2_outputs(12407) <= not (a and b);
    layer2_outputs(12408) <= b;
    layer2_outputs(12409) <= '1';
    layer2_outputs(12410) <= not b;
    layer2_outputs(12411) <= not a;
    layer2_outputs(12412) <= a and b;
    layer2_outputs(12413) <= not (a or b);
    layer2_outputs(12414) <= a or b;
    layer2_outputs(12415) <= b;
    layer2_outputs(12416) <= a and not b;
    layer2_outputs(12417) <= not (a and b);
    layer2_outputs(12418) <= a;
    layer2_outputs(12419) <= a or b;
    layer2_outputs(12420) <= a and b;
    layer2_outputs(12421) <= not a;
    layer2_outputs(12422) <= not (a xor b);
    layer2_outputs(12423) <= a and b;
    layer2_outputs(12424) <= b and not a;
    layer2_outputs(12425) <= b;
    layer2_outputs(12426) <= not a or b;
    layer2_outputs(12427) <= a or b;
    layer2_outputs(12428) <= not (a or b);
    layer2_outputs(12429) <= a or b;
    layer2_outputs(12430) <= a;
    layer2_outputs(12431) <= '1';
    layer2_outputs(12432) <= not b or a;
    layer2_outputs(12433) <= not a or b;
    layer2_outputs(12434) <= a;
    layer2_outputs(12435) <= not (a and b);
    layer2_outputs(12436) <= a;
    layer2_outputs(12437) <= a;
    layer2_outputs(12438) <= a or b;
    layer2_outputs(12439) <= not (a and b);
    layer2_outputs(12440) <= not b or a;
    layer2_outputs(12441) <= not b;
    layer2_outputs(12442) <= b and not a;
    layer2_outputs(12443) <= not b;
    layer2_outputs(12444) <= b and not a;
    layer2_outputs(12445) <= a or b;
    layer2_outputs(12446) <= not b;
    layer2_outputs(12447) <= b;
    layer2_outputs(12448) <= a;
    layer2_outputs(12449) <= not a;
    layer2_outputs(12450) <= a or b;
    layer2_outputs(12451) <= not a;
    layer2_outputs(12452) <= a and b;
    layer2_outputs(12453) <= not (a or b);
    layer2_outputs(12454) <= a and b;
    layer2_outputs(12455) <= not a;
    layer2_outputs(12456) <= a;
    layer2_outputs(12457) <= a xor b;
    layer2_outputs(12458) <= b and not a;
    layer2_outputs(12459) <= not (a xor b);
    layer2_outputs(12460) <= not a;
    layer2_outputs(12461) <= not b or a;
    layer2_outputs(12462) <= a or b;
    layer2_outputs(12463) <= a and not b;
    layer2_outputs(12464) <= b and not a;
    layer2_outputs(12465) <= a and not b;
    layer2_outputs(12466) <= not (a or b);
    layer2_outputs(12467) <= not (a xor b);
    layer2_outputs(12468) <= a and b;
    layer2_outputs(12469) <= a and not b;
    layer2_outputs(12470) <= '1';
    layer2_outputs(12471) <= not a or b;
    layer2_outputs(12472) <= a;
    layer2_outputs(12473) <= not (a or b);
    layer2_outputs(12474) <= not b or a;
    layer2_outputs(12475) <= not a;
    layer2_outputs(12476) <= '0';
    layer2_outputs(12477) <= not (a xor b);
    layer2_outputs(12478) <= '1';
    layer2_outputs(12479) <= not (a or b);
    layer2_outputs(12480) <= a and b;
    layer2_outputs(12481) <= not (a or b);
    layer2_outputs(12482) <= not (a and b);
    layer2_outputs(12483) <= a and b;
    layer2_outputs(12484) <= a or b;
    layer2_outputs(12485) <= not b or a;
    layer2_outputs(12486) <= not b;
    layer2_outputs(12487) <= a and b;
    layer2_outputs(12488) <= not a;
    layer2_outputs(12489) <= not (a or b);
    layer2_outputs(12490) <= not a;
    layer2_outputs(12491) <= not (a xor b);
    layer2_outputs(12492) <= '1';
    layer2_outputs(12493) <= b;
    layer2_outputs(12494) <= not b;
    layer2_outputs(12495) <= not (a and b);
    layer2_outputs(12496) <= b and not a;
    layer2_outputs(12497) <= b;
    layer2_outputs(12498) <= a and not b;
    layer2_outputs(12499) <= a;
    layer2_outputs(12500) <= a and not b;
    layer2_outputs(12501) <= a and not b;
    layer2_outputs(12502) <= b;
    layer2_outputs(12503) <= '1';
    layer2_outputs(12504) <= not a;
    layer2_outputs(12505) <= '1';
    layer2_outputs(12506) <= b;
    layer2_outputs(12507) <= not a;
    layer2_outputs(12508) <= not a;
    layer2_outputs(12509) <= not (a and b);
    layer2_outputs(12510) <= '0';
    layer2_outputs(12511) <= not b or a;
    layer2_outputs(12512) <= a and not b;
    layer2_outputs(12513) <= b;
    layer2_outputs(12514) <= b and not a;
    layer2_outputs(12515) <= not b or a;
    layer2_outputs(12516) <= not b or a;
    layer2_outputs(12517) <= a and b;
    layer2_outputs(12518) <= not b or a;
    layer2_outputs(12519) <= not a;
    layer2_outputs(12520) <= not (a and b);
    layer2_outputs(12521) <= not a;
    layer2_outputs(12522) <= a xor b;
    layer2_outputs(12523) <= not b or a;
    layer2_outputs(12524) <= b and not a;
    layer2_outputs(12525) <= '0';
    layer2_outputs(12526) <= a and not b;
    layer2_outputs(12527) <= not (a or b);
    layer2_outputs(12528) <= not b or a;
    layer2_outputs(12529) <= '0';
    layer2_outputs(12530) <= '1';
    layer2_outputs(12531) <= a or b;
    layer2_outputs(12532) <= not a;
    layer2_outputs(12533) <= not a or b;
    layer2_outputs(12534) <= a and not b;
    layer2_outputs(12535) <= a and not b;
    layer2_outputs(12536) <= b;
    layer2_outputs(12537) <= not a;
    layer2_outputs(12538) <= a;
    layer2_outputs(12539) <= a and b;
    layer2_outputs(12540) <= not b;
    layer2_outputs(12541) <= '0';
    layer2_outputs(12542) <= a or b;
    layer2_outputs(12543) <= '0';
    layer2_outputs(12544) <= not b;
    layer2_outputs(12545) <= not a;
    layer2_outputs(12546) <= b and not a;
    layer2_outputs(12547) <= a or b;
    layer2_outputs(12548) <= b;
    layer2_outputs(12549) <= a and b;
    layer2_outputs(12550) <= a;
    layer2_outputs(12551) <= not (a or b);
    layer2_outputs(12552) <= '0';
    layer2_outputs(12553) <= b and not a;
    layer2_outputs(12554) <= not (a and b);
    layer2_outputs(12555) <= a and not b;
    layer2_outputs(12556) <= not b;
    layer2_outputs(12557) <= not (a or b);
    layer2_outputs(12558) <= a;
    layer2_outputs(12559) <= not (a xor b);
    layer2_outputs(12560) <= a;
    layer2_outputs(12561) <= not (a or b);
    layer2_outputs(12562) <= not a;
    layer2_outputs(12563) <= a;
    layer2_outputs(12564) <= b;
    layer2_outputs(12565) <= a and b;
    layer2_outputs(12566) <= not (a and b);
    layer2_outputs(12567) <= a and not b;
    layer2_outputs(12568) <= a and b;
    layer2_outputs(12569) <= '1';
    layer2_outputs(12570) <= a and not b;
    layer2_outputs(12571) <= not b or a;
    layer2_outputs(12572) <= not a;
    layer2_outputs(12573) <= a and not b;
    layer2_outputs(12574) <= not (a or b);
    layer2_outputs(12575) <= not a;
    layer2_outputs(12576) <= a xor b;
    layer2_outputs(12577) <= not a;
    layer2_outputs(12578) <= not (a or b);
    layer2_outputs(12579) <= not a or b;
    layer2_outputs(12580) <= a xor b;
    layer2_outputs(12581) <= not (a and b);
    layer2_outputs(12582) <= a and not b;
    layer2_outputs(12583) <= b and not a;
    layer2_outputs(12584) <= '1';
    layer2_outputs(12585) <= a xor b;
    layer2_outputs(12586) <= a;
    layer2_outputs(12587) <= not b;
    layer2_outputs(12588) <= not (a or b);
    layer2_outputs(12589) <= b;
    layer2_outputs(12590) <= a;
    layer2_outputs(12591) <= b;
    layer2_outputs(12592) <= '1';
    layer2_outputs(12593) <= not a or b;
    layer2_outputs(12594) <= a;
    layer2_outputs(12595) <= not a;
    layer2_outputs(12596) <= b;
    layer2_outputs(12597) <= a;
    layer2_outputs(12598) <= a and b;
    layer2_outputs(12599) <= a and b;
    layer2_outputs(12600) <= not b;
    layer2_outputs(12601) <= a and not b;
    layer2_outputs(12602) <= not a or b;
    layer2_outputs(12603) <= not (a or b);
    layer2_outputs(12604) <= a and b;
    layer2_outputs(12605) <= a xor b;
    layer2_outputs(12606) <= not b;
    layer2_outputs(12607) <= a xor b;
    layer2_outputs(12608) <= not (a xor b);
    layer2_outputs(12609) <= not b;
    layer2_outputs(12610) <= not (a or b);
    layer2_outputs(12611) <= not a or b;
    layer2_outputs(12612) <= not a;
    layer2_outputs(12613) <= a and not b;
    layer2_outputs(12614) <= a and b;
    layer2_outputs(12615) <= a;
    layer2_outputs(12616) <= not a or b;
    layer2_outputs(12617) <= a xor b;
    layer2_outputs(12618) <= a and not b;
    layer2_outputs(12619) <= not (a and b);
    layer2_outputs(12620) <= '1';
    layer2_outputs(12621) <= not (a xor b);
    layer2_outputs(12622) <= a;
    layer2_outputs(12623) <= b and not a;
    layer2_outputs(12624) <= a or b;
    layer2_outputs(12625) <= not a;
    layer2_outputs(12626) <= '1';
    layer2_outputs(12627) <= b;
    layer2_outputs(12628) <= not (a or b);
    layer2_outputs(12629) <= not (a and b);
    layer2_outputs(12630) <= not b;
    layer2_outputs(12631) <= not a;
    layer2_outputs(12632) <= a or b;
    layer2_outputs(12633) <= not a or b;
    layer2_outputs(12634) <= b;
    layer2_outputs(12635) <= not b;
    layer2_outputs(12636) <= b;
    layer2_outputs(12637) <= b and not a;
    layer2_outputs(12638) <= '1';
    layer2_outputs(12639) <= not (a or b);
    layer2_outputs(12640) <= not b or a;
    layer2_outputs(12641) <= a;
    layer2_outputs(12642) <= not b;
    layer2_outputs(12643) <= not (a and b);
    layer2_outputs(12644) <= not a or b;
    layer2_outputs(12645) <= not a;
    layer2_outputs(12646) <= not b or a;
    layer2_outputs(12647) <= a and not b;
    layer2_outputs(12648) <= a or b;
    layer2_outputs(12649) <= not (a or b);
    layer2_outputs(12650) <= a;
    layer2_outputs(12651) <= a;
    layer2_outputs(12652) <= a xor b;
    layer2_outputs(12653) <= not (a or b);
    layer2_outputs(12654) <= a and b;
    layer2_outputs(12655) <= '0';
    layer2_outputs(12656) <= a;
    layer2_outputs(12657) <= b and not a;
    layer2_outputs(12658) <= not (a xor b);
    layer2_outputs(12659) <= not b;
    layer2_outputs(12660) <= '0';
    layer2_outputs(12661) <= not a or b;
    layer2_outputs(12662) <= b and not a;
    layer2_outputs(12663) <= not a;
    layer2_outputs(12664) <= not a;
    layer2_outputs(12665) <= not (a and b);
    layer2_outputs(12666) <= not b or a;
    layer2_outputs(12667) <= '1';
    layer2_outputs(12668) <= not a or b;
    layer2_outputs(12669) <= a;
    layer2_outputs(12670) <= not a or b;
    layer2_outputs(12671) <= a;
    layer2_outputs(12672) <= a or b;
    layer2_outputs(12673) <= not b or a;
    layer2_outputs(12674) <= a;
    layer2_outputs(12675) <= b;
    layer2_outputs(12676) <= not (a and b);
    layer2_outputs(12677) <= a and b;
    layer2_outputs(12678) <= not b;
    layer2_outputs(12679) <= b;
    layer2_outputs(12680) <= not (a xor b);
    layer2_outputs(12681) <= a and not b;
    layer2_outputs(12682) <= a;
    layer2_outputs(12683) <= b and not a;
    layer2_outputs(12684) <= not b or a;
    layer2_outputs(12685) <= a and not b;
    layer2_outputs(12686) <= a and not b;
    layer2_outputs(12687) <= a and not b;
    layer2_outputs(12688) <= a;
    layer2_outputs(12689) <= not a;
    layer2_outputs(12690) <= a and b;
    layer2_outputs(12691) <= a;
    layer2_outputs(12692) <= a xor b;
    layer2_outputs(12693) <= '1';
    layer2_outputs(12694) <= '1';
    layer2_outputs(12695) <= b and not a;
    layer2_outputs(12696) <= not a or b;
    layer2_outputs(12697) <= not (a and b);
    layer2_outputs(12698) <= not a;
    layer2_outputs(12699) <= '0';
    layer2_outputs(12700) <= a and b;
    layer2_outputs(12701) <= not a;
    layer2_outputs(12702) <= a and not b;
    layer2_outputs(12703) <= b;
    layer2_outputs(12704) <= a xor b;
    layer2_outputs(12705) <= a;
    layer2_outputs(12706) <= not b;
    layer2_outputs(12707) <= not b;
    layer2_outputs(12708) <= b;
    layer2_outputs(12709) <= not b;
    layer2_outputs(12710) <= not a or b;
    layer2_outputs(12711) <= b;
    layer2_outputs(12712) <= b;
    layer2_outputs(12713) <= a and not b;
    layer2_outputs(12714) <= not a;
    layer2_outputs(12715) <= not (a and b);
    layer2_outputs(12716) <= a and b;
    layer2_outputs(12717) <= not (a or b);
    layer2_outputs(12718) <= '0';
    layer2_outputs(12719) <= not (a or b);
    layer2_outputs(12720) <= not b or a;
    layer2_outputs(12721) <= a;
    layer2_outputs(12722) <= not b;
    layer2_outputs(12723) <= a or b;
    layer2_outputs(12724) <= a xor b;
    layer2_outputs(12725) <= not b;
    layer2_outputs(12726) <= not b or a;
    layer2_outputs(12727) <= a and not b;
    layer2_outputs(12728) <= not (a or b);
    layer2_outputs(12729) <= not (a or b);
    layer2_outputs(12730) <= not (a or b);
    layer2_outputs(12731) <= not b;
    layer2_outputs(12732) <= a and b;
    layer2_outputs(12733) <= not (a and b);
    layer2_outputs(12734) <= '0';
    layer2_outputs(12735) <= a and b;
    layer2_outputs(12736) <= a;
    layer2_outputs(12737) <= a and b;
    layer2_outputs(12738) <= not b or a;
    layer2_outputs(12739) <= not b;
    layer2_outputs(12740) <= a;
    layer2_outputs(12741) <= not (a xor b);
    layer2_outputs(12742) <= a or b;
    layer2_outputs(12743) <= a or b;
    layer2_outputs(12744) <= a and not b;
    layer2_outputs(12745) <= not (a xor b);
    layer2_outputs(12746) <= b;
    layer2_outputs(12747) <= b;
    layer2_outputs(12748) <= a or b;
    layer2_outputs(12749) <= a;
    layer2_outputs(12750) <= '1';
    layer2_outputs(12751) <= '0';
    layer2_outputs(12752) <= not (a xor b);
    layer2_outputs(12753) <= not (a or b);
    layer2_outputs(12754) <= a or b;
    layer2_outputs(12755) <= not (a xor b);
    layer2_outputs(12756) <= b;
    layer2_outputs(12757) <= b;
    layer2_outputs(12758) <= a;
    layer2_outputs(12759) <= not (a and b);
    layer2_outputs(12760) <= a and not b;
    layer2_outputs(12761) <= a;
    layer2_outputs(12762) <= b and not a;
    layer2_outputs(12763) <= not b;
    layer2_outputs(12764) <= not b;
    layer2_outputs(12765) <= not (a or b);
    layer2_outputs(12766) <= not (a or b);
    layer2_outputs(12767) <= a or b;
    layer2_outputs(12768) <= b;
    layer2_outputs(12769) <= not a;
    layer2_outputs(12770) <= not (a or b);
    layer2_outputs(12771) <= not a;
    layer2_outputs(12772) <= b and not a;
    layer2_outputs(12773) <= not (a or b);
    layer2_outputs(12774) <= a and not b;
    layer2_outputs(12775) <= not (a and b);
    layer2_outputs(12776) <= not b or a;
    layer2_outputs(12777) <= not a or b;
    layer2_outputs(12778) <= not b;
    layer2_outputs(12779) <= not b or a;
    layer2_outputs(12780) <= b;
    layer2_outputs(12781) <= not a or b;
    layer2_outputs(12782) <= a and b;
    layer2_outputs(12783) <= not a or b;
    layer2_outputs(12784) <= '0';
    layer2_outputs(12785) <= a xor b;
    layer2_outputs(12786) <= b;
    layer2_outputs(12787) <= '0';
    layer2_outputs(12788) <= not (a or b);
    layer2_outputs(12789) <= not (a xor b);
    layer2_outputs(12790) <= not (a and b);
    layer2_outputs(12791) <= not a or b;
    layer2_outputs(12792) <= a;
    layer2_outputs(12793) <= b;
    layer2_outputs(12794) <= a and b;
    layer2_outputs(12795) <= '0';
    layer2_outputs(12796) <= b and not a;
    layer2_outputs(12797) <= b;
    layer2_outputs(12798) <= not a or b;
    layer2_outputs(12799) <= a and b;
    layer3_outputs(0) <= not a;
    layer3_outputs(1) <= b and not a;
    layer3_outputs(2) <= a;
    layer3_outputs(3) <= not b or a;
    layer3_outputs(4) <= a and not b;
    layer3_outputs(5) <= not b;
    layer3_outputs(6) <= not a;
    layer3_outputs(7) <= '0';
    layer3_outputs(8) <= b;
    layer3_outputs(9) <= a and b;
    layer3_outputs(10) <= a and not b;
    layer3_outputs(11) <= not a;
    layer3_outputs(12) <= b and not a;
    layer3_outputs(13) <= b and not a;
    layer3_outputs(14) <= a and b;
    layer3_outputs(15) <= not (a and b);
    layer3_outputs(16) <= not (a xor b);
    layer3_outputs(17) <= a and not b;
    layer3_outputs(18) <= a or b;
    layer3_outputs(19) <= a and b;
    layer3_outputs(20) <= not a;
    layer3_outputs(21) <= '0';
    layer3_outputs(22) <= a xor b;
    layer3_outputs(23) <= not b or a;
    layer3_outputs(24) <= not (a and b);
    layer3_outputs(25) <= b;
    layer3_outputs(26) <= not a;
    layer3_outputs(27) <= not (a xor b);
    layer3_outputs(28) <= not a;
    layer3_outputs(29) <= a and b;
    layer3_outputs(30) <= not a;
    layer3_outputs(31) <= b;
    layer3_outputs(32) <= not a;
    layer3_outputs(33) <= '1';
    layer3_outputs(34) <= not b;
    layer3_outputs(35) <= b and not a;
    layer3_outputs(36) <= b;
    layer3_outputs(37) <= not b;
    layer3_outputs(38) <= a and not b;
    layer3_outputs(39) <= a and b;
    layer3_outputs(40) <= not (a and b);
    layer3_outputs(41) <= not b or a;
    layer3_outputs(42) <= a and not b;
    layer3_outputs(43) <= b and not a;
    layer3_outputs(44) <= b;
    layer3_outputs(45) <= not b;
    layer3_outputs(46) <= b;
    layer3_outputs(47) <= b;
    layer3_outputs(48) <= '0';
    layer3_outputs(49) <= a or b;
    layer3_outputs(50) <= '0';
    layer3_outputs(51) <= not a;
    layer3_outputs(52) <= not (a and b);
    layer3_outputs(53) <= not b or a;
    layer3_outputs(54) <= a;
    layer3_outputs(55) <= not b;
    layer3_outputs(56) <= not b;
    layer3_outputs(57) <= a and not b;
    layer3_outputs(58) <= not a;
    layer3_outputs(59) <= a;
    layer3_outputs(60) <= not b;
    layer3_outputs(61) <= b;
    layer3_outputs(62) <= not b;
    layer3_outputs(63) <= b and not a;
    layer3_outputs(64) <= not b or a;
    layer3_outputs(65) <= not (a and b);
    layer3_outputs(66) <= not (a xor b);
    layer3_outputs(67) <= not a or b;
    layer3_outputs(68) <= a;
    layer3_outputs(69) <= not a or b;
    layer3_outputs(70) <= not a or b;
    layer3_outputs(71) <= a;
    layer3_outputs(72) <= a and b;
    layer3_outputs(73) <= b;
    layer3_outputs(74) <= not (a or b);
    layer3_outputs(75) <= a or b;
    layer3_outputs(76) <= '1';
    layer3_outputs(77) <= not a or b;
    layer3_outputs(78) <= not b;
    layer3_outputs(79) <= not (a or b);
    layer3_outputs(80) <= a or b;
    layer3_outputs(81) <= a and not b;
    layer3_outputs(82) <= not a;
    layer3_outputs(83) <= not b;
    layer3_outputs(84) <= a or b;
    layer3_outputs(85) <= b and not a;
    layer3_outputs(86) <= a xor b;
    layer3_outputs(87) <= not b;
    layer3_outputs(88) <= a xor b;
    layer3_outputs(89) <= not (a xor b);
    layer3_outputs(90) <= not (a xor b);
    layer3_outputs(91) <= b;
    layer3_outputs(92) <= not (a or b);
    layer3_outputs(93) <= a or b;
    layer3_outputs(94) <= b;
    layer3_outputs(95) <= b;
    layer3_outputs(96) <= not a;
    layer3_outputs(97) <= a;
    layer3_outputs(98) <= '1';
    layer3_outputs(99) <= not a;
    layer3_outputs(100) <= not a;
    layer3_outputs(101) <= not a;
    layer3_outputs(102) <= '0';
    layer3_outputs(103) <= not b;
    layer3_outputs(104) <= b;
    layer3_outputs(105) <= not (a and b);
    layer3_outputs(106) <= not (a or b);
    layer3_outputs(107) <= a;
    layer3_outputs(108) <= '0';
    layer3_outputs(109) <= not b;
    layer3_outputs(110) <= not (a and b);
    layer3_outputs(111) <= not b;
    layer3_outputs(112) <= a and not b;
    layer3_outputs(113) <= not a or b;
    layer3_outputs(114) <= b and not a;
    layer3_outputs(115) <= b and not a;
    layer3_outputs(116) <= not b;
    layer3_outputs(117) <= not b or a;
    layer3_outputs(118) <= not b;
    layer3_outputs(119) <= not (a or b);
    layer3_outputs(120) <= a xor b;
    layer3_outputs(121) <= not b;
    layer3_outputs(122) <= not b;
    layer3_outputs(123) <= b;
    layer3_outputs(124) <= not (a or b);
    layer3_outputs(125) <= not (a or b);
    layer3_outputs(126) <= not a or b;
    layer3_outputs(127) <= '1';
    layer3_outputs(128) <= not a;
    layer3_outputs(129) <= b;
    layer3_outputs(130) <= a and b;
    layer3_outputs(131) <= a;
    layer3_outputs(132) <= not b;
    layer3_outputs(133) <= not (a xor b);
    layer3_outputs(134) <= not b;
    layer3_outputs(135) <= not a;
    layer3_outputs(136) <= not b;
    layer3_outputs(137) <= not a;
    layer3_outputs(138) <= '1';
    layer3_outputs(139) <= not b;
    layer3_outputs(140) <= a or b;
    layer3_outputs(141) <= not a;
    layer3_outputs(142) <= b;
    layer3_outputs(143) <= a xor b;
    layer3_outputs(144) <= b and not a;
    layer3_outputs(145) <= not (a or b);
    layer3_outputs(146) <= a xor b;
    layer3_outputs(147) <= a and not b;
    layer3_outputs(148) <= not (a xor b);
    layer3_outputs(149) <= not b;
    layer3_outputs(150) <= not b;
    layer3_outputs(151) <= a and not b;
    layer3_outputs(152) <= a and not b;
    layer3_outputs(153) <= not b;
    layer3_outputs(154) <= not a;
    layer3_outputs(155) <= a and b;
    layer3_outputs(156) <= '0';
    layer3_outputs(157) <= not b;
    layer3_outputs(158) <= not a;
    layer3_outputs(159) <= a and b;
    layer3_outputs(160) <= not b;
    layer3_outputs(161) <= not b;
    layer3_outputs(162) <= '1';
    layer3_outputs(163) <= not (a or b);
    layer3_outputs(164) <= a and b;
    layer3_outputs(165) <= a;
    layer3_outputs(166) <= a;
    layer3_outputs(167) <= not (a xor b);
    layer3_outputs(168) <= not (a or b);
    layer3_outputs(169) <= not b;
    layer3_outputs(170) <= '0';
    layer3_outputs(171) <= not (a xor b);
    layer3_outputs(172) <= not b or a;
    layer3_outputs(173) <= not (a or b);
    layer3_outputs(174) <= not b;
    layer3_outputs(175) <= a;
    layer3_outputs(176) <= '1';
    layer3_outputs(177) <= not a;
    layer3_outputs(178) <= not a;
    layer3_outputs(179) <= a;
    layer3_outputs(180) <= not b;
    layer3_outputs(181) <= not (a and b);
    layer3_outputs(182) <= not b or a;
    layer3_outputs(183) <= not b;
    layer3_outputs(184) <= b;
    layer3_outputs(185) <= not a;
    layer3_outputs(186) <= a or b;
    layer3_outputs(187) <= a;
    layer3_outputs(188) <= not b or a;
    layer3_outputs(189) <= not b;
    layer3_outputs(190) <= not b;
    layer3_outputs(191) <= a;
    layer3_outputs(192) <= a and b;
    layer3_outputs(193) <= a xor b;
    layer3_outputs(194) <= b;
    layer3_outputs(195) <= a xor b;
    layer3_outputs(196) <= not (a and b);
    layer3_outputs(197) <= not b or a;
    layer3_outputs(198) <= a and not b;
    layer3_outputs(199) <= not b or a;
    layer3_outputs(200) <= a;
    layer3_outputs(201) <= a and not b;
    layer3_outputs(202) <= a and not b;
    layer3_outputs(203) <= not a;
    layer3_outputs(204) <= not a or b;
    layer3_outputs(205) <= a and b;
    layer3_outputs(206) <= b;
    layer3_outputs(207) <= '0';
    layer3_outputs(208) <= not b;
    layer3_outputs(209) <= '1';
    layer3_outputs(210) <= not b;
    layer3_outputs(211) <= a;
    layer3_outputs(212) <= not (a or b);
    layer3_outputs(213) <= b and not a;
    layer3_outputs(214) <= not b;
    layer3_outputs(215) <= not b;
    layer3_outputs(216) <= b and not a;
    layer3_outputs(217) <= a or b;
    layer3_outputs(218) <= not a or b;
    layer3_outputs(219) <= a;
    layer3_outputs(220) <= '0';
    layer3_outputs(221) <= a;
    layer3_outputs(222) <= not b or a;
    layer3_outputs(223) <= a;
    layer3_outputs(224) <= '0';
    layer3_outputs(225) <= a and b;
    layer3_outputs(226) <= a and not b;
    layer3_outputs(227) <= a and not b;
    layer3_outputs(228) <= b;
    layer3_outputs(229) <= a or b;
    layer3_outputs(230) <= not a;
    layer3_outputs(231) <= b and not a;
    layer3_outputs(232) <= not a or b;
    layer3_outputs(233) <= b;
    layer3_outputs(234) <= not (a and b);
    layer3_outputs(235) <= not b;
    layer3_outputs(236) <= a;
    layer3_outputs(237) <= not b;
    layer3_outputs(238) <= a;
    layer3_outputs(239) <= not (a and b);
    layer3_outputs(240) <= a;
    layer3_outputs(241) <= not b or a;
    layer3_outputs(242) <= not a or b;
    layer3_outputs(243) <= not b or a;
    layer3_outputs(244) <= a and b;
    layer3_outputs(245) <= not a;
    layer3_outputs(246) <= a;
    layer3_outputs(247) <= not a;
    layer3_outputs(248) <= b and not a;
    layer3_outputs(249) <= a and not b;
    layer3_outputs(250) <= a and b;
    layer3_outputs(251) <= a;
    layer3_outputs(252) <= b;
    layer3_outputs(253) <= a and not b;
    layer3_outputs(254) <= b and not a;
    layer3_outputs(255) <= not b;
    layer3_outputs(256) <= not a;
    layer3_outputs(257) <= not (a and b);
    layer3_outputs(258) <= a and b;
    layer3_outputs(259) <= a and not b;
    layer3_outputs(260) <= a;
    layer3_outputs(261) <= a xor b;
    layer3_outputs(262) <= not b;
    layer3_outputs(263) <= a;
    layer3_outputs(264) <= a or b;
    layer3_outputs(265) <= not (a and b);
    layer3_outputs(266) <= '0';
    layer3_outputs(267) <= not (a or b);
    layer3_outputs(268) <= not b;
    layer3_outputs(269) <= a or b;
    layer3_outputs(270) <= a and not b;
    layer3_outputs(271) <= not a;
    layer3_outputs(272) <= b and not a;
    layer3_outputs(273) <= b and not a;
    layer3_outputs(274) <= a;
    layer3_outputs(275) <= not a or b;
    layer3_outputs(276) <= '0';
    layer3_outputs(277) <= a and not b;
    layer3_outputs(278) <= not (a and b);
    layer3_outputs(279) <= not (a or b);
    layer3_outputs(280) <= not b;
    layer3_outputs(281) <= not a or b;
    layer3_outputs(282) <= a;
    layer3_outputs(283) <= not (a or b);
    layer3_outputs(284) <= a xor b;
    layer3_outputs(285) <= not (a or b);
    layer3_outputs(286) <= not (a xor b);
    layer3_outputs(287) <= not (a and b);
    layer3_outputs(288) <= a;
    layer3_outputs(289) <= b;
    layer3_outputs(290) <= a and b;
    layer3_outputs(291) <= '0';
    layer3_outputs(292) <= not (a and b);
    layer3_outputs(293) <= not b;
    layer3_outputs(294) <= b and not a;
    layer3_outputs(295) <= a and not b;
    layer3_outputs(296) <= a and b;
    layer3_outputs(297) <= a or b;
    layer3_outputs(298) <= not (a or b);
    layer3_outputs(299) <= not a;
    layer3_outputs(300) <= b;
    layer3_outputs(301) <= not b or a;
    layer3_outputs(302) <= a;
    layer3_outputs(303) <= not (a and b);
    layer3_outputs(304) <= not a;
    layer3_outputs(305) <= not a or b;
    layer3_outputs(306) <= not (a xor b);
    layer3_outputs(307) <= not a or b;
    layer3_outputs(308) <= not (a and b);
    layer3_outputs(309) <= not b or a;
    layer3_outputs(310) <= a;
    layer3_outputs(311) <= a xor b;
    layer3_outputs(312) <= not a;
    layer3_outputs(313) <= a or b;
    layer3_outputs(314) <= '1';
    layer3_outputs(315) <= '1';
    layer3_outputs(316) <= b;
    layer3_outputs(317) <= b;
    layer3_outputs(318) <= not (a and b);
    layer3_outputs(319) <= a and not b;
    layer3_outputs(320) <= not b or a;
    layer3_outputs(321) <= a;
    layer3_outputs(322) <= a or b;
    layer3_outputs(323) <= b;
    layer3_outputs(324) <= not (a and b);
    layer3_outputs(325) <= not (a xor b);
    layer3_outputs(326) <= a;
    layer3_outputs(327) <= b and not a;
    layer3_outputs(328) <= not a;
    layer3_outputs(329) <= not (a or b);
    layer3_outputs(330) <= a or b;
    layer3_outputs(331) <= a;
    layer3_outputs(332) <= b and not a;
    layer3_outputs(333) <= '0';
    layer3_outputs(334) <= b;
    layer3_outputs(335) <= a;
    layer3_outputs(336) <= b;
    layer3_outputs(337) <= not (a and b);
    layer3_outputs(338) <= not b;
    layer3_outputs(339) <= a;
    layer3_outputs(340) <= not b;
    layer3_outputs(341) <= not (a and b);
    layer3_outputs(342) <= a and not b;
    layer3_outputs(343) <= not (a and b);
    layer3_outputs(344) <= a and not b;
    layer3_outputs(345) <= b and not a;
    layer3_outputs(346) <= not (a or b);
    layer3_outputs(347) <= not b or a;
    layer3_outputs(348) <= not a or b;
    layer3_outputs(349) <= a and b;
    layer3_outputs(350) <= a;
    layer3_outputs(351) <= a or b;
    layer3_outputs(352) <= '1';
    layer3_outputs(353) <= a or b;
    layer3_outputs(354) <= a;
    layer3_outputs(355) <= a and b;
    layer3_outputs(356) <= b and not a;
    layer3_outputs(357) <= b;
    layer3_outputs(358) <= b;
    layer3_outputs(359) <= not (a and b);
    layer3_outputs(360) <= not a;
    layer3_outputs(361) <= a;
    layer3_outputs(362) <= not b;
    layer3_outputs(363) <= not b or a;
    layer3_outputs(364) <= not (a or b);
    layer3_outputs(365) <= not b;
    layer3_outputs(366) <= b;
    layer3_outputs(367) <= a and not b;
    layer3_outputs(368) <= a and b;
    layer3_outputs(369) <= b;
    layer3_outputs(370) <= a and b;
    layer3_outputs(371) <= a and not b;
    layer3_outputs(372) <= not a;
    layer3_outputs(373) <= not b;
    layer3_outputs(374) <= not a;
    layer3_outputs(375) <= '1';
    layer3_outputs(376) <= '0';
    layer3_outputs(377) <= '0';
    layer3_outputs(378) <= b;
    layer3_outputs(379) <= not (a xor b);
    layer3_outputs(380) <= '0';
    layer3_outputs(381) <= a;
    layer3_outputs(382) <= not b or a;
    layer3_outputs(383) <= b and not a;
    layer3_outputs(384) <= b and not a;
    layer3_outputs(385) <= a and not b;
    layer3_outputs(386) <= b;
    layer3_outputs(387) <= not b;
    layer3_outputs(388) <= a or b;
    layer3_outputs(389) <= a or b;
    layer3_outputs(390) <= a or b;
    layer3_outputs(391) <= not (a or b);
    layer3_outputs(392) <= a or b;
    layer3_outputs(393) <= not (a or b);
    layer3_outputs(394) <= '1';
    layer3_outputs(395) <= a;
    layer3_outputs(396) <= not b;
    layer3_outputs(397) <= b;
    layer3_outputs(398) <= not b or a;
    layer3_outputs(399) <= a and b;
    layer3_outputs(400) <= not b or a;
    layer3_outputs(401) <= '0';
    layer3_outputs(402) <= not a or b;
    layer3_outputs(403) <= b;
    layer3_outputs(404) <= a or b;
    layer3_outputs(405) <= a;
    layer3_outputs(406) <= not a;
    layer3_outputs(407) <= a and b;
    layer3_outputs(408) <= not (a and b);
    layer3_outputs(409) <= a and not b;
    layer3_outputs(410) <= b and not a;
    layer3_outputs(411) <= a and not b;
    layer3_outputs(412) <= not b;
    layer3_outputs(413) <= b;
    layer3_outputs(414) <= a and b;
    layer3_outputs(415) <= not a or b;
    layer3_outputs(416) <= b;
    layer3_outputs(417) <= not b;
    layer3_outputs(418) <= a;
    layer3_outputs(419) <= not b;
    layer3_outputs(420) <= a xor b;
    layer3_outputs(421) <= a xor b;
    layer3_outputs(422) <= not a or b;
    layer3_outputs(423) <= a and b;
    layer3_outputs(424) <= not b;
    layer3_outputs(425) <= b and not a;
    layer3_outputs(426) <= b;
    layer3_outputs(427) <= not b or a;
    layer3_outputs(428) <= not a or b;
    layer3_outputs(429) <= not b or a;
    layer3_outputs(430) <= not b or a;
    layer3_outputs(431) <= not (a xor b);
    layer3_outputs(432) <= b;
    layer3_outputs(433) <= b;
    layer3_outputs(434) <= b and not a;
    layer3_outputs(435) <= not (a or b);
    layer3_outputs(436) <= not b or a;
    layer3_outputs(437) <= not (a xor b);
    layer3_outputs(438) <= not b;
    layer3_outputs(439) <= a or b;
    layer3_outputs(440) <= a or b;
    layer3_outputs(441) <= not b;
    layer3_outputs(442) <= not a;
    layer3_outputs(443) <= not a;
    layer3_outputs(444) <= not (a or b);
    layer3_outputs(445) <= not (a or b);
    layer3_outputs(446) <= a or b;
    layer3_outputs(447) <= not b;
    layer3_outputs(448) <= b;
    layer3_outputs(449) <= not (a or b);
    layer3_outputs(450) <= a or b;
    layer3_outputs(451) <= b and not a;
    layer3_outputs(452) <= b;
    layer3_outputs(453) <= a and b;
    layer3_outputs(454) <= not b;
    layer3_outputs(455) <= not (a xor b);
    layer3_outputs(456) <= b and not a;
    layer3_outputs(457) <= a and b;
    layer3_outputs(458) <= '0';
    layer3_outputs(459) <= not b;
    layer3_outputs(460) <= not a;
    layer3_outputs(461) <= not (a or b);
    layer3_outputs(462) <= b;
    layer3_outputs(463) <= not a;
    layer3_outputs(464) <= not b;
    layer3_outputs(465) <= not b or a;
    layer3_outputs(466) <= not b or a;
    layer3_outputs(467) <= b and not a;
    layer3_outputs(468) <= not (a or b);
    layer3_outputs(469) <= b;
    layer3_outputs(470) <= not b;
    layer3_outputs(471) <= not b;
    layer3_outputs(472) <= a or b;
    layer3_outputs(473) <= a and not b;
    layer3_outputs(474) <= a;
    layer3_outputs(475) <= not b;
    layer3_outputs(476) <= not b;
    layer3_outputs(477) <= not b or a;
    layer3_outputs(478) <= a;
    layer3_outputs(479) <= not b;
    layer3_outputs(480) <= not (a or b);
    layer3_outputs(481) <= not b;
    layer3_outputs(482) <= a and b;
    layer3_outputs(483) <= b and not a;
    layer3_outputs(484) <= not (a or b);
    layer3_outputs(485) <= not a or b;
    layer3_outputs(486) <= not (a and b);
    layer3_outputs(487) <= not b;
    layer3_outputs(488) <= a or b;
    layer3_outputs(489) <= b and not a;
    layer3_outputs(490) <= not a or b;
    layer3_outputs(491) <= a and not b;
    layer3_outputs(492) <= not b;
    layer3_outputs(493) <= a and b;
    layer3_outputs(494) <= b;
    layer3_outputs(495) <= b and not a;
    layer3_outputs(496) <= a xor b;
    layer3_outputs(497) <= a or b;
    layer3_outputs(498) <= a and b;
    layer3_outputs(499) <= not b;
    layer3_outputs(500) <= a;
    layer3_outputs(501) <= not b or a;
    layer3_outputs(502) <= not b or a;
    layer3_outputs(503) <= a;
    layer3_outputs(504) <= not b;
    layer3_outputs(505) <= a or b;
    layer3_outputs(506) <= not b;
    layer3_outputs(507) <= not b or a;
    layer3_outputs(508) <= not a;
    layer3_outputs(509) <= not (a and b);
    layer3_outputs(510) <= b;
    layer3_outputs(511) <= a;
    layer3_outputs(512) <= b;
    layer3_outputs(513) <= not a or b;
    layer3_outputs(514) <= not (a or b);
    layer3_outputs(515) <= a and b;
    layer3_outputs(516) <= not b;
    layer3_outputs(517) <= not b or a;
    layer3_outputs(518) <= b;
    layer3_outputs(519) <= a;
    layer3_outputs(520) <= '1';
    layer3_outputs(521) <= a;
    layer3_outputs(522) <= not a;
    layer3_outputs(523) <= not (a xor b);
    layer3_outputs(524) <= a;
    layer3_outputs(525) <= a and b;
    layer3_outputs(526) <= a and not b;
    layer3_outputs(527) <= not (a or b);
    layer3_outputs(528) <= not a;
    layer3_outputs(529) <= a;
    layer3_outputs(530) <= not a;
    layer3_outputs(531) <= a or b;
    layer3_outputs(532) <= a or b;
    layer3_outputs(533) <= a or b;
    layer3_outputs(534) <= not (a or b);
    layer3_outputs(535) <= b;
    layer3_outputs(536) <= b;
    layer3_outputs(537) <= not (a or b);
    layer3_outputs(538) <= not b;
    layer3_outputs(539) <= b;
    layer3_outputs(540) <= a or b;
    layer3_outputs(541) <= a and not b;
    layer3_outputs(542) <= b and not a;
    layer3_outputs(543) <= not a or b;
    layer3_outputs(544) <= not b;
    layer3_outputs(545) <= b;
    layer3_outputs(546) <= a xor b;
    layer3_outputs(547) <= a;
    layer3_outputs(548) <= not (a or b);
    layer3_outputs(549) <= not (a xor b);
    layer3_outputs(550) <= a xor b;
    layer3_outputs(551) <= b and not a;
    layer3_outputs(552) <= not (a xor b);
    layer3_outputs(553) <= not b;
    layer3_outputs(554) <= a xor b;
    layer3_outputs(555) <= not b;
    layer3_outputs(556) <= a xor b;
    layer3_outputs(557) <= not (a and b);
    layer3_outputs(558) <= not b;
    layer3_outputs(559) <= not (a or b);
    layer3_outputs(560) <= not b;
    layer3_outputs(561) <= '1';
    layer3_outputs(562) <= not a;
    layer3_outputs(563) <= not b;
    layer3_outputs(564) <= b;
    layer3_outputs(565) <= a;
    layer3_outputs(566) <= a;
    layer3_outputs(567) <= b;
    layer3_outputs(568) <= not b or a;
    layer3_outputs(569) <= b and not a;
    layer3_outputs(570) <= not b or a;
    layer3_outputs(571) <= '0';
    layer3_outputs(572) <= not (a xor b);
    layer3_outputs(573) <= not a or b;
    layer3_outputs(574) <= a and b;
    layer3_outputs(575) <= a xor b;
    layer3_outputs(576) <= not (a and b);
    layer3_outputs(577) <= not a or b;
    layer3_outputs(578) <= not a or b;
    layer3_outputs(579) <= not (a xor b);
    layer3_outputs(580) <= a and not b;
    layer3_outputs(581) <= a and b;
    layer3_outputs(582) <= not a or b;
    layer3_outputs(583) <= not b;
    layer3_outputs(584) <= not a or b;
    layer3_outputs(585) <= a or b;
    layer3_outputs(586) <= not b;
    layer3_outputs(587) <= not a or b;
    layer3_outputs(588) <= a and not b;
    layer3_outputs(589) <= a;
    layer3_outputs(590) <= not a or b;
    layer3_outputs(591) <= a;
    layer3_outputs(592) <= a and not b;
    layer3_outputs(593) <= b;
    layer3_outputs(594) <= not a;
    layer3_outputs(595) <= b;
    layer3_outputs(596) <= not b or a;
    layer3_outputs(597) <= b and not a;
    layer3_outputs(598) <= not a or b;
    layer3_outputs(599) <= b and not a;
    layer3_outputs(600) <= a or b;
    layer3_outputs(601) <= not a or b;
    layer3_outputs(602) <= a and not b;
    layer3_outputs(603) <= not (a or b);
    layer3_outputs(604) <= not b;
    layer3_outputs(605) <= a or b;
    layer3_outputs(606) <= not (a or b);
    layer3_outputs(607) <= b and not a;
    layer3_outputs(608) <= '1';
    layer3_outputs(609) <= a or b;
    layer3_outputs(610) <= a;
    layer3_outputs(611) <= not (a or b);
    layer3_outputs(612) <= not (a or b);
    layer3_outputs(613) <= not (a or b);
    layer3_outputs(614) <= a;
    layer3_outputs(615) <= b;
    layer3_outputs(616) <= a;
    layer3_outputs(617) <= b;
    layer3_outputs(618) <= a;
    layer3_outputs(619) <= not b;
    layer3_outputs(620) <= b;
    layer3_outputs(621) <= b;
    layer3_outputs(622) <= a or b;
    layer3_outputs(623) <= not a;
    layer3_outputs(624) <= not b or a;
    layer3_outputs(625) <= a;
    layer3_outputs(626) <= not b;
    layer3_outputs(627) <= not a;
    layer3_outputs(628) <= not b or a;
    layer3_outputs(629) <= b and not a;
    layer3_outputs(630) <= '0';
    layer3_outputs(631) <= '0';
    layer3_outputs(632) <= a or b;
    layer3_outputs(633) <= '1';
    layer3_outputs(634) <= a;
    layer3_outputs(635) <= b and not a;
    layer3_outputs(636) <= not b or a;
    layer3_outputs(637) <= not b or a;
    layer3_outputs(638) <= a;
    layer3_outputs(639) <= not b;
    layer3_outputs(640) <= b;
    layer3_outputs(641) <= not b;
    layer3_outputs(642) <= not b or a;
    layer3_outputs(643) <= not b;
    layer3_outputs(644) <= '1';
    layer3_outputs(645) <= not b;
    layer3_outputs(646) <= not a or b;
    layer3_outputs(647) <= a xor b;
    layer3_outputs(648) <= b;
    layer3_outputs(649) <= a and not b;
    layer3_outputs(650) <= a and b;
    layer3_outputs(651) <= b;
    layer3_outputs(652) <= not b;
    layer3_outputs(653) <= not (a xor b);
    layer3_outputs(654) <= not a or b;
    layer3_outputs(655) <= not a;
    layer3_outputs(656) <= not a;
    layer3_outputs(657) <= a;
    layer3_outputs(658) <= not a or b;
    layer3_outputs(659) <= b;
    layer3_outputs(660) <= b;
    layer3_outputs(661) <= not b;
    layer3_outputs(662) <= not a or b;
    layer3_outputs(663) <= '0';
    layer3_outputs(664) <= not a;
    layer3_outputs(665) <= a;
    layer3_outputs(666) <= not b;
    layer3_outputs(667) <= not b;
    layer3_outputs(668) <= b;
    layer3_outputs(669) <= a and b;
    layer3_outputs(670) <= not a or b;
    layer3_outputs(671) <= not (a and b);
    layer3_outputs(672) <= b and not a;
    layer3_outputs(673) <= a and not b;
    layer3_outputs(674) <= '0';
    layer3_outputs(675) <= not b;
    layer3_outputs(676) <= b;
    layer3_outputs(677) <= not a or b;
    layer3_outputs(678) <= a or b;
    layer3_outputs(679) <= '1';
    layer3_outputs(680) <= '0';
    layer3_outputs(681) <= b and not a;
    layer3_outputs(682) <= a and not b;
    layer3_outputs(683) <= a or b;
    layer3_outputs(684) <= a or b;
    layer3_outputs(685) <= not (a and b);
    layer3_outputs(686) <= not a;
    layer3_outputs(687) <= b and not a;
    layer3_outputs(688) <= not a;
    layer3_outputs(689) <= not b;
    layer3_outputs(690) <= b and not a;
    layer3_outputs(691) <= not b;
    layer3_outputs(692) <= a or b;
    layer3_outputs(693) <= b;
    layer3_outputs(694) <= not a;
    layer3_outputs(695) <= not (a xor b);
    layer3_outputs(696) <= not a or b;
    layer3_outputs(697) <= a;
    layer3_outputs(698) <= a;
    layer3_outputs(699) <= not b or a;
    layer3_outputs(700) <= not b;
    layer3_outputs(701) <= not a;
    layer3_outputs(702) <= not (a and b);
    layer3_outputs(703) <= b and not a;
    layer3_outputs(704) <= not b or a;
    layer3_outputs(705) <= a and not b;
    layer3_outputs(706) <= not (a or b);
    layer3_outputs(707) <= not a or b;
    layer3_outputs(708) <= '0';
    layer3_outputs(709) <= b;
    layer3_outputs(710) <= a and not b;
    layer3_outputs(711) <= '1';
    layer3_outputs(712) <= a and b;
    layer3_outputs(713) <= not (a or b);
    layer3_outputs(714) <= a;
    layer3_outputs(715) <= a;
    layer3_outputs(716) <= not a;
    layer3_outputs(717) <= b;
    layer3_outputs(718) <= not b or a;
    layer3_outputs(719) <= not a or b;
    layer3_outputs(720) <= a or b;
    layer3_outputs(721) <= a and b;
    layer3_outputs(722) <= b;
    layer3_outputs(723) <= a;
    layer3_outputs(724) <= b;
    layer3_outputs(725) <= '1';
    layer3_outputs(726) <= a and b;
    layer3_outputs(727) <= b and not a;
    layer3_outputs(728) <= a xor b;
    layer3_outputs(729) <= not b;
    layer3_outputs(730) <= a;
    layer3_outputs(731) <= not b;
    layer3_outputs(732) <= not b;
    layer3_outputs(733) <= a and not b;
    layer3_outputs(734) <= b;
    layer3_outputs(735) <= not a;
    layer3_outputs(736) <= b and not a;
    layer3_outputs(737) <= not a or b;
    layer3_outputs(738) <= a;
    layer3_outputs(739) <= a;
    layer3_outputs(740) <= not b;
    layer3_outputs(741) <= b and not a;
    layer3_outputs(742) <= not b;
    layer3_outputs(743) <= a or b;
    layer3_outputs(744) <= not a;
    layer3_outputs(745) <= not (a and b);
    layer3_outputs(746) <= '0';
    layer3_outputs(747) <= not b or a;
    layer3_outputs(748) <= b;
    layer3_outputs(749) <= b;
    layer3_outputs(750) <= not a;
    layer3_outputs(751) <= a and not b;
    layer3_outputs(752) <= a;
    layer3_outputs(753) <= not (a xor b);
    layer3_outputs(754) <= a;
    layer3_outputs(755) <= a or b;
    layer3_outputs(756) <= '0';
    layer3_outputs(757) <= not b;
    layer3_outputs(758) <= a xor b;
    layer3_outputs(759) <= not a or b;
    layer3_outputs(760) <= not (a and b);
    layer3_outputs(761) <= a xor b;
    layer3_outputs(762) <= not b;
    layer3_outputs(763) <= not a;
    layer3_outputs(764) <= a and b;
    layer3_outputs(765) <= not (a and b);
    layer3_outputs(766) <= a;
    layer3_outputs(767) <= a;
    layer3_outputs(768) <= not b;
    layer3_outputs(769) <= b and not a;
    layer3_outputs(770) <= not (a or b);
    layer3_outputs(771) <= a and b;
    layer3_outputs(772) <= a and not b;
    layer3_outputs(773) <= not a;
    layer3_outputs(774) <= a and not b;
    layer3_outputs(775) <= not a;
    layer3_outputs(776) <= not b or a;
    layer3_outputs(777) <= not a;
    layer3_outputs(778) <= a and b;
    layer3_outputs(779) <= '0';
    layer3_outputs(780) <= not (a or b);
    layer3_outputs(781) <= not b;
    layer3_outputs(782) <= a and not b;
    layer3_outputs(783) <= a and b;
    layer3_outputs(784) <= a or b;
    layer3_outputs(785) <= a and b;
    layer3_outputs(786) <= a;
    layer3_outputs(787) <= not b;
    layer3_outputs(788) <= not (a and b);
    layer3_outputs(789) <= b;
    layer3_outputs(790) <= a xor b;
    layer3_outputs(791) <= not a;
    layer3_outputs(792) <= not (a or b);
    layer3_outputs(793) <= b and not a;
    layer3_outputs(794) <= a xor b;
    layer3_outputs(795) <= not (a and b);
    layer3_outputs(796) <= not b or a;
    layer3_outputs(797) <= '1';
    layer3_outputs(798) <= not b;
    layer3_outputs(799) <= a;
    layer3_outputs(800) <= b;
    layer3_outputs(801) <= not b;
    layer3_outputs(802) <= b and not a;
    layer3_outputs(803) <= a and b;
    layer3_outputs(804) <= a xor b;
    layer3_outputs(805) <= a;
    layer3_outputs(806) <= not b;
    layer3_outputs(807) <= not (a or b);
    layer3_outputs(808) <= '0';
    layer3_outputs(809) <= a xor b;
    layer3_outputs(810) <= a or b;
    layer3_outputs(811) <= not (a xor b);
    layer3_outputs(812) <= not (a and b);
    layer3_outputs(813) <= not (a and b);
    layer3_outputs(814) <= b;
    layer3_outputs(815) <= a and not b;
    layer3_outputs(816) <= not a;
    layer3_outputs(817) <= not a;
    layer3_outputs(818) <= a xor b;
    layer3_outputs(819) <= not a;
    layer3_outputs(820) <= a and b;
    layer3_outputs(821) <= not (a or b);
    layer3_outputs(822) <= not a;
    layer3_outputs(823) <= b and not a;
    layer3_outputs(824) <= a and b;
    layer3_outputs(825) <= a;
    layer3_outputs(826) <= not (a or b);
    layer3_outputs(827) <= not b or a;
    layer3_outputs(828) <= not (a xor b);
    layer3_outputs(829) <= a and not b;
    layer3_outputs(830) <= not a;
    layer3_outputs(831) <= not a or b;
    layer3_outputs(832) <= not (a and b);
    layer3_outputs(833) <= a or b;
    layer3_outputs(834) <= a;
    layer3_outputs(835) <= b;
    layer3_outputs(836) <= '0';
    layer3_outputs(837) <= b and not a;
    layer3_outputs(838) <= not b;
    layer3_outputs(839) <= not b;
    layer3_outputs(840) <= b and not a;
    layer3_outputs(841) <= not a;
    layer3_outputs(842) <= not a or b;
    layer3_outputs(843) <= a and b;
    layer3_outputs(844) <= a;
    layer3_outputs(845) <= a and b;
    layer3_outputs(846) <= b and not a;
    layer3_outputs(847) <= not a or b;
    layer3_outputs(848) <= b and not a;
    layer3_outputs(849) <= not b;
    layer3_outputs(850) <= not a;
    layer3_outputs(851) <= a or b;
    layer3_outputs(852) <= not a;
    layer3_outputs(853) <= b;
    layer3_outputs(854) <= a and not b;
    layer3_outputs(855) <= not (a and b);
    layer3_outputs(856) <= '0';
    layer3_outputs(857) <= not (a and b);
    layer3_outputs(858) <= not a;
    layer3_outputs(859) <= b and not a;
    layer3_outputs(860) <= a;
    layer3_outputs(861) <= not a or b;
    layer3_outputs(862) <= b;
    layer3_outputs(863) <= a and b;
    layer3_outputs(864) <= a xor b;
    layer3_outputs(865) <= b;
    layer3_outputs(866) <= not b or a;
    layer3_outputs(867) <= b;
    layer3_outputs(868) <= '1';
    layer3_outputs(869) <= a xor b;
    layer3_outputs(870) <= not a or b;
    layer3_outputs(871) <= not (a or b);
    layer3_outputs(872) <= a;
    layer3_outputs(873) <= a and b;
    layer3_outputs(874) <= not a or b;
    layer3_outputs(875) <= a xor b;
    layer3_outputs(876) <= b and not a;
    layer3_outputs(877) <= not (a xor b);
    layer3_outputs(878) <= not (a or b);
    layer3_outputs(879) <= a;
    layer3_outputs(880) <= not a;
    layer3_outputs(881) <= not (a xor b);
    layer3_outputs(882) <= not a or b;
    layer3_outputs(883) <= not (a xor b);
    layer3_outputs(884) <= not (a and b);
    layer3_outputs(885) <= not a;
    layer3_outputs(886) <= not b;
    layer3_outputs(887) <= not (a xor b);
    layer3_outputs(888) <= a and b;
    layer3_outputs(889) <= b;
    layer3_outputs(890) <= not (a and b);
    layer3_outputs(891) <= '0';
    layer3_outputs(892) <= not b or a;
    layer3_outputs(893) <= not (a or b);
    layer3_outputs(894) <= not b;
    layer3_outputs(895) <= '1';
    layer3_outputs(896) <= a;
    layer3_outputs(897) <= a and not b;
    layer3_outputs(898) <= not a or b;
    layer3_outputs(899) <= not b;
    layer3_outputs(900) <= not b;
    layer3_outputs(901) <= not a or b;
    layer3_outputs(902) <= not a;
    layer3_outputs(903) <= not a;
    layer3_outputs(904) <= b and not a;
    layer3_outputs(905) <= not b;
    layer3_outputs(906) <= not b or a;
    layer3_outputs(907) <= a or b;
    layer3_outputs(908) <= not b or a;
    layer3_outputs(909) <= not a;
    layer3_outputs(910) <= not b or a;
    layer3_outputs(911) <= b and not a;
    layer3_outputs(912) <= a and b;
    layer3_outputs(913) <= '1';
    layer3_outputs(914) <= not (a xor b);
    layer3_outputs(915) <= not (a xor b);
    layer3_outputs(916) <= a;
    layer3_outputs(917) <= not a;
    layer3_outputs(918) <= not b;
    layer3_outputs(919) <= b and not a;
    layer3_outputs(920) <= not b;
    layer3_outputs(921) <= a xor b;
    layer3_outputs(922) <= not a;
    layer3_outputs(923) <= not a or b;
    layer3_outputs(924) <= a and b;
    layer3_outputs(925) <= '1';
    layer3_outputs(926) <= not (a or b);
    layer3_outputs(927) <= a;
    layer3_outputs(928) <= a or b;
    layer3_outputs(929) <= not a;
    layer3_outputs(930) <= not a or b;
    layer3_outputs(931) <= not a;
    layer3_outputs(932) <= not a or b;
    layer3_outputs(933) <= not (a and b);
    layer3_outputs(934) <= not (a and b);
    layer3_outputs(935) <= a and not b;
    layer3_outputs(936) <= b and not a;
    layer3_outputs(937) <= not (a or b);
    layer3_outputs(938) <= not (a or b);
    layer3_outputs(939) <= not (a and b);
    layer3_outputs(940) <= not a or b;
    layer3_outputs(941) <= not b;
    layer3_outputs(942) <= '0';
    layer3_outputs(943) <= '1';
    layer3_outputs(944) <= not b;
    layer3_outputs(945) <= not a or b;
    layer3_outputs(946) <= a and not b;
    layer3_outputs(947) <= a and not b;
    layer3_outputs(948) <= not b or a;
    layer3_outputs(949) <= a and b;
    layer3_outputs(950) <= not (a or b);
    layer3_outputs(951) <= not a;
    layer3_outputs(952) <= not b;
    layer3_outputs(953) <= a and b;
    layer3_outputs(954) <= not b or a;
    layer3_outputs(955) <= a and b;
    layer3_outputs(956) <= not a;
    layer3_outputs(957) <= a;
    layer3_outputs(958) <= b;
    layer3_outputs(959) <= b;
    layer3_outputs(960) <= not (a and b);
    layer3_outputs(961) <= '1';
    layer3_outputs(962) <= a;
    layer3_outputs(963) <= not (a and b);
    layer3_outputs(964) <= not a;
    layer3_outputs(965) <= a and b;
    layer3_outputs(966) <= b and not a;
    layer3_outputs(967) <= not a;
    layer3_outputs(968) <= not a or b;
    layer3_outputs(969) <= a and not b;
    layer3_outputs(970) <= b;
    layer3_outputs(971) <= not (a and b);
    layer3_outputs(972) <= not (a and b);
    layer3_outputs(973) <= not b;
    layer3_outputs(974) <= not a or b;
    layer3_outputs(975) <= not a or b;
    layer3_outputs(976) <= not b;
    layer3_outputs(977) <= not b;
    layer3_outputs(978) <= a and not b;
    layer3_outputs(979) <= a;
    layer3_outputs(980) <= '0';
    layer3_outputs(981) <= a;
    layer3_outputs(982) <= not b;
    layer3_outputs(983) <= a;
    layer3_outputs(984) <= not a;
    layer3_outputs(985) <= '1';
    layer3_outputs(986) <= not b or a;
    layer3_outputs(987) <= a or b;
    layer3_outputs(988) <= not a;
    layer3_outputs(989) <= not (a or b);
    layer3_outputs(990) <= not a or b;
    layer3_outputs(991) <= not a or b;
    layer3_outputs(992) <= a and b;
    layer3_outputs(993) <= not (a and b);
    layer3_outputs(994) <= b and not a;
    layer3_outputs(995) <= b;
    layer3_outputs(996) <= '0';
    layer3_outputs(997) <= a and b;
    layer3_outputs(998) <= not b;
    layer3_outputs(999) <= a and not b;
    layer3_outputs(1000) <= a xor b;
    layer3_outputs(1001) <= a;
    layer3_outputs(1002) <= not b;
    layer3_outputs(1003) <= '0';
    layer3_outputs(1004) <= a and not b;
    layer3_outputs(1005) <= a and not b;
    layer3_outputs(1006) <= a and b;
    layer3_outputs(1007) <= b and not a;
    layer3_outputs(1008) <= a or b;
    layer3_outputs(1009) <= a and not b;
    layer3_outputs(1010) <= a and not b;
    layer3_outputs(1011) <= not b or a;
    layer3_outputs(1012) <= b;
    layer3_outputs(1013) <= not (a and b);
    layer3_outputs(1014) <= a;
    layer3_outputs(1015) <= a;
    layer3_outputs(1016) <= not a;
    layer3_outputs(1017) <= not (a xor b);
    layer3_outputs(1018) <= not (a and b);
    layer3_outputs(1019) <= a and b;
    layer3_outputs(1020) <= '1';
    layer3_outputs(1021) <= a and b;
    layer3_outputs(1022) <= b;
    layer3_outputs(1023) <= not (a and b);
    layer3_outputs(1024) <= b and not a;
    layer3_outputs(1025) <= not (a xor b);
    layer3_outputs(1026) <= b;
    layer3_outputs(1027) <= b and not a;
    layer3_outputs(1028) <= not (a xor b);
    layer3_outputs(1029) <= not (a or b);
    layer3_outputs(1030) <= not b or a;
    layer3_outputs(1031) <= a and not b;
    layer3_outputs(1032) <= not b;
    layer3_outputs(1033) <= not (a and b);
    layer3_outputs(1034) <= not a;
    layer3_outputs(1035) <= not (a and b);
    layer3_outputs(1036) <= not a;
    layer3_outputs(1037) <= '1';
    layer3_outputs(1038) <= not (a or b);
    layer3_outputs(1039) <= not a;
    layer3_outputs(1040) <= a or b;
    layer3_outputs(1041) <= not a;
    layer3_outputs(1042) <= a xor b;
    layer3_outputs(1043) <= b and not a;
    layer3_outputs(1044) <= b and not a;
    layer3_outputs(1045) <= not (a or b);
    layer3_outputs(1046) <= b and not a;
    layer3_outputs(1047) <= b and not a;
    layer3_outputs(1048) <= a or b;
    layer3_outputs(1049) <= a and b;
    layer3_outputs(1050) <= a or b;
    layer3_outputs(1051) <= b and not a;
    layer3_outputs(1052) <= not b;
    layer3_outputs(1053) <= b and not a;
    layer3_outputs(1054) <= not (a or b);
    layer3_outputs(1055) <= not (a and b);
    layer3_outputs(1056) <= a and b;
    layer3_outputs(1057) <= a;
    layer3_outputs(1058) <= not a;
    layer3_outputs(1059) <= not a;
    layer3_outputs(1060) <= b;
    layer3_outputs(1061) <= not (a and b);
    layer3_outputs(1062) <= a and not b;
    layer3_outputs(1063) <= a and not b;
    layer3_outputs(1064) <= b and not a;
    layer3_outputs(1065) <= b;
    layer3_outputs(1066) <= b and not a;
    layer3_outputs(1067) <= b;
    layer3_outputs(1068) <= not b or a;
    layer3_outputs(1069) <= b and not a;
    layer3_outputs(1070) <= not (a or b);
    layer3_outputs(1071) <= a xor b;
    layer3_outputs(1072) <= a or b;
    layer3_outputs(1073) <= not a or b;
    layer3_outputs(1074) <= '0';
    layer3_outputs(1075) <= b and not a;
    layer3_outputs(1076) <= not b or a;
    layer3_outputs(1077) <= b;
    layer3_outputs(1078) <= a and b;
    layer3_outputs(1079) <= a or b;
    layer3_outputs(1080) <= not a;
    layer3_outputs(1081) <= not (a xor b);
    layer3_outputs(1082) <= not b;
    layer3_outputs(1083) <= not a;
    layer3_outputs(1084) <= not b;
    layer3_outputs(1085) <= not a;
    layer3_outputs(1086) <= not a;
    layer3_outputs(1087) <= a;
    layer3_outputs(1088) <= a and b;
    layer3_outputs(1089) <= not (a xor b);
    layer3_outputs(1090) <= b;
    layer3_outputs(1091) <= a and b;
    layer3_outputs(1092) <= a and not b;
    layer3_outputs(1093) <= b;
    layer3_outputs(1094) <= a xor b;
    layer3_outputs(1095) <= a and not b;
    layer3_outputs(1096) <= b and not a;
    layer3_outputs(1097) <= a and b;
    layer3_outputs(1098) <= not (a xor b);
    layer3_outputs(1099) <= a or b;
    layer3_outputs(1100) <= not (a and b);
    layer3_outputs(1101) <= b;
    layer3_outputs(1102) <= not (a and b);
    layer3_outputs(1103) <= not (a and b);
    layer3_outputs(1104) <= not (a or b);
    layer3_outputs(1105) <= a and b;
    layer3_outputs(1106) <= not (a xor b);
    layer3_outputs(1107) <= not b;
    layer3_outputs(1108) <= not b;
    layer3_outputs(1109) <= b and not a;
    layer3_outputs(1110) <= a;
    layer3_outputs(1111) <= a or b;
    layer3_outputs(1112) <= not a;
    layer3_outputs(1113) <= b;
    layer3_outputs(1114) <= not b;
    layer3_outputs(1115) <= '0';
    layer3_outputs(1116) <= a;
    layer3_outputs(1117) <= not a or b;
    layer3_outputs(1118) <= not (a and b);
    layer3_outputs(1119) <= not b or a;
    layer3_outputs(1120) <= a or b;
    layer3_outputs(1121) <= not (a and b);
    layer3_outputs(1122) <= b;
    layer3_outputs(1123) <= not b;
    layer3_outputs(1124) <= not (a and b);
    layer3_outputs(1125) <= not b;
    layer3_outputs(1126) <= not a or b;
    layer3_outputs(1127) <= not (a or b);
    layer3_outputs(1128) <= '0';
    layer3_outputs(1129) <= not a;
    layer3_outputs(1130) <= a and b;
    layer3_outputs(1131) <= a;
    layer3_outputs(1132) <= not b;
    layer3_outputs(1133) <= b;
    layer3_outputs(1134) <= not a;
    layer3_outputs(1135) <= not b;
    layer3_outputs(1136) <= not (a and b);
    layer3_outputs(1137) <= not a or b;
    layer3_outputs(1138) <= not (a or b);
    layer3_outputs(1139) <= not (a and b);
    layer3_outputs(1140) <= not (a or b);
    layer3_outputs(1141) <= not a;
    layer3_outputs(1142) <= a or b;
    layer3_outputs(1143) <= not a;
    layer3_outputs(1144) <= not b;
    layer3_outputs(1145) <= not (a or b);
    layer3_outputs(1146) <= a and b;
    layer3_outputs(1147) <= b;
    layer3_outputs(1148) <= not a or b;
    layer3_outputs(1149) <= not a;
    layer3_outputs(1150) <= not (a xor b);
    layer3_outputs(1151) <= not a;
    layer3_outputs(1152) <= b and not a;
    layer3_outputs(1153) <= not (a or b);
    layer3_outputs(1154) <= not a or b;
    layer3_outputs(1155) <= not b or a;
    layer3_outputs(1156) <= not b or a;
    layer3_outputs(1157) <= not (a and b);
    layer3_outputs(1158) <= a;
    layer3_outputs(1159) <= not (a or b);
    layer3_outputs(1160) <= not (a xor b);
    layer3_outputs(1161) <= a and b;
    layer3_outputs(1162) <= not (a xor b);
    layer3_outputs(1163) <= not b;
    layer3_outputs(1164) <= not a or b;
    layer3_outputs(1165) <= a;
    layer3_outputs(1166) <= b;
    layer3_outputs(1167) <= not (a xor b);
    layer3_outputs(1168) <= '0';
    layer3_outputs(1169) <= not (a or b);
    layer3_outputs(1170) <= b;
    layer3_outputs(1171) <= not a or b;
    layer3_outputs(1172) <= not b;
    layer3_outputs(1173) <= not (a and b);
    layer3_outputs(1174) <= not b;
    layer3_outputs(1175) <= '0';
    layer3_outputs(1176) <= a;
    layer3_outputs(1177) <= b;
    layer3_outputs(1178) <= a;
    layer3_outputs(1179) <= b;
    layer3_outputs(1180) <= not (a and b);
    layer3_outputs(1181) <= not b;
    layer3_outputs(1182) <= not (a or b);
    layer3_outputs(1183) <= b;
    layer3_outputs(1184) <= not b;
    layer3_outputs(1185) <= '1';
    layer3_outputs(1186) <= not (a or b);
    layer3_outputs(1187) <= '1';
    layer3_outputs(1188) <= not a;
    layer3_outputs(1189) <= not (a and b);
    layer3_outputs(1190) <= a;
    layer3_outputs(1191) <= not b or a;
    layer3_outputs(1192) <= b;
    layer3_outputs(1193) <= b and not a;
    layer3_outputs(1194) <= not a;
    layer3_outputs(1195) <= a;
    layer3_outputs(1196) <= not (a xor b);
    layer3_outputs(1197) <= a;
    layer3_outputs(1198) <= b;
    layer3_outputs(1199) <= a or b;
    layer3_outputs(1200) <= not b;
    layer3_outputs(1201) <= a;
    layer3_outputs(1202) <= not (a and b);
    layer3_outputs(1203) <= not (a or b);
    layer3_outputs(1204) <= not a or b;
    layer3_outputs(1205) <= not (a xor b);
    layer3_outputs(1206) <= a and not b;
    layer3_outputs(1207) <= not b;
    layer3_outputs(1208) <= a and b;
    layer3_outputs(1209) <= not b;
    layer3_outputs(1210) <= not (a or b);
    layer3_outputs(1211) <= not (a or b);
    layer3_outputs(1212) <= not b;
    layer3_outputs(1213) <= not b;
    layer3_outputs(1214) <= '1';
    layer3_outputs(1215) <= b and not a;
    layer3_outputs(1216) <= not b;
    layer3_outputs(1217) <= '1';
    layer3_outputs(1218) <= a and b;
    layer3_outputs(1219) <= a xor b;
    layer3_outputs(1220) <= a;
    layer3_outputs(1221) <= a and not b;
    layer3_outputs(1222) <= not a;
    layer3_outputs(1223) <= a and not b;
    layer3_outputs(1224) <= a and not b;
    layer3_outputs(1225) <= not a;
    layer3_outputs(1226) <= not b;
    layer3_outputs(1227) <= a and not b;
    layer3_outputs(1228) <= a and b;
    layer3_outputs(1229) <= not b;
    layer3_outputs(1230) <= not b;
    layer3_outputs(1231) <= not (a or b);
    layer3_outputs(1232) <= b and not a;
    layer3_outputs(1233) <= b and not a;
    layer3_outputs(1234) <= b and not a;
    layer3_outputs(1235) <= not a;
    layer3_outputs(1236) <= a and b;
    layer3_outputs(1237) <= not a;
    layer3_outputs(1238) <= '0';
    layer3_outputs(1239) <= not (a and b);
    layer3_outputs(1240) <= not a or b;
    layer3_outputs(1241) <= a and b;
    layer3_outputs(1242) <= b;
    layer3_outputs(1243) <= not (a and b);
    layer3_outputs(1244) <= not (a or b);
    layer3_outputs(1245) <= a or b;
    layer3_outputs(1246) <= '0';
    layer3_outputs(1247) <= a;
    layer3_outputs(1248) <= a and b;
    layer3_outputs(1249) <= not (a or b);
    layer3_outputs(1250) <= not a or b;
    layer3_outputs(1251) <= a and b;
    layer3_outputs(1252) <= a or b;
    layer3_outputs(1253) <= not a or b;
    layer3_outputs(1254) <= not (a xor b);
    layer3_outputs(1255) <= not (a and b);
    layer3_outputs(1256) <= not a or b;
    layer3_outputs(1257) <= not (a or b);
    layer3_outputs(1258) <= a xor b;
    layer3_outputs(1259) <= not a;
    layer3_outputs(1260) <= not (a xor b);
    layer3_outputs(1261) <= a or b;
    layer3_outputs(1262) <= '1';
    layer3_outputs(1263) <= not b;
    layer3_outputs(1264) <= not b;
    layer3_outputs(1265) <= '0';
    layer3_outputs(1266) <= a or b;
    layer3_outputs(1267) <= not (a and b);
    layer3_outputs(1268) <= b;
    layer3_outputs(1269) <= a and not b;
    layer3_outputs(1270) <= a xor b;
    layer3_outputs(1271) <= b;
    layer3_outputs(1272) <= not b;
    layer3_outputs(1273) <= not a;
    layer3_outputs(1274) <= a and not b;
    layer3_outputs(1275) <= '1';
    layer3_outputs(1276) <= a and b;
    layer3_outputs(1277) <= a and not b;
    layer3_outputs(1278) <= not (a or b);
    layer3_outputs(1279) <= a and not b;
    layer3_outputs(1280) <= not b;
    layer3_outputs(1281) <= not a;
    layer3_outputs(1282) <= a and b;
    layer3_outputs(1283) <= not (a xor b);
    layer3_outputs(1284) <= not a;
    layer3_outputs(1285) <= not (a and b);
    layer3_outputs(1286) <= a;
    layer3_outputs(1287) <= not b or a;
    layer3_outputs(1288) <= not b;
    layer3_outputs(1289) <= not b;
    layer3_outputs(1290) <= a and not b;
    layer3_outputs(1291) <= not a;
    layer3_outputs(1292) <= not b;
    layer3_outputs(1293) <= not (a and b);
    layer3_outputs(1294) <= a;
    layer3_outputs(1295) <= not (a or b);
    layer3_outputs(1296) <= a;
    layer3_outputs(1297) <= b;
    layer3_outputs(1298) <= not a;
    layer3_outputs(1299) <= not b or a;
    layer3_outputs(1300) <= a or b;
    layer3_outputs(1301) <= '1';
    layer3_outputs(1302) <= a or b;
    layer3_outputs(1303) <= '0';
    layer3_outputs(1304) <= not (a xor b);
    layer3_outputs(1305) <= not (a or b);
    layer3_outputs(1306) <= b;
    layer3_outputs(1307) <= a or b;
    layer3_outputs(1308) <= not (a xor b);
    layer3_outputs(1309) <= '1';
    layer3_outputs(1310) <= not a or b;
    layer3_outputs(1311) <= not (a or b);
    layer3_outputs(1312) <= a xor b;
    layer3_outputs(1313) <= '1';
    layer3_outputs(1314) <= a and not b;
    layer3_outputs(1315) <= a;
    layer3_outputs(1316) <= not a;
    layer3_outputs(1317) <= a xor b;
    layer3_outputs(1318) <= a or b;
    layer3_outputs(1319) <= not b;
    layer3_outputs(1320) <= not b;
    layer3_outputs(1321) <= b;
    layer3_outputs(1322) <= not (a and b);
    layer3_outputs(1323) <= not b;
    layer3_outputs(1324) <= a xor b;
    layer3_outputs(1325) <= not a;
    layer3_outputs(1326) <= not (a or b);
    layer3_outputs(1327) <= not b or a;
    layer3_outputs(1328) <= '1';
    layer3_outputs(1329) <= b;
    layer3_outputs(1330) <= not a;
    layer3_outputs(1331) <= a;
    layer3_outputs(1332) <= a and b;
    layer3_outputs(1333) <= not a;
    layer3_outputs(1334) <= a or b;
    layer3_outputs(1335) <= a and not b;
    layer3_outputs(1336) <= not a;
    layer3_outputs(1337) <= b and not a;
    layer3_outputs(1338) <= not a or b;
    layer3_outputs(1339) <= '1';
    layer3_outputs(1340) <= a;
    layer3_outputs(1341) <= a and not b;
    layer3_outputs(1342) <= a xor b;
    layer3_outputs(1343) <= not (a xor b);
    layer3_outputs(1344) <= not b or a;
    layer3_outputs(1345) <= b and not a;
    layer3_outputs(1346) <= b;
    layer3_outputs(1347) <= not b;
    layer3_outputs(1348) <= b;
    layer3_outputs(1349) <= '1';
    layer3_outputs(1350) <= a;
    layer3_outputs(1351) <= not (a and b);
    layer3_outputs(1352) <= not (a and b);
    layer3_outputs(1353) <= b;
    layer3_outputs(1354) <= not b or a;
    layer3_outputs(1355) <= not b;
    layer3_outputs(1356) <= '1';
    layer3_outputs(1357) <= b and not a;
    layer3_outputs(1358) <= b;
    layer3_outputs(1359) <= b;
    layer3_outputs(1360) <= a xor b;
    layer3_outputs(1361) <= not b or a;
    layer3_outputs(1362) <= not b;
    layer3_outputs(1363) <= not (a or b);
    layer3_outputs(1364) <= '1';
    layer3_outputs(1365) <= not a or b;
    layer3_outputs(1366) <= not a or b;
    layer3_outputs(1367) <= '1';
    layer3_outputs(1368) <= not a;
    layer3_outputs(1369) <= b;
    layer3_outputs(1370) <= not (a and b);
    layer3_outputs(1371) <= a;
    layer3_outputs(1372) <= not (a xor b);
    layer3_outputs(1373) <= a and b;
    layer3_outputs(1374) <= not (a and b);
    layer3_outputs(1375) <= not b;
    layer3_outputs(1376) <= a or b;
    layer3_outputs(1377) <= a;
    layer3_outputs(1378) <= '0';
    layer3_outputs(1379) <= b;
    layer3_outputs(1380) <= not a;
    layer3_outputs(1381) <= not a;
    layer3_outputs(1382) <= not b;
    layer3_outputs(1383) <= not a;
    layer3_outputs(1384) <= a or b;
    layer3_outputs(1385) <= a;
    layer3_outputs(1386) <= b;
    layer3_outputs(1387) <= not b;
    layer3_outputs(1388) <= not a;
    layer3_outputs(1389) <= b and not a;
    layer3_outputs(1390) <= b;
    layer3_outputs(1391) <= a xor b;
    layer3_outputs(1392) <= not b or a;
    layer3_outputs(1393) <= a and not b;
    layer3_outputs(1394) <= b and not a;
    layer3_outputs(1395) <= a and b;
    layer3_outputs(1396) <= not a or b;
    layer3_outputs(1397) <= not b or a;
    layer3_outputs(1398) <= not (a and b);
    layer3_outputs(1399) <= b and not a;
    layer3_outputs(1400) <= not b;
    layer3_outputs(1401) <= a;
    layer3_outputs(1402) <= '1';
    layer3_outputs(1403) <= not b or a;
    layer3_outputs(1404) <= a and b;
    layer3_outputs(1405) <= a;
    layer3_outputs(1406) <= not b;
    layer3_outputs(1407) <= a;
    layer3_outputs(1408) <= a and not b;
    layer3_outputs(1409) <= b;
    layer3_outputs(1410) <= not b or a;
    layer3_outputs(1411) <= b;
    layer3_outputs(1412) <= not (a and b);
    layer3_outputs(1413) <= a xor b;
    layer3_outputs(1414) <= not a or b;
    layer3_outputs(1415) <= a or b;
    layer3_outputs(1416) <= a or b;
    layer3_outputs(1417) <= a;
    layer3_outputs(1418) <= '0';
    layer3_outputs(1419) <= b;
    layer3_outputs(1420) <= b;
    layer3_outputs(1421) <= not b;
    layer3_outputs(1422) <= not a;
    layer3_outputs(1423) <= not (a and b);
    layer3_outputs(1424) <= not b;
    layer3_outputs(1425) <= a;
    layer3_outputs(1426) <= a and not b;
    layer3_outputs(1427) <= b and not a;
    layer3_outputs(1428) <= not (a xor b);
    layer3_outputs(1429) <= '0';
    layer3_outputs(1430) <= a;
    layer3_outputs(1431) <= not (a and b);
    layer3_outputs(1432) <= '0';
    layer3_outputs(1433) <= b;
    layer3_outputs(1434) <= not (a and b);
    layer3_outputs(1435) <= a or b;
    layer3_outputs(1436) <= not (a and b);
    layer3_outputs(1437) <= not b or a;
    layer3_outputs(1438) <= '1';
    layer3_outputs(1439) <= a;
    layer3_outputs(1440) <= b;
    layer3_outputs(1441) <= not (a or b);
    layer3_outputs(1442) <= a;
    layer3_outputs(1443) <= not b;
    layer3_outputs(1444) <= b and not a;
    layer3_outputs(1445) <= not (a xor b);
    layer3_outputs(1446) <= not b;
    layer3_outputs(1447) <= a and not b;
    layer3_outputs(1448) <= b;
    layer3_outputs(1449) <= a and b;
    layer3_outputs(1450) <= not a;
    layer3_outputs(1451) <= a and not b;
    layer3_outputs(1452) <= a or b;
    layer3_outputs(1453) <= a;
    layer3_outputs(1454) <= not b;
    layer3_outputs(1455) <= a and not b;
    layer3_outputs(1456) <= b and not a;
    layer3_outputs(1457) <= not a;
    layer3_outputs(1458) <= a or b;
    layer3_outputs(1459) <= b;
    layer3_outputs(1460) <= not b;
    layer3_outputs(1461) <= b;
    layer3_outputs(1462) <= b and not a;
    layer3_outputs(1463) <= b and not a;
    layer3_outputs(1464) <= a or b;
    layer3_outputs(1465) <= b;
    layer3_outputs(1466) <= not b;
    layer3_outputs(1467) <= not a;
    layer3_outputs(1468) <= not a or b;
    layer3_outputs(1469) <= not b;
    layer3_outputs(1470) <= a xor b;
    layer3_outputs(1471) <= '0';
    layer3_outputs(1472) <= not b or a;
    layer3_outputs(1473) <= not a;
    layer3_outputs(1474) <= not (a or b);
    layer3_outputs(1475) <= '1';
    layer3_outputs(1476) <= a and not b;
    layer3_outputs(1477) <= a and b;
    layer3_outputs(1478) <= a and b;
    layer3_outputs(1479) <= a and not b;
    layer3_outputs(1480) <= a and not b;
    layer3_outputs(1481) <= b;
    layer3_outputs(1482) <= not b;
    layer3_outputs(1483) <= not (a and b);
    layer3_outputs(1484) <= a;
    layer3_outputs(1485) <= a or b;
    layer3_outputs(1486) <= a xor b;
    layer3_outputs(1487) <= not b or a;
    layer3_outputs(1488) <= not b;
    layer3_outputs(1489) <= a;
    layer3_outputs(1490) <= not (a xor b);
    layer3_outputs(1491) <= not b or a;
    layer3_outputs(1492) <= not b or a;
    layer3_outputs(1493) <= not a or b;
    layer3_outputs(1494) <= b and not a;
    layer3_outputs(1495) <= '0';
    layer3_outputs(1496) <= not a;
    layer3_outputs(1497) <= not b;
    layer3_outputs(1498) <= a xor b;
    layer3_outputs(1499) <= not b;
    layer3_outputs(1500) <= not a or b;
    layer3_outputs(1501) <= not (a or b);
    layer3_outputs(1502) <= b and not a;
    layer3_outputs(1503) <= a and not b;
    layer3_outputs(1504) <= a and not b;
    layer3_outputs(1505) <= not b;
    layer3_outputs(1506) <= a;
    layer3_outputs(1507) <= b;
    layer3_outputs(1508) <= not (a xor b);
    layer3_outputs(1509) <= b;
    layer3_outputs(1510) <= a;
    layer3_outputs(1511) <= not b;
    layer3_outputs(1512) <= a and not b;
    layer3_outputs(1513) <= a and b;
    layer3_outputs(1514) <= not (a or b);
    layer3_outputs(1515) <= a or b;
    layer3_outputs(1516) <= not b;
    layer3_outputs(1517) <= not a;
    layer3_outputs(1518) <= '0';
    layer3_outputs(1519) <= b;
    layer3_outputs(1520) <= a and not b;
    layer3_outputs(1521) <= '0';
    layer3_outputs(1522) <= not a;
    layer3_outputs(1523) <= a;
    layer3_outputs(1524) <= a and not b;
    layer3_outputs(1525) <= not (a and b);
    layer3_outputs(1526) <= '1';
    layer3_outputs(1527) <= not (a or b);
    layer3_outputs(1528) <= not a;
    layer3_outputs(1529) <= '1';
    layer3_outputs(1530) <= not a;
    layer3_outputs(1531) <= b;
    layer3_outputs(1532) <= a or b;
    layer3_outputs(1533) <= not b or a;
    layer3_outputs(1534) <= not (a or b);
    layer3_outputs(1535) <= a and not b;
    layer3_outputs(1536) <= a;
    layer3_outputs(1537) <= a;
    layer3_outputs(1538) <= not b;
    layer3_outputs(1539) <= not (a or b);
    layer3_outputs(1540) <= a xor b;
    layer3_outputs(1541) <= a xor b;
    layer3_outputs(1542) <= a and b;
    layer3_outputs(1543) <= not a;
    layer3_outputs(1544) <= '1';
    layer3_outputs(1545) <= a;
    layer3_outputs(1546) <= a or b;
    layer3_outputs(1547) <= b;
    layer3_outputs(1548) <= not a;
    layer3_outputs(1549) <= not b or a;
    layer3_outputs(1550) <= a;
    layer3_outputs(1551) <= not a;
    layer3_outputs(1552) <= not a or b;
    layer3_outputs(1553) <= not (a or b);
    layer3_outputs(1554) <= not (a and b);
    layer3_outputs(1555) <= a and b;
    layer3_outputs(1556) <= not b;
    layer3_outputs(1557) <= a and b;
    layer3_outputs(1558) <= a;
    layer3_outputs(1559) <= not b;
    layer3_outputs(1560) <= not a;
    layer3_outputs(1561) <= not b;
    layer3_outputs(1562) <= b and not a;
    layer3_outputs(1563) <= a and not b;
    layer3_outputs(1564) <= not a or b;
    layer3_outputs(1565) <= not a;
    layer3_outputs(1566) <= not a or b;
    layer3_outputs(1567) <= a or b;
    layer3_outputs(1568) <= a and not b;
    layer3_outputs(1569) <= not a or b;
    layer3_outputs(1570) <= '1';
    layer3_outputs(1571) <= a and b;
    layer3_outputs(1572) <= '1';
    layer3_outputs(1573) <= not (a and b);
    layer3_outputs(1574) <= not (a or b);
    layer3_outputs(1575) <= not a or b;
    layer3_outputs(1576) <= not a;
    layer3_outputs(1577) <= a;
    layer3_outputs(1578) <= not (a and b);
    layer3_outputs(1579) <= a or b;
    layer3_outputs(1580) <= b and not a;
    layer3_outputs(1581) <= a or b;
    layer3_outputs(1582) <= not (a xor b);
    layer3_outputs(1583) <= a and b;
    layer3_outputs(1584) <= not (a xor b);
    layer3_outputs(1585) <= a and not b;
    layer3_outputs(1586) <= a or b;
    layer3_outputs(1587) <= not (a xor b);
    layer3_outputs(1588) <= not a;
    layer3_outputs(1589) <= a or b;
    layer3_outputs(1590) <= not a;
    layer3_outputs(1591) <= a;
    layer3_outputs(1592) <= b;
    layer3_outputs(1593) <= a;
    layer3_outputs(1594) <= not a;
    layer3_outputs(1595) <= a;
    layer3_outputs(1596) <= '0';
    layer3_outputs(1597) <= not a;
    layer3_outputs(1598) <= a;
    layer3_outputs(1599) <= not (a xor b);
    layer3_outputs(1600) <= a;
    layer3_outputs(1601) <= not a;
    layer3_outputs(1602) <= not b;
    layer3_outputs(1603) <= not b;
    layer3_outputs(1604) <= not (a and b);
    layer3_outputs(1605) <= b;
    layer3_outputs(1606) <= '0';
    layer3_outputs(1607) <= not (a and b);
    layer3_outputs(1608) <= not (a xor b);
    layer3_outputs(1609) <= not b or a;
    layer3_outputs(1610) <= '0';
    layer3_outputs(1611) <= a or b;
    layer3_outputs(1612) <= b;
    layer3_outputs(1613) <= not b;
    layer3_outputs(1614) <= a xor b;
    layer3_outputs(1615) <= not b;
    layer3_outputs(1616) <= not (a and b);
    layer3_outputs(1617) <= not a or b;
    layer3_outputs(1618) <= not (a xor b);
    layer3_outputs(1619) <= not (a xor b);
    layer3_outputs(1620) <= not a or b;
    layer3_outputs(1621) <= a xor b;
    layer3_outputs(1622) <= not (a and b);
    layer3_outputs(1623) <= a and b;
    layer3_outputs(1624) <= not a or b;
    layer3_outputs(1625) <= b;
    layer3_outputs(1626) <= '1';
    layer3_outputs(1627) <= a or b;
    layer3_outputs(1628) <= a;
    layer3_outputs(1629) <= not a or b;
    layer3_outputs(1630) <= not b;
    layer3_outputs(1631) <= not a;
    layer3_outputs(1632) <= a or b;
    layer3_outputs(1633) <= a and not b;
    layer3_outputs(1634) <= b;
    layer3_outputs(1635) <= not b;
    layer3_outputs(1636) <= a or b;
    layer3_outputs(1637) <= '0';
    layer3_outputs(1638) <= not (a and b);
    layer3_outputs(1639) <= not a;
    layer3_outputs(1640) <= a;
    layer3_outputs(1641) <= not (a and b);
    layer3_outputs(1642) <= not (a or b);
    layer3_outputs(1643) <= a;
    layer3_outputs(1644) <= a and b;
    layer3_outputs(1645) <= not (a or b);
    layer3_outputs(1646) <= not (a xor b);
    layer3_outputs(1647) <= a or b;
    layer3_outputs(1648) <= not (a and b);
    layer3_outputs(1649) <= a and b;
    layer3_outputs(1650) <= not b or a;
    layer3_outputs(1651) <= not b;
    layer3_outputs(1652) <= b and not a;
    layer3_outputs(1653) <= a and b;
    layer3_outputs(1654) <= not b or a;
    layer3_outputs(1655) <= b and not a;
    layer3_outputs(1656) <= not (a xor b);
    layer3_outputs(1657) <= a xor b;
    layer3_outputs(1658) <= not (a or b);
    layer3_outputs(1659) <= a and not b;
    layer3_outputs(1660) <= a;
    layer3_outputs(1661) <= b;
    layer3_outputs(1662) <= a;
    layer3_outputs(1663) <= a;
    layer3_outputs(1664) <= not b;
    layer3_outputs(1665) <= a and b;
    layer3_outputs(1666) <= not b;
    layer3_outputs(1667) <= a or b;
    layer3_outputs(1668) <= b;
    layer3_outputs(1669) <= not b;
    layer3_outputs(1670) <= not (a or b);
    layer3_outputs(1671) <= not (a and b);
    layer3_outputs(1672) <= a;
    layer3_outputs(1673) <= a and not b;
    layer3_outputs(1674) <= not a;
    layer3_outputs(1675) <= a and not b;
    layer3_outputs(1676) <= not b or a;
    layer3_outputs(1677) <= a and b;
    layer3_outputs(1678) <= b;
    layer3_outputs(1679) <= a or b;
    layer3_outputs(1680) <= a;
    layer3_outputs(1681) <= a;
    layer3_outputs(1682) <= b;
    layer3_outputs(1683) <= not b;
    layer3_outputs(1684) <= b and not a;
    layer3_outputs(1685) <= a and b;
    layer3_outputs(1686) <= a xor b;
    layer3_outputs(1687) <= not (a and b);
    layer3_outputs(1688) <= '0';
    layer3_outputs(1689) <= a and not b;
    layer3_outputs(1690) <= not (a or b);
    layer3_outputs(1691) <= '1';
    layer3_outputs(1692) <= a xor b;
    layer3_outputs(1693) <= b;
    layer3_outputs(1694) <= not (a and b);
    layer3_outputs(1695) <= not (a and b);
    layer3_outputs(1696) <= a and b;
    layer3_outputs(1697) <= a or b;
    layer3_outputs(1698) <= a;
    layer3_outputs(1699) <= not b or a;
    layer3_outputs(1700) <= b;
    layer3_outputs(1701) <= not (a or b);
    layer3_outputs(1702) <= b and not a;
    layer3_outputs(1703) <= not a or b;
    layer3_outputs(1704) <= not b;
    layer3_outputs(1705) <= a;
    layer3_outputs(1706) <= '1';
    layer3_outputs(1707) <= not b or a;
    layer3_outputs(1708) <= not a or b;
    layer3_outputs(1709) <= '1';
    layer3_outputs(1710) <= a and not b;
    layer3_outputs(1711) <= a and b;
    layer3_outputs(1712) <= not (a xor b);
    layer3_outputs(1713) <= a xor b;
    layer3_outputs(1714) <= not a or b;
    layer3_outputs(1715) <= a and not b;
    layer3_outputs(1716) <= not b;
    layer3_outputs(1717) <= a xor b;
    layer3_outputs(1718) <= b;
    layer3_outputs(1719) <= not b;
    layer3_outputs(1720) <= not (a and b);
    layer3_outputs(1721) <= a or b;
    layer3_outputs(1722) <= a and not b;
    layer3_outputs(1723) <= not b;
    layer3_outputs(1724) <= b and not a;
    layer3_outputs(1725) <= '1';
    layer3_outputs(1726) <= not a or b;
    layer3_outputs(1727) <= a and not b;
    layer3_outputs(1728) <= not b;
    layer3_outputs(1729) <= b and not a;
    layer3_outputs(1730) <= a and b;
    layer3_outputs(1731) <= a and not b;
    layer3_outputs(1732) <= a and not b;
    layer3_outputs(1733) <= '1';
    layer3_outputs(1734) <= b;
    layer3_outputs(1735) <= a;
    layer3_outputs(1736) <= b;
    layer3_outputs(1737) <= b and not a;
    layer3_outputs(1738) <= not b;
    layer3_outputs(1739) <= not a;
    layer3_outputs(1740) <= a and b;
    layer3_outputs(1741) <= b;
    layer3_outputs(1742) <= '1';
    layer3_outputs(1743) <= not b;
    layer3_outputs(1744) <= not b or a;
    layer3_outputs(1745) <= not (a and b);
    layer3_outputs(1746) <= not b;
    layer3_outputs(1747) <= not (a or b);
    layer3_outputs(1748) <= a or b;
    layer3_outputs(1749) <= not b;
    layer3_outputs(1750) <= a xor b;
    layer3_outputs(1751) <= not b;
    layer3_outputs(1752) <= b and not a;
    layer3_outputs(1753) <= b and not a;
    layer3_outputs(1754) <= not b;
    layer3_outputs(1755) <= not b;
    layer3_outputs(1756) <= not a;
    layer3_outputs(1757) <= not b;
    layer3_outputs(1758) <= not a;
    layer3_outputs(1759) <= not a;
    layer3_outputs(1760) <= '1';
    layer3_outputs(1761) <= a;
    layer3_outputs(1762) <= not b or a;
    layer3_outputs(1763) <= a or b;
    layer3_outputs(1764) <= not a;
    layer3_outputs(1765) <= a xor b;
    layer3_outputs(1766) <= a and b;
    layer3_outputs(1767) <= not a;
    layer3_outputs(1768) <= a and not b;
    layer3_outputs(1769) <= not b;
    layer3_outputs(1770) <= a and not b;
    layer3_outputs(1771) <= b;
    layer3_outputs(1772) <= not b or a;
    layer3_outputs(1773) <= b;
    layer3_outputs(1774) <= a and b;
    layer3_outputs(1775) <= a;
    layer3_outputs(1776) <= not (a and b);
    layer3_outputs(1777) <= not b;
    layer3_outputs(1778) <= a xor b;
    layer3_outputs(1779) <= a;
    layer3_outputs(1780) <= not b;
    layer3_outputs(1781) <= not (a or b);
    layer3_outputs(1782) <= a and not b;
    layer3_outputs(1783) <= a;
    layer3_outputs(1784) <= not (a or b);
    layer3_outputs(1785) <= not a;
    layer3_outputs(1786) <= not (a or b);
    layer3_outputs(1787) <= not a;
    layer3_outputs(1788) <= b and not a;
    layer3_outputs(1789) <= not b or a;
    layer3_outputs(1790) <= a and not b;
    layer3_outputs(1791) <= a and b;
    layer3_outputs(1792) <= not a;
    layer3_outputs(1793) <= not b or a;
    layer3_outputs(1794) <= '1';
    layer3_outputs(1795) <= '0';
    layer3_outputs(1796) <= not b;
    layer3_outputs(1797) <= not a or b;
    layer3_outputs(1798) <= not b;
    layer3_outputs(1799) <= b;
    layer3_outputs(1800) <= not a;
    layer3_outputs(1801) <= a xor b;
    layer3_outputs(1802) <= a and b;
    layer3_outputs(1803) <= not (a and b);
    layer3_outputs(1804) <= b;
    layer3_outputs(1805) <= b;
    layer3_outputs(1806) <= not b;
    layer3_outputs(1807) <= not b or a;
    layer3_outputs(1808) <= b and not a;
    layer3_outputs(1809) <= a or b;
    layer3_outputs(1810) <= not a or b;
    layer3_outputs(1811) <= '1';
    layer3_outputs(1812) <= not b or a;
    layer3_outputs(1813) <= a and not b;
    layer3_outputs(1814) <= not a or b;
    layer3_outputs(1815) <= a or b;
    layer3_outputs(1816) <= a;
    layer3_outputs(1817) <= a;
    layer3_outputs(1818) <= b;
    layer3_outputs(1819) <= not a;
    layer3_outputs(1820) <= not (a and b);
    layer3_outputs(1821) <= not a;
    layer3_outputs(1822) <= not a or b;
    layer3_outputs(1823) <= a;
    layer3_outputs(1824) <= not b;
    layer3_outputs(1825) <= not (a xor b);
    layer3_outputs(1826) <= a or b;
    layer3_outputs(1827) <= not a or b;
    layer3_outputs(1828) <= not (a or b);
    layer3_outputs(1829) <= not b;
    layer3_outputs(1830) <= not b;
    layer3_outputs(1831) <= not b;
    layer3_outputs(1832) <= not b;
    layer3_outputs(1833) <= a or b;
    layer3_outputs(1834) <= a and b;
    layer3_outputs(1835) <= a and b;
    layer3_outputs(1836) <= a or b;
    layer3_outputs(1837) <= not a;
    layer3_outputs(1838) <= not b;
    layer3_outputs(1839) <= not a;
    layer3_outputs(1840) <= not b;
    layer3_outputs(1841) <= not b;
    layer3_outputs(1842) <= not (a and b);
    layer3_outputs(1843) <= not b;
    layer3_outputs(1844) <= not (a and b);
    layer3_outputs(1845) <= b and not a;
    layer3_outputs(1846) <= a;
    layer3_outputs(1847) <= a and b;
    layer3_outputs(1848) <= a or b;
    layer3_outputs(1849) <= not a;
    layer3_outputs(1850) <= not (a xor b);
    layer3_outputs(1851) <= a and not b;
    layer3_outputs(1852) <= b and not a;
    layer3_outputs(1853) <= not b;
    layer3_outputs(1854) <= a and b;
    layer3_outputs(1855) <= not a or b;
    layer3_outputs(1856) <= '1';
    layer3_outputs(1857) <= b and not a;
    layer3_outputs(1858) <= not a;
    layer3_outputs(1859) <= b and not a;
    layer3_outputs(1860) <= '0';
    layer3_outputs(1861) <= a and not b;
    layer3_outputs(1862) <= a;
    layer3_outputs(1863) <= a and b;
    layer3_outputs(1864) <= b and not a;
    layer3_outputs(1865) <= b and not a;
    layer3_outputs(1866) <= not b;
    layer3_outputs(1867) <= '1';
    layer3_outputs(1868) <= not (a and b);
    layer3_outputs(1869) <= '0';
    layer3_outputs(1870) <= b;
    layer3_outputs(1871) <= a xor b;
    layer3_outputs(1872) <= not b or a;
    layer3_outputs(1873) <= not b;
    layer3_outputs(1874) <= a and not b;
    layer3_outputs(1875) <= a;
    layer3_outputs(1876) <= not (a or b);
    layer3_outputs(1877) <= b and not a;
    layer3_outputs(1878) <= not (a and b);
    layer3_outputs(1879) <= a or b;
    layer3_outputs(1880) <= a and not b;
    layer3_outputs(1881) <= '0';
    layer3_outputs(1882) <= not (a and b);
    layer3_outputs(1883) <= not b;
    layer3_outputs(1884) <= not (a and b);
    layer3_outputs(1885) <= not (a xor b);
    layer3_outputs(1886) <= a and b;
    layer3_outputs(1887) <= a or b;
    layer3_outputs(1888) <= b and not a;
    layer3_outputs(1889) <= not a;
    layer3_outputs(1890) <= not (a or b);
    layer3_outputs(1891) <= b;
    layer3_outputs(1892) <= b;
    layer3_outputs(1893) <= a;
    layer3_outputs(1894) <= '1';
    layer3_outputs(1895) <= a or b;
    layer3_outputs(1896) <= not b;
    layer3_outputs(1897) <= not b;
    layer3_outputs(1898) <= b;
    layer3_outputs(1899) <= a and not b;
    layer3_outputs(1900) <= a and b;
    layer3_outputs(1901) <= a xor b;
    layer3_outputs(1902) <= a and b;
    layer3_outputs(1903) <= a;
    layer3_outputs(1904) <= a and b;
    layer3_outputs(1905) <= '1';
    layer3_outputs(1906) <= not b;
    layer3_outputs(1907) <= not a or b;
    layer3_outputs(1908) <= not b or a;
    layer3_outputs(1909) <= b and not a;
    layer3_outputs(1910) <= b;
    layer3_outputs(1911) <= a and not b;
    layer3_outputs(1912) <= a and b;
    layer3_outputs(1913) <= a or b;
    layer3_outputs(1914) <= not a or b;
    layer3_outputs(1915) <= b;
    layer3_outputs(1916) <= not (a and b);
    layer3_outputs(1917) <= a and not b;
    layer3_outputs(1918) <= b;
    layer3_outputs(1919) <= '1';
    layer3_outputs(1920) <= b;
    layer3_outputs(1921) <= not (a xor b);
    layer3_outputs(1922) <= b;
    layer3_outputs(1923) <= not a;
    layer3_outputs(1924) <= not b or a;
    layer3_outputs(1925) <= not (a and b);
    layer3_outputs(1926) <= not b;
    layer3_outputs(1927) <= a or b;
    layer3_outputs(1928) <= b and not a;
    layer3_outputs(1929) <= not b or a;
    layer3_outputs(1930) <= not a or b;
    layer3_outputs(1931) <= a;
    layer3_outputs(1932) <= '1';
    layer3_outputs(1933) <= b;
    layer3_outputs(1934) <= '1';
    layer3_outputs(1935) <= not a or b;
    layer3_outputs(1936) <= '1';
    layer3_outputs(1937) <= a or b;
    layer3_outputs(1938) <= '1';
    layer3_outputs(1939) <= not a;
    layer3_outputs(1940) <= a xor b;
    layer3_outputs(1941) <= not a;
    layer3_outputs(1942) <= b and not a;
    layer3_outputs(1943) <= a;
    layer3_outputs(1944) <= b and not a;
    layer3_outputs(1945) <= a;
    layer3_outputs(1946) <= not (a or b);
    layer3_outputs(1947) <= not (a or b);
    layer3_outputs(1948) <= b;
    layer3_outputs(1949) <= not b or a;
    layer3_outputs(1950) <= not b or a;
    layer3_outputs(1951) <= a and not b;
    layer3_outputs(1952) <= not a or b;
    layer3_outputs(1953) <= not a;
    layer3_outputs(1954) <= not (a or b);
    layer3_outputs(1955) <= not a;
    layer3_outputs(1956) <= a and not b;
    layer3_outputs(1957) <= a xor b;
    layer3_outputs(1958) <= b;
    layer3_outputs(1959) <= not (a and b);
    layer3_outputs(1960) <= a or b;
    layer3_outputs(1961) <= not (a xor b);
    layer3_outputs(1962) <= a;
    layer3_outputs(1963) <= a;
    layer3_outputs(1964) <= not a;
    layer3_outputs(1965) <= a;
    layer3_outputs(1966) <= b;
    layer3_outputs(1967) <= a;
    layer3_outputs(1968) <= not (a xor b);
    layer3_outputs(1969) <= a;
    layer3_outputs(1970) <= a and not b;
    layer3_outputs(1971) <= not a;
    layer3_outputs(1972) <= not (a and b);
    layer3_outputs(1973) <= a or b;
    layer3_outputs(1974) <= not (a and b);
    layer3_outputs(1975) <= a and not b;
    layer3_outputs(1976) <= a or b;
    layer3_outputs(1977) <= b and not a;
    layer3_outputs(1978) <= a;
    layer3_outputs(1979) <= b and not a;
    layer3_outputs(1980) <= '1';
    layer3_outputs(1981) <= b and not a;
    layer3_outputs(1982) <= not b;
    layer3_outputs(1983) <= a xor b;
    layer3_outputs(1984) <= '1';
    layer3_outputs(1985) <= a;
    layer3_outputs(1986) <= not (a and b);
    layer3_outputs(1987) <= not (a and b);
    layer3_outputs(1988) <= not a;
    layer3_outputs(1989) <= a or b;
    layer3_outputs(1990) <= not (a and b);
    layer3_outputs(1991) <= not (a or b);
    layer3_outputs(1992) <= not a or b;
    layer3_outputs(1993) <= b and not a;
    layer3_outputs(1994) <= a;
    layer3_outputs(1995) <= a;
    layer3_outputs(1996) <= a and b;
    layer3_outputs(1997) <= b and not a;
    layer3_outputs(1998) <= not b or a;
    layer3_outputs(1999) <= not b;
    layer3_outputs(2000) <= not a;
    layer3_outputs(2001) <= '1';
    layer3_outputs(2002) <= a;
    layer3_outputs(2003) <= a and b;
    layer3_outputs(2004) <= a;
    layer3_outputs(2005) <= not (a or b);
    layer3_outputs(2006) <= not (a and b);
    layer3_outputs(2007) <= not (a or b);
    layer3_outputs(2008) <= a and b;
    layer3_outputs(2009) <= not a;
    layer3_outputs(2010) <= a;
    layer3_outputs(2011) <= not a;
    layer3_outputs(2012) <= b and not a;
    layer3_outputs(2013) <= not (a xor b);
    layer3_outputs(2014) <= not (a and b);
    layer3_outputs(2015) <= a or b;
    layer3_outputs(2016) <= b;
    layer3_outputs(2017) <= not b or a;
    layer3_outputs(2018) <= not a or b;
    layer3_outputs(2019) <= not b;
    layer3_outputs(2020) <= not (a or b);
    layer3_outputs(2021) <= '1';
    layer3_outputs(2022) <= '0';
    layer3_outputs(2023) <= a or b;
    layer3_outputs(2024) <= not b;
    layer3_outputs(2025) <= b and not a;
    layer3_outputs(2026) <= not b;
    layer3_outputs(2027) <= b;
    layer3_outputs(2028) <= not a or b;
    layer3_outputs(2029) <= a xor b;
    layer3_outputs(2030) <= not a;
    layer3_outputs(2031) <= a or b;
    layer3_outputs(2032) <= not (a and b);
    layer3_outputs(2033) <= a;
    layer3_outputs(2034) <= not b;
    layer3_outputs(2035) <= a or b;
    layer3_outputs(2036) <= a and b;
    layer3_outputs(2037) <= a;
    layer3_outputs(2038) <= a xor b;
    layer3_outputs(2039) <= not (a and b);
    layer3_outputs(2040) <= b and not a;
    layer3_outputs(2041) <= b and not a;
    layer3_outputs(2042) <= not b or a;
    layer3_outputs(2043) <= '1';
    layer3_outputs(2044) <= not b;
    layer3_outputs(2045) <= not (a and b);
    layer3_outputs(2046) <= not (a or b);
    layer3_outputs(2047) <= b;
    layer3_outputs(2048) <= not a;
    layer3_outputs(2049) <= not (a xor b);
    layer3_outputs(2050) <= a;
    layer3_outputs(2051) <= a;
    layer3_outputs(2052) <= not a;
    layer3_outputs(2053) <= b and not a;
    layer3_outputs(2054) <= not b;
    layer3_outputs(2055) <= not b;
    layer3_outputs(2056) <= not b;
    layer3_outputs(2057) <= not (a and b);
    layer3_outputs(2058) <= '0';
    layer3_outputs(2059) <= not b or a;
    layer3_outputs(2060) <= not b or a;
    layer3_outputs(2061) <= not a;
    layer3_outputs(2062) <= '0';
    layer3_outputs(2063) <= a;
    layer3_outputs(2064) <= a xor b;
    layer3_outputs(2065) <= a and b;
    layer3_outputs(2066) <= not (a xor b);
    layer3_outputs(2067) <= not (a or b);
    layer3_outputs(2068) <= a;
    layer3_outputs(2069) <= not b;
    layer3_outputs(2070) <= b and not a;
    layer3_outputs(2071) <= a;
    layer3_outputs(2072) <= a and b;
    layer3_outputs(2073) <= a or b;
    layer3_outputs(2074) <= not a;
    layer3_outputs(2075) <= not (a and b);
    layer3_outputs(2076) <= not (a or b);
    layer3_outputs(2077) <= b;
    layer3_outputs(2078) <= a;
    layer3_outputs(2079) <= not b or a;
    layer3_outputs(2080) <= b;
    layer3_outputs(2081) <= a xor b;
    layer3_outputs(2082) <= not b;
    layer3_outputs(2083) <= not a or b;
    layer3_outputs(2084) <= a and b;
    layer3_outputs(2085) <= not (a or b);
    layer3_outputs(2086) <= a;
    layer3_outputs(2087) <= not b;
    layer3_outputs(2088) <= not a;
    layer3_outputs(2089) <= a;
    layer3_outputs(2090) <= not a;
    layer3_outputs(2091) <= a and b;
    layer3_outputs(2092) <= not a or b;
    layer3_outputs(2093) <= b;
    layer3_outputs(2094) <= a and b;
    layer3_outputs(2095) <= a or b;
    layer3_outputs(2096) <= b;
    layer3_outputs(2097) <= '0';
    layer3_outputs(2098) <= not a or b;
    layer3_outputs(2099) <= '0';
    layer3_outputs(2100) <= not a or b;
    layer3_outputs(2101) <= '1';
    layer3_outputs(2102) <= a or b;
    layer3_outputs(2103) <= not a;
    layer3_outputs(2104) <= a and b;
    layer3_outputs(2105) <= a and not b;
    layer3_outputs(2106) <= not (a or b);
    layer3_outputs(2107) <= '0';
    layer3_outputs(2108) <= b;
    layer3_outputs(2109) <= not (a xor b);
    layer3_outputs(2110) <= a;
    layer3_outputs(2111) <= b;
    layer3_outputs(2112) <= a;
    layer3_outputs(2113) <= not a;
    layer3_outputs(2114) <= '0';
    layer3_outputs(2115) <= not b or a;
    layer3_outputs(2116) <= b and not a;
    layer3_outputs(2117) <= not (a or b);
    layer3_outputs(2118) <= a;
    layer3_outputs(2119) <= not a;
    layer3_outputs(2120) <= not (a xor b);
    layer3_outputs(2121) <= a and not b;
    layer3_outputs(2122) <= a or b;
    layer3_outputs(2123) <= a xor b;
    layer3_outputs(2124) <= a xor b;
    layer3_outputs(2125) <= not (a and b);
    layer3_outputs(2126) <= not a or b;
    layer3_outputs(2127) <= a;
    layer3_outputs(2128) <= not (a and b);
    layer3_outputs(2129) <= a and b;
    layer3_outputs(2130) <= a and not b;
    layer3_outputs(2131) <= a xor b;
    layer3_outputs(2132) <= not b;
    layer3_outputs(2133) <= a and b;
    layer3_outputs(2134) <= not a;
    layer3_outputs(2135) <= '0';
    layer3_outputs(2136) <= b and not a;
    layer3_outputs(2137) <= a or b;
    layer3_outputs(2138) <= a;
    layer3_outputs(2139) <= b;
    layer3_outputs(2140) <= not (a or b);
    layer3_outputs(2141) <= a;
    layer3_outputs(2142) <= '1';
    layer3_outputs(2143) <= not a;
    layer3_outputs(2144) <= not b;
    layer3_outputs(2145) <= a;
    layer3_outputs(2146) <= a;
    layer3_outputs(2147) <= a and b;
    layer3_outputs(2148) <= b;
    layer3_outputs(2149) <= not (a xor b);
    layer3_outputs(2150) <= a;
    layer3_outputs(2151) <= not (a xor b);
    layer3_outputs(2152) <= a and b;
    layer3_outputs(2153) <= not b or a;
    layer3_outputs(2154) <= not a or b;
    layer3_outputs(2155) <= not (a or b);
    layer3_outputs(2156) <= a;
    layer3_outputs(2157) <= '1';
    layer3_outputs(2158) <= not a;
    layer3_outputs(2159) <= a;
    layer3_outputs(2160) <= b;
    layer3_outputs(2161) <= not (a and b);
    layer3_outputs(2162) <= b;
    layer3_outputs(2163) <= not a or b;
    layer3_outputs(2164) <= a or b;
    layer3_outputs(2165) <= b;
    layer3_outputs(2166) <= a or b;
    layer3_outputs(2167) <= not b;
    layer3_outputs(2168) <= not b or a;
    layer3_outputs(2169) <= a and b;
    layer3_outputs(2170) <= a and not b;
    layer3_outputs(2171) <= a;
    layer3_outputs(2172) <= not b or a;
    layer3_outputs(2173) <= a or b;
    layer3_outputs(2174) <= '0';
    layer3_outputs(2175) <= '0';
    layer3_outputs(2176) <= not (a xor b);
    layer3_outputs(2177) <= not b;
    layer3_outputs(2178) <= a;
    layer3_outputs(2179) <= not a;
    layer3_outputs(2180) <= a or b;
    layer3_outputs(2181) <= not a;
    layer3_outputs(2182) <= a;
    layer3_outputs(2183) <= not (a or b);
    layer3_outputs(2184) <= b and not a;
    layer3_outputs(2185) <= a and b;
    layer3_outputs(2186) <= not a or b;
    layer3_outputs(2187) <= a;
    layer3_outputs(2188) <= not (a or b);
    layer3_outputs(2189) <= '0';
    layer3_outputs(2190) <= a;
    layer3_outputs(2191) <= not a or b;
    layer3_outputs(2192) <= not a or b;
    layer3_outputs(2193) <= a;
    layer3_outputs(2194) <= a and b;
    layer3_outputs(2195) <= not b;
    layer3_outputs(2196) <= not a or b;
    layer3_outputs(2197) <= a and b;
    layer3_outputs(2198) <= not (a or b);
    layer3_outputs(2199) <= not b;
    layer3_outputs(2200) <= not (a or b);
    layer3_outputs(2201) <= a and b;
    layer3_outputs(2202) <= a;
    layer3_outputs(2203) <= a or b;
    layer3_outputs(2204) <= not (a and b);
    layer3_outputs(2205) <= '1';
    layer3_outputs(2206) <= a;
    layer3_outputs(2207) <= a and not b;
    layer3_outputs(2208) <= b;
    layer3_outputs(2209) <= not a or b;
    layer3_outputs(2210) <= '1';
    layer3_outputs(2211) <= a and not b;
    layer3_outputs(2212) <= a;
    layer3_outputs(2213) <= not a;
    layer3_outputs(2214) <= a and b;
    layer3_outputs(2215) <= not (a xor b);
    layer3_outputs(2216) <= not (a and b);
    layer3_outputs(2217) <= not a or b;
    layer3_outputs(2218) <= b;
    layer3_outputs(2219) <= b;
    layer3_outputs(2220) <= a and b;
    layer3_outputs(2221) <= not a or b;
    layer3_outputs(2222) <= not (a or b);
    layer3_outputs(2223) <= not (a and b);
    layer3_outputs(2224) <= not b;
    layer3_outputs(2225) <= not a;
    layer3_outputs(2226) <= a and b;
    layer3_outputs(2227) <= a or b;
    layer3_outputs(2228) <= b;
    layer3_outputs(2229) <= not b;
    layer3_outputs(2230) <= not b or a;
    layer3_outputs(2231) <= '1';
    layer3_outputs(2232) <= not (a and b);
    layer3_outputs(2233) <= b;
    layer3_outputs(2234) <= '1';
    layer3_outputs(2235) <= a;
    layer3_outputs(2236) <= a and not b;
    layer3_outputs(2237) <= a or b;
    layer3_outputs(2238) <= a and b;
    layer3_outputs(2239) <= not (a xor b);
    layer3_outputs(2240) <= not a;
    layer3_outputs(2241) <= b;
    layer3_outputs(2242) <= not a;
    layer3_outputs(2243) <= not b;
    layer3_outputs(2244) <= a and not b;
    layer3_outputs(2245) <= a or b;
    layer3_outputs(2246) <= b;
    layer3_outputs(2247) <= not (a and b);
    layer3_outputs(2248) <= not b;
    layer3_outputs(2249) <= a xor b;
    layer3_outputs(2250) <= a or b;
    layer3_outputs(2251) <= a xor b;
    layer3_outputs(2252) <= not a;
    layer3_outputs(2253) <= b and not a;
    layer3_outputs(2254) <= not a;
    layer3_outputs(2255) <= not a or b;
    layer3_outputs(2256) <= b;
    layer3_outputs(2257) <= a;
    layer3_outputs(2258) <= not (a xor b);
    layer3_outputs(2259) <= '0';
    layer3_outputs(2260) <= a and b;
    layer3_outputs(2261) <= a;
    layer3_outputs(2262) <= not a;
    layer3_outputs(2263) <= not (a or b);
    layer3_outputs(2264) <= '1';
    layer3_outputs(2265) <= a or b;
    layer3_outputs(2266) <= not b or a;
    layer3_outputs(2267) <= not (a or b);
    layer3_outputs(2268) <= not b;
    layer3_outputs(2269) <= not (a or b);
    layer3_outputs(2270) <= b and not a;
    layer3_outputs(2271) <= b;
    layer3_outputs(2272) <= not b;
    layer3_outputs(2273) <= not a;
    layer3_outputs(2274) <= not a or b;
    layer3_outputs(2275) <= b;
    layer3_outputs(2276) <= not a;
    layer3_outputs(2277) <= a;
    layer3_outputs(2278) <= not b;
    layer3_outputs(2279) <= a;
    layer3_outputs(2280) <= a;
    layer3_outputs(2281) <= '1';
    layer3_outputs(2282) <= b and not a;
    layer3_outputs(2283) <= not (a xor b);
    layer3_outputs(2284) <= not (a and b);
    layer3_outputs(2285) <= a and b;
    layer3_outputs(2286) <= a;
    layer3_outputs(2287) <= a and b;
    layer3_outputs(2288) <= not (a xor b);
    layer3_outputs(2289) <= a;
    layer3_outputs(2290) <= a or b;
    layer3_outputs(2291) <= not a;
    layer3_outputs(2292) <= not (a or b);
    layer3_outputs(2293) <= not a;
    layer3_outputs(2294) <= not (a xor b);
    layer3_outputs(2295) <= not b;
    layer3_outputs(2296) <= b;
    layer3_outputs(2297) <= not a;
    layer3_outputs(2298) <= a or b;
    layer3_outputs(2299) <= not b or a;
    layer3_outputs(2300) <= not (a xor b);
    layer3_outputs(2301) <= a and not b;
    layer3_outputs(2302) <= not (a or b);
    layer3_outputs(2303) <= b;
    layer3_outputs(2304) <= a and b;
    layer3_outputs(2305) <= not b;
    layer3_outputs(2306) <= a xor b;
    layer3_outputs(2307) <= a or b;
    layer3_outputs(2308) <= not (a or b);
    layer3_outputs(2309) <= a and not b;
    layer3_outputs(2310) <= a or b;
    layer3_outputs(2311) <= not a;
    layer3_outputs(2312) <= a;
    layer3_outputs(2313) <= a and b;
    layer3_outputs(2314) <= not (a and b);
    layer3_outputs(2315) <= not a or b;
    layer3_outputs(2316) <= b and not a;
    layer3_outputs(2317) <= b;
    layer3_outputs(2318) <= not (a or b);
    layer3_outputs(2319) <= b;
    layer3_outputs(2320) <= a xor b;
    layer3_outputs(2321) <= not (a xor b);
    layer3_outputs(2322) <= '0';
    layer3_outputs(2323) <= not b or a;
    layer3_outputs(2324) <= not a;
    layer3_outputs(2325) <= not (a and b);
    layer3_outputs(2326) <= not a or b;
    layer3_outputs(2327) <= not (a or b);
    layer3_outputs(2328) <= a and not b;
    layer3_outputs(2329) <= a;
    layer3_outputs(2330) <= b and not a;
    layer3_outputs(2331) <= b;
    layer3_outputs(2332) <= a and not b;
    layer3_outputs(2333) <= a or b;
    layer3_outputs(2334) <= not (a xor b);
    layer3_outputs(2335) <= a and not b;
    layer3_outputs(2336) <= '0';
    layer3_outputs(2337) <= not b;
    layer3_outputs(2338) <= a and b;
    layer3_outputs(2339) <= a and not b;
    layer3_outputs(2340) <= a or b;
    layer3_outputs(2341) <= not (a or b);
    layer3_outputs(2342) <= a;
    layer3_outputs(2343) <= a xor b;
    layer3_outputs(2344) <= not (a xor b);
    layer3_outputs(2345) <= a xor b;
    layer3_outputs(2346) <= a xor b;
    layer3_outputs(2347) <= not (a and b);
    layer3_outputs(2348) <= a and b;
    layer3_outputs(2349) <= a and b;
    layer3_outputs(2350) <= a and not b;
    layer3_outputs(2351) <= a or b;
    layer3_outputs(2352) <= not a;
    layer3_outputs(2353) <= b;
    layer3_outputs(2354) <= b;
    layer3_outputs(2355) <= not a;
    layer3_outputs(2356) <= a;
    layer3_outputs(2357) <= not b or a;
    layer3_outputs(2358) <= not a;
    layer3_outputs(2359) <= a or b;
    layer3_outputs(2360) <= '0';
    layer3_outputs(2361) <= b;
    layer3_outputs(2362) <= not (a and b);
    layer3_outputs(2363) <= not b or a;
    layer3_outputs(2364) <= not a;
    layer3_outputs(2365) <= '0';
    layer3_outputs(2366) <= a or b;
    layer3_outputs(2367) <= not a;
    layer3_outputs(2368) <= not b;
    layer3_outputs(2369) <= not (a or b);
    layer3_outputs(2370) <= b;
    layer3_outputs(2371) <= not b;
    layer3_outputs(2372) <= not b;
    layer3_outputs(2373) <= '1';
    layer3_outputs(2374) <= not a;
    layer3_outputs(2375) <= not b;
    layer3_outputs(2376) <= a and not b;
    layer3_outputs(2377) <= a and not b;
    layer3_outputs(2378) <= not a;
    layer3_outputs(2379) <= not b;
    layer3_outputs(2380) <= a and not b;
    layer3_outputs(2381) <= not b;
    layer3_outputs(2382) <= not (a or b);
    layer3_outputs(2383) <= a and b;
    layer3_outputs(2384) <= a;
    layer3_outputs(2385) <= not (a or b);
    layer3_outputs(2386) <= b;
    layer3_outputs(2387) <= not a;
    layer3_outputs(2388) <= not b or a;
    layer3_outputs(2389) <= a;
    layer3_outputs(2390) <= a and not b;
    layer3_outputs(2391) <= not b;
    layer3_outputs(2392) <= b;
    layer3_outputs(2393) <= not b;
    layer3_outputs(2394) <= not (a xor b);
    layer3_outputs(2395) <= not b;
    layer3_outputs(2396) <= a and not b;
    layer3_outputs(2397) <= not (a and b);
    layer3_outputs(2398) <= not b;
    layer3_outputs(2399) <= a and b;
    layer3_outputs(2400) <= a or b;
    layer3_outputs(2401) <= a and not b;
    layer3_outputs(2402) <= b;
    layer3_outputs(2403) <= not a or b;
    layer3_outputs(2404) <= a;
    layer3_outputs(2405) <= not b;
    layer3_outputs(2406) <= '1';
    layer3_outputs(2407) <= a and not b;
    layer3_outputs(2408) <= not a or b;
    layer3_outputs(2409) <= not b or a;
    layer3_outputs(2410) <= b;
    layer3_outputs(2411) <= not b;
    layer3_outputs(2412) <= not b;
    layer3_outputs(2413) <= not a;
    layer3_outputs(2414) <= not b;
    layer3_outputs(2415) <= '1';
    layer3_outputs(2416) <= b and not a;
    layer3_outputs(2417) <= a;
    layer3_outputs(2418) <= b;
    layer3_outputs(2419) <= not (a or b);
    layer3_outputs(2420) <= a and not b;
    layer3_outputs(2421) <= not b;
    layer3_outputs(2422) <= a xor b;
    layer3_outputs(2423) <= a xor b;
    layer3_outputs(2424) <= not b;
    layer3_outputs(2425) <= not b or a;
    layer3_outputs(2426) <= a xor b;
    layer3_outputs(2427) <= a xor b;
    layer3_outputs(2428) <= not b;
    layer3_outputs(2429) <= a;
    layer3_outputs(2430) <= a and not b;
    layer3_outputs(2431) <= b;
    layer3_outputs(2432) <= not (a and b);
    layer3_outputs(2433) <= a or b;
    layer3_outputs(2434) <= not b;
    layer3_outputs(2435) <= not a or b;
    layer3_outputs(2436) <= b and not a;
    layer3_outputs(2437) <= '0';
    layer3_outputs(2438) <= not (a xor b);
    layer3_outputs(2439) <= a;
    layer3_outputs(2440) <= b;
    layer3_outputs(2441) <= not a;
    layer3_outputs(2442) <= '1';
    layer3_outputs(2443) <= not a;
    layer3_outputs(2444) <= a or b;
    layer3_outputs(2445) <= not (a or b);
    layer3_outputs(2446) <= a;
    layer3_outputs(2447) <= a;
    layer3_outputs(2448) <= a and not b;
    layer3_outputs(2449) <= not b or a;
    layer3_outputs(2450) <= b and not a;
    layer3_outputs(2451) <= a and not b;
    layer3_outputs(2452) <= a and b;
    layer3_outputs(2453) <= not a;
    layer3_outputs(2454) <= a;
    layer3_outputs(2455) <= '0';
    layer3_outputs(2456) <= a;
    layer3_outputs(2457) <= not (a and b);
    layer3_outputs(2458) <= not a;
    layer3_outputs(2459) <= not b or a;
    layer3_outputs(2460) <= '0';
    layer3_outputs(2461) <= a xor b;
    layer3_outputs(2462) <= not (a and b);
    layer3_outputs(2463) <= '1';
    layer3_outputs(2464) <= a and not b;
    layer3_outputs(2465) <= a and b;
    layer3_outputs(2466) <= b;
    layer3_outputs(2467) <= not b;
    layer3_outputs(2468) <= not a;
    layer3_outputs(2469) <= a and not b;
    layer3_outputs(2470) <= not b or a;
    layer3_outputs(2471) <= '0';
    layer3_outputs(2472) <= a;
    layer3_outputs(2473) <= not b or a;
    layer3_outputs(2474) <= a;
    layer3_outputs(2475) <= not b;
    layer3_outputs(2476) <= a and b;
    layer3_outputs(2477) <= a and b;
    layer3_outputs(2478) <= not b or a;
    layer3_outputs(2479) <= not (a and b);
    layer3_outputs(2480) <= a;
    layer3_outputs(2481) <= not a;
    layer3_outputs(2482) <= '0';
    layer3_outputs(2483) <= a and b;
    layer3_outputs(2484) <= not (a xor b);
    layer3_outputs(2485) <= not (a and b);
    layer3_outputs(2486) <= a xor b;
    layer3_outputs(2487) <= b;
    layer3_outputs(2488) <= not a;
    layer3_outputs(2489) <= a;
    layer3_outputs(2490) <= not b or a;
    layer3_outputs(2491) <= not b;
    layer3_outputs(2492) <= a;
    layer3_outputs(2493) <= b;
    layer3_outputs(2494) <= not a;
    layer3_outputs(2495) <= b;
    layer3_outputs(2496) <= a and not b;
    layer3_outputs(2497) <= '1';
    layer3_outputs(2498) <= a xor b;
    layer3_outputs(2499) <= not (a and b);
    layer3_outputs(2500) <= b and not a;
    layer3_outputs(2501) <= b and not a;
    layer3_outputs(2502) <= not (a and b);
    layer3_outputs(2503) <= not b or a;
    layer3_outputs(2504) <= a;
    layer3_outputs(2505) <= not a or b;
    layer3_outputs(2506) <= a;
    layer3_outputs(2507) <= '0';
    layer3_outputs(2508) <= not b;
    layer3_outputs(2509) <= b and not a;
    layer3_outputs(2510) <= not b;
    layer3_outputs(2511) <= not (a xor b);
    layer3_outputs(2512) <= not b;
    layer3_outputs(2513) <= not a or b;
    layer3_outputs(2514) <= b;
    layer3_outputs(2515) <= a;
    layer3_outputs(2516) <= not a;
    layer3_outputs(2517) <= a and b;
    layer3_outputs(2518) <= b and not a;
    layer3_outputs(2519) <= not b or a;
    layer3_outputs(2520) <= a or b;
    layer3_outputs(2521) <= a and b;
    layer3_outputs(2522) <= a;
    layer3_outputs(2523) <= not a or b;
    layer3_outputs(2524) <= a and b;
    layer3_outputs(2525) <= not a or b;
    layer3_outputs(2526) <= a;
    layer3_outputs(2527) <= a xor b;
    layer3_outputs(2528) <= '1';
    layer3_outputs(2529) <= a and b;
    layer3_outputs(2530) <= b;
    layer3_outputs(2531) <= not b or a;
    layer3_outputs(2532) <= not b;
    layer3_outputs(2533) <= not (a and b);
    layer3_outputs(2534) <= not (a or b);
    layer3_outputs(2535) <= not b;
    layer3_outputs(2536) <= b;
    layer3_outputs(2537) <= not a;
    layer3_outputs(2538) <= not (a and b);
    layer3_outputs(2539) <= a xor b;
    layer3_outputs(2540) <= not (a or b);
    layer3_outputs(2541) <= not b;
    layer3_outputs(2542) <= not (a and b);
    layer3_outputs(2543) <= not (a or b);
    layer3_outputs(2544) <= b and not a;
    layer3_outputs(2545) <= not a;
    layer3_outputs(2546) <= b and not a;
    layer3_outputs(2547) <= not a or b;
    layer3_outputs(2548) <= a and b;
    layer3_outputs(2549) <= not (a or b);
    layer3_outputs(2550) <= a or b;
    layer3_outputs(2551) <= a or b;
    layer3_outputs(2552) <= b;
    layer3_outputs(2553) <= not a;
    layer3_outputs(2554) <= not a or b;
    layer3_outputs(2555) <= a;
    layer3_outputs(2556) <= not (a and b);
    layer3_outputs(2557) <= not (a xor b);
    layer3_outputs(2558) <= not b or a;
    layer3_outputs(2559) <= not a;
    layer3_outputs(2560) <= b and not a;
    layer3_outputs(2561) <= b;
    layer3_outputs(2562) <= a and not b;
    layer3_outputs(2563) <= not b;
    layer3_outputs(2564) <= not b or a;
    layer3_outputs(2565) <= b and not a;
    layer3_outputs(2566) <= not (a or b);
    layer3_outputs(2567) <= not (a or b);
    layer3_outputs(2568) <= a;
    layer3_outputs(2569) <= not b;
    layer3_outputs(2570) <= not (a or b);
    layer3_outputs(2571) <= '0';
    layer3_outputs(2572) <= '0';
    layer3_outputs(2573) <= '1';
    layer3_outputs(2574) <= b and not a;
    layer3_outputs(2575) <= not b;
    layer3_outputs(2576) <= b;
    layer3_outputs(2577) <= b;
    layer3_outputs(2578) <= not b;
    layer3_outputs(2579) <= not a or b;
    layer3_outputs(2580) <= a and not b;
    layer3_outputs(2581) <= not (a xor b);
    layer3_outputs(2582) <= not (a and b);
    layer3_outputs(2583) <= '1';
    layer3_outputs(2584) <= a and b;
    layer3_outputs(2585) <= b;
    layer3_outputs(2586) <= '1';
    layer3_outputs(2587) <= not a or b;
    layer3_outputs(2588) <= not (a and b);
    layer3_outputs(2589) <= not b or a;
    layer3_outputs(2590) <= not a or b;
    layer3_outputs(2591) <= not (a and b);
    layer3_outputs(2592) <= b and not a;
    layer3_outputs(2593) <= not (a or b);
    layer3_outputs(2594) <= a and b;
    layer3_outputs(2595) <= not a;
    layer3_outputs(2596) <= not b;
    layer3_outputs(2597) <= not (a and b);
    layer3_outputs(2598) <= not b or a;
    layer3_outputs(2599) <= a or b;
    layer3_outputs(2600) <= not b;
    layer3_outputs(2601) <= a;
    layer3_outputs(2602) <= not a or b;
    layer3_outputs(2603) <= not (a and b);
    layer3_outputs(2604) <= a;
    layer3_outputs(2605) <= not (a or b);
    layer3_outputs(2606) <= not (a xor b);
    layer3_outputs(2607) <= not b;
    layer3_outputs(2608) <= not a or b;
    layer3_outputs(2609) <= not (a and b);
    layer3_outputs(2610) <= a or b;
    layer3_outputs(2611) <= not b;
    layer3_outputs(2612) <= not a or b;
    layer3_outputs(2613) <= b and not a;
    layer3_outputs(2614) <= not a;
    layer3_outputs(2615) <= not (a or b);
    layer3_outputs(2616) <= not (a or b);
    layer3_outputs(2617) <= not a;
    layer3_outputs(2618) <= not b or a;
    layer3_outputs(2619) <= not b or a;
    layer3_outputs(2620) <= a;
    layer3_outputs(2621) <= not (a xor b);
    layer3_outputs(2622) <= a or b;
    layer3_outputs(2623) <= not a;
    layer3_outputs(2624) <= b and not a;
    layer3_outputs(2625) <= not (a or b);
    layer3_outputs(2626) <= a;
    layer3_outputs(2627) <= not a;
    layer3_outputs(2628) <= '1';
    layer3_outputs(2629) <= not a;
    layer3_outputs(2630) <= a and b;
    layer3_outputs(2631) <= not b or a;
    layer3_outputs(2632) <= not a;
    layer3_outputs(2633) <= not (a and b);
    layer3_outputs(2634) <= b;
    layer3_outputs(2635) <= b and not a;
    layer3_outputs(2636) <= not (a xor b);
    layer3_outputs(2637) <= not a;
    layer3_outputs(2638) <= not (a or b);
    layer3_outputs(2639) <= not a;
    layer3_outputs(2640) <= a and b;
    layer3_outputs(2641) <= a and not b;
    layer3_outputs(2642) <= b and not a;
    layer3_outputs(2643) <= b and not a;
    layer3_outputs(2644) <= a and not b;
    layer3_outputs(2645) <= not (a xor b);
    layer3_outputs(2646) <= not (a and b);
    layer3_outputs(2647) <= b and not a;
    layer3_outputs(2648) <= not a or b;
    layer3_outputs(2649) <= not b or a;
    layer3_outputs(2650) <= not a;
    layer3_outputs(2651) <= b and not a;
    layer3_outputs(2652) <= not a;
    layer3_outputs(2653) <= a and b;
    layer3_outputs(2654) <= '0';
    layer3_outputs(2655) <= '0';
    layer3_outputs(2656) <= not b or a;
    layer3_outputs(2657) <= a;
    layer3_outputs(2658) <= not b;
    layer3_outputs(2659) <= not (a or b);
    layer3_outputs(2660) <= a xor b;
    layer3_outputs(2661) <= not b or a;
    layer3_outputs(2662) <= b;
    layer3_outputs(2663) <= a or b;
    layer3_outputs(2664) <= a and not b;
    layer3_outputs(2665) <= not b;
    layer3_outputs(2666) <= not (a xor b);
    layer3_outputs(2667) <= not (a and b);
    layer3_outputs(2668) <= not b;
    layer3_outputs(2669) <= not (a and b);
    layer3_outputs(2670) <= a;
    layer3_outputs(2671) <= a;
    layer3_outputs(2672) <= not a;
    layer3_outputs(2673) <= '0';
    layer3_outputs(2674) <= not b or a;
    layer3_outputs(2675) <= a;
    layer3_outputs(2676) <= not (a or b);
    layer3_outputs(2677) <= not (a and b);
    layer3_outputs(2678) <= '1';
    layer3_outputs(2679) <= '1';
    layer3_outputs(2680) <= '1';
    layer3_outputs(2681) <= b and not a;
    layer3_outputs(2682) <= '0';
    layer3_outputs(2683) <= a;
    layer3_outputs(2684) <= not b;
    layer3_outputs(2685) <= b;
    layer3_outputs(2686) <= b;
    layer3_outputs(2687) <= not a;
    layer3_outputs(2688) <= a;
    layer3_outputs(2689) <= not a;
    layer3_outputs(2690) <= not (a and b);
    layer3_outputs(2691) <= a or b;
    layer3_outputs(2692) <= not a;
    layer3_outputs(2693) <= not a;
    layer3_outputs(2694) <= b and not a;
    layer3_outputs(2695) <= not (a and b);
    layer3_outputs(2696) <= '0';
    layer3_outputs(2697) <= not (a or b);
    layer3_outputs(2698) <= a xor b;
    layer3_outputs(2699) <= not b;
    layer3_outputs(2700) <= b;
    layer3_outputs(2701) <= not b or a;
    layer3_outputs(2702) <= not (a xor b);
    layer3_outputs(2703) <= not a or b;
    layer3_outputs(2704) <= not (a or b);
    layer3_outputs(2705) <= a and not b;
    layer3_outputs(2706) <= b and not a;
    layer3_outputs(2707) <= '0';
    layer3_outputs(2708) <= '0';
    layer3_outputs(2709) <= not a;
    layer3_outputs(2710) <= a;
    layer3_outputs(2711) <= a and b;
    layer3_outputs(2712) <= a xor b;
    layer3_outputs(2713) <= not (a xor b);
    layer3_outputs(2714) <= '0';
    layer3_outputs(2715) <= a and not b;
    layer3_outputs(2716) <= a and not b;
    layer3_outputs(2717) <= not a;
    layer3_outputs(2718) <= not b;
    layer3_outputs(2719) <= not b;
    layer3_outputs(2720) <= not (a and b);
    layer3_outputs(2721) <= not a;
    layer3_outputs(2722) <= not a;
    layer3_outputs(2723) <= a or b;
    layer3_outputs(2724) <= a;
    layer3_outputs(2725) <= '0';
    layer3_outputs(2726) <= a xor b;
    layer3_outputs(2727) <= a or b;
    layer3_outputs(2728) <= a and b;
    layer3_outputs(2729) <= not a or b;
    layer3_outputs(2730) <= not b;
    layer3_outputs(2731) <= a and b;
    layer3_outputs(2732) <= not a;
    layer3_outputs(2733) <= '1';
    layer3_outputs(2734) <= not a;
    layer3_outputs(2735) <= a xor b;
    layer3_outputs(2736) <= a and b;
    layer3_outputs(2737) <= not (a or b);
    layer3_outputs(2738) <= a and not b;
    layer3_outputs(2739) <= not (a or b);
    layer3_outputs(2740) <= not (a xor b);
    layer3_outputs(2741) <= not a;
    layer3_outputs(2742) <= b;
    layer3_outputs(2743) <= b;
    layer3_outputs(2744) <= a;
    layer3_outputs(2745) <= a or b;
    layer3_outputs(2746) <= not b or a;
    layer3_outputs(2747) <= not (a or b);
    layer3_outputs(2748) <= a xor b;
    layer3_outputs(2749) <= not (a and b);
    layer3_outputs(2750) <= '0';
    layer3_outputs(2751) <= not (a and b);
    layer3_outputs(2752) <= not b;
    layer3_outputs(2753) <= a;
    layer3_outputs(2754) <= a and not b;
    layer3_outputs(2755) <= not a or b;
    layer3_outputs(2756) <= not a;
    layer3_outputs(2757) <= b;
    layer3_outputs(2758) <= b and not a;
    layer3_outputs(2759) <= a;
    layer3_outputs(2760) <= not (a xor b);
    layer3_outputs(2761) <= not a or b;
    layer3_outputs(2762) <= not a;
    layer3_outputs(2763) <= b and not a;
    layer3_outputs(2764) <= b and not a;
    layer3_outputs(2765) <= not (a and b);
    layer3_outputs(2766) <= a;
    layer3_outputs(2767) <= a and b;
    layer3_outputs(2768) <= not a;
    layer3_outputs(2769) <= a xor b;
    layer3_outputs(2770) <= b;
    layer3_outputs(2771) <= not b;
    layer3_outputs(2772) <= a and not b;
    layer3_outputs(2773) <= a and not b;
    layer3_outputs(2774) <= not (a or b);
    layer3_outputs(2775) <= a and b;
    layer3_outputs(2776) <= a and not b;
    layer3_outputs(2777) <= b;
    layer3_outputs(2778) <= not (a xor b);
    layer3_outputs(2779) <= not b;
    layer3_outputs(2780) <= a and not b;
    layer3_outputs(2781) <= not a;
    layer3_outputs(2782) <= a;
    layer3_outputs(2783) <= not (a xor b);
    layer3_outputs(2784) <= a or b;
    layer3_outputs(2785) <= not (a and b);
    layer3_outputs(2786) <= not a or b;
    layer3_outputs(2787) <= b and not a;
    layer3_outputs(2788) <= b and not a;
    layer3_outputs(2789) <= not a or b;
    layer3_outputs(2790) <= not b or a;
    layer3_outputs(2791) <= not b;
    layer3_outputs(2792) <= not b or a;
    layer3_outputs(2793) <= '1';
    layer3_outputs(2794) <= not b;
    layer3_outputs(2795) <= not (a and b);
    layer3_outputs(2796) <= not (a or b);
    layer3_outputs(2797) <= '0';
    layer3_outputs(2798) <= b and not a;
    layer3_outputs(2799) <= not a or b;
    layer3_outputs(2800) <= not b;
    layer3_outputs(2801) <= not (a or b);
    layer3_outputs(2802) <= not (a and b);
    layer3_outputs(2803) <= a;
    layer3_outputs(2804) <= not (a and b);
    layer3_outputs(2805) <= not a or b;
    layer3_outputs(2806) <= a or b;
    layer3_outputs(2807) <= a and b;
    layer3_outputs(2808) <= a;
    layer3_outputs(2809) <= not a or b;
    layer3_outputs(2810) <= b and not a;
    layer3_outputs(2811) <= a and b;
    layer3_outputs(2812) <= a;
    layer3_outputs(2813) <= a;
    layer3_outputs(2814) <= a and b;
    layer3_outputs(2815) <= a and b;
    layer3_outputs(2816) <= a and b;
    layer3_outputs(2817) <= not b or a;
    layer3_outputs(2818) <= b and not a;
    layer3_outputs(2819) <= a and not b;
    layer3_outputs(2820) <= b and not a;
    layer3_outputs(2821) <= a or b;
    layer3_outputs(2822) <= not a;
    layer3_outputs(2823) <= b;
    layer3_outputs(2824) <= a and not b;
    layer3_outputs(2825) <= not a;
    layer3_outputs(2826) <= b;
    layer3_outputs(2827) <= '1';
    layer3_outputs(2828) <= b;
    layer3_outputs(2829) <= a and not b;
    layer3_outputs(2830) <= '1';
    layer3_outputs(2831) <= not a;
    layer3_outputs(2832) <= b;
    layer3_outputs(2833) <= a or b;
    layer3_outputs(2834) <= b;
    layer3_outputs(2835) <= a and b;
    layer3_outputs(2836) <= a and b;
    layer3_outputs(2837) <= not (a or b);
    layer3_outputs(2838) <= a;
    layer3_outputs(2839) <= '1';
    layer3_outputs(2840) <= a xor b;
    layer3_outputs(2841) <= a;
    layer3_outputs(2842) <= not b;
    layer3_outputs(2843) <= b;
    layer3_outputs(2844) <= not b or a;
    layer3_outputs(2845) <= b and not a;
    layer3_outputs(2846) <= a;
    layer3_outputs(2847) <= a;
    layer3_outputs(2848) <= a or b;
    layer3_outputs(2849) <= b;
    layer3_outputs(2850) <= not a;
    layer3_outputs(2851) <= not a;
    layer3_outputs(2852) <= a;
    layer3_outputs(2853) <= '0';
    layer3_outputs(2854) <= b;
    layer3_outputs(2855) <= a and b;
    layer3_outputs(2856) <= b;
    layer3_outputs(2857) <= a and not b;
    layer3_outputs(2858) <= a;
    layer3_outputs(2859) <= a;
    layer3_outputs(2860) <= b;
    layer3_outputs(2861) <= a;
    layer3_outputs(2862) <= not a or b;
    layer3_outputs(2863) <= not a;
    layer3_outputs(2864) <= not (a or b);
    layer3_outputs(2865) <= b;
    layer3_outputs(2866) <= not a;
    layer3_outputs(2867) <= not b;
    layer3_outputs(2868) <= a or b;
    layer3_outputs(2869) <= b;
    layer3_outputs(2870) <= not (a xor b);
    layer3_outputs(2871) <= not b;
    layer3_outputs(2872) <= a;
    layer3_outputs(2873) <= not b or a;
    layer3_outputs(2874) <= a and not b;
    layer3_outputs(2875) <= not (a or b);
    layer3_outputs(2876) <= not b or a;
    layer3_outputs(2877) <= b and not a;
    layer3_outputs(2878) <= not b;
    layer3_outputs(2879) <= not (a and b);
    layer3_outputs(2880) <= b;
    layer3_outputs(2881) <= not (a and b);
    layer3_outputs(2882) <= not a;
    layer3_outputs(2883) <= not (a or b);
    layer3_outputs(2884) <= b and not a;
    layer3_outputs(2885) <= not (a and b);
    layer3_outputs(2886) <= not b or a;
    layer3_outputs(2887) <= not b;
    layer3_outputs(2888) <= a or b;
    layer3_outputs(2889) <= not (a or b);
    layer3_outputs(2890) <= not (a xor b);
    layer3_outputs(2891) <= b and not a;
    layer3_outputs(2892) <= a;
    layer3_outputs(2893) <= not (a and b);
    layer3_outputs(2894) <= not (a or b);
    layer3_outputs(2895) <= not (a or b);
    layer3_outputs(2896) <= not b or a;
    layer3_outputs(2897) <= b;
    layer3_outputs(2898) <= b and not a;
    layer3_outputs(2899) <= not b;
    layer3_outputs(2900) <= '0';
    layer3_outputs(2901) <= not (a xor b);
    layer3_outputs(2902) <= not b;
    layer3_outputs(2903) <= '0';
    layer3_outputs(2904) <= a and b;
    layer3_outputs(2905) <= not b;
    layer3_outputs(2906) <= a and not b;
    layer3_outputs(2907) <= b;
    layer3_outputs(2908) <= b and not a;
    layer3_outputs(2909) <= b and not a;
    layer3_outputs(2910) <= not a;
    layer3_outputs(2911) <= not a;
    layer3_outputs(2912) <= not b;
    layer3_outputs(2913) <= a and b;
    layer3_outputs(2914) <= a and not b;
    layer3_outputs(2915) <= '0';
    layer3_outputs(2916) <= not a;
    layer3_outputs(2917) <= not (a or b);
    layer3_outputs(2918) <= not b;
    layer3_outputs(2919) <= not (a or b);
    layer3_outputs(2920) <= b;
    layer3_outputs(2921) <= b;
    layer3_outputs(2922) <= '0';
    layer3_outputs(2923) <= a;
    layer3_outputs(2924) <= '0';
    layer3_outputs(2925) <= a;
    layer3_outputs(2926) <= not b;
    layer3_outputs(2927) <= a and not b;
    layer3_outputs(2928) <= '0';
    layer3_outputs(2929) <= '0';
    layer3_outputs(2930) <= a or b;
    layer3_outputs(2931) <= b;
    layer3_outputs(2932) <= b;
    layer3_outputs(2933) <= a;
    layer3_outputs(2934) <= not (a or b);
    layer3_outputs(2935) <= not (a xor b);
    layer3_outputs(2936) <= a and b;
    layer3_outputs(2937) <= b and not a;
    layer3_outputs(2938) <= not b or a;
    layer3_outputs(2939) <= not b;
    layer3_outputs(2940) <= a;
    layer3_outputs(2941) <= a;
    layer3_outputs(2942) <= not a or b;
    layer3_outputs(2943) <= not a;
    layer3_outputs(2944) <= a;
    layer3_outputs(2945) <= not b;
    layer3_outputs(2946) <= not (a and b);
    layer3_outputs(2947) <= not a;
    layer3_outputs(2948) <= a xor b;
    layer3_outputs(2949) <= not a;
    layer3_outputs(2950) <= not (a and b);
    layer3_outputs(2951) <= not (a and b);
    layer3_outputs(2952) <= not b;
    layer3_outputs(2953) <= '1';
    layer3_outputs(2954) <= a xor b;
    layer3_outputs(2955) <= a;
    layer3_outputs(2956) <= b;
    layer3_outputs(2957) <= b and not a;
    layer3_outputs(2958) <= not a or b;
    layer3_outputs(2959) <= a;
    layer3_outputs(2960) <= not b;
    layer3_outputs(2961) <= '1';
    layer3_outputs(2962) <= a;
    layer3_outputs(2963) <= b;
    layer3_outputs(2964) <= b;
    layer3_outputs(2965) <= a and b;
    layer3_outputs(2966) <= not a;
    layer3_outputs(2967) <= a and not b;
    layer3_outputs(2968) <= a or b;
    layer3_outputs(2969) <= a;
    layer3_outputs(2970) <= b;
    layer3_outputs(2971) <= a;
    layer3_outputs(2972) <= a xor b;
    layer3_outputs(2973) <= '1';
    layer3_outputs(2974) <= a xor b;
    layer3_outputs(2975) <= a and not b;
    layer3_outputs(2976) <= a or b;
    layer3_outputs(2977) <= not b;
    layer3_outputs(2978) <= not b;
    layer3_outputs(2979) <= a or b;
    layer3_outputs(2980) <= a;
    layer3_outputs(2981) <= b;
    layer3_outputs(2982) <= not b;
    layer3_outputs(2983) <= a and b;
    layer3_outputs(2984) <= not a or b;
    layer3_outputs(2985) <= not (a and b);
    layer3_outputs(2986) <= not a;
    layer3_outputs(2987) <= not b or a;
    layer3_outputs(2988) <= not a or b;
    layer3_outputs(2989) <= a or b;
    layer3_outputs(2990) <= a xor b;
    layer3_outputs(2991) <= not (a and b);
    layer3_outputs(2992) <= not b;
    layer3_outputs(2993) <= a;
    layer3_outputs(2994) <= a;
    layer3_outputs(2995) <= b;
    layer3_outputs(2996) <= a;
    layer3_outputs(2997) <= a;
    layer3_outputs(2998) <= not a;
    layer3_outputs(2999) <= not (a and b);
    layer3_outputs(3000) <= not (a xor b);
    layer3_outputs(3001) <= not b or a;
    layer3_outputs(3002) <= not b;
    layer3_outputs(3003) <= a;
    layer3_outputs(3004) <= not (a xor b);
    layer3_outputs(3005) <= not a or b;
    layer3_outputs(3006) <= a and not b;
    layer3_outputs(3007) <= not a;
    layer3_outputs(3008) <= not (a and b);
    layer3_outputs(3009) <= a;
    layer3_outputs(3010) <= not a;
    layer3_outputs(3011) <= b;
    layer3_outputs(3012) <= a;
    layer3_outputs(3013) <= a or b;
    layer3_outputs(3014) <= not a;
    layer3_outputs(3015) <= '1';
    layer3_outputs(3016) <= a and b;
    layer3_outputs(3017) <= b;
    layer3_outputs(3018) <= b;
    layer3_outputs(3019) <= not (a and b);
    layer3_outputs(3020) <= b and not a;
    layer3_outputs(3021) <= not (a and b);
    layer3_outputs(3022) <= a xor b;
    layer3_outputs(3023) <= b;
    layer3_outputs(3024) <= not b;
    layer3_outputs(3025) <= not (a and b);
    layer3_outputs(3026) <= a or b;
    layer3_outputs(3027) <= a xor b;
    layer3_outputs(3028) <= not a or b;
    layer3_outputs(3029) <= not (a and b);
    layer3_outputs(3030) <= not a;
    layer3_outputs(3031) <= a and not b;
    layer3_outputs(3032) <= not a;
    layer3_outputs(3033) <= not (a or b);
    layer3_outputs(3034) <= not a;
    layer3_outputs(3035) <= not b;
    layer3_outputs(3036) <= a xor b;
    layer3_outputs(3037) <= not b;
    layer3_outputs(3038) <= a and b;
    layer3_outputs(3039) <= not a;
    layer3_outputs(3040) <= a;
    layer3_outputs(3041) <= a;
    layer3_outputs(3042) <= a or b;
    layer3_outputs(3043) <= not a;
    layer3_outputs(3044) <= '0';
    layer3_outputs(3045) <= not b;
    layer3_outputs(3046) <= b and not a;
    layer3_outputs(3047) <= a or b;
    layer3_outputs(3048) <= '0';
    layer3_outputs(3049) <= a;
    layer3_outputs(3050) <= a;
    layer3_outputs(3051) <= not a or b;
    layer3_outputs(3052) <= not b;
    layer3_outputs(3053) <= not a or b;
    layer3_outputs(3054) <= a or b;
    layer3_outputs(3055) <= b and not a;
    layer3_outputs(3056) <= not a;
    layer3_outputs(3057) <= a;
    layer3_outputs(3058) <= b;
    layer3_outputs(3059) <= '0';
    layer3_outputs(3060) <= b and not a;
    layer3_outputs(3061) <= a and b;
    layer3_outputs(3062) <= not (a and b);
    layer3_outputs(3063) <= b;
    layer3_outputs(3064) <= not b or a;
    layer3_outputs(3065) <= not (a xor b);
    layer3_outputs(3066) <= not b or a;
    layer3_outputs(3067) <= a;
    layer3_outputs(3068) <= not a;
    layer3_outputs(3069) <= not a or b;
    layer3_outputs(3070) <= a;
    layer3_outputs(3071) <= not b;
    layer3_outputs(3072) <= a and b;
    layer3_outputs(3073) <= a and not b;
    layer3_outputs(3074) <= a and b;
    layer3_outputs(3075) <= not b;
    layer3_outputs(3076) <= not (a xor b);
    layer3_outputs(3077) <= not (a or b);
    layer3_outputs(3078) <= not b;
    layer3_outputs(3079) <= b;
    layer3_outputs(3080) <= a or b;
    layer3_outputs(3081) <= b;
    layer3_outputs(3082) <= b;
    layer3_outputs(3083) <= not a or b;
    layer3_outputs(3084) <= '0';
    layer3_outputs(3085) <= '0';
    layer3_outputs(3086) <= not (a or b);
    layer3_outputs(3087) <= not (a xor b);
    layer3_outputs(3088) <= b;
    layer3_outputs(3089) <= b and not a;
    layer3_outputs(3090) <= not a;
    layer3_outputs(3091) <= a xor b;
    layer3_outputs(3092) <= not (a or b);
    layer3_outputs(3093) <= not (a and b);
    layer3_outputs(3094) <= a and not b;
    layer3_outputs(3095) <= a and b;
    layer3_outputs(3096) <= b;
    layer3_outputs(3097) <= a or b;
    layer3_outputs(3098) <= a;
    layer3_outputs(3099) <= not b;
    layer3_outputs(3100) <= b;
    layer3_outputs(3101) <= not (a and b);
    layer3_outputs(3102) <= a and b;
    layer3_outputs(3103) <= not (a xor b);
    layer3_outputs(3104) <= a or b;
    layer3_outputs(3105) <= not (a xor b);
    layer3_outputs(3106) <= a or b;
    layer3_outputs(3107) <= a;
    layer3_outputs(3108) <= '0';
    layer3_outputs(3109) <= a;
    layer3_outputs(3110) <= '0';
    layer3_outputs(3111) <= a;
    layer3_outputs(3112) <= b and not a;
    layer3_outputs(3113) <= not (a and b);
    layer3_outputs(3114) <= not a;
    layer3_outputs(3115) <= not a or b;
    layer3_outputs(3116) <= a or b;
    layer3_outputs(3117) <= not b;
    layer3_outputs(3118) <= not b or a;
    layer3_outputs(3119) <= '1';
    layer3_outputs(3120) <= not (a and b);
    layer3_outputs(3121) <= not b or a;
    layer3_outputs(3122) <= not (a or b);
    layer3_outputs(3123) <= a;
    layer3_outputs(3124) <= not a;
    layer3_outputs(3125) <= not a;
    layer3_outputs(3126) <= not a or b;
    layer3_outputs(3127) <= '0';
    layer3_outputs(3128) <= '0';
    layer3_outputs(3129) <= a or b;
    layer3_outputs(3130) <= a;
    layer3_outputs(3131) <= b and not a;
    layer3_outputs(3132) <= b and not a;
    layer3_outputs(3133) <= '0';
    layer3_outputs(3134) <= not (a and b);
    layer3_outputs(3135) <= a xor b;
    layer3_outputs(3136) <= not (a or b);
    layer3_outputs(3137) <= not a or b;
    layer3_outputs(3138) <= not (a xor b);
    layer3_outputs(3139) <= '0';
    layer3_outputs(3140) <= not (a and b);
    layer3_outputs(3141) <= a and b;
    layer3_outputs(3142) <= b and not a;
    layer3_outputs(3143) <= not (a xor b);
    layer3_outputs(3144) <= not b or a;
    layer3_outputs(3145) <= b;
    layer3_outputs(3146) <= not (a and b);
    layer3_outputs(3147) <= not b;
    layer3_outputs(3148) <= a;
    layer3_outputs(3149) <= not (a and b);
    layer3_outputs(3150) <= a and not b;
    layer3_outputs(3151) <= not b or a;
    layer3_outputs(3152) <= a and not b;
    layer3_outputs(3153) <= a xor b;
    layer3_outputs(3154) <= not a or b;
    layer3_outputs(3155) <= a;
    layer3_outputs(3156) <= not (a or b);
    layer3_outputs(3157) <= not a or b;
    layer3_outputs(3158) <= not b;
    layer3_outputs(3159) <= not (a and b);
    layer3_outputs(3160) <= a or b;
    layer3_outputs(3161) <= not b;
    layer3_outputs(3162) <= not (a and b);
    layer3_outputs(3163) <= not a;
    layer3_outputs(3164) <= not (a xor b);
    layer3_outputs(3165) <= not (a and b);
    layer3_outputs(3166) <= not b;
    layer3_outputs(3167) <= a or b;
    layer3_outputs(3168) <= '0';
    layer3_outputs(3169) <= b and not a;
    layer3_outputs(3170) <= not b or a;
    layer3_outputs(3171) <= b;
    layer3_outputs(3172) <= a or b;
    layer3_outputs(3173) <= a or b;
    layer3_outputs(3174) <= a and b;
    layer3_outputs(3175) <= not (a and b);
    layer3_outputs(3176) <= a and b;
    layer3_outputs(3177) <= a xor b;
    layer3_outputs(3178) <= b;
    layer3_outputs(3179) <= b and not a;
    layer3_outputs(3180) <= '0';
    layer3_outputs(3181) <= a;
    layer3_outputs(3182) <= not b;
    layer3_outputs(3183) <= a or b;
    layer3_outputs(3184) <= not (a xor b);
    layer3_outputs(3185) <= a;
    layer3_outputs(3186) <= b;
    layer3_outputs(3187) <= a and not b;
    layer3_outputs(3188) <= a xor b;
    layer3_outputs(3189) <= not a;
    layer3_outputs(3190) <= a and b;
    layer3_outputs(3191) <= a or b;
    layer3_outputs(3192) <= not a or b;
    layer3_outputs(3193) <= a and not b;
    layer3_outputs(3194) <= not (a and b);
    layer3_outputs(3195) <= a or b;
    layer3_outputs(3196) <= a and not b;
    layer3_outputs(3197) <= '1';
    layer3_outputs(3198) <= a and not b;
    layer3_outputs(3199) <= not b;
    layer3_outputs(3200) <= a;
    layer3_outputs(3201) <= not b;
    layer3_outputs(3202) <= not a;
    layer3_outputs(3203) <= '1';
    layer3_outputs(3204) <= a and b;
    layer3_outputs(3205) <= a;
    layer3_outputs(3206) <= '0';
    layer3_outputs(3207) <= b;
    layer3_outputs(3208) <= a xor b;
    layer3_outputs(3209) <= a;
    layer3_outputs(3210) <= not b;
    layer3_outputs(3211) <= b;
    layer3_outputs(3212) <= '0';
    layer3_outputs(3213) <= not a;
    layer3_outputs(3214) <= not a;
    layer3_outputs(3215) <= not (a xor b);
    layer3_outputs(3216) <= not a;
    layer3_outputs(3217) <= a and b;
    layer3_outputs(3218) <= not b or a;
    layer3_outputs(3219) <= not (a xor b);
    layer3_outputs(3220) <= '1';
    layer3_outputs(3221) <= not b;
    layer3_outputs(3222) <= a and not b;
    layer3_outputs(3223) <= b;
    layer3_outputs(3224) <= not a;
    layer3_outputs(3225) <= a and b;
    layer3_outputs(3226) <= not (a or b);
    layer3_outputs(3227) <= not (a or b);
    layer3_outputs(3228) <= not a or b;
    layer3_outputs(3229) <= '0';
    layer3_outputs(3230) <= not (a xor b);
    layer3_outputs(3231) <= a and b;
    layer3_outputs(3232) <= b;
    layer3_outputs(3233) <= '1';
    layer3_outputs(3234) <= a and not b;
    layer3_outputs(3235) <= a;
    layer3_outputs(3236) <= not b;
    layer3_outputs(3237) <= b;
    layer3_outputs(3238) <= a and not b;
    layer3_outputs(3239) <= not a;
    layer3_outputs(3240) <= not b;
    layer3_outputs(3241) <= a;
    layer3_outputs(3242) <= a or b;
    layer3_outputs(3243) <= a;
    layer3_outputs(3244) <= not a or b;
    layer3_outputs(3245) <= not a;
    layer3_outputs(3246) <= a and b;
    layer3_outputs(3247) <= not b;
    layer3_outputs(3248) <= not b or a;
    layer3_outputs(3249) <= not b;
    layer3_outputs(3250) <= not a;
    layer3_outputs(3251) <= a;
    layer3_outputs(3252) <= not (a xor b);
    layer3_outputs(3253) <= not b;
    layer3_outputs(3254) <= not b or a;
    layer3_outputs(3255) <= b and not a;
    layer3_outputs(3256) <= not (a and b);
    layer3_outputs(3257) <= a and not b;
    layer3_outputs(3258) <= a;
    layer3_outputs(3259) <= b;
    layer3_outputs(3260) <= not (a and b);
    layer3_outputs(3261) <= a and not b;
    layer3_outputs(3262) <= a;
    layer3_outputs(3263) <= not b or a;
    layer3_outputs(3264) <= a;
    layer3_outputs(3265) <= '1';
    layer3_outputs(3266) <= not (a or b);
    layer3_outputs(3267) <= not a;
    layer3_outputs(3268) <= a and b;
    layer3_outputs(3269) <= b and not a;
    layer3_outputs(3270) <= b and not a;
    layer3_outputs(3271) <= a and b;
    layer3_outputs(3272) <= '1';
    layer3_outputs(3273) <= not a;
    layer3_outputs(3274) <= a and b;
    layer3_outputs(3275) <= b;
    layer3_outputs(3276) <= '0';
    layer3_outputs(3277) <= a;
    layer3_outputs(3278) <= not a;
    layer3_outputs(3279) <= not a;
    layer3_outputs(3280) <= a;
    layer3_outputs(3281) <= not b or a;
    layer3_outputs(3282) <= not (a or b);
    layer3_outputs(3283) <= a or b;
    layer3_outputs(3284) <= a and b;
    layer3_outputs(3285) <= b;
    layer3_outputs(3286) <= not b or a;
    layer3_outputs(3287) <= not (a xor b);
    layer3_outputs(3288) <= not a or b;
    layer3_outputs(3289) <= a or b;
    layer3_outputs(3290) <= a;
    layer3_outputs(3291) <= b;
    layer3_outputs(3292) <= not (a or b);
    layer3_outputs(3293) <= a and not b;
    layer3_outputs(3294) <= a or b;
    layer3_outputs(3295) <= a and b;
    layer3_outputs(3296) <= not b;
    layer3_outputs(3297) <= not b;
    layer3_outputs(3298) <= a;
    layer3_outputs(3299) <= b;
    layer3_outputs(3300) <= not (a and b);
    layer3_outputs(3301) <= not b;
    layer3_outputs(3302) <= not a;
    layer3_outputs(3303) <= a;
    layer3_outputs(3304) <= '0';
    layer3_outputs(3305) <= a;
    layer3_outputs(3306) <= a and b;
    layer3_outputs(3307) <= not a;
    layer3_outputs(3308) <= a and b;
    layer3_outputs(3309) <= not (a and b);
    layer3_outputs(3310) <= b;
    layer3_outputs(3311) <= a and not b;
    layer3_outputs(3312) <= not b;
    layer3_outputs(3313) <= a xor b;
    layer3_outputs(3314) <= b and not a;
    layer3_outputs(3315) <= not a;
    layer3_outputs(3316) <= b and not a;
    layer3_outputs(3317) <= '1';
    layer3_outputs(3318) <= not a;
    layer3_outputs(3319) <= not a;
    layer3_outputs(3320) <= b;
    layer3_outputs(3321) <= b and not a;
    layer3_outputs(3322) <= not (a or b);
    layer3_outputs(3323) <= b;
    layer3_outputs(3324) <= a;
    layer3_outputs(3325) <= a;
    layer3_outputs(3326) <= a or b;
    layer3_outputs(3327) <= b and not a;
    layer3_outputs(3328) <= b and not a;
    layer3_outputs(3329) <= a xor b;
    layer3_outputs(3330) <= a or b;
    layer3_outputs(3331) <= not a;
    layer3_outputs(3332) <= b;
    layer3_outputs(3333) <= not b or a;
    layer3_outputs(3334) <= a and not b;
    layer3_outputs(3335) <= not a;
    layer3_outputs(3336) <= '0';
    layer3_outputs(3337) <= b;
    layer3_outputs(3338) <= a;
    layer3_outputs(3339) <= b;
    layer3_outputs(3340) <= not b;
    layer3_outputs(3341) <= not b;
    layer3_outputs(3342) <= '1';
    layer3_outputs(3343) <= not a;
    layer3_outputs(3344) <= '0';
    layer3_outputs(3345) <= not b;
    layer3_outputs(3346) <= not b or a;
    layer3_outputs(3347) <= a or b;
    layer3_outputs(3348) <= not a;
    layer3_outputs(3349) <= not a;
    layer3_outputs(3350) <= b and not a;
    layer3_outputs(3351) <= not b;
    layer3_outputs(3352) <= a or b;
    layer3_outputs(3353) <= not (a or b);
    layer3_outputs(3354) <= a;
    layer3_outputs(3355) <= not b;
    layer3_outputs(3356) <= not a;
    layer3_outputs(3357) <= not a or b;
    layer3_outputs(3358) <= not b or a;
    layer3_outputs(3359) <= b and not a;
    layer3_outputs(3360) <= not a;
    layer3_outputs(3361) <= a or b;
    layer3_outputs(3362) <= not a;
    layer3_outputs(3363) <= not b;
    layer3_outputs(3364) <= not a or b;
    layer3_outputs(3365) <= b;
    layer3_outputs(3366) <= a and b;
    layer3_outputs(3367) <= b and not a;
    layer3_outputs(3368) <= a;
    layer3_outputs(3369) <= not a or b;
    layer3_outputs(3370) <= a xor b;
    layer3_outputs(3371) <= b and not a;
    layer3_outputs(3372) <= a;
    layer3_outputs(3373) <= not (a and b);
    layer3_outputs(3374) <= not (a and b);
    layer3_outputs(3375) <= not b;
    layer3_outputs(3376) <= not a or b;
    layer3_outputs(3377) <= '1';
    layer3_outputs(3378) <= not a;
    layer3_outputs(3379) <= not (a and b);
    layer3_outputs(3380) <= not b or a;
    layer3_outputs(3381) <= '1';
    layer3_outputs(3382) <= b and not a;
    layer3_outputs(3383) <= b and not a;
    layer3_outputs(3384) <= b;
    layer3_outputs(3385) <= b;
    layer3_outputs(3386) <= '1';
    layer3_outputs(3387) <= not a;
    layer3_outputs(3388) <= not b or a;
    layer3_outputs(3389) <= b;
    layer3_outputs(3390) <= b;
    layer3_outputs(3391) <= '1';
    layer3_outputs(3392) <= '0';
    layer3_outputs(3393) <= a or b;
    layer3_outputs(3394) <= b;
    layer3_outputs(3395) <= a;
    layer3_outputs(3396) <= a;
    layer3_outputs(3397) <= not (a or b);
    layer3_outputs(3398) <= not (a xor b);
    layer3_outputs(3399) <= not a or b;
    layer3_outputs(3400) <= not (a or b);
    layer3_outputs(3401) <= a;
    layer3_outputs(3402) <= a or b;
    layer3_outputs(3403) <= not b or a;
    layer3_outputs(3404) <= not (a and b);
    layer3_outputs(3405) <= not b;
    layer3_outputs(3406) <= b and not a;
    layer3_outputs(3407) <= not b;
    layer3_outputs(3408) <= b and not a;
    layer3_outputs(3409) <= a;
    layer3_outputs(3410) <= a;
    layer3_outputs(3411) <= '1';
    layer3_outputs(3412) <= a;
    layer3_outputs(3413) <= b;
    layer3_outputs(3414) <= a;
    layer3_outputs(3415) <= not b;
    layer3_outputs(3416) <= a and not b;
    layer3_outputs(3417) <= a;
    layer3_outputs(3418) <= a xor b;
    layer3_outputs(3419) <= a or b;
    layer3_outputs(3420) <= not b;
    layer3_outputs(3421) <= not (a xor b);
    layer3_outputs(3422) <= '1';
    layer3_outputs(3423) <= not (a xor b);
    layer3_outputs(3424) <= not a;
    layer3_outputs(3425) <= not (a and b);
    layer3_outputs(3426) <= a and not b;
    layer3_outputs(3427) <= '1';
    layer3_outputs(3428) <= a or b;
    layer3_outputs(3429) <= not a;
    layer3_outputs(3430) <= not b or a;
    layer3_outputs(3431) <= a;
    layer3_outputs(3432) <= '0';
    layer3_outputs(3433) <= not (a xor b);
    layer3_outputs(3434) <= not b;
    layer3_outputs(3435) <= not (a and b);
    layer3_outputs(3436) <= a and not b;
    layer3_outputs(3437) <= a;
    layer3_outputs(3438) <= not a or b;
    layer3_outputs(3439) <= not a;
    layer3_outputs(3440) <= not b;
    layer3_outputs(3441) <= a xor b;
    layer3_outputs(3442) <= not b;
    layer3_outputs(3443) <= '0';
    layer3_outputs(3444) <= a or b;
    layer3_outputs(3445) <= '1';
    layer3_outputs(3446) <= '1';
    layer3_outputs(3447) <= b;
    layer3_outputs(3448) <= '1';
    layer3_outputs(3449) <= a;
    layer3_outputs(3450) <= not b or a;
    layer3_outputs(3451) <= a and b;
    layer3_outputs(3452) <= not a;
    layer3_outputs(3453) <= '0';
    layer3_outputs(3454) <= not a;
    layer3_outputs(3455) <= a and not b;
    layer3_outputs(3456) <= not a;
    layer3_outputs(3457) <= not b;
    layer3_outputs(3458) <= b and not a;
    layer3_outputs(3459) <= not a;
    layer3_outputs(3460) <= not a or b;
    layer3_outputs(3461) <= not a;
    layer3_outputs(3462) <= not (a xor b);
    layer3_outputs(3463) <= a;
    layer3_outputs(3464) <= b and not a;
    layer3_outputs(3465) <= '0';
    layer3_outputs(3466) <= '1';
    layer3_outputs(3467) <= not b or a;
    layer3_outputs(3468) <= not a or b;
    layer3_outputs(3469) <= not b;
    layer3_outputs(3470) <= b and not a;
    layer3_outputs(3471) <= not b;
    layer3_outputs(3472) <= a;
    layer3_outputs(3473) <= a;
    layer3_outputs(3474) <= not b or a;
    layer3_outputs(3475) <= a;
    layer3_outputs(3476) <= not b;
    layer3_outputs(3477) <= '1';
    layer3_outputs(3478) <= b;
    layer3_outputs(3479) <= b;
    layer3_outputs(3480) <= not (a or b);
    layer3_outputs(3481) <= b;
    layer3_outputs(3482) <= a xor b;
    layer3_outputs(3483) <= a and not b;
    layer3_outputs(3484) <= b;
    layer3_outputs(3485) <= not b or a;
    layer3_outputs(3486) <= b;
    layer3_outputs(3487) <= not a;
    layer3_outputs(3488) <= not b or a;
    layer3_outputs(3489) <= a and b;
    layer3_outputs(3490) <= not a;
    layer3_outputs(3491) <= a or b;
    layer3_outputs(3492) <= a and not b;
    layer3_outputs(3493) <= not (a xor b);
    layer3_outputs(3494) <= a and not b;
    layer3_outputs(3495) <= not (a or b);
    layer3_outputs(3496) <= not a or b;
    layer3_outputs(3497) <= not (a xor b);
    layer3_outputs(3498) <= not a;
    layer3_outputs(3499) <= not b or a;
    layer3_outputs(3500) <= not b;
    layer3_outputs(3501) <= b;
    layer3_outputs(3502) <= not (a xor b);
    layer3_outputs(3503) <= not (a and b);
    layer3_outputs(3504) <= not b;
    layer3_outputs(3505) <= a;
    layer3_outputs(3506) <= a and b;
    layer3_outputs(3507) <= not b or a;
    layer3_outputs(3508) <= a or b;
    layer3_outputs(3509) <= a and b;
    layer3_outputs(3510) <= not (a or b);
    layer3_outputs(3511) <= a;
    layer3_outputs(3512) <= not a or b;
    layer3_outputs(3513) <= a and b;
    layer3_outputs(3514) <= not (a or b);
    layer3_outputs(3515) <= not (a or b);
    layer3_outputs(3516) <= not (a xor b);
    layer3_outputs(3517) <= not (a and b);
    layer3_outputs(3518) <= not (a and b);
    layer3_outputs(3519) <= a and b;
    layer3_outputs(3520) <= a and not b;
    layer3_outputs(3521) <= not b or a;
    layer3_outputs(3522) <= not a;
    layer3_outputs(3523) <= a and not b;
    layer3_outputs(3524) <= b;
    layer3_outputs(3525) <= not a;
    layer3_outputs(3526) <= not (a or b);
    layer3_outputs(3527) <= not (a and b);
    layer3_outputs(3528) <= not b;
    layer3_outputs(3529) <= not a;
    layer3_outputs(3530) <= a;
    layer3_outputs(3531) <= not b;
    layer3_outputs(3532) <= not a or b;
    layer3_outputs(3533) <= not a;
    layer3_outputs(3534) <= not (a or b);
    layer3_outputs(3535) <= a and not b;
    layer3_outputs(3536) <= a or b;
    layer3_outputs(3537) <= a;
    layer3_outputs(3538) <= not a or b;
    layer3_outputs(3539) <= not b;
    layer3_outputs(3540) <= b and not a;
    layer3_outputs(3541) <= b and not a;
    layer3_outputs(3542) <= a and not b;
    layer3_outputs(3543) <= not b;
    layer3_outputs(3544) <= a;
    layer3_outputs(3545) <= a or b;
    layer3_outputs(3546) <= b;
    layer3_outputs(3547) <= not b;
    layer3_outputs(3548) <= b;
    layer3_outputs(3549) <= not b;
    layer3_outputs(3550) <= a;
    layer3_outputs(3551) <= not a;
    layer3_outputs(3552) <= '0';
    layer3_outputs(3553) <= a;
    layer3_outputs(3554) <= b;
    layer3_outputs(3555) <= not (a and b);
    layer3_outputs(3556) <= not a;
    layer3_outputs(3557) <= not (a or b);
    layer3_outputs(3558) <= not (a and b);
    layer3_outputs(3559) <= a;
    layer3_outputs(3560) <= not a;
    layer3_outputs(3561) <= a xor b;
    layer3_outputs(3562) <= a and b;
    layer3_outputs(3563) <= not a or b;
    layer3_outputs(3564) <= a and b;
    layer3_outputs(3565) <= not (a or b);
    layer3_outputs(3566) <= a and b;
    layer3_outputs(3567) <= not (a or b);
    layer3_outputs(3568) <= a;
    layer3_outputs(3569) <= '0';
    layer3_outputs(3570) <= a or b;
    layer3_outputs(3571) <= a and not b;
    layer3_outputs(3572) <= b and not a;
    layer3_outputs(3573) <= '0';
    layer3_outputs(3574) <= b;
    layer3_outputs(3575) <= not (a or b);
    layer3_outputs(3576) <= '1';
    layer3_outputs(3577) <= b and not a;
    layer3_outputs(3578) <= a xor b;
    layer3_outputs(3579) <= not (a or b);
    layer3_outputs(3580) <= b and not a;
    layer3_outputs(3581) <= b;
    layer3_outputs(3582) <= not (a and b);
    layer3_outputs(3583) <= not (a and b);
    layer3_outputs(3584) <= a;
    layer3_outputs(3585) <= '1';
    layer3_outputs(3586) <= not (a and b);
    layer3_outputs(3587) <= not (a or b);
    layer3_outputs(3588) <= b and not a;
    layer3_outputs(3589) <= not b;
    layer3_outputs(3590) <= b;
    layer3_outputs(3591) <= not (a or b);
    layer3_outputs(3592) <= not b;
    layer3_outputs(3593) <= a and b;
    layer3_outputs(3594) <= a and b;
    layer3_outputs(3595) <= '0';
    layer3_outputs(3596) <= a;
    layer3_outputs(3597) <= not b or a;
    layer3_outputs(3598) <= not (a xor b);
    layer3_outputs(3599) <= not a or b;
    layer3_outputs(3600) <= not a;
    layer3_outputs(3601) <= not a or b;
    layer3_outputs(3602) <= not (a and b);
    layer3_outputs(3603) <= not b;
    layer3_outputs(3604) <= a and not b;
    layer3_outputs(3605) <= a and b;
    layer3_outputs(3606) <= b and not a;
    layer3_outputs(3607) <= a xor b;
    layer3_outputs(3608) <= a;
    layer3_outputs(3609) <= '1';
    layer3_outputs(3610) <= not (a or b);
    layer3_outputs(3611) <= '0';
    layer3_outputs(3612) <= not a or b;
    layer3_outputs(3613) <= not a or b;
    layer3_outputs(3614) <= not a;
    layer3_outputs(3615) <= a or b;
    layer3_outputs(3616) <= not a;
    layer3_outputs(3617) <= '0';
    layer3_outputs(3618) <= not b;
    layer3_outputs(3619) <= a xor b;
    layer3_outputs(3620) <= not a or b;
    layer3_outputs(3621) <= not (a and b);
    layer3_outputs(3622) <= a xor b;
    layer3_outputs(3623) <= '0';
    layer3_outputs(3624) <= '0';
    layer3_outputs(3625) <= not a;
    layer3_outputs(3626) <= not b;
    layer3_outputs(3627) <= b;
    layer3_outputs(3628) <= not b;
    layer3_outputs(3629) <= not b;
    layer3_outputs(3630) <= '0';
    layer3_outputs(3631) <= a and not b;
    layer3_outputs(3632) <= not (a and b);
    layer3_outputs(3633) <= '1';
    layer3_outputs(3634) <= not b;
    layer3_outputs(3635) <= '1';
    layer3_outputs(3636) <= a;
    layer3_outputs(3637) <= not b;
    layer3_outputs(3638) <= a and b;
    layer3_outputs(3639) <= '1';
    layer3_outputs(3640) <= a and not b;
    layer3_outputs(3641) <= a and not b;
    layer3_outputs(3642) <= not b or a;
    layer3_outputs(3643) <= not a;
    layer3_outputs(3644) <= a and not b;
    layer3_outputs(3645) <= b and not a;
    layer3_outputs(3646) <= a and not b;
    layer3_outputs(3647) <= b and not a;
    layer3_outputs(3648) <= not b;
    layer3_outputs(3649) <= a;
    layer3_outputs(3650) <= '1';
    layer3_outputs(3651) <= a and b;
    layer3_outputs(3652) <= a or b;
    layer3_outputs(3653) <= not (a or b);
    layer3_outputs(3654) <= b;
    layer3_outputs(3655) <= not a or b;
    layer3_outputs(3656) <= a and not b;
    layer3_outputs(3657) <= '0';
    layer3_outputs(3658) <= a and b;
    layer3_outputs(3659) <= a;
    layer3_outputs(3660) <= '1';
    layer3_outputs(3661) <= a and b;
    layer3_outputs(3662) <= b and not a;
    layer3_outputs(3663) <= '0';
    layer3_outputs(3664) <= not a;
    layer3_outputs(3665) <= a and not b;
    layer3_outputs(3666) <= a;
    layer3_outputs(3667) <= not (a or b);
    layer3_outputs(3668) <= '0';
    layer3_outputs(3669) <= not (a or b);
    layer3_outputs(3670) <= not a or b;
    layer3_outputs(3671) <= not a;
    layer3_outputs(3672) <= '0';
    layer3_outputs(3673) <= b;
    layer3_outputs(3674) <= not (a xor b);
    layer3_outputs(3675) <= a;
    layer3_outputs(3676) <= not b or a;
    layer3_outputs(3677) <= '0';
    layer3_outputs(3678) <= a and b;
    layer3_outputs(3679) <= not a;
    layer3_outputs(3680) <= b;
    layer3_outputs(3681) <= not b;
    layer3_outputs(3682) <= a or b;
    layer3_outputs(3683) <= not (a and b);
    layer3_outputs(3684) <= not a;
    layer3_outputs(3685) <= not b;
    layer3_outputs(3686) <= not b;
    layer3_outputs(3687) <= a and b;
    layer3_outputs(3688) <= not b;
    layer3_outputs(3689) <= not (a xor b);
    layer3_outputs(3690) <= a;
    layer3_outputs(3691) <= '0';
    layer3_outputs(3692) <= not a or b;
    layer3_outputs(3693) <= not (a or b);
    layer3_outputs(3694) <= not (a xor b);
    layer3_outputs(3695) <= not a;
    layer3_outputs(3696) <= a or b;
    layer3_outputs(3697) <= not a or b;
    layer3_outputs(3698) <= '0';
    layer3_outputs(3699) <= a;
    layer3_outputs(3700) <= not a or b;
    layer3_outputs(3701) <= not b;
    layer3_outputs(3702) <= not b;
    layer3_outputs(3703) <= a;
    layer3_outputs(3704) <= b and not a;
    layer3_outputs(3705) <= not b or a;
    layer3_outputs(3706) <= not b;
    layer3_outputs(3707) <= not a or b;
    layer3_outputs(3708) <= a and not b;
    layer3_outputs(3709) <= a;
    layer3_outputs(3710) <= not a or b;
    layer3_outputs(3711) <= not a;
    layer3_outputs(3712) <= not (a and b);
    layer3_outputs(3713) <= b;
    layer3_outputs(3714) <= b;
    layer3_outputs(3715) <= not (a xor b);
    layer3_outputs(3716) <= a and b;
    layer3_outputs(3717) <= not (a and b);
    layer3_outputs(3718) <= not a;
    layer3_outputs(3719) <= not a;
    layer3_outputs(3720) <= '1';
    layer3_outputs(3721) <= not b;
    layer3_outputs(3722) <= not (a or b);
    layer3_outputs(3723) <= not b or a;
    layer3_outputs(3724) <= a and b;
    layer3_outputs(3725) <= not (a or b);
    layer3_outputs(3726) <= a;
    layer3_outputs(3727) <= a and not b;
    layer3_outputs(3728) <= not a;
    layer3_outputs(3729) <= a;
    layer3_outputs(3730) <= '1';
    layer3_outputs(3731) <= not a;
    layer3_outputs(3732) <= not b;
    layer3_outputs(3733) <= not (a and b);
    layer3_outputs(3734) <= b;
    layer3_outputs(3735) <= a;
    layer3_outputs(3736) <= a;
    layer3_outputs(3737) <= not b;
    layer3_outputs(3738) <= not (a and b);
    layer3_outputs(3739) <= not a or b;
    layer3_outputs(3740) <= not a;
    layer3_outputs(3741) <= '0';
    layer3_outputs(3742) <= b;
    layer3_outputs(3743) <= a xor b;
    layer3_outputs(3744) <= not b;
    layer3_outputs(3745) <= a;
    layer3_outputs(3746) <= not b;
    layer3_outputs(3747) <= a xor b;
    layer3_outputs(3748) <= b;
    layer3_outputs(3749) <= not b;
    layer3_outputs(3750) <= a and not b;
    layer3_outputs(3751) <= not (a or b);
    layer3_outputs(3752) <= not b;
    layer3_outputs(3753) <= not a or b;
    layer3_outputs(3754) <= not (a and b);
    layer3_outputs(3755) <= a xor b;
    layer3_outputs(3756) <= b and not a;
    layer3_outputs(3757) <= '0';
    layer3_outputs(3758) <= '1';
    layer3_outputs(3759) <= b and not a;
    layer3_outputs(3760) <= not a;
    layer3_outputs(3761) <= not (a xor b);
    layer3_outputs(3762) <= '0';
    layer3_outputs(3763) <= not (a xor b);
    layer3_outputs(3764) <= not a;
    layer3_outputs(3765) <= b;
    layer3_outputs(3766) <= a;
    layer3_outputs(3767) <= not b;
    layer3_outputs(3768) <= b;
    layer3_outputs(3769) <= b and not a;
    layer3_outputs(3770) <= a;
    layer3_outputs(3771) <= not a;
    layer3_outputs(3772) <= not a or b;
    layer3_outputs(3773) <= b;
    layer3_outputs(3774) <= not b or a;
    layer3_outputs(3775) <= not (a and b);
    layer3_outputs(3776) <= not a;
    layer3_outputs(3777) <= not (a xor b);
    layer3_outputs(3778) <= a or b;
    layer3_outputs(3779) <= not (a or b);
    layer3_outputs(3780) <= a xor b;
    layer3_outputs(3781) <= b;
    layer3_outputs(3782) <= a and not b;
    layer3_outputs(3783) <= b;
    layer3_outputs(3784) <= not (a or b);
    layer3_outputs(3785) <= not b;
    layer3_outputs(3786) <= a;
    layer3_outputs(3787) <= not b;
    layer3_outputs(3788) <= a or b;
    layer3_outputs(3789) <= not b or a;
    layer3_outputs(3790) <= b and not a;
    layer3_outputs(3791) <= not a or b;
    layer3_outputs(3792) <= not (a and b);
    layer3_outputs(3793) <= not a;
    layer3_outputs(3794) <= '1';
    layer3_outputs(3795) <= not a;
    layer3_outputs(3796) <= b;
    layer3_outputs(3797) <= not a or b;
    layer3_outputs(3798) <= not (a and b);
    layer3_outputs(3799) <= a;
    layer3_outputs(3800) <= not b;
    layer3_outputs(3801) <= b and not a;
    layer3_outputs(3802) <= not a;
    layer3_outputs(3803) <= not a;
    layer3_outputs(3804) <= not b;
    layer3_outputs(3805) <= '0';
    layer3_outputs(3806) <= a;
    layer3_outputs(3807) <= '0';
    layer3_outputs(3808) <= not b;
    layer3_outputs(3809) <= a;
    layer3_outputs(3810) <= not b;
    layer3_outputs(3811) <= a and b;
    layer3_outputs(3812) <= not (a and b);
    layer3_outputs(3813) <= not b;
    layer3_outputs(3814) <= b and not a;
    layer3_outputs(3815) <= a or b;
    layer3_outputs(3816) <= not (a and b);
    layer3_outputs(3817) <= not b;
    layer3_outputs(3818) <= b and not a;
    layer3_outputs(3819) <= a or b;
    layer3_outputs(3820) <= a;
    layer3_outputs(3821) <= not (a or b);
    layer3_outputs(3822) <= not (a xor b);
    layer3_outputs(3823) <= not b or a;
    layer3_outputs(3824) <= a and b;
    layer3_outputs(3825) <= a and b;
    layer3_outputs(3826) <= '0';
    layer3_outputs(3827) <= not (a or b);
    layer3_outputs(3828) <= not a or b;
    layer3_outputs(3829) <= a and b;
    layer3_outputs(3830) <= a and not b;
    layer3_outputs(3831) <= b and not a;
    layer3_outputs(3832) <= a or b;
    layer3_outputs(3833) <= b and not a;
    layer3_outputs(3834) <= not b;
    layer3_outputs(3835) <= not a or b;
    layer3_outputs(3836) <= a and b;
    layer3_outputs(3837) <= b and not a;
    layer3_outputs(3838) <= not b;
    layer3_outputs(3839) <= a xor b;
    layer3_outputs(3840) <= b and not a;
    layer3_outputs(3841) <= a;
    layer3_outputs(3842) <= a or b;
    layer3_outputs(3843) <= a;
    layer3_outputs(3844) <= not a;
    layer3_outputs(3845) <= a and b;
    layer3_outputs(3846) <= a;
    layer3_outputs(3847) <= not a or b;
    layer3_outputs(3848) <= a xor b;
    layer3_outputs(3849) <= not (a or b);
    layer3_outputs(3850) <= b;
    layer3_outputs(3851) <= not (a and b);
    layer3_outputs(3852) <= b and not a;
    layer3_outputs(3853) <= b;
    layer3_outputs(3854) <= a;
    layer3_outputs(3855) <= a;
    layer3_outputs(3856) <= a or b;
    layer3_outputs(3857) <= b and not a;
    layer3_outputs(3858) <= not b or a;
    layer3_outputs(3859) <= not a;
    layer3_outputs(3860) <= not a;
    layer3_outputs(3861) <= b;
    layer3_outputs(3862) <= not b;
    layer3_outputs(3863) <= not b;
    layer3_outputs(3864) <= a;
    layer3_outputs(3865) <= '1';
    layer3_outputs(3866) <= not b;
    layer3_outputs(3867) <= not (a and b);
    layer3_outputs(3868) <= a xor b;
    layer3_outputs(3869) <= not b or a;
    layer3_outputs(3870) <= not a or b;
    layer3_outputs(3871) <= '1';
    layer3_outputs(3872) <= not a or b;
    layer3_outputs(3873) <= b and not a;
    layer3_outputs(3874) <= b;
    layer3_outputs(3875) <= not (a or b);
    layer3_outputs(3876) <= a and b;
    layer3_outputs(3877) <= not (a or b);
    layer3_outputs(3878) <= a or b;
    layer3_outputs(3879) <= a;
    layer3_outputs(3880) <= b;
    layer3_outputs(3881) <= not a;
    layer3_outputs(3882) <= '1';
    layer3_outputs(3883) <= not b;
    layer3_outputs(3884) <= not a or b;
    layer3_outputs(3885) <= a xor b;
    layer3_outputs(3886) <= not (a xor b);
    layer3_outputs(3887) <= '0';
    layer3_outputs(3888) <= not a;
    layer3_outputs(3889) <= not (a xor b);
    layer3_outputs(3890) <= b;
    layer3_outputs(3891) <= b and not a;
    layer3_outputs(3892) <= not a or b;
    layer3_outputs(3893) <= b;
    layer3_outputs(3894) <= '1';
    layer3_outputs(3895) <= a or b;
    layer3_outputs(3896) <= a;
    layer3_outputs(3897) <= a and b;
    layer3_outputs(3898) <= not a;
    layer3_outputs(3899) <= not (a and b);
    layer3_outputs(3900) <= not b;
    layer3_outputs(3901) <= '1';
    layer3_outputs(3902) <= not b or a;
    layer3_outputs(3903) <= a and not b;
    layer3_outputs(3904) <= '0';
    layer3_outputs(3905) <= a or b;
    layer3_outputs(3906) <= '0';
    layer3_outputs(3907) <= not (a and b);
    layer3_outputs(3908) <= not (a or b);
    layer3_outputs(3909) <= a or b;
    layer3_outputs(3910) <= not (a xor b);
    layer3_outputs(3911) <= '1';
    layer3_outputs(3912) <= a and not b;
    layer3_outputs(3913) <= not b or a;
    layer3_outputs(3914) <= '1';
    layer3_outputs(3915) <= not a or b;
    layer3_outputs(3916) <= not a;
    layer3_outputs(3917) <= b and not a;
    layer3_outputs(3918) <= not a or b;
    layer3_outputs(3919) <= not a;
    layer3_outputs(3920) <= '1';
    layer3_outputs(3921) <= not a;
    layer3_outputs(3922) <= a and not b;
    layer3_outputs(3923) <= b;
    layer3_outputs(3924) <= a;
    layer3_outputs(3925) <= not (a or b);
    layer3_outputs(3926) <= b;
    layer3_outputs(3927) <= not b;
    layer3_outputs(3928) <= a and b;
    layer3_outputs(3929) <= a or b;
    layer3_outputs(3930) <= '0';
    layer3_outputs(3931) <= not b;
    layer3_outputs(3932) <= not a or b;
    layer3_outputs(3933) <= not a;
    layer3_outputs(3934) <= a or b;
    layer3_outputs(3935) <= not (a and b);
    layer3_outputs(3936) <= a and not b;
    layer3_outputs(3937) <= a xor b;
    layer3_outputs(3938) <= b;
    layer3_outputs(3939) <= '1';
    layer3_outputs(3940) <= not (a and b);
    layer3_outputs(3941) <= a and b;
    layer3_outputs(3942) <= a or b;
    layer3_outputs(3943) <= not a;
    layer3_outputs(3944) <= b;
    layer3_outputs(3945) <= not b;
    layer3_outputs(3946) <= not (a or b);
    layer3_outputs(3947) <= not a;
    layer3_outputs(3948) <= not a or b;
    layer3_outputs(3949) <= a;
    layer3_outputs(3950) <= not b or a;
    layer3_outputs(3951) <= not (a or b);
    layer3_outputs(3952) <= not a;
    layer3_outputs(3953) <= b;
    layer3_outputs(3954) <= b;
    layer3_outputs(3955) <= not (a or b);
    layer3_outputs(3956) <= '0';
    layer3_outputs(3957) <= b;
    layer3_outputs(3958) <= not (a and b);
    layer3_outputs(3959) <= a or b;
    layer3_outputs(3960) <= not (a or b);
    layer3_outputs(3961) <= a and not b;
    layer3_outputs(3962) <= '1';
    layer3_outputs(3963) <= a xor b;
    layer3_outputs(3964) <= '1';
    layer3_outputs(3965) <= not (a and b);
    layer3_outputs(3966) <= '0';
    layer3_outputs(3967) <= not b or a;
    layer3_outputs(3968) <= '0';
    layer3_outputs(3969) <= not b or a;
    layer3_outputs(3970) <= not (a xor b);
    layer3_outputs(3971) <= b;
    layer3_outputs(3972) <= a;
    layer3_outputs(3973) <= b;
    layer3_outputs(3974) <= not (a and b);
    layer3_outputs(3975) <= not a;
    layer3_outputs(3976) <= not (a or b);
    layer3_outputs(3977) <= a and not b;
    layer3_outputs(3978) <= '1';
    layer3_outputs(3979) <= b;
    layer3_outputs(3980) <= not b or a;
    layer3_outputs(3981) <= a and b;
    layer3_outputs(3982) <= not (a xor b);
    layer3_outputs(3983) <= b;
    layer3_outputs(3984) <= a or b;
    layer3_outputs(3985) <= a;
    layer3_outputs(3986) <= not a;
    layer3_outputs(3987) <= b;
    layer3_outputs(3988) <= not (a xor b);
    layer3_outputs(3989) <= not a;
    layer3_outputs(3990) <= '1';
    layer3_outputs(3991) <= a;
    layer3_outputs(3992) <= not a;
    layer3_outputs(3993) <= not b;
    layer3_outputs(3994) <= not (a xor b);
    layer3_outputs(3995) <= not b or a;
    layer3_outputs(3996) <= a xor b;
    layer3_outputs(3997) <= not (a and b);
    layer3_outputs(3998) <= a and b;
    layer3_outputs(3999) <= a xor b;
    layer3_outputs(4000) <= a xor b;
    layer3_outputs(4001) <= a or b;
    layer3_outputs(4002) <= b and not a;
    layer3_outputs(4003) <= a and b;
    layer3_outputs(4004) <= b;
    layer3_outputs(4005) <= b and not a;
    layer3_outputs(4006) <= not a;
    layer3_outputs(4007) <= a xor b;
    layer3_outputs(4008) <= a xor b;
    layer3_outputs(4009) <= not a or b;
    layer3_outputs(4010) <= not b;
    layer3_outputs(4011) <= a;
    layer3_outputs(4012) <= b;
    layer3_outputs(4013) <= b;
    layer3_outputs(4014) <= not (a or b);
    layer3_outputs(4015) <= a or b;
    layer3_outputs(4016) <= not (a and b);
    layer3_outputs(4017) <= b;
    layer3_outputs(4018) <= not b or a;
    layer3_outputs(4019) <= not a or b;
    layer3_outputs(4020) <= not a or b;
    layer3_outputs(4021) <= b;
    layer3_outputs(4022) <= b and not a;
    layer3_outputs(4023) <= not (a or b);
    layer3_outputs(4024) <= a and b;
    layer3_outputs(4025) <= not (a xor b);
    layer3_outputs(4026) <= b;
    layer3_outputs(4027) <= not b;
    layer3_outputs(4028) <= a or b;
    layer3_outputs(4029) <= not b;
    layer3_outputs(4030) <= a;
    layer3_outputs(4031) <= not (a and b);
    layer3_outputs(4032) <= b and not a;
    layer3_outputs(4033) <= not b;
    layer3_outputs(4034) <= not b or a;
    layer3_outputs(4035) <= a;
    layer3_outputs(4036) <= b;
    layer3_outputs(4037) <= a;
    layer3_outputs(4038) <= not b or a;
    layer3_outputs(4039) <= not a;
    layer3_outputs(4040) <= not (a or b);
    layer3_outputs(4041) <= '0';
    layer3_outputs(4042) <= a;
    layer3_outputs(4043) <= '0';
    layer3_outputs(4044) <= a xor b;
    layer3_outputs(4045) <= a;
    layer3_outputs(4046) <= not a or b;
    layer3_outputs(4047) <= not b;
    layer3_outputs(4048) <= not (a or b);
    layer3_outputs(4049) <= b;
    layer3_outputs(4050) <= not a;
    layer3_outputs(4051) <= a;
    layer3_outputs(4052) <= not a or b;
    layer3_outputs(4053) <= a xor b;
    layer3_outputs(4054) <= not b;
    layer3_outputs(4055) <= not a;
    layer3_outputs(4056) <= a;
    layer3_outputs(4057) <= not (a and b);
    layer3_outputs(4058) <= not (a and b);
    layer3_outputs(4059) <= a;
    layer3_outputs(4060) <= a or b;
    layer3_outputs(4061) <= a;
    layer3_outputs(4062) <= a xor b;
    layer3_outputs(4063) <= b and not a;
    layer3_outputs(4064) <= a and not b;
    layer3_outputs(4065) <= not (a or b);
    layer3_outputs(4066) <= '1';
    layer3_outputs(4067) <= a or b;
    layer3_outputs(4068) <= a xor b;
    layer3_outputs(4069) <= not (a or b);
    layer3_outputs(4070) <= a xor b;
    layer3_outputs(4071) <= not (a and b);
    layer3_outputs(4072) <= not (a and b);
    layer3_outputs(4073) <= a and not b;
    layer3_outputs(4074) <= a and b;
    layer3_outputs(4075) <= not (a or b);
    layer3_outputs(4076) <= not b;
    layer3_outputs(4077) <= not (a or b);
    layer3_outputs(4078) <= a and b;
    layer3_outputs(4079) <= not (a or b);
    layer3_outputs(4080) <= not (a and b);
    layer3_outputs(4081) <= not a;
    layer3_outputs(4082) <= a and not b;
    layer3_outputs(4083) <= a and b;
    layer3_outputs(4084) <= not (a and b);
    layer3_outputs(4085) <= b;
    layer3_outputs(4086) <= not (a and b);
    layer3_outputs(4087) <= not b;
    layer3_outputs(4088) <= not (a xor b);
    layer3_outputs(4089) <= a;
    layer3_outputs(4090) <= a or b;
    layer3_outputs(4091) <= not a or b;
    layer3_outputs(4092) <= b and not a;
    layer3_outputs(4093) <= a xor b;
    layer3_outputs(4094) <= a;
    layer3_outputs(4095) <= not a or b;
    layer3_outputs(4096) <= a;
    layer3_outputs(4097) <= b;
    layer3_outputs(4098) <= a xor b;
    layer3_outputs(4099) <= a or b;
    layer3_outputs(4100) <= a;
    layer3_outputs(4101) <= not (a and b);
    layer3_outputs(4102) <= not a or b;
    layer3_outputs(4103) <= b;
    layer3_outputs(4104) <= not a;
    layer3_outputs(4105) <= a;
    layer3_outputs(4106) <= a;
    layer3_outputs(4107) <= not (a xor b);
    layer3_outputs(4108) <= not b;
    layer3_outputs(4109) <= a and not b;
    layer3_outputs(4110) <= a and b;
    layer3_outputs(4111) <= '0';
    layer3_outputs(4112) <= a xor b;
    layer3_outputs(4113) <= not a;
    layer3_outputs(4114) <= b;
    layer3_outputs(4115) <= not b;
    layer3_outputs(4116) <= not b;
    layer3_outputs(4117) <= not (a and b);
    layer3_outputs(4118) <= not a or b;
    layer3_outputs(4119) <= b;
    layer3_outputs(4120) <= not b;
    layer3_outputs(4121) <= b;
    layer3_outputs(4122) <= a and not b;
    layer3_outputs(4123) <= '1';
    layer3_outputs(4124) <= b and not a;
    layer3_outputs(4125) <= not (a or b);
    layer3_outputs(4126) <= b;
    layer3_outputs(4127) <= a and b;
    layer3_outputs(4128) <= not a;
    layer3_outputs(4129) <= a or b;
    layer3_outputs(4130) <= not a;
    layer3_outputs(4131) <= a;
    layer3_outputs(4132) <= not b;
    layer3_outputs(4133) <= a and b;
    layer3_outputs(4134) <= not (a and b);
    layer3_outputs(4135) <= a or b;
    layer3_outputs(4136) <= not b or a;
    layer3_outputs(4137) <= not a;
    layer3_outputs(4138) <= '0';
    layer3_outputs(4139) <= a and not b;
    layer3_outputs(4140) <= not b or a;
    layer3_outputs(4141) <= not a or b;
    layer3_outputs(4142) <= not a;
    layer3_outputs(4143) <= b and not a;
    layer3_outputs(4144) <= not b;
    layer3_outputs(4145) <= not (a xor b);
    layer3_outputs(4146) <= b;
    layer3_outputs(4147) <= b;
    layer3_outputs(4148) <= a or b;
    layer3_outputs(4149) <= a;
    layer3_outputs(4150) <= '0';
    layer3_outputs(4151) <= a and not b;
    layer3_outputs(4152) <= b and not a;
    layer3_outputs(4153) <= b and not a;
    layer3_outputs(4154) <= a and b;
    layer3_outputs(4155) <= b;
    layer3_outputs(4156) <= a and b;
    layer3_outputs(4157) <= not a;
    layer3_outputs(4158) <= not (a and b);
    layer3_outputs(4159) <= a or b;
    layer3_outputs(4160) <= b and not a;
    layer3_outputs(4161) <= b;
    layer3_outputs(4162) <= '0';
    layer3_outputs(4163) <= a and b;
    layer3_outputs(4164) <= not b;
    layer3_outputs(4165) <= not b;
    layer3_outputs(4166) <= a and not b;
    layer3_outputs(4167) <= a xor b;
    layer3_outputs(4168) <= not a;
    layer3_outputs(4169) <= a or b;
    layer3_outputs(4170) <= a or b;
    layer3_outputs(4171) <= a and not b;
    layer3_outputs(4172) <= not b;
    layer3_outputs(4173) <= a xor b;
    layer3_outputs(4174) <= not b;
    layer3_outputs(4175) <= not (a and b);
    layer3_outputs(4176) <= a or b;
    layer3_outputs(4177) <= not (a and b);
    layer3_outputs(4178) <= '1';
    layer3_outputs(4179) <= a and not b;
    layer3_outputs(4180) <= not b or a;
    layer3_outputs(4181) <= b and not a;
    layer3_outputs(4182) <= not a or b;
    layer3_outputs(4183) <= b;
    layer3_outputs(4184) <= a;
    layer3_outputs(4185) <= '1';
    layer3_outputs(4186) <= a;
    layer3_outputs(4187) <= '0';
    layer3_outputs(4188) <= b and not a;
    layer3_outputs(4189) <= not b;
    layer3_outputs(4190) <= '1';
    layer3_outputs(4191) <= a or b;
    layer3_outputs(4192) <= '0';
    layer3_outputs(4193) <= a;
    layer3_outputs(4194) <= not a;
    layer3_outputs(4195) <= a;
    layer3_outputs(4196) <= not b;
    layer3_outputs(4197) <= a or b;
    layer3_outputs(4198) <= not a or b;
    layer3_outputs(4199) <= not (a and b);
    layer3_outputs(4200) <= not b;
    layer3_outputs(4201) <= '1';
    layer3_outputs(4202) <= b;
    layer3_outputs(4203) <= not (a and b);
    layer3_outputs(4204) <= a and not b;
    layer3_outputs(4205) <= not b;
    layer3_outputs(4206) <= not a or b;
    layer3_outputs(4207) <= not b or a;
    layer3_outputs(4208) <= not (a xor b);
    layer3_outputs(4209) <= a;
    layer3_outputs(4210) <= not (a and b);
    layer3_outputs(4211) <= a and not b;
    layer3_outputs(4212) <= a;
    layer3_outputs(4213) <= a;
    layer3_outputs(4214) <= not b;
    layer3_outputs(4215) <= not b or a;
    layer3_outputs(4216) <= not b or a;
    layer3_outputs(4217) <= '0';
    layer3_outputs(4218) <= '1';
    layer3_outputs(4219) <= b;
    layer3_outputs(4220) <= not (a and b);
    layer3_outputs(4221) <= not b;
    layer3_outputs(4222) <= a and b;
    layer3_outputs(4223) <= a;
    layer3_outputs(4224) <= a;
    layer3_outputs(4225) <= not b or a;
    layer3_outputs(4226) <= a or b;
    layer3_outputs(4227) <= not b or a;
    layer3_outputs(4228) <= b;
    layer3_outputs(4229) <= b and not a;
    layer3_outputs(4230) <= '0';
    layer3_outputs(4231) <= not (a xor b);
    layer3_outputs(4232) <= not a or b;
    layer3_outputs(4233) <= a xor b;
    layer3_outputs(4234) <= not b;
    layer3_outputs(4235) <= a;
    layer3_outputs(4236) <= not (a and b);
    layer3_outputs(4237) <= a;
    layer3_outputs(4238) <= not a or b;
    layer3_outputs(4239) <= not a or b;
    layer3_outputs(4240) <= a;
    layer3_outputs(4241) <= a and b;
    layer3_outputs(4242) <= a;
    layer3_outputs(4243) <= b;
    layer3_outputs(4244) <= not b or a;
    layer3_outputs(4245) <= a and not b;
    layer3_outputs(4246) <= not b;
    layer3_outputs(4247) <= b and not a;
    layer3_outputs(4248) <= a or b;
    layer3_outputs(4249) <= a xor b;
    layer3_outputs(4250) <= a;
    layer3_outputs(4251) <= not (a and b);
    layer3_outputs(4252) <= a;
    layer3_outputs(4253) <= not (a and b);
    layer3_outputs(4254) <= b;
    layer3_outputs(4255) <= not b or a;
    layer3_outputs(4256) <= a and b;
    layer3_outputs(4257) <= b;
    layer3_outputs(4258) <= a or b;
    layer3_outputs(4259) <= a or b;
    layer3_outputs(4260) <= a and b;
    layer3_outputs(4261) <= not (a or b);
    layer3_outputs(4262) <= a xor b;
    layer3_outputs(4263) <= not b;
    layer3_outputs(4264) <= a and b;
    layer3_outputs(4265) <= not a;
    layer3_outputs(4266) <= b;
    layer3_outputs(4267) <= a;
    layer3_outputs(4268) <= b;
    layer3_outputs(4269) <= a or b;
    layer3_outputs(4270) <= b;
    layer3_outputs(4271) <= not b or a;
    layer3_outputs(4272) <= b and not a;
    layer3_outputs(4273) <= a or b;
    layer3_outputs(4274) <= not a or b;
    layer3_outputs(4275) <= '1';
    layer3_outputs(4276) <= not a or b;
    layer3_outputs(4277) <= not (a and b);
    layer3_outputs(4278) <= not (a or b);
    layer3_outputs(4279) <= not b;
    layer3_outputs(4280) <= '1';
    layer3_outputs(4281) <= b;
    layer3_outputs(4282) <= not (a and b);
    layer3_outputs(4283) <= a and not b;
    layer3_outputs(4284) <= b;
    layer3_outputs(4285) <= a and b;
    layer3_outputs(4286) <= a xor b;
    layer3_outputs(4287) <= a and b;
    layer3_outputs(4288) <= a;
    layer3_outputs(4289) <= not b;
    layer3_outputs(4290) <= not b or a;
    layer3_outputs(4291) <= not b;
    layer3_outputs(4292) <= not b;
    layer3_outputs(4293) <= not b;
    layer3_outputs(4294) <= not (a and b);
    layer3_outputs(4295) <= b;
    layer3_outputs(4296) <= '0';
    layer3_outputs(4297) <= b;
    layer3_outputs(4298) <= a;
    layer3_outputs(4299) <= a and not b;
    layer3_outputs(4300) <= b;
    layer3_outputs(4301) <= not a or b;
    layer3_outputs(4302) <= not b;
    layer3_outputs(4303) <= not (a and b);
    layer3_outputs(4304) <= not (a xor b);
    layer3_outputs(4305) <= b and not a;
    layer3_outputs(4306) <= not a;
    layer3_outputs(4307) <= not a;
    layer3_outputs(4308) <= not b or a;
    layer3_outputs(4309) <= not a;
    layer3_outputs(4310) <= b;
    layer3_outputs(4311) <= b and not a;
    layer3_outputs(4312) <= a and not b;
    layer3_outputs(4313) <= not (a xor b);
    layer3_outputs(4314) <= not a;
    layer3_outputs(4315) <= not b;
    layer3_outputs(4316) <= not b;
    layer3_outputs(4317) <= not a or b;
    layer3_outputs(4318) <= b and not a;
    layer3_outputs(4319) <= not b;
    layer3_outputs(4320) <= not b or a;
    layer3_outputs(4321) <= b and not a;
    layer3_outputs(4322) <= b;
    layer3_outputs(4323) <= a and not b;
    layer3_outputs(4324) <= b and not a;
    layer3_outputs(4325) <= not (a or b);
    layer3_outputs(4326) <= not a;
    layer3_outputs(4327) <= not (a and b);
    layer3_outputs(4328) <= a;
    layer3_outputs(4329) <= not b or a;
    layer3_outputs(4330) <= a and not b;
    layer3_outputs(4331) <= a;
    layer3_outputs(4332) <= not b or a;
    layer3_outputs(4333) <= b and not a;
    layer3_outputs(4334) <= not a;
    layer3_outputs(4335) <= not b;
    layer3_outputs(4336) <= '0';
    layer3_outputs(4337) <= not a;
    layer3_outputs(4338) <= b;
    layer3_outputs(4339) <= a;
    layer3_outputs(4340) <= not a;
    layer3_outputs(4341) <= b and not a;
    layer3_outputs(4342) <= b;
    layer3_outputs(4343) <= not a;
    layer3_outputs(4344) <= not b;
    layer3_outputs(4345) <= a;
    layer3_outputs(4346) <= b;
    layer3_outputs(4347) <= b and not a;
    layer3_outputs(4348) <= b;
    layer3_outputs(4349) <= a or b;
    layer3_outputs(4350) <= b;
    layer3_outputs(4351) <= a xor b;
    layer3_outputs(4352) <= b;
    layer3_outputs(4353) <= b;
    layer3_outputs(4354) <= not (a xor b);
    layer3_outputs(4355) <= not b;
    layer3_outputs(4356) <= not (a or b);
    layer3_outputs(4357) <= not a;
    layer3_outputs(4358) <= a and not b;
    layer3_outputs(4359) <= '0';
    layer3_outputs(4360) <= a;
    layer3_outputs(4361) <= not (a or b);
    layer3_outputs(4362) <= b and not a;
    layer3_outputs(4363) <= '0';
    layer3_outputs(4364) <= a or b;
    layer3_outputs(4365) <= not (a xor b);
    layer3_outputs(4366) <= not a or b;
    layer3_outputs(4367) <= not (a or b);
    layer3_outputs(4368) <= not a;
    layer3_outputs(4369) <= a;
    layer3_outputs(4370) <= not b;
    layer3_outputs(4371) <= b and not a;
    layer3_outputs(4372) <= '1';
    layer3_outputs(4373) <= not (a xor b);
    layer3_outputs(4374) <= a and not b;
    layer3_outputs(4375) <= not (a or b);
    layer3_outputs(4376) <= a;
    layer3_outputs(4377) <= not a;
    layer3_outputs(4378) <= '1';
    layer3_outputs(4379) <= not a or b;
    layer3_outputs(4380) <= not b or a;
    layer3_outputs(4381) <= not b or a;
    layer3_outputs(4382) <= not (a or b);
    layer3_outputs(4383) <= a or b;
    layer3_outputs(4384) <= not a;
    layer3_outputs(4385) <= a xor b;
    layer3_outputs(4386) <= b;
    layer3_outputs(4387) <= not (a or b);
    layer3_outputs(4388) <= a and not b;
    layer3_outputs(4389) <= a or b;
    layer3_outputs(4390) <= not b;
    layer3_outputs(4391) <= a;
    layer3_outputs(4392) <= not a;
    layer3_outputs(4393) <= not (a and b);
    layer3_outputs(4394) <= not (a and b);
    layer3_outputs(4395) <= not a;
    layer3_outputs(4396) <= not a or b;
    layer3_outputs(4397) <= not b;
    layer3_outputs(4398) <= b;
    layer3_outputs(4399) <= a xor b;
    layer3_outputs(4400) <= a xor b;
    layer3_outputs(4401) <= a and not b;
    layer3_outputs(4402) <= a or b;
    layer3_outputs(4403) <= not (a and b);
    layer3_outputs(4404) <= a;
    layer3_outputs(4405) <= a and not b;
    layer3_outputs(4406) <= a or b;
    layer3_outputs(4407) <= not a or b;
    layer3_outputs(4408) <= not a;
    layer3_outputs(4409) <= not a or b;
    layer3_outputs(4410) <= a or b;
    layer3_outputs(4411) <= a;
    layer3_outputs(4412) <= not a;
    layer3_outputs(4413) <= not (a or b);
    layer3_outputs(4414) <= b;
    layer3_outputs(4415) <= a or b;
    layer3_outputs(4416) <= a and b;
    layer3_outputs(4417) <= not (a xor b);
    layer3_outputs(4418) <= not a;
    layer3_outputs(4419) <= not (a and b);
    layer3_outputs(4420) <= not b;
    layer3_outputs(4421) <= b and not a;
    layer3_outputs(4422) <= not b;
    layer3_outputs(4423) <= not a or b;
    layer3_outputs(4424) <= '0';
    layer3_outputs(4425) <= not b or a;
    layer3_outputs(4426) <= b;
    layer3_outputs(4427) <= a or b;
    layer3_outputs(4428) <= a and b;
    layer3_outputs(4429) <= not a;
    layer3_outputs(4430) <= a or b;
    layer3_outputs(4431) <= b and not a;
    layer3_outputs(4432) <= a or b;
    layer3_outputs(4433) <= a;
    layer3_outputs(4434) <= not a;
    layer3_outputs(4435) <= a or b;
    layer3_outputs(4436) <= '0';
    layer3_outputs(4437) <= not b or a;
    layer3_outputs(4438) <= not a;
    layer3_outputs(4439) <= '1';
    layer3_outputs(4440) <= a or b;
    layer3_outputs(4441) <= not (a and b);
    layer3_outputs(4442) <= not a;
    layer3_outputs(4443) <= b and not a;
    layer3_outputs(4444) <= not (a or b);
    layer3_outputs(4445) <= not b;
    layer3_outputs(4446) <= b;
    layer3_outputs(4447) <= b and not a;
    layer3_outputs(4448) <= '1';
    layer3_outputs(4449) <= a or b;
    layer3_outputs(4450) <= not b;
    layer3_outputs(4451) <= not (a and b);
    layer3_outputs(4452) <= b;
    layer3_outputs(4453) <= not (a and b);
    layer3_outputs(4454) <= '1';
    layer3_outputs(4455) <= '0';
    layer3_outputs(4456) <= not b or a;
    layer3_outputs(4457) <= not b;
    layer3_outputs(4458) <= not (a or b);
    layer3_outputs(4459) <= '0';
    layer3_outputs(4460) <= a or b;
    layer3_outputs(4461) <= not a or b;
    layer3_outputs(4462) <= not a or b;
    layer3_outputs(4463) <= b and not a;
    layer3_outputs(4464) <= b;
    layer3_outputs(4465) <= not (a and b);
    layer3_outputs(4466) <= '1';
    layer3_outputs(4467) <= '1';
    layer3_outputs(4468) <= a;
    layer3_outputs(4469) <= a;
    layer3_outputs(4470) <= not (a and b);
    layer3_outputs(4471) <= b;
    layer3_outputs(4472) <= not b;
    layer3_outputs(4473) <= b;
    layer3_outputs(4474) <= a;
    layer3_outputs(4475) <= a;
    layer3_outputs(4476) <= a and b;
    layer3_outputs(4477) <= not a;
    layer3_outputs(4478) <= a or b;
    layer3_outputs(4479) <= not b or a;
    layer3_outputs(4480) <= not (a or b);
    layer3_outputs(4481) <= a or b;
    layer3_outputs(4482) <= a;
    layer3_outputs(4483) <= a and not b;
    layer3_outputs(4484) <= not b or a;
    layer3_outputs(4485) <= a or b;
    layer3_outputs(4486) <= b;
    layer3_outputs(4487) <= a or b;
    layer3_outputs(4488) <= not b;
    layer3_outputs(4489) <= not b or a;
    layer3_outputs(4490) <= not b or a;
    layer3_outputs(4491) <= a and b;
    layer3_outputs(4492) <= not b;
    layer3_outputs(4493) <= b;
    layer3_outputs(4494) <= b;
    layer3_outputs(4495) <= not b or a;
    layer3_outputs(4496) <= b;
    layer3_outputs(4497) <= not (a xor b);
    layer3_outputs(4498) <= not b;
    layer3_outputs(4499) <= '1';
    layer3_outputs(4500) <= b;
    layer3_outputs(4501) <= '1';
    layer3_outputs(4502) <= not a or b;
    layer3_outputs(4503) <= not (a or b);
    layer3_outputs(4504) <= b;
    layer3_outputs(4505) <= b and not a;
    layer3_outputs(4506) <= not (a or b);
    layer3_outputs(4507) <= not (a xor b);
    layer3_outputs(4508) <= a;
    layer3_outputs(4509) <= not b or a;
    layer3_outputs(4510) <= b and not a;
    layer3_outputs(4511) <= b;
    layer3_outputs(4512) <= not a or b;
    layer3_outputs(4513) <= a and b;
    layer3_outputs(4514) <= not b;
    layer3_outputs(4515) <= a;
    layer3_outputs(4516) <= a;
    layer3_outputs(4517) <= a and b;
    layer3_outputs(4518) <= not a;
    layer3_outputs(4519) <= b;
    layer3_outputs(4520) <= not a;
    layer3_outputs(4521) <= a xor b;
    layer3_outputs(4522) <= a and not b;
    layer3_outputs(4523) <= not (a and b);
    layer3_outputs(4524) <= b and not a;
    layer3_outputs(4525) <= '0';
    layer3_outputs(4526) <= not a;
    layer3_outputs(4527) <= not (a or b);
    layer3_outputs(4528) <= b and not a;
    layer3_outputs(4529) <= not a or b;
    layer3_outputs(4530) <= not a;
    layer3_outputs(4531) <= b;
    layer3_outputs(4532) <= not b or a;
    layer3_outputs(4533) <= '0';
    layer3_outputs(4534) <= not a;
    layer3_outputs(4535) <= b;
    layer3_outputs(4536) <= a or b;
    layer3_outputs(4537) <= not (a xor b);
    layer3_outputs(4538) <= not b;
    layer3_outputs(4539) <= b and not a;
    layer3_outputs(4540) <= not a;
    layer3_outputs(4541) <= a or b;
    layer3_outputs(4542) <= not b;
    layer3_outputs(4543) <= a and not b;
    layer3_outputs(4544) <= a and b;
    layer3_outputs(4545) <= not a or b;
    layer3_outputs(4546) <= a;
    layer3_outputs(4547) <= a;
    layer3_outputs(4548) <= not (a or b);
    layer3_outputs(4549) <= not b;
    layer3_outputs(4550) <= a xor b;
    layer3_outputs(4551) <= not b or a;
    layer3_outputs(4552) <= not a or b;
    layer3_outputs(4553) <= a;
    layer3_outputs(4554) <= not a;
    layer3_outputs(4555) <= a and not b;
    layer3_outputs(4556) <= not a;
    layer3_outputs(4557) <= not (a or b);
    layer3_outputs(4558) <= not b;
    layer3_outputs(4559) <= not b;
    layer3_outputs(4560) <= '0';
    layer3_outputs(4561) <= not a or b;
    layer3_outputs(4562) <= not a or b;
    layer3_outputs(4563) <= not a;
    layer3_outputs(4564) <= not b;
    layer3_outputs(4565) <= b;
    layer3_outputs(4566) <= not b;
    layer3_outputs(4567) <= a;
    layer3_outputs(4568) <= a or b;
    layer3_outputs(4569) <= '0';
    layer3_outputs(4570) <= '1';
    layer3_outputs(4571) <= a xor b;
    layer3_outputs(4572) <= a or b;
    layer3_outputs(4573) <= not (a xor b);
    layer3_outputs(4574) <= not b;
    layer3_outputs(4575) <= '0';
    layer3_outputs(4576) <= a or b;
    layer3_outputs(4577) <= not (a and b);
    layer3_outputs(4578) <= '1';
    layer3_outputs(4579) <= b;
    layer3_outputs(4580) <= a or b;
    layer3_outputs(4581) <= not b or a;
    layer3_outputs(4582) <= not (a and b);
    layer3_outputs(4583) <= not (a and b);
    layer3_outputs(4584) <= not a;
    layer3_outputs(4585) <= b;
    layer3_outputs(4586) <= not a;
    layer3_outputs(4587) <= a and not b;
    layer3_outputs(4588) <= a;
    layer3_outputs(4589) <= a xor b;
    layer3_outputs(4590) <= not b or a;
    layer3_outputs(4591) <= b and not a;
    layer3_outputs(4592) <= '0';
    layer3_outputs(4593) <= b and not a;
    layer3_outputs(4594) <= a xor b;
    layer3_outputs(4595) <= not b or a;
    layer3_outputs(4596) <= not a;
    layer3_outputs(4597) <= not b;
    layer3_outputs(4598) <= not (a xor b);
    layer3_outputs(4599) <= a;
    layer3_outputs(4600) <= not a or b;
    layer3_outputs(4601) <= a;
    layer3_outputs(4602) <= a and b;
    layer3_outputs(4603) <= a and b;
    layer3_outputs(4604) <= '1';
    layer3_outputs(4605) <= b;
    layer3_outputs(4606) <= '1';
    layer3_outputs(4607) <= not (a or b);
    layer3_outputs(4608) <= not (a and b);
    layer3_outputs(4609) <= a or b;
    layer3_outputs(4610) <= a;
    layer3_outputs(4611) <= not a;
    layer3_outputs(4612) <= not (a or b);
    layer3_outputs(4613) <= not (a and b);
    layer3_outputs(4614) <= not b or a;
    layer3_outputs(4615) <= b;
    layer3_outputs(4616) <= a and b;
    layer3_outputs(4617) <= b;
    layer3_outputs(4618) <= a and b;
    layer3_outputs(4619) <= a;
    layer3_outputs(4620) <= not a;
    layer3_outputs(4621) <= a and b;
    layer3_outputs(4622) <= not (a and b);
    layer3_outputs(4623) <= not (a or b);
    layer3_outputs(4624) <= a and b;
    layer3_outputs(4625) <= a and not b;
    layer3_outputs(4626) <= not b or a;
    layer3_outputs(4627) <= b;
    layer3_outputs(4628) <= a and b;
    layer3_outputs(4629) <= '1';
    layer3_outputs(4630) <= not (a and b);
    layer3_outputs(4631) <= not (a and b);
    layer3_outputs(4632) <= a and not b;
    layer3_outputs(4633) <= not (a and b);
    layer3_outputs(4634) <= a and b;
    layer3_outputs(4635) <= '0';
    layer3_outputs(4636) <= a;
    layer3_outputs(4637) <= not a;
    layer3_outputs(4638) <= not b or a;
    layer3_outputs(4639) <= a and not b;
    layer3_outputs(4640) <= '0';
    layer3_outputs(4641) <= a and b;
    layer3_outputs(4642) <= not a;
    layer3_outputs(4643) <= a and not b;
    layer3_outputs(4644) <= a xor b;
    layer3_outputs(4645) <= a;
    layer3_outputs(4646) <= a or b;
    layer3_outputs(4647) <= a or b;
    layer3_outputs(4648) <= not b;
    layer3_outputs(4649) <= b and not a;
    layer3_outputs(4650) <= b;
    layer3_outputs(4651) <= b;
    layer3_outputs(4652) <= not a;
    layer3_outputs(4653) <= not b;
    layer3_outputs(4654) <= not a or b;
    layer3_outputs(4655) <= not b or a;
    layer3_outputs(4656) <= not (a xor b);
    layer3_outputs(4657) <= not b;
    layer3_outputs(4658) <= not a;
    layer3_outputs(4659) <= not b or a;
    layer3_outputs(4660) <= a and not b;
    layer3_outputs(4661) <= a and b;
    layer3_outputs(4662) <= '0';
    layer3_outputs(4663) <= not (a xor b);
    layer3_outputs(4664) <= b and not a;
    layer3_outputs(4665) <= not b;
    layer3_outputs(4666) <= not a;
    layer3_outputs(4667) <= not b or a;
    layer3_outputs(4668) <= a or b;
    layer3_outputs(4669) <= not (a and b);
    layer3_outputs(4670) <= not b or a;
    layer3_outputs(4671) <= not b or a;
    layer3_outputs(4672) <= not (a and b);
    layer3_outputs(4673) <= a;
    layer3_outputs(4674) <= b and not a;
    layer3_outputs(4675) <= not (a or b);
    layer3_outputs(4676) <= a and not b;
    layer3_outputs(4677) <= not (a and b);
    layer3_outputs(4678) <= not (a or b);
    layer3_outputs(4679) <= b;
    layer3_outputs(4680) <= a or b;
    layer3_outputs(4681) <= b;
    layer3_outputs(4682) <= not a or b;
    layer3_outputs(4683) <= not a or b;
    layer3_outputs(4684) <= not b or a;
    layer3_outputs(4685) <= b;
    layer3_outputs(4686) <= a or b;
    layer3_outputs(4687) <= b and not a;
    layer3_outputs(4688) <= a;
    layer3_outputs(4689) <= not a;
    layer3_outputs(4690) <= a xor b;
    layer3_outputs(4691) <= b;
    layer3_outputs(4692) <= not b or a;
    layer3_outputs(4693) <= not (a xor b);
    layer3_outputs(4694) <= not b or a;
    layer3_outputs(4695) <= '1';
    layer3_outputs(4696) <= not b or a;
    layer3_outputs(4697) <= a xor b;
    layer3_outputs(4698) <= not (a and b);
    layer3_outputs(4699) <= not a;
    layer3_outputs(4700) <= b;
    layer3_outputs(4701) <= not a;
    layer3_outputs(4702) <= b;
    layer3_outputs(4703) <= b and not a;
    layer3_outputs(4704) <= b and not a;
    layer3_outputs(4705) <= b and not a;
    layer3_outputs(4706) <= a;
    layer3_outputs(4707) <= a;
    layer3_outputs(4708) <= a;
    layer3_outputs(4709) <= not (a or b);
    layer3_outputs(4710) <= not (a xor b);
    layer3_outputs(4711) <= a or b;
    layer3_outputs(4712) <= not a or b;
    layer3_outputs(4713) <= not b;
    layer3_outputs(4714) <= '0';
    layer3_outputs(4715) <= a and not b;
    layer3_outputs(4716) <= b and not a;
    layer3_outputs(4717) <= a or b;
    layer3_outputs(4718) <= a;
    layer3_outputs(4719) <= not a;
    layer3_outputs(4720) <= '0';
    layer3_outputs(4721) <= a;
    layer3_outputs(4722) <= a and not b;
    layer3_outputs(4723) <= not a;
    layer3_outputs(4724) <= a;
    layer3_outputs(4725) <= a xor b;
    layer3_outputs(4726) <= not (a and b);
    layer3_outputs(4727) <= '1';
    layer3_outputs(4728) <= a and b;
    layer3_outputs(4729) <= '0';
    layer3_outputs(4730) <= not b;
    layer3_outputs(4731) <= a and b;
    layer3_outputs(4732) <= not (a or b);
    layer3_outputs(4733) <= not a;
    layer3_outputs(4734) <= a and not b;
    layer3_outputs(4735) <= a and b;
    layer3_outputs(4736) <= b;
    layer3_outputs(4737) <= a or b;
    layer3_outputs(4738) <= b;
    layer3_outputs(4739) <= not a or b;
    layer3_outputs(4740) <= not (a and b);
    layer3_outputs(4741) <= not (a or b);
    layer3_outputs(4742) <= not a;
    layer3_outputs(4743) <= b;
    layer3_outputs(4744) <= not (a xor b);
    layer3_outputs(4745) <= a and not b;
    layer3_outputs(4746) <= '0';
    layer3_outputs(4747) <= a;
    layer3_outputs(4748) <= '1';
    layer3_outputs(4749) <= not (a and b);
    layer3_outputs(4750) <= a;
    layer3_outputs(4751) <= a and b;
    layer3_outputs(4752) <= b;
    layer3_outputs(4753) <= not b;
    layer3_outputs(4754) <= not a or b;
    layer3_outputs(4755) <= b and not a;
    layer3_outputs(4756) <= a or b;
    layer3_outputs(4757) <= not b or a;
    layer3_outputs(4758) <= b and not a;
    layer3_outputs(4759) <= a or b;
    layer3_outputs(4760) <= '1';
    layer3_outputs(4761) <= not b or a;
    layer3_outputs(4762) <= a;
    layer3_outputs(4763) <= a and not b;
    layer3_outputs(4764) <= not (a and b);
    layer3_outputs(4765) <= a or b;
    layer3_outputs(4766) <= a and not b;
    layer3_outputs(4767) <= not a;
    layer3_outputs(4768) <= b and not a;
    layer3_outputs(4769) <= not (a xor b);
    layer3_outputs(4770) <= a;
    layer3_outputs(4771) <= not b;
    layer3_outputs(4772) <= not b;
    layer3_outputs(4773) <= a;
    layer3_outputs(4774) <= not (a and b);
    layer3_outputs(4775) <= '1';
    layer3_outputs(4776) <= a;
    layer3_outputs(4777) <= a or b;
    layer3_outputs(4778) <= a and b;
    layer3_outputs(4779) <= not b or a;
    layer3_outputs(4780) <= a and not b;
    layer3_outputs(4781) <= a or b;
    layer3_outputs(4782) <= not b or a;
    layer3_outputs(4783) <= a;
    layer3_outputs(4784) <= not (a xor b);
    layer3_outputs(4785) <= not b or a;
    layer3_outputs(4786) <= a or b;
    layer3_outputs(4787) <= not (a or b);
    layer3_outputs(4788) <= b;
    layer3_outputs(4789) <= not b or a;
    layer3_outputs(4790) <= not b or a;
    layer3_outputs(4791) <= not a;
    layer3_outputs(4792) <= b;
    layer3_outputs(4793) <= not a or b;
    layer3_outputs(4794) <= not (a or b);
    layer3_outputs(4795) <= a;
    layer3_outputs(4796) <= not a;
    layer3_outputs(4797) <= not (a or b);
    layer3_outputs(4798) <= not a or b;
    layer3_outputs(4799) <= not (a and b);
    layer3_outputs(4800) <= b;
    layer3_outputs(4801) <= not b or a;
    layer3_outputs(4802) <= not a or b;
    layer3_outputs(4803) <= not a;
    layer3_outputs(4804) <= a xor b;
    layer3_outputs(4805) <= '0';
    layer3_outputs(4806) <= not a;
    layer3_outputs(4807) <= not b;
    layer3_outputs(4808) <= not (a or b);
    layer3_outputs(4809) <= not b or a;
    layer3_outputs(4810) <= a and b;
    layer3_outputs(4811) <= '0';
    layer3_outputs(4812) <= not b;
    layer3_outputs(4813) <= '0';
    layer3_outputs(4814) <= not a or b;
    layer3_outputs(4815) <= not a;
    layer3_outputs(4816) <= not b or a;
    layer3_outputs(4817) <= not b;
    layer3_outputs(4818) <= not b or a;
    layer3_outputs(4819) <= a and b;
    layer3_outputs(4820) <= not b or a;
    layer3_outputs(4821) <= not a or b;
    layer3_outputs(4822) <= b;
    layer3_outputs(4823) <= not (a and b);
    layer3_outputs(4824) <= a;
    layer3_outputs(4825) <= a and not b;
    layer3_outputs(4826) <= a xor b;
    layer3_outputs(4827) <= not b;
    layer3_outputs(4828) <= not b or a;
    layer3_outputs(4829) <= '1';
    layer3_outputs(4830) <= a xor b;
    layer3_outputs(4831) <= not (a and b);
    layer3_outputs(4832) <= '0';
    layer3_outputs(4833) <= not (a or b);
    layer3_outputs(4834) <= b;
    layer3_outputs(4835) <= a and b;
    layer3_outputs(4836) <= not (a or b);
    layer3_outputs(4837) <= b;
    layer3_outputs(4838) <= a xor b;
    layer3_outputs(4839) <= a;
    layer3_outputs(4840) <= a xor b;
    layer3_outputs(4841) <= not a or b;
    layer3_outputs(4842) <= not (a xor b);
    layer3_outputs(4843) <= not a or b;
    layer3_outputs(4844) <= not (a or b);
    layer3_outputs(4845) <= b;
    layer3_outputs(4846) <= a xor b;
    layer3_outputs(4847) <= b and not a;
    layer3_outputs(4848) <= not b;
    layer3_outputs(4849) <= not a;
    layer3_outputs(4850) <= b and not a;
    layer3_outputs(4851) <= b;
    layer3_outputs(4852) <= not a;
    layer3_outputs(4853) <= not b or a;
    layer3_outputs(4854) <= a or b;
    layer3_outputs(4855) <= a xor b;
    layer3_outputs(4856) <= a and b;
    layer3_outputs(4857) <= a xor b;
    layer3_outputs(4858) <= not b or a;
    layer3_outputs(4859) <= not (a and b);
    layer3_outputs(4860) <= a and b;
    layer3_outputs(4861) <= not b;
    layer3_outputs(4862) <= a and not b;
    layer3_outputs(4863) <= not a;
    layer3_outputs(4864) <= a;
    layer3_outputs(4865) <= a and b;
    layer3_outputs(4866) <= '1';
    layer3_outputs(4867) <= not a or b;
    layer3_outputs(4868) <= b and not a;
    layer3_outputs(4869) <= not (a xor b);
    layer3_outputs(4870) <= a and not b;
    layer3_outputs(4871) <= a or b;
    layer3_outputs(4872) <= not b;
    layer3_outputs(4873) <= a;
    layer3_outputs(4874) <= b and not a;
    layer3_outputs(4875) <= a and not b;
    layer3_outputs(4876) <= not b;
    layer3_outputs(4877) <= a;
    layer3_outputs(4878) <= not b;
    layer3_outputs(4879) <= not b;
    layer3_outputs(4880) <= b and not a;
    layer3_outputs(4881) <= a;
    layer3_outputs(4882) <= a or b;
    layer3_outputs(4883) <= not (a or b);
    layer3_outputs(4884) <= not b;
    layer3_outputs(4885) <= b;
    layer3_outputs(4886) <= not a or b;
    layer3_outputs(4887) <= '0';
    layer3_outputs(4888) <= not b or a;
    layer3_outputs(4889) <= a or b;
    layer3_outputs(4890) <= not (a and b);
    layer3_outputs(4891) <= '1';
    layer3_outputs(4892) <= not b or a;
    layer3_outputs(4893) <= not (a or b);
    layer3_outputs(4894) <= b;
    layer3_outputs(4895) <= not (a xor b);
    layer3_outputs(4896) <= not b;
    layer3_outputs(4897) <= not a or b;
    layer3_outputs(4898) <= b;
    layer3_outputs(4899) <= not a or b;
    layer3_outputs(4900) <= b;
    layer3_outputs(4901) <= not (a or b);
    layer3_outputs(4902) <= a and not b;
    layer3_outputs(4903) <= not a;
    layer3_outputs(4904) <= a and b;
    layer3_outputs(4905) <= a;
    layer3_outputs(4906) <= b;
    layer3_outputs(4907) <= b;
    layer3_outputs(4908) <= not (a xor b);
    layer3_outputs(4909) <= a and b;
    layer3_outputs(4910) <= b and not a;
    layer3_outputs(4911) <= a;
    layer3_outputs(4912) <= a xor b;
    layer3_outputs(4913) <= not a;
    layer3_outputs(4914) <= a xor b;
    layer3_outputs(4915) <= b and not a;
    layer3_outputs(4916) <= b and not a;
    layer3_outputs(4917) <= not b;
    layer3_outputs(4918) <= a xor b;
    layer3_outputs(4919) <= not a or b;
    layer3_outputs(4920) <= not b;
    layer3_outputs(4921) <= not b;
    layer3_outputs(4922) <= not a or b;
    layer3_outputs(4923) <= not b;
    layer3_outputs(4924) <= not b or a;
    layer3_outputs(4925) <= a xor b;
    layer3_outputs(4926) <= a and b;
    layer3_outputs(4927) <= not b or a;
    layer3_outputs(4928) <= a and b;
    layer3_outputs(4929) <= not (a and b);
    layer3_outputs(4930) <= not a or b;
    layer3_outputs(4931) <= a and not b;
    layer3_outputs(4932) <= b;
    layer3_outputs(4933) <= not (a or b);
    layer3_outputs(4934) <= b;
    layer3_outputs(4935) <= '0';
    layer3_outputs(4936) <= not b or a;
    layer3_outputs(4937) <= not a;
    layer3_outputs(4938) <= not (a or b);
    layer3_outputs(4939) <= b and not a;
    layer3_outputs(4940) <= a and b;
    layer3_outputs(4941) <= not (a or b);
    layer3_outputs(4942) <= not (a or b);
    layer3_outputs(4943) <= not (a or b);
    layer3_outputs(4944) <= a or b;
    layer3_outputs(4945) <= b and not a;
    layer3_outputs(4946) <= a;
    layer3_outputs(4947) <= a xor b;
    layer3_outputs(4948) <= not b;
    layer3_outputs(4949) <= '0';
    layer3_outputs(4950) <= b;
    layer3_outputs(4951) <= not a or b;
    layer3_outputs(4952) <= a and b;
    layer3_outputs(4953) <= a or b;
    layer3_outputs(4954) <= not a;
    layer3_outputs(4955) <= '0';
    layer3_outputs(4956) <= not a;
    layer3_outputs(4957) <= not b;
    layer3_outputs(4958) <= not (a and b);
    layer3_outputs(4959) <= not (a and b);
    layer3_outputs(4960) <= a or b;
    layer3_outputs(4961) <= not a or b;
    layer3_outputs(4962) <= not a;
    layer3_outputs(4963) <= not b;
    layer3_outputs(4964) <= not b or a;
    layer3_outputs(4965) <= not (a xor b);
    layer3_outputs(4966) <= not b;
    layer3_outputs(4967) <= a;
    layer3_outputs(4968) <= not a or b;
    layer3_outputs(4969) <= b and not a;
    layer3_outputs(4970) <= not (a and b);
    layer3_outputs(4971) <= b and not a;
    layer3_outputs(4972) <= b;
    layer3_outputs(4973) <= not (a or b);
    layer3_outputs(4974) <= not a;
    layer3_outputs(4975) <= not (a and b);
    layer3_outputs(4976) <= not a or b;
    layer3_outputs(4977) <= not b;
    layer3_outputs(4978) <= not b or a;
    layer3_outputs(4979) <= a;
    layer3_outputs(4980) <= not b or a;
    layer3_outputs(4981) <= not (a xor b);
    layer3_outputs(4982) <= a or b;
    layer3_outputs(4983) <= not b;
    layer3_outputs(4984) <= a and not b;
    layer3_outputs(4985) <= a;
    layer3_outputs(4986) <= a;
    layer3_outputs(4987) <= not b;
    layer3_outputs(4988) <= a and not b;
    layer3_outputs(4989) <= a;
    layer3_outputs(4990) <= not b;
    layer3_outputs(4991) <= not a;
    layer3_outputs(4992) <= not a or b;
    layer3_outputs(4993) <= a xor b;
    layer3_outputs(4994) <= not (a xor b);
    layer3_outputs(4995) <= a;
    layer3_outputs(4996) <= not (a and b);
    layer3_outputs(4997) <= not b or a;
    layer3_outputs(4998) <= not (a or b);
    layer3_outputs(4999) <= a and not b;
    layer3_outputs(5000) <= not (a or b);
    layer3_outputs(5001) <= not a or b;
    layer3_outputs(5002) <= b;
    layer3_outputs(5003) <= not a;
    layer3_outputs(5004) <= a and not b;
    layer3_outputs(5005) <= not (a or b);
    layer3_outputs(5006) <= b;
    layer3_outputs(5007) <= not (a and b);
    layer3_outputs(5008) <= a or b;
    layer3_outputs(5009) <= '0';
    layer3_outputs(5010) <= b and not a;
    layer3_outputs(5011) <= not b;
    layer3_outputs(5012) <= '0';
    layer3_outputs(5013) <= '1';
    layer3_outputs(5014) <= not (a or b);
    layer3_outputs(5015) <= not a;
    layer3_outputs(5016) <= not (a or b);
    layer3_outputs(5017) <= '1';
    layer3_outputs(5018) <= not b;
    layer3_outputs(5019) <= a and not b;
    layer3_outputs(5020) <= not a;
    layer3_outputs(5021) <= not (a and b);
    layer3_outputs(5022) <= not a or b;
    layer3_outputs(5023) <= a and not b;
    layer3_outputs(5024) <= b;
    layer3_outputs(5025) <= not a or b;
    layer3_outputs(5026) <= b;
    layer3_outputs(5027) <= not (a xor b);
    layer3_outputs(5028) <= not (a and b);
    layer3_outputs(5029) <= b;
    layer3_outputs(5030) <= not b or a;
    layer3_outputs(5031) <= b and not a;
    layer3_outputs(5032) <= b;
    layer3_outputs(5033) <= not a;
    layer3_outputs(5034) <= not b;
    layer3_outputs(5035) <= not (a xor b);
    layer3_outputs(5036) <= a or b;
    layer3_outputs(5037) <= not b or a;
    layer3_outputs(5038) <= b and not a;
    layer3_outputs(5039) <= a;
    layer3_outputs(5040) <= '0';
    layer3_outputs(5041) <= not b or a;
    layer3_outputs(5042) <= a and not b;
    layer3_outputs(5043) <= b;
    layer3_outputs(5044) <= a and b;
    layer3_outputs(5045) <= a;
    layer3_outputs(5046) <= not b;
    layer3_outputs(5047) <= not a;
    layer3_outputs(5048) <= not a;
    layer3_outputs(5049) <= not a;
    layer3_outputs(5050) <= '0';
    layer3_outputs(5051) <= a;
    layer3_outputs(5052) <= not (a or b);
    layer3_outputs(5053) <= a or b;
    layer3_outputs(5054) <= not (a or b);
    layer3_outputs(5055) <= not b or a;
    layer3_outputs(5056) <= not a;
    layer3_outputs(5057) <= b;
    layer3_outputs(5058) <= a xor b;
    layer3_outputs(5059) <= a xor b;
    layer3_outputs(5060) <= '1';
    layer3_outputs(5061) <= not b;
    layer3_outputs(5062) <= not a;
    layer3_outputs(5063) <= not a or b;
    layer3_outputs(5064) <= '1';
    layer3_outputs(5065) <= '0';
    layer3_outputs(5066) <= a;
    layer3_outputs(5067) <= not (a and b);
    layer3_outputs(5068) <= a;
    layer3_outputs(5069) <= not a or b;
    layer3_outputs(5070) <= '0';
    layer3_outputs(5071) <= not (a and b);
    layer3_outputs(5072) <= b;
    layer3_outputs(5073) <= not b;
    layer3_outputs(5074) <= b and not a;
    layer3_outputs(5075) <= not b;
    layer3_outputs(5076) <= not (a or b);
    layer3_outputs(5077) <= not a or b;
    layer3_outputs(5078) <= a or b;
    layer3_outputs(5079) <= not a or b;
    layer3_outputs(5080) <= not (a xor b);
    layer3_outputs(5081) <= not (a and b);
    layer3_outputs(5082) <= not (a and b);
    layer3_outputs(5083) <= a or b;
    layer3_outputs(5084) <= not a or b;
    layer3_outputs(5085) <= b;
    layer3_outputs(5086) <= b;
    layer3_outputs(5087) <= not (a xor b);
    layer3_outputs(5088) <= b and not a;
    layer3_outputs(5089) <= '1';
    layer3_outputs(5090) <= not a or b;
    layer3_outputs(5091) <= '0';
    layer3_outputs(5092) <= a and b;
    layer3_outputs(5093) <= a and b;
    layer3_outputs(5094) <= not (a or b);
    layer3_outputs(5095) <= not (a or b);
    layer3_outputs(5096) <= not a or b;
    layer3_outputs(5097) <= b;
    layer3_outputs(5098) <= a or b;
    layer3_outputs(5099) <= b and not a;
    layer3_outputs(5100) <= a xor b;
    layer3_outputs(5101) <= a xor b;
    layer3_outputs(5102) <= a and not b;
    layer3_outputs(5103) <= not b;
    layer3_outputs(5104) <= not (a and b);
    layer3_outputs(5105) <= not a;
    layer3_outputs(5106) <= b;
    layer3_outputs(5107) <= not a;
    layer3_outputs(5108) <= a and b;
    layer3_outputs(5109) <= '0';
    layer3_outputs(5110) <= a;
    layer3_outputs(5111) <= not b;
    layer3_outputs(5112) <= a xor b;
    layer3_outputs(5113) <= b and not a;
    layer3_outputs(5114) <= not (a and b);
    layer3_outputs(5115) <= not (a or b);
    layer3_outputs(5116) <= a;
    layer3_outputs(5117) <= not (a or b);
    layer3_outputs(5118) <= b and not a;
    layer3_outputs(5119) <= a and not b;
    layer3_outputs(5120) <= a xor b;
    layer3_outputs(5121) <= a and not b;
    layer3_outputs(5122) <= not b or a;
    layer3_outputs(5123) <= a;
    layer3_outputs(5124) <= a or b;
    layer3_outputs(5125) <= b and not a;
    layer3_outputs(5126) <= not a;
    layer3_outputs(5127) <= a and b;
    layer3_outputs(5128) <= not a;
    layer3_outputs(5129) <= not b;
    layer3_outputs(5130) <= not a;
    layer3_outputs(5131) <= not (a or b);
    layer3_outputs(5132) <= a and not b;
    layer3_outputs(5133) <= not b or a;
    layer3_outputs(5134) <= not a;
    layer3_outputs(5135) <= a;
    layer3_outputs(5136) <= a;
    layer3_outputs(5137) <= b;
    layer3_outputs(5138) <= a and b;
    layer3_outputs(5139) <= not (a or b);
    layer3_outputs(5140) <= b;
    layer3_outputs(5141) <= not a;
    layer3_outputs(5142) <= b;
    layer3_outputs(5143) <= b and not a;
    layer3_outputs(5144) <= b;
    layer3_outputs(5145) <= b;
    layer3_outputs(5146) <= not b or a;
    layer3_outputs(5147) <= not (a and b);
    layer3_outputs(5148) <= not a;
    layer3_outputs(5149) <= not a;
    layer3_outputs(5150) <= a and not b;
    layer3_outputs(5151) <= a;
    layer3_outputs(5152) <= not a or b;
    layer3_outputs(5153) <= not (a and b);
    layer3_outputs(5154) <= not (a and b);
    layer3_outputs(5155) <= a;
    layer3_outputs(5156) <= a xor b;
    layer3_outputs(5157) <= '1';
    layer3_outputs(5158) <= not a or b;
    layer3_outputs(5159) <= a xor b;
    layer3_outputs(5160) <= b;
    layer3_outputs(5161) <= b;
    layer3_outputs(5162) <= not (a and b);
    layer3_outputs(5163) <= not a or b;
    layer3_outputs(5164) <= a;
    layer3_outputs(5165) <= not b or a;
    layer3_outputs(5166) <= a or b;
    layer3_outputs(5167) <= a or b;
    layer3_outputs(5168) <= not (a xor b);
    layer3_outputs(5169) <= not b;
    layer3_outputs(5170) <= a and not b;
    layer3_outputs(5171) <= not (a or b);
    layer3_outputs(5172) <= a and not b;
    layer3_outputs(5173) <= a xor b;
    layer3_outputs(5174) <= not (a xor b);
    layer3_outputs(5175) <= a xor b;
    layer3_outputs(5176) <= not (a xor b);
    layer3_outputs(5177) <= b;
    layer3_outputs(5178) <= not a or b;
    layer3_outputs(5179) <= b;
    layer3_outputs(5180) <= not a;
    layer3_outputs(5181) <= a and b;
    layer3_outputs(5182) <= a;
    layer3_outputs(5183) <= not (a or b);
    layer3_outputs(5184) <= not b;
    layer3_outputs(5185) <= b and not a;
    layer3_outputs(5186) <= a and not b;
    layer3_outputs(5187) <= a xor b;
    layer3_outputs(5188) <= a and b;
    layer3_outputs(5189) <= a or b;
    layer3_outputs(5190) <= not a or b;
    layer3_outputs(5191) <= not (a or b);
    layer3_outputs(5192) <= a;
    layer3_outputs(5193) <= not (a and b);
    layer3_outputs(5194) <= b;
    layer3_outputs(5195) <= not a or b;
    layer3_outputs(5196) <= not b;
    layer3_outputs(5197) <= b;
    layer3_outputs(5198) <= a or b;
    layer3_outputs(5199) <= not b or a;
    layer3_outputs(5200) <= not (a xor b);
    layer3_outputs(5201) <= b;
    layer3_outputs(5202) <= not (a and b);
    layer3_outputs(5203) <= not a;
    layer3_outputs(5204) <= a or b;
    layer3_outputs(5205) <= b and not a;
    layer3_outputs(5206) <= a;
    layer3_outputs(5207) <= not a;
    layer3_outputs(5208) <= '0';
    layer3_outputs(5209) <= a xor b;
    layer3_outputs(5210) <= '0';
    layer3_outputs(5211) <= a;
    layer3_outputs(5212) <= not b;
    layer3_outputs(5213) <= '0';
    layer3_outputs(5214) <= a and b;
    layer3_outputs(5215) <= not b;
    layer3_outputs(5216) <= not b;
    layer3_outputs(5217) <= not (a or b);
    layer3_outputs(5218) <= not (a or b);
    layer3_outputs(5219) <= not b or a;
    layer3_outputs(5220) <= not (a or b);
    layer3_outputs(5221) <= not a;
    layer3_outputs(5222) <= not b or a;
    layer3_outputs(5223) <= a or b;
    layer3_outputs(5224) <= b;
    layer3_outputs(5225) <= not (a and b);
    layer3_outputs(5226) <= a;
    layer3_outputs(5227) <= not a;
    layer3_outputs(5228) <= not b;
    layer3_outputs(5229) <= a or b;
    layer3_outputs(5230) <= not (a or b);
    layer3_outputs(5231) <= not a;
    layer3_outputs(5232) <= a xor b;
    layer3_outputs(5233) <= a;
    layer3_outputs(5234) <= not (a and b);
    layer3_outputs(5235) <= a or b;
    layer3_outputs(5236) <= not a or b;
    layer3_outputs(5237) <= b and not a;
    layer3_outputs(5238) <= not (a and b);
    layer3_outputs(5239) <= b and not a;
    layer3_outputs(5240) <= not (a or b);
    layer3_outputs(5241) <= a and b;
    layer3_outputs(5242) <= not a or b;
    layer3_outputs(5243) <= a xor b;
    layer3_outputs(5244) <= b and not a;
    layer3_outputs(5245) <= not (a or b);
    layer3_outputs(5246) <= not (a xor b);
    layer3_outputs(5247) <= a and b;
    layer3_outputs(5248) <= a or b;
    layer3_outputs(5249) <= b and not a;
    layer3_outputs(5250) <= a;
    layer3_outputs(5251) <= not b or a;
    layer3_outputs(5252) <= a xor b;
    layer3_outputs(5253) <= a or b;
    layer3_outputs(5254) <= not b;
    layer3_outputs(5255) <= not a;
    layer3_outputs(5256) <= not a;
    layer3_outputs(5257) <= '0';
    layer3_outputs(5258) <= b;
    layer3_outputs(5259) <= b and not a;
    layer3_outputs(5260) <= a or b;
    layer3_outputs(5261) <= a;
    layer3_outputs(5262) <= not a;
    layer3_outputs(5263) <= not b;
    layer3_outputs(5264) <= a;
    layer3_outputs(5265) <= not a;
    layer3_outputs(5266) <= '1';
    layer3_outputs(5267) <= a xor b;
    layer3_outputs(5268) <= not a;
    layer3_outputs(5269) <= not b;
    layer3_outputs(5270) <= not a;
    layer3_outputs(5271) <= not b or a;
    layer3_outputs(5272) <= not (a or b);
    layer3_outputs(5273) <= b and not a;
    layer3_outputs(5274) <= '0';
    layer3_outputs(5275) <= not (a or b);
    layer3_outputs(5276) <= a or b;
    layer3_outputs(5277) <= a and b;
    layer3_outputs(5278) <= a xor b;
    layer3_outputs(5279) <= not a;
    layer3_outputs(5280) <= not b;
    layer3_outputs(5281) <= '0';
    layer3_outputs(5282) <= a and not b;
    layer3_outputs(5283) <= '0';
    layer3_outputs(5284) <= not (a or b);
    layer3_outputs(5285) <= a or b;
    layer3_outputs(5286) <= a and b;
    layer3_outputs(5287) <= a and b;
    layer3_outputs(5288) <= a and b;
    layer3_outputs(5289) <= a and b;
    layer3_outputs(5290) <= not a;
    layer3_outputs(5291) <= not a;
    layer3_outputs(5292) <= a or b;
    layer3_outputs(5293) <= not a;
    layer3_outputs(5294) <= b;
    layer3_outputs(5295) <= '1';
    layer3_outputs(5296) <= a and b;
    layer3_outputs(5297) <= a xor b;
    layer3_outputs(5298) <= not (a xor b);
    layer3_outputs(5299) <= not b;
    layer3_outputs(5300) <= a or b;
    layer3_outputs(5301) <= b and not a;
    layer3_outputs(5302) <= not b;
    layer3_outputs(5303) <= b;
    layer3_outputs(5304) <= not a or b;
    layer3_outputs(5305) <= not a or b;
    layer3_outputs(5306) <= not a or b;
    layer3_outputs(5307) <= not (a and b);
    layer3_outputs(5308) <= not a or b;
    layer3_outputs(5309) <= a;
    layer3_outputs(5310) <= not b or a;
    layer3_outputs(5311) <= a and not b;
    layer3_outputs(5312) <= a xor b;
    layer3_outputs(5313) <= b;
    layer3_outputs(5314) <= a and b;
    layer3_outputs(5315) <= a or b;
    layer3_outputs(5316) <= not b;
    layer3_outputs(5317) <= not a;
    layer3_outputs(5318) <= a and not b;
    layer3_outputs(5319) <= not b;
    layer3_outputs(5320) <= not b or a;
    layer3_outputs(5321) <= not (a or b);
    layer3_outputs(5322) <= a or b;
    layer3_outputs(5323) <= not a or b;
    layer3_outputs(5324) <= '0';
    layer3_outputs(5325) <= not (a and b);
    layer3_outputs(5326) <= not a;
    layer3_outputs(5327) <= not a;
    layer3_outputs(5328) <= a;
    layer3_outputs(5329) <= b;
    layer3_outputs(5330) <= a and b;
    layer3_outputs(5331) <= b;
    layer3_outputs(5332) <= a;
    layer3_outputs(5333) <= not b;
    layer3_outputs(5334) <= b;
    layer3_outputs(5335) <= a and not b;
    layer3_outputs(5336) <= not (a or b);
    layer3_outputs(5337) <= b and not a;
    layer3_outputs(5338) <= a xor b;
    layer3_outputs(5339) <= not (a and b);
    layer3_outputs(5340) <= not b or a;
    layer3_outputs(5341) <= not b or a;
    layer3_outputs(5342) <= a and not b;
    layer3_outputs(5343) <= a and b;
    layer3_outputs(5344) <= b and not a;
    layer3_outputs(5345) <= not b;
    layer3_outputs(5346) <= a;
    layer3_outputs(5347) <= b;
    layer3_outputs(5348) <= a or b;
    layer3_outputs(5349) <= not a or b;
    layer3_outputs(5350) <= not b or a;
    layer3_outputs(5351) <= a and not b;
    layer3_outputs(5352) <= a xor b;
    layer3_outputs(5353) <= '0';
    layer3_outputs(5354) <= b and not a;
    layer3_outputs(5355) <= a and not b;
    layer3_outputs(5356) <= not b;
    layer3_outputs(5357) <= b and not a;
    layer3_outputs(5358) <= not a;
    layer3_outputs(5359) <= not (a and b);
    layer3_outputs(5360) <= a;
    layer3_outputs(5361) <= not b or a;
    layer3_outputs(5362) <= '0';
    layer3_outputs(5363) <= '0';
    layer3_outputs(5364) <= a or b;
    layer3_outputs(5365) <= b;
    layer3_outputs(5366) <= not b;
    layer3_outputs(5367) <= a;
    layer3_outputs(5368) <= not a;
    layer3_outputs(5369) <= not b;
    layer3_outputs(5370) <= a and not b;
    layer3_outputs(5371) <= b and not a;
    layer3_outputs(5372) <= not a;
    layer3_outputs(5373) <= not a;
    layer3_outputs(5374) <= not a or b;
    layer3_outputs(5375) <= not b or a;
    layer3_outputs(5376) <= b and not a;
    layer3_outputs(5377) <= not a or b;
    layer3_outputs(5378) <= not b or a;
    layer3_outputs(5379) <= a or b;
    layer3_outputs(5380) <= a;
    layer3_outputs(5381) <= not (a or b);
    layer3_outputs(5382) <= not a;
    layer3_outputs(5383) <= b;
    layer3_outputs(5384) <= a and b;
    layer3_outputs(5385) <= b;
    layer3_outputs(5386) <= b;
    layer3_outputs(5387) <= not b;
    layer3_outputs(5388) <= b;
    layer3_outputs(5389) <= a and b;
    layer3_outputs(5390) <= not (a xor b);
    layer3_outputs(5391) <= b and not a;
    layer3_outputs(5392) <= not (a xor b);
    layer3_outputs(5393) <= not b or a;
    layer3_outputs(5394) <= not b;
    layer3_outputs(5395) <= a or b;
    layer3_outputs(5396) <= not b;
    layer3_outputs(5397) <= b and not a;
    layer3_outputs(5398) <= a;
    layer3_outputs(5399) <= b;
    layer3_outputs(5400) <= a or b;
    layer3_outputs(5401) <= b;
    layer3_outputs(5402) <= not a;
    layer3_outputs(5403) <= a or b;
    layer3_outputs(5404) <= a or b;
    layer3_outputs(5405) <= a and b;
    layer3_outputs(5406) <= not b;
    layer3_outputs(5407) <= a;
    layer3_outputs(5408) <= a;
    layer3_outputs(5409) <= not a;
    layer3_outputs(5410) <= not a;
    layer3_outputs(5411) <= not (a xor b);
    layer3_outputs(5412) <= '0';
    layer3_outputs(5413) <= not b;
    layer3_outputs(5414) <= not (a and b);
    layer3_outputs(5415) <= not a;
    layer3_outputs(5416) <= a or b;
    layer3_outputs(5417) <= a and not b;
    layer3_outputs(5418) <= not b or a;
    layer3_outputs(5419) <= a and b;
    layer3_outputs(5420) <= a xor b;
    layer3_outputs(5421) <= not a;
    layer3_outputs(5422) <= b;
    layer3_outputs(5423) <= not (a and b);
    layer3_outputs(5424) <= not (a xor b);
    layer3_outputs(5425) <= not (a or b);
    layer3_outputs(5426) <= a and not b;
    layer3_outputs(5427) <= b and not a;
    layer3_outputs(5428) <= a xor b;
    layer3_outputs(5429) <= not a;
    layer3_outputs(5430) <= a or b;
    layer3_outputs(5431) <= '0';
    layer3_outputs(5432) <= '0';
    layer3_outputs(5433) <= a;
    layer3_outputs(5434) <= a and b;
    layer3_outputs(5435) <= a xor b;
    layer3_outputs(5436) <= a;
    layer3_outputs(5437) <= a;
    layer3_outputs(5438) <= '0';
    layer3_outputs(5439) <= not (a or b);
    layer3_outputs(5440) <= b and not a;
    layer3_outputs(5441) <= not b;
    layer3_outputs(5442) <= a and b;
    layer3_outputs(5443) <= not (a and b);
    layer3_outputs(5444) <= a xor b;
    layer3_outputs(5445) <= a;
    layer3_outputs(5446) <= not b or a;
    layer3_outputs(5447) <= not (a or b);
    layer3_outputs(5448) <= b and not a;
    layer3_outputs(5449) <= not (a xor b);
    layer3_outputs(5450) <= a;
    layer3_outputs(5451) <= '0';
    layer3_outputs(5452) <= not a or b;
    layer3_outputs(5453) <= a or b;
    layer3_outputs(5454) <= not (a and b);
    layer3_outputs(5455) <= b;
    layer3_outputs(5456) <= not a or b;
    layer3_outputs(5457) <= a and b;
    layer3_outputs(5458) <= a;
    layer3_outputs(5459) <= not b;
    layer3_outputs(5460) <= not (a or b);
    layer3_outputs(5461) <= not a or b;
    layer3_outputs(5462) <= not a;
    layer3_outputs(5463) <= b and not a;
    layer3_outputs(5464) <= not (a or b);
    layer3_outputs(5465) <= not a;
    layer3_outputs(5466) <= not b or a;
    layer3_outputs(5467) <= '1';
    layer3_outputs(5468) <= not b;
    layer3_outputs(5469) <= a and not b;
    layer3_outputs(5470) <= a and b;
    layer3_outputs(5471) <= a or b;
    layer3_outputs(5472) <= a and b;
    layer3_outputs(5473) <= not a or b;
    layer3_outputs(5474) <= not b;
    layer3_outputs(5475) <= a and not b;
    layer3_outputs(5476) <= b;
    layer3_outputs(5477) <= not a;
    layer3_outputs(5478) <= not b or a;
    layer3_outputs(5479) <= not a;
    layer3_outputs(5480) <= not a or b;
    layer3_outputs(5481) <= a and not b;
    layer3_outputs(5482) <= b and not a;
    layer3_outputs(5483) <= a and b;
    layer3_outputs(5484) <= not b or a;
    layer3_outputs(5485) <= not b or a;
    layer3_outputs(5486) <= not b or a;
    layer3_outputs(5487) <= not b;
    layer3_outputs(5488) <= a or b;
    layer3_outputs(5489) <= not b or a;
    layer3_outputs(5490) <= not a;
    layer3_outputs(5491) <= not a;
    layer3_outputs(5492) <= not (a and b);
    layer3_outputs(5493) <= b;
    layer3_outputs(5494) <= not a;
    layer3_outputs(5495) <= not (a and b);
    layer3_outputs(5496) <= b and not a;
    layer3_outputs(5497) <= a;
    layer3_outputs(5498) <= not a or b;
    layer3_outputs(5499) <= not (a and b);
    layer3_outputs(5500) <= b and not a;
    layer3_outputs(5501) <= a;
    layer3_outputs(5502) <= not (a and b);
    layer3_outputs(5503) <= not a;
    layer3_outputs(5504) <= a and b;
    layer3_outputs(5505) <= a or b;
    layer3_outputs(5506) <= b;
    layer3_outputs(5507) <= a;
    layer3_outputs(5508) <= not (a and b);
    layer3_outputs(5509) <= '1';
    layer3_outputs(5510) <= not (a or b);
    layer3_outputs(5511) <= not b;
    layer3_outputs(5512) <= a and b;
    layer3_outputs(5513) <= not a;
    layer3_outputs(5514) <= not b;
    layer3_outputs(5515) <= not b;
    layer3_outputs(5516) <= not b;
    layer3_outputs(5517) <= not a or b;
    layer3_outputs(5518) <= b;
    layer3_outputs(5519) <= not (a or b);
    layer3_outputs(5520) <= not (a xor b);
    layer3_outputs(5521) <= a and b;
    layer3_outputs(5522) <= not b or a;
    layer3_outputs(5523) <= a xor b;
    layer3_outputs(5524) <= not (a and b);
    layer3_outputs(5525) <= '0';
    layer3_outputs(5526) <= not (a or b);
    layer3_outputs(5527) <= a or b;
    layer3_outputs(5528) <= a xor b;
    layer3_outputs(5529) <= not b;
    layer3_outputs(5530) <= a and b;
    layer3_outputs(5531) <= not a;
    layer3_outputs(5532) <= not (a and b);
    layer3_outputs(5533) <= not (a xor b);
    layer3_outputs(5534) <= a xor b;
    layer3_outputs(5535) <= a and b;
    layer3_outputs(5536) <= b;
    layer3_outputs(5537) <= a xor b;
    layer3_outputs(5538) <= '1';
    layer3_outputs(5539) <= not b;
    layer3_outputs(5540) <= not a or b;
    layer3_outputs(5541) <= a and b;
    layer3_outputs(5542) <= '0';
    layer3_outputs(5543) <= '0';
    layer3_outputs(5544) <= not (a and b);
    layer3_outputs(5545) <= not (a or b);
    layer3_outputs(5546) <= not b or a;
    layer3_outputs(5547) <= a and b;
    layer3_outputs(5548) <= not (a or b);
    layer3_outputs(5549) <= b and not a;
    layer3_outputs(5550) <= a xor b;
    layer3_outputs(5551) <= '0';
    layer3_outputs(5552) <= a xor b;
    layer3_outputs(5553) <= b and not a;
    layer3_outputs(5554) <= a;
    layer3_outputs(5555) <= not (a xor b);
    layer3_outputs(5556) <= a xor b;
    layer3_outputs(5557) <= not b;
    layer3_outputs(5558) <= a or b;
    layer3_outputs(5559) <= not (a and b);
    layer3_outputs(5560) <= not a;
    layer3_outputs(5561) <= '1';
    layer3_outputs(5562) <= not a;
    layer3_outputs(5563) <= a and b;
    layer3_outputs(5564) <= a or b;
    layer3_outputs(5565) <= a;
    layer3_outputs(5566) <= '1';
    layer3_outputs(5567) <= not (a or b);
    layer3_outputs(5568) <= a xor b;
    layer3_outputs(5569) <= not a;
    layer3_outputs(5570) <= a xor b;
    layer3_outputs(5571) <= b;
    layer3_outputs(5572) <= not b or a;
    layer3_outputs(5573) <= b;
    layer3_outputs(5574) <= not b;
    layer3_outputs(5575) <= b;
    layer3_outputs(5576) <= not b;
    layer3_outputs(5577) <= not b or a;
    layer3_outputs(5578) <= b;
    layer3_outputs(5579) <= b and not a;
    layer3_outputs(5580) <= b;
    layer3_outputs(5581) <= a;
    layer3_outputs(5582) <= a;
    layer3_outputs(5583) <= not (a and b);
    layer3_outputs(5584) <= not (a xor b);
    layer3_outputs(5585) <= a and not b;
    layer3_outputs(5586) <= '0';
    layer3_outputs(5587) <= not (a and b);
    layer3_outputs(5588) <= a and b;
    layer3_outputs(5589) <= a and not b;
    layer3_outputs(5590) <= a;
    layer3_outputs(5591) <= a xor b;
    layer3_outputs(5592) <= not a;
    layer3_outputs(5593) <= '0';
    layer3_outputs(5594) <= a and b;
    layer3_outputs(5595) <= a and b;
    layer3_outputs(5596) <= a or b;
    layer3_outputs(5597) <= a and b;
    layer3_outputs(5598) <= b and not a;
    layer3_outputs(5599) <= a and not b;
    layer3_outputs(5600) <= not a;
    layer3_outputs(5601) <= a and b;
    layer3_outputs(5602) <= not b or a;
    layer3_outputs(5603) <= b and not a;
    layer3_outputs(5604) <= not (a or b);
    layer3_outputs(5605) <= a;
    layer3_outputs(5606) <= a or b;
    layer3_outputs(5607) <= a or b;
    layer3_outputs(5608) <= '1';
    layer3_outputs(5609) <= a or b;
    layer3_outputs(5610) <= not a or b;
    layer3_outputs(5611) <= a xor b;
    layer3_outputs(5612) <= a;
    layer3_outputs(5613) <= b and not a;
    layer3_outputs(5614) <= a or b;
    layer3_outputs(5615) <= '1';
    layer3_outputs(5616) <= not a or b;
    layer3_outputs(5617) <= b and not a;
    layer3_outputs(5618) <= a and not b;
    layer3_outputs(5619) <= '1';
    layer3_outputs(5620) <= not b;
    layer3_outputs(5621) <= not b;
    layer3_outputs(5622) <= b;
    layer3_outputs(5623) <= '1';
    layer3_outputs(5624) <= not b;
    layer3_outputs(5625) <= '1';
    layer3_outputs(5626) <= not a;
    layer3_outputs(5627) <= not b;
    layer3_outputs(5628) <= '0';
    layer3_outputs(5629) <= a and not b;
    layer3_outputs(5630) <= not (a and b);
    layer3_outputs(5631) <= not a;
    layer3_outputs(5632) <= not (a and b);
    layer3_outputs(5633) <= not a;
    layer3_outputs(5634) <= '1';
    layer3_outputs(5635) <= not a;
    layer3_outputs(5636) <= not (a or b);
    layer3_outputs(5637) <= not a;
    layer3_outputs(5638) <= not a or b;
    layer3_outputs(5639) <= '0';
    layer3_outputs(5640) <= b and not a;
    layer3_outputs(5641) <= not b;
    layer3_outputs(5642) <= a or b;
    layer3_outputs(5643) <= b;
    layer3_outputs(5644) <= a and b;
    layer3_outputs(5645) <= a xor b;
    layer3_outputs(5646) <= a;
    layer3_outputs(5647) <= not b;
    layer3_outputs(5648) <= a and b;
    layer3_outputs(5649) <= not (a or b);
    layer3_outputs(5650) <= a;
    layer3_outputs(5651) <= a and b;
    layer3_outputs(5652) <= '0';
    layer3_outputs(5653) <= a or b;
    layer3_outputs(5654) <= '1';
    layer3_outputs(5655) <= not a;
    layer3_outputs(5656) <= not (a or b);
    layer3_outputs(5657) <= not (a xor b);
    layer3_outputs(5658) <= a and b;
    layer3_outputs(5659) <= b;
    layer3_outputs(5660) <= not (a or b);
    layer3_outputs(5661) <= not b or a;
    layer3_outputs(5662) <= a xor b;
    layer3_outputs(5663) <= a or b;
    layer3_outputs(5664) <= a xor b;
    layer3_outputs(5665) <= not (a xor b);
    layer3_outputs(5666) <= a and not b;
    layer3_outputs(5667) <= '1';
    layer3_outputs(5668) <= a;
    layer3_outputs(5669) <= not (a xor b);
    layer3_outputs(5670) <= b;
    layer3_outputs(5671) <= not a or b;
    layer3_outputs(5672) <= '0';
    layer3_outputs(5673) <= a and not b;
    layer3_outputs(5674) <= not (a and b);
    layer3_outputs(5675) <= not a or b;
    layer3_outputs(5676) <= a and b;
    layer3_outputs(5677) <= not (a or b);
    layer3_outputs(5678) <= not (a and b);
    layer3_outputs(5679) <= not b;
    layer3_outputs(5680) <= a and b;
    layer3_outputs(5681) <= '0';
    layer3_outputs(5682) <= not b;
    layer3_outputs(5683) <= not b;
    layer3_outputs(5684) <= a and b;
    layer3_outputs(5685) <= a and not b;
    layer3_outputs(5686) <= not (a and b);
    layer3_outputs(5687) <= not a or b;
    layer3_outputs(5688) <= not (a or b);
    layer3_outputs(5689) <= not b;
    layer3_outputs(5690) <= not a or b;
    layer3_outputs(5691) <= not (a xor b);
    layer3_outputs(5692) <= not (a and b);
    layer3_outputs(5693) <= not b;
    layer3_outputs(5694) <= b;
    layer3_outputs(5695) <= a and not b;
    layer3_outputs(5696) <= not a or b;
    layer3_outputs(5697) <= not (a or b);
    layer3_outputs(5698) <= not (a xor b);
    layer3_outputs(5699) <= b;
    layer3_outputs(5700) <= '0';
    layer3_outputs(5701) <= a and not b;
    layer3_outputs(5702) <= a and b;
    layer3_outputs(5703) <= not (a or b);
    layer3_outputs(5704) <= b and not a;
    layer3_outputs(5705) <= a and not b;
    layer3_outputs(5706) <= not (a and b);
    layer3_outputs(5707) <= not a;
    layer3_outputs(5708) <= not b;
    layer3_outputs(5709) <= a;
    layer3_outputs(5710) <= not (a and b);
    layer3_outputs(5711) <= b;
    layer3_outputs(5712) <= b;
    layer3_outputs(5713) <= a and not b;
    layer3_outputs(5714) <= a xor b;
    layer3_outputs(5715) <= a;
    layer3_outputs(5716) <= a xor b;
    layer3_outputs(5717) <= a;
    layer3_outputs(5718) <= a and b;
    layer3_outputs(5719) <= b;
    layer3_outputs(5720) <= not a;
    layer3_outputs(5721) <= not (a or b);
    layer3_outputs(5722) <= b;
    layer3_outputs(5723) <= b and not a;
    layer3_outputs(5724) <= not a;
    layer3_outputs(5725) <= not (a xor b);
    layer3_outputs(5726) <= not b;
    layer3_outputs(5727) <= a;
    layer3_outputs(5728) <= b;
    layer3_outputs(5729) <= not a or b;
    layer3_outputs(5730) <= not b or a;
    layer3_outputs(5731) <= b and not a;
    layer3_outputs(5732) <= not a or b;
    layer3_outputs(5733) <= not a;
    layer3_outputs(5734) <= a or b;
    layer3_outputs(5735) <= not b;
    layer3_outputs(5736) <= not (a or b);
    layer3_outputs(5737) <= a or b;
    layer3_outputs(5738) <= not b or a;
    layer3_outputs(5739) <= not b;
    layer3_outputs(5740) <= not (a and b);
    layer3_outputs(5741) <= not (a xor b);
    layer3_outputs(5742) <= b;
    layer3_outputs(5743) <= not b or a;
    layer3_outputs(5744) <= a and b;
    layer3_outputs(5745) <= not a or b;
    layer3_outputs(5746) <= b;
    layer3_outputs(5747) <= '0';
    layer3_outputs(5748) <= not (a or b);
    layer3_outputs(5749) <= not b or a;
    layer3_outputs(5750) <= a or b;
    layer3_outputs(5751) <= '1';
    layer3_outputs(5752) <= a or b;
    layer3_outputs(5753) <= a and not b;
    layer3_outputs(5754) <= b;
    layer3_outputs(5755) <= not (a xor b);
    layer3_outputs(5756) <= not (a and b);
    layer3_outputs(5757) <= not b;
    layer3_outputs(5758) <= b;
    layer3_outputs(5759) <= b and not a;
    layer3_outputs(5760) <= not (a xor b);
    layer3_outputs(5761) <= not b;
    layer3_outputs(5762) <= '1';
    layer3_outputs(5763) <= b;
    layer3_outputs(5764) <= not a;
    layer3_outputs(5765) <= a and b;
    layer3_outputs(5766) <= b;
    layer3_outputs(5767) <= not b;
    layer3_outputs(5768) <= b;
    layer3_outputs(5769) <= not b;
    layer3_outputs(5770) <= a and b;
    layer3_outputs(5771) <= a;
    layer3_outputs(5772) <= not b or a;
    layer3_outputs(5773) <= b;
    layer3_outputs(5774) <= a;
    layer3_outputs(5775) <= '1';
    layer3_outputs(5776) <= not (a and b);
    layer3_outputs(5777) <= not (a and b);
    layer3_outputs(5778) <= not (a and b);
    layer3_outputs(5779) <= not b or a;
    layer3_outputs(5780) <= b;
    layer3_outputs(5781) <= '1';
    layer3_outputs(5782) <= b;
    layer3_outputs(5783) <= not a;
    layer3_outputs(5784) <= not a or b;
    layer3_outputs(5785) <= not (a and b);
    layer3_outputs(5786) <= not b or a;
    layer3_outputs(5787) <= not (a or b);
    layer3_outputs(5788) <= b and not a;
    layer3_outputs(5789) <= not a or b;
    layer3_outputs(5790) <= not a;
    layer3_outputs(5791) <= '0';
    layer3_outputs(5792) <= b and not a;
    layer3_outputs(5793) <= not a;
    layer3_outputs(5794) <= not b or a;
    layer3_outputs(5795) <= a xor b;
    layer3_outputs(5796) <= not (a or b);
    layer3_outputs(5797) <= not (a or b);
    layer3_outputs(5798) <= b;
    layer3_outputs(5799) <= a or b;
    layer3_outputs(5800) <= '0';
    layer3_outputs(5801) <= a and not b;
    layer3_outputs(5802) <= a or b;
    layer3_outputs(5803) <= b;
    layer3_outputs(5804) <= a;
    layer3_outputs(5805) <= not (a and b);
    layer3_outputs(5806) <= a or b;
    layer3_outputs(5807) <= b and not a;
    layer3_outputs(5808) <= a and b;
    layer3_outputs(5809) <= a and b;
    layer3_outputs(5810) <= not a or b;
    layer3_outputs(5811) <= not (a or b);
    layer3_outputs(5812) <= a and b;
    layer3_outputs(5813) <= not a;
    layer3_outputs(5814) <= a and b;
    layer3_outputs(5815) <= a or b;
    layer3_outputs(5816) <= b;
    layer3_outputs(5817) <= b and not a;
    layer3_outputs(5818) <= a xor b;
    layer3_outputs(5819) <= not (a and b);
    layer3_outputs(5820) <= not a;
    layer3_outputs(5821) <= not (a xor b);
    layer3_outputs(5822) <= not b;
    layer3_outputs(5823) <= a and not b;
    layer3_outputs(5824) <= a;
    layer3_outputs(5825) <= not a;
    layer3_outputs(5826) <= not b;
    layer3_outputs(5827) <= not (a or b);
    layer3_outputs(5828) <= a and not b;
    layer3_outputs(5829) <= not b or a;
    layer3_outputs(5830) <= not a;
    layer3_outputs(5831) <= not a;
    layer3_outputs(5832) <= a and not b;
    layer3_outputs(5833) <= a and not b;
    layer3_outputs(5834) <= not b;
    layer3_outputs(5835) <= not (a and b);
    layer3_outputs(5836) <= '1';
    layer3_outputs(5837) <= a;
    layer3_outputs(5838) <= b;
    layer3_outputs(5839) <= not (a and b);
    layer3_outputs(5840) <= a or b;
    layer3_outputs(5841) <= a and b;
    layer3_outputs(5842) <= a;
    layer3_outputs(5843) <= a and b;
    layer3_outputs(5844) <= a;
    layer3_outputs(5845) <= a and not b;
    layer3_outputs(5846) <= not (a xor b);
    layer3_outputs(5847) <= b;
    layer3_outputs(5848) <= not a or b;
    layer3_outputs(5849) <= not b;
    layer3_outputs(5850) <= b and not a;
    layer3_outputs(5851) <= a and b;
    layer3_outputs(5852) <= a;
    layer3_outputs(5853) <= b and not a;
    layer3_outputs(5854) <= a and b;
    layer3_outputs(5855) <= not a;
    layer3_outputs(5856) <= not (a or b);
    layer3_outputs(5857) <= a or b;
    layer3_outputs(5858) <= b;
    layer3_outputs(5859) <= b;
    layer3_outputs(5860) <= not b or a;
    layer3_outputs(5861) <= not a;
    layer3_outputs(5862) <= not a;
    layer3_outputs(5863) <= '0';
    layer3_outputs(5864) <= a and not b;
    layer3_outputs(5865) <= b;
    layer3_outputs(5866) <= '1';
    layer3_outputs(5867) <= not b;
    layer3_outputs(5868) <= a and b;
    layer3_outputs(5869) <= a and not b;
    layer3_outputs(5870) <= not a;
    layer3_outputs(5871) <= not (a and b);
    layer3_outputs(5872) <= a;
    layer3_outputs(5873) <= not a;
    layer3_outputs(5874) <= '1';
    layer3_outputs(5875) <= b and not a;
    layer3_outputs(5876) <= not b or a;
    layer3_outputs(5877) <= a and not b;
    layer3_outputs(5878) <= b;
    layer3_outputs(5879) <= a or b;
    layer3_outputs(5880) <= not b;
    layer3_outputs(5881) <= not a or b;
    layer3_outputs(5882) <= not (a xor b);
    layer3_outputs(5883) <= b;
    layer3_outputs(5884) <= a;
    layer3_outputs(5885) <= '0';
    layer3_outputs(5886) <= not b or a;
    layer3_outputs(5887) <= b;
    layer3_outputs(5888) <= a and not b;
    layer3_outputs(5889) <= b and not a;
    layer3_outputs(5890) <= b;
    layer3_outputs(5891) <= '0';
    layer3_outputs(5892) <= not b;
    layer3_outputs(5893) <= b and not a;
    layer3_outputs(5894) <= a and not b;
    layer3_outputs(5895) <= not (a and b);
    layer3_outputs(5896) <= b;
    layer3_outputs(5897) <= a and not b;
    layer3_outputs(5898) <= not (a xor b);
    layer3_outputs(5899) <= '0';
    layer3_outputs(5900) <= not (a or b);
    layer3_outputs(5901) <= a;
    layer3_outputs(5902) <= a and not b;
    layer3_outputs(5903) <= not (a xor b);
    layer3_outputs(5904) <= '1';
    layer3_outputs(5905) <= b;
    layer3_outputs(5906) <= a and b;
    layer3_outputs(5907) <= a;
    layer3_outputs(5908) <= a and not b;
    layer3_outputs(5909) <= a;
    layer3_outputs(5910) <= b;
    layer3_outputs(5911) <= not (a or b);
    layer3_outputs(5912) <= not (a and b);
    layer3_outputs(5913) <= not (a xor b);
    layer3_outputs(5914) <= '1';
    layer3_outputs(5915) <= a xor b;
    layer3_outputs(5916) <= a and not b;
    layer3_outputs(5917) <= a;
    layer3_outputs(5918) <= not a;
    layer3_outputs(5919) <= a xor b;
    layer3_outputs(5920) <= not a or b;
    layer3_outputs(5921) <= b;
    layer3_outputs(5922) <= not a;
    layer3_outputs(5923) <= not a or b;
    layer3_outputs(5924) <= not a;
    layer3_outputs(5925) <= b;
    layer3_outputs(5926) <= b and not a;
    layer3_outputs(5927) <= not b or a;
    layer3_outputs(5928) <= a;
    layer3_outputs(5929) <= a;
    layer3_outputs(5930) <= not (a and b);
    layer3_outputs(5931) <= b;
    layer3_outputs(5932) <= a or b;
    layer3_outputs(5933) <= not (a and b);
    layer3_outputs(5934) <= b;
    layer3_outputs(5935) <= not b;
    layer3_outputs(5936) <= not (a xor b);
    layer3_outputs(5937) <= not (a and b);
    layer3_outputs(5938) <= not b;
    layer3_outputs(5939) <= b and not a;
    layer3_outputs(5940) <= a or b;
    layer3_outputs(5941) <= a;
    layer3_outputs(5942) <= not (a and b);
    layer3_outputs(5943) <= b;
    layer3_outputs(5944) <= not b or a;
    layer3_outputs(5945) <= not b or a;
    layer3_outputs(5946) <= b;
    layer3_outputs(5947) <= '1';
    layer3_outputs(5948) <= not (a and b);
    layer3_outputs(5949) <= not (a or b);
    layer3_outputs(5950) <= '1';
    layer3_outputs(5951) <= not a;
    layer3_outputs(5952) <= b and not a;
    layer3_outputs(5953) <= a;
    layer3_outputs(5954) <= not b;
    layer3_outputs(5955) <= b and not a;
    layer3_outputs(5956) <= a and b;
    layer3_outputs(5957) <= not (a or b);
    layer3_outputs(5958) <= not a or b;
    layer3_outputs(5959) <= not a or b;
    layer3_outputs(5960) <= a xor b;
    layer3_outputs(5961) <= not b;
    layer3_outputs(5962) <= '1';
    layer3_outputs(5963) <= not (a and b);
    layer3_outputs(5964) <= a;
    layer3_outputs(5965) <= a or b;
    layer3_outputs(5966) <= '1';
    layer3_outputs(5967) <= not b;
    layer3_outputs(5968) <= not a;
    layer3_outputs(5969) <= '1';
    layer3_outputs(5970) <= not (a and b);
    layer3_outputs(5971) <= '1';
    layer3_outputs(5972) <= '0';
    layer3_outputs(5973) <= not a;
    layer3_outputs(5974) <= a xor b;
    layer3_outputs(5975) <= not (a and b);
    layer3_outputs(5976) <= a and not b;
    layer3_outputs(5977) <= b;
    layer3_outputs(5978) <= not (a and b);
    layer3_outputs(5979) <= not b or a;
    layer3_outputs(5980) <= not (a or b);
    layer3_outputs(5981) <= a or b;
    layer3_outputs(5982) <= not b;
    layer3_outputs(5983) <= not b;
    layer3_outputs(5984) <= b;
    layer3_outputs(5985) <= a;
    layer3_outputs(5986) <= not (a xor b);
    layer3_outputs(5987) <= not a;
    layer3_outputs(5988) <= a and b;
    layer3_outputs(5989) <= not (a and b);
    layer3_outputs(5990) <= a and b;
    layer3_outputs(5991) <= a xor b;
    layer3_outputs(5992) <= not (a or b);
    layer3_outputs(5993) <= not a or b;
    layer3_outputs(5994) <= not a;
    layer3_outputs(5995) <= a;
    layer3_outputs(5996) <= a and b;
    layer3_outputs(5997) <= not (a and b);
    layer3_outputs(5998) <= a or b;
    layer3_outputs(5999) <= '1';
    layer3_outputs(6000) <= not b or a;
    layer3_outputs(6001) <= a and b;
    layer3_outputs(6002) <= not b or a;
    layer3_outputs(6003) <= b;
    layer3_outputs(6004) <= b;
    layer3_outputs(6005) <= a;
    layer3_outputs(6006) <= not b;
    layer3_outputs(6007) <= a and not b;
    layer3_outputs(6008) <= a;
    layer3_outputs(6009) <= a;
    layer3_outputs(6010) <= not a;
    layer3_outputs(6011) <= b;
    layer3_outputs(6012) <= not b;
    layer3_outputs(6013) <= b and not a;
    layer3_outputs(6014) <= b and not a;
    layer3_outputs(6015) <= a or b;
    layer3_outputs(6016) <= not b or a;
    layer3_outputs(6017) <= b;
    layer3_outputs(6018) <= a and not b;
    layer3_outputs(6019) <= '1';
    layer3_outputs(6020) <= '1';
    layer3_outputs(6021) <= b;
    layer3_outputs(6022) <= not b or a;
    layer3_outputs(6023) <= a or b;
    layer3_outputs(6024) <= a and b;
    layer3_outputs(6025) <= not b or a;
    layer3_outputs(6026) <= a xor b;
    layer3_outputs(6027) <= b and not a;
    layer3_outputs(6028) <= not a;
    layer3_outputs(6029) <= not b or a;
    layer3_outputs(6030) <= not (a xor b);
    layer3_outputs(6031) <= not (a and b);
    layer3_outputs(6032) <= not b or a;
    layer3_outputs(6033) <= a xor b;
    layer3_outputs(6034) <= b and not a;
    layer3_outputs(6035) <= not a;
    layer3_outputs(6036) <= b;
    layer3_outputs(6037) <= b;
    layer3_outputs(6038) <= not b;
    layer3_outputs(6039) <= not (a and b);
    layer3_outputs(6040) <= a or b;
    layer3_outputs(6041) <= b;
    layer3_outputs(6042) <= a xor b;
    layer3_outputs(6043) <= not a;
    layer3_outputs(6044) <= b;
    layer3_outputs(6045) <= a and b;
    layer3_outputs(6046) <= not (a and b);
    layer3_outputs(6047) <= a or b;
    layer3_outputs(6048) <= '1';
    layer3_outputs(6049) <= not b;
    layer3_outputs(6050) <= '0';
    layer3_outputs(6051) <= not a;
    layer3_outputs(6052) <= a and b;
    layer3_outputs(6053) <= not (a or b);
    layer3_outputs(6054) <= a or b;
    layer3_outputs(6055) <= a and not b;
    layer3_outputs(6056) <= b;
    layer3_outputs(6057) <= '0';
    layer3_outputs(6058) <= not a;
    layer3_outputs(6059) <= a or b;
    layer3_outputs(6060) <= not (a or b);
    layer3_outputs(6061) <= not (a xor b);
    layer3_outputs(6062) <= not a or b;
    layer3_outputs(6063) <= not b or a;
    layer3_outputs(6064) <= a and not b;
    layer3_outputs(6065) <= a and b;
    layer3_outputs(6066) <= not (a and b);
    layer3_outputs(6067) <= a and b;
    layer3_outputs(6068) <= a and b;
    layer3_outputs(6069) <= b and not a;
    layer3_outputs(6070) <= a and not b;
    layer3_outputs(6071) <= not a or b;
    layer3_outputs(6072) <= b;
    layer3_outputs(6073) <= a;
    layer3_outputs(6074) <= b;
    layer3_outputs(6075) <= not (a or b);
    layer3_outputs(6076) <= not a;
    layer3_outputs(6077) <= b;
    layer3_outputs(6078) <= a or b;
    layer3_outputs(6079) <= not (a or b);
    layer3_outputs(6080) <= not b;
    layer3_outputs(6081) <= not b;
    layer3_outputs(6082) <= b;
    layer3_outputs(6083) <= a;
    layer3_outputs(6084) <= not a;
    layer3_outputs(6085) <= not b or a;
    layer3_outputs(6086) <= b;
    layer3_outputs(6087) <= a;
    layer3_outputs(6088) <= '1';
    layer3_outputs(6089) <= a and b;
    layer3_outputs(6090) <= a and b;
    layer3_outputs(6091) <= b and not a;
    layer3_outputs(6092) <= not (a xor b);
    layer3_outputs(6093) <= not (a or b);
    layer3_outputs(6094) <= not a or b;
    layer3_outputs(6095) <= b;
    layer3_outputs(6096) <= not a or b;
    layer3_outputs(6097) <= '1';
    layer3_outputs(6098) <= a and not b;
    layer3_outputs(6099) <= not (a and b);
    layer3_outputs(6100) <= a;
    layer3_outputs(6101) <= '1';
    layer3_outputs(6102) <= not a;
    layer3_outputs(6103) <= b and not a;
    layer3_outputs(6104) <= not (a and b);
    layer3_outputs(6105) <= a and not b;
    layer3_outputs(6106) <= '1';
    layer3_outputs(6107) <= not a;
    layer3_outputs(6108) <= not a;
    layer3_outputs(6109) <= b;
    layer3_outputs(6110) <= b and not a;
    layer3_outputs(6111) <= b;
    layer3_outputs(6112) <= not b;
    layer3_outputs(6113) <= b;
    layer3_outputs(6114) <= a or b;
    layer3_outputs(6115) <= not b or a;
    layer3_outputs(6116) <= not a;
    layer3_outputs(6117) <= not b;
    layer3_outputs(6118) <= a;
    layer3_outputs(6119) <= a and b;
    layer3_outputs(6120) <= not a or b;
    layer3_outputs(6121) <= not a;
    layer3_outputs(6122) <= a and not b;
    layer3_outputs(6123) <= not (a xor b);
    layer3_outputs(6124) <= not b;
    layer3_outputs(6125) <= a;
    layer3_outputs(6126) <= a and b;
    layer3_outputs(6127) <= a xor b;
    layer3_outputs(6128) <= b and not a;
    layer3_outputs(6129) <= b;
    layer3_outputs(6130) <= '0';
    layer3_outputs(6131) <= not b;
    layer3_outputs(6132) <= a;
    layer3_outputs(6133) <= '1';
    layer3_outputs(6134) <= b;
    layer3_outputs(6135) <= not b;
    layer3_outputs(6136) <= not a or b;
    layer3_outputs(6137) <= a and not b;
    layer3_outputs(6138) <= a and b;
    layer3_outputs(6139) <= a and b;
    layer3_outputs(6140) <= not b;
    layer3_outputs(6141) <= a and not b;
    layer3_outputs(6142) <= not b;
    layer3_outputs(6143) <= '0';
    layer3_outputs(6144) <= b;
    layer3_outputs(6145) <= not (a and b);
    layer3_outputs(6146) <= '0';
    layer3_outputs(6147) <= not (a or b);
    layer3_outputs(6148) <= not b or a;
    layer3_outputs(6149) <= not (a xor b);
    layer3_outputs(6150) <= b and not a;
    layer3_outputs(6151) <= a xor b;
    layer3_outputs(6152) <= not (a or b);
    layer3_outputs(6153) <= not (a or b);
    layer3_outputs(6154) <= not a;
    layer3_outputs(6155) <= a;
    layer3_outputs(6156) <= b;
    layer3_outputs(6157) <= not (a xor b);
    layer3_outputs(6158) <= b;
    layer3_outputs(6159) <= not (a or b);
    layer3_outputs(6160) <= b;
    layer3_outputs(6161) <= a xor b;
    layer3_outputs(6162) <= not (a or b);
    layer3_outputs(6163) <= not (a or b);
    layer3_outputs(6164) <= b and not a;
    layer3_outputs(6165) <= not b or a;
    layer3_outputs(6166) <= a;
    layer3_outputs(6167) <= a and not b;
    layer3_outputs(6168) <= a;
    layer3_outputs(6169) <= b;
    layer3_outputs(6170) <= not (a or b);
    layer3_outputs(6171) <= not (a and b);
    layer3_outputs(6172) <= not b;
    layer3_outputs(6173) <= a and b;
    layer3_outputs(6174) <= not a;
    layer3_outputs(6175) <= not a or b;
    layer3_outputs(6176) <= '0';
    layer3_outputs(6177) <= not a or b;
    layer3_outputs(6178) <= b and not a;
    layer3_outputs(6179) <= a and not b;
    layer3_outputs(6180) <= a;
    layer3_outputs(6181) <= '1';
    layer3_outputs(6182) <= not b;
    layer3_outputs(6183) <= a or b;
    layer3_outputs(6184) <= a;
    layer3_outputs(6185) <= not a;
    layer3_outputs(6186) <= not (a and b);
    layer3_outputs(6187) <= not a;
    layer3_outputs(6188) <= a or b;
    layer3_outputs(6189) <= not a;
    layer3_outputs(6190) <= a;
    layer3_outputs(6191) <= b;
    layer3_outputs(6192) <= not a or b;
    layer3_outputs(6193) <= not a;
    layer3_outputs(6194) <= a;
    layer3_outputs(6195) <= a;
    layer3_outputs(6196) <= a;
    layer3_outputs(6197) <= not (a or b);
    layer3_outputs(6198) <= not b or a;
    layer3_outputs(6199) <= not (a or b);
    layer3_outputs(6200) <= not b or a;
    layer3_outputs(6201) <= '1';
    layer3_outputs(6202) <= b;
    layer3_outputs(6203) <= a;
    layer3_outputs(6204) <= not b or a;
    layer3_outputs(6205) <= not b;
    layer3_outputs(6206) <= b and not a;
    layer3_outputs(6207) <= not (a or b);
    layer3_outputs(6208) <= not b or a;
    layer3_outputs(6209) <= not (a and b);
    layer3_outputs(6210) <= b;
    layer3_outputs(6211) <= not a;
    layer3_outputs(6212) <= not a;
    layer3_outputs(6213) <= not b;
    layer3_outputs(6214) <= not b or a;
    layer3_outputs(6215) <= a and not b;
    layer3_outputs(6216) <= '1';
    layer3_outputs(6217) <= b and not a;
    layer3_outputs(6218) <= not (a or b);
    layer3_outputs(6219) <= not b or a;
    layer3_outputs(6220) <= a xor b;
    layer3_outputs(6221) <= a and b;
    layer3_outputs(6222) <= not (a xor b);
    layer3_outputs(6223) <= b and not a;
    layer3_outputs(6224) <= not a or b;
    layer3_outputs(6225) <= b and not a;
    layer3_outputs(6226) <= a;
    layer3_outputs(6227) <= a xor b;
    layer3_outputs(6228) <= not b or a;
    layer3_outputs(6229) <= not b;
    layer3_outputs(6230) <= '0';
    layer3_outputs(6231) <= a;
    layer3_outputs(6232) <= '0';
    layer3_outputs(6233) <= not b;
    layer3_outputs(6234) <= not a;
    layer3_outputs(6235) <= b;
    layer3_outputs(6236) <= a;
    layer3_outputs(6237) <= not (a or b);
    layer3_outputs(6238) <= b;
    layer3_outputs(6239) <= not a;
    layer3_outputs(6240) <= b and not a;
    layer3_outputs(6241) <= not a or b;
    layer3_outputs(6242) <= b;
    layer3_outputs(6243) <= a xor b;
    layer3_outputs(6244) <= a;
    layer3_outputs(6245) <= not a or b;
    layer3_outputs(6246) <= '0';
    layer3_outputs(6247) <= not a;
    layer3_outputs(6248) <= a or b;
    layer3_outputs(6249) <= not (a xor b);
    layer3_outputs(6250) <= a;
    layer3_outputs(6251) <= not a or b;
    layer3_outputs(6252) <= not a or b;
    layer3_outputs(6253) <= '1';
    layer3_outputs(6254) <= a or b;
    layer3_outputs(6255) <= a and b;
    layer3_outputs(6256) <= not b;
    layer3_outputs(6257) <= not a;
    layer3_outputs(6258) <= not (a xor b);
    layer3_outputs(6259) <= not (a and b);
    layer3_outputs(6260) <= b and not a;
    layer3_outputs(6261) <= not (a or b);
    layer3_outputs(6262) <= not a or b;
    layer3_outputs(6263) <= b;
    layer3_outputs(6264) <= not (a or b);
    layer3_outputs(6265) <= not b;
    layer3_outputs(6266) <= not a or b;
    layer3_outputs(6267) <= a;
    layer3_outputs(6268) <= not b or a;
    layer3_outputs(6269) <= not b;
    layer3_outputs(6270) <= a or b;
    layer3_outputs(6271) <= not b;
    layer3_outputs(6272) <= a;
    layer3_outputs(6273) <= a xor b;
    layer3_outputs(6274) <= not a;
    layer3_outputs(6275) <= '0';
    layer3_outputs(6276) <= '1';
    layer3_outputs(6277) <= not b or a;
    layer3_outputs(6278) <= not (a and b);
    layer3_outputs(6279) <= not b;
    layer3_outputs(6280) <= not a;
    layer3_outputs(6281) <= a and b;
    layer3_outputs(6282) <= not a;
    layer3_outputs(6283) <= not b;
    layer3_outputs(6284) <= a;
    layer3_outputs(6285) <= not b or a;
    layer3_outputs(6286) <= '0';
    layer3_outputs(6287) <= not (a and b);
    layer3_outputs(6288) <= not (a and b);
    layer3_outputs(6289) <= a;
    layer3_outputs(6290) <= a or b;
    layer3_outputs(6291) <= not b or a;
    layer3_outputs(6292) <= a;
    layer3_outputs(6293) <= a and b;
    layer3_outputs(6294) <= not (a xor b);
    layer3_outputs(6295) <= b;
    layer3_outputs(6296) <= not a;
    layer3_outputs(6297) <= not b;
    layer3_outputs(6298) <= not a;
    layer3_outputs(6299) <= not a or b;
    layer3_outputs(6300) <= not a;
    layer3_outputs(6301) <= '1';
    layer3_outputs(6302) <= a;
    layer3_outputs(6303) <= not (a xor b);
    layer3_outputs(6304) <= not a;
    layer3_outputs(6305) <= a;
    layer3_outputs(6306) <= not a;
    layer3_outputs(6307) <= a;
    layer3_outputs(6308) <= not a;
    layer3_outputs(6309) <= a and b;
    layer3_outputs(6310) <= not a or b;
    layer3_outputs(6311) <= '1';
    layer3_outputs(6312) <= not a;
    layer3_outputs(6313) <= a and not b;
    layer3_outputs(6314) <= not (a and b);
    layer3_outputs(6315) <= a;
    layer3_outputs(6316) <= not b;
    layer3_outputs(6317) <= not a or b;
    layer3_outputs(6318) <= a;
    layer3_outputs(6319) <= not (a or b);
    layer3_outputs(6320) <= a and not b;
    layer3_outputs(6321) <= a;
    layer3_outputs(6322) <= b;
    layer3_outputs(6323) <= not b;
    layer3_outputs(6324) <= b;
    layer3_outputs(6325) <= not b;
    layer3_outputs(6326) <= not (a or b);
    layer3_outputs(6327) <= a;
    layer3_outputs(6328) <= not a;
    layer3_outputs(6329) <= '1';
    layer3_outputs(6330) <= b;
    layer3_outputs(6331) <= b;
    layer3_outputs(6332) <= b;
    layer3_outputs(6333) <= not b or a;
    layer3_outputs(6334) <= not (a and b);
    layer3_outputs(6335) <= a and b;
    layer3_outputs(6336) <= a;
    layer3_outputs(6337) <= a and b;
    layer3_outputs(6338) <= a and not b;
    layer3_outputs(6339) <= a xor b;
    layer3_outputs(6340) <= not (a and b);
    layer3_outputs(6341) <= not a;
    layer3_outputs(6342) <= not b;
    layer3_outputs(6343) <= a or b;
    layer3_outputs(6344) <= '1';
    layer3_outputs(6345) <= not b or a;
    layer3_outputs(6346) <= b;
    layer3_outputs(6347) <= a and not b;
    layer3_outputs(6348) <= not (a or b);
    layer3_outputs(6349) <= not (a or b);
    layer3_outputs(6350) <= not a or b;
    layer3_outputs(6351) <= '1';
    layer3_outputs(6352) <= not a;
    layer3_outputs(6353) <= not (a or b);
    layer3_outputs(6354) <= a and b;
    layer3_outputs(6355) <= not a;
    layer3_outputs(6356) <= a or b;
    layer3_outputs(6357) <= a and b;
    layer3_outputs(6358) <= not (a and b);
    layer3_outputs(6359) <= not b;
    layer3_outputs(6360) <= not (a or b);
    layer3_outputs(6361) <= not (a or b);
    layer3_outputs(6362) <= not a or b;
    layer3_outputs(6363) <= not a or b;
    layer3_outputs(6364) <= a;
    layer3_outputs(6365) <= '0';
    layer3_outputs(6366) <= not b;
    layer3_outputs(6367) <= b and not a;
    layer3_outputs(6368) <= b;
    layer3_outputs(6369) <= not b;
    layer3_outputs(6370) <= not b or a;
    layer3_outputs(6371) <= not b;
    layer3_outputs(6372) <= not a or b;
    layer3_outputs(6373) <= a or b;
    layer3_outputs(6374) <= a and not b;
    layer3_outputs(6375) <= b and not a;
    layer3_outputs(6376) <= not b;
    layer3_outputs(6377) <= not b or a;
    layer3_outputs(6378) <= a;
    layer3_outputs(6379) <= b and not a;
    layer3_outputs(6380) <= not (a xor b);
    layer3_outputs(6381) <= not a;
    layer3_outputs(6382) <= '1';
    layer3_outputs(6383) <= not b;
    layer3_outputs(6384) <= not a or b;
    layer3_outputs(6385) <= not a or b;
    layer3_outputs(6386) <= b;
    layer3_outputs(6387) <= a and not b;
    layer3_outputs(6388) <= not b;
    layer3_outputs(6389) <= b and not a;
    layer3_outputs(6390) <= not (a or b);
    layer3_outputs(6391) <= not b;
    layer3_outputs(6392) <= not (a or b);
    layer3_outputs(6393) <= a xor b;
    layer3_outputs(6394) <= a;
    layer3_outputs(6395) <= a and not b;
    layer3_outputs(6396) <= not (a or b);
    layer3_outputs(6397) <= b;
    layer3_outputs(6398) <= '1';
    layer3_outputs(6399) <= a xor b;
    layer3_outputs(6400) <= not (a or b);
    layer3_outputs(6401) <= a and not b;
    layer3_outputs(6402) <= a and b;
    layer3_outputs(6403) <= a and b;
    layer3_outputs(6404) <= not b;
    layer3_outputs(6405) <= not b;
    layer3_outputs(6406) <= not (a and b);
    layer3_outputs(6407) <= '0';
    layer3_outputs(6408) <= '0';
    layer3_outputs(6409) <= not (a xor b);
    layer3_outputs(6410) <= not b;
    layer3_outputs(6411) <= not b;
    layer3_outputs(6412) <= not a or b;
    layer3_outputs(6413) <= not a or b;
    layer3_outputs(6414) <= not (a or b);
    layer3_outputs(6415) <= a;
    layer3_outputs(6416) <= a and b;
    layer3_outputs(6417) <= a or b;
    layer3_outputs(6418) <= b;
    layer3_outputs(6419) <= '0';
    layer3_outputs(6420) <= a;
    layer3_outputs(6421) <= not a;
    layer3_outputs(6422) <= a and b;
    layer3_outputs(6423) <= not b;
    layer3_outputs(6424) <= not b;
    layer3_outputs(6425) <= not b;
    layer3_outputs(6426) <= not a or b;
    layer3_outputs(6427) <= not a or b;
    layer3_outputs(6428) <= not (a xor b);
    layer3_outputs(6429) <= a or b;
    layer3_outputs(6430) <= '1';
    layer3_outputs(6431) <= b;
    layer3_outputs(6432) <= b;
    layer3_outputs(6433) <= not (a or b);
    layer3_outputs(6434) <= b;
    layer3_outputs(6435) <= not b;
    layer3_outputs(6436) <= '0';
    layer3_outputs(6437) <= a and not b;
    layer3_outputs(6438) <= a and b;
    layer3_outputs(6439) <= a and not b;
    layer3_outputs(6440) <= not (a xor b);
    layer3_outputs(6441) <= not b;
    layer3_outputs(6442) <= not (a or b);
    layer3_outputs(6443) <= b;
    layer3_outputs(6444) <= a or b;
    layer3_outputs(6445) <= b;
    layer3_outputs(6446) <= b;
    layer3_outputs(6447) <= not a or b;
    layer3_outputs(6448) <= not a;
    layer3_outputs(6449) <= not (a xor b);
    layer3_outputs(6450) <= not a or b;
    layer3_outputs(6451) <= not (a or b);
    layer3_outputs(6452) <= b;
    layer3_outputs(6453) <= a and not b;
    layer3_outputs(6454) <= '1';
    layer3_outputs(6455) <= a;
    layer3_outputs(6456) <= b;
    layer3_outputs(6457) <= a and not b;
    layer3_outputs(6458) <= '1';
    layer3_outputs(6459) <= b;
    layer3_outputs(6460) <= not b;
    layer3_outputs(6461) <= b and not a;
    layer3_outputs(6462) <= not (a xor b);
    layer3_outputs(6463) <= not b or a;
    layer3_outputs(6464) <= a and b;
    layer3_outputs(6465) <= not b or a;
    layer3_outputs(6466) <= b and not a;
    layer3_outputs(6467) <= not b;
    layer3_outputs(6468) <= b and not a;
    layer3_outputs(6469) <= a;
    layer3_outputs(6470) <= b;
    layer3_outputs(6471) <= b;
    layer3_outputs(6472) <= b and not a;
    layer3_outputs(6473) <= not b;
    layer3_outputs(6474) <= b;
    layer3_outputs(6475) <= b and not a;
    layer3_outputs(6476) <= not a;
    layer3_outputs(6477) <= '1';
    layer3_outputs(6478) <= not b;
    layer3_outputs(6479) <= not a or b;
    layer3_outputs(6480) <= a and not b;
    layer3_outputs(6481) <= not b;
    layer3_outputs(6482) <= not a or b;
    layer3_outputs(6483) <= a;
    layer3_outputs(6484) <= not (a or b);
    layer3_outputs(6485) <= a and b;
    layer3_outputs(6486) <= not (a and b);
    layer3_outputs(6487) <= a;
    layer3_outputs(6488) <= b and not a;
    layer3_outputs(6489) <= not a or b;
    layer3_outputs(6490) <= not (a xor b);
    layer3_outputs(6491) <= b and not a;
    layer3_outputs(6492) <= not (a and b);
    layer3_outputs(6493) <= '0';
    layer3_outputs(6494) <= not a;
    layer3_outputs(6495) <= a and not b;
    layer3_outputs(6496) <= a xor b;
    layer3_outputs(6497) <= not b;
    layer3_outputs(6498) <= not (a or b);
    layer3_outputs(6499) <= not (a or b);
    layer3_outputs(6500) <= a and b;
    layer3_outputs(6501) <= b;
    layer3_outputs(6502) <= not b;
    layer3_outputs(6503) <= not (a and b);
    layer3_outputs(6504) <= not a;
    layer3_outputs(6505) <= '1';
    layer3_outputs(6506) <= not a;
    layer3_outputs(6507) <= not b;
    layer3_outputs(6508) <= not a;
    layer3_outputs(6509) <= a and b;
    layer3_outputs(6510) <= b;
    layer3_outputs(6511) <= not (a and b);
    layer3_outputs(6512) <= a;
    layer3_outputs(6513) <= not a or b;
    layer3_outputs(6514) <= not b or a;
    layer3_outputs(6515) <= b;
    layer3_outputs(6516) <= b;
    layer3_outputs(6517) <= '0';
    layer3_outputs(6518) <= not (a or b);
    layer3_outputs(6519) <= not b or a;
    layer3_outputs(6520) <= a and not b;
    layer3_outputs(6521) <= a;
    layer3_outputs(6522) <= b;
    layer3_outputs(6523) <= a xor b;
    layer3_outputs(6524) <= a;
    layer3_outputs(6525) <= not b or a;
    layer3_outputs(6526) <= '0';
    layer3_outputs(6527) <= not (a and b);
    layer3_outputs(6528) <= not a or b;
    layer3_outputs(6529) <= not (a and b);
    layer3_outputs(6530) <= not b;
    layer3_outputs(6531) <= a;
    layer3_outputs(6532) <= not b;
    layer3_outputs(6533) <= not (a or b);
    layer3_outputs(6534) <= '1';
    layer3_outputs(6535) <= b and not a;
    layer3_outputs(6536) <= not a;
    layer3_outputs(6537) <= b;
    layer3_outputs(6538) <= b and not a;
    layer3_outputs(6539) <= not (a xor b);
    layer3_outputs(6540) <= not (a and b);
    layer3_outputs(6541) <= a and b;
    layer3_outputs(6542) <= a or b;
    layer3_outputs(6543) <= not b;
    layer3_outputs(6544) <= not b or a;
    layer3_outputs(6545) <= a;
    layer3_outputs(6546) <= not b or a;
    layer3_outputs(6547) <= b and not a;
    layer3_outputs(6548) <= not (a and b);
    layer3_outputs(6549) <= b and not a;
    layer3_outputs(6550) <= b and not a;
    layer3_outputs(6551) <= not a;
    layer3_outputs(6552) <= not b;
    layer3_outputs(6553) <= b and not a;
    layer3_outputs(6554) <= not (a xor b);
    layer3_outputs(6555) <= a and b;
    layer3_outputs(6556) <= not b or a;
    layer3_outputs(6557) <= '1';
    layer3_outputs(6558) <= a and not b;
    layer3_outputs(6559) <= not (a or b);
    layer3_outputs(6560) <= a and not b;
    layer3_outputs(6561) <= a and not b;
    layer3_outputs(6562) <= a and not b;
    layer3_outputs(6563) <= not b or a;
    layer3_outputs(6564) <= b and not a;
    layer3_outputs(6565) <= b;
    layer3_outputs(6566) <= not (a and b);
    layer3_outputs(6567) <= not (a or b);
    layer3_outputs(6568) <= not (a xor b);
    layer3_outputs(6569) <= a or b;
    layer3_outputs(6570) <= b and not a;
    layer3_outputs(6571) <= not b;
    layer3_outputs(6572) <= b and not a;
    layer3_outputs(6573) <= not (a and b);
    layer3_outputs(6574) <= not (a and b);
    layer3_outputs(6575) <= not b;
    layer3_outputs(6576) <= not (a xor b);
    layer3_outputs(6577) <= not a or b;
    layer3_outputs(6578) <= a;
    layer3_outputs(6579) <= not a;
    layer3_outputs(6580) <= a xor b;
    layer3_outputs(6581) <= not a;
    layer3_outputs(6582) <= not a;
    layer3_outputs(6583) <= b;
    layer3_outputs(6584) <= a;
    layer3_outputs(6585) <= not (a and b);
    layer3_outputs(6586) <= not (a or b);
    layer3_outputs(6587) <= not b;
    layer3_outputs(6588) <= a and not b;
    layer3_outputs(6589) <= not (a xor b);
    layer3_outputs(6590) <= not b;
    layer3_outputs(6591) <= not (a and b);
    layer3_outputs(6592) <= not (a and b);
    layer3_outputs(6593) <= a;
    layer3_outputs(6594) <= not a or b;
    layer3_outputs(6595) <= not b;
    layer3_outputs(6596) <= b and not a;
    layer3_outputs(6597) <= a and not b;
    layer3_outputs(6598) <= not b or a;
    layer3_outputs(6599) <= '0';
    layer3_outputs(6600) <= a or b;
    layer3_outputs(6601) <= b;
    layer3_outputs(6602) <= not b;
    layer3_outputs(6603) <= not b or a;
    layer3_outputs(6604) <= a;
    layer3_outputs(6605) <= not b;
    layer3_outputs(6606) <= not b;
    layer3_outputs(6607) <= b and not a;
    layer3_outputs(6608) <= '0';
    layer3_outputs(6609) <= a;
    layer3_outputs(6610) <= not b;
    layer3_outputs(6611) <= not b;
    layer3_outputs(6612) <= not a;
    layer3_outputs(6613) <= not a;
    layer3_outputs(6614) <= a;
    layer3_outputs(6615) <= a and b;
    layer3_outputs(6616) <= not a or b;
    layer3_outputs(6617) <= a;
    layer3_outputs(6618) <= not b;
    layer3_outputs(6619) <= '0';
    layer3_outputs(6620) <= b;
    layer3_outputs(6621) <= not a or b;
    layer3_outputs(6622) <= a or b;
    layer3_outputs(6623) <= not (a or b);
    layer3_outputs(6624) <= a and not b;
    layer3_outputs(6625) <= a xor b;
    layer3_outputs(6626) <= not b;
    layer3_outputs(6627) <= b;
    layer3_outputs(6628) <= not (a and b);
    layer3_outputs(6629) <= a and not b;
    layer3_outputs(6630) <= b and not a;
    layer3_outputs(6631) <= not a;
    layer3_outputs(6632) <= a and b;
    layer3_outputs(6633) <= a;
    layer3_outputs(6634) <= b;
    layer3_outputs(6635) <= a xor b;
    layer3_outputs(6636) <= a or b;
    layer3_outputs(6637) <= not b or a;
    layer3_outputs(6638) <= b;
    layer3_outputs(6639) <= a xor b;
    layer3_outputs(6640) <= not b or a;
    layer3_outputs(6641) <= a and b;
    layer3_outputs(6642) <= not (a or b);
    layer3_outputs(6643) <= a and not b;
    layer3_outputs(6644) <= not b or a;
    layer3_outputs(6645) <= not (a xor b);
    layer3_outputs(6646) <= b and not a;
    layer3_outputs(6647) <= a;
    layer3_outputs(6648) <= b;
    layer3_outputs(6649) <= a;
    layer3_outputs(6650) <= a;
    layer3_outputs(6651) <= not (a xor b);
    layer3_outputs(6652) <= not b;
    layer3_outputs(6653) <= a;
    layer3_outputs(6654) <= not (a and b);
    layer3_outputs(6655) <= not b;
    layer3_outputs(6656) <= not (a or b);
    layer3_outputs(6657) <= '1';
    layer3_outputs(6658) <= a and not b;
    layer3_outputs(6659) <= a and b;
    layer3_outputs(6660) <= not (a or b);
    layer3_outputs(6661) <= a;
    layer3_outputs(6662) <= not b or a;
    layer3_outputs(6663) <= not (a or b);
    layer3_outputs(6664) <= not a;
    layer3_outputs(6665) <= not (a or b);
    layer3_outputs(6666) <= not b;
    layer3_outputs(6667) <= b;
    layer3_outputs(6668) <= a and not b;
    layer3_outputs(6669) <= not b or a;
    layer3_outputs(6670) <= not a;
    layer3_outputs(6671) <= not (a or b);
    layer3_outputs(6672) <= b;
    layer3_outputs(6673) <= a or b;
    layer3_outputs(6674) <= not a or b;
    layer3_outputs(6675) <= a;
    layer3_outputs(6676) <= not a or b;
    layer3_outputs(6677) <= b;
    layer3_outputs(6678) <= not b or a;
    layer3_outputs(6679) <= not (a or b);
    layer3_outputs(6680) <= a or b;
    layer3_outputs(6681) <= a or b;
    layer3_outputs(6682) <= b;
    layer3_outputs(6683) <= not a or b;
    layer3_outputs(6684) <= not (a and b);
    layer3_outputs(6685) <= not b;
    layer3_outputs(6686) <= a and not b;
    layer3_outputs(6687) <= not (a and b);
    layer3_outputs(6688) <= not (a xor b);
    layer3_outputs(6689) <= b and not a;
    layer3_outputs(6690) <= a and not b;
    layer3_outputs(6691) <= a xor b;
    layer3_outputs(6692) <= not a or b;
    layer3_outputs(6693) <= not a;
    layer3_outputs(6694) <= not (a or b);
    layer3_outputs(6695) <= a and b;
    layer3_outputs(6696) <= not a;
    layer3_outputs(6697) <= not a;
    layer3_outputs(6698) <= b;
    layer3_outputs(6699) <= '1';
    layer3_outputs(6700) <= a;
    layer3_outputs(6701) <= a xor b;
    layer3_outputs(6702) <= a xor b;
    layer3_outputs(6703) <= '1';
    layer3_outputs(6704) <= a;
    layer3_outputs(6705) <= not b;
    layer3_outputs(6706) <= not a or b;
    layer3_outputs(6707) <= b and not a;
    layer3_outputs(6708) <= a and b;
    layer3_outputs(6709) <= not b or a;
    layer3_outputs(6710) <= a;
    layer3_outputs(6711) <= not (a and b);
    layer3_outputs(6712) <= not a or b;
    layer3_outputs(6713) <= not b or a;
    layer3_outputs(6714) <= a and not b;
    layer3_outputs(6715) <= a;
    layer3_outputs(6716) <= not b;
    layer3_outputs(6717) <= '1';
    layer3_outputs(6718) <= b;
    layer3_outputs(6719) <= not b;
    layer3_outputs(6720) <= not a;
    layer3_outputs(6721) <= not b;
    layer3_outputs(6722) <= a xor b;
    layer3_outputs(6723) <= not b;
    layer3_outputs(6724) <= not (a xor b);
    layer3_outputs(6725) <= a;
    layer3_outputs(6726) <= a or b;
    layer3_outputs(6727) <= '1';
    layer3_outputs(6728) <= not a;
    layer3_outputs(6729) <= not (a or b);
    layer3_outputs(6730) <= not (a or b);
    layer3_outputs(6731) <= not b;
    layer3_outputs(6732) <= not a;
    layer3_outputs(6733) <= not a or b;
    layer3_outputs(6734) <= '1';
    layer3_outputs(6735) <= not (a or b);
    layer3_outputs(6736) <= a and not b;
    layer3_outputs(6737) <= b and not a;
    layer3_outputs(6738) <= b;
    layer3_outputs(6739) <= a and b;
    layer3_outputs(6740) <= b;
    layer3_outputs(6741) <= not (a and b);
    layer3_outputs(6742) <= a;
    layer3_outputs(6743) <= '0';
    layer3_outputs(6744) <= not b or a;
    layer3_outputs(6745) <= a and b;
    layer3_outputs(6746) <= not a;
    layer3_outputs(6747) <= '0';
    layer3_outputs(6748) <= b;
    layer3_outputs(6749) <= b;
    layer3_outputs(6750) <= b;
    layer3_outputs(6751) <= not a;
    layer3_outputs(6752) <= not b or a;
    layer3_outputs(6753) <= a xor b;
    layer3_outputs(6754) <= '1';
    layer3_outputs(6755) <= a and not b;
    layer3_outputs(6756) <= b;
    layer3_outputs(6757) <= not b;
    layer3_outputs(6758) <= not b;
    layer3_outputs(6759) <= not b or a;
    layer3_outputs(6760) <= not (a xor b);
    layer3_outputs(6761) <= not b;
    layer3_outputs(6762) <= not a or b;
    layer3_outputs(6763) <= a or b;
    layer3_outputs(6764) <= a and not b;
    layer3_outputs(6765) <= a and b;
    layer3_outputs(6766) <= not (a and b);
    layer3_outputs(6767) <= a;
    layer3_outputs(6768) <= not a;
    layer3_outputs(6769) <= not (a and b);
    layer3_outputs(6770) <= b;
    layer3_outputs(6771) <= a or b;
    layer3_outputs(6772) <= not b;
    layer3_outputs(6773) <= '0';
    layer3_outputs(6774) <= not a or b;
    layer3_outputs(6775) <= b;
    layer3_outputs(6776) <= b;
    layer3_outputs(6777) <= not (a or b);
    layer3_outputs(6778) <= a;
    layer3_outputs(6779) <= not b;
    layer3_outputs(6780) <= not (a or b);
    layer3_outputs(6781) <= b;
    layer3_outputs(6782) <= a;
    layer3_outputs(6783) <= '0';
    layer3_outputs(6784) <= b and not a;
    layer3_outputs(6785) <= not (a or b);
    layer3_outputs(6786) <= '0';
    layer3_outputs(6787) <= a;
    layer3_outputs(6788) <= not a;
    layer3_outputs(6789) <= not a;
    layer3_outputs(6790) <= b;
    layer3_outputs(6791) <= not (a and b);
    layer3_outputs(6792) <= a;
    layer3_outputs(6793) <= not a or b;
    layer3_outputs(6794) <= b;
    layer3_outputs(6795) <= not (a or b);
    layer3_outputs(6796) <= not a or b;
    layer3_outputs(6797) <= not a or b;
    layer3_outputs(6798) <= a and not b;
    layer3_outputs(6799) <= b;
    layer3_outputs(6800) <= not b;
    layer3_outputs(6801) <= a or b;
    layer3_outputs(6802) <= not a;
    layer3_outputs(6803) <= a or b;
    layer3_outputs(6804) <= not b;
    layer3_outputs(6805) <= not a;
    layer3_outputs(6806) <= b;
    layer3_outputs(6807) <= not b;
    layer3_outputs(6808) <= not (a and b);
    layer3_outputs(6809) <= not a;
    layer3_outputs(6810) <= a and b;
    layer3_outputs(6811) <= '1';
    layer3_outputs(6812) <= a and not b;
    layer3_outputs(6813) <= not (a xor b);
    layer3_outputs(6814) <= not (a or b);
    layer3_outputs(6815) <= a;
    layer3_outputs(6816) <= not a;
    layer3_outputs(6817) <= not (a or b);
    layer3_outputs(6818) <= not b or a;
    layer3_outputs(6819) <= a and b;
    layer3_outputs(6820) <= not b;
    layer3_outputs(6821) <= b;
    layer3_outputs(6822) <= not b;
    layer3_outputs(6823) <= b and not a;
    layer3_outputs(6824) <= not (a or b);
    layer3_outputs(6825) <= a and not b;
    layer3_outputs(6826) <= a;
    layer3_outputs(6827) <= not a;
    layer3_outputs(6828) <= not a;
    layer3_outputs(6829) <= a and not b;
    layer3_outputs(6830) <= not (a and b);
    layer3_outputs(6831) <= '0';
    layer3_outputs(6832) <= not b or a;
    layer3_outputs(6833) <= a;
    layer3_outputs(6834) <= b and not a;
    layer3_outputs(6835) <= not (a or b);
    layer3_outputs(6836) <= not (a xor b);
    layer3_outputs(6837) <= b;
    layer3_outputs(6838) <= not b or a;
    layer3_outputs(6839) <= b and not a;
    layer3_outputs(6840) <= not b;
    layer3_outputs(6841) <= b;
    layer3_outputs(6842) <= b;
    layer3_outputs(6843) <= not (a or b);
    layer3_outputs(6844) <= not (a xor b);
    layer3_outputs(6845) <= '0';
    layer3_outputs(6846) <= b;
    layer3_outputs(6847) <= not (a or b);
    layer3_outputs(6848) <= not (a or b);
    layer3_outputs(6849) <= b;
    layer3_outputs(6850) <= a and not b;
    layer3_outputs(6851) <= not (a or b);
    layer3_outputs(6852) <= not (a or b);
    layer3_outputs(6853) <= b and not a;
    layer3_outputs(6854) <= not a or b;
    layer3_outputs(6855) <= a or b;
    layer3_outputs(6856) <= not (a or b);
    layer3_outputs(6857) <= not (a or b);
    layer3_outputs(6858) <= not b;
    layer3_outputs(6859) <= not a;
    layer3_outputs(6860) <= not b or a;
    layer3_outputs(6861) <= a or b;
    layer3_outputs(6862) <= b;
    layer3_outputs(6863) <= a xor b;
    layer3_outputs(6864) <= a xor b;
    layer3_outputs(6865) <= b;
    layer3_outputs(6866) <= a;
    layer3_outputs(6867) <= b;
    layer3_outputs(6868) <= b and not a;
    layer3_outputs(6869) <= '1';
    layer3_outputs(6870) <= not b or a;
    layer3_outputs(6871) <= not (a or b);
    layer3_outputs(6872) <= not (a and b);
    layer3_outputs(6873) <= not a;
    layer3_outputs(6874) <= not a;
    layer3_outputs(6875) <= a;
    layer3_outputs(6876) <= '0';
    layer3_outputs(6877) <= not (a or b);
    layer3_outputs(6878) <= b;
    layer3_outputs(6879) <= b and not a;
    layer3_outputs(6880) <= not (a and b);
    layer3_outputs(6881) <= '0';
    layer3_outputs(6882) <= not b;
    layer3_outputs(6883) <= not (a or b);
    layer3_outputs(6884) <= not b;
    layer3_outputs(6885) <= a;
    layer3_outputs(6886) <= b;
    layer3_outputs(6887) <= not b or a;
    layer3_outputs(6888) <= b;
    layer3_outputs(6889) <= not b;
    layer3_outputs(6890) <= b;
    layer3_outputs(6891) <= not a;
    layer3_outputs(6892) <= a xor b;
    layer3_outputs(6893) <= not a;
    layer3_outputs(6894) <= not b;
    layer3_outputs(6895) <= a xor b;
    layer3_outputs(6896) <= not a;
    layer3_outputs(6897) <= not b;
    layer3_outputs(6898) <= not a or b;
    layer3_outputs(6899) <= not (a or b);
    layer3_outputs(6900) <= a and b;
    layer3_outputs(6901) <= not (a xor b);
    layer3_outputs(6902) <= '1';
    layer3_outputs(6903) <= a;
    layer3_outputs(6904) <= not (a and b);
    layer3_outputs(6905) <= not b or a;
    layer3_outputs(6906) <= not b;
    layer3_outputs(6907) <= not a or b;
    layer3_outputs(6908) <= a and not b;
    layer3_outputs(6909) <= not a or b;
    layer3_outputs(6910) <= not a;
    layer3_outputs(6911) <= '1';
    layer3_outputs(6912) <= not b or a;
    layer3_outputs(6913) <= a or b;
    layer3_outputs(6914) <= not (a and b);
    layer3_outputs(6915) <= not b;
    layer3_outputs(6916) <= not b or a;
    layer3_outputs(6917) <= a and b;
    layer3_outputs(6918) <= a and b;
    layer3_outputs(6919) <= '0';
    layer3_outputs(6920) <= not (a or b);
    layer3_outputs(6921) <= not b;
    layer3_outputs(6922) <= b;
    layer3_outputs(6923) <= a or b;
    layer3_outputs(6924) <= b;
    layer3_outputs(6925) <= not (a xor b);
    layer3_outputs(6926) <= a xor b;
    layer3_outputs(6927) <= a;
    layer3_outputs(6928) <= '1';
    layer3_outputs(6929) <= not (a or b);
    layer3_outputs(6930) <= a;
    layer3_outputs(6931) <= b;
    layer3_outputs(6932) <= b;
    layer3_outputs(6933) <= b;
    layer3_outputs(6934) <= b;
    layer3_outputs(6935) <= b;
    layer3_outputs(6936) <= not a or b;
    layer3_outputs(6937) <= not b;
    layer3_outputs(6938) <= not a;
    layer3_outputs(6939) <= a or b;
    layer3_outputs(6940) <= not a or b;
    layer3_outputs(6941) <= '0';
    layer3_outputs(6942) <= '0';
    layer3_outputs(6943) <= a or b;
    layer3_outputs(6944) <= not a;
    layer3_outputs(6945) <= not a;
    layer3_outputs(6946) <= not a or b;
    layer3_outputs(6947) <= a;
    layer3_outputs(6948) <= not b;
    layer3_outputs(6949) <= not b or a;
    layer3_outputs(6950) <= not (a and b);
    layer3_outputs(6951) <= a xor b;
    layer3_outputs(6952) <= a;
    layer3_outputs(6953) <= not b or a;
    layer3_outputs(6954) <= b and not a;
    layer3_outputs(6955) <= not (a xor b);
    layer3_outputs(6956) <= not a;
    layer3_outputs(6957) <= b and not a;
    layer3_outputs(6958) <= '0';
    layer3_outputs(6959) <= not a or b;
    layer3_outputs(6960) <= not (a or b);
    layer3_outputs(6961) <= '0';
    layer3_outputs(6962) <= a;
    layer3_outputs(6963) <= a and not b;
    layer3_outputs(6964) <= b;
    layer3_outputs(6965) <= not (a and b);
    layer3_outputs(6966) <= a and b;
    layer3_outputs(6967) <= a xor b;
    layer3_outputs(6968) <= not b;
    layer3_outputs(6969) <= '0';
    layer3_outputs(6970) <= b;
    layer3_outputs(6971) <= b;
    layer3_outputs(6972) <= a and b;
    layer3_outputs(6973) <= a and not b;
    layer3_outputs(6974) <= a xor b;
    layer3_outputs(6975) <= a or b;
    layer3_outputs(6976) <= not (a or b);
    layer3_outputs(6977) <= b;
    layer3_outputs(6978) <= b;
    layer3_outputs(6979) <= a and b;
    layer3_outputs(6980) <= not a;
    layer3_outputs(6981) <= not b;
    layer3_outputs(6982) <= '1';
    layer3_outputs(6983) <= not (a and b);
    layer3_outputs(6984) <= a;
    layer3_outputs(6985) <= not a;
    layer3_outputs(6986) <= not (a or b);
    layer3_outputs(6987) <= not a;
    layer3_outputs(6988) <= b;
    layer3_outputs(6989) <= '1';
    layer3_outputs(6990) <= a and b;
    layer3_outputs(6991) <= not b;
    layer3_outputs(6992) <= not a or b;
    layer3_outputs(6993) <= '1';
    layer3_outputs(6994) <= not b;
    layer3_outputs(6995) <= not (a xor b);
    layer3_outputs(6996) <= a or b;
    layer3_outputs(6997) <= not (a or b);
    layer3_outputs(6998) <= a or b;
    layer3_outputs(6999) <= not b;
    layer3_outputs(7000) <= a or b;
    layer3_outputs(7001) <= not (a or b);
    layer3_outputs(7002) <= a xor b;
    layer3_outputs(7003) <= not (a and b);
    layer3_outputs(7004) <= b and not a;
    layer3_outputs(7005) <= a;
    layer3_outputs(7006) <= not b;
    layer3_outputs(7007) <= not (a or b);
    layer3_outputs(7008) <= '0';
    layer3_outputs(7009) <= not b;
    layer3_outputs(7010) <= a;
    layer3_outputs(7011) <= a;
    layer3_outputs(7012) <= b and not a;
    layer3_outputs(7013) <= not (a and b);
    layer3_outputs(7014) <= not (a and b);
    layer3_outputs(7015) <= a or b;
    layer3_outputs(7016) <= a xor b;
    layer3_outputs(7017) <= a;
    layer3_outputs(7018) <= '1';
    layer3_outputs(7019) <= '1';
    layer3_outputs(7020) <= not a or b;
    layer3_outputs(7021) <= not b;
    layer3_outputs(7022) <= not (a and b);
    layer3_outputs(7023) <= b;
    layer3_outputs(7024) <= not a;
    layer3_outputs(7025) <= not (a and b);
    layer3_outputs(7026) <= a and b;
    layer3_outputs(7027) <= a and not b;
    layer3_outputs(7028) <= not a;
    layer3_outputs(7029) <= not (a or b);
    layer3_outputs(7030) <= b;
    layer3_outputs(7031) <= not a;
    layer3_outputs(7032) <= not b;
    layer3_outputs(7033) <= a;
    layer3_outputs(7034) <= not b;
    layer3_outputs(7035) <= not (a or b);
    layer3_outputs(7036) <= a and not b;
    layer3_outputs(7037) <= not (a and b);
    layer3_outputs(7038) <= not b;
    layer3_outputs(7039) <= not b or a;
    layer3_outputs(7040) <= not b;
    layer3_outputs(7041) <= not a or b;
    layer3_outputs(7042) <= not a;
    layer3_outputs(7043) <= not a;
    layer3_outputs(7044) <= b;
    layer3_outputs(7045) <= not (a or b);
    layer3_outputs(7046) <= b and not a;
    layer3_outputs(7047) <= not (a and b);
    layer3_outputs(7048) <= not b;
    layer3_outputs(7049) <= not (a xor b);
    layer3_outputs(7050) <= not (a xor b);
    layer3_outputs(7051) <= a;
    layer3_outputs(7052) <= '1';
    layer3_outputs(7053) <= a;
    layer3_outputs(7054) <= b;
    layer3_outputs(7055) <= not (a or b);
    layer3_outputs(7056) <= not (a and b);
    layer3_outputs(7057) <= not a or b;
    layer3_outputs(7058) <= not a;
    layer3_outputs(7059) <= not b or a;
    layer3_outputs(7060) <= not b;
    layer3_outputs(7061) <= a and not b;
    layer3_outputs(7062) <= a or b;
    layer3_outputs(7063) <= b and not a;
    layer3_outputs(7064) <= not (a or b);
    layer3_outputs(7065) <= b;
    layer3_outputs(7066) <= a and b;
    layer3_outputs(7067) <= a xor b;
    layer3_outputs(7068) <= a;
    layer3_outputs(7069) <= '0';
    layer3_outputs(7070) <= '0';
    layer3_outputs(7071) <= a;
    layer3_outputs(7072) <= a;
    layer3_outputs(7073) <= not a or b;
    layer3_outputs(7074) <= b;
    layer3_outputs(7075) <= not (a and b);
    layer3_outputs(7076) <= not b or a;
    layer3_outputs(7077) <= not (a xor b);
    layer3_outputs(7078) <= a;
    layer3_outputs(7079) <= not a;
    layer3_outputs(7080) <= not b or a;
    layer3_outputs(7081) <= a or b;
    layer3_outputs(7082) <= not a;
    layer3_outputs(7083) <= not a or b;
    layer3_outputs(7084) <= b and not a;
    layer3_outputs(7085) <= not (a or b);
    layer3_outputs(7086) <= a and b;
    layer3_outputs(7087) <= not a or b;
    layer3_outputs(7088) <= not (a xor b);
    layer3_outputs(7089) <= a or b;
    layer3_outputs(7090) <= b and not a;
    layer3_outputs(7091) <= not a;
    layer3_outputs(7092) <= not (a xor b);
    layer3_outputs(7093) <= a and not b;
    layer3_outputs(7094) <= b;
    layer3_outputs(7095) <= a and not b;
    layer3_outputs(7096) <= not (a xor b);
    layer3_outputs(7097) <= not a;
    layer3_outputs(7098) <= a or b;
    layer3_outputs(7099) <= not a;
    layer3_outputs(7100) <= not (a or b);
    layer3_outputs(7101) <= b and not a;
    layer3_outputs(7102) <= not (a xor b);
    layer3_outputs(7103) <= not a;
    layer3_outputs(7104) <= not a;
    layer3_outputs(7105) <= not b or a;
    layer3_outputs(7106) <= a and not b;
    layer3_outputs(7107) <= not b or a;
    layer3_outputs(7108) <= a or b;
    layer3_outputs(7109) <= '0';
    layer3_outputs(7110) <= '1';
    layer3_outputs(7111) <= not a;
    layer3_outputs(7112) <= a xor b;
    layer3_outputs(7113) <= b;
    layer3_outputs(7114) <= b;
    layer3_outputs(7115) <= not (a and b);
    layer3_outputs(7116) <= not (a and b);
    layer3_outputs(7117) <= '0';
    layer3_outputs(7118) <= a or b;
    layer3_outputs(7119) <= a and not b;
    layer3_outputs(7120) <= b and not a;
    layer3_outputs(7121) <= '1';
    layer3_outputs(7122) <= not a or b;
    layer3_outputs(7123) <= a and b;
    layer3_outputs(7124) <= a or b;
    layer3_outputs(7125) <= a;
    layer3_outputs(7126) <= a and b;
    layer3_outputs(7127) <= b;
    layer3_outputs(7128) <= not a;
    layer3_outputs(7129) <= not a;
    layer3_outputs(7130) <= not b or a;
    layer3_outputs(7131) <= a and b;
    layer3_outputs(7132) <= '0';
    layer3_outputs(7133) <= not a or b;
    layer3_outputs(7134) <= not (a xor b);
    layer3_outputs(7135) <= not a;
    layer3_outputs(7136) <= not b;
    layer3_outputs(7137) <= not (a and b);
    layer3_outputs(7138) <= '1';
    layer3_outputs(7139) <= '1';
    layer3_outputs(7140) <= b and not a;
    layer3_outputs(7141) <= b;
    layer3_outputs(7142) <= '0';
    layer3_outputs(7143) <= not b;
    layer3_outputs(7144) <= not (a or b);
    layer3_outputs(7145) <= b;
    layer3_outputs(7146) <= not b;
    layer3_outputs(7147) <= not a;
    layer3_outputs(7148) <= not a or b;
    layer3_outputs(7149) <= b and not a;
    layer3_outputs(7150) <= a;
    layer3_outputs(7151) <= a xor b;
    layer3_outputs(7152) <= not a or b;
    layer3_outputs(7153) <= a and b;
    layer3_outputs(7154) <= not b or a;
    layer3_outputs(7155) <= a or b;
    layer3_outputs(7156) <= a;
    layer3_outputs(7157) <= a;
    layer3_outputs(7158) <= not b or a;
    layer3_outputs(7159) <= '0';
    layer3_outputs(7160) <= not (a and b);
    layer3_outputs(7161) <= b and not a;
    layer3_outputs(7162) <= '1';
    layer3_outputs(7163) <= a xor b;
    layer3_outputs(7164) <= not b or a;
    layer3_outputs(7165) <= not (a or b);
    layer3_outputs(7166) <= not (a xor b);
    layer3_outputs(7167) <= a and b;
    layer3_outputs(7168) <= not b;
    layer3_outputs(7169) <= not (a and b);
    layer3_outputs(7170) <= not (a or b);
    layer3_outputs(7171) <= b;
    layer3_outputs(7172) <= not b or a;
    layer3_outputs(7173) <= not a or b;
    layer3_outputs(7174) <= not a;
    layer3_outputs(7175) <= not (a and b);
    layer3_outputs(7176) <= not (a or b);
    layer3_outputs(7177) <= not a;
    layer3_outputs(7178) <= a;
    layer3_outputs(7179) <= not b or a;
    layer3_outputs(7180) <= not (a xor b);
    layer3_outputs(7181) <= not (a and b);
    layer3_outputs(7182) <= '0';
    layer3_outputs(7183) <= not b;
    layer3_outputs(7184) <= not (a and b);
    layer3_outputs(7185) <= b and not a;
    layer3_outputs(7186) <= a xor b;
    layer3_outputs(7187) <= not (a or b);
    layer3_outputs(7188) <= '0';
    layer3_outputs(7189) <= b and not a;
    layer3_outputs(7190) <= a and not b;
    layer3_outputs(7191) <= '0';
    layer3_outputs(7192) <= '1';
    layer3_outputs(7193) <= not a;
    layer3_outputs(7194) <= '0';
    layer3_outputs(7195) <= not a;
    layer3_outputs(7196) <= '0';
    layer3_outputs(7197) <= not a;
    layer3_outputs(7198) <= not a;
    layer3_outputs(7199) <= not b;
    layer3_outputs(7200) <= a or b;
    layer3_outputs(7201) <= a;
    layer3_outputs(7202) <= not (a or b);
    layer3_outputs(7203) <= a;
    layer3_outputs(7204) <= not a or b;
    layer3_outputs(7205) <= not a or b;
    layer3_outputs(7206) <= '0';
    layer3_outputs(7207) <= not a or b;
    layer3_outputs(7208) <= not (a and b);
    layer3_outputs(7209) <= a and not b;
    layer3_outputs(7210) <= '0';
    layer3_outputs(7211) <= a;
    layer3_outputs(7212) <= b and not a;
    layer3_outputs(7213) <= a or b;
    layer3_outputs(7214) <= not a;
    layer3_outputs(7215) <= a or b;
    layer3_outputs(7216) <= not (a or b);
    layer3_outputs(7217) <= a;
    layer3_outputs(7218) <= not b;
    layer3_outputs(7219) <= a;
    layer3_outputs(7220) <= '1';
    layer3_outputs(7221) <= b and not a;
    layer3_outputs(7222) <= a;
    layer3_outputs(7223) <= not a or b;
    layer3_outputs(7224) <= not a;
    layer3_outputs(7225) <= not a or b;
    layer3_outputs(7226) <= not a;
    layer3_outputs(7227) <= a and not b;
    layer3_outputs(7228) <= not a;
    layer3_outputs(7229) <= not b;
    layer3_outputs(7230) <= not (a and b);
    layer3_outputs(7231) <= a and b;
    layer3_outputs(7232) <= not a or b;
    layer3_outputs(7233) <= not a;
    layer3_outputs(7234) <= a and b;
    layer3_outputs(7235) <= a xor b;
    layer3_outputs(7236) <= not (a and b);
    layer3_outputs(7237) <= not b;
    layer3_outputs(7238) <= a;
    layer3_outputs(7239) <= a and b;
    layer3_outputs(7240) <= not b;
    layer3_outputs(7241) <= '1';
    layer3_outputs(7242) <= not a;
    layer3_outputs(7243) <= not (a xor b);
    layer3_outputs(7244) <= b;
    layer3_outputs(7245) <= a and not b;
    layer3_outputs(7246) <= b;
    layer3_outputs(7247) <= not b or a;
    layer3_outputs(7248) <= a and b;
    layer3_outputs(7249) <= '0';
    layer3_outputs(7250) <= a and not b;
    layer3_outputs(7251) <= a or b;
    layer3_outputs(7252) <= a and not b;
    layer3_outputs(7253) <= not b;
    layer3_outputs(7254) <= not (a or b);
    layer3_outputs(7255) <= a;
    layer3_outputs(7256) <= not (a or b);
    layer3_outputs(7257) <= not (a or b);
    layer3_outputs(7258) <= not (a or b);
    layer3_outputs(7259) <= not a;
    layer3_outputs(7260) <= not b or a;
    layer3_outputs(7261) <= not (a xor b);
    layer3_outputs(7262) <= a;
    layer3_outputs(7263) <= not (a and b);
    layer3_outputs(7264) <= not b or a;
    layer3_outputs(7265) <= '1';
    layer3_outputs(7266) <= not b or a;
    layer3_outputs(7267) <= not a;
    layer3_outputs(7268) <= a and b;
    layer3_outputs(7269) <= not b;
    layer3_outputs(7270) <= not b or a;
    layer3_outputs(7271) <= a and not b;
    layer3_outputs(7272) <= not a;
    layer3_outputs(7273) <= '0';
    layer3_outputs(7274) <= a xor b;
    layer3_outputs(7275) <= a and not b;
    layer3_outputs(7276) <= '0';
    layer3_outputs(7277) <= not (a xor b);
    layer3_outputs(7278) <= not b or a;
    layer3_outputs(7279) <= '0';
    layer3_outputs(7280) <= a and not b;
    layer3_outputs(7281) <= not a or b;
    layer3_outputs(7282) <= not a;
    layer3_outputs(7283) <= not (a or b);
    layer3_outputs(7284) <= b;
    layer3_outputs(7285) <= not a;
    layer3_outputs(7286) <= '0';
    layer3_outputs(7287) <= a or b;
    layer3_outputs(7288) <= b;
    layer3_outputs(7289) <= not a or b;
    layer3_outputs(7290) <= b and not a;
    layer3_outputs(7291) <= not (a and b);
    layer3_outputs(7292) <= b;
    layer3_outputs(7293) <= a or b;
    layer3_outputs(7294) <= a xor b;
    layer3_outputs(7295) <= a or b;
    layer3_outputs(7296) <= not a;
    layer3_outputs(7297) <= not b or a;
    layer3_outputs(7298) <= a and not b;
    layer3_outputs(7299) <= a;
    layer3_outputs(7300) <= a;
    layer3_outputs(7301) <= not (a and b);
    layer3_outputs(7302) <= not a;
    layer3_outputs(7303) <= not (a and b);
    layer3_outputs(7304) <= b and not a;
    layer3_outputs(7305) <= '1';
    layer3_outputs(7306) <= not (a xor b);
    layer3_outputs(7307) <= not (a and b);
    layer3_outputs(7308) <= not b or a;
    layer3_outputs(7309) <= not b;
    layer3_outputs(7310) <= b;
    layer3_outputs(7311) <= not b;
    layer3_outputs(7312) <= not a;
    layer3_outputs(7313) <= not a;
    layer3_outputs(7314) <= a;
    layer3_outputs(7315) <= a;
    layer3_outputs(7316) <= b;
    layer3_outputs(7317) <= a;
    layer3_outputs(7318) <= b;
    layer3_outputs(7319) <= a;
    layer3_outputs(7320) <= not b;
    layer3_outputs(7321) <= '0';
    layer3_outputs(7322) <= not a;
    layer3_outputs(7323) <= not a or b;
    layer3_outputs(7324) <= b;
    layer3_outputs(7325) <= a;
    layer3_outputs(7326) <= b;
    layer3_outputs(7327) <= a;
    layer3_outputs(7328) <= not a or b;
    layer3_outputs(7329) <= not a or b;
    layer3_outputs(7330) <= a xor b;
    layer3_outputs(7331) <= a and b;
    layer3_outputs(7332) <= not (a xor b);
    layer3_outputs(7333) <= b;
    layer3_outputs(7334) <= a or b;
    layer3_outputs(7335) <= a or b;
    layer3_outputs(7336) <= a xor b;
    layer3_outputs(7337) <= a and b;
    layer3_outputs(7338) <= not (a xor b);
    layer3_outputs(7339) <= not (a and b);
    layer3_outputs(7340) <= not (a and b);
    layer3_outputs(7341) <= not (a xor b);
    layer3_outputs(7342) <= b;
    layer3_outputs(7343) <= not (a or b);
    layer3_outputs(7344) <= a;
    layer3_outputs(7345) <= a;
    layer3_outputs(7346) <= a;
    layer3_outputs(7347) <= not (a and b);
    layer3_outputs(7348) <= a and b;
    layer3_outputs(7349) <= not (a or b);
    layer3_outputs(7350) <= a and b;
    layer3_outputs(7351) <= not (a and b);
    layer3_outputs(7352) <= not a;
    layer3_outputs(7353) <= b;
    layer3_outputs(7354) <= not a or b;
    layer3_outputs(7355) <= b;
    layer3_outputs(7356) <= b;
    layer3_outputs(7357) <= b;
    layer3_outputs(7358) <= b and not a;
    layer3_outputs(7359) <= not b;
    layer3_outputs(7360) <= '1';
    layer3_outputs(7361) <= not b or a;
    layer3_outputs(7362) <= not b or a;
    layer3_outputs(7363) <= not a or b;
    layer3_outputs(7364) <= not b;
    layer3_outputs(7365) <= a or b;
    layer3_outputs(7366) <= not (a or b);
    layer3_outputs(7367) <= not b;
    layer3_outputs(7368) <= '1';
    layer3_outputs(7369) <= a;
    layer3_outputs(7370) <= a xor b;
    layer3_outputs(7371) <= not a;
    layer3_outputs(7372) <= b and not a;
    layer3_outputs(7373) <= '1';
    layer3_outputs(7374) <= b;
    layer3_outputs(7375) <= not (a xor b);
    layer3_outputs(7376) <= a;
    layer3_outputs(7377) <= not a;
    layer3_outputs(7378) <= a;
    layer3_outputs(7379) <= not b;
    layer3_outputs(7380) <= not (a xor b);
    layer3_outputs(7381) <= a or b;
    layer3_outputs(7382) <= a and b;
    layer3_outputs(7383) <= a and b;
    layer3_outputs(7384) <= not a or b;
    layer3_outputs(7385) <= not (a or b);
    layer3_outputs(7386) <= '1';
    layer3_outputs(7387) <= a;
    layer3_outputs(7388) <= not a;
    layer3_outputs(7389) <= a or b;
    layer3_outputs(7390) <= b;
    layer3_outputs(7391) <= a;
    layer3_outputs(7392) <= not b;
    layer3_outputs(7393) <= b and not a;
    layer3_outputs(7394) <= '0';
    layer3_outputs(7395) <= not b or a;
    layer3_outputs(7396) <= not (a or b);
    layer3_outputs(7397) <= not a;
    layer3_outputs(7398) <= a;
    layer3_outputs(7399) <= a;
    layer3_outputs(7400) <= b and not a;
    layer3_outputs(7401) <= a;
    layer3_outputs(7402) <= not (a and b);
    layer3_outputs(7403) <= a and not b;
    layer3_outputs(7404) <= a;
    layer3_outputs(7405) <= not a;
    layer3_outputs(7406) <= not (a and b);
    layer3_outputs(7407) <= b;
    layer3_outputs(7408) <= b and not a;
    layer3_outputs(7409) <= b and not a;
    layer3_outputs(7410) <= a;
    layer3_outputs(7411) <= b;
    layer3_outputs(7412) <= a and not b;
    layer3_outputs(7413) <= '0';
    layer3_outputs(7414) <= not a or b;
    layer3_outputs(7415) <= not b;
    layer3_outputs(7416) <= a or b;
    layer3_outputs(7417) <= not (a or b);
    layer3_outputs(7418) <= a and b;
    layer3_outputs(7419) <= a or b;
    layer3_outputs(7420) <= a and not b;
    layer3_outputs(7421) <= not (a or b);
    layer3_outputs(7422) <= not a;
    layer3_outputs(7423) <= b and not a;
    layer3_outputs(7424) <= not b or a;
    layer3_outputs(7425) <= b and not a;
    layer3_outputs(7426) <= not a or b;
    layer3_outputs(7427) <= not b;
    layer3_outputs(7428) <= not (a or b);
    layer3_outputs(7429) <= not (a xor b);
    layer3_outputs(7430) <= b;
    layer3_outputs(7431) <= not (a xor b);
    layer3_outputs(7432) <= not a;
    layer3_outputs(7433) <= not (a or b);
    layer3_outputs(7434) <= not a;
    layer3_outputs(7435) <= a;
    layer3_outputs(7436) <= not (a and b);
    layer3_outputs(7437) <= not a or b;
    layer3_outputs(7438) <= not b or a;
    layer3_outputs(7439) <= not a;
    layer3_outputs(7440) <= not b;
    layer3_outputs(7441) <= not a;
    layer3_outputs(7442) <= not (a xor b);
    layer3_outputs(7443) <= a or b;
    layer3_outputs(7444) <= b and not a;
    layer3_outputs(7445) <= not (a xor b);
    layer3_outputs(7446) <= a;
    layer3_outputs(7447) <= not b or a;
    layer3_outputs(7448) <= a and not b;
    layer3_outputs(7449) <= a or b;
    layer3_outputs(7450) <= b;
    layer3_outputs(7451) <= not (a or b);
    layer3_outputs(7452) <= a or b;
    layer3_outputs(7453) <= '1';
    layer3_outputs(7454) <= b and not a;
    layer3_outputs(7455) <= a and b;
    layer3_outputs(7456) <= a or b;
    layer3_outputs(7457) <= not a or b;
    layer3_outputs(7458) <= a and not b;
    layer3_outputs(7459) <= not (a and b);
    layer3_outputs(7460) <= not b or a;
    layer3_outputs(7461) <= a and not b;
    layer3_outputs(7462) <= a xor b;
    layer3_outputs(7463) <= not a;
    layer3_outputs(7464) <= a;
    layer3_outputs(7465) <= a xor b;
    layer3_outputs(7466) <= not b or a;
    layer3_outputs(7467) <= not b or a;
    layer3_outputs(7468) <= a and not b;
    layer3_outputs(7469) <= not b;
    layer3_outputs(7470) <= a and b;
    layer3_outputs(7471) <= b;
    layer3_outputs(7472) <= '0';
    layer3_outputs(7473) <= not b;
    layer3_outputs(7474) <= not b or a;
    layer3_outputs(7475) <= not a;
    layer3_outputs(7476) <= b;
    layer3_outputs(7477) <= not a or b;
    layer3_outputs(7478) <= not a or b;
    layer3_outputs(7479) <= not b;
    layer3_outputs(7480) <= a and not b;
    layer3_outputs(7481) <= a or b;
    layer3_outputs(7482) <= a and b;
    layer3_outputs(7483) <= a and b;
    layer3_outputs(7484) <= b;
    layer3_outputs(7485) <= not a or b;
    layer3_outputs(7486) <= a;
    layer3_outputs(7487) <= not (a and b);
    layer3_outputs(7488) <= a xor b;
    layer3_outputs(7489) <= a or b;
    layer3_outputs(7490) <= not (a or b);
    layer3_outputs(7491) <= a and b;
    layer3_outputs(7492) <= a;
    layer3_outputs(7493) <= a;
    layer3_outputs(7494) <= b;
    layer3_outputs(7495) <= not a or b;
    layer3_outputs(7496) <= a;
    layer3_outputs(7497) <= not (a and b);
    layer3_outputs(7498) <= not b or a;
    layer3_outputs(7499) <= a and not b;
    layer3_outputs(7500) <= a and not b;
    layer3_outputs(7501) <= a or b;
    layer3_outputs(7502) <= not b;
    layer3_outputs(7503) <= not b;
    layer3_outputs(7504) <= a and b;
    layer3_outputs(7505) <= b;
    layer3_outputs(7506) <= '1';
    layer3_outputs(7507) <= a and not b;
    layer3_outputs(7508) <= a and b;
    layer3_outputs(7509) <= a and not b;
    layer3_outputs(7510) <= b;
    layer3_outputs(7511) <= not b;
    layer3_outputs(7512) <= not b;
    layer3_outputs(7513) <= not (a or b);
    layer3_outputs(7514) <= b and not a;
    layer3_outputs(7515) <= b and not a;
    layer3_outputs(7516) <= a;
    layer3_outputs(7517) <= a;
    layer3_outputs(7518) <= not (a xor b);
    layer3_outputs(7519) <= not (a or b);
    layer3_outputs(7520) <= '1';
    layer3_outputs(7521) <= not a;
    layer3_outputs(7522) <= not (a or b);
    layer3_outputs(7523) <= a xor b;
    layer3_outputs(7524) <= a xor b;
    layer3_outputs(7525) <= not b or a;
    layer3_outputs(7526) <= b;
    layer3_outputs(7527) <= not a or b;
    layer3_outputs(7528) <= not b;
    layer3_outputs(7529) <= not (a or b);
    layer3_outputs(7530) <= a or b;
    layer3_outputs(7531) <= a;
    layer3_outputs(7532) <= a;
    layer3_outputs(7533) <= not a;
    layer3_outputs(7534) <= b;
    layer3_outputs(7535) <= b;
    layer3_outputs(7536) <= '0';
    layer3_outputs(7537) <= '0';
    layer3_outputs(7538) <= not b or a;
    layer3_outputs(7539) <= not a;
    layer3_outputs(7540) <= a;
    layer3_outputs(7541) <= not a;
    layer3_outputs(7542) <= a or b;
    layer3_outputs(7543) <= a and b;
    layer3_outputs(7544) <= b;
    layer3_outputs(7545) <= not b or a;
    layer3_outputs(7546) <= b;
    layer3_outputs(7547) <= b;
    layer3_outputs(7548) <= b and not a;
    layer3_outputs(7549) <= '0';
    layer3_outputs(7550) <= b;
    layer3_outputs(7551) <= not a;
    layer3_outputs(7552) <= a and b;
    layer3_outputs(7553) <= a and b;
    layer3_outputs(7554) <= a xor b;
    layer3_outputs(7555) <= a and not b;
    layer3_outputs(7556) <= not b or a;
    layer3_outputs(7557) <= not (a xor b);
    layer3_outputs(7558) <= b;
    layer3_outputs(7559) <= not a or b;
    layer3_outputs(7560) <= a xor b;
    layer3_outputs(7561) <= not b;
    layer3_outputs(7562) <= not a or b;
    layer3_outputs(7563) <= a or b;
    layer3_outputs(7564) <= b and not a;
    layer3_outputs(7565) <= a;
    layer3_outputs(7566) <= not (a or b);
    layer3_outputs(7567) <= not a;
    layer3_outputs(7568) <= not (a or b);
    layer3_outputs(7569) <= a or b;
    layer3_outputs(7570) <= not b;
    layer3_outputs(7571) <= b and not a;
    layer3_outputs(7572) <= not b;
    layer3_outputs(7573) <= not (a xor b);
    layer3_outputs(7574) <= a and b;
    layer3_outputs(7575) <= a;
    layer3_outputs(7576) <= not (a or b);
    layer3_outputs(7577) <= not a;
    layer3_outputs(7578) <= a and b;
    layer3_outputs(7579) <= b and not a;
    layer3_outputs(7580) <= a or b;
    layer3_outputs(7581) <= not a or b;
    layer3_outputs(7582) <= not (a and b);
    layer3_outputs(7583) <= a;
    layer3_outputs(7584) <= not b;
    layer3_outputs(7585) <= a and not b;
    layer3_outputs(7586) <= not (a or b);
    layer3_outputs(7587) <= not a;
    layer3_outputs(7588) <= b;
    layer3_outputs(7589) <= a;
    layer3_outputs(7590) <= a or b;
    layer3_outputs(7591) <= not b;
    layer3_outputs(7592) <= not (a xor b);
    layer3_outputs(7593) <= a xor b;
    layer3_outputs(7594) <= not a;
    layer3_outputs(7595) <= not (a xor b);
    layer3_outputs(7596) <= a and b;
    layer3_outputs(7597) <= not (a or b);
    layer3_outputs(7598) <= '0';
    layer3_outputs(7599) <= b;
    layer3_outputs(7600) <= not (a or b);
    layer3_outputs(7601) <= not b or a;
    layer3_outputs(7602) <= b;
    layer3_outputs(7603) <= b;
    layer3_outputs(7604) <= not b or a;
    layer3_outputs(7605) <= a;
    layer3_outputs(7606) <= a and b;
    layer3_outputs(7607) <= a and b;
    layer3_outputs(7608) <= not b or a;
    layer3_outputs(7609) <= a;
    layer3_outputs(7610) <= not b;
    layer3_outputs(7611) <= not b or a;
    layer3_outputs(7612) <= a and b;
    layer3_outputs(7613) <= b;
    layer3_outputs(7614) <= a or b;
    layer3_outputs(7615) <= a xor b;
    layer3_outputs(7616) <= not (a and b);
    layer3_outputs(7617) <= a;
    layer3_outputs(7618) <= a and b;
    layer3_outputs(7619) <= '1';
    layer3_outputs(7620) <= not b or a;
    layer3_outputs(7621) <= not (a and b);
    layer3_outputs(7622) <= not (a and b);
    layer3_outputs(7623) <= not b;
    layer3_outputs(7624) <= a and not b;
    layer3_outputs(7625) <= '0';
    layer3_outputs(7626) <= not (a and b);
    layer3_outputs(7627) <= not (a xor b);
    layer3_outputs(7628) <= not (a and b);
    layer3_outputs(7629) <= '1';
    layer3_outputs(7630) <= not b;
    layer3_outputs(7631) <= not a;
    layer3_outputs(7632) <= not b;
    layer3_outputs(7633) <= not b;
    layer3_outputs(7634) <= not (a and b);
    layer3_outputs(7635) <= not a;
    layer3_outputs(7636) <= not b;
    layer3_outputs(7637) <= a and not b;
    layer3_outputs(7638) <= '0';
    layer3_outputs(7639) <= b and not a;
    layer3_outputs(7640) <= not (a xor b);
    layer3_outputs(7641) <= '1';
    layer3_outputs(7642) <= not b;
    layer3_outputs(7643) <= a and b;
    layer3_outputs(7644) <= '1';
    layer3_outputs(7645) <= a and not b;
    layer3_outputs(7646) <= not b;
    layer3_outputs(7647) <= a or b;
    layer3_outputs(7648) <= not (a or b);
    layer3_outputs(7649) <= a and not b;
    layer3_outputs(7650) <= a;
    layer3_outputs(7651) <= not a;
    layer3_outputs(7652) <= b;
    layer3_outputs(7653) <= not a or b;
    layer3_outputs(7654) <= '0';
    layer3_outputs(7655) <= a and not b;
    layer3_outputs(7656) <= a and not b;
    layer3_outputs(7657) <= '1';
    layer3_outputs(7658) <= b and not a;
    layer3_outputs(7659) <= not (a or b);
    layer3_outputs(7660) <= not (a and b);
    layer3_outputs(7661) <= not (a or b);
    layer3_outputs(7662) <= not (a xor b);
    layer3_outputs(7663) <= not (a and b);
    layer3_outputs(7664) <= b and not a;
    layer3_outputs(7665) <= b;
    layer3_outputs(7666) <= not a;
    layer3_outputs(7667) <= not b;
    layer3_outputs(7668) <= not b or a;
    layer3_outputs(7669) <= a xor b;
    layer3_outputs(7670) <= not (a or b);
    layer3_outputs(7671) <= b;
    layer3_outputs(7672) <= a;
    layer3_outputs(7673) <= not (a and b);
    layer3_outputs(7674) <= not a or b;
    layer3_outputs(7675) <= not a or b;
    layer3_outputs(7676) <= a xor b;
    layer3_outputs(7677) <= a and b;
    layer3_outputs(7678) <= not a;
    layer3_outputs(7679) <= b and not a;
    layer3_outputs(7680) <= '1';
    layer3_outputs(7681) <= not b;
    layer3_outputs(7682) <= '0';
    layer3_outputs(7683) <= a;
    layer3_outputs(7684) <= not b;
    layer3_outputs(7685) <= not (a and b);
    layer3_outputs(7686) <= not a;
    layer3_outputs(7687) <= not a;
    layer3_outputs(7688) <= a and not b;
    layer3_outputs(7689) <= not (a xor b);
    layer3_outputs(7690) <= b and not a;
    layer3_outputs(7691) <= not a;
    layer3_outputs(7692) <= not b or a;
    layer3_outputs(7693) <= a;
    layer3_outputs(7694) <= not (a xor b);
    layer3_outputs(7695) <= '1';
    layer3_outputs(7696) <= not a or b;
    layer3_outputs(7697) <= a and not b;
    layer3_outputs(7698) <= not a;
    layer3_outputs(7699) <= a;
    layer3_outputs(7700) <= '1';
    layer3_outputs(7701) <= a;
    layer3_outputs(7702) <= a;
    layer3_outputs(7703) <= b;
    layer3_outputs(7704) <= not a or b;
    layer3_outputs(7705) <= not b or a;
    layer3_outputs(7706) <= not b;
    layer3_outputs(7707) <= b;
    layer3_outputs(7708) <= not b or a;
    layer3_outputs(7709) <= a and b;
    layer3_outputs(7710) <= not a;
    layer3_outputs(7711) <= a;
    layer3_outputs(7712) <= a xor b;
    layer3_outputs(7713) <= a or b;
    layer3_outputs(7714) <= a;
    layer3_outputs(7715) <= not b;
    layer3_outputs(7716) <= a and b;
    layer3_outputs(7717) <= b and not a;
    layer3_outputs(7718) <= b and not a;
    layer3_outputs(7719) <= not a;
    layer3_outputs(7720) <= a and b;
    layer3_outputs(7721) <= not a;
    layer3_outputs(7722) <= not (a and b);
    layer3_outputs(7723) <= b;
    layer3_outputs(7724) <= a or b;
    layer3_outputs(7725) <= '0';
    layer3_outputs(7726) <= not a or b;
    layer3_outputs(7727) <= b;
    layer3_outputs(7728) <= b and not a;
    layer3_outputs(7729) <= not b or a;
    layer3_outputs(7730) <= not a;
    layer3_outputs(7731) <= not a;
    layer3_outputs(7732) <= a;
    layer3_outputs(7733) <= '1';
    layer3_outputs(7734) <= not b;
    layer3_outputs(7735) <= not b;
    layer3_outputs(7736) <= not b or a;
    layer3_outputs(7737) <= not b or a;
    layer3_outputs(7738) <= '1';
    layer3_outputs(7739) <= not a or b;
    layer3_outputs(7740) <= not (a or b);
    layer3_outputs(7741) <= '1';
    layer3_outputs(7742) <= a;
    layer3_outputs(7743) <= a or b;
    layer3_outputs(7744) <= not (a or b);
    layer3_outputs(7745) <= not (a or b);
    layer3_outputs(7746) <= a or b;
    layer3_outputs(7747) <= a and not b;
    layer3_outputs(7748) <= a xor b;
    layer3_outputs(7749) <= b and not a;
    layer3_outputs(7750) <= not b;
    layer3_outputs(7751) <= not b;
    layer3_outputs(7752) <= not a;
    layer3_outputs(7753) <= not (a xor b);
    layer3_outputs(7754) <= not b or a;
    layer3_outputs(7755) <= not a;
    layer3_outputs(7756) <= not a;
    layer3_outputs(7757) <= b;
    layer3_outputs(7758) <= b;
    layer3_outputs(7759) <= not b;
    layer3_outputs(7760) <= '1';
    layer3_outputs(7761) <= a xor b;
    layer3_outputs(7762) <= not a;
    layer3_outputs(7763) <= not (a or b);
    layer3_outputs(7764) <= not b;
    layer3_outputs(7765) <= a;
    layer3_outputs(7766) <= '1';
    layer3_outputs(7767) <= b;
    layer3_outputs(7768) <= a or b;
    layer3_outputs(7769) <= a;
    layer3_outputs(7770) <= not a;
    layer3_outputs(7771) <= a;
    layer3_outputs(7772) <= not b or a;
    layer3_outputs(7773) <= a;
    layer3_outputs(7774) <= not a or b;
    layer3_outputs(7775) <= not b;
    layer3_outputs(7776) <= not b;
    layer3_outputs(7777) <= not (a xor b);
    layer3_outputs(7778) <= not b;
    layer3_outputs(7779) <= not (a and b);
    layer3_outputs(7780) <= b and not a;
    layer3_outputs(7781) <= a;
    layer3_outputs(7782) <= a and b;
    layer3_outputs(7783) <= b and not a;
    layer3_outputs(7784) <= not (a or b);
    layer3_outputs(7785) <= not (a xor b);
    layer3_outputs(7786) <= a;
    layer3_outputs(7787) <= not (a xor b);
    layer3_outputs(7788) <= not b or a;
    layer3_outputs(7789) <= not a or b;
    layer3_outputs(7790) <= not a;
    layer3_outputs(7791) <= a or b;
    layer3_outputs(7792) <= not (a xor b);
    layer3_outputs(7793) <= a;
    layer3_outputs(7794) <= not a or b;
    layer3_outputs(7795) <= a and not b;
    layer3_outputs(7796) <= not (a or b);
    layer3_outputs(7797) <= a and not b;
    layer3_outputs(7798) <= not a or b;
    layer3_outputs(7799) <= not (a and b);
    layer3_outputs(7800) <= b;
    layer3_outputs(7801) <= not b or a;
    layer3_outputs(7802) <= a xor b;
    layer3_outputs(7803) <= a or b;
    layer3_outputs(7804) <= not a;
    layer3_outputs(7805) <= b and not a;
    layer3_outputs(7806) <= '1';
    layer3_outputs(7807) <= a and b;
    layer3_outputs(7808) <= b;
    layer3_outputs(7809) <= '1';
    layer3_outputs(7810) <= a and b;
    layer3_outputs(7811) <= not b;
    layer3_outputs(7812) <= a;
    layer3_outputs(7813) <= b;
    layer3_outputs(7814) <= b;
    layer3_outputs(7815) <= not (a xor b);
    layer3_outputs(7816) <= not (a or b);
    layer3_outputs(7817) <= a and not b;
    layer3_outputs(7818) <= not (a xor b);
    layer3_outputs(7819) <= a;
    layer3_outputs(7820) <= not (a xor b);
    layer3_outputs(7821) <= b;
    layer3_outputs(7822) <= b and not a;
    layer3_outputs(7823) <= b;
    layer3_outputs(7824) <= a and not b;
    layer3_outputs(7825) <= not (a and b);
    layer3_outputs(7826) <= not (a or b);
    layer3_outputs(7827) <= b and not a;
    layer3_outputs(7828) <= not b;
    layer3_outputs(7829) <= not b;
    layer3_outputs(7830) <= not (a or b);
    layer3_outputs(7831) <= '0';
    layer3_outputs(7832) <= '1';
    layer3_outputs(7833) <= a;
    layer3_outputs(7834) <= not a;
    layer3_outputs(7835) <= a and b;
    layer3_outputs(7836) <= not a or b;
    layer3_outputs(7837) <= not (a and b);
    layer3_outputs(7838) <= a xor b;
    layer3_outputs(7839) <= b;
    layer3_outputs(7840) <= a and b;
    layer3_outputs(7841) <= not b;
    layer3_outputs(7842) <= a or b;
    layer3_outputs(7843) <= a or b;
    layer3_outputs(7844) <= b;
    layer3_outputs(7845) <= '0';
    layer3_outputs(7846) <= not b or a;
    layer3_outputs(7847) <= not b;
    layer3_outputs(7848) <= a and b;
    layer3_outputs(7849) <= not b;
    layer3_outputs(7850) <= a xor b;
    layer3_outputs(7851) <= not (a and b);
    layer3_outputs(7852) <= b and not a;
    layer3_outputs(7853) <= a or b;
    layer3_outputs(7854) <= a or b;
    layer3_outputs(7855) <= b and not a;
    layer3_outputs(7856) <= a;
    layer3_outputs(7857) <= a;
    layer3_outputs(7858) <= a;
    layer3_outputs(7859) <= not (a or b);
    layer3_outputs(7860) <= a;
    layer3_outputs(7861) <= not b or a;
    layer3_outputs(7862) <= a;
    layer3_outputs(7863) <= not a;
    layer3_outputs(7864) <= b;
    layer3_outputs(7865) <= not b;
    layer3_outputs(7866) <= b and not a;
    layer3_outputs(7867) <= not a;
    layer3_outputs(7868) <= not a;
    layer3_outputs(7869) <= a;
    layer3_outputs(7870) <= '0';
    layer3_outputs(7871) <= a;
    layer3_outputs(7872) <= not (a and b);
    layer3_outputs(7873) <= not (a and b);
    layer3_outputs(7874) <= a and not b;
    layer3_outputs(7875) <= not a;
    layer3_outputs(7876) <= not (a and b);
    layer3_outputs(7877) <= not b or a;
    layer3_outputs(7878) <= a or b;
    layer3_outputs(7879) <= not b;
    layer3_outputs(7880) <= a xor b;
    layer3_outputs(7881) <= '1';
    layer3_outputs(7882) <= a and b;
    layer3_outputs(7883) <= not a or b;
    layer3_outputs(7884) <= not b or a;
    layer3_outputs(7885) <= not b;
    layer3_outputs(7886) <= not (a and b);
    layer3_outputs(7887) <= a;
    layer3_outputs(7888) <= a;
    layer3_outputs(7889) <= a and not b;
    layer3_outputs(7890) <= not (a and b);
    layer3_outputs(7891) <= not (a or b);
    layer3_outputs(7892) <= b;
    layer3_outputs(7893) <= a and b;
    layer3_outputs(7894) <= b;
    layer3_outputs(7895) <= not a;
    layer3_outputs(7896) <= not a or b;
    layer3_outputs(7897) <= not (a xor b);
    layer3_outputs(7898) <= a and not b;
    layer3_outputs(7899) <= '0';
    layer3_outputs(7900) <= b and not a;
    layer3_outputs(7901) <= not b;
    layer3_outputs(7902) <= not (a and b);
    layer3_outputs(7903) <= not b;
    layer3_outputs(7904) <= a;
    layer3_outputs(7905) <= not a;
    layer3_outputs(7906) <= b;
    layer3_outputs(7907) <= b;
    layer3_outputs(7908) <= b;
    layer3_outputs(7909) <= not b;
    layer3_outputs(7910) <= a xor b;
    layer3_outputs(7911) <= not (a and b);
    layer3_outputs(7912) <= not a;
    layer3_outputs(7913) <= a or b;
    layer3_outputs(7914) <= b and not a;
    layer3_outputs(7915) <= a;
    layer3_outputs(7916) <= not a;
    layer3_outputs(7917) <= not (a xor b);
    layer3_outputs(7918) <= a and b;
    layer3_outputs(7919) <= not (a xor b);
    layer3_outputs(7920) <= not a;
    layer3_outputs(7921) <= not b or a;
    layer3_outputs(7922) <= not (a or b);
    layer3_outputs(7923) <= a xor b;
    layer3_outputs(7924) <= b and not a;
    layer3_outputs(7925) <= a and not b;
    layer3_outputs(7926) <= '0';
    layer3_outputs(7927) <= not a;
    layer3_outputs(7928) <= not (a and b);
    layer3_outputs(7929) <= a and not b;
    layer3_outputs(7930) <= a;
    layer3_outputs(7931) <= not b;
    layer3_outputs(7932) <= b;
    layer3_outputs(7933) <= a and b;
    layer3_outputs(7934) <= '1';
    layer3_outputs(7935) <= a and not b;
    layer3_outputs(7936) <= not b or a;
    layer3_outputs(7937) <= a or b;
    layer3_outputs(7938) <= a;
    layer3_outputs(7939) <= a;
    layer3_outputs(7940) <= not b;
    layer3_outputs(7941) <= not b;
    layer3_outputs(7942) <= '0';
    layer3_outputs(7943) <= b;
    layer3_outputs(7944) <= not b;
    layer3_outputs(7945) <= a;
    layer3_outputs(7946) <= b and not a;
    layer3_outputs(7947) <= a and not b;
    layer3_outputs(7948) <= a and b;
    layer3_outputs(7949) <= a xor b;
    layer3_outputs(7950) <= b;
    layer3_outputs(7951) <= not (a xor b);
    layer3_outputs(7952) <= '1';
    layer3_outputs(7953) <= a and b;
    layer3_outputs(7954) <= not (a xor b);
    layer3_outputs(7955) <= not b or a;
    layer3_outputs(7956) <= not a;
    layer3_outputs(7957) <= a or b;
    layer3_outputs(7958) <= not a;
    layer3_outputs(7959) <= b;
    layer3_outputs(7960) <= not (a and b);
    layer3_outputs(7961) <= b;
    layer3_outputs(7962) <= not b;
    layer3_outputs(7963) <= a;
    layer3_outputs(7964) <= b;
    layer3_outputs(7965) <= a and b;
    layer3_outputs(7966) <= a or b;
    layer3_outputs(7967) <= b;
    layer3_outputs(7968) <= a;
    layer3_outputs(7969) <= not (a xor b);
    layer3_outputs(7970) <= b;
    layer3_outputs(7971) <= not (a and b);
    layer3_outputs(7972) <= a and not b;
    layer3_outputs(7973) <= '0';
    layer3_outputs(7974) <= not a;
    layer3_outputs(7975) <= not a;
    layer3_outputs(7976) <= not b;
    layer3_outputs(7977) <= a;
    layer3_outputs(7978) <= a and not b;
    layer3_outputs(7979) <= not (a xor b);
    layer3_outputs(7980) <= not b;
    layer3_outputs(7981) <= not b;
    layer3_outputs(7982) <= a and b;
    layer3_outputs(7983) <= not (a and b);
    layer3_outputs(7984) <= b and not a;
    layer3_outputs(7985) <= not (a or b);
    layer3_outputs(7986) <= not (a or b);
    layer3_outputs(7987) <= a xor b;
    layer3_outputs(7988) <= b;
    layer3_outputs(7989) <= not b or a;
    layer3_outputs(7990) <= not (a and b);
    layer3_outputs(7991) <= not b;
    layer3_outputs(7992) <= b and not a;
    layer3_outputs(7993) <= a;
    layer3_outputs(7994) <= not (a or b);
    layer3_outputs(7995) <= a and b;
    layer3_outputs(7996) <= not b or a;
    layer3_outputs(7997) <= not (a or b);
    layer3_outputs(7998) <= not a or b;
    layer3_outputs(7999) <= b and not a;
    layer3_outputs(8000) <= b and not a;
    layer3_outputs(8001) <= not a;
    layer3_outputs(8002) <= not a or b;
    layer3_outputs(8003) <= b and not a;
    layer3_outputs(8004) <= a;
    layer3_outputs(8005) <= not (a or b);
    layer3_outputs(8006) <= not (a or b);
    layer3_outputs(8007) <= a and not b;
    layer3_outputs(8008) <= b;
    layer3_outputs(8009) <= a;
    layer3_outputs(8010) <= not a;
    layer3_outputs(8011) <= not b or a;
    layer3_outputs(8012) <= '0';
    layer3_outputs(8013) <= not a;
    layer3_outputs(8014) <= a;
    layer3_outputs(8015) <= a;
    layer3_outputs(8016) <= not (a xor b);
    layer3_outputs(8017) <= a;
    layer3_outputs(8018) <= not a;
    layer3_outputs(8019) <= not (a xor b);
    layer3_outputs(8020) <= b and not a;
    layer3_outputs(8021) <= not a;
    layer3_outputs(8022) <= not b or a;
    layer3_outputs(8023) <= a and b;
    layer3_outputs(8024) <= a or b;
    layer3_outputs(8025) <= not (a and b);
    layer3_outputs(8026) <= a;
    layer3_outputs(8027) <= not (a and b);
    layer3_outputs(8028) <= a or b;
    layer3_outputs(8029) <= not (a or b);
    layer3_outputs(8030) <= b;
    layer3_outputs(8031) <= b and not a;
    layer3_outputs(8032) <= not b or a;
    layer3_outputs(8033) <= not b;
    layer3_outputs(8034) <= not b;
    layer3_outputs(8035) <= not a or b;
    layer3_outputs(8036) <= a;
    layer3_outputs(8037) <= b;
    layer3_outputs(8038) <= not a;
    layer3_outputs(8039) <= not (a and b);
    layer3_outputs(8040) <= a;
    layer3_outputs(8041) <= b;
    layer3_outputs(8042) <= a;
    layer3_outputs(8043) <= b;
    layer3_outputs(8044) <= not (a or b);
    layer3_outputs(8045) <= not b or a;
    layer3_outputs(8046) <= not a;
    layer3_outputs(8047) <= b;
    layer3_outputs(8048) <= '1';
    layer3_outputs(8049) <= not a or b;
    layer3_outputs(8050) <= a and not b;
    layer3_outputs(8051) <= not (a xor b);
    layer3_outputs(8052) <= '1';
    layer3_outputs(8053) <= a;
    layer3_outputs(8054) <= a;
    layer3_outputs(8055) <= not (a or b);
    layer3_outputs(8056) <= a;
    layer3_outputs(8057) <= not a;
    layer3_outputs(8058) <= not a or b;
    layer3_outputs(8059) <= '0';
    layer3_outputs(8060) <= not (a and b);
    layer3_outputs(8061) <= a and not b;
    layer3_outputs(8062) <= a and not b;
    layer3_outputs(8063) <= b;
    layer3_outputs(8064) <= not (a xor b);
    layer3_outputs(8065) <= b;
    layer3_outputs(8066) <= a or b;
    layer3_outputs(8067) <= not a;
    layer3_outputs(8068) <= not b;
    layer3_outputs(8069) <= b;
    layer3_outputs(8070) <= b;
    layer3_outputs(8071) <= not b;
    layer3_outputs(8072) <= a;
    layer3_outputs(8073) <= not (a xor b);
    layer3_outputs(8074) <= not a;
    layer3_outputs(8075) <= not (a or b);
    layer3_outputs(8076) <= not a or b;
    layer3_outputs(8077) <= '0';
    layer3_outputs(8078) <= a and b;
    layer3_outputs(8079) <= a;
    layer3_outputs(8080) <= b;
    layer3_outputs(8081) <= a and not b;
    layer3_outputs(8082) <= not a;
    layer3_outputs(8083) <= not (a or b);
    layer3_outputs(8084) <= b and not a;
    layer3_outputs(8085) <= a;
    layer3_outputs(8086) <= a and b;
    layer3_outputs(8087) <= not (a or b);
    layer3_outputs(8088) <= a;
    layer3_outputs(8089) <= a;
    layer3_outputs(8090) <= b and not a;
    layer3_outputs(8091) <= a and b;
    layer3_outputs(8092) <= a;
    layer3_outputs(8093) <= a;
    layer3_outputs(8094) <= not b;
    layer3_outputs(8095) <= a and not b;
    layer3_outputs(8096) <= not b or a;
    layer3_outputs(8097) <= b;
    layer3_outputs(8098) <= a;
    layer3_outputs(8099) <= b;
    layer3_outputs(8100) <= not (a or b);
    layer3_outputs(8101) <= not a or b;
    layer3_outputs(8102) <= '0';
    layer3_outputs(8103) <= not (a xor b);
    layer3_outputs(8104) <= a or b;
    layer3_outputs(8105) <= not a or b;
    layer3_outputs(8106) <= not (a or b);
    layer3_outputs(8107) <= not b or a;
    layer3_outputs(8108) <= not b;
    layer3_outputs(8109) <= not b or a;
    layer3_outputs(8110) <= not a or b;
    layer3_outputs(8111) <= b;
    layer3_outputs(8112) <= a and b;
    layer3_outputs(8113) <= b;
    layer3_outputs(8114) <= a and not b;
    layer3_outputs(8115) <= not b;
    layer3_outputs(8116) <= a and b;
    layer3_outputs(8117) <= a and not b;
    layer3_outputs(8118) <= a and not b;
    layer3_outputs(8119) <= not b;
    layer3_outputs(8120) <= a or b;
    layer3_outputs(8121) <= b;
    layer3_outputs(8122) <= not (a xor b);
    layer3_outputs(8123) <= a or b;
    layer3_outputs(8124) <= not (a and b);
    layer3_outputs(8125) <= not b or a;
    layer3_outputs(8126) <= a;
    layer3_outputs(8127) <= not b or a;
    layer3_outputs(8128) <= b;
    layer3_outputs(8129) <= not (a and b);
    layer3_outputs(8130) <= a and not b;
    layer3_outputs(8131) <= a and not b;
    layer3_outputs(8132) <= a or b;
    layer3_outputs(8133) <= '0';
    layer3_outputs(8134) <= not a;
    layer3_outputs(8135) <= not (a or b);
    layer3_outputs(8136) <= '1';
    layer3_outputs(8137) <= a;
    layer3_outputs(8138) <= '1';
    layer3_outputs(8139) <= a and b;
    layer3_outputs(8140) <= not a;
    layer3_outputs(8141) <= a xor b;
    layer3_outputs(8142) <= b;
    layer3_outputs(8143) <= not a or b;
    layer3_outputs(8144) <= not b or a;
    layer3_outputs(8145) <= b;
    layer3_outputs(8146) <= not b;
    layer3_outputs(8147) <= not (a or b);
    layer3_outputs(8148) <= not a or b;
    layer3_outputs(8149) <= b and not a;
    layer3_outputs(8150) <= not (a xor b);
    layer3_outputs(8151) <= a and not b;
    layer3_outputs(8152) <= a;
    layer3_outputs(8153) <= a and b;
    layer3_outputs(8154) <= not (a xor b);
    layer3_outputs(8155) <= a and not b;
    layer3_outputs(8156) <= not a;
    layer3_outputs(8157) <= b;
    layer3_outputs(8158) <= b and not a;
    layer3_outputs(8159) <= not b;
    layer3_outputs(8160) <= a;
    layer3_outputs(8161) <= not a or b;
    layer3_outputs(8162) <= a;
    layer3_outputs(8163) <= a;
    layer3_outputs(8164) <= not b or a;
    layer3_outputs(8165) <= a and not b;
    layer3_outputs(8166) <= not b or a;
    layer3_outputs(8167) <= a and b;
    layer3_outputs(8168) <= a;
    layer3_outputs(8169) <= b and not a;
    layer3_outputs(8170) <= a;
    layer3_outputs(8171) <= not a;
    layer3_outputs(8172) <= not b;
    layer3_outputs(8173) <= not (a or b);
    layer3_outputs(8174) <= not (a or b);
    layer3_outputs(8175) <= not b;
    layer3_outputs(8176) <= not (a or b);
    layer3_outputs(8177) <= not a or b;
    layer3_outputs(8178) <= not a or b;
    layer3_outputs(8179) <= not b or a;
    layer3_outputs(8180) <= a and not b;
    layer3_outputs(8181) <= a and not b;
    layer3_outputs(8182) <= '0';
    layer3_outputs(8183) <= a and b;
    layer3_outputs(8184) <= not a or b;
    layer3_outputs(8185) <= a;
    layer3_outputs(8186) <= not b or a;
    layer3_outputs(8187) <= b and not a;
    layer3_outputs(8188) <= not b;
    layer3_outputs(8189) <= not a;
    layer3_outputs(8190) <= a or b;
    layer3_outputs(8191) <= not (a or b);
    layer3_outputs(8192) <= not a or b;
    layer3_outputs(8193) <= not b or a;
    layer3_outputs(8194) <= a and b;
    layer3_outputs(8195) <= a;
    layer3_outputs(8196) <= not (a and b);
    layer3_outputs(8197) <= b;
    layer3_outputs(8198) <= b;
    layer3_outputs(8199) <= not a;
    layer3_outputs(8200) <= a;
    layer3_outputs(8201) <= a and b;
    layer3_outputs(8202) <= not (a and b);
    layer3_outputs(8203) <= a;
    layer3_outputs(8204) <= not b;
    layer3_outputs(8205) <= '0';
    layer3_outputs(8206) <= not a or b;
    layer3_outputs(8207) <= a or b;
    layer3_outputs(8208) <= not (a and b);
    layer3_outputs(8209) <= b;
    layer3_outputs(8210) <= not (a and b);
    layer3_outputs(8211) <= not b;
    layer3_outputs(8212) <= a or b;
    layer3_outputs(8213) <= not (a and b);
    layer3_outputs(8214) <= b and not a;
    layer3_outputs(8215) <= not b;
    layer3_outputs(8216) <= '0';
    layer3_outputs(8217) <= a and not b;
    layer3_outputs(8218) <= a or b;
    layer3_outputs(8219) <= a;
    layer3_outputs(8220) <= b and not a;
    layer3_outputs(8221) <= a and not b;
    layer3_outputs(8222) <= not a;
    layer3_outputs(8223) <= a or b;
    layer3_outputs(8224) <= a and b;
    layer3_outputs(8225) <= not a;
    layer3_outputs(8226) <= b and not a;
    layer3_outputs(8227) <= a or b;
    layer3_outputs(8228) <= a and b;
    layer3_outputs(8229) <= not b;
    layer3_outputs(8230) <= not (a or b);
    layer3_outputs(8231) <= not b;
    layer3_outputs(8232) <= a or b;
    layer3_outputs(8233) <= not (a or b);
    layer3_outputs(8234) <= a xor b;
    layer3_outputs(8235) <= not b or a;
    layer3_outputs(8236) <= a;
    layer3_outputs(8237) <= not b or a;
    layer3_outputs(8238) <= '1';
    layer3_outputs(8239) <= not a;
    layer3_outputs(8240) <= b and not a;
    layer3_outputs(8241) <= b;
    layer3_outputs(8242) <= not a;
    layer3_outputs(8243) <= a;
    layer3_outputs(8244) <= not (a xor b);
    layer3_outputs(8245) <= a and not b;
    layer3_outputs(8246) <= not a;
    layer3_outputs(8247) <= not a;
    layer3_outputs(8248) <= b and not a;
    layer3_outputs(8249) <= not b or a;
    layer3_outputs(8250) <= a and b;
    layer3_outputs(8251) <= a or b;
    layer3_outputs(8252) <= b;
    layer3_outputs(8253) <= '0';
    layer3_outputs(8254) <= a xor b;
    layer3_outputs(8255) <= not a or b;
    layer3_outputs(8256) <= a;
    layer3_outputs(8257) <= not a;
    layer3_outputs(8258) <= a or b;
    layer3_outputs(8259) <= a;
    layer3_outputs(8260) <= a;
    layer3_outputs(8261) <= b and not a;
    layer3_outputs(8262) <= b;
    layer3_outputs(8263) <= a and not b;
    layer3_outputs(8264) <= not b or a;
    layer3_outputs(8265) <= b;
    layer3_outputs(8266) <= b;
    layer3_outputs(8267) <= not (a or b);
    layer3_outputs(8268) <= not b or a;
    layer3_outputs(8269) <= b and not a;
    layer3_outputs(8270) <= not a or b;
    layer3_outputs(8271) <= not a;
    layer3_outputs(8272) <= not (a or b);
    layer3_outputs(8273) <= a or b;
    layer3_outputs(8274) <= not a or b;
    layer3_outputs(8275) <= not b;
    layer3_outputs(8276) <= '1';
    layer3_outputs(8277) <= not a;
    layer3_outputs(8278) <= a;
    layer3_outputs(8279) <= a;
    layer3_outputs(8280) <= a;
    layer3_outputs(8281) <= not (a or b);
    layer3_outputs(8282) <= not (a and b);
    layer3_outputs(8283) <= not (a and b);
    layer3_outputs(8284) <= not b;
    layer3_outputs(8285) <= not a;
    layer3_outputs(8286) <= not (a or b);
    layer3_outputs(8287) <= a and b;
    layer3_outputs(8288) <= a and b;
    layer3_outputs(8289) <= b and not a;
    layer3_outputs(8290) <= not b or a;
    layer3_outputs(8291) <= b and not a;
    layer3_outputs(8292) <= not (a or b);
    layer3_outputs(8293) <= not b or a;
    layer3_outputs(8294) <= a xor b;
    layer3_outputs(8295) <= not b;
    layer3_outputs(8296) <= b;
    layer3_outputs(8297) <= b and not a;
    layer3_outputs(8298) <= a and not b;
    layer3_outputs(8299) <= not a;
    layer3_outputs(8300) <= not (a and b);
    layer3_outputs(8301) <= not a;
    layer3_outputs(8302) <= '0';
    layer3_outputs(8303) <= '1';
    layer3_outputs(8304) <= b;
    layer3_outputs(8305) <= a;
    layer3_outputs(8306) <= '1';
    layer3_outputs(8307) <= a and b;
    layer3_outputs(8308) <= a and b;
    layer3_outputs(8309) <= b;
    layer3_outputs(8310) <= '1';
    layer3_outputs(8311) <= '0';
    layer3_outputs(8312) <= b and not a;
    layer3_outputs(8313) <= b;
    layer3_outputs(8314) <= '1';
    layer3_outputs(8315) <= not b;
    layer3_outputs(8316) <= not a;
    layer3_outputs(8317) <= a and not b;
    layer3_outputs(8318) <= not (a xor b);
    layer3_outputs(8319) <= b and not a;
    layer3_outputs(8320) <= not (a or b);
    layer3_outputs(8321) <= a and not b;
    layer3_outputs(8322) <= b;
    layer3_outputs(8323) <= a and b;
    layer3_outputs(8324) <= not b or a;
    layer3_outputs(8325) <= not a or b;
    layer3_outputs(8326) <= not a or b;
    layer3_outputs(8327) <= a;
    layer3_outputs(8328) <= '1';
    layer3_outputs(8329) <= a or b;
    layer3_outputs(8330) <= not b;
    layer3_outputs(8331) <= b;
    layer3_outputs(8332) <= b;
    layer3_outputs(8333) <= b;
    layer3_outputs(8334) <= a;
    layer3_outputs(8335) <= a or b;
    layer3_outputs(8336) <= not a or b;
    layer3_outputs(8337) <= b;
    layer3_outputs(8338) <= not b;
    layer3_outputs(8339) <= a and not b;
    layer3_outputs(8340) <= a and not b;
    layer3_outputs(8341) <= b and not a;
    layer3_outputs(8342) <= b;
    layer3_outputs(8343) <= not a;
    layer3_outputs(8344) <= a;
    layer3_outputs(8345) <= a;
    layer3_outputs(8346) <= not b;
    layer3_outputs(8347) <= a and b;
    layer3_outputs(8348) <= not b;
    layer3_outputs(8349) <= not b;
    layer3_outputs(8350) <= not b or a;
    layer3_outputs(8351) <= a and not b;
    layer3_outputs(8352) <= not (a or b);
    layer3_outputs(8353) <= b and not a;
    layer3_outputs(8354) <= not b or a;
    layer3_outputs(8355) <= a;
    layer3_outputs(8356) <= not b;
    layer3_outputs(8357) <= '0';
    layer3_outputs(8358) <= not a;
    layer3_outputs(8359) <= '1';
    layer3_outputs(8360) <= not a or b;
    layer3_outputs(8361) <= b;
    layer3_outputs(8362) <= not a;
    layer3_outputs(8363) <= b;
    layer3_outputs(8364) <= not (a or b);
    layer3_outputs(8365) <= not a or b;
    layer3_outputs(8366) <= '1';
    layer3_outputs(8367) <= b;
    layer3_outputs(8368) <= b and not a;
    layer3_outputs(8369) <= not (a or b);
    layer3_outputs(8370) <= not a;
    layer3_outputs(8371) <= not a or b;
    layer3_outputs(8372) <= a or b;
    layer3_outputs(8373) <= b and not a;
    layer3_outputs(8374) <= not b;
    layer3_outputs(8375) <= a or b;
    layer3_outputs(8376) <= a and b;
    layer3_outputs(8377) <= not a;
    layer3_outputs(8378) <= a and b;
    layer3_outputs(8379) <= not b;
    layer3_outputs(8380) <= a xor b;
    layer3_outputs(8381) <= not b;
    layer3_outputs(8382) <= a xor b;
    layer3_outputs(8383) <= not (a xor b);
    layer3_outputs(8384) <= a or b;
    layer3_outputs(8385) <= a and b;
    layer3_outputs(8386) <= not (a xor b);
    layer3_outputs(8387) <= a or b;
    layer3_outputs(8388) <= '0';
    layer3_outputs(8389) <= not a;
    layer3_outputs(8390) <= b;
    layer3_outputs(8391) <= '1';
    layer3_outputs(8392) <= a xor b;
    layer3_outputs(8393) <= b;
    layer3_outputs(8394) <= a and b;
    layer3_outputs(8395) <= '0';
    layer3_outputs(8396) <= a;
    layer3_outputs(8397) <= not (a or b);
    layer3_outputs(8398) <= not b;
    layer3_outputs(8399) <= a;
    layer3_outputs(8400) <= a and not b;
    layer3_outputs(8401) <= '0';
    layer3_outputs(8402) <= not a;
    layer3_outputs(8403) <= not (a or b);
    layer3_outputs(8404) <= a and b;
    layer3_outputs(8405) <= not b;
    layer3_outputs(8406) <= not b;
    layer3_outputs(8407) <= a;
    layer3_outputs(8408) <= a;
    layer3_outputs(8409) <= a or b;
    layer3_outputs(8410) <= not b;
    layer3_outputs(8411) <= b and not a;
    layer3_outputs(8412) <= not (a xor b);
    layer3_outputs(8413) <= not (a xor b);
    layer3_outputs(8414) <= not (a or b);
    layer3_outputs(8415) <= not a or b;
    layer3_outputs(8416) <= not (a and b);
    layer3_outputs(8417) <= not a;
    layer3_outputs(8418) <= a and b;
    layer3_outputs(8419) <= not (a and b);
    layer3_outputs(8420) <= a and b;
    layer3_outputs(8421) <= a xor b;
    layer3_outputs(8422) <= a;
    layer3_outputs(8423) <= '1';
    layer3_outputs(8424) <= a and b;
    layer3_outputs(8425) <= b;
    layer3_outputs(8426) <= a and b;
    layer3_outputs(8427) <= not b;
    layer3_outputs(8428) <= not (a or b);
    layer3_outputs(8429) <= a xor b;
    layer3_outputs(8430) <= not a or b;
    layer3_outputs(8431) <= a and not b;
    layer3_outputs(8432) <= not (a and b);
    layer3_outputs(8433) <= a and not b;
    layer3_outputs(8434) <= a;
    layer3_outputs(8435) <= not a;
    layer3_outputs(8436) <= not (a or b);
    layer3_outputs(8437) <= '1';
    layer3_outputs(8438) <= a and not b;
    layer3_outputs(8439) <= b;
    layer3_outputs(8440) <= not (a and b);
    layer3_outputs(8441) <= not a;
    layer3_outputs(8442) <= not (a and b);
    layer3_outputs(8443) <= b and not a;
    layer3_outputs(8444) <= not a or b;
    layer3_outputs(8445) <= a;
    layer3_outputs(8446) <= not b;
    layer3_outputs(8447) <= a;
    layer3_outputs(8448) <= not b or a;
    layer3_outputs(8449) <= not a;
    layer3_outputs(8450) <= not (a or b);
    layer3_outputs(8451) <= a or b;
    layer3_outputs(8452) <= a;
    layer3_outputs(8453) <= b and not a;
    layer3_outputs(8454) <= a;
    layer3_outputs(8455) <= a and b;
    layer3_outputs(8456) <= not (a or b);
    layer3_outputs(8457) <= b;
    layer3_outputs(8458) <= not b;
    layer3_outputs(8459) <= not b;
    layer3_outputs(8460) <= b;
    layer3_outputs(8461) <= b;
    layer3_outputs(8462) <= b;
    layer3_outputs(8463) <= not (a or b);
    layer3_outputs(8464) <= b;
    layer3_outputs(8465) <= b and not a;
    layer3_outputs(8466) <= b and not a;
    layer3_outputs(8467) <= a and not b;
    layer3_outputs(8468) <= a and b;
    layer3_outputs(8469) <= a or b;
    layer3_outputs(8470) <= not (a and b);
    layer3_outputs(8471) <= a;
    layer3_outputs(8472) <= a or b;
    layer3_outputs(8473) <= not a or b;
    layer3_outputs(8474) <= not b or a;
    layer3_outputs(8475) <= not (a and b);
    layer3_outputs(8476) <= b;
    layer3_outputs(8477) <= a xor b;
    layer3_outputs(8478) <= a xor b;
    layer3_outputs(8479) <= not a;
    layer3_outputs(8480) <= a xor b;
    layer3_outputs(8481) <= a or b;
    layer3_outputs(8482) <= b;
    layer3_outputs(8483) <= not b;
    layer3_outputs(8484) <= a or b;
    layer3_outputs(8485) <= not (a and b);
    layer3_outputs(8486) <= a;
    layer3_outputs(8487) <= not (a xor b);
    layer3_outputs(8488) <= a or b;
    layer3_outputs(8489) <= not (a and b);
    layer3_outputs(8490) <= a xor b;
    layer3_outputs(8491) <= not a;
    layer3_outputs(8492) <= not (a xor b);
    layer3_outputs(8493) <= not b;
    layer3_outputs(8494) <= not (a and b);
    layer3_outputs(8495) <= a and b;
    layer3_outputs(8496) <= a or b;
    layer3_outputs(8497) <= not b;
    layer3_outputs(8498) <= b and not a;
    layer3_outputs(8499) <= not (a or b);
    layer3_outputs(8500) <= b;
    layer3_outputs(8501) <= a or b;
    layer3_outputs(8502) <= not b;
    layer3_outputs(8503) <= not (a and b);
    layer3_outputs(8504) <= b;
    layer3_outputs(8505) <= a;
    layer3_outputs(8506) <= not (a or b);
    layer3_outputs(8507) <= b;
    layer3_outputs(8508) <= a;
    layer3_outputs(8509) <= not (a or b);
    layer3_outputs(8510) <= b and not a;
    layer3_outputs(8511) <= '0';
    layer3_outputs(8512) <= not a or b;
    layer3_outputs(8513) <= a and not b;
    layer3_outputs(8514) <= a xor b;
    layer3_outputs(8515) <= a;
    layer3_outputs(8516) <= not b or a;
    layer3_outputs(8517) <= a;
    layer3_outputs(8518) <= not (a xor b);
    layer3_outputs(8519) <= not (a and b);
    layer3_outputs(8520) <= not a;
    layer3_outputs(8521) <= not (a xor b);
    layer3_outputs(8522) <= b;
    layer3_outputs(8523) <= not b;
    layer3_outputs(8524) <= a or b;
    layer3_outputs(8525) <= '1';
    layer3_outputs(8526) <= not (a xor b);
    layer3_outputs(8527) <= '0';
    layer3_outputs(8528) <= '0';
    layer3_outputs(8529) <= b and not a;
    layer3_outputs(8530) <= a;
    layer3_outputs(8531) <= a and b;
    layer3_outputs(8532) <= '1';
    layer3_outputs(8533) <= a;
    layer3_outputs(8534) <= a;
    layer3_outputs(8535) <= not (a or b);
    layer3_outputs(8536) <= not a or b;
    layer3_outputs(8537) <= not b or a;
    layer3_outputs(8538) <= a;
    layer3_outputs(8539) <= a and not b;
    layer3_outputs(8540) <= a and not b;
    layer3_outputs(8541) <= not b or a;
    layer3_outputs(8542) <= a or b;
    layer3_outputs(8543) <= not b;
    layer3_outputs(8544) <= a or b;
    layer3_outputs(8545) <= a and b;
    layer3_outputs(8546) <= not b;
    layer3_outputs(8547) <= a or b;
    layer3_outputs(8548) <= a;
    layer3_outputs(8549) <= not b;
    layer3_outputs(8550) <= b and not a;
    layer3_outputs(8551) <= not b;
    layer3_outputs(8552) <= a and not b;
    layer3_outputs(8553) <= a and b;
    layer3_outputs(8554) <= not (a and b);
    layer3_outputs(8555) <= a or b;
    layer3_outputs(8556) <= not b or a;
    layer3_outputs(8557) <= b;
    layer3_outputs(8558) <= a and b;
    layer3_outputs(8559) <= not (a or b);
    layer3_outputs(8560) <= b and not a;
    layer3_outputs(8561) <= a and b;
    layer3_outputs(8562) <= not b or a;
    layer3_outputs(8563) <= b and not a;
    layer3_outputs(8564) <= not a;
    layer3_outputs(8565) <= not (a xor b);
    layer3_outputs(8566) <= not (a or b);
    layer3_outputs(8567) <= not (a or b);
    layer3_outputs(8568) <= b;
    layer3_outputs(8569) <= b;
    layer3_outputs(8570) <= not b or a;
    layer3_outputs(8571) <= not (a and b);
    layer3_outputs(8572) <= not a;
    layer3_outputs(8573) <= a and not b;
    layer3_outputs(8574) <= a or b;
    layer3_outputs(8575) <= a and not b;
    layer3_outputs(8576) <= a;
    layer3_outputs(8577) <= a or b;
    layer3_outputs(8578) <= a or b;
    layer3_outputs(8579) <= not b;
    layer3_outputs(8580) <= b;
    layer3_outputs(8581) <= a;
    layer3_outputs(8582) <= '1';
    layer3_outputs(8583) <= b;
    layer3_outputs(8584) <= a xor b;
    layer3_outputs(8585) <= not a;
    layer3_outputs(8586) <= '0';
    layer3_outputs(8587) <= a or b;
    layer3_outputs(8588) <= b;
    layer3_outputs(8589) <= not a;
    layer3_outputs(8590) <= a and not b;
    layer3_outputs(8591) <= a;
    layer3_outputs(8592) <= not a;
    layer3_outputs(8593) <= not b;
    layer3_outputs(8594) <= not b;
    layer3_outputs(8595) <= not (a xor b);
    layer3_outputs(8596) <= not b;
    layer3_outputs(8597) <= not (a or b);
    layer3_outputs(8598) <= a and not b;
    layer3_outputs(8599) <= a;
    layer3_outputs(8600) <= b;
    layer3_outputs(8601) <= not (a xor b);
    layer3_outputs(8602) <= not a;
    layer3_outputs(8603) <= not a;
    layer3_outputs(8604) <= a or b;
    layer3_outputs(8605) <= b;
    layer3_outputs(8606) <= '1';
    layer3_outputs(8607) <= a and b;
    layer3_outputs(8608) <= not (a or b);
    layer3_outputs(8609) <= not b;
    layer3_outputs(8610) <= not (a xor b);
    layer3_outputs(8611) <= a and not b;
    layer3_outputs(8612) <= not (a and b);
    layer3_outputs(8613) <= not a or b;
    layer3_outputs(8614) <= a and not b;
    layer3_outputs(8615) <= '1';
    layer3_outputs(8616) <= a or b;
    layer3_outputs(8617) <= a or b;
    layer3_outputs(8618) <= '1';
    layer3_outputs(8619) <= a or b;
    layer3_outputs(8620) <= not (a and b);
    layer3_outputs(8621) <= b;
    layer3_outputs(8622) <= a;
    layer3_outputs(8623) <= not b;
    layer3_outputs(8624) <= a or b;
    layer3_outputs(8625) <= not a or b;
    layer3_outputs(8626) <= b;
    layer3_outputs(8627) <= not b;
    layer3_outputs(8628) <= not a;
    layer3_outputs(8629) <= not (a and b);
    layer3_outputs(8630) <= b;
    layer3_outputs(8631) <= b;
    layer3_outputs(8632) <= '0';
    layer3_outputs(8633) <= not a;
    layer3_outputs(8634) <= a xor b;
    layer3_outputs(8635) <= b and not a;
    layer3_outputs(8636) <= a;
    layer3_outputs(8637) <= not b or a;
    layer3_outputs(8638) <= not b;
    layer3_outputs(8639) <= a;
    layer3_outputs(8640) <= b and not a;
    layer3_outputs(8641) <= not b;
    layer3_outputs(8642) <= a or b;
    layer3_outputs(8643) <= b;
    layer3_outputs(8644) <= not b or a;
    layer3_outputs(8645) <= not a;
    layer3_outputs(8646) <= a;
    layer3_outputs(8647) <= not b;
    layer3_outputs(8648) <= b and not a;
    layer3_outputs(8649) <= a;
    layer3_outputs(8650) <= a;
    layer3_outputs(8651) <= not b or a;
    layer3_outputs(8652) <= b;
    layer3_outputs(8653) <= a;
    layer3_outputs(8654) <= a xor b;
    layer3_outputs(8655) <= not a or b;
    layer3_outputs(8656) <= b and not a;
    layer3_outputs(8657) <= b;
    layer3_outputs(8658) <= not b or a;
    layer3_outputs(8659) <= '1';
    layer3_outputs(8660) <= not b or a;
    layer3_outputs(8661) <= a xor b;
    layer3_outputs(8662) <= '1';
    layer3_outputs(8663) <= '1';
    layer3_outputs(8664) <= a;
    layer3_outputs(8665) <= not b;
    layer3_outputs(8666) <= a and not b;
    layer3_outputs(8667) <= not (a xor b);
    layer3_outputs(8668) <= not a or b;
    layer3_outputs(8669) <= not a or b;
    layer3_outputs(8670) <= a and b;
    layer3_outputs(8671) <= a xor b;
    layer3_outputs(8672) <= '1';
    layer3_outputs(8673) <= not a;
    layer3_outputs(8674) <= b and not a;
    layer3_outputs(8675) <= not (a and b);
    layer3_outputs(8676) <= a xor b;
    layer3_outputs(8677) <= '1';
    layer3_outputs(8678) <= '1';
    layer3_outputs(8679) <= a or b;
    layer3_outputs(8680) <= a;
    layer3_outputs(8681) <= a or b;
    layer3_outputs(8682) <= a or b;
    layer3_outputs(8683) <= not (a and b);
    layer3_outputs(8684) <= not (a or b);
    layer3_outputs(8685) <= not b;
    layer3_outputs(8686) <= a;
    layer3_outputs(8687) <= b;
    layer3_outputs(8688) <= a or b;
    layer3_outputs(8689) <= b;
    layer3_outputs(8690) <= not b;
    layer3_outputs(8691) <= not a;
    layer3_outputs(8692) <= not a or b;
    layer3_outputs(8693) <= not a or b;
    layer3_outputs(8694) <= not a;
    layer3_outputs(8695) <= b;
    layer3_outputs(8696) <= a or b;
    layer3_outputs(8697) <= a or b;
    layer3_outputs(8698) <= not a;
    layer3_outputs(8699) <= a xor b;
    layer3_outputs(8700) <= '1';
    layer3_outputs(8701) <= a or b;
    layer3_outputs(8702) <= not b;
    layer3_outputs(8703) <= a;
    layer3_outputs(8704) <= '0';
    layer3_outputs(8705) <= b;
    layer3_outputs(8706) <= a and not b;
    layer3_outputs(8707) <= a;
    layer3_outputs(8708) <= '1';
    layer3_outputs(8709) <= b and not a;
    layer3_outputs(8710) <= b;
    layer3_outputs(8711) <= b and not a;
    layer3_outputs(8712) <= b;
    layer3_outputs(8713) <= a or b;
    layer3_outputs(8714) <= b and not a;
    layer3_outputs(8715) <= not a or b;
    layer3_outputs(8716) <= not (a or b);
    layer3_outputs(8717) <= a;
    layer3_outputs(8718) <= a;
    layer3_outputs(8719) <= not a;
    layer3_outputs(8720) <= '0';
    layer3_outputs(8721) <= not a or b;
    layer3_outputs(8722) <= not a or b;
    layer3_outputs(8723) <= not b or a;
    layer3_outputs(8724) <= a and b;
    layer3_outputs(8725) <= a or b;
    layer3_outputs(8726) <= not (a xor b);
    layer3_outputs(8727) <= '0';
    layer3_outputs(8728) <= a or b;
    layer3_outputs(8729) <= '1';
    layer3_outputs(8730) <= b and not a;
    layer3_outputs(8731) <= a and not b;
    layer3_outputs(8732) <= a and b;
    layer3_outputs(8733) <= not b;
    layer3_outputs(8734) <= not (a or b);
    layer3_outputs(8735) <= a and not b;
    layer3_outputs(8736) <= not b;
    layer3_outputs(8737) <= a and not b;
    layer3_outputs(8738) <= a and b;
    layer3_outputs(8739) <= a;
    layer3_outputs(8740) <= not b or a;
    layer3_outputs(8741) <= a;
    layer3_outputs(8742) <= a;
    layer3_outputs(8743) <= not (a or b);
    layer3_outputs(8744) <= not b or a;
    layer3_outputs(8745) <= not b;
    layer3_outputs(8746) <= not a or b;
    layer3_outputs(8747) <= not b;
    layer3_outputs(8748) <= a and not b;
    layer3_outputs(8749) <= a or b;
    layer3_outputs(8750) <= b;
    layer3_outputs(8751) <= a;
    layer3_outputs(8752) <= not (a and b);
    layer3_outputs(8753) <= '0';
    layer3_outputs(8754) <= a xor b;
    layer3_outputs(8755) <= b;
    layer3_outputs(8756) <= not b;
    layer3_outputs(8757) <= a;
    layer3_outputs(8758) <= '0';
    layer3_outputs(8759) <= b;
    layer3_outputs(8760) <= a and b;
    layer3_outputs(8761) <= b and not a;
    layer3_outputs(8762) <= a and b;
    layer3_outputs(8763) <= not a;
    layer3_outputs(8764) <= not a or b;
    layer3_outputs(8765) <= not (a or b);
    layer3_outputs(8766) <= a and not b;
    layer3_outputs(8767) <= '0';
    layer3_outputs(8768) <= a and b;
    layer3_outputs(8769) <= not b;
    layer3_outputs(8770) <= not a or b;
    layer3_outputs(8771) <= a;
    layer3_outputs(8772) <= a and b;
    layer3_outputs(8773) <= a and b;
    layer3_outputs(8774) <= b;
    layer3_outputs(8775) <= not b;
    layer3_outputs(8776) <= not a;
    layer3_outputs(8777) <= not a or b;
    layer3_outputs(8778) <= a and b;
    layer3_outputs(8779) <= b;
    layer3_outputs(8780) <= not b;
    layer3_outputs(8781) <= a or b;
    layer3_outputs(8782) <= not b;
    layer3_outputs(8783) <= not (a or b);
    layer3_outputs(8784) <= b;
    layer3_outputs(8785) <= not (a and b);
    layer3_outputs(8786) <= not b or a;
    layer3_outputs(8787) <= '0';
    layer3_outputs(8788) <= not a or b;
    layer3_outputs(8789) <= b and not a;
    layer3_outputs(8790) <= '1';
    layer3_outputs(8791) <= not (a xor b);
    layer3_outputs(8792) <= not (a or b);
    layer3_outputs(8793) <= '0';
    layer3_outputs(8794) <= not (a or b);
    layer3_outputs(8795) <= not a;
    layer3_outputs(8796) <= a and b;
    layer3_outputs(8797) <= '1';
    layer3_outputs(8798) <= not b;
    layer3_outputs(8799) <= a and b;
    layer3_outputs(8800) <= not (a or b);
    layer3_outputs(8801) <= a and not b;
    layer3_outputs(8802) <= a and not b;
    layer3_outputs(8803) <= not (a and b);
    layer3_outputs(8804) <= a;
    layer3_outputs(8805) <= not (a or b);
    layer3_outputs(8806) <= not (a and b);
    layer3_outputs(8807) <= a or b;
    layer3_outputs(8808) <= not a or b;
    layer3_outputs(8809) <= '0';
    layer3_outputs(8810) <= b and not a;
    layer3_outputs(8811) <= not b;
    layer3_outputs(8812) <= a;
    layer3_outputs(8813) <= not (a and b);
    layer3_outputs(8814) <= a and b;
    layer3_outputs(8815) <= '0';
    layer3_outputs(8816) <= b;
    layer3_outputs(8817) <= a and b;
    layer3_outputs(8818) <= b;
    layer3_outputs(8819) <= not (a xor b);
    layer3_outputs(8820) <= not b;
    layer3_outputs(8821) <= not b or a;
    layer3_outputs(8822) <= a and not b;
    layer3_outputs(8823) <= a;
    layer3_outputs(8824) <= not b or a;
    layer3_outputs(8825) <= b;
    layer3_outputs(8826) <= not (a or b);
    layer3_outputs(8827) <= not (a xor b);
    layer3_outputs(8828) <= '0';
    layer3_outputs(8829) <= not (a xor b);
    layer3_outputs(8830) <= b;
    layer3_outputs(8831) <= not b or a;
    layer3_outputs(8832) <= a and b;
    layer3_outputs(8833) <= not (a and b);
    layer3_outputs(8834) <= a or b;
    layer3_outputs(8835) <= '0';
    layer3_outputs(8836) <= a;
    layer3_outputs(8837) <= not b;
    layer3_outputs(8838) <= a;
    layer3_outputs(8839) <= not a or b;
    layer3_outputs(8840) <= b and not a;
    layer3_outputs(8841) <= not (a or b);
    layer3_outputs(8842) <= '1';
    layer3_outputs(8843) <= a and b;
    layer3_outputs(8844) <= '1';
    layer3_outputs(8845) <= a and b;
    layer3_outputs(8846) <= a;
    layer3_outputs(8847) <= not b;
    layer3_outputs(8848) <= a and b;
    layer3_outputs(8849) <= not a;
    layer3_outputs(8850) <= not b;
    layer3_outputs(8851) <= '1';
    layer3_outputs(8852) <= a or b;
    layer3_outputs(8853) <= not a or b;
    layer3_outputs(8854) <= '1';
    layer3_outputs(8855) <= not b;
    layer3_outputs(8856) <= b and not a;
    layer3_outputs(8857) <= a or b;
    layer3_outputs(8858) <= not a or b;
    layer3_outputs(8859) <= a;
    layer3_outputs(8860) <= not (a and b);
    layer3_outputs(8861) <= not a;
    layer3_outputs(8862) <= a;
    layer3_outputs(8863) <= a;
    layer3_outputs(8864) <= a or b;
    layer3_outputs(8865) <= not (a xor b);
    layer3_outputs(8866) <= not a;
    layer3_outputs(8867) <= a and b;
    layer3_outputs(8868) <= '0';
    layer3_outputs(8869) <= a and not b;
    layer3_outputs(8870) <= not b;
    layer3_outputs(8871) <= b;
    layer3_outputs(8872) <= a and b;
    layer3_outputs(8873) <= a;
    layer3_outputs(8874) <= a xor b;
    layer3_outputs(8875) <= not b or a;
    layer3_outputs(8876) <= b and not a;
    layer3_outputs(8877) <= not a;
    layer3_outputs(8878) <= not b or a;
    layer3_outputs(8879) <= not b;
    layer3_outputs(8880) <= a and not b;
    layer3_outputs(8881) <= not b;
    layer3_outputs(8882) <= a or b;
    layer3_outputs(8883) <= a;
    layer3_outputs(8884) <= not a or b;
    layer3_outputs(8885) <= not a or b;
    layer3_outputs(8886) <= not b;
    layer3_outputs(8887) <= a and b;
    layer3_outputs(8888) <= not (a or b);
    layer3_outputs(8889) <= a and b;
    layer3_outputs(8890) <= not a;
    layer3_outputs(8891) <= b;
    layer3_outputs(8892) <= a and not b;
    layer3_outputs(8893) <= a and b;
    layer3_outputs(8894) <= not b or a;
    layer3_outputs(8895) <= not a;
    layer3_outputs(8896) <= not (a and b);
    layer3_outputs(8897) <= not b or a;
    layer3_outputs(8898) <= '0';
    layer3_outputs(8899) <= not (a xor b);
    layer3_outputs(8900) <= not a or b;
    layer3_outputs(8901) <= not a;
    layer3_outputs(8902) <= a;
    layer3_outputs(8903) <= b;
    layer3_outputs(8904) <= a or b;
    layer3_outputs(8905) <= a and b;
    layer3_outputs(8906) <= a;
    layer3_outputs(8907) <= a and not b;
    layer3_outputs(8908) <= a and b;
    layer3_outputs(8909) <= a and not b;
    layer3_outputs(8910) <= a;
    layer3_outputs(8911) <= b;
    layer3_outputs(8912) <= not a or b;
    layer3_outputs(8913) <= not (a xor b);
    layer3_outputs(8914) <= not a;
    layer3_outputs(8915) <= '1';
    layer3_outputs(8916) <= a;
    layer3_outputs(8917) <= a;
    layer3_outputs(8918) <= not (a or b);
    layer3_outputs(8919) <= b and not a;
    layer3_outputs(8920) <= a and b;
    layer3_outputs(8921) <= a;
    layer3_outputs(8922) <= not a;
    layer3_outputs(8923) <= '0';
    layer3_outputs(8924) <= a and not b;
    layer3_outputs(8925) <= a xor b;
    layer3_outputs(8926) <= not (a and b);
    layer3_outputs(8927) <= a and not b;
    layer3_outputs(8928) <= b;
    layer3_outputs(8929) <= a;
    layer3_outputs(8930) <= a;
    layer3_outputs(8931) <= a;
    layer3_outputs(8932) <= not (a or b);
    layer3_outputs(8933) <= not (a or b);
    layer3_outputs(8934) <= not a;
    layer3_outputs(8935) <= '1';
    layer3_outputs(8936) <= b and not a;
    layer3_outputs(8937) <= b;
    layer3_outputs(8938) <= not b;
    layer3_outputs(8939) <= a and not b;
    layer3_outputs(8940) <= not b;
    layer3_outputs(8941) <= a and not b;
    layer3_outputs(8942) <= not a;
    layer3_outputs(8943) <= not b;
    layer3_outputs(8944) <= b and not a;
    layer3_outputs(8945) <= '0';
    layer3_outputs(8946) <= not (a and b);
    layer3_outputs(8947) <= a xor b;
    layer3_outputs(8948) <= '0';
    layer3_outputs(8949) <= not b or a;
    layer3_outputs(8950) <= '0';
    layer3_outputs(8951) <= not (a and b);
    layer3_outputs(8952) <= a and b;
    layer3_outputs(8953) <= not (a or b);
    layer3_outputs(8954) <= a;
    layer3_outputs(8955) <= b;
    layer3_outputs(8956) <= b and not a;
    layer3_outputs(8957) <= b;
    layer3_outputs(8958) <= not a or b;
    layer3_outputs(8959) <= a or b;
    layer3_outputs(8960) <= not (a or b);
    layer3_outputs(8961) <= not b;
    layer3_outputs(8962) <= a and not b;
    layer3_outputs(8963) <= '0';
    layer3_outputs(8964) <= a xor b;
    layer3_outputs(8965) <= b;
    layer3_outputs(8966) <= not a or b;
    layer3_outputs(8967) <= not a;
    layer3_outputs(8968) <= not b;
    layer3_outputs(8969) <= b;
    layer3_outputs(8970) <= a;
    layer3_outputs(8971) <= a;
    layer3_outputs(8972) <= not b or a;
    layer3_outputs(8973) <= not a;
    layer3_outputs(8974) <= not b;
    layer3_outputs(8975) <= a and b;
    layer3_outputs(8976) <= a;
    layer3_outputs(8977) <= not (a and b);
    layer3_outputs(8978) <= b and not a;
    layer3_outputs(8979) <= not a;
    layer3_outputs(8980) <= not a or b;
    layer3_outputs(8981) <= a and not b;
    layer3_outputs(8982) <= a and b;
    layer3_outputs(8983) <= a or b;
    layer3_outputs(8984) <= not (a xor b);
    layer3_outputs(8985) <= a and not b;
    layer3_outputs(8986) <= b;
    layer3_outputs(8987) <= not b or a;
    layer3_outputs(8988) <= not (a and b);
    layer3_outputs(8989) <= b and not a;
    layer3_outputs(8990) <= '0';
    layer3_outputs(8991) <= b;
    layer3_outputs(8992) <= '0';
    layer3_outputs(8993) <= not a;
    layer3_outputs(8994) <= b;
    layer3_outputs(8995) <= '1';
    layer3_outputs(8996) <= a and b;
    layer3_outputs(8997) <= not a or b;
    layer3_outputs(8998) <= b and not a;
    layer3_outputs(8999) <= not b;
    layer3_outputs(9000) <= b;
    layer3_outputs(9001) <= not (a and b);
    layer3_outputs(9002) <= not b;
    layer3_outputs(9003) <= not (a or b);
    layer3_outputs(9004) <= not a or b;
    layer3_outputs(9005) <= a and b;
    layer3_outputs(9006) <= b;
    layer3_outputs(9007) <= not a or b;
    layer3_outputs(9008) <= not b;
    layer3_outputs(9009) <= b;
    layer3_outputs(9010) <= a;
    layer3_outputs(9011) <= b;
    layer3_outputs(9012) <= not b or a;
    layer3_outputs(9013) <= a;
    layer3_outputs(9014) <= b;
    layer3_outputs(9015) <= '0';
    layer3_outputs(9016) <= not b or a;
    layer3_outputs(9017) <= not a;
    layer3_outputs(9018) <= a or b;
    layer3_outputs(9019) <= a;
    layer3_outputs(9020) <= a;
    layer3_outputs(9021) <= not (a xor b);
    layer3_outputs(9022) <= not b;
    layer3_outputs(9023) <= a;
    layer3_outputs(9024) <= a and not b;
    layer3_outputs(9025) <= a xor b;
    layer3_outputs(9026) <= b;
    layer3_outputs(9027) <= '0';
    layer3_outputs(9028) <= '0';
    layer3_outputs(9029) <= not (a and b);
    layer3_outputs(9030) <= not a or b;
    layer3_outputs(9031) <= a and b;
    layer3_outputs(9032) <= not (a or b);
    layer3_outputs(9033) <= a and b;
    layer3_outputs(9034) <= b and not a;
    layer3_outputs(9035) <= a and not b;
    layer3_outputs(9036) <= not b;
    layer3_outputs(9037) <= not b;
    layer3_outputs(9038) <= a and not b;
    layer3_outputs(9039) <= a;
    layer3_outputs(9040) <= not b;
    layer3_outputs(9041) <= not (a and b);
    layer3_outputs(9042) <= not a;
    layer3_outputs(9043) <= b and not a;
    layer3_outputs(9044) <= not (a and b);
    layer3_outputs(9045) <= a or b;
    layer3_outputs(9046) <= not a;
    layer3_outputs(9047) <= not a;
    layer3_outputs(9048) <= b and not a;
    layer3_outputs(9049) <= a;
    layer3_outputs(9050) <= not b or a;
    layer3_outputs(9051) <= a and b;
    layer3_outputs(9052) <= not a or b;
    layer3_outputs(9053) <= not a or b;
    layer3_outputs(9054) <= not a;
    layer3_outputs(9055) <= not b;
    layer3_outputs(9056) <= a and b;
    layer3_outputs(9057) <= a or b;
    layer3_outputs(9058) <= not (a and b);
    layer3_outputs(9059) <= '0';
    layer3_outputs(9060) <= not (a and b);
    layer3_outputs(9061) <= not a;
    layer3_outputs(9062) <= b;
    layer3_outputs(9063) <= not a or b;
    layer3_outputs(9064) <= a xor b;
    layer3_outputs(9065) <= not a or b;
    layer3_outputs(9066) <= not b;
    layer3_outputs(9067) <= b;
    layer3_outputs(9068) <= not b;
    layer3_outputs(9069) <= a and not b;
    layer3_outputs(9070) <= not b;
    layer3_outputs(9071) <= not (a and b);
    layer3_outputs(9072) <= not a or b;
    layer3_outputs(9073) <= not a or b;
    layer3_outputs(9074) <= not b;
    layer3_outputs(9075) <= b;
    layer3_outputs(9076) <= b and not a;
    layer3_outputs(9077) <= b and not a;
    layer3_outputs(9078) <= not (a and b);
    layer3_outputs(9079) <= a or b;
    layer3_outputs(9080) <= b;
    layer3_outputs(9081) <= not b or a;
    layer3_outputs(9082) <= not b;
    layer3_outputs(9083) <= a;
    layer3_outputs(9084) <= '0';
    layer3_outputs(9085) <= not a or b;
    layer3_outputs(9086) <= not (a xor b);
    layer3_outputs(9087) <= b;
    layer3_outputs(9088) <= not a;
    layer3_outputs(9089) <= a;
    layer3_outputs(9090) <= not (a or b);
    layer3_outputs(9091) <= not b or a;
    layer3_outputs(9092) <= not b;
    layer3_outputs(9093) <= not a or b;
    layer3_outputs(9094) <= not a or b;
    layer3_outputs(9095) <= a and b;
    layer3_outputs(9096) <= a xor b;
    layer3_outputs(9097) <= a or b;
    layer3_outputs(9098) <= not (a xor b);
    layer3_outputs(9099) <= not (a and b);
    layer3_outputs(9100) <= a and b;
    layer3_outputs(9101) <= not b;
    layer3_outputs(9102) <= '1';
    layer3_outputs(9103) <= b;
    layer3_outputs(9104) <= a and b;
    layer3_outputs(9105) <= a or b;
    layer3_outputs(9106) <= b;
    layer3_outputs(9107) <= not (a xor b);
    layer3_outputs(9108) <= '1';
    layer3_outputs(9109) <= b and not a;
    layer3_outputs(9110) <= not b or a;
    layer3_outputs(9111) <= a and not b;
    layer3_outputs(9112) <= b and not a;
    layer3_outputs(9113) <= not b;
    layer3_outputs(9114) <= a;
    layer3_outputs(9115) <= b and not a;
    layer3_outputs(9116) <= not a;
    layer3_outputs(9117) <= a and not b;
    layer3_outputs(9118) <= not b;
    layer3_outputs(9119) <= not b;
    layer3_outputs(9120) <= b and not a;
    layer3_outputs(9121) <= not b;
    layer3_outputs(9122) <= '1';
    layer3_outputs(9123) <= not a;
    layer3_outputs(9124) <= a or b;
    layer3_outputs(9125) <= a and not b;
    layer3_outputs(9126) <= not b or a;
    layer3_outputs(9127) <= a or b;
    layer3_outputs(9128) <= not a;
    layer3_outputs(9129) <= not b;
    layer3_outputs(9130) <= not b;
    layer3_outputs(9131) <= a and b;
    layer3_outputs(9132) <= b and not a;
    layer3_outputs(9133) <= not b;
    layer3_outputs(9134) <= b and not a;
    layer3_outputs(9135) <= '1';
    layer3_outputs(9136) <= b and not a;
    layer3_outputs(9137) <= not b;
    layer3_outputs(9138) <= not b;
    layer3_outputs(9139) <= '0';
    layer3_outputs(9140) <= a;
    layer3_outputs(9141) <= a and not b;
    layer3_outputs(9142) <= a or b;
    layer3_outputs(9143) <= not (a and b);
    layer3_outputs(9144) <= a and b;
    layer3_outputs(9145) <= not (a and b);
    layer3_outputs(9146) <= a and b;
    layer3_outputs(9147) <= not (a or b);
    layer3_outputs(9148) <= '0';
    layer3_outputs(9149) <= '1';
    layer3_outputs(9150) <= '1';
    layer3_outputs(9151) <= b;
    layer3_outputs(9152) <= not (a or b);
    layer3_outputs(9153) <= a and not b;
    layer3_outputs(9154) <= not b;
    layer3_outputs(9155) <= a and not b;
    layer3_outputs(9156) <= not (a xor b);
    layer3_outputs(9157) <= a and not b;
    layer3_outputs(9158) <= b;
    layer3_outputs(9159) <= not b;
    layer3_outputs(9160) <= not (a and b);
    layer3_outputs(9161) <= a and b;
    layer3_outputs(9162) <= b;
    layer3_outputs(9163) <= not (a xor b);
    layer3_outputs(9164) <= b and not a;
    layer3_outputs(9165) <= a and not b;
    layer3_outputs(9166) <= b and not a;
    layer3_outputs(9167) <= not a;
    layer3_outputs(9168) <= a xor b;
    layer3_outputs(9169) <= a;
    layer3_outputs(9170) <= b;
    layer3_outputs(9171) <= not b;
    layer3_outputs(9172) <= not b;
    layer3_outputs(9173) <= a or b;
    layer3_outputs(9174) <= a;
    layer3_outputs(9175) <= not (a and b);
    layer3_outputs(9176) <= not (a xor b);
    layer3_outputs(9177) <= '0';
    layer3_outputs(9178) <= not b;
    layer3_outputs(9179) <= b;
    layer3_outputs(9180) <= a;
    layer3_outputs(9181) <= a and b;
    layer3_outputs(9182) <= b;
    layer3_outputs(9183) <= not a;
    layer3_outputs(9184) <= not (a and b);
    layer3_outputs(9185) <= not b or a;
    layer3_outputs(9186) <= '0';
    layer3_outputs(9187) <= not b;
    layer3_outputs(9188) <= b and not a;
    layer3_outputs(9189) <= b;
    layer3_outputs(9190) <= not a;
    layer3_outputs(9191) <= a and not b;
    layer3_outputs(9192) <= b;
    layer3_outputs(9193) <= b and not a;
    layer3_outputs(9194) <= not a;
    layer3_outputs(9195) <= a and not b;
    layer3_outputs(9196) <= not a;
    layer3_outputs(9197) <= '1';
    layer3_outputs(9198) <= '0';
    layer3_outputs(9199) <= b;
    layer3_outputs(9200) <= '0';
    layer3_outputs(9201) <= b;
    layer3_outputs(9202) <= b;
    layer3_outputs(9203) <= not a;
    layer3_outputs(9204) <= '1';
    layer3_outputs(9205) <= not a;
    layer3_outputs(9206) <= a and b;
    layer3_outputs(9207) <= '0';
    layer3_outputs(9208) <= b and not a;
    layer3_outputs(9209) <= a or b;
    layer3_outputs(9210) <= not (a or b);
    layer3_outputs(9211) <= a or b;
    layer3_outputs(9212) <= not a;
    layer3_outputs(9213) <= not (a or b);
    layer3_outputs(9214) <= b;
    layer3_outputs(9215) <= a xor b;
    layer3_outputs(9216) <= not (a and b);
    layer3_outputs(9217) <= not a or b;
    layer3_outputs(9218) <= not (a and b);
    layer3_outputs(9219) <= not b or a;
    layer3_outputs(9220) <= not (a and b);
    layer3_outputs(9221) <= b and not a;
    layer3_outputs(9222) <= not (a and b);
    layer3_outputs(9223) <= a or b;
    layer3_outputs(9224) <= b and not a;
    layer3_outputs(9225) <= a;
    layer3_outputs(9226) <= not b or a;
    layer3_outputs(9227) <= b and not a;
    layer3_outputs(9228) <= not b;
    layer3_outputs(9229) <= '0';
    layer3_outputs(9230) <= b;
    layer3_outputs(9231) <= a and b;
    layer3_outputs(9232) <= a xor b;
    layer3_outputs(9233) <= a and not b;
    layer3_outputs(9234) <= not a or b;
    layer3_outputs(9235) <= a xor b;
    layer3_outputs(9236) <= a;
    layer3_outputs(9237) <= '1';
    layer3_outputs(9238) <= a;
    layer3_outputs(9239) <= not (a or b);
    layer3_outputs(9240) <= a;
    layer3_outputs(9241) <= '1';
    layer3_outputs(9242) <= not (a and b);
    layer3_outputs(9243) <= not (a and b);
    layer3_outputs(9244) <= not (a or b);
    layer3_outputs(9245) <= a and not b;
    layer3_outputs(9246) <= not b or a;
    layer3_outputs(9247) <= '1';
    layer3_outputs(9248) <= not (a or b);
    layer3_outputs(9249) <= a and b;
    layer3_outputs(9250) <= a or b;
    layer3_outputs(9251) <= not a;
    layer3_outputs(9252) <= not b;
    layer3_outputs(9253) <= '1';
    layer3_outputs(9254) <= a;
    layer3_outputs(9255) <= '0';
    layer3_outputs(9256) <= not a;
    layer3_outputs(9257) <= b and not a;
    layer3_outputs(9258) <= a and not b;
    layer3_outputs(9259) <= not b;
    layer3_outputs(9260) <= '0';
    layer3_outputs(9261) <= a or b;
    layer3_outputs(9262) <= not (a xor b);
    layer3_outputs(9263) <= not (a and b);
    layer3_outputs(9264) <= not (a and b);
    layer3_outputs(9265) <= not (a or b);
    layer3_outputs(9266) <= a and b;
    layer3_outputs(9267) <= a or b;
    layer3_outputs(9268) <= b and not a;
    layer3_outputs(9269) <= not a;
    layer3_outputs(9270) <= a and not b;
    layer3_outputs(9271) <= not (a or b);
    layer3_outputs(9272) <= b;
    layer3_outputs(9273) <= b;
    layer3_outputs(9274) <= a and b;
    layer3_outputs(9275) <= b;
    layer3_outputs(9276) <= not (a and b);
    layer3_outputs(9277) <= not b;
    layer3_outputs(9278) <= not b;
    layer3_outputs(9279) <= not (a or b);
    layer3_outputs(9280) <= a and b;
    layer3_outputs(9281) <= a xor b;
    layer3_outputs(9282) <= b and not a;
    layer3_outputs(9283) <= not (a xor b);
    layer3_outputs(9284) <= b;
    layer3_outputs(9285) <= not b or a;
    layer3_outputs(9286) <= not a or b;
    layer3_outputs(9287) <= not b or a;
    layer3_outputs(9288) <= not (a and b);
    layer3_outputs(9289) <= not a;
    layer3_outputs(9290) <= '0';
    layer3_outputs(9291) <= not b or a;
    layer3_outputs(9292) <= not a;
    layer3_outputs(9293) <= b and not a;
    layer3_outputs(9294) <= b;
    layer3_outputs(9295) <= not b or a;
    layer3_outputs(9296) <= not a;
    layer3_outputs(9297) <= a;
    layer3_outputs(9298) <= b;
    layer3_outputs(9299) <= a or b;
    layer3_outputs(9300) <= not (a or b);
    layer3_outputs(9301) <= not (a or b);
    layer3_outputs(9302) <= not (a or b);
    layer3_outputs(9303) <= not b;
    layer3_outputs(9304) <= not (a and b);
    layer3_outputs(9305) <= not (a or b);
    layer3_outputs(9306) <= not b or a;
    layer3_outputs(9307) <= not (a and b);
    layer3_outputs(9308) <= not a;
    layer3_outputs(9309) <= not (a xor b);
    layer3_outputs(9310) <= not b;
    layer3_outputs(9311) <= '0';
    layer3_outputs(9312) <= a and not b;
    layer3_outputs(9313) <= not b;
    layer3_outputs(9314) <= not a;
    layer3_outputs(9315) <= b;
    layer3_outputs(9316) <= not b;
    layer3_outputs(9317) <= not a;
    layer3_outputs(9318) <= not (a xor b);
    layer3_outputs(9319) <= not b or a;
    layer3_outputs(9320) <= a;
    layer3_outputs(9321) <= b;
    layer3_outputs(9322) <= a and b;
    layer3_outputs(9323) <= a;
    layer3_outputs(9324) <= not a;
    layer3_outputs(9325) <= a and b;
    layer3_outputs(9326) <= b;
    layer3_outputs(9327) <= a;
    layer3_outputs(9328) <= a or b;
    layer3_outputs(9329) <= a;
    layer3_outputs(9330) <= b and not a;
    layer3_outputs(9331) <= not (a xor b);
    layer3_outputs(9332) <= not b;
    layer3_outputs(9333) <= not a;
    layer3_outputs(9334) <= a and b;
    layer3_outputs(9335) <= '1';
    layer3_outputs(9336) <= not b;
    layer3_outputs(9337) <= b;
    layer3_outputs(9338) <= not a or b;
    layer3_outputs(9339) <= not a;
    layer3_outputs(9340) <= not b;
    layer3_outputs(9341) <= not b;
    layer3_outputs(9342) <= not b or a;
    layer3_outputs(9343) <= a and b;
    layer3_outputs(9344) <= not b or a;
    layer3_outputs(9345) <= a or b;
    layer3_outputs(9346) <= not a;
    layer3_outputs(9347) <= '1';
    layer3_outputs(9348) <= b and not a;
    layer3_outputs(9349) <= not (a or b);
    layer3_outputs(9350) <= not b or a;
    layer3_outputs(9351) <= b;
    layer3_outputs(9352) <= not a;
    layer3_outputs(9353) <= a xor b;
    layer3_outputs(9354) <= not b;
    layer3_outputs(9355) <= a and not b;
    layer3_outputs(9356) <= '0';
    layer3_outputs(9357) <= b and not a;
    layer3_outputs(9358) <= not b or a;
    layer3_outputs(9359) <= a and not b;
    layer3_outputs(9360) <= b and not a;
    layer3_outputs(9361) <= not a or b;
    layer3_outputs(9362) <= a;
    layer3_outputs(9363) <= not a;
    layer3_outputs(9364) <= not (a or b);
    layer3_outputs(9365) <= a xor b;
    layer3_outputs(9366) <= '1';
    layer3_outputs(9367) <= not a;
    layer3_outputs(9368) <= b;
    layer3_outputs(9369) <= not (a and b);
    layer3_outputs(9370) <= b;
    layer3_outputs(9371) <= a;
    layer3_outputs(9372) <= not a or b;
    layer3_outputs(9373) <= '0';
    layer3_outputs(9374) <= b;
    layer3_outputs(9375) <= b;
    layer3_outputs(9376) <= not b;
    layer3_outputs(9377) <= a;
    layer3_outputs(9378) <= not b;
    layer3_outputs(9379) <= b and not a;
    layer3_outputs(9380) <= not a or b;
    layer3_outputs(9381) <= not a or b;
    layer3_outputs(9382) <= not (a xor b);
    layer3_outputs(9383) <= a and not b;
    layer3_outputs(9384) <= a;
    layer3_outputs(9385) <= not b;
    layer3_outputs(9386) <= not b or a;
    layer3_outputs(9387) <= a and b;
    layer3_outputs(9388) <= not (a or b);
    layer3_outputs(9389) <= a and b;
    layer3_outputs(9390) <= not (a and b);
    layer3_outputs(9391) <= a;
    layer3_outputs(9392) <= b;
    layer3_outputs(9393) <= not (a or b);
    layer3_outputs(9394) <= not a or b;
    layer3_outputs(9395) <= not a or b;
    layer3_outputs(9396) <= not b or a;
    layer3_outputs(9397) <= a or b;
    layer3_outputs(9398) <= not b or a;
    layer3_outputs(9399) <= not a or b;
    layer3_outputs(9400) <= a;
    layer3_outputs(9401) <= b;
    layer3_outputs(9402) <= a;
    layer3_outputs(9403) <= '1';
    layer3_outputs(9404) <= b;
    layer3_outputs(9405) <= not b;
    layer3_outputs(9406) <= not b or a;
    layer3_outputs(9407) <= not b;
    layer3_outputs(9408) <= not a;
    layer3_outputs(9409) <= b and not a;
    layer3_outputs(9410) <= not a;
    layer3_outputs(9411) <= b;
    layer3_outputs(9412) <= not (a xor b);
    layer3_outputs(9413) <= a or b;
    layer3_outputs(9414) <= not (a and b);
    layer3_outputs(9415) <= not b;
    layer3_outputs(9416) <= b and not a;
    layer3_outputs(9417) <= b;
    layer3_outputs(9418) <= not (a or b);
    layer3_outputs(9419) <= not b;
    layer3_outputs(9420) <= b;
    layer3_outputs(9421) <= a and not b;
    layer3_outputs(9422) <= b;
    layer3_outputs(9423) <= a and not b;
    layer3_outputs(9424) <= a and b;
    layer3_outputs(9425) <= a and not b;
    layer3_outputs(9426) <= b and not a;
    layer3_outputs(9427) <= a and b;
    layer3_outputs(9428) <= a;
    layer3_outputs(9429) <= not a or b;
    layer3_outputs(9430) <= not a;
    layer3_outputs(9431) <= not (a xor b);
    layer3_outputs(9432) <= not a or b;
    layer3_outputs(9433) <= b and not a;
    layer3_outputs(9434) <= '0';
    layer3_outputs(9435) <= not a;
    layer3_outputs(9436) <= a and b;
    layer3_outputs(9437) <= not a or b;
    layer3_outputs(9438) <= a and not b;
    layer3_outputs(9439) <= '0';
    layer3_outputs(9440) <= not a or b;
    layer3_outputs(9441) <= a xor b;
    layer3_outputs(9442) <= not a or b;
    layer3_outputs(9443) <= not b or a;
    layer3_outputs(9444) <= b;
    layer3_outputs(9445) <= not b or a;
    layer3_outputs(9446) <= not b;
    layer3_outputs(9447) <= not a or b;
    layer3_outputs(9448) <= not a;
    layer3_outputs(9449) <= not a;
    layer3_outputs(9450) <= b and not a;
    layer3_outputs(9451) <= b;
    layer3_outputs(9452) <= b;
    layer3_outputs(9453) <= b;
    layer3_outputs(9454) <= a;
    layer3_outputs(9455) <= not b or a;
    layer3_outputs(9456) <= not (a or b);
    layer3_outputs(9457) <= '0';
    layer3_outputs(9458) <= not (a and b);
    layer3_outputs(9459) <= b;
    layer3_outputs(9460) <= not (a and b);
    layer3_outputs(9461) <= not b or a;
    layer3_outputs(9462) <= not b;
    layer3_outputs(9463) <= not b;
    layer3_outputs(9464) <= not a;
    layer3_outputs(9465) <= not a;
    layer3_outputs(9466) <= a xor b;
    layer3_outputs(9467) <= not (a and b);
    layer3_outputs(9468) <= not (a xor b);
    layer3_outputs(9469) <= a and b;
    layer3_outputs(9470) <= not a;
    layer3_outputs(9471) <= not b or a;
    layer3_outputs(9472) <= b;
    layer3_outputs(9473) <= not b or a;
    layer3_outputs(9474) <= a and not b;
    layer3_outputs(9475) <= not a;
    layer3_outputs(9476) <= not (a and b);
    layer3_outputs(9477) <= not b;
    layer3_outputs(9478) <= b and not a;
    layer3_outputs(9479) <= a;
    layer3_outputs(9480) <= not b;
    layer3_outputs(9481) <= not b;
    layer3_outputs(9482) <= not (a xor b);
    layer3_outputs(9483) <= not b;
    layer3_outputs(9484) <= a and b;
    layer3_outputs(9485) <= not a;
    layer3_outputs(9486) <= not (a or b);
    layer3_outputs(9487) <= not (a or b);
    layer3_outputs(9488) <= not b or a;
    layer3_outputs(9489) <= not a;
    layer3_outputs(9490) <= not a or b;
    layer3_outputs(9491) <= b and not a;
    layer3_outputs(9492) <= not a;
    layer3_outputs(9493) <= a xor b;
    layer3_outputs(9494) <= not a or b;
    layer3_outputs(9495) <= a;
    layer3_outputs(9496) <= not a;
    layer3_outputs(9497) <= not a or b;
    layer3_outputs(9498) <= not (a or b);
    layer3_outputs(9499) <= '0';
    layer3_outputs(9500) <= b and not a;
    layer3_outputs(9501) <= a and not b;
    layer3_outputs(9502) <= b;
    layer3_outputs(9503) <= not (a and b);
    layer3_outputs(9504) <= not a or b;
    layer3_outputs(9505) <= a xor b;
    layer3_outputs(9506) <= not a or b;
    layer3_outputs(9507) <= not (a or b);
    layer3_outputs(9508) <= not (a and b);
    layer3_outputs(9509) <= not (a or b);
    layer3_outputs(9510) <= b and not a;
    layer3_outputs(9511) <= not a or b;
    layer3_outputs(9512) <= b and not a;
    layer3_outputs(9513) <= not b;
    layer3_outputs(9514) <= a and b;
    layer3_outputs(9515) <= not b;
    layer3_outputs(9516) <= b;
    layer3_outputs(9517) <= not b;
    layer3_outputs(9518) <= not (a or b);
    layer3_outputs(9519) <= not b;
    layer3_outputs(9520) <= a and not b;
    layer3_outputs(9521) <= '0';
    layer3_outputs(9522) <= not b or a;
    layer3_outputs(9523) <= not b;
    layer3_outputs(9524) <= not b;
    layer3_outputs(9525) <= a;
    layer3_outputs(9526) <= b;
    layer3_outputs(9527) <= a xor b;
    layer3_outputs(9528) <= not b;
    layer3_outputs(9529) <= a;
    layer3_outputs(9530) <= not b or a;
    layer3_outputs(9531) <= a;
    layer3_outputs(9532) <= not a or b;
    layer3_outputs(9533) <= not a;
    layer3_outputs(9534) <= a;
    layer3_outputs(9535) <= not b;
    layer3_outputs(9536) <= a;
    layer3_outputs(9537) <= not b;
    layer3_outputs(9538) <= a or b;
    layer3_outputs(9539) <= a;
    layer3_outputs(9540) <= not b;
    layer3_outputs(9541) <= a xor b;
    layer3_outputs(9542) <= not a;
    layer3_outputs(9543) <= a and not b;
    layer3_outputs(9544) <= b and not a;
    layer3_outputs(9545) <= not (a or b);
    layer3_outputs(9546) <= not b;
    layer3_outputs(9547) <= not (a or b);
    layer3_outputs(9548) <= b;
    layer3_outputs(9549) <= a and not b;
    layer3_outputs(9550) <= not b;
    layer3_outputs(9551) <= not b;
    layer3_outputs(9552) <= a and b;
    layer3_outputs(9553) <= not (a or b);
    layer3_outputs(9554) <= b;
    layer3_outputs(9555) <= a;
    layer3_outputs(9556) <= not (a or b);
    layer3_outputs(9557) <= not (a or b);
    layer3_outputs(9558) <= b;
    layer3_outputs(9559) <= a or b;
    layer3_outputs(9560) <= not a;
    layer3_outputs(9561) <= b;
    layer3_outputs(9562) <= a xor b;
    layer3_outputs(9563) <= not (a or b);
    layer3_outputs(9564) <= a and not b;
    layer3_outputs(9565) <= '0';
    layer3_outputs(9566) <= '1';
    layer3_outputs(9567) <= b and not a;
    layer3_outputs(9568) <= not a;
    layer3_outputs(9569) <= b and not a;
    layer3_outputs(9570) <= not b;
    layer3_outputs(9571) <= a;
    layer3_outputs(9572) <= not a;
    layer3_outputs(9573) <= b;
    layer3_outputs(9574) <= '1';
    layer3_outputs(9575) <= not (a xor b);
    layer3_outputs(9576) <= a;
    layer3_outputs(9577) <= not b;
    layer3_outputs(9578) <= b;
    layer3_outputs(9579) <= not a;
    layer3_outputs(9580) <= not (a and b);
    layer3_outputs(9581) <= a xor b;
    layer3_outputs(9582) <= a and not b;
    layer3_outputs(9583) <= b;
    layer3_outputs(9584) <= '0';
    layer3_outputs(9585) <= b and not a;
    layer3_outputs(9586) <= b and not a;
    layer3_outputs(9587) <= not (a xor b);
    layer3_outputs(9588) <= a;
    layer3_outputs(9589) <= a and not b;
    layer3_outputs(9590) <= not a;
    layer3_outputs(9591) <= a xor b;
    layer3_outputs(9592) <= b;
    layer3_outputs(9593) <= a;
    layer3_outputs(9594) <= a and b;
    layer3_outputs(9595) <= b;
    layer3_outputs(9596) <= not (a xor b);
    layer3_outputs(9597) <= not a;
    layer3_outputs(9598) <= not (a or b);
    layer3_outputs(9599) <= not b;
    layer3_outputs(9600) <= a or b;
    layer3_outputs(9601) <= a or b;
    layer3_outputs(9602) <= not a or b;
    layer3_outputs(9603) <= '1';
    layer3_outputs(9604) <= '0';
    layer3_outputs(9605) <= a;
    layer3_outputs(9606) <= b;
    layer3_outputs(9607) <= a or b;
    layer3_outputs(9608) <= not b or a;
    layer3_outputs(9609) <= b and not a;
    layer3_outputs(9610) <= not (a or b);
    layer3_outputs(9611) <= b;
    layer3_outputs(9612) <= b;
    layer3_outputs(9613) <= not a or b;
    layer3_outputs(9614) <= a and b;
    layer3_outputs(9615) <= a and b;
    layer3_outputs(9616) <= not b;
    layer3_outputs(9617) <= a or b;
    layer3_outputs(9618) <= b;
    layer3_outputs(9619) <= not (a or b);
    layer3_outputs(9620) <= not (a and b);
    layer3_outputs(9621) <= a or b;
    layer3_outputs(9622) <= a xor b;
    layer3_outputs(9623) <= not (a and b);
    layer3_outputs(9624) <= not a;
    layer3_outputs(9625) <= a;
    layer3_outputs(9626) <= b;
    layer3_outputs(9627) <= not (a and b);
    layer3_outputs(9628) <= a or b;
    layer3_outputs(9629) <= a and not b;
    layer3_outputs(9630) <= b;
    layer3_outputs(9631) <= not (a and b);
    layer3_outputs(9632) <= not (a xor b);
    layer3_outputs(9633) <= not b or a;
    layer3_outputs(9634) <= not a;
    layer3_outputs(9635) <= '1';
    layer3_outputs(9636) <= a or b;
    layer3_outputs(9637) <= not b or a;
    layer3_outputs(9638) <= not a;
    layer3_outputs(9639) <= not (a and b);
    layer3_outputs(9640) <= '0';
    layer3_outputs(9641) <= not a or b;
    layer3_outputs(9642) <= not a;
    layer3_outputs(9643) <= not (a and b);
    layer3_outputs(9644) <= not a;
    layer3_outputs(9645) <= not a;
    layer3_outputs(9646) <= not a;
    layer3_outputs(9647) <= a and b;
    layer3_outputs(9648) <= a and not b;
    layer3_outputs(9649) <= not b or a;
    layer3_outputs(9650) <= not (a xor b);
    layer3_outputs(9651) <= not b;
    layer3_outputs(9652) <= not b;
    layer3_outputs(9653) <= not (a xor b);
    layer3_outputs(9654) <= not (a or b);
    layer3_outputs(9655) <= not a or b;
    layer3_outputs(9656) <= a or b;
    layer3_outputs(9657) <= a xor b;
    layer3_outputs(9658) <= b;
    layer3_outputs(9659) <= not a;
    layer3_outputs(9660) <= not (a or b);
    layer3_outputs(9661) <= not b;
    layer3_outputs(9662) <= b;
    layer3_outputs(9663) <= a xor b;
    layer3_outputs(9664) <= a and b;
    layer3_outputs(9665) <= a and not b;
    layer3_outputs(9666) <= b;
    layer3_outputs(9667) <= not (a and b);
    layer3_outputs(9668) <= b;
    layer3_outputs(9669) <= a or b;
    layer3_outputs(9670) <= a;
    layer3_outputs(9671) <= a and b;
    layer3_outputs(9672) <= '1';
    layer3_outputs(9673) <= a or b;
    layer3_outputs(9674) <= not a;
    layer3_outputs(9675) <= b;
    layer3_outputs(9676) <= not b or a;
    layer3_outputs(9677) <= b;
    layer3_outputs(9678) <= not b;
    layer3_outputs(9679) <= not a;
    layer3_outputs(9680) <= '1';
    layer3_outputs(9681) <= a and not b;
    layer3_outputs(9682) <= b and not a;
    layer3_outputs(9683) <= a;
    layer3_outputs(9684) <= a and not b;
    layer3_outputs(9685) <= b and not a;
    layer3_outputs(9686) <= not a;
    layer3_outputs(9687) <= a;
    layer3_outputs(9688) <= a and not b;
    layer3_outputs(9689) <= not a;
    layer3_outputs(9690) <= not b;
    layer3_outputs(9691) <= a;
    layer3_outputs(9692) <= a or b;
    layer3_outputs(9693) <= a and b;
    layer3_outputs(9694) <= not b or a;
    layer3_outputs(9695) <= not (a and b);
    layer3_outputs(9696) <= b and not a;
    layer3_outputs(9697) <= not b;
    layer3_outputs(9698) <= b;
    layer3_outputs(9699) <= a xor b;
    layer3_outputs(9700) <= '1';
    layer3_outputs(9701) <= b and not a;
    layer3_outputs(9702) <= not b;
    layer3_outputs(9703) <= not b or a;
    layer3_outputs(9704) <= not a;
    layer3_outputs(9705) <= a xor b;
    layer3_outputs(9706) <= not a;
    layer3_outputs(9707) <= not (a and b);
    layer3_outputs(9708) <= not (a and b);
    layer3_outputs(9709) <= a and b;
    layer3_outputs(9710) <= b;
    layer3_outputs(9711) <= a or b;
    layer3_outputs(9712) <= not b;
    layer3_outputs(9713) <= a and not b;
    layer3_outputs(9714) <= b and not a;
    layer3_outputs(9715) <= a and b;
    layer3_outputs(9716) <= not b or a;
    layer3_outputs(9717) <= not b or a;
    layer3_outputs(9718) <= a or b;
    layer3_outputs(9719) <= not a;
    layer3_outputs(9720) <= not b;
    layer3_outputs(9721) <= not a;
    layer3_outputs(9722) <= not a or b;
    layer3_outputs(9723) <= b;
    layer3_outputs(9724) <= not b;
    layer3_outputs(9725) <= a and b;
    layer3_outputs(9726) <= not a;
    layer3_outputs(9727) <= a and not b;
    layer3_outputs(9728) <= not (a xor b);
    layer3_outputs(9729) <= a and not b;
    layer3_outputs(9730) <= a;
    layer3_outputs(9731) <= b;
    layer3_outputs(9732) <= a and not b;
    layer3_outputs(9733) <= not b or a;
    layer3_outputs(9734) <= not b or a;
    layer3_outputs(9735) <= not (a and b);
    layer3_outputs(9736) <= b and not a;
    layer3_outputs(9737) <= not b;
    layer3_outputs(9738) <= a and b;
    layer3_outputs(9739) <= a or b;
    layer3_outputs(9740) <= not b;
    layer3_outputs(9741) <= not a or b;
    layer3_outputs(9742) <= '1';
    layer3_outputs(9743) <= not (a xor b);
    layer3_outputs(9744) <= a xor b;
    layer3_outputs(9745) <= b;
    layer3_outputs(9746) <= a and b;
    layer3_outputs(9747) <= b and not a;
    layer3_outputs(9748) <= not a;
    layer3_outputs(9749) <= not (a and b);
    layer3_outputs(9750) <= not (a or b);
    layer3_outputs(9751) <= not b or a;
    layer3_outputs(9752) <= not (a xor b);
    layer3_outputs(9753) <= not b or a;
    layer3_outputs(9754) <= a and not b;
    layer3_outputs(9755) <= a and not b;
    layer3_outputs(9756) <= not b;
    layer3_outputs(9757) <= not b;
    layer3_outputs(9758) <= a and b;
    layer3_outputs(9759) <= not a or b;
    layer3_outputs(9760) <= a and b;
    layer3_outputs(9761) <= not a;
    layer3_outputs(9762) <= not b;
    layer3_outputs(9763) <= '1';
    layer3_outputs(9764) <= not a;
    layer3_outputs(9765) <= '0';
    layer3_outputs(9766) <= a and b;
    layer3_outputs(9767) <= a or b;
    layer3_outputs(9768) <= a and not b;
    layer3_outputs(9769) <= a xor b;
    layer3_outputs(9770) <= a;
    layer3_outputs(9771) <= not b;
    layer3_outputs(9772) <= not b;
    layer3_outputs(9773) <= not b;
    layer3_outputs(9774) <= a;
    layer3_outputs(9775) <= a or b;
    layer3_outputs(9776) <= not a;
    layer3_outputs(9777) <= not (a or b);
    layer3_outputs(9778) <= a;
    layer3_outputs(9779) <= a;
    layer3_outputs(9780) <= '0';
    layer3_outputs(9781) <= not b or a;
    layer3_outputs(9782) <= b and not a;
    layer3_outputs(9783) <= a or b;
    layer3_outputs(9784) <= '1';
    layer3_outputs(9785) <= a and b;
    layer3_outputs(9786) <= not a or b;
    layer3_outputs(9787) <= b and not a;
    layer3_outputs(9788) <= a or b;
    layer3_outputs(9789) <= a or b;
    layer3_outputs(9790) <= b;
    layer3_outputs(9791) <= a;
    layer3_outputs(9792) <= not (a or b);
    layer3_outputs(9793) <= not b or a;
    layer3_outputs(9794) <= a;
    layer3_outputs(9795) <= not a;
    layer3_outputs(9796) <= b and not a;
    layer3_outputs(9797) <= a xor b;
    layer3_outputs(9798) <= not a or b;
    layer3_outputs(9799) <= a or b;
    layer3_outputs(9800) <= b;
    layer3_outputs(9801) <= not (a xor b);
    layer3_outputs(9802) <= a;
    layer3_outputs(9803) <= a;
    layer3_outputs(9804) <= a and b;
    layer3_outputs(9805) <= not a;
    layer3_outputs(9806) <= not (a or b);
    layer3_outputs(9807) <= not (a xor b);
    layer3_outputs(9808) <= not (a xor b);
    layer3_outputs(9809) <= not b or a;
    layer3_outputs(9810) <= not a;
    layer3_outputs(9811) <= '0';
    layer3_outputs(9812) <= a and b;
    layer3_outputs(9813) <= not (a and b);
    layer3_outputs(9814) <= not a;
    layer3_outputs(9815) <= not b or a;
    layer3_outputs(9816) <= not a;
    layer3_outputs(9817) <= a or b;
    layer3_outputs(9818) <= not (a xor b);
    layer3_outputs(9819) <= a or b;
    layer3_outputs(9820) <= b;
    layer3_outputs(9821) <= '0';
    layer3_outputs(9822) <= not b;
    layer3_outputs(9823) <= not (a or b);
    layer3_outputs(9824) <= a and not b;
    layer3_outputs(9825) <= not a or b;
    layer3_outputs(9826) <= not b or a;
    layer3_outputs(9827) <= not (a xor b);
    layer3_outputs(9828) <= not b;
    layer3_outputs(9829) <= a and b;
    layer3_outputs(9830) <= a xor b;
    layer3_outputs(9831) <= not (a or b);
    layer3_outputs(9832) <= not b or a;
    layer3_outputs(9833) <= not a or b;
    layer3_outputs(9834) <= '0';
    layer3_outputs(9835) <= a and b;
    layer3_outputs(9836) <= not b;
    layer3_outputs(9837) <= not (a xor b);
    layer3_outputs(9838) <= a xor b;
    layer3_outputs(9839) <= a and not b;
    layer3_outputs(9840) <= '0';
    layer3_outputs(9841) <= '1';
    layer3_outputs(9842) <= not a;
    layer3_outputs(9843) <= not (a or b);
    layer3_outputs(9844) <= not (a or b);
    layer3_outputs(9845) <= a and not b;
    layer3_outputs(9846) <= '0';
    layer3_outputs(9847) <= not (a and b);
    layer3_outputs(9848) <= not b;
    layer3_outputs(9849) <= a and b;
    layer3_outputs(9850) <= b;
    layer3_outputs(9851) <= a and b;
    layer3_outputs(9852) <= a and not b;
    layer3_outputs(9853) <= not (a or b);
    layer3_outputs(9854) <= a and b;
    layer3_outputs(9855) <= b and not a;
    layer3_outputs(9856) <= not (a or b);
    layer3_outputs(9857) <= not (a xor b);
    layer3_outputs(9858) <= not b or a;
    layer3_outputs(9859) <= '0';
    layer3_outputs(9860) <= b;
    layer3_outputs(9861) <= b and not a;
    layer3_outputs(9862) <= not (a or b);
    layer3_outputs(9863) <= b;
    layer3_outputs(9864) <= not a;
    layer3_outputs(9865) <= not a;
    layer3_outputs(9866) <= not b;
    layer3_outputs(9867) <= a and not b;
    layer3_outputs(9868) <= a xor b;
    layer3_outputs(9869) <= not a;
    layer3_outputs(9870) <= a and b;
    layer3_outputs(9871) <= a or b;
    layer3_outputs(9872) <= a and not b;
    layer3_outputs(9873) <= not a;
    layer3_outputs(9874) <= not a;
    layer3_outputs(9875) <= a;
    layer3_outputs(9876) <= not b or a;
    layer3_outputs(9877) <= '0';
    layer3_outputs(9878) <= not b;
    layer3_outputs(9879) <= a or b;
    layer3_outputs(9880) <= not b;
    layer3_outputs(9881) <= not (a xor b);
    layer3_outputs(9882) <= not a or b;
    layer3_outputs(9883) <= not b;
    layer3_outputs(9884) <= not (a or b);
    layer3_outputs(9885) <= b and not a;
    layer3_outputs(9886) <= a and not b;
    layer3_outputs(9887) <= a xor b;
    layer3_outputs(9888) <= '1';
    layer3_outputs(9889) <= not a;
    layer3_outputs(9890) <= b and not a;
    layer3_outputs(9891) <= a or b;
    layer3_outputs(9892) <= '0';
    layer3_outputs(9893) <= a and not b;
    layer3_outputs(9894) <= b and not a;
    layer3_outputs(9895) <= not b;
    layer3_outputs(9896) <= not a;
    layer3_outputs(9897) <= not (a or b);
    layer3_outputs(9898) <= not b or a;
    layer3_outputs(9899) <= a or b;
    layer3_outputs(9900) <= a xor b;
    layer3_outputs(9901) <= not (a or b);
    layer3_outputs(9902) <= a and b;
    layer3_outputs(9903) <= a and b;
    layer3_outputs(9904) <= not b;
    layer3_outputs(9905) <= not a;
    layer3_outputs(9906) <= b and not a;
    layer3_outputs(9907) <= a and b;
    layer3_outputs(9908) <= not b;
    layer3_outputs(9909) <= a;
    layer3_outputs(9910) <= b;
    layer3_outputs(9911) <= not (a xor b);
    layer3_outputs(9912) <= b and not a;
    layer3_outputs(9913) <= b;
    layer3_outputs(9914) <= not b;
    layer3_outputs(9915) <= a and not b;
    layer3_outputs(9916) <= '1';
    layer3_outputs(9917) <= not a or b;
    layer3_outputs(9918) <= not a;
    layer3_outputs(9919) <= not b;
    layer3_outputs(9920) <= not b;
    layer3_outputs(9921) <= not a;
    layer3_outputs(9922) <= not a or b;
    layer3_outputs(9923) <= a and b;
    layer3_outputs(9924) <= a;
    layer3_outputs(9925) <= not (a and b);
    layer3_outputs(9926) <= not b or a;
    layer3_outputs(9927) <= b;
    layer3_outputs(9928) <= not a or b;
    layer3_outputs(9929) <= a and not b;
    layer3_outputs(9930) <= '1';
    layer3_outputs(9931) <= not (a and b);
    layer3_outputs(9932) <= a and not b;
    layer3_outputs(9933) <= b;
    layer3_outputs(9934) <= a xor b;
    layer3_outputs(9935) <= not a or b;
    layer3_outputs(9936) <= '0';
    layer3_outputs(9937) <= not (a xor b);
    layer3_outputs(9938) <= not a or b;
    layer3_outputs(9939) <= not b or a;
    layer3_outputs(9940) <= a and b;
    layer3_outputs(9941) <= '1';
    layer3_outputs(9942) <= not b;
    layer3_outputs(9943) <= not b or a;
    layer3_outputs(9944) <= '0';
    layer3_outputs(9945) <= not (a xor b);
    layer3_outputs(9946) <= a and not b;
    layer3_outputs(9947) <= not b or a;
    layer3_outputs(9948) <= a or b;
    layer3_outputs(9949) <= not b;
    layer3_outputs(9950) <= not a;
    layer3_outputs(9951) <= '1';
    layer3_outputs(9952) <= '0';
    layer3_outputs(9953) <= b and not a;
    layer3_outputs(9954) <= not a or b;
    layer3_outputs(9955) <= '0';
    layer3_outputs(9956) <= '1';
    layer3_outputs(9957) <= not a;
    layer3_outputs(9958) <= not (a or b);
    layer3_outputs(9959) <= b;
    layer3_outputs(9960) <= '0';
    layer3_outputs(9961) <= not b;
    layer3_outputs(9962) <= not (a and b);
    layer3_outputs(9963) <= not a or b;
    layer3_outputs(9964) <= not a or b;
    layer3_outputs(9965) <= b;
    layer3_outputs(9966) <= '0';
    layer3_outputs(9967) <= b;
    layer3_outputs(9968) <= a;
    layer3_outputs(9969) <= not b;
    layer3_outputs(9970) <= not (a or b);
    layer3_outputs(9971) <= not a or b;
    layer3_outputs(9972) <= b;
    layer3_outputs(9973) <= not a;
    layer3_outputs(9974) <= a;
    layer3_outputs(9975) <= a;
    layer3_outputs(9976) <= '0';
    layer3_outputs(9977) <= not (a and b);
    layer3_outputs(9978) <= not (a and b);
    layer3_outputs(9979) <= a;
    layer3_outputs(9980) <= a;
    layer3_outputs(9981) <= not b;
    layer3_outputs(9982) <= a;
    layer3_outputs(9983) <= not b or a;
    layer3_outputs(9984) <= not b or a;
    layer3_outputs(9985) <= b and not a;
    layer3_outputs(9986) <= a xor b;
    layer3_outputs(9987) <= b;
    layer3_outputs(9988) <= not b;
    layer3_outputs(9989) <= b and not a;
    layer3_outputs(9990) <= a and b;
    layer3_outputs(9991) <= a xor b;
    layer3_outputs(9992) <= a xor b;
    layer3_outputs(9993) <= b;
    layer3_outputs(9994) <= '1';
    layer3_outputs(9995) <= not b;
    layer3_outputs(9996) <= not b or a;
    layer3_outputs(9997) <= '1';
    layer3_outputs(9998) <= not a or b;
    layer3_outputs(9999) <= '1';
    layer3_outputs(10000) <= not (a and b);
    layer3_outputs(10001) <= not a or b;
    layer3_outputs(10002) <= b and not a;
    layer3_outputs(10003) <= a xor b;
    layer3_outputs(10004) <= not b;
    layer3_outputs(10005) <= not (a xor b);
    layer3_outputs(10006) <= not a;
    layer3_outputs(10007) <= not b;
    layer3_outputs(10008) <= not (a and b);
    layer3_outputs(10009) <= a and b;
    layer3_outputs(10010) <= a xor b;
    layer3_outputs(10011) <= a;
    layer3_outputs(10012) <= a;
    layer3_outputs(10013) <= not b or a;
    layer3_outputs(10014) <= '1';
    layer3_outputs(10015) <= a;
    layer3_outputs(10016) <= a or b;
    layer3_outputs(10017) <= not a;
    layer3_outputs(10018) <= not b;
    layer3_outputs(10019) <= not (a xor b);
    layer3_outputs(10020) <= a and b;
    layer3_outputs(10021) <= not b;
    layer3_outputs(10022) <= b;
    layer3_outputs(10023) <= a and b;
    layer3_outputs(10024) <= a;
    layer3_outputs(10025) <= not a or b;
    layer3_outputs(10026) <= a and b;
    layer3_outputs(10027) <= not a;
    layer3_outputs(10028) <= a;
    layer3_outputs(10029) <= not a;
    layer3_outputs(10030) <= not a;
    layer3_outputs(10031) <= a and not b;
    layer3_outputs(10032) <= a or b;
    layer3_outputs(10033) <= a;
    layer3_outputs(10034) <= a;
    layer3_outputs(10035) <= a and not b;
    layer3_outputs(10036) <= not b;
    layer3_outputs(10037) <= not b;
    layer3_outputs(10038) <= '1';
    layer3_outputs(10039) <= a or b;
    layer3_outputs(10040) <= '1';
    layer3_outputs(10041) <= a xor b;
    layer3_outputs(10042) <= '0';
    layer3_outputs(10043) <= a;
    layer3_outputs(10044) <= '0';
    layer3_outputs(10045) <= not (a or b);
    layer3_outputs(10046) <= '1';
    layer3_outputs(10047) <= a;
    layer3_outputs(10048) <= a xor b;
    layer3_outputs(10049) <= b and not a;
    layer3_outputs(10050) <= not b;
    layer3_outputs(10051) <= not b or a;
    layer3_outputs(10052) <= not a;
    layer3_outputs(10053) <= not a;
    layer3_outputs(10054) <= '0';
    layer3_outputs(10055) <= not (a and b);
    layer3_outputs(10056) <= a and b;
    layer3_outputs(10057) <= a;
    layer3_outputs(10058) <= a;
    layer3_outputs(10059) <= not (a or b);
    layer3_outputs(10060) <= b;
    layer3_outputs(10061) <= a and not b;
    layer3_outputs(10062) <= not (a xor b);
    layer3_outputs(10063) <= b;
    layer3_outputs(10064) <= not (a xor b);
    layer3_outputs(10065) <= not (a or b);
    layer3_outputs(10066) <= a and b;
    layer3_outputs(10067) <= '1';
    layer3_outputs(10068) <= not (a xor b);
    layer3_outputs(10069) <= a or b;
    layer3_outputs(10070) <= b and not a;
    layer3_outputs(10071) <= a;
    layer3_outputs(10072) <= b;
    layer3_outputs(10073) <= a and not b;
    layer3_outputs(10074) <= a;
    layer3_outputs(10075) <= not b;
    layer3_outputs(10076) <= a;
    layer3_outputs(10077) <= not (a or b);
    layer3_outputs(10078) <= a;
    layer3_outputs(10079) <= a xor b;
    layer3_outputs(10080) <= a or b;
    layer3_outputs(10081) <= not (a or b);
    layer3_outputs(10082) <= not (a and b);
    layer3_outputs(10083) <= a and b;
    layer3_outputs(10084) <= b and not a;
    layer3_outputs(10085) <= a xor b;
    layer3_outputs(10086) <= not a;
    layer3_outputs(10087) <= b;
    layer3_outputs(10088) <= not a or b;
    layer3_outputs(10089) <= a and b;
    layer3_outputs(10090) <= a or b;
    layer3_outputs(10091) <= not a;
    layer3_outputs(10092) <= a xor b;
    layer3_outputs(10093) <= not b;
    layer3_outputs(10094) <= a;
    layer3_outputs(10095) <= a;
    layer3_outputs(10096) <= not a or b;
    layer3_outputs(10097) <= '0';
    layer3_outputs(10098) <= a and b;
    layer3_outputs(10099) <= a and not b;
    layer3_outputs(10100) <= a;
    layer3_outputs(10101) <= a;
    layer3_outputs(10102) <= '1';
    layer3_outputs(10103) <= a or b;
    layer3_outputs(10104) <= not a;
    layer3_outputs(10105) <= not (a or b);
    layer3_outputs(10106) <= b;
    layer3_outputs(10107) <= not b;
    layer3_outputs(10108) <= a;
    layer3_outputs(10109) <= '0';
    layer3_outputs(10110) <= not (a or b);
    layer3_outputs(10111) <= not a;
    layer3_outputs(10112) <= not (a and b);
    layer3_outputs(10113) <= not (a or b);
    layer3_outputs(10114) <= not b;
    layer3_outputs(10115) <= a and b;
    layer3_outputs(10116) <= b;
    layer3_outputs(10117) <= not a;
    layer3_outputs(10118) <= not a;
    layer3_outputs(10119) <= b;
    layer3_outputs(10120) <= b;
    layer3_outputs(10121) <= not (a and b);
    layer3_outputs(10122) <= not (a and b);
    layer3_outputs(10123) <= not b or a;
    layer3_outputs(10124) <= a or b;
    layer3_outputs(10125) <= a;
    layer3_outputs(10126) <= not b;
    layer3_outputs(10127) <= not (a or b);
    layer3_outputs(10128) <= b;
    layer3_outputs(10129) <= a and b;
    layer3_outputs(10130) <= '0';
    layer3_outputs(10131) <= not b;
    layer3_outputs(10132) <= a;
    layer3_outputs(10133) <= b;
    layer3_outputs(10134) <= not a or b;
    layer3_outputs(10135) <= a;
    layer3_outputs(10136) <= not (a or b);
    layer3_outputs(10137) <= a and b;
    layer3_outputs(10138) <= b and not a;
    layer3_outputs(10139) <= a;
    layer3_outputs(10140) <= a xor b;
    layer3_outputs(10141) <= a and b;
    layer3_outputs(10142) <= a xor b;
    layer3_outputs(10143) <= not (a or b);
    layer3_outputs(10144) <= not b;
    layer3_outputs(10145) <= not b;
    layer3_outputs(10146) <= '0';
    layer3_outputs(10147) <= not (a xor b);
    layer3_outputs(10148) <= a and not b;
    layer3_outputs(10149) <= a;
    layer3_outputs(10150) <= a;
    layer3_outputs(10151) <= not b;
    layer3_outputs(10152) <= a;
    layer3_outputs(10153) <= '1';
    layer3_outputs(10154) <= not b or a;
    layer3_outputs(10155) <= b;
    layer3_outputs(10156) <= not a;
    layer3_outputs(10157) <= a and not b;
    layer3_outputs(10158) <= not a or b;
    layer3_outputs(10159) <= not b;
    layer3_outputs(10160) <= not (a and b);
    layer3_outputs(10161) <= not b or a;
    layer3_outputs(10162) <= b;
    layer3_outputs(10163) <= a xor b;
    layer3_outputs(10164) <= a;
    layer3_outputs(10165) <= not (a xor b);
    layer3_outputs(10166) <= b and not a;
    layer3_outputs(10167) <= not (a or b);
    layer3_outputs(10168) <= a and b;
    layer3_outputs(10169) <= a;
    layer3_outputs(10170) <= not (a and b);
    layer3_outputs(10171) <= '1';
    layer3_outputs(10172) <= not a;
    layer3_outputs(10173) <= b;
    layer3_outputs(10174) <= not a;
    layer3_outputs(10175) <= b;
    layer3_outputs(10176) <= a and b;
    layer3_outputs(10177) <= b and not a;
    layer3_outputs(10178) <= a;
    layer3_outputs(10179) <= not (a or b);
    layer3_outputs(10180) <= a xor b;
    layer3_outputs(10181) <= not b;
    layer3_outputs(10182) <= a and b;
    layer3_outputs(10183) <= b and not a;
    layer3_outputs(10184) <= not (a or b);
    layer3_outputs(10185) <= b;
    layer3_outputs(10186) <= not a;
    layer3_outputs(10187) <= not a;
    layer3_outputs(10188) <= not b;
    layer3_outputs(10189) <= not b;
    layer3_outputs(10190) <= a;
    layer3_outputs(10191) <= '1';
    layer3_outputs(10192) <= not (a or b);
    layer3_outputs(10193) <= a;
    layer3_outputs(10194) <= '1';
    layer3_outputs(10195) <= not a;
    layer3_outputs(10196) <= a;
    layer3_outputs(10197) <= b and not a;
    layer3_outputs(10198) <= not b;
    layer3_outputs(10199) <= a;
    layer3_outputs(10200) <= not a;
    layer3_outputs(10201) <= not (a xor b);
    layer3_outputs(10202) <= a and not b;
    layer3_outputs(10203) <= b;
    layer3_outputs(10204) <= a;
    layer3_outputs(10205) <= not (a or b);
    layer3_outputs(10206) <= not (a xor b);
    layer3_outputs(10207) <= a and b;
    layer3_outputs(10208) <= a and not b;
    layer3_outputs(10209) <= b;
    layer3_outputs(10210) <= a;
    layer3_outputs(10211) <= not b;
    layer3_outputs(10212) <= a and not b;
    layer3_outputs(10213) <= a and b;
    layer3_outputs(10214) <= a and not b;
    layer3_outputs(10215) <= not a or b;
    layer3_outputs(10216) <= not a or b;
    layer3_outputs(10217) <= not a;
    layer3_outputs(10218) <= b and not a;
    layer3_outputs(10219) <= not a;
    layer3_outputs(10220) <= not (a and b);
    layer3_outputs(10221) <= not a;
    layer3_outputs(10222) <= not b;
    layer3_outputs(10223) <= a and b;
    layer3_outputs(10224) <= not b;
    layer3_outputs(10225) <= a and b;
    layer3_outputs(10226) <= not (a and b);
    layer3_outputs(10227) <= '1';
    layer3_outputs(10228) <= a or b;
    layer3_outputs(10229) <= '0';
    layer3_outputs(10230) <= not b;
    layer3_outputs(10231) <= not a;
    layer3_outputs(10232) <= b and not a;
    layer3_outputs(10233) <= not (a or b);
    layer3_outputs(10234) <= b and not a;
    layer3_outputs(10235) <= not a;
    layer3_outputs(10236) <= '0';
    layer3_outputs(10237) <= '0';
    layer3_outputs(10238) <= a xor b;
    layer3_outputs(10239) <= a;
    layer3_outputs(10240) <= not (a and b);
    layer3_outputs(10241) <= not (a and b);
    layer3_outputs(10242) <= a and not b;
    layer3_outputs(10243) <= b;
    layer3_outputs(10244) <= a and not b;
    layer3_outputs(10245) <= a and b;
    layer3_outputs(10246) <= not (a and b);
    layer3_outputs(10247) <= a or b;
    layer3_outputs(10248) <= not (a xor b);
    layer3_outputs(10249) <= a;
    layer3_outputs(10250) <= not a or b;
    layer3_outputs(10251) <= a and b;
    layer3_outputs(10252) <= not a or b;
    layer3_outputs(10253) <= not b;
    layer3_outputs(10254) <= not b or a;
    layer3_outputs(10255) <= a;
    layer3_outputs(10256) <= not a;
    layer3_outputs(10257) <= not a;
    layer3_outputs(10258) <= not a or b;
    layer3_outputs(10259) <= not (a or b);
    layer3_outputs(10260) <= a or b;
    layer3_outputs(10261) <= a and b;
    layer3_outputs(10262) <= b;
    layer3_outputs(10263) <= not b or a;
    layer3_outputs(10264) <= not a or b;
    layer3_outputs(10265) <= not (a xor b);
    layer3_outputs(10266) <= not (a xor b);
    layer3_outputs(10267) <= b and not a;
    layer3_outputs(10268) <= not b;
    layer3_outputs(10269) <= not a or b;
    layer3_outputs(10270) <= b;
    layer3_outputs(10271) <= not a;
    layer3_outputs(10272) <= not a or b;
    layer3_outputs(10273) <= not b;
    layer3_outputs(10274) <= a xor b;
    layer3_outputs(10275) <= a or b;
    layer3_outputs(10276) <= not b;
    layer3_outputs(10277) <= not b;
    layer3_outputs(10278) <= not b or a;
    layer3_outputs(10279) <= a and not b;
    layer3_outputs(10280) <= not a;
    layer3_outputs(10281) <= not (a xor b);
    layer3_outputs(10282) <= b;
    layer3_outputs(10283) <= not a;
    layer3_outputs(10284) <= b;
    layer3_outputs(10285) <= a;
    layer3_outputs(10286) <= not b;
    layer3_outputs(10287) <= a and b;
    layer3_outputs(10288) <= not (a or b);
    layer3_outputs(10289) <= '1';
    layer3_outputs(10290) <= not a;
    layer3_outputs(10291) <= not (a or b);
    layer3_outputs(10292) <= not (a and b);
    layer3_outputs(10293) <= not b;
    layer3_outputs(10294) <= not (a or b);
    layer3_outputs(10295) <= not a or b;
    layer3_outputs(10296) <= not (a and b);
    layer3_outputs(10297) <= not a;
    layer3_outputs(10298) <= not (a or b);
    layer3_outputs(10299) <= a or b;
    layer3_outputs(10300) <= a xor b;
    layer3_outputs(10301) <= '0';
    layer3_outputs(10302) <= not a;
    layer3_outputs(10303) <= a or b;
    layer3_outputs(10304) <= a and not b;
    layer3_outputs(10305) <= a;
    layer3_outputs(10306) <= a and not b;
    layer3_outputs(10307) <= not (a or b);
    layer3_outputs(10308) <= a or b;
    layer3_outputs(10309) <= a;
    layer3_outputs(10310) <= a or b;
    layer3_outputs(10311) <= a;
    layer3_outputs(10312) <= a or b;
    layer3_outputs(10313) <= not (a and b);
    layer3_outputs(10314) <= a and b;
    layer3_outputs(10315) <= not (a or b);
    layer3_outputs(10316) <= a;
    layer3_outputs(10317) <= a and not b;
    layer3_outputs(10318) <= not b;
    layer3_outputs(10319) <= not a or b;
    layer3_outputs(10320) <= not a;
    layer3_outputs(10321) <= b;
    layer3_outputs(10322) <= not (a and b);
    layer3_outputs(10323) <= not b or a;
    layer3_outputs(10324) <= b;
    layer3_outputs(10325) <= '1';
    layer3_outputs(10326) <= a xor b;
    layer3_outputs(10327) <= not a or b;
    layer3_outputs(10328) <= a and b;
    layer3_outputs(10329) <= b and not a;
    layer3_outputs(10330) <= b and not a;
    layer3_outputs(10331) <= a;
    layer3_outputs(10332) <= not b;
    layer3_outputs(10333) <= a and not b;
    layer3_outputs(10334) <= not (a xor b);
    layer3_outputs(10335) <= b;
    layer3_outputs(10336) <= not a;
    layer3_outputs(10337) <= a;
    layer3_outputs(10338) <= b;
    layer3_outputs(10339) <= not b or a;
    layer3_outputs(10340) <= b;
    layer3_outputs(10341) <= a;
    layer3_outputs(10342) <= not a or b;
    layer3_outputs(10343) <= a;
    layer3_outputs(10344) <= a or b;
    layer3_outputs(10345) <= '0';
    layer3_outputs(10346) <= a xor b;
    layer3_outputs(10347) <= not b or a;
    layer3_outputs(10348) <= a and b;
    layer3_outputs(10349) <= not a;
    layer3_outputs(10350) <= not a;
    layer3_outputs(10351) <= not (a or b);
    layer3_outputs(10352) <= not a;
    layer3_outputs(10353) <= b and not a;
    layer3_outputs(10354) <= not (a and b);
    layer3_outputs(10355) <= not a;
    layer3_outputs(10356) <= not a;
    layer3_outputs(10357) <= a and b;
    layer3_outputs(10358) <= b;
    layer3_outputs(10359) <= not (a and b);
    layer3_outputs(10360) <= not a or b;
    layer3_outputs(10361) <= a xor b;
    layer3_outputs(10362) <= not b or a;
    layer3_outputs(10363) <= b;
    layer3_outputs(10364) <= a xor b;
    layer3_outputs(10365) <= '0';
    layer3_outputs(10366) <= a or b;
    layer3_outputs(10367) <= '1';
    layer3_outputs(10368) <= a or b;
    layer3_outputs(10369) <= not b;
    layer3_outputs(10370) <= not a or b;
    layer3_outputs(10371) <= b;
    layer3_outputs(10372) <= not b;
    layer3_outputs(10373) <= a and b;
    layer3_outputs(10374) <= not b;
    layer3_outputs(10375) <= not (a or b);
    layer3_outputs(10376) <= not a;
    layer3_outputs(10377) <= a;
    layer3_outputs(10378) <= not b;
    layer3_outputs(10379) <= b and not a;
    layer3_outputs(10380) <= not (a or b);
    layer3_outputs(10381) <= a or b;
    layer3_outputs(10382) <= not b or a;
    layer3_outputs(10383) <= not (a xor b);
    layer3_outputs(10384) <= not (a and b);
    layer3_outputs(10385) <= not a;
    layer3_outputs(10386) <= a;
    layer3_outputs(10387) <= a;
    layer3_outputs(10388) <= not (a or b);
    layer3_outputs(10389) <= a and not b;
    layer3_outputs(10390) <= b;
    layer3_outputs(10391) <= not b;
    layer3_outputs(10392) <= not b;
    layer3_outputs(10393) <= a;
    layer3_outputs(10394) <= not (a xor b);
    layer3_outputs(10395) <= not (a or b);
    layer3_outputs(10396) <= b and not a;
    layer3_outputs(10397) <= not a;
    layer3_outputs(10398) <= b;
    layer3_outputs(10399) <= not a or b;
    layer3_outputs(10400) <= b and not a;
    layer3_outputs(10401) <= a;
    layer3_outputs(10402) <= b;
    layer3_outputs(10403) <= a or b;
    layer3_outputs(10404) <= a xor b;
    layer3_outputs(10405) <= a;
    layer3_outputs(10406) <= not a;
    layer3_outputs(10407) <= a;
    layer3_outputs(10408) <= not (a and b);
    layer3_outputs(10409) <= not a;
    layer3_outputs(10410) <= b;
    layer3_outputs(10411) <= not (a xor b);
    layer3_outputs(10412) <= not a;
    layer3_outputs(10413) <= b and not a;
    layer3_outputs(10414) <= a;
    layer3_outputs(10415) <= not b;
    layer3_outputs(10416) <= a and b;
    layer3_outputs(10417) <= b;
    layer3_outputs(10418) <= not a or b;
    layer3_outputs(10419) <= b;
    layer3_outputs(10420) <= not (a and b);
    layer3_outputs(10421) <= a and b;
    layer3_outputs(10422) <= not a;
    layer3_outputs(10423) <= a and b;
    layer3_outputs(10424) <= b and not a;
    layer3_outputs(10425) <= a;
    layer3_outputs(10426) <= a;
    layer3_outputs(10427) <= b and not a;
    layer3_outputs(10428) <= not b;
    layer3_outputs(10429) <= b;
    layer3_outputs(10430) <= not a or b;
    layer3_outputs(10431) <= not b;
    layer3_outputs(10432) <= a;
    layer3_outputs(10433) <= not b;
    layer3_outputs(10434) <= b;
    layer3_outputs(10435) <= not (a and b);
    layer3_outputs(10436) <= a and b;
    layer3_outputs(10437) <= not (a or b);
    layer3_outputs(10438) <= '1';
    layer3_outputs(10439) <= not a;
    layer3_outputs(10440) <= a xor b;
    layer3_outputs(10441) <= a and b;
    layer3_outputs(10442) <= not a;
    layer3_outputs(10443) <= not b;
    layer3_outputs(10444) <= b;
    layer3_outputs(10445) <= not (a and b);
    layer3_outputs(10446) <= b and not a;
    layer3_outputs(10447) <= not (a and b);
    layer3_outputs(10448) <= not a or b;
    layer3_outputs(10449) <= not a;
    layer3_outputs(10450) <= not a;
    layer3_outputs(10451) <= not b;
    layer3_outputs(10452) <= b and not a;
    layer3_outputs(10453) <= not a;
    layer3_outputs(10454) <= b and not a;
    layer3_outputs(10455) <= a and b;
    layer3_outputs(10456) <= b;
    layer3_outputs(10457) <= not (a and b);
    layer3_outputs(10458) <= a and b;
    layer3_outputs(10459) <= b and not a;
    layer3_outputs(10460) <= not b or a;
    layer3_outputs(10461) <= not (a or b);
    layer3_outputs(10462) <= not (a xor b);
    layer3_outputs(10463) <= b;
    layer3_outputs(10464) <= not (a xor b);
    layer3_outputs(10465) <= not a;
    layer3_outputs(10466) <= not b or a;
    layer3_outputs(10467) <= not a;
    layer3_outputs(10468) <= a;
    layer3_outputs(10469) <= not (a or b);
    layer3_outputs(10470) <= not (a or b);
    layer3_outputs(10471) <= a;
    layer3_outputs(10472) <= not (a or b);
    layer3_outputs(10473) <= a;
    layer3_outputs(10474) <= not a;
    layer3_outputs(10475) <= not b;
    layer3_outputs(10476) <= not b or a;
    layer3_outputs(10477) <= not (a and b);
    layer3_outputs(10478) <= not (a or b);
    layer3_outputs(10479) <= a or b;
    layer3_outputs(10480) <= a xor b;
    layer3_outputs(10481) <= a;
    layer3_outputs(10482) <= a;
    layer3_outputs(10483) <= not (a and b);
    layer3_outputs(10484) <= not a or b;
    layer3_outputs(10485) <= not a;
    layer3_outputs(10486) <= not a;
    layer3_outputs(10487) <= b;
    layer3_outputs(10488) <= not (a or b);
    layer3_outputs(10489) <= a or b;
    layer3_outputs(10490) <= a xor b;
    layer3_outputs(10491) <= not (a and b);
    layer3_outputs(10492) <= not b or a;
    layer3_outputs(10493) <= a;
    layer3_outputs(10494) <= not (a xor b);
    layer3_outputs(10495) <= a;
    layer3_outputs(10496) <= b;
    layer3_outputs(10497) <= b;
    layer3_outputs(10498) <= not b or a;
    layer3_outputs(10499) <= a xor b;
    layer3_outputs(10500) <= b and not a;
    layer3_outputs(10501) <= a and not b;
    layer3_outputs(10502) <= a and not b;
    layer3_outputs(10503) <= a or b;
    layer3_outputs(10504) <= a and b;
    layer3_outputs(10505) <= b and not a;
    layer3_outputs(10506) <= not b;
    layer3_outputs(10507) <= a xor b;
    layer3_outputs(10508) <= not a;
    layer3_outputs(10509) <= a;
    layer3_outputs(10510) <= not b;
    layer3_outputs(10511) <= a and b;
    layer3_outputs(10512) <= a;
    layer3_outputs(10513) <= a or b;
    layer3_outputs(10514) <= not a or b;
    layer3_outputs(10515) <= not (a and b);
    layer3_outputs(10516) <= not a or b;
    layer3_outputs(10517) <= not (a and b);
    layer3_outputs(10518) <= not a or b;
    layer3_outputs(10519) <= a;
    layer3_outputs(10520) <= not b;
    layer3_outputs(10521) <= a xor b;
    layer3_outputs(10522) <= not (a xor b);
    layer3_outputs(10523) <= not a or b;
    layer3_outputs(10524) <= a;
    layer3_outputs(10525) <= b;
    layer3_outputs(10526) <= a;
    layer3_outputs(10527) <= '0';
    layer3_outputs(10528) <= '1';
    layer3_outputs(10529) <= not (a or b);
    layer3_outputs(10530) <= b and not a;
    layer3_outputs(10531) <= not (a and b);
    layer3_outputs(10532) <= a;
    layer3_outputs(10533) <= not b;
    layer3_outputs(10534) <= a and b;
    layer3_outputs(10535) <= a or b;
    layer3_outputs(10536) <= a and b;
    layer3_outputs(10537) <= b;
    layer3_outputs(10538) <= a and b;
    layer3_outputs(10539) <= not b or a;
    layer3_outputs(10540) <= b and not a;
    layer3_outputs(10541) <= not a or b;
    layer3_outputs(10542) <= not b;
    layer3_outputs(10543) <= b;
    layer3_outputs(10544) <= '1';
    layer3_outputs(10545) <= not (a or b);
    layer3_outputs(10546) <= a;
    layer3_outputs(10547) <= b;
    layer3_outputs(10548) <= a or b;
    layer3_outputs(10549) <= b;
    layer3_outputs(10550) <= b and not a;
    layer3_outputs(10551) <= not b;
    layer3_outputs(10552) <= b;
    layer3_outputs(10553) <= '1';
    layer3_outputs(10554) <= a and not b;
    layer3_outputs(10555) <= not b or a;
    layer3_outputs(10556) <= a;
    layer3_outputs(10557) <= not a or b;
    layer3_outputs(10558) <= a and not b;
    layer3_outputs(10559) <= a and b;
    layer3_outputs(10560) <= not b;
    layer3_outputs(10561) <= not (a or b);
    layer3_outputs(10562) <= b;
    layer3_outputs(10563) <= b and not a;
    layer3_outputs(10564) <= not (a or b);
    layer3_outputs(10565) <= '1';
    layer3_outputs(10566) <= a or b;
    layer3_outputs(10567) <= a xor b;
    layer3_outputs(10568) <= b;
    layer3_outputs(10569) <= not a;
    layer3_outputs(10570) <= not a or b;
    layer3_outputs(10571) <= a;
    layer3_outputs(10572) <= b;
    layer3_outputs(10573) <= not (a or b);
    layer3_outputs(10574) <= b and not a;
    layer3_outputs(10575) <= a or b;
    layer3_outputs(10576) <= a or b;
    layer3_outputs(10577) <= not b;
    layer3_outputs(10578) <= not b;
    layer3_outputs(10579) <= not a;
    layer3_outputs(10580) <= not a;
    layer3_outputs(10581) <= not (a or b);
    layer3_outputs(10582) <= not (a or b);
    layer3_outputs(10583) <= not b;
    layer3_outputs(10584) <= a;
    layer3_outputs(10585) <= not b or a;
    layer3_outputs(10586) <= a and b;
    layer3_outputs(10587) <= not (a xor b);
    layer3_outputs(10588) <= not a or b;
    layer3_outputs(10589) <= a and not b;
    layer3_outputs(10590) <= a;
    layer3_outputs(10591) <= not (a or b);
    layer3_outputs(10592) <= not a;
    layer3_outputs(10593) <= not b;
    layer3_outputs(10594) <= not b;
    layer3_outputs(10595) <= '1';
    layer3_outputs(10596) <= a and b;
    layer3_outputs(10597) <= a and b;
    layer3_outputs(10598) <= a;
    layer3_outputs(10599) <= not b;
    layer3_outputs(10600) <= b;
    layer3_outputs(10601) <= not a;
    layer3_outputs(10602) <= '1';
    layer3_outputs(10603) <= not b;
    layer3_outputs(10604) <= a and b;
    layer3_outputs(10605) <= not (a xor b);
    layer3_outputs(10606) <= not a or b;
    layer3_outputs(10607) <= not a;
    layer3_outputs(10608) <= not (a and b);
    layer3_outputs(10609) <= a;
    layer3_outputs(10610) <= a;
    layer3_outputs(10611) <= not b;
    layer3_outputs(10612) <= a and b;
    layer3_outputs(10613) <= not (a and b);
    layer3_outputs(10614) <= a and not b;
    layer3_outputs(10615) <= not a or b;
    layer3_outputs(10616) <= not b or a;
    layer3_outputs(10617) <= a;
    layer3_outputs(10618) <= not a or b;
    layer3_outputs(10619) <= not a;
    layer3_outputs(10620) <= b and not a;
    layer3_outputs(10621) <= not a;
    layer3_outputs(10622) <= not a or b;
    layer3_outputs(10623) <= '1';
    layer3_outputs(10624) <= not a;
    layer3_outputs(10625) <= not (a and b);
    layer3_outputs(10626) <= not (a or b);
    layer3_outputs(10627) <= a and b;
    layer3_outputs(10628) <= not b;
    layer3_outputs(10629) <= not a;
    layer3_outputs(10630) <= not a;
    layer3_outputs(10631) <= a xor b;
    layer3_outputs(10632) <= b;
    layer3_outputs(10633) <= a;
    layer3_outputs(10634) <= a or b;
    layer3_outputs(10635) <= not b or a;
    layer3_outputs(10636) <= not a;
    layer3_outputs(10637) <= a;
    layer3_outputs(10638) <= not a;
    layer3_outputs(10639) <= '0';
    layer3_outputs(10640) <= not b or a;
    layer3_outputs(10641) <= a;
    layer3_outputs(10642) <= a and not b;
    layer3_outputs(10643) <= '0';
    layer3_outputs(10644) <= a and b;
    layer3_outputs(10645) <= not (a xor b);
    layer3_outputs(10646) <= not b or a;
    layer3_outputs(10647) <= a or b;
    layer3_outputs(10648) <= a or b;
    layer3_outputs(10649) <= a and not b;
    layer3_outputs(10650) <= not b;
    layer3_outputs(10651) <= not b or a;
    layer3_outputs(10652) <= not (a or b);
    layer3_outputs(10653) <= not b;
    layer3_outputs(10654) <= b;
    layer3_outputs(10655) <= not a;
    layer3_outputs(10656) <= not a;
    layer3_outputs(10657) <= a or b;
    layer3_outputs(10658) <= a and b;
    layer3_outputs(10659) <= b;
    layer3_outputs(10660) <= not (a or b);
    layer3_outputs(10661) <= a;
    layer3_outputs(10662) <= not b or a;
    layer3_outputs(10663) <= not b;
    layer3_outputs(10664) <= not (a xor b);
    layer3_outputs(10665) <= '0';
    layer3_outputs(10666) <= not a;
    layer3_outputs(10667) <= a and not b;
    layer3_outputs(10668) <= b and not a;
    layer3_outputs(10669) <= not b;
    layer3_outputs(10670) <= a and not b;
    layer3_outputs(10671) <= a;
    layer3_outputs(10672) <= '1';
    layer3_outputs(10673) <= '0';
    layer3_outputs(10674) <= not b or a;
    layer3_outputs(10675) <= a and b;
    layer3_outputs(10676) <= not a;
    layer3_outputs(10677) <= not (a and b);
    layer3_outputs(10678) <= a or b;
    layer3_outputs(10679) <= a;
    layer3_outputs(10680) <= '0';
    layer3_outputs(10681) <= not a;
    layer3_outputs(10682) <= not b;
    layer3_outputs(10683) <= a;
    layer3_outputs(10684) <= not (a or b);
    layer3_outputs(10685) <= not b;
    layer3_outputs(10686) <= a and b;
    layer3_outputs(10687) <= b;
    layer3_outputs(10688) <= not (a and b);
    layer3_outputs(10689) <= not (a and b);
    layer3_outputs(10690) <= b and not a;
    layer3_outputs(10691) <= '1';
    layer3_outputs(10692) <= not b or a;
    layer3_outputs(10693) <= a xor b;
    layer3_outputs(10694) <= a;
    layer3_outputs(10695) <= a;
    layer3_outputs(10696) <= b and not a;
    layer3_outputs(10697) <= a xor b;
    layer3_outputs(10698) <= not (a and b);
    layer3_outputs(10699) <= '1';
    layer3_outputs(10700) <= not (a and b);
    layer3_outputs(10701) <= not a;
    layer3_outputs(10702) <= a;
    layer3_outputs(10703) <= not (a xor b);
    layer3_outputs(10704) <= a or b;
    layer3_outputs(10705) <= a;
    layer3_outputs(10706) <= not b or a;
    layer3_outputs(10707) <= not b or a;
    layer3_outputs(10708) <= a;
    layer3_outputs(10709) <= not (a or b);
    layer3_outputs(10710) <= not a;
    layer3_outputs(10711) <= '1';
    layer3_outputs(10712) <= b;
    layer3_outputs(10713) <= b;
    layer3_outputs(10714) <= '0';
    layer3_outputs(10715) <= a;
    layer3_outputs(10716) <= a xor b;
    layer3_outputs(10717) <= b and not a;
    layer3_outputs(10718) <= a and not b;
    layer3_outputs(10719) <= '1';
    layer3_outputs(10720) <= not a;
    layer3_outputs(10721) <= not a;
    layer3_outputs(10722) <= b;
    layer3_outputs(10723) <= '1';
    layer3_outputs(10724) <= not b or a;
    layer3_outputs(10725) <= not a;
    layer3_outputs(10726) <= not b;
    layer3_outputs(10727) <= not a;
    layer3_outputs(10728) <= '0';
    layer3_outputs(10729) <= not (a and b);
    layer3_outputs(10730) <= a xor b;
    layer3_outputs(10731) <= b and not a;
    layer3_outputs(10732) <= '1';
    layer3_outputs(10733) <= not b;
    layer3_outputs(10734) <= a or b;
    layer3_outputs(10735) <= not a;
    layer3_outputs(10736) <= a and b;
    layer3_outputs(10737) <= not (a or b);
    layer3_outputs(10738) <= b and not a;
    layer3_outputs(10739) <= b;
    layer3_outputs(10740) <= not (a xor b);
    layer3_outputs(10741) <= not (a or b);
    layer3_outputs(10742) <= not b;
    layer3_outputs(10743) <= a and not b;
    layer3_outputs(10744) <= not a;
    layer3_outputs(10745) <= a and not b;
    layer3_outputs(10746) <= not a or b;
    layer3_outputs(10747) <= a and b;
    layer3_outputs(10748) <= not b;
    layer3_outputs(10749) <= a or b;
    layer3_outputs(10750) <= not (a xor b);
    layer3_outputs(10751) <= not (a xor b);
    layer3_outputs(10752) <= not b or a;
    layer3_outputs(10753) <= a and b;
    layer3_outputs(10754) <= '1';
    layer3_outputs(10755) <= b;
    layer3_outputs(10756) <= not b or a;
    layer3_outputs(10757) <= b;
    layer3_outputs(10758) <= not b;
    layer3_outputs(10759) <= '1';
    layer3_outputs(10760) <= a and b;
    layer3_outputs(10761) <= b and not a;
    layer3_outputs(10762) <= not (a or b);
    layer3_outputs(10763) <= b;
    layer3_outputs(10764) <= not (a and b);
    layer3_outputs(10765) <= a and not b;
    layer3_outputs(10766) <= '0';
    layer3_outputs(10767) <= b and not a;
    layer3_outputs(10768) <= not (a or b);
    layer3_outputs(10769) <= a and b;
    layer3_outputs(10770) <= b and not a;
    layer3_outputs(10771) <= not b;
    layer3_outputs(10772) <= a and not b;
    layer3_outputs(10773) <= not b;
    layer3_outputs(10774) <= a;
    layer3_outputs(10775) <= not a;
    layer3_outputs(10776) <= a;
    layer3_outputs(10777) <= b;
    layer3_outputs(10778) <= not b;
    layer3_outputs(10779) <= '0';
    layer3_outputs(10780) <= not b;
    layer3_outputs(10781) <= not b or a;
    layer3_outputs(10782) <= a and b;
    layer3_outputs(10783) <= b;
    layer3_outputs(10784) <= a and not b;
    layer3_outputs(10785) <= '0';
    layer3_outputs(10786) <= '1';
    layer3_outputs(10787) <= not (a or b);
    layer3_outputs(10788) <= not a or b;
    layer3_outputs(10789) <= not b;
    layer3_outputs(10790) <= not b;
    layer3_outputs(10791) <= b and not a;
    layer3_outputs(10792) <= b;
    layer3_outputs(10793) <= not (a or b);
    layer3_outputs(10794) <= a and not b;
    layer3_outputs(10795) <= not (a or b);
    layer3_outputs(10796) <= not b;
    layer3_outputs(10797) <= not a;
    layer3_outputs(10798) <= not (a and b);
    layer3_outputs(10799) <= not a or b;
    layer3_outputs(10800) <= b;
    layer3_outputs(10801) <= not a;
    layer3_outputs(10802) <= b;
    layer3_outputs(10803) <= a xor b;
    layer3_outputs(10804) <= not b;
    layer3_outputs(10805) <= '1';
    layer3_outputs(10806) <= not (a xor b);
    layer3_outputs(10807) <= not b;
    layer3_outputs(10808) <= a and b;
    layer3_outputs(10809) <= b and not a;
    layer3_outputs(10810) <= b;
    layer3_outputs(10811) <= not b or a;
    layer3_outputs(10812) <= not b;
    layer3_outputs(10813) <= '1';
    layer3_outputs(10814) <= b and not a;
    layer3_outputs(10815) <= a;
    layer3_outputs(10816) <= a xor b;
    layer3_outputs(10817) <= not b or a;
    layer3_outputs(10818) <= not (a or b);
    layer3_outputs(10819) <= not b;
    layer3_outputs(10820) <= b;
    layer3_outputs(10821) <= not a;
    layer3_outputs(10822) <= a and not b;
    layer3_outputs(10823) <= not (a or b);
    layer3_outputs(10824) <= a and b;
    layer3_outputs(10825) <= a or b;
    layer3_outputs(10826) <= not b or a;
    layer3_outputs(10827) <= not (a or b);
    layer3_outputs(10828) <= not b or a;
    layer3_outputs(10829) <= a or b;
    layer3_outputs(10830) <= b and not a;
    layer3_outputs(10831) <= not b;
    layer3_outputs(10832) <= not (a xor b);
    layer3_outputs(10833) <= not (a and b);
    layer3_outputs(10834) <= a;
    layer3_outputs(10835) <= b;
    layer3_outputs(10836) <= a;
    layer3_outputs(10837) <= a and b;
    layer3_outputs(10838) <= not b;
    layer3_outputs(10839) <= a and b;
    layer3_outputs(10840) <= not a;
    layer3_outputs(10841) <= not b;
    layer3_outputs(10842) <= not b;
    layer3_outputs(10843) <= not (a or b);
    layer3_outputs(10844) <= not b;
    layer3_outputs(10845) <= b;
    layer3_outputs(10846) <= not a or b;
    layer3_outputs(10847) <= '1';
    layer3_outputs(10848) <= a xor b;
    layer3_outputs(10849) <= not b;
    layer3_outputs(10850) <= a and not b;
    layer3_outputs(10851) <= a and not b;
    layer3_outputs(10852) <= not a;
    layer3_outputs(10853) <= a and not b;
    layer3_outputs(10854) <= a;
    layer3_outputs(10855) <= b;
    layer3_outputs(10856) <= b;
    layer3_outputs(10857) <= not b or a;
    layer3_outputs(10858) <= a and b;
    layer3_outputs(10859) <= not a or b;
    layer3_outputs(10860) <= not b;
    layer3_outputs(10861) <= a xor b;
    layer3_outputs(10862) <= a;
    layer3_outputs(10863) <= not (a or b);
    layer3_outputs(10864) <= not (a or b);
    layer3_outputs(10865) <= not a or b;
    layer3_outputs(10866) <= not b;
    layer3_outputs(10867) <= not a;
    layer3_outputs(10868) <= not (a or b);
    layer3_outputs(10869) <= a or b;
    layer3_outputs(10870) <= '0';
    layer3_outputs(10871) <= a and not b;
    layer3_outputs(10872) <= not (a and b);
    layer3_outputs(10873) <= not (a xor b);
    layer3_outputs(10874) <= a;
    layer3_outputs(10875) <= a or b;
    layer3_outputs(10876) <= not a;
    layer3_outputs(10877) <= not a;
    layer3_outputs(10878) <= a xor b;
    layer3_outputs(10879) <= not a;
    layer3_outputs(10880) <= a or b;
    layer3_outputs(10881) <= b and not a;
    layer3_outputs(10882) <= a;
    layer3_outputs(10883) <= not (a xor b);
    layer3_outputs(10884) <= '0';
    layer3_outputs(10885) <= not b;
    layer3_outputs(10886) <= '0';
    layer3_outputs(10887) <= a;
    layer3_outputs(10888) <= '0';
    layer3_outputs(10889) <= not (a and b);
    layer3_outputs(10890) <= not (a xor b);
    layer3_outputs(10891) <= a and b;
    layer3_outputs(10892) <= a and not b;
    layer3_outputs(10893) <= a and not b;
    layer3_outputs(10894) <= a;
    layer3_outputs(10895) <= not a or b;
    layer3_outputs(10896) <= not (a and b);
    layer3_outputs(10897) <= not a or b;
    layer3_outputs(10898) <= a xor b;
    layer3_outputs(10899) <= not a;
    layer3_outputs(10900) <= b and not a;
    layer3_outputs(10901) <= a xor b;
    layer3_outputs(10902) <= a and not b;
    layer3_outputs(10903) <= not (a or b);
    layer3_outputs(10904) <= '0';
    layer3_outputs(10905) <= not (a or b);
    layer3_outputs(10906) <= a or b;
    layer3_outputs(10907) <= a and b;
    layer3_outputs(10908) <= '0';
    layer3_outputs(10909) <= not a;
    layer3_outputs(10910) <= '1';
    layer3_outputs(10911) <= not a;
    layer3_outputs(10912) <= a;
    layer3_outputs(10913) <= not (a or b);
    layer3_outputs(10914) <= a or b;
    layer3_outputs(10915) <= a and b;
    layer3_outputs(10916) <= not b or a;
    layer3_outputs(10917) <= a or b;
    layer3_outputs(10918) <= a or b;
    layer3_outputs(10919) <= not a;
    layer3_outputs(10920) <= a;
    layer3_outputs(10921) <= b and not a;
    layer3_outputs(10922) <= b;
    layer3_outputs(10923) <= b and not a;
    layer3_outputs(10924) <= '0';
    layer3_outputs(10925) <= not (a or b);
    layer3_outputs(10926) <= not b or a;
    layer3_outputs(10927) <= not b or a;
    layer3_outputs(10928) <= not b;
    layer3_outputs(10929) <= not (a and b);
    layer3_outputs(10930) <= not b;
    layer3_outputs(10931) <= b;
    layer3_outputs(10932) <= a and b;
    layer3_outputs(10933) <= a and b;
    layer3_outputs(10934) <= not a;
    layer3_outputs(10935) <= b;
    layer3_outputs(10936) <= not a;
    layer3_outputs(10937) <= b;
    layer3_outputs(10938) <= not (a and b);
    layer3_outputs(10939) <= not a;
    layer3_outputs(10940) <= a;
    layer3_outputs(10941) <= b;
    layer3_outputs(10942) <= b;
    layer3_outputs(10943) <= not (a xor b);
    layer3_outputs(10944) <= b;
    layer3_outputs(10945) <= not a;
    layer3_outputs(10946) <= a or b;
    layer3_outputs(10947) <= not b or a;
    layer3_outputs(10948) <= not (a and b);
    layer3_outputs(10949) <= a;
    layer3_outputs(10950) <= not b;
    layer3_outputs(10951) <= not (a xor b);
    layer3_outputs(10952) <= a;
    layer3_outputs(10953) <= '0';
    layer3_outputs(10954) <= a and b;
    layer3_outputs(10955) <= not a;
    layer3_outputs(10956) <= a or b;
    layer3_outputs(10957) <= a;
    layer3_outputs(10958) <= not (a or b);
    layer3_outputs(10959) <= not b or a;
    layer3_outputs(10960) <= not a or b;
    layer3_outputs(10961) <= not (a and b);
    layer3_outputs(10962) <= a;
    layer3_outputs(10963) <= not b;
    layer3_outputs(10964) <= b and not a;
    layer3_outputs(10965) <= a or b;
    layer3_outputs(10966) <= '1';
    layer3_outputs(10967) <= a and not b;
    layer3_outputs(10968) <= a and b;
    layer3_outputs(10969) <= a or b;
    layer3_outputs(10970) <= b and not a;
    layer3_outputs(10971) <= not a or b;
    layer3_outputs(10972) <= '0';
    layer3_outputs(10973) <= a and not b;
    layer3_outputs(10974) <= a and not b;
    layer3_outputs(10975) <= not a or b;
    layer3_outputs(10976) <= '1';
    layer3_outputs(10977) <= a and b;
    layer3_outputs(10978) <= not a or b;
    layer3_outputs(10979) <= a xor b;
    layer3_outputs(10980) <= not b or a;
    layer3_outputs(10981) <= not b;
    layer3_outputs(10982) <= a and b;
    layer3_outputs(10983) <= not a;
    layer3_outputs(10984) <= '0';
    layer3_outputs(10985) <= not (a xor b);
    layer3_outputs(10986) <= a;
    layer3_outputs(10987) <= not b;
    layer3_outputs(10988) <= a and not b;
    layer3_outputs(10989) <= not (a and b);
    layer3_outputs(10990) <= not a or b;
    layer3_outputs(10991) <= b;
    layer3_outputs(10992) <= not b or a;
    layer3_outputs(10993) <= '0';
    layer3_outputs(10994) <= a and b;
    layer3_outputs(10995) <= not b;
    layer3_outputs(10996) <= a and not b;
    layer3_outputs(10997) <= b and not a;
    layer3_outputs(10998) <= not a;
    layer3_outputs(10999) <= a or b;
    layer3_outputs(11000) <= not b;
    layer3_outputs(11001) <= a and not b;
    layer3_outputs(11002) <= not a or b;
    layer3_outputs(11003) <= a and not b;
    layer3_outputs(11004) <= a xor b;
    layer3_outputs(11005) <= not a or b;
    layer3_outputs(11006) <= b;
    layer3_outputs(11007) <= not (a and b);
    layer3_outputs(11008) <= a xor b;
    layer3_outputs(11009) <= b;
    layer3_outputs(11010) <= b and not a;
    layer3_outputs(11011) <= a or b;
    layer3_outputs(11012) <= '1';
    layer3_outputs(11013) <= not a or b;
    layer3_outputs(11014) <= a;
    layer3_outputs(11015) <= not (a and b);
    layer3_outputs(11016) <= not (a and b);
    layer3_outputs(11017) <= '0';
    layer3_outputs(11018) <= not b;
    layer3_outputs(11019) <= b;
    layer3_outputs(11020) <= b;
    layer3_outputs(11021) <= not (a and b);
    layer3_outputs(11022) <= not (a or b);
    layer3_outputs(11023) <= a or b;
    layer3_outputs(11024) <= not a;
    layer3_outputs(11025) <= not (a or b);
    layer3_outputs(11026) <= a;
    layer3_outputs(11027) <= not b;
    layer3_outputs(11028) <= not b;
    layer3_outputs(11029) <= a;
    layer3_outputs(11030) <= a and not b;
    layer3_outputs(11031) <= a xor b;
    layer3_outputs(11032) <= b and not a;
    layer3_outputs(11033) <= not a;
    layer3_outputs(11034) <= a and not b;
    layer3_outputs(11035) <= not b or a;
    layer3_outputs(11036) <= a xor b;
    layer3_outputs(11037) <= b;
    layer3_outputs(11038) <= not (a or b);
    layer3_outputs(11039) <= not b or a;
    layer3_outputs(11040) <= a and b;
    layer3_outputs(11041) <= not (a or b);
    layer3_outputs(11042) <= a and not b;
    layer3_outputs(11043) <= a;
    layer3_outputs(11044) <= '0';
    layer3_outputs(11045) <= a and b;
    layer3_outputs(11046) <= '0';
    layer3_outputs(11047) <= not a;
    layer3_outputs(11048) <= a;
    layer3_outputs(11049) <= a;
    layer3_outputs(11050) <= a and not b;
    layer3_outputs(11051) <= not (a and b);
    layer3_outputs(11052) <= not b;
    layer3_outputs(11053) <= b;
    layer3_outputs(11054) <= not b;
    layer3_outputs(11055) <= not a or b;
    layer3_outputs(11056) <= a or b;
    layer3_outputs(11057) <= not a;
    layer3_outputs(11058) <= not (a or b);
    layer3_outputs(11059) <= a and not b;
    layer3_outputs(11060) <= b;
    layer3_outputs(11061) <= not b;
    layer3_outputs(11062) <= not b;
    layer3_outputs(11063) <= a;
    layer3_outputs(11064) <= not (a and b);
    layer3_outputs(11065) <= a and b;
    layer3_outputs(11066) <= b;
    layer3_outputs(11067) <= a xor b;
    layer3_outputs(11068) <= not b or a;
    layer3_outputs(11069) <= b and not a;
    layer3_outputs(11070) <= not a;
    layer3_outputs(11071) <= a and b;
    layer3_outputs(11072) <= a xor b;
    layer3_outputs(11073) <= not (a xor b);
    layer3_outputs(11074) <= a and b;
    layer3_outputs(11075) <= not (a or b);
    layer3_outputs(11076) <= a xor b;
    layer3_outputs(11077) <= not (a or b);
    layer3_outputs(11078) <= a xor b;
    layer3_outputs(11079) <= a or b;
    layer3_outputs(11080) <= not a;
    layer3_outputs(11081) <= a;
    layer3_outputs(11082) <= a xor b;
    layer3_outputs(11083) <= b;
    layer3_outputs(11084) <= not (a or b);
    layer3_outputs(11085) <= not (a or b);
    layer3_outputs(11086) <= not (a and b);
    layer3_outputs(11087) <= not b;
    layer3_outputs(11088) <= '0';
    layer3_outputs(11089) <= a and b;
    layer3_outputs(11090) <= not (a and b);
    layer3_outputs(11091) <= b and not a;
    layer3_outputs(11092) <= not b;
    layer3_outputs(11093) <= not b;
    layer3_outputs(11094) <= a xor b;
    layer3_outputs(11095) <= not b or a;
    layer3_outputs(11096) <= a xor b;
    layer3_outputs(11097) <= a;
    layer3_outputs(11098) <= b;
    layer3_outputs(11099) <= not (a and b);
    layer3_outputs(11100) <= not (a or b);
    layer3_outputs(11101) <= not a;
    layer3_outputs(11102) <= not (a and b);
    layer3_outputs(11103) <= not a or b;
    layer3_outputs(11104) <= not (a and b);
    layer3_outputs(11105) <= b;
    layer3_outputs(11106) <= '0';
    layer3_outputs(11107) <= a;
    layer3_outputs(11108) <= not b or a;
    layer3_outputs(11109) <= not a;
    layer3_outputs(11110) <= not (a xor b);
    layer3_outputs(11111) <= not (a xor b);
    layer3_outputs(11112) <= a and b;
    layer3_outputs(11113) <= not a;
    layer3_outputs(11114) <= a;
    layer3_outputs(11115) <= not b;
    layer3_outputs(11116) <= not (a xor b);
    layer3_outputs(11117) <= a and not b;
    layer3_outputs(11118) <= not a or b;
    layer3_outputs(11119) <= not (a xor b);
    layer3_outputs(11120) <= b;
    layer3_outputs(11121) <= a and not b;
    layer3_outputs(11122) <= not (a xor b);
    layer3_outputs(11123) <= not b;
    layer3_outputs(11124) <= a xor b;
    layer3_outputs(11125) <= not b or a;
    layer3_outputs(11126) <= not (a xor b);
    layer3_outputs(11127) <= not (a or b);
    layer3_outputs(11128) <= not a;
    layer3_outputs(11129) <= not a or b;
    layer3_outputs(11130) <= not a or b;
    layer3_outputs(11131) <= not (a xor b);
    layer3_outputs(11132) <= not a;
    layer3_outputs(11133) <= not (a and b);
    layer3_outputs(11134) <= not (a or b);
    layer3_outputs(11135) <= a xor b;
    layer3_outputs(11136) <= not (a or b);
    layer3_outputs(11137) <= '1';
    layer3_outputs(11138) <= a or b;
    layer3_outputs(11139) <= '1';
    layer3_outputs(11140) <= not b;
    layer3_outputs(11141) <= b and not a;
    layer3_outputs(11142) <= a and not b;
    layer3_outputs(11143) <= b;
    layer3_outputs(11144) <= b;
    layer3_outputs(11145) <= not a;
    layer3_outputs(11146) <= not b or a;
    layer3_outputs(11147) <= a and b;
    layer3_outputs(11148) <= not b or a;
    layer3_outputs(11149) <= b;
    layer3_outputs(11150) <= '1';
    layer3_outputs(11151) <= a and b;
    layer3_outputs(11152) <= not b;
    layer3_outputs(11153) <= a;
    layer3_outputs(11154) <= not (a and b);
    layer3_outputs(11155) <= not (a and b);
    layer3_outputs(11156) <= a and b;
    layer3_outputs(11157) <= b and not a;
    layer3_outputs(11158) <= not (a and b);
    layer3_outputs(11159) <= a and b;
    layer3_outputs(11160) <= not b;
    layer3_outputs(11161) <= b;
    layer3_outputs(11162) <= not b or a;
    layer3_outputs(11163) <= b;
    layer3_outputs(11164) <= a xor b;
    layer3_outputs(11165) <= not (a and b);
    layer3_outputs(11166) <= a and not b;
    layer3_outputs(11167) <= not (a or b);
    layer3_outputs(11168) <= a or b;
    layer3_outputs(11169) <= not b or a;
    layer3_outputs(11170) <= not b or a;
    layer3_outputs(11171) <= a xor b;
    layer3_outputs(11172) <= a xor b;
    layer3_outputs(11173) <= not b;
    layer3_outputs(11174) <= a;
    layer3_outputs(11175) <= b and not a;
    layer3_outputs(11176) <= b and not a;
    layer3_outputs(11177) <= not b or a;
    layer3_outputs(11178) <= b;
    layer3_outputs(11179) <= '0';
    layer3_outputs(11180) <= a xor b;
    layer3_outputs(11181) <= a and not b;
    layer3_outputs(11182) <= not a or b;
    layer3_outputs(11183) <= b;
    layer3_outputs(11184) <= not a or b;
    layer3_outputs(11185) <= not (a xor b);
    layer3_outputs(11186) <= not (a or b);
    layer3_outputs(11187) <= a or b;
    layer3_outputs(11188) <= not (a or b);
    layer3_outputs(11189) <= b;
    layer3_outputs(11190) <= not a or b;
    layer3_outputs(11191) <= not b;
    layer3_outputs(11192) <= not b or a;
    layer3_outputs(11193) <= not b or a;
    layer3_outputs(11194) <= not a or b;
    layer3_outputs(11195) <= a and not b;
    layer3_outputs(11196) <= not a or b;
    layer3_outputs(11197) <= a and not b;
    layer3_outputs(11198) <= not b or a;
    layer3_outputs(11199) <= a;
    layer3_outputs(11200) <= '0';
    layer3_outputs(11201) <= a;
    layer3_outputs(11202) <= a or b;
    layer3_outputs(11203) <= not (a or b);
    layer3_outputs(11204) <= not a;
    layer3_outputs(11205) <= not b or a;
    layer3_outputs(11206) <= not b or a;
    layer3_outputs(11207) <= not (a and b);
    layer3_outputs(11208) <= not (a or b);
    layer3_outputs(11209) <= not (a and b);
    layer3_outputs(11210) <= a;
    layer3_outputs(11211) <= not a;
    layer3_outputs(11212) <= a and not b;
    layer3_outputs(11213) <= b and not a;
    layer3_outputs(11214) <= a or b;
    layer3_outputs(11215) <= not (a xor b);
    layer3_outputs(11216) <= b;
    layer3_outputs(11217) <= a and not b;
    layer3_outputs(11218) <= b and not a;
    layer3_outputs(11219) <= a or b;
    layer3_outputs(11220) <= b;
    layer3_outputs(11221) <= not a;
    layer3_outputs(11222) <= not (a xor b);
    layer3_outputs(11223) <= not (a or b);
    layer3_outputs(11224) <= b;
    layer3_outputs(11225) <= a and not b;
    layer3_outputs(11226) <= not a or b;
    layer3_outputs(11227) <= not (a and b);
    layer3_outputs(11228) <= a and not b;
    layer3_outputs(11229) <= not a;
    layer3_outputs(11230) <= '0';
    layer3_outputs(11231) <= a;
    layer3_outputs(11232) <= a;
    layer3_outputs(11233) <= not b or a;
    layer3_outputs(11234) <= not (a or b);
    layer3_outputs(11235) <= not (a and b);
    layer3_outputs(11236) <= b;
    layer3_outputs(11237) <= '1';
    layer3_outputs(11238) <= a;
    layer3_outputs(11239) <= a or b;
    layer3_outputs(11240) <= a;
    layer3_outputs(11241) <= a and b;
    layer3_outputs(11242) <= not (a and b);
    layer3_outputs(11243) <= a;
    layer3_outputs(11244) <= a;
    layer3_outputs(11245) <= not a;
    layer3_outputs(11246) <= a;
    layer3_outputs(11247) <= not (a and b);
    layer3_outputs(11248) <= a and b;
    layer3_outputs(11249) <= not a or b;
    layer3_outputs(11250) <= a;
    layer3_outputs(11251) <= a or b;
    layer3_outputs(11252) <= not (a and b);
    layer3_outputs(11253) <= not b or a;
    layer3_outputs(11254) <= not (a xor b);
    layer3_outputs(11255) <= not b;
    layer3_outputs(11256) <= a;
    layer3_outputs(11257) <= not a;
    layer3_outputs(11258) <= not b;
    layer3_outputs(11259) <= b;
    layer3_outputs(11260) <= not a or b;
    layer3_outputs(11261) <= not (a xor b);
    layer3_outputs(11262) <= not b;
    layer3_outputs(11263) <= a;
    layer3_outputs(11264) <= b;
    layer3_outputs(11265) <= b and not a;
    layer3_outputs(11266) <= b;
    layer3_outputs(11267) <= a and b;
    layer3_outputs(11268) <= not (a or b);
    layer3_outputs(11269) <= '0';
    layer3_outputs(11270) <= b;
    layer3_outputs(11271) <= not (a and b);
    layer3_outputs(11272) <= a;
    layer3_outputs(11273) <= not b or a;
    layer3_outputs(11274) <= not b;
    layer3_outputs(11275) <= not b or a;
    layer3_outputs(11276) <= not b;
    layer3_outputs(11277) <= a;
    layer3_outputs(11278) <= '0';
    layer3_outputs(11279) <= a and b;
    layer3_outputs(11280) <= a and b;
    layer3_outputs(11281) <= a and not b;
    layer3_outputs(11282) <= not a;
    layer3_outputs(11283) <= '1';
    layer3_outputs(11284) <= not b;
    layer3_outputs(11285) <= '1';
    layer3_outputs(11286) <= a xor b;
    layer3_outputs(11287) <= not b;
    layer3_outputs(11288) <= a;
    layer3_outputs(11289) <= a and b;
    layer3_outputs(11290) <= b;
    layer3_outputs(11291) <= a;
    layer3_outputs(11292) <= a;
    layer3_outputs(11293) <= a;
    layer3_outputs(11294) <= not a or b;
    layer3_outputs(11295) <= b;
    layer3_outputs(11296) <= b;
    layer3_outputs(11297) <= not b or a;
    layer3_outputs(11298) <= not b or a;
    layer3_outputs(11299) <= '1';
    layer3_outputs(11300) <= not a;
    layer3_outputs(11301) <= a and b;
    layer3_outputs(11302) <= not (a and b);
    layer3_outputs(11303) <= '0';
    layer3_outputs(11304) <= not b;
    layer3_outputs(11305) <= not b;
    layer3_outputs(11306) <= '1';
    layer3_outputs(11307) <= a or b;
    layer3_outputs(11308) <= a and not b;
    layer3_outputs(11309) <= not (a or b);
    layer3_outputs(11310) <= b;
    layer3_outputs(11311) <= a or b;
    layer3_outputs(11312) <= a;
    layer3_outputs(11313) <= a and not b;
    layer3_outputs(11314) <= not (a and b);
    layer3_outputs(11315) <= a;
    layer3_outputs(11316) <= a;
    layer3_outputs(11317) <= '0';
    layer3_outputs(11318) <= a and b;
    layer3_outputs(11319) <= b;
    layer3_outputs(11320) <= not (a or b);
    layer3_outputs(11321) <= a and not b;
    layer3_outputs(11322) <= not (a or b);
    layer3_outputs(11323) <= b and not a;
    layer3_outputs(11324) <= not (a and b);
    layer3_outputs(11325) <= b and not a;
    layer3_outputs(11326) <= not b or a;
    layer3_outputs(11327) <= b;
    layer3_outputs(11328) <= b and not a;
    layer3_outputs(11329) <= not b;
    layer3_outputs(11330) <= a;
    layer3_outputs(11331) <= not a;
    layer3_outputs(11332) <= not a or b;
    layer3_outputs(11333) <= not a or b;
    layer3_outputs(11334) <= not b;
    layer3_outputs(11335) <= '1';
    layer3_outputs(11336) <= not (a xor b);
    layer3_outputs(11337) <= not a;
    layer3_outputs(11338) <= not b;
    layer3_outputs(11339) <= not (a or b);
    layer3_outputs(11340) <= not (a and b);
    layer3_outputs(11341) <= not a;
    layer3_outputs(11342) <= not a or b;
    layer3_outputs(11343) <= not a;
    layer3_outputs(11344) <= not (a or b);
    layer3_outputs(11345) <= a;
    layer3_outputs(11346) <= b;
    layer3_outputs(11347) <= b;
    layer3_outputs(11348) <= not a;
    layer3_outputs(11349) <= not a;
    layer3_outputs(11350) <= a;
    layer3_outputs(11351) <= not b or a;
    layer3_outputs(11352) <= a or b;
    layer3_outputs(11353) <= a and not b;
    layer3_outputs(11354) <= a and not b;
    layer3_outputs(11355) <= not a or b;
    layer3_outputs(11356) <= a;
    layer3_outputs(11357) <= not a;
    layer3_outputs(11358) <= not (a and b);
    layer3_outputs(11359) <= not (a and b);
    layer3_outputs(11360) <= not b;
    layer3_outputs(11361) <= not b;
    layer3_outputs(11362) <= not a;
    layer3_outputs(11363) <= not b;
    layer3_outputs(11364) <= not (a and b);
    layer3_outputs(11365) <= not a or b;
    layer3_outputs(11366) <= b;
    layer3_outputs(11367) <= b and not a;
    layer3_outputs(11368) <= not (a and b);
    layer3_outputs(11369) <= a and not b;
    layer3_outputs(11370) <= '0';
    layer3_outputs(11371) <= a and b;
    layer3_outputs(11372) <= not b;
    layer3_outputs(11373) <= a and not b;
    layer3_outputs(11374) <= not a;
    layer3_outputs(11375) <= a or b;
    layer3_outputs(11376) <= a and not b;
    layer3_outputs(11377) <= b;
    layer3_outputs(11378) <= b;
    layer3_outputs(11379) <= not (a xor b);
    layer3_outputs(11380) <= '1';
    layer3_outputs(11381) <= not b or a;
    layer3_outputs(11382) <= not a or b;
    layer3_outputs(11383) <= not a or b;
    layer3_outputs(11384) <= a and not b;
    layer3_outputs(11385) <= b and not a;
    layer3_outputs(11386) <= not (a or b);
    layer3_outputs(11387) <= not b or a;
    layer3_outputs(11388) <= b;
    layer3_outputs(11389) <= not a;
    layer3_outputs(11390) <= not b;
    layer3_outputs(11391) <= not b or a;
    layer3_outputs(11392) <= a and b;
    layer3_outputs(11393) <= a xor b;
    layer3_outputs(11394) <= not b;
    layer3_outputs(11395) <= not (a and b);
    layer3_outputs(11396) <= not b;
    layer3_outputs(11397) <= a and not b;
    layer3_outputs(11398) <= not a;
    layer3_outputs(11399) <= a;
    layer3_outputs(11400) <= not b;
    layer3_outputs(11401) <= not a;
    layer3_outputs(11402) <= a xor b;
    layer3_outputs(11403) <= a and not b;
    layer3_outputs(11404) <= a xor b;
    layer3_outputs(11405) <= '1';
    layer3_outputs(11406) <= not b;
    layer3_outputs(11407) <= not a or b;
    layer3_outputs(11408) <= not (a or b);
    layer3_outputs(11409) <= a or b;
    layer3_outputs(11410) <= not b or a;
    layer3_outputs(11411) <= a and not b;
    layer3_outputs(11412) <= b and not a;
    layer3_outputs(11413) <= a;
    layer3_outputs(11414) <= not b;
    layer3_outputs(11415) <= not b or a;
    layer3_outputs(11416) <= a and b;
    layer3_outputs(11417) <= '0';
    layer3_outputs(11418) <= not a;
    layer3_outputs(11419) <= not a;
    layer3_outputs(11420) <= b;
    layer3_outputs(11421) <= a;
    layer3_outputs(11422) <= not (a xor b);
    layer3_outputs(11423) <= a;
    layer3_outputs(11424) <= a xor b;
    layer3_outputs(11425) <= a or b;
    layer3_outputs(11426) <= not b;
    layer3_outputs(11427) <= a xor b;
    layer3_outputs(11428) <= b;
    layer3_outputs(11429) <= b;
    layer3_outputs(11430) <= a or b;
    layer3_outputs(11431) <= b;
    layer3_outputs(11432) <= '1';
    layer3_outputs(11433) <= '0';
    layer3_outputs(11434) <= not b;
    layer3_outputs(11435) <= a and not b;
    layer3_outputs(11436) <= not b or a;
    layer3_outputs(11437) <= not b;
    layer3_outputs(11438) <= '1';
    layer3_outputs(11439) <= not b;
    layer3_outputs(11440) <= not a or b;
    layer3_outputs(11441) <= not b;
    layer3_outputs(11442) <= not (a and b);
    layer3_outputs(11443) <= not b;
    layer3_outputs(11444) <= b and not a;
    layer3_outputs(11445) <= a xor b;
    layer3_outputs(11446) <= not a;
    layer3_outputs(11447) <= not (a xor b);
    layer3_outputs(11448) <= not a or b;
    layer3_outputs(11449) <= not b;
    layer3_outputs(11450) <= a and not b;
    layer3_outputs(11451) <= b and not a;
    layer3_outputs(11452) <= '1';
    layer3_outputs(11453) <= a or b;
    layer3_outputs(11454) <= a;
    layer3_outputs(11455) <= '0';
    layer3_outputs(11456) <= a and b;
    layer3_outputs(11457) <= a xor b;
    layer3_outputs(11458) <= not (a and b);
    layer3_outputs(11459) <= not (a or b);
    layer3_outputs(11460) <= not (a and b);
    layer3_outputs(11461) <= b and not a;
    layer3_outputs(11462) <= a or b;
    layer3_outputs(11463) <= not b or a;
    layer3_outputs(11464) <= a;
    layer3_outputs(11465) <= '1';
    layer3_outputs(11466) <= a;
    layer3_outputs(11467) <= not a;
    layer3_outputs(11468) <= not b or a;
    layer3_outputs(11469) <= a;
    layer3_outputs(11470) <= not (a and b);
    layer3_outputs(11471) <= a and not b;
    layer3_outputs(11472) <= a and not b;
    layer3_outputs(11473) <= not (a or b);
    layer3_outputs(11474) <= a;
    layer3_outputs(11475) <= a;
    layer3_outputs(11476) <= b;
    layer3_outputs(11477) <= not b;
    layer3_outputs(11478) <= not a;
    layer3_outputs(11479) <= not a or b;
    layer3_outputs(11480) <= a;
    layer3_outputs(11481) <= not a or b;
    layer3_outputs(11482) <= not (a and b);
    layer3_outputs(11483) <= not a or b;
    layer3_outputs(11484) <= a or b;
    layer3_outputs(11485) <= not a;
    layer3_outputs(11486) <= not a;
    layer3_outputs(11487) <= not b;
    layer3_outputs(11488) <= b and not a;
    layer3_outputs(11489) <= not b;
    layer3_outputs(11490) <= '1';
    layer3_outputs(11491) <= not b or a;
    layer3_outputs(11492) <= not (a or b);
    layer3_outputs(11493) <= a;
    layer3_outputs(11494) <= not (a or b);
    layer3_outputs(11495) <= not b;
    layer3_outputs(11496) <= not a;
    layer3_outputs(11497) <= not a or b;
    layer3_outputs(11498) <= b;
    layer3_outputs(11499) <= a;
    layer3_outputs(11500) <= not a or b;
    layer3_outputs(11501) <= a and not b;
    layer3_outputs(11502) <= not b;
    layer3_outputs(11503) <= b and not a;
    layer3_outputs(11504) <= a;
    layer3_outputs(11505) <= not b;
    layer3_outputs(11506) <= not a or b;
    layer3_outputs(11507) <= a;
    layer3_outputs(11508) <= a;
    layer3_outputs(11509) <= not a;
    layer3_outputs(11510) <= '1';
    layer3_outputs(11511) <= b;
    layer3_outputs(11512) <= not (a and b);
    layer3_outputs(11513) <= not a;
    layer3_outputs(11514) <= not b;
    layer3_outputs(11515) <= not (a or b);
    layer3_outputs(11516) <= not (a and b);
    layer3_outputs(11517) <= a;
    layer3_outputs(11518) <= b;
    layer3_outputs(11519) <= not (a or b);
    layer3_outputs(11520) <= '0';
    layer3_outputs(11521) <= not a;
    layer3_outputs(11522) <= not a or b;
    layer3_outputs(11523) <= a and b;
    layer3_outputs(11524) <= b;
    layer3_outputs(11525) <= b;
    layer3_outputs(11526) <= not (a and b);
    layer3_outputs(11527) <= a;
    layer3_outputs(11528) <= a;
    layer3_outputs(11529) <= b;
    layer3_outputs(11530) <= not b;
    layer3_outputs(11531) <= b and not a;
    layer3_outputs(11532) <= a;
    layer3_outputs(11533) <= '0';
    layer3_outputs(11534) <= not a or b;
    layer3_outputs(11535) <= not (a and b);
    layer3_outputs(11536) <= a and not b;
    layer3_outputs(11537) <= a xor b;
    layer3_outputs(11538) <= not (a or b);
    layer3_outputs(11539) <= b and not a;
    layer3_outputs(11540) <= not (a or b);
    layer3_outputs(11541) <= a;
    layer3_outputs(11542) <= not a;
    layer3_outputs(11543) <= a;
    layer3_outputs(11544) <= '0';
    layer3_outputs(11545) <= '1';
    layer3_outputs(11546) <= not a;
    layer3_outputs(11547) <= a and not b;
    layer3_outputs(11548) <= not (a xor b);
    layer3_outputs(11549) <= b;
    layer3_outputs(11550) <= not a;
    layer3_outputs(11551) <= b and not a;
    layer3_outputs(11552) <= not b;
    layer3_outputs(11553) <= not b;
    layer3_outputs(11554) <= not a;
    layer3_outputs(11555) <= b and not a;
    layer3_outputs(11556) <= a and not b;
    layer3_outputs(11557) <= a xor b;
    layer3_outputs(11558) <= b;
    layer3_outputs(11559) <= not (a and b);
    layer3_outputs(11560) <= not (a xor b);
    layer3_outputs(11561) <= not b;
    layer3_outputs(11562) <= not (a xor b);
    layer3_outputs(11563) <= not (a or b);
    layer3_outputs(11564) <= a and b;
    layer3_outputs(11565) <= not a or b;
    layer3_outputs(11566) <= not b;
    layer3_outputs(11567) <= not (a or b);
    layer3_outputs(11568) <= not b or a;
    layer3_outputs(11569) <= '1';
    layer3_outputs(11570) <= not a or b;
    layer3_outputs(11571) <= b;
    layer3_outputs(11572) <= not b or a;
    layer3_outputs(11573) <= not b or a;
    layer3_outputs(11574) <= b;
    layer3_outputs(11575) <= a;
    layer3_outputs(11576) <= not b;
    layer3_outputs(11577) <= not b;
    layer3_outputs(11578) <= a and b;
    layer3_outputs(11579) <= b;
    layer3_outputs(11580) <= a or b;
    layer3_outputs(11581) <= '1';
    layer3_outputs(11582) <= a and not b;
    layer3_outputs(11583) <= not (a and b);
    layer3_outputs(11584) <= not (a or b);
    layer3_outputs(11585) <= not a;
    layer3_outputs(11586) <= not b;
    layer3_outputs(11587) <= not a;
    layer3_outputs(11588) <= not (a or b);
    layer3_outputs(11589) <= not b or a;
    layer3_outputs(11590) <= b;
    layer3_outputs(11591) <= not a;
    layer3_outputs(11592) <= not (a and b);
    layer3_outputs(11593) <= not (a and b);
    layer3_outputs(11594) <= not (a or b);
    layer3_outputs(11595) <= not b;
    layer3_outputs(11596) <= b;
    layer3_outputs(11597) <= b;
    layer3_outputs(11598) <= not a or b;
    layer3_outputs(11599) <= not a;
    layer3_outputs(11600) <= '0';
    layer3_outputs(11601) <= not b or a;
    layer3_outputs(11602) <= not (a or b);
    layer3_outputs(11603) <= b and not a;
    layer3_outputs(11604) <= not (a xor b);
    layer3_outputs(11605) <= '0';
    layer3_outputs(11606) <= '1';
    layer3_outputs(11607) <= not a;
    layer3_outputs(11608) <= not (a xor b);
    layer3_outputs(11609) <= a;
    layer3_outputs(11610) <= a or b;
    layer3_outputs(11611) <= not (a or b);
    layer3_outputs(11612) <= not a or b;
    layer3_outputs(11613) <= a or b;
    layer3_outputs(11614) <= not a or b;
    layer3_outputs(11615) <= not a or b;
    layer3_outputs(11616) <= not a;
    layer3_outputs(11617) <= a;
    layer3_outputs(11618) <= not b or a;
    layer3_outputs(11619) <= a or b;
    layer3_outputs(11620) <= a and not b;
    layer3_outputs(11621) <= b;
    layer3_outputs(11622) <= not b or a;
    layer3_outputs(11623) <= not b;
    layer3_outputs(11624) <= not a or b;
    layer3_outputs(11625) <= b and not a;
    layer3_outputs(11626) <= a;
    layer3_outputs(11627) <= a or b;
    layer3_outputs(11628) <= a and b;
    layer3_outputs(11629) <= not a or b;
    layer3_outputs(11630) <= b;
    layer3_outputs(11631) <= not (a and b);
    layer3_outputs(11632) <= not b;
    layer3_outputs(11633) <= not b;
    layer3_outputs(11634) <= not (a xor b);
    layer3_outputs(11635) <= a and b;
    layer3_outputs(11636) <= not a;
    layer3_outputs(11637) <= not a;
    layer3_outputs(11638) <= a;
    layer3_outputs(11639) <= b;
    layer3_outputs(11640) <= a or b;
    layer3_outputs(11641) <= a;
    layer3_outputs(11642) <= not b;
    layer3_outputs(11643) <= a xor b;
    layer3_outputs(11644) <= not a or b;
    layer3_outputs(11645) <= not a or b;
    layer3_outputs(11646) <= b and not a;
    layer3_outputs(11647) <= b;
    layer3_outputs(11648) <= a;
    layer3_outputs(11649) <= b and not a;
    layer3_outputs(11650) <= not a;
    layer3_outputs(11651) <= b and not a;
    layer3_outputs(11652) <= a and not b;
    layer3_outputs(11653) <= not (a xor b);
    layer3_outputs(11654) <= b and not a;
    layer3_outputs(11655) <= a;
    layer3_outputs(11656) <= not b;
    layer3_outputs(11657) <= not a;
    layer3_outputs(11658) <= a xor b;
    layer3_outputs(11659) <= b;
    layer3_outputs(11660) <= '0';
    layer3_outputs(11661) <= b and not a;
    layer3_outputs(11662) <= b and not a;
    layer3_outputs(11663) <= not (a or b);
    layer3_outputs(11664) <= a xor b;
    layer3_outputs(11665) <= a and not b;
    layer3_outputs(11666) <= a xor b;
    layer3_outputs(11667) <= not (a xor b);
    layer3_outputs(11668) <= not a or b;
    layer3_outputs(11669) <= a or b;
    layer3_outputs(11670) <= b and not a;
    layer3_outputs(11671) <= not (a xor b);
    layer3_outputs(11672) <= not b;
    layer3_outputs(11673) <= '1';
    layer3_outputs(11674) <= not b or a;
    layer3_outputs(11675) <= a and not b;
    layer3_outputs(11676) <= a;
    layer3_outputs(11677) <= a and not b;
    layer3_outputs(11678) <= not (a xor b);
    layer3_outputs(11679) <= a;
    layer3_outputs(11680) <= not a;
    layer3_outputs(11681) <= not b;
    layer3_outputs(11682) <= not a;
    layer3_outputs(11683) <= b;
    layer3_outputs(11684) <= not b;
    layer3_outputs(11685) <= not a;
    layer3_outputs(11686) <= a or b;
    layer3_outputs(11687) <= not b;
    layer3_outputs(11688) <= a and not b;
    layer3_outputs(11689) <= '1';
    layer3_outputs(11690) <= not b or a;
    layer3_outputs(11691) <= a;
    layer3_outputs(11692) <= a and not b;
    layer3_outputs(11693) <= b;
    layer3_outputs(11694) <= a xor b;
    layer3_outputs(11695) <= '1';
    layer3_outputs(11696) <= not b;
    layer3_outputs(11697) <= not a;
    layer3_outputs(11698) <= not b or a;
    layer3_outputs(11699) <= not a or b;
    layer3_outputs(11700) <= not b;
    layer3_outputs(11701) <= a xor b;
    layer3_outputs(11702) <= not b;
    layer3_outputs(11703) <= b and not a;
    layer3_outputs(11704) <= not b or a;
    layer3_outputs(11705) <= not a or b;
    layer3_outputs(11706) <= not (a and b);
    layer3_outputs(11707) <= not (a and b);
    layer3_outputs(11708) <= not b;
    layer3_outputs(11709) <= not a;
    layer3_outputs(11710) <= a or b;
    layer3_outputs(11711) <= not a or b;
    layer3_outputs(11712) <= not (a and b);
    layer3_outputs(11713) <= not a;
    layer3_outputs(11714) <= a;
    layer3_outputs(11715) <= not b;
    layer3_outputs(11716) <= not b;
    layer3_outputs(11717) <= a;
    layer3_outputs(11718) <= '1';
    layer3_outputs(11719) <= not (a or b);
    layer3_outputs(11720) <= '0';
    layer3_outputs(11721) <= not a or b;
    layer3_outputs(11722) <= a and b;
    layer3_outputs(11723) <= not a or b;
    layer3_outputs(11724) <= a and not b;
    layer3_outputs(11725) <= b and not a;
    layer3_outputs(11726) <= not a or b;
    layer3_outputs(11727) <= b and not a;
    layer3_outputs(11728) <= not (a and b);
    layer3_outputs(11729) <= not a or b;
    layer3_outputs(11730) <= a or b;
    layer3_outputs(11731) <= a and b;
    layer3_outputs(11732) <= '1';
    layer3_outputs(11733) <= not a or b;
    layer3_outputs(11734) <= not a or b;
    layer3_outputs(11735) <= not a or b;
    layer3_outputs(11736) <= a;
    layer3_outputs(11737) <= not (a and b);
    layer3_outputs(11738) <= a and not b;
    layer3_outputs(11739) <= a or b;
    layer3_outputs(11740) <= not a;
    layer3_outputs(11741) <= b and not a;
    layer3_outputs(11742) <= not (a and b);
    layer3_outputs(11743) <= a and b;
    layer3_outputs(11744) <= b;
    layer3_outputs(11745) <= a;
    layer3_outputs(11746) <= b and not a;
    layer3_outputs(11747) <= a;
    layer3_outputs(11748) <= a or b;
    layer3_outputs(11749) <= a;
    layer3_outputs(11750) <= a;
    layer3_outputs(11751) <= '0';
    layer3_outputs(11752) <= not a;
    layer3_outputs(11753) <= not a;
    layer3_outputs(11754) <= a and not b;
    layer3_outputs(11755) <= '0';
    layer3_outputs(11756) <= not a or b;
    layer3_outputs(11757) <= not (a and b);
    layer3_outputs(11758) <= a xor b;
    layer3_outputs(11759) <= '0';
    layer3_outputs(11760) <= not a;
    layer3_outputs(11761) <= a and not b;
    layer3_outputs(11762) <= b and not a;
    layer3_outputs(11763) <= not (a and b);
    layer3_outputs(11764) <= not b;
    layer3_outputs(11765) <= a and not b;
    layer3_outputs(11766) <= '1';
    layer3_outputs(11767) <= not (a xor b);
    layer3_outputs(11768) <= not b;
    layer3_outputs(11769) <= b;
    layer3_outputs(11770) <= '1';
    layer3_outputs(11771) <= a;
    layer3_outputs(11772) <= not b or a;
    layer3_outputs(11773) <= not (a or b);
    layer3_outputs(11774) <= not (a and b);
    layer3_outputs(11775) <= a or b;
    layer3_outputs(11776) <= not b or a;
    layer3_outputs(11777) <= b and not a;
    layer3_outputs(11778) <= not a;
    layer3_outputs(11779) <= not b or a;
    layer3_outputs(11780) <= b;
    layer3_outputs(11781) <= not b or a;
    layer3_outputs(11782) <= a and not b;
    layer3_outputs(11783) <= b and not a;
    layer3_outputs(11784) <= '1';
    layer3_outputs(11785) <= a;
    layer3_outputs(11786) <= not b or a;
    layer3_outputs(11787) <= not (a or b);
    layer3_outputs(11788) <= a or b;
    layer3_outputs(11789) <= a or b;
    layer3_outputs(11790) <= not b or a;
    layer3_outputs(11791) <= b;
    layer3_outputs(11792) <= b and not a;
    layer3_outputs(11793) <= not a or b;
    layer3_outputs(11794) <= not a;
    layer3_outputs(11795) <= b;
    layer3_outputs(11796) <= a xor b;
    layer3_outputs(11797) <= '0';
    layer3_outputs(11798) <= '0';
    layer3_outputs(11799) <= a;
    layer3_outputs(11800) <= a;
    layer3_outputs(11801) <= b;
    layer3_outputs(11802) <= a;
    layer3_outputs(11803) <= a and b;
    layer3_outputs(11804) <= a and b;
    layer3_outputs(11805) <= not b;
    layer3_outputs(11806) <= not a or b;
    layer3_outputs(11807) <= a xor b;
    layer3_outputs(11808) <= b;
    layer3_outputs(11809) <= b;
    layer3_outputs(11810) <= not a;
    layer3_outputs(11811) <= not (a or b);
    layer3_outputs(11812) <= '0';
    layer3_outputs(11813) <= not a or b;
    layer3_outputs(11814) <= not b or a;
    layer3_outputs(11815) <= a;
    layer3_outputs(11816) <= b and not a;
    layer3_outputs(11817) <= a and not b;
    layer3_outputs(11818) <= not (a or b);
    layer3_outputs(11819) <= not (a and b);
    layer3_outputs(11820) <= b and not a;
    layer3_outputs(11821) <= not (a or b);
    layer3_outputs(11822) <= not (a and b);
    layer3_outputs(11823) <= not (a and b);
    layer3_outputs(11824) <= not (a or b);
    layer3_outputs(11825) <= '0';
    layer3_outputs(11826) <= a and b;
    layer3_outputs(11827) <= a or b;
    layer3_outputs(11828) <= b;
    layer3_outputs(11829) <= not b or a;
    layer3_outputs(11830) <= not b or a;
    layer3_outputs(11831) <= not a or b;
    layer3_outputs(11832) <= not (a or b);
    layer3_outputs(11833) <= a or b;
    layer3_outputs(11834) <= '0';
    layer3_outputs(11835) <= b;
    layer3_outputs(11836) <= not (a xor b);
    layer3_outputs(11837) <= b;
    layer3_outputs(11838) <= a;
    layer3_outputs(11839) <= not b;
    layer3_outputs(11840) <= not b or a;
    layer3_outputs(11841) <= a and b;
    layer3_outputs(11842) <= not (a or b);
    layer3_outputs(11843) <= a and not b;
    layer3_outputs(11844) <= not (a xor b);
    layer3_outputs(11845) <= not b or a;
    layer3_outputs(11846) <= a or b;
    layer3_outputs(11847) <= a and b;
    layer3_outputs(11848) <= not a or b;
    layer3_outputs(11849) <= a and b;
    layer3_outputs(11850) <= b;
    layer3_outputs(11851) <= b;
    layer3_outputs(11852) <= a;
    layer3_outputs(11853) <= not a or b;
    layer3_outputs(11854) <= '1';
    layer3_outputs(11855) <= b and not a;
    layer3_outputs(11856) <= not b or a;
    layer3_outputs(11857) <= b;
    layer3_outputs(11858) <= not (a or b);
    layer3_outputs(11859) <= not (a and b);
    layer3_outputs(11860) <= a or b;
    layer3_outputs(11861) <= a;
    layer3_outputs(11862) <= a;
    layer3_outputs(11863) <= a;
    layer3_outputs(11864) <= not a;
    layer3_outputs(11865) <= not (a and b);
    layer3_outputs(11866) <= not (a or b);
    layer3_outputs(11867) <= '1';
    layer3_outputs(11868) <= not b;
    layer3_outputs(11869) <= b and not a;
    layer3_outputs(11870) <= not a;
    layer3_outputs(11871) <= b and not a;
    layer3_outputs(11872) <= not (a xor b);
    layer3_outputs(11873) <= not a;
    layer3_outputs(11874) <= not b;
    layer3_outputs(11875) <= not b;
    layer3_outputs(11876) <= a or b;
    layer3_outputs(11877) <= a;
    layer3_outputs(11878) <= not b;
    layer3_outputs(11879) <= not (a or b);
    layer3_outputs(11880) <= not b;
    layer3_outputs(11881) <= a or b;
    layer3_outputs(11882) <= not b;
    layer3_outputs(11883) <= not b;
    layer3_outputs(11884) <= a xor b;
    layer3_outputs(11885) <= b;
    layer3_outputs(11886) <= not b or a;
    layer3_outputs(11887) <= a;
    layer3_outputs(11888) <= a and b;
    layer3_outputs(11889) <= not (a xor b);
    layer3_outputs(11890) <= not (a or b);
    layer3_outputs(11891) <= not (a xor b);
    layer3_outputs(11892) <= a and b;
    layer3_outputs(11893) <= not b;
    layer3_outputs(11894) <= b and not a;
    layer3_outputs(11895) <= a and b;
    layer3_outputs(11896) <= a xor b;
    layer3_outputs(11897) <= not (a or b);
    layer3_outputs(11898) <= not (a xor b);
    layer3_outputs(11899) <= not (a xor b);
    layer3_outputs(11900) <= a;
    layer3_outputs(11901) <= not b;
    layer3_outputs(11902) <= not (a xor b);
    layer3_outputs(11903) <= b and not a;
    layer3_outputs(11904) <= not a or b;
    layer3_outputs(11905) <= not a;
    layer3_outputs(11906) <= a or b;
    layer3_outputs(11907) <= a;
    layer3_outputs(11908) <= b;
    layer3_outputs(11909) <= not b;
    layer3_outputs(11910) <= not (a or b);
    layer3_outputs(11911) <= b;
    layer3_outputs(11912) <= not (a or b);
    layer3_outputs(11913) <= not (a xor b);
    layer3_outputs(11914) <= not b;
    layer3_outputs(11915) <= a and not b;
    layer3_outputs(11916) <= not a or b;
    layer3_outputs(11917) <= not a or b;
    layer3_outputs(11918) <= a;
    layer3_outputs(11919) <= a or b;
    layer3_outputs(11920) <= not (a xor b);
    layer3_outputs(11921) <= a xor b;
    layer3_outputs(11922) <= not a or b;
    layer3_outputs(11923) <= not b;
    layer3_outputs(11924) <= not b or a;
    layer3_outputs(11925) <= not a;
    layer3_outputs(11926) <= not a;
    layer3_outputs(11927) <= not b or a;
    layer3_outputs(11928) <= b;
    layer3_outputs(11929) <= not b;
    layer3_outputs(11930) <= not b;
    layer3_outputs(11931) <= a or b;
    layer3_outputs(11932) <= not b;
    layer3_outputs(11933) <= '0';
    layer3_outputs(11934) <= not a;
    layer3_outputs(11935) <= b;
    layer3_outputs(11936) <= not b;
    layer3_outputs(11937) <= b;
    layer3_outputs(11938) <= not a;
    layer3_outputs(11939) <= b;
    layer3_outputs(11940) <= a;
    layer3_outputs(11941) <= '1';
    layer3_outputs(11942) <= not b or a;
    layer3_outputs(11943) <= '0';
    layer3_outputs(11944) <= a and not b;
    layer3_outputs(11945) <= a and b;
    layer3_outputs(11946) <= b;
    layer3_outputs(11947) <= a and not b;
    layer3_outputs(11948) <= a;
    layer3_outputs(11949) <= not a;
    layer3_outputs(11950) <= not (a xor b);
    layer3_outputs(11951) <= not a;
    layer3_outputs(11952) <= not b or a;
    layer3_outputs(11953) <= a and b;
    layer3_outputs(11954) <= b;
    layer3_outputs(11955) <= not a;
    layer3_outputs(11956) <= a or b;
    layer3_outputs(11957) <= not b or a;
    layer3_outputs(11958) <= a;
    layer3_outputs(11959) <= not a or b;
    layer3_outputs(11960) <= a;
    layer3_outputs(11961) <= not b;
    layer3_outputs(11962) <= not a;
    layer3_outputs(11963) <= '1';
    layer3_outputs(11964) <= not a or b;
    layer3_outputs(11965) <= b and not a;
    layer3_outputs(11966) <= '1';
    layer3_outputs(11967) <= not a;
    layer3_outputs(11968) <= not b or a;
    layer3_outputs(11969) <= '1';
    layer3_outputs(11970) <= not b;
    layer3_outputs(11971) <= not a;
    layer3_outputs(11972) <= not a;
    layer3_outputs(11973) <= not b;
    layer3_outputs(11974) <= '0';
    layer3_outputs(11975) <= b and not a;
    layer3_outputs(11976) <= a or b;
    layer3_outputs(11977) <= not (a xor b);
    layer3_outputs(11978) <= not (a or b);
    layer3_outputs(11979) <= a xor b;
    layer3_outputs(11980) <= b;
    layer3_outputs(11981) <= not b;
    layer3_outputs(11982) <= b;
    layer3_outputs(11983) <= b;
    layer3_outputs(11984) <= '1';
    layer3_outputs(11985) <= a;
    layer3_outputs(11986) <= not b;
    layer3_outputs(11987) <= not b or a;
    layer3_outputs(11988) <= not (a and b);
    layer3_outputs(11989) <= a xor b;
    layer3_outputs(11990) <= a and not b;
    layer3_outputs(11991) <= a xor b;
    layer3_outputs(11992) <= not b;
    layer3_outputs(11993) <= not (a and b);
    layer3_outputs(11994) <= not a;
    layer3_outputs(11995) <= a;
    layer3_outputs(11996) <= not (a xor b);
    layer3_outputs(11997) <= a xor b;
    layer3_outputs(11998) <= '1';
    layer3_outputs(11999) <= a and not b;
    layer3_outputs(12000) <= not (a and b);
    layer3_outputs(12001) <= not b or a;
    layer3_outputs(12002) <= b;
    layer3_outputs(12003) <= b;
    layer3_outputs(12004) <= '1';
    layer3_outputs(12005) <= a;
    layer3_outputs(12006) <= not (a xor b);
    layer3_outputs(12007) <= a or b;
    layer3_outputs(12008) <= a and b;
    layer3_outputs(12009) <= a and not b;
    layer3_outputs(12010) <= not (a or b);
    layer3_outputs(12011) <= '0';
    layer3_outputs(12012) <= not b or a;
    layer3_outputs(12013) <= not (a or b);
    layer3_outputs(12014) <= not b;
    layer3_outputs(12015) <= '0';
    layer3_outputs(12016) <= b;
    layer3_outputs(12017) <= a;
    layer3_outputs(12018) <= b;
    layer3_outputs(12019) <= not (a xor b);
    layer3_outputs(12020) <= b;
    layer3_outputs(12021) <= a;
    layer3_outputs(12022) <= not a or b;
    layer3_outputs(12023) <= a xor b;
    layer3_outputs(12024) <= not b or a;
    layer3_outputs(12025) <= a xor b;
    layer3_outputs(12026) <= a and b;
    layer3_outputs(12027) <= not b or a;
    layer3_outputs(12028) <= not b or a;
    layer3_outputs(12029) <= not a;
    layer3_outputs(12030) <= a;
    layer3_outputs(12031) <= a and not b;
    layer3_outputs(12032) <= not a or b;
    layer3_outputs(12033) <= not (a or b);
    layer3_outputs(12034) <= not b;
    layer3_outputs(12035) <= not b or a;
    layer3_outputs(12036) <= a and not b;
    layer3_outputs(12037) <= not a;
    layer3_outputs(12038) <= not a or b;
    layer3_outputs(12039) <= not b;
    layer3_outputs(12040) <= b and not a;
    layer3_outputs(12041) <= not a;
    layer3_outputs(12042) <= a;
    layer3_outputs(12043) <= not b or a;
    layer3_outputs(12044) <= a and b;
    layer3_outputs(12045) <= not b;
    layer3_outputs(12046) <= a;
    layer3_outputs(12047) <= b and not a;
    layer3_outputs(12048) <= '0';
    layer3_outputs(12049) <= a;
    layer3_outputs(12050) <= a;
    layer3_outputs(12051) <= '0';
    layer3_outputs(12052) <= not b or a;
    layer3_outputs(12053) <= b and not a;
    layer3_outputs(12054) <= a and not b;
    layer3_outputs(12055) <= a;
    layer3_outputs(12056) <= a;
    layer3_outputs(12057) <= not a;
    layer3_outputs(12058) <= not a;
    layer3_outputs(12059) <= a;
    layer3_outputs(12060) <= b and not a;
    layer3_outputs(12061) <= a;
    layer3_outputs(12062) <= not b or a;
    layer3_outputs(12063) <= not (a or b);
    layer3_outputs(12064) <= not (a or b);
    layer3_outputs(12065) <= not (a or b);
    layer3_outputs(12066) <= b and not a;
    layer3_outputs(12067) <= a;
    layer3_outputs(12068) <= a and b;
    layer3_outputs(12069) <= not (a or b);
    layer3_outputs(12070) <= not a or b;
    layer3_outputs(12071) <= not b;
    layer3_outputs(12072) <= not a;
    layer3_outputs(12073) <= b and not a;
    layer3_outputs(12074) <= a or b;
    layer3_outputs(12075) <= '0';
    layer3_outputs(12076) <= not b or a;
    layer3_outputs(12077) <= not (a xor b);
    layer3_outputs(12078) <= a xor b;
    layer3_outputs(12079) <= a;
    layer3_outputs(12080) <= a and not b;
    layer3_outputs(12081) <= '0';
    layer3_outputs(12082) <= not (a or b);
    layer3_outputs(12083) <= not b or a;
    layer3_outputs(12084) <= a and not b;
    layer3_outputs(12085) <= a xor b;
    layer3_outputs(12086) <= a;
    layer3_outputs(12087) <= b and not a;
    layer3_outputs(12088) <= '0';
    layer3_outputs(12089) <= not (a or b);
    layer3_outputs(12090) <= a or b;
    layer3_outputs(12091) <= not a or b;
    layer3_outputs(12092) <= b;
    layer3_outputs(12093) <= not b or a;
    layer3_outputs(12094) <= a;
    layer3_outputs(12095) <= not a;
    layer3_outputs(12096) <= a xor b;
    layer3_outputs(12097) <= not a;
    layer3_outputs(12098) <= a;
    layer3_outputs(12099) <= b;
    layer3_outputs(12100) <= a and b;
    layer3_outputs(12101) <= not a;
    layer3_outputs(12102) <= not a;
    layer3_outputs(12103) <= a;
    layer3_outputs(12104) <= b and not a;
    layer3_outputs(12105) <= a and not b;
    layer3_outputs(12106) <= a;
    layer3_outputs(12107) <= not a;
    layer3_outputs(12108) <= b;
    layer3_outputs(12109) <= not a;
    layer3_outputs(12110) <= '1';
    layer3_outputs(12111) <= b and not a;
    layer3_outputs(12112) <= b and not a;
    layer3_outputs(12113) <= a;
    layer3_outputs(12114) <= not (a or b);
    layer3_outputs(12115) <= not b or a;
    layer3_outputs(12116) <= b;
    layer3_outputs(12117) <= not a;
    layer3_outputs(12118) <= a and b;
    layer3_outputs(12119) <= b;
    layer3_outputs(12120) <= '0';
    layer3_outputs(12121) <= not b or a;
    layer3_outputs(12122) <= not a;
    layer3_outputs(12123) <= a and b;
    layer3_outputs(12124) <= a;
    layer3_outputs(12125) <= not b;
    layer3_outputs(12126) <= b;
    layer3_outputs(12127) <= not (a and b);
    layer3_outputs(12128) <= not (a and b);
    layer3_outputs(12129) <= not a;
    layer3_outputs(12130) <= a or b;
    layer3_outputs(12131) <= a and not b;
    layer3_outputs(12132) <= a;
    layer3_outputs(12133) <= b and not a;
    layer3_outputs(12134) <= not (a or b);
    layer3_outputs(12135) <= a and not b;
    layer3_outputs(12136) <= '1';
    layer3_outputs(12137) <= b and not a;
    layer3_outputs(12138) <= '0';
    layer3_outputs(12139) <= not b;
    layer3_outputs(12140) <= a and b;
    layer3_outputs(12141) <= not a;
    layer3_outputs(12142) <= b and not a;
    layer3_outputs(12143) <= not (a and b);
    layer3_outputs(12144) <= not b or a;
    layer3_outputs(12145) <= not b or a;
    layer3_outputs(12146) <= not (a or b);
    layer3_outputs(12147) <= not b;
    layer3_outputs(12148) <= not a or b;
    layer3_outputs(12149) <= not b or a;
    layer3_outputs(12150) <= a and b;
    layer3_outputs(12151) <= not b or a;
    layer3_outputs(12152) <= a;
    layer3_outputs(12153) <= a xor b;
    layer3_outputs(12154) <= a and not b;
    layer3_outputs(12155) <= a and b;
    layer3_outputs(12156) <= b;
    layer3_outputs(12157) <= a;
    layer3_outputs(12158) <= not a;
    layer3_outputs(12159) <= not a;
    layer3_outputs(12160) <= not (a or b);
    layer3_outputs(12161) <= a xor b;
    layer3_outputs(12162) <= not b or a;
    layer3_outputs(12163) <= '0';
    layer3_outputs(12164) <= '1';
    layer3_outputs(12165) <= not b or a;
    layer3_outputs(12166) <= not b or a;
    layer3_outputs(12167) <= not (a or b);
    layer3_outputs(12168) <= b;
    layer3_outputs(12169) <= b;
    layer3_outputs(12170) <= b;
    layer3_outputs(12171) <= b;
    layer3_outputs(12172) <= '0';
    layer3_outputs(12173) <= a or b;
    layer3_outputs(12174) <= not b or a;
    layer3_outputs(12175) <= not (a xor b);
    layer3_outputs(12176) <= b and not a;
    layer3_outputs(12177) <= b;
    layer3_outputs(12178) <= a xor b;
    layer3_outputs(12179) <= not b;
    layer3_outputs(12180) <= not a or b;
    layer3_outputs(12181) <= not a or b;
    layer3_outputs(12182) <= not a or b;
    layer3_outputs(12183) <= not a;
    layer3_outputs(12184) <= a and not b;
    layer3_outputs(12185) <= not (a and b);
    layer3_outputs(12186) <= not a;
    layer3_outputs(12187) <= a;
    layer3_outputs(12188) <= not (a or b);
    layer3_outputs(12189) <= not b or a;
    layer3_outputs(12190) <= a;
    layer3_outputs(12191) <= b;
    layer3_outputs(12192) <= a;
    layer3_outputs(12193) <= not (a and b);
    layer3_outputs(12194) <= not a or b;
    layer3_outputs(12195) <= not a;
    layer3_outputs(12196) <= not a or b;
    layer3_outputs(12197) <= not b;
    layer3_outputs(12198) <= not (a xor b);
    layer3_outputs(12199) <= a and not b;
    layer3_outputs(12200) <= not a or b;
    layer3_outputs(12201) <= not (a and b);
    layer3_outputs(12202) <= not (a xor b);
    layer3_outputs(12203) <= not (a and b);
    layer3_outputs(12204) <= '1';
    layer3_outputs(12205) <= '0';
    layer3_outputs(12206) <= not a or b;
    layer3_outputs(12207) <= a or b;
    layer3_outputs(12208) <= b;
    layer3_outputs(12209) <= not b;
    layer3_outputs(12210) <= not b;
    layer3_outputs(12211) <= a and b;
    layer3_outputs(12212) <= not b or a;
    layer3_outputs(12213) <= not (a and b);
    layer3_outputs(12214) <= not a or b;
    layer3_outputs(12215) <= b and not a;
    layer3_outputs(12216) <= not (a xor b);
    layer3_outputs(12217) <= a and b;
    layer3_outputs(12218) <= a and b;
    layer3_outputs(12219) <= a or b;
    layer3_outputs(12220) <= b;
    layer3_outputs(12221) <= not (a xor b);
    layer3_outputs(12222) <= not a;
    layer3_outputs(12223) <= '1';
    layer3_outputs(12224) <= not (a and b);
    layer3_outputs(12225) <= b;
    layer3_outputs(12226) <= b and not a;
    layer3_outputs(12227) <= not a;
    layer3_outputs(12228) <= a or b;
    layer3_outputs(12229) <= a or b;
    layer3_outputs(12230) <= a xor b;
    layer3_outputs(12231) <= b;
    layer3_outputs(12232) <= not (a or b);
    layer3_outputs(12233) <= b;
    layer3_outputs(12234) <= not a;
    layer3_outputs(12235) <= not (a xor b);
    layer3_outputs(12236) <= not (a or b);
    layer3_outputs(12237) <= not b or a;
    layer3_outputs(12238) <= not b;
    layer3_outputs(12239) <= '0';
    layer3_outputs(12240) <= not b or a;
    layer3_outputs(12241) <= not (a and b);
    layer3_outputs(12242) <= b;
    layer3_outputs(12243) <= not a;
    layer3_outputs(12244) <= a xor b;
    layer3_outputs(12245) <= '1';
    layer3_outputs(12246) <= b;
    layer3_outputs(12247) <= a xor b;
    layer3_outputs(12248) <= b;
    layer3_outputs(12249) <= not a;
    layer3_outputs(12250) <= not a or b;
    layer3_outputs(12251) <= not b;
    layer3_outputs(12252) <= not a or b;
    layer3_outputs(12253) <= not b or a;
    layer3_outputs(12254) <= not b;
    layer3_outputs(12255) <= b;
    layer3_outputs(12256) <= a or b;
    layer3_outputs(12257) <= a;
    layer3_outputs(12258) <= not a or b;
    layer3_outputs(12259) <= a or b;
    layer3_outputs(12260) <= not b;
    layer3_outputs(12261) <= b and not a;
    layer3_outputs(12262) <= a and b;
    layer3_outputs(12263) <= not (a and b);
    layer3_outputs(12264) <= a and b;
    layer3_outputs(12265) <= not (a xor b);
    layer3_outputs(12266) <= not (a or b);
    layer3_outputs(12267) <= a xor b;
    layer3_outputs(12268) <= not (a or b);
    layer3_outputs(12269) <= a;
    layer3_outputs(12270) <= a;
    layer3_outputs(12271) <= not (a xor b);
    layer3_outputs(12272) <= not (a xor b);
    layer3_outputs(12273) <= a and b;
    layer3_outputs(12274) <= not a or b;
    layer3_outputs(12275) <= not a;
    layer3_outputs(12276) <= not b;
    layer3_outputs(12277) <= a;
    layer3_outputs(12278) <= '1';
    layer3_outputs(12279) <= not (a and b);
    layer3_outputs(12280) <= a;
    layer3_outputs(12281) <= b;
    layer3_outputs(12282) <= a and b;
    layer3_outputs(12283) <= not (a or b);
    layer3_outputs(12284) <= not (a xor b);
    layer3_outputs(12285) <= not a or b;
    layer3_outputs(12286) <= b;
    layer3_outputs(12287) <= not (a or b);
    layer3_outputs(12288) <= not (a xor b);
    layer3_outputs(12289) <= not b;
    layer3_outputs(12290) <= not (a and b);
    layer3_outputs(12291) <= b;
    layer3_outputs(12292) <= a;
    layer3_outputs(12293) <= a or b;
    layer3_outputs(12294) <= '1';
    layer3_outputs(12295) <= a;
    layer3_outputs(12296) <= a or b;
    layer3_outputs(12297) <= a or b;
    layer3_outputs(12298) <= not (a xor b);
    layer3_outputs(12299) <= a and b;
    layer3_outputs(12300) <= not b or a;
    layer3_outputs(12301) <= not (a xor b);
    layer3_outputs(12302) <= '0';
    layer3_outputs(12303) <= not a;
    layer3_outputs(12304) <= a or b;
    layer3_outputs(12305) <= b;
    layer3_outputs(12306) <= a or b;
    layer3_outputs(12307) <= a and not b;
    layer3_outputs(12308) <= '1';
    layer3_outputs(12309) <= not b;
    layer3_outputs(12310) <= not a;
    layer3_outputs(12311) <= not a or b;
    layer3_outputs(12312) <= not b;
    layer3_outputs(12313) <= b and not a;
    layer3_outputs(12314) <= a or b;
    layer3_outputs(12315) <= not b;
    layer3_outputs(12316) <= '0';
    layer3_outputs(12317) <= a xor b;
    layer3_outputs(12318) <= not a or b;
    layer3_outputs(12319) <= '0';
    layer3_outputs(12320) <= b;
    layer3_outputs(12321) <= a xor b;
    layer3_outputs(12322) <= not b;
    layer3_outputs(12323) <= b;
    layer3_outputs(12324) <= b;
    layer3_outputs(12325) <= b;
    layer3_outputs(12326) <= a;
    layer3_outputs(12327) <= b;
    layer3_outputs(12328) <= not a;
    layer3_outputs(12329) <= '1';
    layer3_outputs(12330) <= '1';
    layer3_outputs(12331) <= a;
    layer3_outputs(12332) <= not b;
    layer3_outputs(12333) <= not a or b;
    layer3_outputs(12334) <= not a or b;
    layer3_outputs(12335) <= a and not b;
    layer3_outputs(12336) <= a and not b;
    layer3_outputs(12337) <= '0';
    layer3_outputs(12338) <= b and not a;
    layer3_outputs(12339) <= not a;
    layer3_outputs(12340) <= b;
    layer3_outputs(12341) <= '0';
    layer3_outputs(12342) <= not (a and b);
    layer3_outputs(12343) <= not b;
    layer3_outputs(12344) <= not (a and b);
    layer3_outputs(12345) <= '0';
    layer3_outputs(12346) <= not b;
    layer3_outputs(12347) <= not b;
    layer3_outputs(12348) <= b;
    layer3_outputs(12349) <= not (a and b);
    layer3_outputs(12350) <= a;
    layer3_outputs(12351) <= not (a or b);
    layer3_outputs(12352) <= not (a xor b);
    layer3_outputs(12353) <= not a;
    layer3_outputs(12354) <= not b;
    layer3_outputs(12355) <= a;
    layer3_outputs(12356) <= '1';
    layer3_outputs(12357) <= not b or a;
    layer3_outputs(12358) <= not a or b;
    layer3_outputs(12359) <= b;
    layer3_outputs(12360) <= not b or a;
    layer3_outputs(12361) <= not a or b;
    layer3_outputs(12362) <= b and not a;
    layer3_outputs(12363) <= a and not b;
    layer3_outputs(12364) <= a and b;
    layer3_outputs(12365) <= b;
    layer3_outputs(12366) <= not (a and b);
    layer3_outputs(12367) <= a;
    layer3_outputs(12368) <= b;
    layer3_outputs(12369) <= b;
    layer3_outputs(12370) <= '0';
    layer3_outputs(12371) <= a;
    layer3_outputs(12372) <= not b or a;
    layer3_outputs(12373) <= a;
    layer3_outputs(12374) <= b;
    layer3_outputs(12375) <= '0';
    layer3_outputs(12376) <= not (a or b);
    layer3_outputs(12377) <= a and b;
    layer3_outputs(12378) <= a xor b;
    layer3_outputs(12379) <= a xor b;
    layer3_outputs(12380) <= a;
    layer3_outputs(12381) <= not b;
    layer3_outputs(12382) <= not a or b;
    layer3_outputs(12383) <= not a;
    layer3_outputs(12384) <= '1';
    layer3_outputs(12385) <= '1';
    layer3_outputs(12386) <= not b or a;
    layer3_outputs(12387) <= not a;
    layer3_outputs(12388) <= '1';
    layer3_outputs(12389) <= b and not a;
    layer3_outputs(12390) <= not (a and b);
    layer3_outputs(12391) <= not b or a;
    layer3_outputs(12392) <= '1';
    layer3_outputs(12393) <= a;
    layer3_outputs(12394) <= not a or b;
    layer3_outputs(12395) <= not b;
    layer3_outputs(12396) <= not (a xor b);
    layer3_outputs(12397) <= not b;
    layer3_outputs(12398) <= b;
    layer3_outputs(12399) <= not b or a;
    layer3_outputs(12400) <= b;
    layer3_outputs(12401) <= a and b;
    layer3_outputs(12402) <= not b or a;
    layer3_outputs(12403) <= not a or b;
    layer3_outputs(12404) <= a and b;
    layer3_outputs(12405) <= not a or b;
    layer3_outputs(12406) <= not a;
    layer3_outputs(12407) <= not a or b;
    layer3_outputs(12408) <= '0';
    layer3_outputs(12409) <= not b;
    layer3_outputs(12410) <= b;
    layer3_outputs(12411) <= not b;
    layer3_outputs(12412) <= not a or b;
    layer3_outputs(12413) <= '0';
    layer3_outputs(12414) <= a or b;
    layer3_outputs(12415) <= not b or a;
    layer3_outputs(12416) <= not (a or b);
    layer3_outputs(12417) <= '0';
    layer3_outputs(12418) <= a and not b;
    layer3_outputs(12419) <= a;
    layer3_outputs(12420) <= b;
    layer3_outputs(12421) <= a and not b;
    layer3_outputs(12422) <= not a or b;
    layer3_outputs(12423) <= a;
    layer3_outputs(12424) <= a and b;
    layer3_outputs(12425) <= not (a or b);
    layer3_outputs(12426) <= a;
    layer3_outputs(12427) <= a xor b;
    layer3_outputs(12428) <= a or b;
    layer3_outputs(12429) <= not b;
    layer3_outputs(12430) <= not (a and b);
    layer3_outputs(12431) <= not (a and b);
    layer3_outputs(12432) <= b and not a;
    layer3_outputs(12433) <= a and not b;
    layer3_outputs(12434) <= b and not a;
    layer3_outputs(12435) <= not (a and b);
    layer3_outputs(12436) <= a or b;
    layer3_outputs(12437) <= '1';
    layer3_outputs(12438) <= a and b;
    layer3_outputs(12439) <= b;
    layer3_outputs(12440) <= a;
    layer3_outputs(12441) <= not a;
    layer3_outputs(12442) <= b;
    layer3_outputs(12443) <= a and b;
    layer3_outputs(12444) <= a or b;
    layer3_outputs(12445) <= a or b;
    layer3_outputs(12446) <= b and not a;
    layer3_outputs(12447) <= not a;
    layer3_outputs(12448) <= a and not b;
    layer3_outputs(12449) <= '1';
    layer3_outputs(12450) <= not a or b;
    layer3_outputs(12451) <= not b;
    layer3_outputs(12452) <= not a or b;
    layer3_outputs(12453) <= not (a and b);
    layer3_outputs(12454) <= a or b;
    layer3_outputs(12455) <= not b;
    layer3_outputs(12456) <= not a;
    layer3_outputs(12457) <= not b or a;
    layer3_outputs(12458) <= not (a or b);
    layer3_outputs(12459) <= not (a or b);
    layer3_outputs(12460) <= b and not a;
    layer3_outputs(12461) <= a and not b;
    layer3_outputs(12462) <= '0';
    layer3_outputs(12463) <= b;
    layer3_outputs(12464) <= a and b;
    layer3_outputs(12465) <= not a;
    layer3_outputs(12466) <= a and b;
    layer3_outputs(12467) <= not a or b;
    layer3_outputs(12468) <= not (a and b);
    layer3_outputs(12469) <= not b;
    layer3_outputs(12470) <= a xor b;
    layer3_outputs(12471) <= a and not b;
    layer3_outputs(12472) <= b and not a;
    layer3_outputs(12473) <= b;
    layer3_outputs(12474) <= a and b;
    layer3_outputs(12475) <= a;
    layer3_outputs(12476) <= b and not a;
    layer3_outputs(12477) <= b and not a;
    layer3_outputs(12478) <= a or b;
    layer3_outputs(12479) <= '0';
    layer3_outputs(12480) <= b;
    layer3_outputs(12481) <= not (a or b);
    layer3_outputs(12482) <= a;
    layer3_outputs(12483) <= not a or b;
    layer3_outputs(12484) <= b;
    layer3_outputs(12485) <= '0';
    layer3_outputs(12486) <= not (a xor b);
    layer3_outputs(12487) <= a and b;
    layer3_outputs(12488) <= b;
    layer3_outputs(12489) <= not a;
    layer3_outputs(12490) <= a;
    layer3_outputs(12491) <= a and b;
    layer3_outputs(12492) <= not b;
    layer3_outputs(12493) <= not (a or b);
    layer3_outputs(12494) <= not (a and b);
    layer3_outputs(12495) <= '0';
    layer3_outputs(12496) <= not a;
    layer3_outputs(12497) <= a and not b;
    layer3_outputs(12498) <= not a;
    layer3_outputs(12499) <= a or b;
    layer3_outputs(12500) <= a;
    layer3_outputs(12501) <= not b or a;
    layer3_outputs(12502) <= b;
    layer3_outputs(12503) <= b;
    layer3_outputs(12504) <= not b;
    layer3_outputs(12505) <= a and b;
    layer3_outputs(12506) <= a or b;
    layer3_outputs(12507) <= b;
    layer3_outputs(12508) <= '0';
    layer3_outputs(12509) <= not a or b;
    layer3_outputs(12510) <= b;
    layer3_outputs(12511) <= not b;
    layer3_outputs(12512) <= a and not b;
    layer3_outputs(12513) <= '0';
    layer3_outputs(12514) <= '1';
    layer3_outputs(12515) <= a;
    layer3_outputs(12516) <= not a or b;
    layer3_outputs(12517) <= a or b;
    layer3_outputs(12518) <= not (a and b);
    layer3_outputs(12519) <= b;
    layer3_outputs(12520) <= not b;
    layer3_outputs(12521) <= not (a and b);
    layer3_outputs(12522) <= a;
    layer3_outputs(12523) <= b and not a;
    layer3_outputs(12524) <= not a;
    layer3_outputs(12525) <= not b or a;
    layer3_outputs(12526) <= not (a or b);
    layer3_outputs(12527) <= not b;
    layer3_outputs(12528) <= b;
    layer3_outputs(12529) <= not b;
    layer3_outputs(12530) <= not b or a;
    layer3_outputs(12531) <= b;
    layer3_outputs(12532) <= not (a or b);
    layer3_outputs(12533) <= a and b;
    layer3_outputs(12534) <= not (a or b);
    layer3_outputs(12535) <= a;
    layer3_outputs(12536) <= a;
    layer3_outputs(12537) <= not (a or b);
    layer3_outputs(12538) <= not (a xor b);
    layer3_outputs(12539) <= b;
    layer3_outputs(12540) <= not (a or b);
    layer3_outputs(12541) <= a xor b;
    layer3_outputs(12542) <= not (a and b);
    layer3_outputs(12543) <= not a;
    layer3_outputs(12544) <= not a;
    layer3_outputs(12545) <= not b;
    layer3_outputs(12546) <= b;
    layer3_outputs(12547) <= a;
    layer3_outputs(12548) <= not b or a;
    layer3_outputs(12549) <= not a;
    layer3_outputs(12550) <= not b;
    layer3_outputs(12551) <= '0';
    layer3_outputs(12552) <= not b or a;
    layer3_outputs(12553) <= b;
    layer3_outputs(12554) <= a xor b;
    layer3_outputs(12555) <= not (a xor b);
    layer3_outputs(12556) <= not a or b;
    layer3_outputs(12557) <= b and not a;
    layer3_outputs(12558) <= not (a xor b);
    layer3_outputs(12559) <= not a or b;
    layer3_outputs(12560) <= a and not b;
    layer3_outputs(12561) <= a;
    layer3_outputs(12562) <= not a;
    layer3_outputs(12563) <= b;
    layer3_outputs(12564) <= a and b;
    layer3_outputs(12565) <= b;
    layer3_outputs(12566) <= a and not b;
    layer3_outputs(12567) <= not (a xor b);
    layer3_outputs(12568) <= a xor b;
    layer3_outputs(12569) <= not a;
    layer3_outputs(12570) <= a and b;
    layer3_outputs(12571) <= a and not b;
    layer3_outputs(12572) <= not (a xor b);
    layer3_outputs(12573) <= not a;
    layer3_outputs(12574) <= b;
    layer3_outputs(12575) <= not a or b;
    layer3_outputs(12576) <= a or b;
    layer3_outputs(12577) <= a and b;
    layer3_outputs(12578) <= a and b;
    layer3_outputs(12579) <= '1';
    layer3_outputs(12580) <= b;
    layer3_outputs(12581) <= not (a or b);
    layer3_outputs(12582) <= not (a and b);
    layer3_outputs(12583) <= not b;
    layer3_outputs(12584) <= not (a xor b);
    layer3_outputs(12585) <= not (a or b);
    layer3_outputs(12586) <= b;
    layer3_outputs(12587) <= b;
    layer3_outputs(12588) <= a and b;
    layer3_outputs(12589) <= b;
    layer3_outputs(12590) <= not (a or b);
    layer3_outputs(12591) <= a;
    layer3_outputs(12592) <= not b;
    layer3_outputs(12593) <= b;
    layer3_outputs(12594) <= not a;
    layer3_outputs(12595) <= b;
    layer3_outputs(12596) <= a and b;
    layer3_outputs(12597) <= a and b;
    layer3_outputs(12598) <= not a;
    layer3_outputs(12599) <= '0';
    layer3_outputs(12600) <= not (a xor b);
    layer3_outputs(12601) <= not (a and b);
    layer3_outputs(12602) <= a xor b;
    layer3_outputs(12603) <= a or b;
    layer3_outputs(12604) <= b;
    layer3_outputs(12605) <= a and not b;
    layer3_outputs(12606) <= not b;
    layer3_outputs(12607) <= not a;
    layer3_outputs(12608) <= a and b;
    layer3_outputs(12609) <= not a;
    layer3_outputs(12610) <= b and not a;
    layer3_outputs(12611) <= b;
    layer3_outputs(12612) <= b and not a;
    layer3_outputs(12613) <= not (a or b);
    layer3_outputs(12614) <= not a;
    layer3_outputs(12615) <= a and not b;
    layer3_outputs(12616) <= not a or b;
    layer3_outputs(12617) <= a and not b;
    layer3_outputs(12618) <= not a;
    layer3_outputs(12619) <= a;
    layer3_outputs(12620) <= not b or a;
    layer3_outputs(12621) <= a and not b;
    layer3_outputs(12622) <= not a;
    layer3_outputs(12623) <= not b;
    layer3_outputs(12624) <= not (a xor b);
    layer3_outputs(12625) <= b;
    layer3_outputs(12626) <= '0';
    layer3_outputs(12627) <= a or b;
    layer3_outputs(12628) <= '0';
    layer3_outputs(12629) <= not a;
    layer3_outputs(12630) <= not a or b;
    layer3_outputs(12631) <= a;
    layer3_outputs(12632) <= a;
    layer3_outputs(12633) <= a;
    layer3_outputs(12634) <= a;
    layer3_outputs(12635) <= not b or a;
    layer3_outputs(12636) <= not b;
    layer3_outputs(12637) <= a;
    layer3_outputs(12638) <= '0';
    layer3_outputs(12639) <= a xor b;
    layer3_outputs(12640) <= '1';
    layer3_outputs(12641) <= not b;
    layer3_outputs(12642) <= not a or b;
    layer3_outputs(12643) <= not b;
    layer3_outputs(12644) <= not a or b;
    layer3_outputs(12645) <= not (a or b);
    layer3_outputs(12646) <= a and not b;
    layer3_outputs(12647) <= not b;
    layer3_outputs(12648) <= a;
    layer3_outputs(12649) <= a and b;
    layer3_outputs(12650) <= a xor b;
    layer3_outputs(12651) <= not b or a;
    layer3_outputs(12652) <= not (a and b);
    layer3_outputs(12653) <= not (a and b);
    layer3_outputs(12654) <= not b or a;
    layer3_outputs(12655) <= not a;
    layer3_outputs(12656) <= not (a xor b);
    layer3_outputs(12657) <= not a;
    layer3_outputs(12658) <= a or b;
    layer3_outputs(12659) <= not a or b;
    layer3_outputs(12660) <= b;
    layer3_outputs(12661) <= a and not b;
    layer3_outputs(12662) <= not (a or b);
    layer3_outputs(12663) <= a and not b;
    layer3_outputs(12664) <= b and not a;
    layer3_outputs(12665) <= a;
    layer3_outputs(12666) <= b and not a;
    layer3_outputs(12667) <= a and b;
    layer3_outputs(12668) <= a or b;
    layer3_outputs(12669) <= a;
    layer3_outputs(12670) <= not a;
    layer3_outputs(12671) <= a;
    layer3_outputs(12672) <= not b;
    layer3_outputs(12673) <= not (a xor b);
    layer3_outputs(12674) <= a and b;
    layer3_outputs(12675) <= a and b;
    layer3_outputs(12676) <= not (a xor b);
    layer3_outputs(12677) <= a or b;
    layer3_outputs(12678) <= a;
    layer3_outputs(12679) <= b and not a;
    layer3_outputs(12680) <= b;
    layer3_outputs(12681) <= '0';
    layer3_outputs(12682) <= '1';
    layer3_outputs(12683) <= a or b;
    layer3_outputs(12684) <= not a or b;
    layer3_outputs(12685) <= a;
    layer3_outputs(12686) <= not (a xor b);
    layer3_outputs(12687) <= b;
    layer3_outputs(12688) <= not a;
    layer3_outputs(12689) <= not b;
    layer3_outputs(12690) <= not b;
    layer3_outputs(12691) <= not b;
    layer3_outputs(12692) <= b and not a;
    layer3_outputs(12693) <= not b;
    layer3_outputs(12694) <= not (a xor b);
    layer3_outputs(12695) <= not a or b;
    layer3_outputs(12696) <= b and not a;
    layer3_outputs(12697) <= not (a and b);
    layer3_outputs(12698) <= not b or a;
    layer3_outputs(12699) <= b;
    layer3_outputs(12700) <= '0';
    layer3_outputs(12701) <= a and b;
    layer3_outputs(12702) <= b;
    layer3_outputs(12703) <= a;
    layer3_outputs(12704) <= a or b;
    layer3_outputs(12705) <= b;
    layer3_outputs(12706) <= not (a and b);
    layer3_outputs(12707) <= not b or a;
    layer3_outputs(12708) <= not a or b;
    layer3_outputs(12709) <= b;
    layer3_outputs(12710) <= b and not a;
    layer3_outputs(12711) <= a xor b;
    layer3_outputs(12712) <= not b;
    layer3_outputs(12713) <= a and b;
    layer3_outputs(12714) <= a and not b;
    layer3_outputs(12715) <= not b or a;
    layer3_outputs(12716) <= a and b;
    layer3_outputs(12717) <= not b;
    layer3_outputs(12718) <= not (a and b);
    layer3_outputs(12719) <= not (a or b);
    layer3_outputs(12720) <= b;
    layer3_outputs(12721) <= a and not b;
    layer3_outputs(12722) <= a and b;
    layer3_outputs(12723) <= a and not b;
    layer3_outputs(12724) <= not (a and b);
    layer3_outputs(12725) <= not (a xor b);
    layer3_outputs(12726) <= not a or b;
    layer3_outputs(12727) <= a;
    layer3_outputs(12728) <= not b;
    layer3_outputs(12729) <= not b;
    layer3_outputs(12730) <= '1';
    layer3_outputs(12731) <= not b or a;
    layer3_outputs(12732) <= not a;
    layer3_outputs(12733) <= a xor b;
    layer3_outputs(12734) <= not (a or b);
    layer3_outputs(12735) <= b;
    layer3_outputs(12736) <= not b;
    layer3_outputs(12737) <= not (a xor b);
    layer3_outputs(12738) <= b;
    layer3_outputs(12739) <= a;
    layer3_outputs(12740) <= b;
    layer3_outputs(12741) <= not a or b;
    layer3_outputs(12742) <= '0';
    layer3_outputs(12743) <= b and not a;
    layer3_outputs(12744) <= not b;
    layer3_outputs(12745) <= not (a or b);
    layer3_outputs(12746) <= a xor b;
    layer3_outputs(12747) <= not b;
    layer3_outputs(12748) <= not (a and b);
    layer3_outputs(12749) <= not a or b;
    layer3_outputs(12750) <= not (a and b);
    layer3_outputs(12751) <= a and b;
    layer3_outputs(12752) <= '0';
    layer3_outputs(12753) <= a and not b;
    layer3_outputs(12754) <= not a;
    layer3_outputs(12755) <= a xor b;
    layer3_outputs(12756) <= '0';
    layer3_outputs(12757) <= not a or b;
    layer3_outputs(12758) <= b;
    layer3_outputs(12759) <= a or b;
    layer3_outputs(12760) <= not b or a;
    layer3_outputs(12761) <= not b or a;
    layer3_outputs(12762) <= a;
    layer3_outputs(12763) <= b and not a;
    layer3_outputs(12764) <= a;
    layer3_outputs(12765) <= not (a or b);
    layer3_outputs(12766) <= not b;
    layer3_outputs(12767) <= a xor b;
    layer3_outputs(12768) <= b;
    layer3_outputs(12769) <= b and not a;
    layer3_outputs(12770) <= not a or b;
    layer3_outputs(12771) <= a;
    layer3_outputs(12772) <= not a or b;
    layer3_outputs(12773) <= not b;
    layer3_outputs(12774) <= b and not a;
    layer3_outputs(12775) <= not (a or b);
    layer3_outputs(12776) <= b;
    layer3_outputs(12777) <= a;
    layer3_outputs(12778) <= not (a or b);
    layer3_outputs(12779) <= not (a and b);
    layer3_outputs(12780) <= b and not a;
    layer3_outputs(12781) <= not b or a;
    layer3_outputs(12782) <= a and b;
    layer3_outputs(12783) <= not (a xor b);
    layer3_outputs(12784) <= not a or b;
    layer3_outputs(12785) <= '1';
    layer3_outputs(12786) <= not b;
    layer3_outputs(12787) <= a and not b;
    layer3_outputs(12788) <= a;
    layer3_outputs(12789) <= not b;
    layer3_outputs(12790) <= a and b;
    layer3_outputs(12791) <= a;
    layer3_outputs(12792) <= a or b;
    layer3_outputs(12793) <= a;
    layer3_outputs(12794) <= not a or b;
    layer3_outputs(12795) <= not b;
    layer3_outputs(12796) <= b;
    layer3_outputs(12797) <= '0';
    layer3_outputs(12798) <= a;
    layer3_outputs(12799) <= not b;
    layer4_outputs(0) <= not (a or b);
    layer4_outputs(1) <= not b;
    layer4_outputs(2) <= a or b;
    layer4_outputs(3) <= not (a or b);
    layer4_outputs(4) <= not a;
    layer4_outputs(5) <= a and b;
    layer4_outputs(6) <= not a or b;
    layer4_outputs(7) <= a and not b;
    layer4_outputs(8) <= b;
    layer4_outputs(9) <= not b or a;
    layer4_outputs(10) <= a xor b;
    layer4_outputs(11) <= not (a xor b);
    layer4_outputs(12) <= a;
    layer4_outputs(13) <= a and b;
    layer4_outputs(14) <= '1';
    layer4_outputs(15) <= not (a or b);
    layer4_outputs(16) <= b;
    layer4_outputs(17) <= b;
    layer4_outputs(18) <= not a;
    layer4_outputs(19) <= b;
    layer4_outputs(20) <= b;
    layer4_outputs(21) <= a;
    layer4_outputs(22) <= not a;
    layer4_outputs(23) <= not a or b;
    layer4_outputs(24) <= not (a and b);
    layer4_outputs(25) <= not (a and b);
    layer4_outputs(26) <= not a;
    layer4_outputs(27) <= b;
    layer4_outputs(28) <= a;
    layer4_outputs(29) <= not (a xor b);
    layer4_outputs(30) <= not (a or b);
    layer4_outputs(31) <= not b;
    layer4_outputs(32) <= a or b;
    layer4_outputs(33) <= '1';
    layer4_outputs(34) <= a or b;
    layer4_outputs(35) <= not a;
    layer4_outputs(36) <= not (a xor b);
    layer4_outputs(37) <= a and b;
    layer4_outputs(38) <= not b;
    layer4_outputs(39) <= a and not b;
    layer4_outputs(40) <= a;
    layer4_outputs(41) <= not a or b;
    layer4_outputs(42) <= '1';
    layer4_outputs(43) <= not (a xor b);
    layer4_outputs(44) <= b;
    layer4_outputs(45) <= b and not a;
    layer4_outputs(46) <= a and not b;
    layer4_outputs(47) <= not a or b;
    layer4_outputs(48) <= not b or a;
    layer4_outputs(49) <= not b;
    layer4_outputs(50) <= a and b;
    layer4_outputs(51) <= a;
    layer4_outputs(52) <= a;
    layer4_outputs(53) <= a and b;
    layer4_outputs(54) <= a;
    layer4_outputs(55) <= b;
    layer4_outputs(56) <= not b;
    layer4_outputs(57) <= a and not b;
    layer4_outputs(58) <= not a;
    layer4_outputs(59) <= a and not b;
    layer4_outputs(60) <= a;
    layer4_outputs(61) <= a;
    layer4_outputs(62) <= b and not a;
    layer4_outputs(63) <= a and not b;
    layer4_outputs(64) <= b and not a;
    layer4_outputs(65) <= a;
    layer4_outputs(66) <= not a or b;
    layer4_outputs(67) <= a xor b;
    layer4_outputs(68) <= not (a or b);
    layer4_outputs(69) <= not a;
    layer4_outputs(70) <= not b;
    layer4_outputs(71) <= not b;
    layer4_outputs(72) <= not (a and b);
    layer4_outputs(73) <= not b;
    layer4_outputs(74) <= b;
    layer4_outputs(75) <= b;
    layer4_outputs(76) <= a xor b;
    layer4_outputs(77) <= a;
    layer4_outputs(78) <= a and b;
    layer4_outputs(79) <= a or b;
    layer4_outputs(80) <= not (a or b);
    layer4_outputs(81) <= not b;
    layer4_outputs(82) <= not a or b;
    layer4_outputs(83) <= a xor b;
    layer4_outputs(84) <= a or b;
    layer4_outputs(85) <= not (a and b);
    layer4_outputs(86) <= '0';
    layer4_outputs(87) <= a;
    layer4_outputs(88) <= a;
    layer4_outputs(89) <= not (a and b);
    layer4_outputs(90) <= not a;
    layer4_outputs(91) <= not b;
    layer4_outputs(92) <= not a or b;
    layer4_outputs(93) <= a and b;
    layer4_outputs(94) <= not a;
    layer4_outputs(95) <= not (a xor b);
    layer4_outputs(96) <= a and not b;
    layer4_outputs(97) <= not a or b;
    layer4_outputs(98) <= not b;
    layer4_outputs(99) <= not a;
    layer4_outputs(100) <= not (a or b);
    layer4_outputs(101) <= not b or a;
    layer4_outputs(102) <= a;
    layer4_outputs(103) <= b and not a;
    layer4_outputs(104) <= not b;
    layer4_outputs(105) <= a or b;
    layer4_outputs(106) <= not a or b;
    layer4_outputs(107) <= not b;
    layer4_outputs(108) <= a or b;
    layer4_outputs(109) <= b;
    layer4_outputs(110) <= a or b;
    layer4_outputs(111) <= not a;
    layer4_outputs(112) <= a and not b;
    layer4_outputs(113) <= not a or b;
    layer4_outputs(114) <= a and b;
    layer4_outputs(115) <= not a;
    layer4_outputs(116) <= a and b;
    layer4_outputs(117) <= not a or b;
    layer4_outputs(118) <= a;
    layer4_outputs(119) <= not (a or b);
    layer4_outputs(120) <= not (a xor b);
    layer4_outputs(121) <= not a or b;
    layer4_outputs(122) <= not (a xor b);
    layer4_outputs(123) <= not (a xor b);
    layer4_outputs(124) <= '0';
    layer4_outputs(125) <= not a or b;
    layer4_outputs(126) <= not a or b;
    layer4_outputs(127) <= a or b;
    layer4_outputs(128) <= not a or b;
    layer4_outputs(129) <= a and not b;
    layer4_outputs(130) <= b;
    layer4_outputs(131) <= not b or a;
    layer4_outputs(132) <= a xor b;
    layer4_outputs(133) <= not b;
    layer4_outputs(134) <= not a;
    layer4_outputs(135) <= not (a or b);
    layer4_outputs(136) <= not (a xor b);
    layer4_outputs(137) <= not b;
    layer4_outputs(138) <= b;
    layer4_outputs(139) <= not b;
    layer4_outputs(140) <= a and not b;
    layer4_outputs(141) <= a and not b;
    layer4_outputs(142) <= not (a or b);
    layer4_outputs(143) <= not a;
    layer4_outputs(144) <= not (a xor b);
    layer4_outputs(145) <= a xor b;
    layer4_outputs(146) <= a;
    layer4_outputs(147) <= b;
    layer4_outputs(148) <= a;
    layer4_outputs(149) <= not (a and b);
    layer4_outputs(150) <= not (a and b);
    layer4_outputs(151) <= b;
    layer4_outputs(152) <= not a or b;
    layer4_outputs(153) <= a and not b;
    layer4_outputs(154) <= b;
    layer4_outputs(155) <= a xor b;
    layer4_outputs(156) <= not a;
    layer4_outputs(157) <= a and b;
    layer4_outputs(158) <= not (a and b);
    layer4_outputs(159) <= a or b;
    layer4_outputs(160) <= not (a or b);
    layer4_outputs(161) <= not a;
    layer4_outputs(162) <= b and not a;
    layer4_outputs(163) <= not (a and b);
    layer4_outputs(164) <= a;
    layer4_outputs(165) <= not a;
    layer4_outputs(166) <= a xor b;
    layer4_outputs(167) <= not (a and b);
    layer4_outputs(168) <= a xor b;
    layer4_outputs(169) <= a and not b;
    layer4_outputs(170) <= a;
    layer4_outputs(171) <= not b;
    layer4_outputs(172) <= not (a or b);
    layer4_outputs(173) <= not b;
    layer4_outputs(174) <= not (a or b);
    layer4_outputs(175) <= b;
    layer4_outputs(176) <= not (a or b);
    layer4_outputs(177) <= not (a or b);
    layer4_outputs(178) <= not b;
    layer4_outputs(179) <= a;
    layer4_outputs(180) <= a;
    layer4_outputs(181) <= b;
    layer4_outputs(182) <= not (a and b);
    layer4_outputs(183) <= not (a and b);
    layer4_outputs(184) <= a;
    layer4_outputs(185) <= not b;
    layer4_outputs(186) <= not (a or b);
    layer4_outputs(187) <= not a;
    layer4_outputs(188) <= a or b;
    layer4_outputs(189) <= b;
    layer4_outputs(190) <= not a;
    layer4_outputs(191) <= not (a and b);
    layer4_outputs(192) <= not a;
    layer4_outputs(193) <= not a or b;
    layer4_outputs(194) <= a and b;
    layer4_outputs(195) <= a xor b;
    layer4_outputs(196) <= not (a xor b);
    layer4_outputs(197) <= a xor b;
    layer4_outputs(198) <= b and not a;
    layer4_outputs(199) <= b;
    layer4_outputs(200) <= a and not b;
    layer4_outputs(201) <= b and not a;
    layer4_outputs(202) <= b and not a;
    layer4_outputs(203) <= b;
    layer4_outputs(204) <= a;
    layer4_outputs(205) <= a;
    layer4_outputs(206) <= not a;
    layer4_outputs(207) <= not a or b;
    layer4_outputs(208) <= a;
    layer4_outputs(209) <= a or b;
    layer4_outputs(210) <= a and b;
    layer4_outputs(211) <= a or b;
    layer4_outputs(212) <= not (a or b);
    layer4_outputs(213) <= '0';
    layer4_outputs(214) <= not b;
    layer4_outputs(215) <= a xor b;
    layer4_outputs(216) <= not a;
    layer4_outputs(217) <= not (a or b);
    layer4_outputs(218) <= a and not b;
    layer4_outputs(219) <= a or b;
    layer4_outputs(220) <= a;
    layer4_outputs(221) <= not a or b;
    layer4_outputs(222) <= not b;
    layer4_outputs(223) <= b and not a;
    layer4_outputs(224) <= not b;
    layer4_outputs(225) <= a or b;
    layer4_outputs(226) <= b and not a;
    layer4_outputs(227) <= not b;
    layer4_outputs(228) <= not a;
    layer4_outputs(229) <= not a;
    layer4_outputs(230) <= a and not b;
    layer4_outputs(231) <= a;
    layer4_outputs(232) <= not a or b;
    layer4_outputs(233) <= not (a xor b);
    layer4_outputs(234) <= not (a or b);
    layer4_outputs(235) <= not (a and b);
    layer4_outputs(236) <= b;
    layer4_outputs(237) <= a;
    layer4_outputs(238) <= not b;
    layer4_outputs(239) <= '1';
    layer4_outputs(240) <= not b or a;
    layer4_outputs(241) <= not (a and b);
    layer4_outputs(242) <= a and b;
    layer4_outputs(243) <= a or b;
    layer4_outputs(244) <= not (a and b);
    layer4_outputs(245) <= b;
    layer4_outputs(246) <= not a;
    layer4_outputs(247) <= not (a and b);
    layer4_outputs(248) <= a;
    layer4_outputs(249) <= not (a xor b);
    layer4_outputs(250) <= a;
    layer4_outputs(251) <= b;
    layer4_outputs(252) <= b and not a;
    layer4_outputs(253) <= not a or b;
    layer4_outputs(254) <= a;
    layer4_outputs(255) <= not (a and b);
    layer4_outputs(256) <= a or b;
    layer4_outputs(257) <= not (a or b);
    layer4_outputs(258) <= not (a or b);
    layer4_outputs(259) <= not (a and b);
    layer4_outputs(260) <= b;
    layer4_outputs(261) <= not b;
    layer4_outputs(262) <= b and not a;
    layer4_outputs(263) <= a xor b;
    layer4_outputs(264) <= not b or a;
    layer4_outputs(265) <= not a;
    layer4_outputs(266) <= a xor b;
    layer4_outputs(267) <= not b;
    layer4_outputs(268) <= not b;
    layer4_outputs(269) <= a and b;
    layer4_outputs(270) <= not b or a;
    layer4_outputs(271) <= b;
    layer4_outputs(272) <= a;
    layer4_outputs(273) <= not b;
    layer4_outputs(274) <= not (a xor b);
    layer4_outputs(275) <= not (a and b);
    layer4_outputs(276) <= b and not a;
    layer4_outputs(277) <= a xor b;
    layer4_outputs(278) <= not (a or b);
    layer4_outputs(279) <= not a;
    layer4_outputs(280) <= a and not b;
    layer4_outputs(281) <= not a;
    layer4_outputs(282) <= not b;
    layer4_outputs(283) <= not (a xor b);
    layer4_outputs(284) <= not a;
    layer4_outputs(285) <= a;
    layer4_outputs(286) <= '1';
    layer4_outputs(287) <= not b or a;
    layer4_outputs(288) <= not a;
    layer4_outputs(289) <= not (a or b);
    layer4_outputs(290) <= a and not b;
    layer4_outputs(291) <= a or b;
    layer4_outputs(292) <= not (a xor b);
    layer4_outputs(293) <= not a or b;
    layer4_outputs(294) <= b and not a;
    layer4_outputs(295) <= a;
    layer4_outputs(296) <= not b;
    layer4_outputs(297) <= a;
    layer4_outputs(298) <= '1';
    layer4_outputs(299) <= not (a and b);
    layer4_outputs(300) <= not a;
    layer4_outputs(301) <= not (a or b);
    layer4_outputs(302) <= b;
    layer4_outputs(303) <= not b;
    layer4_outputs(304) <= not b;
    layer4_outputs(305) <= a;
    layer4_outputs(306) <= not (a and b);
    layer4_outputs(307) <= not b;
    layer4_outputs(308) <= not a;
    layer4_outputs(309) <= not a;
    layer4_outputs(310) <= not (a or b);
    layer4_outputs(311) <= not a;
    layer4_outputs(312) <= b;
    layer4_outputs(313) <= a;
    layer4_outputs(314) <= b;
    layer4_outputs(315) <= not b;
    layer4_outputs(316) <= a;
    layer4_outputs(317) <= a xor b;
    layer4_outputs(318) <= not a;
    layer4_outputs(319) <= not (a xor b);
    layer4_outputs(320) <= a;
    layer4_outputs(321) <= b;
    layer4_outputs(322) <= not (a xor b);
    layer4_outputs(323) <= not a;
    layer4_outputs(324) <= not a;
    layer4_outputs(325) <= not a;
    layer4_outputs(326) <= a xor b;
    layer4_outputs(327) <= '0';
    layer4_outputs(328) <= a xor b;
    layer4_outputs(329) <= b and not a;
    layer4_outputs(330) <= b;
    layer4_outputs(331) <= not a;
    layer4_outputs(332) <= not b;
    layer4_outputs(333) <= b;
    layer4_outputs(334) <= not b or a;
    layer4_outputs(335) <= not b or a;
    layer4_outputs(336) <= not a;
    layer4_outputs(337) <= a;
    layer4_outputs(338) <= not (a and b);
    layer4_outputs(339) <= not b;
    layer4_outputs(340) <= a;
    layer4_outputs(341) <= '1';
    layer4_outputs(342) <= not (a or b);
    layer4_outputs(343) <= not a or b;
    layer4_outputs(344) <= '0';
    layer4_outputs(345) <= not b;
    layer4_outputs(346) <= a;
    layer4_outputs(347) <= not a;
    layer4_outputs(348) <= not a or b;
    layer4_outputs(349) <= a and b;
    layer4_outputs(350) <= b;
    layer4_outputs(351) <= a;
    layer4_outputs(352) <= a xor b;
    layer4_outputs(353) <= not (a or b);
    layer4_outputs(354) <= b;
    layer4_outputs(355) <= b and not a;
    layer4_outputs(356) <= a or b;
    layer4_outputs(357) <= not a or b;
    layer4_outputs(358) <= '1';
    layer4_outputs(359) <= b;
    layer4_outputs(360) <= a xor b;
    layer4_outputs(361) <= a or b;
    layer4_outputs(362) <= b and not a;
    layer4_outputs(363) <= not (a or b);
    layer4_outputs(364) <= not b;
    layer4_outputs(365) <= b and not a;
    layer4_outputs(366) <= a xor b;
    layer4_outputs(367) <= not b or a;
    layer4_outputs(368) <= a and b;
    layer4_outputs(369) <= a;
    layer4_outputs(370) <= not a;
    layer4_outputs(371) <= '1';
    layer4_outputs(372) <= not a or b;
    layer4_outputs(373) <= a and not b;
    layer4_outputs(374) <= a;
    layer4_outputs(375) <= b;
    layer4_outputs(376) <= not a or b;
    layer4_outputs(377) <= not b or a;
    layer4_outputs(378) <= not (a xor b);
    layer4_outputs(379) <= a xor b;
    layer4_outputs(380) <= a;
    layer4_outputs(381) <= not a;
    layer4_outputs(382) <= not a;
    layer4_outputs(383) <= not (a or b);
    layer4_outputs(384) <= b and not a;
    layer4_outputs(385) <= not (a or b);
    layer4_outputs(386) <= a;
    layer4_outputs(387) <= not a;
    layer4_outputs(388) <= a and b;
    layer4_outputs(389) <= a or b;
    layer4_outputs(390) <= b;
    layer4_outputs(391) <= not a;
    layer4_outputs(392) <= not b;
    layer4_outputs(393) <= a and b;
    layer4_outputs(394) <= a xor b;
    layer4_outputs(395) <= a;
    layer4_outputs(396) <= '1';
    layer4_outputs(397) <= not b;
    layer4_outputs(398) <= a or b;
    layer4_outputs(399) <= not (a xor b);
    layer4_outputs(400) <= not b or a;
    layer4_outputs(401) <= not (a xor b);
    layer4_outputs(402) <= '0';
    layer4_outputs(403) <= not a;
    layer4_outputs(404) <= not a or b;
    layer4_outputs(405) <= not a or b;
    layer4_outputs(406) <= b;
    layer4_outputs(407) <= not b;
    layer4_outputs(408) <= a;
    layer4_outputs(409) <= b;
    layer4_outputs(410) <= '0';
    layer4_outputs(411) <= a and b;
    layer4_outputs(412) <= a xor b;
    layer4_outputs(413) <= not a or b;
    layer4_outputs(414) <= not (a and b);
    layer4_outputs(415) <= a or b;
    layer4_outputs(416) <= '0';
    layer4_outputs(417) <= not a or b;
    layer4_outputs(418) <= not (a or b);
    layer4_outputs(419) <= not (a xor b);
    layer4_outputs(420) <= not b;
    layer4_outputs(421) <= not a;
    layer4_outputs(422) <= not b;
    layer4_outputs(423) <= b and not a;
    layer4_outputs(424) <= not (a or b);
    layer4_outputs(425) <= not a or b;
    layer4_outputs(426) <= b;
    layer4_outputs(427) <= not a;
    layer4_outputs(428) <= not a or b;
    layer4_outputs(429) <= not a;
    layer4_outputs(430) <= not (a or b);
    layer4_outputs(431) <= not (a xor b);
    layer4_outputs(432) <= a;
    layer4_outputs(433) <= a;
    layer4_outputs(434) <= a;
    layer4_outputs(435) <= not b;
    layer4_outputs(436) <= not b;
    layer4_outputs(437) <= a and not b;
    layer4_outputs(438) <= not a;
    layer4_outputs(439) <= not b;
    layer4_outputs(440) <= not (a and b);
    layer4_outputs(441) <= not b or a;
    layer4_outputs(442) <= a xor b;
    layer4_outputs(443) <= a or b;
    layer4_outputs(444) <= b;
    layer4_outputs(445) <= b;
    layer4_outputs(446) <= not (a or b);
    layer4_outputs(447) <= b;
    layer4_outputs(448) <= not a;
    layer4_outputs(449) <= not (a and b);
    layer4_outputs(450) <= a or b;
    layer4_outputs(451) <= not (a xor b);
    layer4_outputs(452) <= not a;
    layer4_outputs(453) <= b and not a;
    layer4_outputs(454) <= not a or b;
    layer4_outputs(455) <= a;
    layer4_outputs(456) <= not (a xor b);
    layer4_outputs(457) <= not (a or b);
    layer4_outputs(458) <= a xor b;
    layer4_outputs(459) <= not a;
    layer4_outputs(460) <= not (a and b);
    layer4_outputs(461) <= b and not a;
    layer4_outputs(462) <= a or b;
    layer4_outputs(463) <= not b;
    layer4_outputs(464) <= a and b;
    layer4_outputs(465) <= b;
    layer4_outputs(466) <= not a;
    layer4_outputs(467) <= b;
    layer4_outputs(468) <= a;
    layer4_outputs(469) <= not b;
    layer4_outputs(470) <= a and not b;
    layer4_outputs(471) <= not a;
    layer4_outputs(472) <= not (a xor b);
    layer4_outputs(473) <= not b;
    layer4_outputs(474) <= not (a and b);
    layer4_outputs(475) <= not a;
    layer4_outputs(476) <= a or b;
    layer4_outputs(477) <= b;
    layer4_outputs(478) <= a and not b;
    layer4_outputs(479) <= a and b;
    layer4_outputs(480) <= a;
    layer4_outputs(481) <= a and not b;
    layer4_outputs(482) <= not a;
    layer4_outputs(483) <= b and not a;
    layer4_outputs(484) <= not b;
    layer4_outputs(485) <= not a or b;
    layer4_outputs(486) <= a;
    layer4_outputs(487) <= not (a xor b);
    layer4_outputs(488) <= a;
    layer4_outputs(489) <= b;
    layer4_outputs(490) <= a or b;
    layer4_outputs(491) <= a and not b;
    layer4_outputs(492) <= not (a xor b);
    layer4_outputs(493) <= not b;
    layer4_outputs(494) <= a or b;
    layer4_outputs(495) <= not (a xor b);
    layer4_outputs(496) <= a or b;
    layer4_outputs(497) <= b;
    layer4_outputs(498) <= not (a xor b);
    layer4_outputs(499) <= not a or b;
    layer4_outputs(500) <= not (a and b);
    layer4_outputs(501) <= not (a or b);
    layer4_outputs(502) <= not (a xor b);
    layer4_outputs(503) <= not b;
    layer4_outputs(504) <= b;
    layer4_outputs(505) <= b;
    layer4_outputs(506) <= not (a or b);
    layer4_outputs(507) <= not a;
    layer4_outputs(508) <= not b;
    layer4_outputs(509) <= a and not b;
    layer4_outputs(510) <= not b;
    layer4_outputs(511) <= not (a or b);
    layer4_outputs(512) <= a or b;
    layer4_outputs(513) <= b and not a;
    layer4_outputs(514) <= a or b;
    layer4_outputs(515) <= not a or b;
    layer4_outputs(516) <= not (a xor b);
    layer4_outputs(517) <= not b;
    layer4_outputs(518) <= not a or b;
    layer4_outputs(519) <= not a or b;
    layer4_outputs(520) <= not a or b;
    layer4_outputs(521) <= '0';
    layer4_outputs(522) <= not (a or b);
    layer4_outputs(523) <= a;
    layer4_outputs(524) <= b;
    layer4_outputs(525) <= not b or a;
    layer4_outputs(526) <= not a;
    layer4_outputs(527) <= a or b;
    layer4_outputs(528) <= not a or b;
    layer4_outputs(529) <= b and not a;
    layer4_outputs(530) <= a;
    layer4_outputs(531) <= '1';
    layer4_outputs(532) <= a or b;
    layer4_outputs(533) <= not b;
    layer4_outputs(534) <= a xor b;
    layer4_outputs(535) <= b;
    layer4_outputs(536) <= not a;
    layer4_outputs(537) <= not b;
    layer4_outputs(538) <= not b;
    layer4_outputs(539) <= a xor b;
    layer4_outputs(540) <= a;
    layer4_outputs(541) <= a and b;
    layer4_outputs(542) <= a and b;
    layer4_outputs(543) <= a or b;
    layer4_outputs(544) <= a;
    layer4_outputs(545) <= b and not a;
    layer4_outputs(546) <= a or b;
    layer4_outputs(547) <= a and not b;
    layer4_outputs(548) <= a and not b;
    layer4_outputs(549) <= not (a and b);
    layer4_outputs(550) <= a or b;
    layer4_outputs(551) <= not b;
    layer4_outputs(552) <= not (a and b);
    layer4_outputs(553) <= not b;
    layer4_outputs(554) <= not b or a;
    layer4_outputs(555) <= b;
    layer4_outputs(556) <= not (a and b);
    layer4_outputs(557) <= not b;
    layer4_outputs(558) <= not a;
    layer4_outputs(559) <= not b;
    layer4_outputs(560) <= not b or a;
    layer4_outputs(561) <= b;
    layer4_outputs(562) <= not (a xor b);
    layer4_outputs(563) <= not (a xor b);
    layer4_outputs(564) <= '1';
    layer4_outputs(565) <= b;
    layer4_outputs(566) <= not (a and b);
    layer4_outputs(567) <= not a or b;
    layer4_outputs(568) <= '0';
    layer4_outputs(569) <= not (a xor b);
    layer4_outputs(570) <= not (a or b);
    layer4_outputs(571) <= a and not b;
    layer4_outputs(572) <= not b;
    layer4_outputs(573) <= not (a or b);
    layer4_outputs(574) <= a or b;
    layer4_outputs(575) <= b and not a;
    layer4_outputs(576) <= b;
    layer4_outputs(577) <= a;
    layer4_outputs(578) <= a or b;
    layer4_outputs(579) <= not b;
    layer4_outputs(580) <= not (a and b);
    layer4_outputs(581) <= a or b;
    layer4_outputs(582) <= not (a and b);
    layer4_outputs(583) <= a;
    layer4_outputs(584) <= not a or b;
    layer4_outputs(585) <= not b;
    layer4_outputs(586) <= a and not b;
    layer4_outputs(587) <= not a or b;
    layer4_outputs(588) <= a and b;
    layer4_outputs(589) <= not a or b;
    layer4_outputs(590) <= b and not a;
    layer4_outputs(591) <= not a or b;
    layer4_outputs(592) <= a;
    layer4_outputs(593) <= not (a xor b);
    layer4_outputs(594) <= not a;
    layer4_outputs(595) <= not b;
    layer4_outputs(596) <= not b;
    layer4_outputs(597) <= not b or a;
    layer4_outputs(598) <= a and not b;
    layer4_outputs(599) <= a;
    layer4_outputs(600) <= not a or b;
    layer4_outputs(601) <= a xor b;
    layer4_outputs(602) <= not a or b;
    layer4_outputs(603) <= a and b;
    layer4_outputs(604) <= a or b;
    layer4_outputs(605) <= a;
    layer4_outputs(606) <= not a;
    layer4_outputs(607) <= not b;
    layer4_outputs(608) <= '1';
    layer4_outputs(609) <= a or b;
    layer4_outputs(610) <= a;
    layer4_outputs(611) <= not b or a;
    layer4_outputs(612) <= a and not b;
    layer4_outputs(613) <= not b;
    layer4_outputs(614) <= b and not a;
    layer4_outputs(615) <= a xor b;
    layer4_outputs(616) <= not (a and b);
    layer4_outputs(617) <= a;
    layer4_outputs(618) <= not a;
    layer4_outputs(619) <= a xor b;
    layer4_outputs(620) <= b;
    layer4_outputs(621) <= not a or b;
    layer4_outputs(622) <= not (a xor b);
    layer4_outputs(623) <= a or b;
    layer4_outputs(624) <= b;
    layer4_outputs(625) <= not (a xor b);
    layer4_outputs(626) <= b;
    layer4_outputs(627) <= a and not b;
    layer4_outputs(628) <= a and not b;
    layer4_outputs(629) <= a or b;
    layer4_outputs(630) <= a and not b;
    layer4_outputs(631) <= not b or a;
    layer4_outputs(632) <= a and not b;
    layer4_outputs(633) <= a xor b;
    layer4_outputs(634) <= not b;
    layer4_outputs(635) <= b and not a;
    layer4_outputs(636) <= not b;
    layer4_outputs(637) <= not (a or b);
    layer4_outputs(638) <= not (a or b);
    layer4_outputs(639) <= not (a or b);
    layer4_outputs(640) <= not a;
    layer4_outputs(641) <= a or b;
    layer4_outputs(642) <= b and not a;
    layer4_outputs(643) <= not b;
    layer4_outputs(644) <= not (a or b);
    layer4_outputs(645) <= b;
    layer4_outputs(646) <= not a or b;
    layer4_outputs(647) <= not b;
    layer4_outputs(648) <= b and not a;
    layer4_outputs(649) <= a;
    layer4_outputs(650) <= a and b;
    layer4_outputs(651) <= not (a or b);
    layer4_outputs(652) <= a and b;
    layer4_outputs(653) <= not b or a;
    layer4_outputs(654) <= not a;
    layer4_outputs(655) <= not a or b;
    layer4_outputs(656) <= not a;
    layer4_outputs(657) <= a xor b;
    layer4_outputs(658) <= a;
    layer4_outputs(659) <= b and not a;
    layer4_outputs(660) <= a xor b;
    layer4_outputs(661) <= not b;
    layer4_outputs(662) <= not b;
    layer4_outputs(663) <= not b;
    layer4_outputs(664) <= not a or b;
    layer4_outputs(665) <= not (a or b);
    layer4_outputs(666) <= a;
    layer4_outputs(667) <= not (a xor b);
    layer4_outputs(668) <= a xor b;
    layer4_outputs(669) <= '1';
    layer4_outputs(670) <= '1';
    layer4_outputs(671) <= not (a xor b);
    layer4_outputs(672) <= a and b;
    layer4_outputs(673) <= not b;
    layer4_outputs(674) <= not (a or b);
    layer4_outputs(675) <= not b;
    layer4_outputs(676) <= not a;
    layer4_outputs(677) <= not b;
    layer4_outputs(678) <= b and not a;
    layer4_outputs(679) <= not a;
    layer4_outputs(680) <= not (a xor b);
    layer4_outputs(681) <= not (a and b);
    layer4_outputs(682) <= b;
    layer4_outputs(683) <= a and b;
    layer4_outputs(684) <= a;
    layer4_outputs(685) <= not b;
    layer4_outputs(686) <= not a or b;
    layer4_outputs(687) <= a or b;
    layer4_outputs(688) <= a or b;
    layer4_outputs(689) <= not b;
    layer4_outputs(690) <= not a;
    layer4_outputs(691) <= a xor b;
    layer4_outputs(692) <= not b;
    layer4_outputs(693) <= not b or a;
    layer4_outputs(694) <= not b;
    layer4_outputs(695) <= b and not a;
    layer4_outputs(696) <= a;
    layer4_outputs(697) <= not (a xor b);
    layer4_outputs(698) <= b;
    layer4_outputs(699) <= b;
    layer4_outputs(700) <= '1';
    layer4_outputs(701) <= b and not a;
    layer4_outputs(702) <= a or b;
    layer4_outputs(703) <= a;
    layer4_outputs(704) <= a xor b;
    layer4_outputs(705) <= b;
    layer4_outputs(706) <= not (a xor b);
    layer4_outputs(707) <= a;
    layer4_outputs(708) <= b and not a;
    layer4_outputs(709) <= not a;
    layer4_outputs(710) <= a xor b;
    layer4_outputs(711) <= not (a or b);
    layer4_outputs(712) <= not a;
    layer4_outputs(713) <= not b;
    layer4_outputs(714) <= a;
    layer4_outputs(715) <= '0';
    layer4_outputs(716) <= not b or a;
    layer4_outputs(717) <= not a;
    layer4_outputs(718) <= not a;
    layer4_outputs(719) <= a and not b;
    layer4_outputs(720) <= not a;
    layer4_outputs(721) <= not a;
    layer4_outputs(722) <= a;
    layer4_outputs(723) <= b and not a;
    layer4_outputs(724) <= b;
    layer4_outputs(725) <= not b or a;
    layer4_outputs(726) <= not (a and b);
    layer4_outputs(727) <= not a;
    layer4_outputs(728) <= not a or b;
    layer4_outputs(729) <= not a;
    layer4_outputs(730) <= b;
    layer4_outputs(731) <= b;
    layer4_outputs(732) <= not (a xor b);
    layer4_outputs(733) <= b and not a;
    layer4_outputs(734) <= b;
    layer4_outputs(735) <= not (a and b);
    layer4_outputs(736) <= '0';
    layer4_outputs(737) <= not (a and b);
    layer4_outputs(738) <= not b;
    layer4_outputs(739) <= a xor b;
    layer4_outputs(740) <= a;
    layer4_outputs(741) <= '0';
    layer4_outputs(742) <= a and not b;
    layer4_outputs(743) <= not (a or b);
    layer4_outputs(744) <= not a or b;
    layer4_outputs(745) <= a or b;
    layer4_outputs(746) <= b and not a;
    layer4_outputs(747) <= '1';
    layer4_outputs(748) <= b and not a;
    layer4_outputs(749) <= not (a xor b);
    layer4_outputs(750) <= not b or a;
    layer4_outputs(751) <= not (a xor b);
    layer4_outputs(752) <= not a;
    layer4_outputs(753) <= not a or b;
    layer4_outputs(754) <= not b;
    layer4_outputs(755) <= a and b;
    layer4_outputs(756) <= b;
    layer4_outputs(757) <= a or b;
    layer4_outputs(758) <= not (a and b);
    layer4_outputs(759) <= not b;
    layer4_outputs(760) <= '0';
    layer4_outputs(761) <= not (a and b);
    layer4_outputs(762) <= not (a xor b);
    layer4_outputs(763) <= b;
    layer4_outputs(764) <= not b;
    layer4_outputs(765) <= not (a and b);
    layer4_outputs(766) <= b;
    layer4_outputs(767) <= a or b;
    layer4_outputs(768) <= not b or a;
    layer4_outputs(769) <= not a;
    layer4_outputs(770) <= a or b;
    layer4_outputs(771) <= a or b;
    layer4_outputs(772) <= not a;
    layer4_outputs(773) <= '1';
    layer4_outputs(774) <= not (a and b);
    layer4_outputs(775) <= a and not b;
    layer4_outputs(776) <= not b or a;
    layer4_outputs(777) <= not a;
    layer4_outputs(778) <= not (a or b);
    layer4_outputs(779) <= not b;
    layer4_outputs(780) <= b;
    layer4_outputs(781) <= not b;
    layer4_outputs(782) <= not a;
    layer4_outputs(783) <= a and b;
    layer4_outputs(784) <= not (a or b);
    layer4_outputs(785) <= b;
    layer4_outputs(786) <= a or b;
    layer4_outputs(787) <= a and not b;
    layer4_outputs(788) <= not (a and b);
    layer4_outputs(789) <= a and b;
    layer4_outputs(790) <= a xor b;
    layer4_outputs(791) <= not b;
    layer4_outputs(792) <= a;
    layer4_outputs(793) <= a;
    layer4_outputs(794) <= a or b;
    layer4_outputs(795) <= '1';
    layer4_outputs(796) <= not (a or b);
    layer4_outputs(797) <= b;
    layer4_outputs(798) <= '0';
    layer4_outputs(799) <= not (a and b);
    layer4_outputs(800) <= not a;
    layer4_outputs(801) <= not a;
    layer4_outputs(802) <= a;
    layer4_outputs(803) <= not a or b;
    layer4_outputs(804) <= a and b;
    layer4_outputs(805) <= not a or b;
    layer4_outputs(806) <= '1';
    layer4_outputs(807) <= not (a xor b);
    layer4_outputs(808) <= a and b;
    layer4_outputs(809) <= not a;
    layer4_outputs(810) <= not a;
    layer4_outputs(811) <= not a or b;
    layer4_outputs(812) <= not b;
    layer4_outputs(813) <= not b or a;
    layer4_outputs(814) <= a and not b;
    layer4_outputs(815) <= a xor b;
    layer4_outputs(816) <= not (a and b);
    layer4_outputs(817) <= not a;
    layer4_outputs(818) <= b and not a;
    layer4_outputs(819) <= a xor b;
    layer4_outputs(820) <= a and not b;
    layer4_outputs(821) <= not a;
    layer4_outputs(822) <= not (a and b);
    layer4_outputs(823) <= a or b;
    layer4_outputs(824) <= not a;
    layer4_outputs(825) <= a and b;
    layer4_outputs(826) <= b;
    layer4_outputs(827) <= a and b;
    layer4_outputs(828) <= a and not b;
    layer4_outputs(829) <= a or b;
    layer4_outputs(830) <= a and not b;
    layer4_outputs(831) <= not a;
    layer4_outputs(832) <= b;
    layer4_outputs(833) <= not a or b;
    layer4_outputs(834) <= not b;
    layer4_outputs(835) <= not (a and b);
    layer4_outputs(836) <= not b or a;
    layer4_outputs(837) <= not b;
    layer4_outputs(838) <= b;
    layer4_outputs(839) <= not a;
    layer4_outputs(840) <= not b;
    layer4_outputs(841) <= a and not b;
    layer4_outputs(842) <= a and b;
    layer4_outputs(843) <= not (a or b);
    layer4_outputs(844) <= a xor b;
    layer4_outputs(845) <= not b;
    layer4_outputs(846) <= a;
    layer4_outputs(847) <= not (a and b);
    layer4_outputs(848) <= a and b;
    layer4_outputs(849) <= a and not b;
    layer4_outputs(850) <= not (a or b);
    layer4_outputs(851) <= not a or b;
    layer4_outputs(852) <= not (a and b);
    layer4_outputs(853) <= b;
    layer4_outputs(854) <= not (a and b);
    layer4_outputs(855) <= a;
    layer4_outputs(856) <= not a;
    layer4_outputs(857) <= not (a xor b);
    layer4_outputs(858) <= not b or a;
    layer4_outputs(859) <= not a or b;
    layer4_outputs(860) <= not (a xor b);
    layer4_outputs(861) <= a;
    layer4_outputs(862) <= b;
    layer4_outputs(863) <= not a or b;
    layer4_outputs(864) <= a and b;
    layer4_outputs(865) <= a;
    layer4_outputs(866) <= b;
    layer4_outputs(867) <= not (a xor b);
    layer4_outputs(868) <= not a;
    layer4_outputs(869) <= not a;
    layer4_outputs(870) <= not a;
    layer4_outputs(871) <= not a;
    layer4_outputs(872) <= b;
    layer4_outputs(873) <= a;
    layer4_outputs(874) <= a;
    layer4_outputs(875) <= not a;
    layer4_outputs(876) <= not (a or b);
    layer4_outputs(877) <= b;
    layer4_outputs(878) <= not a;
    layer4_outputs(879) <= not b;
    layer4_outputs(880) <= a;
    layer4_outputs(881) <= a and b;
    layer4_outputs(882) <= a;
    layer4_outputs(883) <= not a;
    layer4_outputs(884) <= not a;
    layer4_outputs(885) <= not (a and b);
    layer4_outputs(886) <= not (a and b);
    layer4_outputs(887) <= a and b;
    layer4_outputs(888) <= not (a and b);
    layer4_outputs(889) <= a and b;
    layer4_outputs(890) <= a and b;
    layer4_outputs(891) <= a and not b;
    layer4_outputs(892) <= b and not a;
    layer4_outputs(893) <= not b;
    layer4_outputs(894) <= a and b;
    layer4_outputs(895) <= not (a and b);
    layer4_outputs(896) <= not a or b;
    layer4_outputs(897) <= not b;
    layer4_outputs(898) <= b;
    layer4_outputs(899) <= not b or a;
    layer4_outputs(900) <= a and b;
    layer4_outputs(901) <= b and not a;
    layer4_outputs(902) <= b and not a;
    layer4_outputs(903) <= b;
    layer4_outputs(904) <= not b;
    layer4_outputs(905) <= not b;
    layer4_outputs(906) <= '0';
    layer4_outputs(907) <= a and not b;
    layer4_outputs(908) <= b and not a;
    layer4_outputs(909) <= a or b;
    layer4_outputs(910) <= not (a or b);
    layer4_outputs(911) <= b;
    layer4_outputs(912) <= b;
    layer4_outputs(913) <= b;
    layer4_outputs(914) <= b;
    layer4_outputs(915) <= not (a and b);
    layer4_outputs(916) <= not (a xor b);
    layer4_outputs(917) <= not a;
    layer4_outputs(918) <= a;
    layer4_outputs(919) <= a xor b;
    layer4_outputs(920) <= not b or a;
    layer4_outputs(921) <= a and b;
    layer4_outputs(922) <= '1';
    layer4_outputs(923) <= a;
    layer4_outputs(924) <= not a;
    layer4_outputs(925) <= a xor b;
    layer4_outputs(926) <= not b;
    layer4_outputs(927) <= not a;
    layer4_outputs(928) <= a;
    layer4_outputs(929) <= '0';
    layer4_outputs(930) <= a and b;
    layer4_outputs(931) <= a;
    layer4_outputs(932) <= not (a or b);
    layer4_outputs(933) <= a;
    layer4_outputs(934) <= a and b;
    layer4_outputs(935) <= a and not b;
    layer4_outputs(936) <= b and not a;
    layer4_outputs(937) <= a and not b;
    layer4_outputs(938) <= '0';
    layer4_outputs(939) <= a and not b;
    layer4_outputs(940) <= not a;
    layer4_outputs(941) <= a;
    layer4_outputs(942) <= not b;
    layer4_outputs(943) <= not b;
    layer4_outputs(944) <= a and not b;
    layer4_outputs(945) <= not a or b;
    layer4_outputs(946) <= b and not a;
    layer4_outputs(947) <= a;
    layer4_outputs(948) <= not b;
    layer4_outputs(949) <= a;
    layer4_outputs(950) <= not a or b;
    layer4_outputs(951) <= a and not b;
    layer4_outputs(952) <= a;
    layer4_outputs(953) <= not a or b;
    layer4_outputs(954) <= not b;
    layer4_outputs(955) <= not b or a;
    layer4_outputs(956) <= not (a and b);
    layer4_outputs(957) <= b;
    layer4_outputs(958) <= b and not a;
    layer4_outputs(959) <= not b;
    layer4_outputs(960) <= a and not b;
    layer4_outputs(961) <= not a;
    layer4_outputs(962) <= a and b;
    layer4_outputs(963) <= not (a or b);
    layer4_outputs(964) <= not (a and b);
    layer4_outputs(965) <= not a or b;
    layer4_outputs(966) <= not a or b;
    layer4_outputs(967) <= '0';
    layer4_outputs(968) <= b;
    layer4_outputs(969) <= not (a and b);
    layer4_outputs(970) <= not (a xor b);
    layer4_outputs(971) <= not a;
    layer4_outputs(972) <= not a or b;
    layer4_outputs(973) <= b;
    layer4_outputs(974) <= not (a or b);
    layer4_outputs(975) <= not (a and b);
    layer4_outputs(976) <= a;
    layer4_outputs(977) <= not (a and b);
    layer4_outputs(978) <= not a;
    layer4_outputs(979) <= b and not a;
    layer4_outputs(980) <= b;
    layer4_outputs(981) <= a or b;
    layer4_outputs(982) <= not a;
    layer4_outputs(983) <= not a;
    layer4_outputs(984) <= a;
    layer4_outputs(985) <= not b;
    layer4_outputs(986) <= a and not b;
    layer4_outputs(987) <= a;
    layer4_outputs(988) <= a and b;
    layer4_outputs(989) <= not a or b;
    layer4_outputs(990) <= a;
    layer4_outputs(991) <= b and not a;
    layer4_outputs(992) <= b;
    layer4_outputs(993) <= b;
    layer4_outputs(994) <= not (a or b);
    layer4_outputs(995) <= not a or b;
    layer4_outputs(996) <= '1';
    layer4_outputs(997) <= a or b;
    layer4_outputs(998) <= not b;
    layer4_outputs(999) <= not b;
    layer4_outputs(1000) <= not (a or b);
    layer4_outputs(1001) <= not (a xor b);
    layer4_outputs(1002) <= b and not a;
    layer4_outputs(1003) <= not (a xor b);
    layer4_outputs(1004) <= a;
    layer4_outputs(1005) <= not b or a;
    layer4_outputs(1006) <= a;
    layer4_outputs(1007) <= a;
    layer4_outputs(1008) <= b;
    layer4_outputs(1009) <= a or b;
    layer4_outputs(1010) <= not a or b;
    layer4_outputs(1011) <= not b or a;
    layer4_outputs(1012) <= not b or a;
    layer4_outputs(1013) <= not b or a;
    layer4_outputs(1014) <= not a;
    layer4_outputs(1015) <= not a;
    layer4_outputs(1016) <= a or b;
    layer4_outputs(1017) <= not a or b;
    layer4_outputs(1018) <= b and not a;
    layer4_outputs(1019) <= not a or b;
    layer4_outputs(1020) <= not b;
    layer4_outputs(1021) <= b;
    layer4_outputs(1022) <= not a;
    layer4_outputs(1023) <= b;
    layer4_outputs(1024) <= a;
    layer4_outputs(1025) <= a or b;
    layer4_outputs(1026) <= not (a xor b);
    layer4_outputs(1027) <= a and not b;
    layer4_outputs(1028) <= a xor b;
    layer4_outputs(1029) <= b and not a;
    layer4_outputs(1030) <= a;
    layer4_outputs(1031) <= a and b;
    layer4_outputs(1032) <= a and b;
    layer4_outputs(1033) <= '0';
    layer4_outputs(1034) <= not (a xor b);
    layer4_outputs(1035) <= a xor b;
    layer4_outputs(1036) <= not b or a;
    layer4_outputs(1037) <= '0';
    layer4_outputs(1038) <= b and not a;
    layer4_outputs(1039) <= not b;
    layer4_outputs(1040) <= b;
    layer4_outputs(1041) <= not a;
    layer4_outputs(1042) <= a;
    layer4_outputs(1043) <= a;
    layer4_outputs(1044) <= not a or b;
    layer4_outputs(1045) <= not a;
    layer4_outputs(1046) <= not b or a;
    layer4_outputs(1047) <= b;
    layer4_outputs(1048) <= '1';
    layer4_outputs(1049) <= b;
    layer4_outputs(1050) <= not a;
    layer4_outputs(1051) <= not (a xor b);
    layer4_outputs(1052) <= '0';
    layer4_outputs(1053) <= a and not b;
    layer4_outputs(1054) <= '1';
    layer4_outputs(1055) <= not (a and b);
    layer4_outputs(1056) <= a;
    layer4_outputs(1057) <= not (a or b);
    layer4_outputs(1058) <= not (a xor b);
    layer4_outputs(1059) <= not (a xor b);
    layer4_outputs(1060) <= a;
    layer4_outputs(1061) <= b;
    layer4_outputs(1062) <= a;
    layer4_outputs(1063) <= not (a xor b);
    layer4_outputs(1064) <= a and b;
    layer4_outputs(1065) <= a;
    layer4_outputs(1066) <= b and not a;
    layer4_outputs(1067) <= not (a xor b);
    layer4_outputs(1068) <= not b or a;
    layer4_outputs(1069) <= b;
    layer4_outputs(1070) <= not b or a;
    layer4_outputs(1071) <= not (a or b);
    layer4_outputs(1072) <= b;
    layer4_outputs(1073) <= not b or a;
    layer4_outputs(1074) <= b;
    layer4_outputs(1075) <= b;
    layer4_outputs(1076) <= a and b;
    layer4_outputs(1077) <= not (a and b);
    layer4_outputs(1078) <= not b or a;
    layer4_outputs(1079) <= not (a xor b);
    layer4_outputs(1080) <= a or b;
    layer4_outputs(1081) <= '1';
    layer4_outputs(1082) <= '1';
    layer4_outputs(1083) <= a;
    layer4_outputs(1084) <= b;
    layer4_outputs(1085) <= not a or b;
    layer4_outputs(1086) <= not a;
    layer4_outputs(1087) <= not a;
    layer4_outputs(1088) <= not (a and b);
    layer4_outputs(1089) <= b;
    layer4_outputs(1090) <= not b;
    layer4_outputs(1091) <= not (a and b);
    layer4_outputs(1092) <= a or b;
    layer4_outputs(1093) <= a and b;
    layer4_outputs(1094) <= not b or a;
    layer4_outputs(1095) <= a xor b;
    layer4_outputs(1096) <= not a;
    layer4_outputs(1097) <= not a or b;
    layer4_outputs(1098) <= a and b;
    layer4_outputs(1099) <= not a;
    layer4_outputs(1100) <= '1';
    layer4_outputs(1101) <= not b;
    layer4_outputs(1102) <= b;
    layer4_outputs(1103) <= not b or a;
    layer4_outputs(1104) <= not b or a;
    layer4_outputs(1105) <= not (a or b);
    layer4_outputs(1106) <= not (a or b);
    layer4_outputs(1107) <= b;
    layer4_outputs(1108) <= '1';
    layer4_outputs(1109) <= not b;
    layer4_outputs(1110) <= a;
    layer4_outputs(1111) <= a;
    layer4_outputs(1112) <= not (a or b);
    layer4_outputs(1113) <= a;
    layer4_outputs(1114) <= not b;
    layer4_outputs(1115) <= not b or a;
    layer4_outputs(1116) <= not a;
    layer4_outputs(1117) <= not a or b;
    layer4_outputs(1118) <= '1';
    layer4_outputs(1119) <= not b or a;
    layer4_outputs(1120) <= a;
    layer4_outputs(1121) <= not (a or b);
    layer4_outputs(1122) <= a;
    layer4_outputs(1123) <= b;
    layer4_outputs(1124) <= a xor b;
    layer4_outputs(1125) <= b;
    layer4_outputs(1126) <= not (a xor b);
    layer4_outputs(1127) <= not (a or b);
    layer4_outputs(1128) <= b and not a;
    layer4_outputs(1129) <= not a;
    layer4_outputs(1130) <= b;
    layer4_outputs(1131) <= not b;
    layer4_outputs(1132) <= not (a xor b);
    layer4_outputs(1133) <= b and not a;
    layer4_outputs(1134) <= a or b;
    layer4_outputs(1135) <= a and not b;
    layer4_outputs(1136) <= not (a and b);
    layer4_outputs(1137) <= a xor b;
    layer4_outputs(1138) <= not b;
    layer4_outputs(1139) <= not b or a;
    layer4_outputs(1140) <= a;
    layer4_outputs(1141) <= b and not a;
    layer4_outputs(1142) <= a and not b;
    layer4_outputs(1143) <= not (a and b);
    layer4_outputs(1144) <= not b;
    layer4_outputs(1145) <= a;
    layer4_outputs(1146) <= b;
    layer4_outputs(1147) <= not (a or b);
    layer4_outputs(1148) <= b;
    layer4_outputs(1149) <= b and not a;
    layer4_outputs(1150) <= a and b;
    layer4_outputs(1151) <= not b;
    layer4_outputs(1152) <= not b;
    layer4_outputs(1153) <= not b;
    layer4_outputs(1154) <= a;
    layer4_outputs(1155) <= a or b;
    layer4_outputs(1156) <= not b or a;
    layer4_outputs(1157) <= not b;
    layer4_outputs(1158) <= a or b;
    layer4_outputs(1159) <= a;
    layer4_outputs(1160) <= a xor b;
    layer4_outputs(1161) <= not b;
    layer4_outputs(1162) <= not (a or b);
    layer4_outputs(1163) <= a;
    layer4_outputs(1164) <= not (a or b);
    layer4_outputs(1165) <= not (a xor b);
    layer4_outputs(1166) <= a xor b;
    layer4_outputs(1167) <= not (a xor b);
    layer4_outputs(1168) <= '1';
    layer4_outputs(1169) <= not b;
    layer4_outputs(1170) <= a and b;
    layer4_outputs(1171) <= a;
    layer4_outputs(1172) <= not b or a;
    layer4_outputs(1173) <= a and not b;
    layer4_outputs(1174) <= a and not b;
    layer4_outputs(1175) <= a and not b;
    layer4_outputs(1176) <= not (a and b);
    layer4_outputs(1177) <= not (a xor b);
    layer4_outputs(1178) <= not b;
    layer4_outputs(1179) <= not b;
    layer4_outputs(1180) <= not (a and b);
    layer4_outputs(1181) <= not b;
    layer4_outputs(1182) <= not b or a;
    layer4_outputs(1183) <= not (a xor b);
    layer4_outputs(1184) <= not b;
    layer4_outputs(1185) <= not b or a;
    layer4_outputs(1186) <= a xor b;
    layer4_outputs(1187) <= b;
    layer4_outputs(1188) <= not a;
    layer4_outputs(1189) <= a or b;
    layer4_outputs(1190) <= not b;
    layer4_outputs(1191) <= not (a and b);
    layer4_outputs(1192) <= a and b;
    layer4_outputs(1193) <= a;
    layer4_outputs(1194) <= not a;
    layer4_outputs(1195) <= a;
    layer4_outputs(1196) <= a;
    layer4_outputs(1197) <= b;
    layer4_outputs(1198) <= not a or b;
    layer4_outputs(1199) <= not (a and b);
    layer4_outputs(1200) <= a;
    layer4_outputs(1201) <= a and b;
    layer4_outputs(1202) <= not b;
    layer4_outputs(1203) <= a;
    layer4_outputs(1204) <= b;
    layer4_outputs(1205) <= not a;
    layer4_outputs(1206) <= a or b;
    layer4_outputs(1207) <= b;
    layer4_outputs(1208) <= b;
    layer4_outputs(1209) <= a or b;
    layer4_outputs(1210) <= not a or b;
    layer4_outputs(1211) <= a and not b;
    layer4_outputs(1212) <= b;
    layer4_outputs(1213) <= not b;
    layer4_outputs(1214) <= not a;
    layer4_outputs(1215) <= not a;
    layer4_outputs(1216) <= not a;
    layer4_outputs(1217) <= a and b;
    layer4_outputs(1218) <= not a;
    layer4_outputs(1219) <= a xor b;
    layer4_outputs(1220) <= not b;
    layer4_outputs(1221) <= b and not a;
    layer4_outputs(1222) <= b and not a;
    layer4_outputs(1223) <= a and not b;
    layer4_outputs(1224) <= not (a or b);
    layer4_outputs(1225) <= not b or a;
    layer4_outputs(1226) <= b;
    layer4_outputs(1227) <= not a;
    layer4_outputs(1228) <= not a;
    layer4_outputs(1229) <= a xor b;
    layer4_outputs(1230) <= not b;
    layer4_outputs(1231) <= not (a and b);
    layer4_outputs(1232) <= not a;
    layer4_outputs(1233) <= a and not b;
    layer4_outputs(1234) <= b;
    layer4_outputs(1235) <= b;
    layer4_outputs(1236) <= b;
    layer4_outputs(1237) <= not b;
    layer4_outputs(1238) <= not a or b;
    layer4_outputs(1239) <= a and not b;
    layer4_outputs(1240) <= a and not b;
    layer4_outputs(1241) <= a or b;
    layer4_outputs(1242) <= not (a xor b);
    layer4_outputs(1243) <= not (a and b);
    layer4_outputs(1244) <= a xor b;
    layer4_outputs(1245) <= not (a or b);
    layer4_outputs(1246) <= not a or b;
    layer4_outputs(1247) <= not b;
    layer4_outputs(1248) <= not (a and b);
    layer4_outputs(1249) <= not (a xor b);
    layer4_outputs(1250) <= b;
    layer4_outputs(1251) <= not a or b;
    layer4_outputs(1252) <= not b or a;
    layer4_outputs(1253) <= b;
    layer4_outputs(1254) <= not a;
    layer4_outputs(1255) <= b;
    layer4_outputs(1256) <= not a;
    layer4_outputs(1257) <= a;
    layer4_outputs(1258) <= not a or b;
    layer4_outputs(1259) <= not a;
    layer4_outputs(1260) <= b;
    layer4_outputs(1261) <= b;
    layer4_outputs(1262) <= a;
    layer4_outputs(1263) <= a and b;
    layer4_outputs(1264) <= not b;
    layer4_outputs(1265) <= not (a and b);
    layer4_outputs(1266) <= not b;
    layer4_outputs(1267) <= a and not b;
    layer4_outputs(1268) <= a and b;
    layer4_outputs(1269) <= b and not a;
    layer4_outputs(1270) <= not a;
    layer4_outputs(1271) <= not b;
    layer4_outputs(1272) <= a xor b;
    layer4_outputs(1273) <= a and not b;
    layer4_outputs(1274) <= b;
    layer4_outputs(1275) <= not a;
    layer4_outputs(1276) <= a;
    layer4_outputs(1277) <= not b;
    layer4_outputs(1278) <= a or b;
    layer4_outputs(1279) <= not b;
    layer4_outputs(1280) <= a;
    layer4_outputs(1281) <= not (a xor b);
    layer4_outputs(1282) <= not (a xor b);
    layer4_outputs(1283) <= b;
    layer4_outputs(1284) <= not a or b;
    layer4_outputs(1285) <= not (a xor b);
    layer4_outputs(1286) <= not b;
    layer4_outputs(1287) <= not a;
    layer4_outputs(1288) <= not b;
    layer4_outputs(1289) <= not b or a;
    layer4_outputs(1290) <= b and not a;
    layer4_outputs(1291) <= not a;
    layer4_outputs(1292) <= b;
    layer4_outputs(1293) <= not a;
    layer4_outputs(1294) <= not (a xor b);
    layer4_outputs(1295) <= a;
    layer4_outputs(1296) <= not a;
    layer4_outputs(1297) <= a and b;
    layer4_outputs(1298) <= not b;
    layer4_outputs(1299) <= a or b;
    layer4_outputs(1300) <= not a or b;
    layer4_outputs(1301) <= not a;
    layer4_outputs(1302) <= b and not a;
    layer4_outputs(1303) <= not a or b;
    layer4_outputs(1304) <= not b;
    layer4_outputs(1305) <= not (a xor b);
    layer4_outputs(1306) <= not (a or b);
    layer4_outputs(1307) <= a and not b;
    layer4_outputs(1308) <= b;
    layer4_outputs(1309) <= '1';
    layer4_outputs(1310) <= a and not b;
    layer4_outputs(1311) <= a xor b;
    layer4_outputs(1312) <= '1';
    layer4_outputs(1313) <= a or b;
    layer4_outputs(1314) <= a;
    layer4_outputs(1315) <= a and b;
    layer4_outputs(1316) <= not a or b;
    layer4_outputs(1317) <= a;
    layer4_outputs(1318) <= not (a and b);
    layer4_outputs(1319) <= a xor b;
    layer4_outputs(1320) <= not a;
    layer4_outputs(1321) <= not (a or b);
    layer4_outputs(1322) <= a xor b;
    layer4_outputs(1323) <= b and not a;
    layer4_outputs(1324) <= not b;
    layer4_outputs(1325) <= not a or b;
    layer4_outputs(1326) <= a and b;
    layer4_outputs(1327) <= not b or a;
    layer4_outputs(1328) <= a;
    layer4_outputs(1329) <= not a;
    layer4_outputs(1330) <= a and b;
    layer4_outputs(1331) <= a and not b;
    layer4_outputs(1332) <= a and b;
    layer4_outputs(1333) <= not a or b;
    layer4_outputs(1334) <= a and not b;
    layer4_outputs(1335) <= not b or a;
    layer4_outputs(1336) <= not (a and b);
    layer4_outputs(1337) <= b and not a;
    layer4_outputs(1338) <= a;
    layer4_outputs(1339) <= not b;
    layer4_outputs(1340) <= b;
    layer4_outputs(1341) <= not a;
    layer4_outputs(1342) <= not a;
    layer4_outputs(1343) <= not (a or b);
    layer4_outputs(1344) <= b;
    layer4_outputs(1345) <= not b;
    layer4_outputs(1346) <= b and not a;
    layer4_outputs(1347) <= a or b;
    layer4_outputs(1348) <= not a;
    layer4_outputs(1349) <= a or b;
    layer4_outputs(1350) <= not b or a;
    layer4_outputs(1351) <= not a;
    layer4_outputs(1352) <= not (a and b);
    layer4_outputs(1353) <= not b;
    layer4_outputs(1354) <= a;
    layer4_outputs(1355) <= b;
    layer4_outputs(1356) <= a xor b;
    layer4_outputs(1357) <= a xor b;
    layer4_outputs(1358) <= a and b;
    layer4_outputs(1359) <= not (a and b);
    layer4_outputs(1360) <= b;
    layer4_outputs(1361) <= a;
    layer4_outputs(1362) <= a xor b;
    layer4_outputs(1363) <= a and not b;
    layer4_outputs(1364) <= a;
    layer4_outputs(1365) <= not a or b;
    layer4_outputs(1366) <= a and b;
    layer4_outputs(1367) <= a or b;
    layer4_outputs(1368) <= a and not b;
    layer4_outputs(1369) <= a;
    layer4_outputs(1370) <= not b;
    layer4_outputs(1371) <= not (a xor b);
    layer4_outputs(1372) <= b;
    layer4_outputs(1373) <= b;
    layer4_outputs(1374) <= not b;
    layer4_outputs(1375) <= a;
    layer4_outputs(1376) <= b;
    layer4_outputs(1377) <= a and b;
    layer4_outputs(1378) <= a and not b;
    layer4_outputs(1379) <= not a;
    layer4_outputs(1380) <= b;
    layer4_outputs(1381) <= not (a and b);
    layer4_outputs(1382) <= not a or b;
    layer4_outputs(1383) <= not b;
    layer4_outputs(1384) <= not b;
    layer4_outputs(1385) <= not a;
    layer4_outputs(1386) <= a and not b;
    layer4_outputs(1387) <= not b;
    layer4_outputs(1388) <= a xor b;
    layer4_outputs(1389) <= not b or a;
    layer4_outputs(1390) <= a and b;
    layer4_outputs(1391) <= not b or a;
    layer4_outputs(1392) <= a and not b;
    layer4_outputs(1393) <= not b;
    layer4_outputs(1394) <= a;
    layer4_outputs(1395) <= a;
    layer4_outputs(1396) <= b;
    layer4_outputs(1397) <= not (a xor b);
    layer4_outputs(1398) <= not (a xor b);
    layer4_outputs(1399) <= not a;
    layer4_outputs(1400) <= not a;
    layer4_outputs(1401) <= a;
    layer4_outputs(1402) <= a and b;
    layer4_outputs(1403) <= not a;
    layer4_outputs(1404) <= b and not a;
    layer4_outputs(1405) <= b;
    layer4_outputs(1406) <= a and not b;
    layer4_outputs(1407) <= not a;
    layer4_outputs(1408) <= a;
    layer4_outputs(1409) <= not b;
    layer4_outputs(1410) <= b;
    layer4_outputs(1411) <= a or b;
    layer4_outputs(1412) <= not a or b;
    layer4_outputs(1413) <= b;
    layer4_outputs(1414) <= not b;
    layer4_outputs(1415) <= b;
    layer4_outputs(1416) <= a and b;
    layer4_outputs(1417) <= a;
    layer4_outputs(1418) <= not a;
    layer4_outputs(1419) <= not (a or b);
    layer4_outputs(1420) <= not b;
    layer4_outputs(1421) <= b;
    layer4_outputs(1422) <= a and b;
    layer4_outputs(1423) <= not (a or b);
    layer4_outputs(1424) <= not a;
    layer4_outputs(1425) <= a xor b;
    layer4_outputs(1426) <= a or b;
    layer4_outputs(1427) <= not a or b;
    layer4_outputs(1428) <= a and not b;
    layer4_outputs(1429) <= not a;
    layer4_outputs(1430) <= not b;
    layer4_outputs(1431) <= a and not b;
    layer4_outputs(1432) <= b;
    layer4_outputs(1433) <= a and not b;
    layer4_outputs(1434) <= b;
    layer4_outputs(1435) <= not b or a;
    layer4_outputs(1436) <= not (a xor b);
    layer4_outputs(1437) <= not a or b;
    layer4_outputs(1438) <= a or b;
    layer4_outputs(1439) <= '0';
    layer4_outputs(1440) <= not b;
    layer4_outputs(1441) <= a or b;
    layer4_outputs(1442) <= not (a xor b);
    layer4_outputs(1443) <= not b or a;
    layer4_outputs(1444) <= a and b;
    layer4_outputs(1445) <= a or b;
    layer4_outputs(1446) <= not (a xor b);
    layer4_outputs(1447) <= not (a xor b);
    layer4_outputs(1448) <= not (a and b);
    layer4_outputs(1449) <= not b;
    layer4_outputs(1450) <= a or b;
    layer4_outputs(1451) <= not a;
    layer4_outputs(1452) <= a or b;
    layer4_outputs(1453) <= not a;
    layer4_outputs(1454) <= not b or a;
    layer4_outputs(1455) <= not b;
    layer4_outputs(1456) <= not (a xor b);
    layer4_outputs(1457) <= not b or a;
    layer4_outputs(1458) <= not b;
    layer4_outputs(1459) <= not a or b;
    layer4_outputs(1460) <= '0';
    layer4_outputs(1461) <= not (a and b);
    layer4_outputs(1462) <= not (a or b);
    layer4_outputs(1463) <= a or b;
    layer4_outputs(1464) <= a or b;
    layer4_outputs(1465) <= a;
    layer4_outputs(1466) <= not (a or b);
    layer4_outputs(1467) <= a and b;
    layer4_outputs(1468) <= not (a and b);
    layer4_outputs(1469) <= not (a xor b);
    layer4_outputs(1470) <= not a;
    layer4_outputs(1471) <= a and b;
    layer4_outputs(1472) <= not b or a;
    layer4_outputs(1473) <= a;
    layer4_outputs(1474) <= not (a xor b);
    layer4_outputs(1475) <= a xor b;
    layer4_outputs(1476) <= a and b;
    layer4_outputs(1477) <= not (a xor b);
    layer4_outputs(1478) <= not a;
    layer4_outputs(1479) <= a and b;
    layer4_outputs(1480) <= a xor b;
    layer4_outputs(1481) <= b;
    layer4_outputs(1482) <= not (a or b);
    layer4_outputs(1483) <= b;
    layer4_outputs(1484) <= not (a xor b);
    layer4_outputs(1485) <= b;
    layer4_outputs(1486) <= a;
    layer4_outputs(1487) <= a and b;
    layer4_outputs(1488) <= not a or b;
    layer4_outputs(1489) <= a and not b;
    layer4_outputs(1490) <= not a;
    layer4_outputs(1491) <= not (a and b);
    layer4_outputs(1492) <= not (a and b);
    layer4_outputs(1493) <= not a or b;
    layer4_outputs(1494) <= not b;
    layer4_outputs(1495) <= a;
    layer4_outputs(1496) <= not (a or b);
    layer4_outputs(1497) <= a;
    layer4_outputs(1498) <= not a or b;
    layer4_outputs(1499) <= not b;
    layer4_outputs(1500) <= not b or a;
    layer4_outputs(1501) <= a xor b;
    layer4_outputs(1502) <= not b or a;
    layer4_outputs(1503) <= not (a or b);
    layer4_outputs(1504) <= b and not a;
    layer4_outputs(1505) <= not a or b;
    layer4_outputs(1506) <= not b or a;
    layer4_outputs(1507) <= not (a and b);
    layer4_outputs(1508) <= not b;
    layer4_outputs(1509) <= a;
    layer4_outputs(1510) <= not b or a;
    layer4_outputs(1511) <= not (a and b);
    layer4_outputs(1512) <= not a;
    layer4_outputs(1513) <= not a;
    layer4_outputs(1514) <= a xor b;
    layer4_outputs(1515) <= a and not b;
    layer4_outputs(1516) <= not (a xor b);
    layer4_outputs(1517) <= '1';
    layer4_outputs(1518) <= a xor b;
    layer4_outputs(1519) <= not b;
    layer4_outputs(1520) <= b and not a;
    layer4_outputs(1521) <= a xor b;
    layer4_outputs(1522) <= not b or a;
    layer4_outputs(1523) <= not (a xor b);
    layer4_outputs(1524) <= not b;
    layer4_outputs(1525) <= b;
    layer4_outputs(1526) <= a;
    layer4_outputs(1527) <= not (a and b);
    layer4_outputs(1528) <= not (a and b);
    layer4_outputs(1529) <= not (a xor b);
    layer4_outputs(1530) <= not (a or b);
    layer4_outputs(1531) <= not a;
    layer4_outputs(1532) <= b and not a;
    layer4_outputs(1533) <= not a or b;
    layer4_outputs(1534) <= a and not b;
    layer4_outputs(1535) <= a;
    layer4_outputs(1536) <= b and not a;
    layer4_outputs(1537) <= not (a or b);
    layer4_outputs(1538) <= not a or b;
    layer4_outputs(1539) <= not b;
    layer4_outputs(1540) <= not a;
    layer4_outputs(1541) <= not (a xor b);
    layer4_outputs(1542) <= a;
    layer4_outputs(1543) <= not b;
    layer4_outputs(1544) <= not (a xor b);
    layer4_outputs(1545) <= b;
    layer4_outputs(1546) <= not (a or b);
    layer4_outputs(1547) <= not a;
    layer4_outputs(1548) <= b and not a;
    layer4_outputs(1549) <= not a;
    layer4_outputs(1550) <= not (a xor b);
    layer4_outputs(1551) <= a;
    layer4_outputs(1552) <= a or b;
    layer4_outputs(1553) <= not (a or b);
    layer4_outputs(1554) <= '1';
    layer4_outputs(1555) <= not (a xor b);
    layer4_outputs(1556) <= not (a or b);
    layer4_outputs(1557) <= b;
    layer4_outputs(1558) <= a;
    layer4_outputs(1559) <= not a;
    layer4_outputs(1560) <= not b;
    layer4_outputs(1561) <= not b;
    layer4_outputs(1562) <= a xor b;
    layer4_outputs(1563) <= not a;
    layer4_outputs(1564) <= not a or b;
    layer4_outputs(1565) <= not (a xor b);
    layer4_outputs(1566) <= not a;
    layer4_outputs(1567) <= not (a or b);
    layer4_outputs(1568) <= a;
    layer4_outputs(1569) <= a and b;
    layer4_outputs(1570) <= b and not a;
    layer4_outputs(1571) <= b;
    layer4_outputs(1572) <= a;
    layer4_outputs(1573) <= a;
    layer4_outputs(1574) <= b;
    layer4_outputs(1575) <= not b or a;
    layer4_outputs(1576) <= a;
    layer4_outputs(1577) <= not a;
    layer4_outputs(1578) <= '1';
    layer4_outputs(1579) <= not a or b;
    layer4_outputs(1580) <= '0';
    layer4_outputs(1581) <= not a;
    layer4_outputs(1582) <= not (a and b);
    layer4_outputs(1583) <= not a;
    layer4_outputs(1584) <= a and b;
    layer4_outputs(1585) <= a;
    layer4_outputs(1586) <= not (a xor b);
    layer4_outputs(1587) <= not a or b;
    layer4_outputs(1588) <= not (a or b);
    layer4_outputs(1589) <= not (a and b);
    layer4_outputs(1590) <= a or b;
    layer4_outputs(1591) <= b;
    layer4_outputs(1592) <= not b or a;
    layer4_outputs(1593) <= '1';
    layer4_outputs(1594) <= a and b;
    layer4_outputs(1595) <= a xor b;
    layer4_outputs(1596) <= a or b;
    layer4_outputs(1597) <= a;
    layer4_outputs(1598) <= not b;
    layer4_outputs(1599) <= a xor b;
    layer4_outputs(1600) <= b;
    layer4_outputs(1601) <= not a;
    layer4_outputs(1602) <= not b;
    layer4_outputs(1603) <= b;
    layer4_outputs(1604) <= '1';
    layer4_outputs(1605) <= a;
    layer4_outputs(1606) <= b and not a;
    layer4_outputs(1607) <= b;
    layer4_outputs(1608) <= a;
    layer4_outputs(1609) <= '1';
    layer4_outputs(1610) <= not (a xor b);
    layer4_outputs(1611) <= a and b;
    layer4_outputs(1612) <= not b;
    layer4_outputs(1613) <= a and not b;
    layer4_outputs(1614) <= '1';
    layer4_outputs(1615) <= not b or a;
    layer4_outputs(1616) <= b;
    layer4_outputs(1617) <= a or b;
    layer4_outputs(1618) <= not a;
    layer4_outputs(1619) <= b and not a;
    layer4_outputs(1620) <= a or b;
    layer4_outputs(1621) <= a and not b;
    layer4_outputs(1622) <= b and not a;
    layer4_outputs(1623) <= not (a or b);
    layer4_outputs(1624) <= not b;
    layer4_outputs(1625) <= not (a or b);
    layer4_outputs(1626) <= a and not b;
    layer4_outputs(1627) <= a;
    layer4_outputs(1628) <= not b;
    layer4_outputs(1629) <= not a or b;
    layer4_outputs(1630) <= not b or a;
    layer4_outputs(1631) <= not (a or b);
    layer4_outputs(1632) <= not (a and b);
    layer4_outputs(1633) <= not (a and b);
    layer4_outputs(1634) <= not b;
    layer4_outputs(1635) <= a and b;
    layer4_outputs(1636) <= not a;
    layer4_outputs(1637) <= not b;
    layer4_outputs(1638) <= not (a and b);
    layer4_outputs(1639) <= a or b;
    layer4_outputs(1640) <= a or b;
    layer4_outputs(1641) <= b;
    layer4_outputs(1642) <= b;
    layer4_outputs(1643) <= not (a xor b);
    layer4_outputs(1644) <= b and not a;
    layer4_outputs(1645) <= not b or a;
    layer4_outputs(1646) <= b;
    layer4_outputs(1647) <= a or b;
    layer4_outputs(1648) <= not a;
    layer4_outputs(1649) <= a xor b;
    layer4_outputs(1650) <= a and not b;
    layer4_outputs(1651) <= not b;
    layer4_outputs(1652) <= a and b;
    layer4_outputs(1653) <= b;
    layer4_outputs(1654) <= not b or a;
    layer4_outputs(1655) <= a and not b;
    layer4_outputs(1656) <= b and not a;
    layer4_outputs(1657) <= b;
    layer4_outputs(1658) <= not b or a;
    layer4_outputs(1659) <= a and not b;
    layer4_outputs(1660) <= not a or b;
    layer4_outputs(1661) <= not b;
    layer4_outputs(1662) <= not b or a;
    layer4_outputs(1663) <= not b;
    layer4_outputs(1664) <= not (a or b);
    layer4_outputs(1665) <= b;
    layer4_outputs(1666) <= a or b;
    layer4_outputs(1667) <= b;
    layer4_outputs(1668) <= not (a xor b);
    layer4_outputs(1669) <= a;
    layer4_outputs(1670) <= not a or b;
    layer4_outputs(1671) <= not b;
    layer4_outputs(1672) <= not b;
    layer4_outputs(1673) <= not (a and b);
    layer4_outputs(1674) <= not (a or b);
    layer4_outputs(1675) <= not (a or b);
    layer4_outputs(1676) <= a xor b;
    layer4_outputs(1677) <= not (a or b);
    layer4_outputs(1678) <= b;
    layer4_outputs(1679) <= a;
    layer4_outputs(1680) <= not (a xor b);
    layer4_outputs(1681) <= not (a or b);
    layer4_outputs(1682) <= not (a xor b);
    layer4_outputs(1683) <= a;
    layer4_outputs(1684) <= not (a or b);
    layer4_outputs(1685) <= not b;
    layer4_outputs(1686) <= not a;
    layer4_outputs(1687) <= not (a xor b);
    layer4_outputs(1688) <= not b or a;
    layer4_outputs(1689) <= not b or a;
    layer4_outputs(1690) <= not (a and b);
    layer4_outputs(1691) <= a;
    layer4_outputs(1692) <= not (a or b);
    layer4_outputs(1693) <= a xor b;
    layer4_outputs(1694) <= a xor b;
    layer4_outputs(1695) <= not (a xor b);
    layer4_outputs(1696) <= a;
    layer4_outputs(1697) <= not a;
    layer4_outputs(1698) <= not (a and b);
    layer4_outputs(1699) <= a;
    layer4_outputs(1700) <= not b;
    layer4_outputs(1701) <= a and b;
    layer4_outputs(1702) <= a and not b;
    layer4_outputs(1703) <= b;
    layer4_outputs(1704) <= not (a or b);
    layer4_outputs(1705) <= a or b;
    layer4_outputs(1706) <= a and b;
    layer4_outputs(1707) <= not b;
    layer4_outputs(1708) <= a xor b;
    layer4_outputs(1709) <= not b or a;
    layer4_outputs(1710) <= a and not b;
    layer4_outputs(1711) <= a and b;
    layer4_outputs(1712) <= not b;
    layer4_outputs(1713) <= not (a or b);
    layer4_outputs(1714) <= not (a or b);
    layer4_outputs(1715) <= not b;
    layer4_outputs(1716) <= a or b;
    layer4_outputs(1717) <= a and not b;
    layer4_outputs(1718) <= b;
    layer4_outputs(1719) <= not (a xor b);
    layer4_outputs(1720) <= a and b;
    layer4_outputs(1721) <= not b;
    layer4_outputs(1722) <= not (a xor b);
    layer4_outputs(1723) <= a xor b;
    layer4_outputs(1724) <= not (a and b);
    layer4_outputs(1725) <= not (a xor b);
    layer4_outputs(1726) <= b;
    layer4_outputs(1727) <= a;
    layer4_outputs(1728) <= a xor b;
    layer4_outputs(1729) <= not (a xor b);
    layer4_outputs(1730) <= not a;
    layer4_outputs(1731) <= a and not b;
    layer4_outputs(1732) <= a;
    layer4_outputs(1733) <= a and b;
    layer4_outputs(1734) <= b and not a;
    layer4_outputs(1735) <= not a;
    layer4_outputs(1736) <= a;
    layer4_outputs(1737) <= not a or b;
    layer4_outputs(1738) <= a or b;
    layer4_outputs(1739) <= not (a or b);
    layer4_outputs(1740) <= not a;
    layer4_outputs(1741) <= not b;
    layer4_outputs(1742) <= not a;
    layer4_outputs(1743) <= b;
    layer4_outputs(1744) <= not b;
    layer4_outputs(1745) <= a and not b;
    layer4_outputs(1746) <= not b or a;
    layer4_outputs(1747) <= b and not a;
    layer4_outputs(1748) <= not (a or b);
    layer4_outputs(1749) <= '1';
    layer4_outputs(1750) <= not (a and b);
    layer4_outputs(1751) <= not (a and b);
    layer4_outputs(1752) <= not b;
    layer4_outputs(1753) <= b;
    layer4_outputs(1754) <= a and not b;
    layer4_outputs(1755) <= a;
    layer4_outputs(1756) <= b;
    layer4_outputs(1757) <= not a;
    layer4_outputs(1758) <= not (a and b);
    layer4_outputs(1759) <= a and not b;
    layer4_outputs(1760) <= b;
    layer4_outputs(1761) <= not (a xor b);
    layer4_outputs(1762) <= not (a and b);
    layer4_outputs(1763) <= a;
    layer4_outputs(1764) <= a;
    layer4_outputs(1765) <= a or b;
    layer4_outputs(1766) <= a and not b;
    layer4_outputs(1767) <= not b;
    layer4_outputs(1768) <= not b;
    layer4_outputs(1769) <= not (a xor b);
    layer4_outputs(1770) <= '1';
    layer4_outputs(1771) <= not (a and b);
    layer4_outputs(1772) <= not a or b;
    layer4_outputs(1773) <= b;
    layer4_outputs(1774) <= not (a xor b);
    layer4_outputs(1775) <= b;
    layer4_outputs(1776) <= not b;
    layer4_outputs(1777) <= not b;
    layer4_outputs(1778) <= b and not a;
    layer4_outputs(1779) <= not b;
    layer4_outputs(1780) <= not b;
    layer4_outputs(1781) <= not a;
    layer4_outputs(1782) <= a;
    layer4_outputs(1783) <= not b;
    layer4_outputs(1784) <= not (a and b);
    layer4_outputs(1785) <= not b;
    layer4_outputs(1786) <= not b;
    layer4_outputs(1787) <= a and b;
    layer4_outputs(1788) <= not (a xor b);
    layer4_outputs(1789) <= not (a or b);
    layer4_outputs(1790) <= a and b;
    layer4_outputs(1791) <= not b;
    layer4_outputs(1792) <= '1';
    layer4_outputs(1793) <= b;
    layer4_outputs(1794) <= not a;
    layer4_outputs(1795) <= not (a or b);
    layer4_outputs(1796) <= a xor b;
    layer4_outputs(1797) <= not b;
    layer4_outputs(1798) <= b and not a;
    layer4_outputs(1799) <= a and b;
    layer4_outputs(1800) <= a and not b;
    layer4_outputs(1801) <= not (a xor b);
    layer4_outputs(1802) <= a and b;
    layer4_outputs(1803) <= not a;
    layer4_outputs(1804) <= b and not a;
    layer4_outputs(1805) <= a and b;
    layer4_outputs(1806) <= not a;
    layer4_outputs(1807) <= a;
    layer4_outputs(1808) <= a xor b;
    layer4_outputs(1809) <= a or b;
    layer4_outputs(1810) <= not b;
    layer4_outputs(1811) <= a and b;
    layer4_outputs(1812) <= not (a and b);
    layer4_outputs(1813) <= b;
    layer4_outputs(1814) <= not a;
    layer4_outputs(1815) <= a xor b;
    layer4_outputs(1816) <= b;
    layer4_outputs(1817) <= a;
    layer4_outputs(1818) <= not (a or b);
    layer4_outputs(1819) <= not a;
    layer4_outputs(1820) <= not (a and b);
    layer4_outputs(1821) <= b;
    layer4_outputs(1822) <= b and not a;
    layer4_outputs(1823) <= not b;
    layer4_outputs(1824) <= a and b;
    layer4_outputs(1825) <= not (a and b);
    layer4_outputs(1826) <= not (a xor b);
    layer4_outputs(1827) <= not a;
    layer4_outputs(1828) <= not a or b;
    layer4_outputs(1829) <= not (a or b);
    layer4_outputs(1830) <= not a;
    layer4_outputs(1831) <= not a;
    layer4_outputs(1832) <= b and not a;
    layer4_outputs(1833) <= b;
    layer4_outputs(1834) <= b;
    layer4_outputs(1835) <= not b or a;
    layer4_outputs(1836) <= b;
    layer4_outputs(1837) <= not (a or b);
    layer4_outputs(1838) <= a or b;
    layer4_outputs(1839) <= not a;
    layer4_outputs(1840) <= not a or b;
    layer4_outputs(1841) <= b and not a;
    layer4_outputs(1842) <= a and not b;
    layer4_outputs(1843) <= '1';
    layer4_outputs(1844) <= '0';
    layer4_outputs(1845) <= '0';
    layer4_outputs(1846) <= a or b;
    layer4_outputs(1847) <= not b or a;
    layer4_outputs(1848) <= not b;
    layer4_outputs(1849) <= not b;
    layer4_outputs(1850) <= not a or b;
    layer4_outputs(1851) <= not (a xor b);
    layer4_outputs(1852) <= not (a or b);
    layer4_outputs(1853) <= not (a and b);
    layer4_outputs(1854) <= not (a xor b);
    layer4_outputs(1855) <= a and not b;
    layer4_outputs(1856) <= not a or b;
    layer4_outputs(1857) <= a;
    layer4_outputs(1858) <= b;
    layer4_outputs(1859) <= not a;
    layer4_outputs(1860) <= not (a and b);
    layer4_outputs(1861) <= not (a xor b);
    layer4_outputs(1862) <= not b;
    layer4_outputs(1863) <= not (a or b);
    layer4_outputs(1864) <= not b or a;
    layer4_outputs(1865) <= not a or b;
    layer4_outputs(1866) <= a and not b;
    layer4_outputs(1867) <= b and not a;
    layer4_outputs(1868) <= not (a or b);
    layer4_outputs(1869) <= b;
    layer4_outputs(1870) <= a xor b;
    layer4_outputs(1871) <= a;
    layer4_outputs(1872) <= not (a xor b);
    layer4_outputs(1873) <= a or b;
    layer4_outputs(1874) <= not a or b;
    layer4_outputs(1875) <= b and not a;
    layer4_outputs(1876) <= a and not b;
    layer4_outputs(1877) <= not (a and b);
    layer4_outputs(1878) <= not (a and b);
    layer4_outputs(1879) <= not b or a;
    layer4_outputs(1880) <= not a;
    layer4_outputs(1881) <= not (a or b);
    layer4_outputs(1882) <= not (a xor b);
    layer4_outputs(1883) <= a and not b;
    layer4_outputs(1884) <= b and not a;
    layer4_outputs(1885) <= not (a or b);
    layer4_outputs(1886) <= a and not b;
    layer4_outputs(1887) <= not a;
    layer4_outputs(1888) <= a xor b;
    layer4_outputs(1889) <= not a or b;
    layer4_outputs(1890) <= not (a xor b);
    layer4_outputs(1891) <= not b;
    layer4_outputs(1892) <= a and not b;
    layer4_outputs(1893) <= b;
    layer4_outputs(1894) <= not a;
    layer4_outputs(1895) <= a;
    layer4_outputs(1896) <= b;
    layer4_outputs(1897) <= a and b;
    layer4_outputs(1898) <= not (a xor b);
    layer4_outputs(1899) <= a;
    layer4_outputs(1900) <= not a or b;
    layer4_outputs(1901) <= b;
    layer4_outputs(1902) <= not a;
    layer4_outputs(1903) <= '1';
    layer4_outputs(1904) <= not b or a;
    layer4_outputs(1905) <= not b or a;
    layer4_outputs(1906) <= not a or b;
    layer4_outputs(1907) <= not (a or b);
    layer4_outputs(1908) <= not b or a;
    layer4_outputs(1909) <= not b;
    layer4_outputs(1910) <= a;
    layer4_outputs(1911) <= not a or b;
    layer4_outputs(1912) <= a xor b;
    layer4_outputs(1913) <= a;
    layer4_outputs(1914) <= a;
    layer4_outputs(1915) <= not b or a;
    layer4_outputs(1916) <= not b;
    layer4_outputs(1917) <= not b;
    layer4_outputs(1918) <= not b or a;
    layer4_outputs(1919) <= a and b;
    layer4_outputs(1920) <= a;
    layer4_outputs(1921) <= b and not a;
    layer4_outputs(1922) <= b and not a;
    layer4_outputs(1923) <= not b;
    layer4_outputs(1924) <= b;
    layer4_outputs(1925) <= not a or b;
    layer4_outputs(1926) <= a xor b;
    layer4_outputs(1927) <= a and not b;
    layer4_outputs(1928) <= not (a xor b);
    layer4_outputs(1929) <= b;
    layer4_outputs(1930) <= not b;
    layer4_outputs(1931) <= a and b;
    layer4_outputs(1932) <= not (a xor b);
    layer4_outputs(1933) <= not (a xor b);
    layer4_outputs(1934) <= not b or a;
    layer4_outputs(1935) <= not b;
    layer4_outputs(1936) <= '1';
    layer4_outputs(1937) <= not b;
    layer4_outputs(1938) <= '0';
    layer4_outputs(1939) <= not b;
    layer4_outputs(1940) <= not b;
    layer4_outputs(1941) <= b and not a;
    layer4_outputs(1942) <= a or b;
    layer4_outputs(1943) <= a;
    layer4_outputs(1944) <= not a or b;
    layer4_outputs(1945) <= not a or b;
    layer4_outputs(1946) <= a and b;
    layer4_outputs(1947) <= not a;
    layer4_outputs(1948) <= not b;
    layer4_outputs(1949) <= b;
    layer4_outputs(1950) <= not a or b;
    layer4_outputs(1951) <= a;
    layer4_outputs(1952) <= b and not a;
    layer4_outputs(1953) <= a or b;
    layer4_outputs(1954) <= not (a and b);
    layer4_outputs(1955) <= not a or b;
    layer4_outputs(1956) <= a and b;
    layer4_outputs(1957) <= not a;
    layer4_outputs(1958) <= not a;
    layer4_outputs(1959) <= b;
    layer4_outputs(1960) <= not b;
    layer4_outputs(1961) <= b;
    layer4_outputs(1962) <= a;
    layer4_outputs(1963) <= a xor b;
    layer4_outputs(1964) <= b and not a;
    layer4_outputs(1965) <= b;
    layer4_outputs(1966) <= a and b;
    layer4_outputs(1967) <= b;
    layer4_outputs(1968) <= not (a and b);
    layer4_outputs(1969) <= a;
    layer4_outputs(1970) <= not (a or b);
    layer4_outputs(1971) <= not b or a;
    layer4_outputs(1972) <= not b;
    layer4_outputs(1973) <= not a;
    layer4_outputs(1974) <= not a or b;
    layer4_outputs(1975) <= not b;
    layer4_outputs(1976) <= not b;
    layer4_outputs(1977) <= not b or a;
    layer4_outputs(1978) <= not (a and b);
    layer4_outputs(1979) <= not a or b;
    layer4_outputs(1980) <= not b;
    layer4_outputs(1981) <= b and not a;
    layer4_outputs(1982) <= not (a or b);
    layer4_outputs(1983) <= b and not a;
    layer4_outputs(1984) <= a and b;
    layer4_outputs(1985) <= not a or b;
    layer4_outputs(1986) <= not b;
    layer4_outputs(1987) <= a and not b;
    layer4_outputs(1988) <= b and not a;
    layer4_outputs(1989) <= a xor b;
    layer4_outputs(1990) <= not (a or b);
    layer4_outputs(1991) <= a and not b;
    layer4_outputs(1992) <= not a or b;
    layer4_outputs(1993) <= not a;
    layer4_outputs(1994) <= not a;
    layer4_outputs(1995) <= not b;
    layer4_outputs(1996) <= b;
    layer4_outputs(1997) <= b;
    layer4_outputs(1998) <= not b or a;
    layer4_outputs(1999) <= not a;
    layer4_outputs(2000) <= not (a and b);
    layer4_outputs(2001) <= not a;
    layer4_outputs(2002) <= b;
    layer4_outputs(2003) <= not (a and b);
    layer4_outputs(2004) <= not b;
    layer4_outputs(2005) <= not a;
    layer4_outputs(2006) <= not b or a;
    layer4_outputs(2007) <= b and not a;
    layer4_outputs(2008) <= a;
    layer4_outputs(2009) <= b;
    layer4_outputs(2010) <= not a;
    layer4_outputs(2011) <= a and not b;
    layer4_outputs(2012) <= b;
    layer4_outputs(2013) <= a;
    layer4_outputs(2014) <= not b;
    layer4_outputs(2015) <= not b;
    layer4_outputs(2016) <= not a;
    layer4_outputs(2017) <= not a or b;
    layer4_outputs(2018) <= not b or a;
    layer4_outputs(2019) <= a xor b;
    layer4_outputs(2020) <= not b;
    layer4_outputs(2021) <= not b;
    layer4_outputs(2022) <= a xor b;
    layer4_outputs(2023) <= not b or a;
    layer4_outputs(2024) <= not a or b;
    layer4_outputs(2025) <= a and b;
    layer4_outputs(2026) <= a xor b;
    layer4_outputs(2027) <= b and not a;
    layer4_outputs(2028) <= not b or a;
    layer4_outputs(2029) <= a;
    layer4_outputs(2030) <= not a;
    layer4_outputs(2031) <= a or b;
    layer4_outputs(2032) <= b and not a;
    layer4_outputs(2033) <= not a;
    layer4_outputs(2034) <= not b;
    layer4_outputs(2035) <= b and not a;
    layer4_outputs(2036) <= a and not b;
    layer4_outputs(2037) <= not (a or b);
    layer4_outputs(2038) <= not a;
    layer4_outputs(2039) <= not (a and b);
    layer4_outputs(2040) <= b;
    layer4_outputs(2041) <= not b or a;
    layer4_outputs(2042) <= not (a and b);
    layer4_outputs(2043) <= a xor b;
    layer4_outputs(2044) <= b;
    layer4_outputs(2045) <= b and not a;
    layer4_outputs(2046) <= a and not b;
    layer4_outputs(2047) <= not b or a;
    layer4_outputs(2048) <= not (a and b);
    layer4_outputs(2049) <= not a;
    layer4_outputs(2050) <= not a;
    layer4_outputs(2051) <= a or b;
    layer4_outputs(2052) <= a;
    layer4_outputs(2053) <= a and not b;
    layer4_outputs(2054) <= b and not a;
    layer4_outputs(2055) <= b and not a;
    layer4_outputs(2056) <= a xor b;
    layer4_outputs(2057) <= not (a xor b);
    layer4_outputs(2058) <= b and not a;
    layer4_outputs(2059) <= not (a and b);
    layer4_outputs(2060) <= a;
    layer4_outputs(2061) <= a or b;
    layer4_outputs(2062) <= not (a or b);
    layer4_outputs(2063) <= a;
    layer4_outputs(2064) <= not b;
    layer4_outputs(2065) <= '0';
    layer4_outputs(2066) <= a and b;
    layer4_outputs(2067) <= a and not b;
    layer4_outputs(2068) <= not (a xor b);
    layer4_outputs(2069) <= not a;
    layer4_outputs(2070) <= b and not a;
    layer4_outputs(2071) <= b;
    layer4_outputs(2072) <= not b or a;
    layer4_outputs(2073) <= a and b;
    layer4_outputs(2074) <= a or b;
    layer4_outputs(2075) <= a or b;
    layer4_outputs(2076) <= a xor b;
    layer4_outputs(2077) <= a;
    layer4_outputs(2078) <= a;
    layer4_outputs(2079) <= not b;
    layer4_outputs(2080) <= a and b;
    layer4_outputs(2081) <= a or b;
    layer4_outputs(2082) <= b;
    layer4_outputs(2083) <= not a or b;
    layer4_outputs(2084) <= not (a or b);
    layer4_outputs(2085) <= a;
    layer4_outputs(2086) <= b;
    layer4_outputs(2087) <= not a or b;
    layer4_outputs(2088) <= not (a and b);
    layer4_outputs(2089) <= b;
    layer4_outputs(2090) <= a or b;
    layer4_outputs(2091) <= a xor b;
    layer4_outputs(2092) <= b;
    layer4_outputs(2093) <= a;
    layer4_outputs(2094) <= not b;
    layer4_outputs(2095) <= a;
    layer4_outputs(2096) <= not (a and b);
    layer4_outputs(2097) <= b;
    layer4_outputs(2098) <= b and not a;
    layer4_outputs(2099) <= a and not b;
    layer4_outputs(2100) <= not b;
    layer4_outputs(2101) <= a or b;
    layer4_outputs(2102) <= a;
    layer4_outputs(2103) <= not a or b;
    layer4_outputs(2104) <= not (a or b);
    layer4_outputs(2105) <= not a or b;
    layer4_outputs(2106) <= a and b;
    layer4_outputs(2107) <= not (a and b);
    layer4_outputs(2108) <= not (a xor b);
    layer4_outputs(2109) <= '1';
    layer4_outputs(2110) <= b;
    layer4_outputs(2111) <= not a or b;
    layer4_outputs(2112) <= not (a and b);
    layer4_outputs(2113) <= not a;
    layer4_outputs(2114) <= '0';
    layer4_outputs(2115) <= not a;
    layer4_outputs(2116) <= b and not a;
    layer4_outputs(2117) <= '0';
    layer4_outputs(2118) <= not a;
    layer4_outputs(2119) <= not a;
    layer4_outputs(2120) <= not a or b;
    layer4_outputs(2121) <= a;
    layer4_outputs(2122) <= b;
    layer4_outputs(2123) <= a xor b;
    layer4_outputs(2124) <= b;
    layer4_outputs(2125) <= a and not b;
    layer4_outputs(2126) <= b;
    layer4_outputs(2127) <= '0';
    layer4_outputs(2128) <= a or b;
    layer4_outputs(2129) <= not (a and b);
    layer4_outputs(2130) <= a xor b;
    layer4_outputs(2131) <= b and not a;
    layer4_outputs(2132) <= b and not a;
    layer4_outputs(2133) <= not b;
    layer4_outputs(2134) <= a;
    layer4_outputs(2135) <= not b;
    layer4_outputs(2136) <= not b or a;
    layer4_outputs(2137) <= not b;
    layer4_outputs(2138) <= not (a xor b);
    layer4_outputs(2139) <= not b or a;
    layer4_outputs(2140) <= not (a and b);
    layer4_outputs(2141) <= a;
    layer4_outputs(2142) <= a;
    layer4_outputs(2143) <= not (a xor b);
    layer4_outputs(2144) <= a and b;
    layer4_outputs(2145) <= a and not b;
    layer4_outputs(2146) <= b and not a;
    layer4_outputs(2147) <= not (a xor b);
    layer4_outputs(2148) <= not a;
    layer4_outputs(2149) <= b and not a;
    layer4_outputs(2150) <= a;
    layer4_outputs(2151) <= a xor b;
    layer4_outputs(2152) <= a and b;
    layer4_outputs(2153) <= b and not a;
    layer4_outputs(2154) <= not (a or b);
    layer4_outputs(2155) <= not a;
    layer4_outputs(2156) <= a and b;
    layer4_outputs(2157) <= a xor b;
    layer4_outputs(2158) <= a or b;
    layer4_outputs(2159) <= a and not b;
    layer4_outputs(2160) <= not b or a;
    layer4_outputs(2161) <= b;
    layer4_outputs(2162) <= a xor b;
    layer4_outputs(2163) <= a xor b;
    layer4_outputs(2164) <= a xor b;
    layer4_outputs(2165) <= not (a and b);
    layer4_outputs(2166) <= a and not b;
    layer4_outputs(2167) <= a or b;
    layer4_outputs(2168) <= b;
    layer4_outputs(2169) <= '1';
    layer4_outputs(2170) <= not a;
    layer4_outputs(2171) <= not (a or b);
    layer4_outputs(2172) <= '1';
    layer4_outputs(2173) <= a and not b;
    layer4_outputs(2174) <= not (a and b);
    layer4_outputs(2175) <= not b or a;
    layer4_outputs(2176) <= b and not a;
    layer4_outputs(2177) <= a xor b;
    layer4_outputs(2178) <= not (a and b);
    layer4_outputs(2179) <= not a or b;
    layer4_outputs(2180) <= b and not a;
    layer4_outputs(2181) <= b and not a;
    layer4_outputs(2182) <= b and not a;
    layer4_outputs(2183) <= not (a or b);
    layer4_outputs(2184) <= '1';
    layer4_outputs(2185) <= not (a xor b);
    layer4_outputs(2186) <= a;
    layer4_outputs(2187) <= a or b;
    layer4_outputs(2188) <= '1';
    layer4_outputs(2189) <= a or b;
    layer4_outputs(2190) <= not b or a;
    layer4_outputs(2191) <= not (a or b);
    layer4_outputs(2192) <= not (a or b);
    layer4_outputs(2193) <= not a;
    layer4_outputs(2194) <= not a;
    layer4_outputs(2195) <= not b;
    layer4_outputs(2196) <= b;
    layer4_outputs(2197) <= b;
    layer4_outputs(2198) <= b;
    layer4_outputs(2199) <= not (a or b);
    layer4_outputs(2200) <= '1';
    layer4_outputs(2201) <= '1';
    layer4_outputs(2202) <= not (a and b);
    layer4_outputs(2203) <= a;
    layer4_outputs(2204) <= not a;
    layer4_outputs(2205) <= not (a or b);
    layer4_outputs(2206) <= '0';
    layer4_outputs(2207) <= a;
    layer4_outputs(2208) <= not a;
    layer4_outputs(2209) <= b and not a;
    layer4_outputs(2210) <= '1';
    layer4_outputs(2211) <= '0';
    layer4_outputs(2212) <= not a;
    layer4_outputs(2213) <= not (a or b);
    layer4_outputs(2214) <= b;
    layer4_outputs(2215) <= not b;
    layer4_outputs(2216) <= not a or b;
    layer4_outputs(2217) <= b;
    layer4_outputs(2218) <= not b or a;
    layer4_outputs(2219) <= not (a or b);
    layer4_outputs(2220) <= a;
    layer4_outputs(2221) <= not (a and b);
    layer4_outputs(2222) <= a xor b;
    layer4_outputs(2223) <= not (a and b);
    layer4_outputs(2224) <= not a;
    layer4_outputs(2225) <= not (a or b);
    layer4_outputs(2226) <= not (a or b);
    layer4_outputs(2227) <= b and not a;
    layer4_outputs(2228) <= not (a and b);
    layer4_outputs(2229) <= a and b;
    layer4_outputs(2230) <= b;
    layer4_outputs(2231) <= a;
    layer4_outputs(2232) <= a;
    layer4_outputs(2233) <= not a;
    layer4_outputs(2234) <= b;
    layer4_outputs(2235) <= not (a and b);
    layer4_outputs(2236) <= not (a xor b);
    layer4_outputs(2237) <= a and b;
    layer4_outputs(2238) <= a;
    layer4_outputs(2239) <= not b or a;
    layer4_outputs(2240) <= not a;
    layer4_outputs(2241) <= not (a or b);
    layer4_outputs(2242) <= b;
    layer4_outputs(2243) <= b;
    layer4_outputs(2244) <= not b;
    layer4_outputs(2245) <= not a;
    layer4_outputs(2246) <= b and not a;
    layer4_outputs(2247) <= a;
    layer4_outputs(2248) <= not (a xor b);
    layer4_outputs(2249) <= b;
    layer4_outputs(2250) <= a;
    layer4_outputs(2251) <= b;
    layer4_outputs(2252) <= not b;
    layer4_outputs(2253) <= a xor b;
    layer4_outputs(2254) <= b;
    layer4_outputs(2255) <= a xor b;
    layer4_outputs(2256) <= not b;
    layer4_outputs(2257) <= b;
    layer4_outputs(2258) <= not a or b;
    layer4_outputs(2259) <= a;
    layer4_outputs(2260) <= '0';
    layer4_outputs(2261) <= b and not a;
    layer4_outputs(2262) <= a and b;
    layer4_outputs(2263) <= b;
    layer4_outputs(2264) <= not a;
    layer4_outputs(2265) <= '0';
    layer4_outputs(2266) <= a;
    layer4_outputs(2267) <= not (a or b);
    layer4_outputs(2268) <= b;
    layer4_outputs(2269) <= a and b;
    layer4_outputs(2270) <= a and not b;
    layer4_outputs(2271) <= not b;
    layer4_outputs(2272) <= '1';
    layer4_outputs(2273) <= not (a xor b);
    layer4_outputs(2274) <= not b or a;
    layer4_outputs(2275) <= '0';
    layer4_outputs(2276) <= a and not b;
    layer4_outputs(2277) <= b and not a;
    layer4_outputs(2278) <= b and not a;
    layer4_outputs(2279) <= not a;
    layer4_outputs(2280) <= b;
    layer4_outputs(2281) <= not (a xor b);
    layer4_outputs(2282) <= b and not a;
    layer4_outputs(2283) <= not a;
    layer4_outputs(2284) <= a xor b;
    layer4_outputs(2285) <= not a;
    layer4_outputs(2286) <= not (a and b);
    layer4_outputs(2287) <= not b or a;
    layer4_outputs(2288) <= '1';
    layer4_outputs(2289) <= not (a and b);
    layer4_outputs(2290) <= b;
    layer4_outputs(2291) <= not b;
    layer4_outputs(2292) <= a;
    layer4_outputs(2293) <= not a;
    layer4_outputs(2294) <= not a;
    layer4_outputs(2295) <= a xor b;
    layer4_outputs(2296) <= b;
    layer4_outputs(2297) <= b and not a;
    layer4_outputs(2298) <= not (a xor b);
    layer4_outputs(2299) <= not b or a;
    layer4_outputs(2300) <= a xor b;
    layer4_outputs(2301) <= a xor b;
    layer4_outputs(2302) <= not (a xor b);
    layer4_outputs(2303) <= a and not b;
    layer4_outputs(2304) <= a;
    layer4_outputs(2305) <= b and not a;
    layer4_outputs(2306) <= a xor b;
    layer4_outputs(2307) <= a and b;
    layer4_outputs(2308) <= a;
    layer4_outputs(2309) <= not (a or b);
    layer4_outputs(2310) <= a or b;
    layer4_outputs(2311) <= b;
    layer4_outputs(2312) <= a and not b;
    layer4_outputs(2313) <= not (a xor b);
    layer4_outputs(2314) <= not (a and b);
    layer4_outputs(2315) <= b;
    layer4_outputs(2316) <= not a;
    layer4_outputs(2317) <= b;
    layer4_outputs(2318) <= b and not a;
    layer4_outputs(2319) <= a or b;
    layer4_outputs(2320) <= b and not a;
    layer4_outputs(2321) <= not b;
    layer4_outputs(2322) <= b;
    layer4_outputs(2323) <= not b;
    layer4_outputs(2324) <= a xor b;
    layer4_outputs(2325) <= a;
    layer4_outputs(2326) <= a or b;
    layer4_outputs(2327) <= not (a or b);
    layer4_outputs(2328) <= a xor b;
    layer4_outputs(2329) <= not a;
    layer4_outputs(2330) <= not b;
    layer4_outputs(2331) <= not a;
    layer4_outputs(2332) <= not b;
    layer4_outputs(2333) <= not a or b;
    layer4_outputs(2334) <= b;
    layer4_outputs(2335) <= b;
    layer4_outputs(2336) <= not a or b;
    layer4_outputs(2337) <= not b;
    layer4_outputs(2338) <= not (a xor b);
    layer4_outputs(2339) <= not a;
    layer4_outputs(2340) <= a;
    layer4_outputs(2341) <= a and not b;
    layer4_outputs(2342) <= not a or b;
    layer4_outputs(2343) <= a;
    layer4_outputs(2344) <= not (a xor b);
    layer4_outputs(2345) <= not (a and b);
    layer4_outputs(2346) <= not b;
    layer4_outputs(2347) <= a;
    layer4_outputs(2348) <= not b;
    layer4_outputs(2349) <= b and not a;
    layer4_outputs(2350) <= a or b;
    layer4_outputs(2351) <= not (a or b);
    layer4_outputs(2352) <= a or b;
    layer4_outputs(2353) <= not b;
    layer4_outputs(2354) <= not (a xor b);
    layer4_outputs(2355) <= a and not b;
    layer4_outputs(2356) <= b;
    layer4_outputs(2357) <= not (a xor b);
    layer4_outputs(2358) <= not (a and b);
    layer4_outputs(2359) <= not a or b;
    layer4_outputs(2360) <= a or b;
    layer4_outputs(2361) <= b;
    layer4_outputs(2362) <= b;
    layer4_outputs(2363) <= not a or b;
    layer4_outputs(2364) <= a;
    layer4_outputs(2365) <= not a;
    layer4_outputs(2366) <= not (a or b);
    layer4_outputs(2367) <= a or b;
    layer4_outputs(2368) <= '1';
    layer4_outputs(2369) <= a;
    layer4_outputs(2370) <= a and not b;
    layer4_outputs(2371) <= not b;
    layer4_outputs(2372) <= not (a xor b);
    layer4_outputs(2373) <= b and not a;
    layer4_outputs(2374) <= a xor b;
    layer4_outputs(2375) <= a;
    layer4_outputs(2376) <= b and not a;
    layer4_outputs(2377) <= a;
    layer4_outputs(2378) <= a and not b;
    layer4_outputs(2379) <= a and not b;
    layer4_outputs(2380) <= not (a or b);
    layer4_outputs(2381) <= not a;
    layer4_outputs(2382) <= '0';
    layer4_outputs(2383) <= a and not b;
    layer4_outputs(2384) <= not b;
    layer4_outputs(2385) <= a or b;
    layer4_outputs(2386) <= not (a xor b);
    layer4_outputs(2387) <= a or b;
    layer4_outputs(2388) <= a or b;
    layer4_outputs(2389) <= a and not b;
    layer4_outputs(2390) <= a xor b;
    layer4_outputs(2391) <= not b or a;
    layer4_outputs(2392) <= a or b;
    layer4_outputs(2393) <= a;
    layer4_outputs(2394) <= not (a and b);
    layer4_outputs(2395) <= a and b;
    layer4_outputs(2396) <= a;
    layer4_outputs(2397) <= a xor b;
    layer4_outputs(2398) <= not b or a;
    layer4_outputs(2399) <= not b;
    layer4_outputs(2400) <= a;
    layer4_outputs(2401) <= not (a or b);
    layer4_outputs(2402) <= a;
    layer4_outputs(2403) <= not a;
    layer4_outputs(2404) <= a;
    layer4_outputs(2405) <= b;
    layer4_outputs(2406) <= not (a and b);
    layer4_outputs(2407) <= not (a and b);
    layer4_outputs(2408) <= not b;
    layer4_outputs(2409) <= a and not b;
    layer4_outputs(2410) <= not a or b;
    layer4_outputs(2411) <= not a;
    layer4_outputs(2412) <= a xor b;
    layer4_outputs(2413) <= a and b;
    layer4_outputs(2414) <= not (a and b);
    layer4_outputs(2415) <= not b or a;
    layer4_outputs(2416) <= a or b;
    layer4_outputs(2417) <= not b;
    layer4_outputs(2418) <= b;
    layer4_outputs(2419) <= not (a or b);
    layer4_outputs(2420) <= a;
    layer4_outputs(2421) <= a and not b;
    layer4_outputs(2422) <= not b or a;
    layer4_outputs(2423) <= not a;
    layer4_outputs(2424) <= not a or b;
    layer4_outputs(2425) <= not b;
    layer4_outputs(2426) <= a and b;
    layer4_outputs(2427) <= a xor b;
    layer4_outputs(2428) <= a;
    layer4_outputs(2429) <= not a or b;
    layer4_outputs(2430) <= not (a xor b);
    layer4_outputs(2431) <= not a;
    layer4_outputs(2432) <= a or b;
    layer4_outputs(2433) <= b;
    layer4_outputs(2434) <= not (a and b);
    layer4_outputs(2435) <= not a;
    layer4_outputs(2436) <= a and not b;
    layer4_outputs(2437) <= a and b;
    layer4_outputs(2438) <= not a or b;
    layer4_outputs(2439) <= a;
    layer4_outputs(2440) <= not b;
    layer4_outputs(2441) <= not b or a;
    layer4_outputs(2442) <= not b;
    layer4_outputs(2443) <= not (a xor b);
    layer4_outputs(2444) <= a;
    layer4_outputs(2445) <= a;
    layer4_outputs(2446) <= '1';
    layer4_outputs(2447) <= not (a xor b);
    layer4_outputs(2448) <= b;
    layer4_outputs(2449) <= b;
    layer4_outputs(2450) <= not (a xor b);
    layer4_outputs(2451) <= not a or b;
    layer4_outputs(2452) <= not b or a;
    layer4_outputs(2453) <= a;
    layer4_outputs(2454) <= not a;
    layer4_outputs(2455) <= '1';
    layer4_outputs(2456) <= a;
    layer4_outputs(2457) <= not a;
    layer4_outputs(2458) <= b;
    layer4_outputs(2459) <= a and not b;
    layer4_outputs(2460) <= not b;
    layer4_outputs(2461) <= a and not b;
    layer4_outputs(2462) <= a xor b;
    layer4_outputs(2463) <= b;
    layer4_outputs(2464) <= not b;
    layer4_outputs(2465) <= a xor b;
    layer4_outputs(2466) <= '1';
    layer4_outputs(2467) <= b;
    layer4_outputs(2468) <= not b or a;
    layer4_outputs(2469) <= not b;
    layer4_outputs(2470) <= not b;
    layer4_outputs(2471) <= a;
    layer4_outputs(2472) <= not a;
    layer4_outputs(2473) <= not a;
    layer4_outputs(2474) <= not b or a;
    layer4_outputs(2475) <= b and not a;
    layer4_outputs(2476) <= b;
    layer4_outputs(2477) <= '1';
    layer4_outputs(2478) <= a xor b;
    layer4_outputs(2479) <= not b;
    layer4_outputs(2480) <= b;
    layer4_outputs(2481) <= '1';
    layer4_outputs(2482) <= not a;
    layer4_outputs(2483) <= '1';
    layer4_outputs(2484) <= not a;
    layer4_outputs(2485) <= not b;
    layer4_outputs(2486) <= a or b;
    layer4_outputs(2487) <= not b;
    layer4_outputs(2488) <= b;
    layer4_outputs(2489) <= a and b;
    layer4_outputs(2490) <= not a;
    layer4_outputs(2491) <= a and not b;
    layer4_outputs(2492) <= not a;
    layer4_outputs(2493) <= a;
    layer4_outputs(2494) <= not a;
    layer4_outputs(2495) <= a;
    layer4_outputs(2496) <= not b;
    layer4_outputs(2497) <= '0';
    layer4_outputs(2498) <= not b;
    layer4_outputs(2499) <= a xor b;
    layer4_outputs(2500) <= a or b;
    layer4_outputs(2501) <= not a;
    layer4_outputs(2502) <= not b;
    layer4_outputs(2503) <= not a or b;
    layer4_outputs(2504) <= a or b;
    layer4_outputs(2505) <= not (a or b);
    layer4_outputs(2506) <= b;
    layer4_outputs(2507) <= not a;
    layer4_outputs(2508) <= a xor b;
    layer4_outputs(2509) <= b;
    layer4_outputs(2510) <= not (a or b);
    layer4_outputs(2511) <= a xor b;
    layer4_outputs(2512) <= not (a and b);
    layer4_outputs(2513) <= b;
    layer4_outputs(2514) <= b;
    layer4_outputs(2515) <= b;
    layer4_outputs(2516) <= b and not a;
    layer4_outputs(2517) <= b;
    layer4_outputs(2518) <= not a or b;
    layer4_outputs(2519) <= a and b;
    layer4_outputs(2520) <= b and not a;
    layer4_outputs(2521) <= a xor b;
    layer4_outputs(2522) <= not a;
    layer4_outputs(2523) <= b;
    layer4_outputs(2524) <= a;
    layer4_outputs(2525) <= a xor b;
    layer4_outputs(2526) <= a;
    layer4_outputs(2527) <= a or b;
    layer4_outputs(2528) <= b and not a;
    layer4_outputs(2529) <= a or b;
    layer4_outputs(2530) <= not b or a;
    layer4_outputs(2531) <= '1';
    layer4_outputs(2532) <= '0';
    layer4_outputs(2533) <= a and b;
    layer4_outputs(2534) <= a;
    layer4_outputs(2535) <= not a or b;
    layer4_outputs(2536) <= a;
    layer4_outputs(2537) <= not (a or b);
    layer4_outputs(2538) <= not a;
    layer4_outputs(2539) <= a;
    layer4_outputs(2540) <= b;
    layer4_outputs(2541) <= a;
    layer4_outputs(2542) <= not (a or b);
    layer4_outputs(2543) <= not b;
    layer4_outputs(2544) <= not b;
    layer4_outputs(2545) <= a;
    layer4_outputs(2546) <= b and not a;
    layer4_outputs(2547) <= not b;
    layer4_outputs(2548) <= b;
    layer4_outputs(2549) <= not b;
    layer4_outputs(2550) <= a and b;
    layer4_outputs(2551) <= not (a or b);
    layer4_outputs(2552) <= a;
    layer4_outputs(2553) <= not b or a;
    layer4_outputs(2554) <= not (a or b);
    layer4_outputs(2555) <= not (a and b);
    layer4_outputs(2556) <= a or b;
    layer4_outputs(2557) <= not b or a;
    layer4_outputs(2558) <= not (a xor b);
    layer4_outputs(2559) <= not (a and b);
    layer4_outputs(2560) <= a and not b;
    layer4_outputs(2561) <= not b;
    layer4_outputs(2562) <= a or b;
    layer4_outputs(2563) <= a and not b;
    layer4_outputs(2564) <= not b or a;
    layer4_outputs(2565) <= not (a or b);
    layer4_outputs(2566) <= b;
    layer4_outputs(2567) <= not (a xor b);
    layer4_outputs(2568) <= '1';
    layer4_outputs(2569) <= a;
    layer4_outputs(2570) <= not (a xor b);
    layer4_outputs(2571) <= not a;
    layer4_outputs(2572) <= '1';
    layer4_outputs(2573) <= a;
    layer4_outputs(2574) <= a xor b;
    layer4_outputs(2575) <= not a;
    layer4_outputs(2576) <= b and not a;
    layer4_outputs(2577) <= a or b;
    layer4_outputs(2578) <= not (a and b);
    layer4_outputs(2579) <= a or b;
    layer4_outputs(2580) <= '1';
    layer4_outputs(2581) <= not a or b;
    layer4_outputs(2582) <= b;
    layer4_outputs(2583) <= a and not b;
    layer4_outputs(2584) <= b;
    layer4_outputs(2585) <= '1';
    layer4_outputs(2586) <= not (a or b);
    layer4_outputs(2587) <= a;
    layer4_outputs(2588) <= a or b;
    layer4_outputs(2589) <= not a or b;
    layer4_outputs(2590) <= not a;
    layer4_outputs(2591) <= b and not a;
    layer4_outputs(2592) <= b;
    layer4_outputs(2593) <= a xor b;
    layer4_outputs(2594) <= not (a xor b);
    layer4_outputs(2595) <= a and not b;
    layer4_outputs(2596) <= not (a or b);
    layer4_outputs(2597) <= '0';
    layer4_outputs(2598) <= b;
    layer4_outputs(2599) <= not a;
    layer4_outputs(2600) <= not b or a;
    layer4_outputs(2601) <= b;
    layer4_outputs(2602) <= a and b;
    layer4_outputs(2603) <= not b or a;
    layer4_outputs(2604) <= a and not b;
    layer4_outputs(2605) <= not a;
    layer4_outputs(2606) <= b;
    layer4_outputs(2607) <= not (a or b);
    layer4_outputs(2608) <= not (a xor b);
    layer4_outputs(2609) <= a;
    layer4_outputs(2610) <= not b;
    layer4_outputs(2611) <= not (a xor b);
    layer4_outputs(2612) <= a;
    layer4_outputs(2613) <= not a or b;
    layer4_outputs(2614) <= not b or a;
    layer4_outputs(2615) <= b;
    layer4_outputs(2616) <= b;
    layer4_outputs(2617) <= not (a or b);
    layer4_outputs(2618) <= not b;
    layer4_outputs(2619) <= a;
    layer4_outputs(2620) <= not (a or b);
    layer4_outputs(2621) <= not (a xor b);
    layer4_outputs(2622) <= a and b;
    layer4_outputs(2623) <= not (a xor b);
    layer4_outputs(2624) <= not a or b;
    layer4_outputs(2625) <= not (a and b);
    layer4_outputs(2626) <= not (a xor b);
    layer4_outputs(2627) <= not b or a;
    layer4_outputs(2628) <= not (a xor b);
    layer4_outputs(2629) <= a and not b;
    layer4_outputs(2630) <= a or b;
    layer4_outputs(2631) <= a;
    layer4_outputs(2632) <= a;
    layer4_outputs(2633) <= a and not b;
    layer4_outputs(2634) <= not a or b;
    layer4_outputs(2635) <= '0';
    layer4_outputs(2636) <= not (a xor b);
    layer4_outputs(2637) <= not b;
    layer4_outputs(2638) <= not b;
    layer4_outputs(2639) <= not a;
    layer4_outputs(2640) <= a and not b;
    layer4_outputs(2641) <= not (a xor b);
    layer4_outputs(2642) <= not a;
    layer4_outputs(2643) <= a xor b;
    layer4_outputs(2644) <= not (a and b);
    layer4_outputs(2645) <= '0';
    layer4_outputs(2646) <= not b or a;
    layer4_outputs(2647) <= not a or b;
    layer4_outputs(2648) <= a or b;
    layer4_outputs(2649) <= not b;
    layer4_outputs(2650) <= not b;
    layer4_outputs(2651) <= a xor b;
    layer4_outputs(2652) <= a;
    layer4_outputs(2653) <= not a;
    layer4_outputs(2654) <= b;
    layer4_outputs(2655) <= not a;
    layer4_outputs(2656) <= not b;
    layer4_outputs(2657) <= a or b;
    layer4_outputs(2658) <= a and b;
    layer4_outputs(2659) <= not a;
    layer4_outputs(2660) <= not a;
    layer4_outputs(2661) <= b;
    layer4_outputs(2662) <= not a;
    layer4_outputs(2663) <= not a;
    layer4_outputs(2664) <= a or b;
    layer4_outputs(2665) <= a xor b;
    layer4_outputs(2666) <= a xor b;
    layer4_outputs(2667) <= not a or b;
    layer4_outputs(2668) <= not (a xor b);
    layer4_outputs(2669) <= b and not a;
    layer4_outputs(2670) <= a or b;
    layer4_outputs(2671) <= a;
    layer4_outputs(2672) <= '1';
    layer4_outputs(2673) <= a and not b;
    layer4_outputs(2674) <= '1';
    layer4_outputs(2675) <= not b;
    layer4_outputs(2676) <= a and b;
    layer4_outputs(2677) <= a or b;
    layer4_outputs(2678) <= b;
    layer4_outputs(2679) <= b and not a;
    layer4_outputs(2680) <= not a or b;
    layer4_outputs(2681) <= not b;
    layer4_outputs(2682) <= a;
    layer4_outputs(2683) <= not (a or b);
    layer4_outputs(2684) <= b;
    layer4_outputs(2685) <= a and b;
    layer4_outputs(2686) <= a and b;
    layer4_outputs(2687) <= a and not b;
    layer4_outputs(2688) <= not b or a;
    layer4_outputs(2689) <= a;
    layer4_outputs(2690) <= not b;
    layer4_outputs(2691) <= not b;
    layer4_outputs(2692) <= not b;
    layer4_outputs(2693) <= a xor b;
    layer4_outputs(2694) <= not b;
    layer4_outputs(2695) <= not b;
    layer4_outputs(2696) <= a;
    layer4_outputs(2697) <= not a;
    layer4_outputs(2698) <= not (a xor b);
    layer4_outputs(2699) <= a or b;
    layer4_outputs(2700) <= a and b;
    layer4_outputs(2701) <= a and not b;
    layer4_outputs(2702) <= '0';
    layer4_outputs(2703) <= a;
    layer4_outputs(2704) <= a;
    layer4_outputs(2705) <= not a or b;
    layer4_outputs(2706) <= a;
    layer4_outputs(2707) <= not a;
    layer4_outputs(2708) <= b;
    layer4_outputs(2709) <= a and not b;
    layer4_outputs(2710) <= not (a xor b);
    layer4_outputs(2711) <= not b;
    layer4_outputs(2712) <= not b;
    layer4_outputs(2713) <= a or b;
    layer4_outputs(2714) <= b and not a;
    layer4_outputs(2715) <= not a;
    layer4_outputs(2716) <= not a or b;
    layer4_outputs(2717) <= a;
    layer4_outputs(2718) <= not (a or b);
    layer4_outputs(2719) <= b;
    layer4_outputs(2720) <= not a;
    layer4_outputs(2721) <= b;
    layer4_outputs(2722) <= not b;
    layer4_outputs(2723) <= not a or b;
    layer4_outputs(2724) <= a and not b;
    layer4_outputs(2725) <= b and not a;
    layer4_outputs(2726) <= not b or a;
    layer4_outputs(2727) <= not b;
    layer4_outputs(2728) <= b;
    layer4_outputs(2729) <= not b;
    layer4_outputs(2730) <= '0';
    layer4_outputs(2731) <= not (a xor b);
    layer4_outputs(2732) <= a and b;
    layer4_outputs(2733) <= not b or a;
    layer4_outputs(2734) <= not a;
    layer4_outputs(2735) <= not (a or b);
    layer4_outputs(2736) <= a and not b;
    layer4_outputs(2737) <= a and b;
    layer4_outputs(2738) <= not a;
    layer4_outputs(2739) <= not b or a;
    layer4_outputs(2740) <= not (a xor b);
    layer4_outputs(2741) <= not a;
    layer4_outputs(2742) <= a and b;
    layer4_outputs(2743) <= b;
    layer4_outputs(2744) <= a and not b;
    layer4_outputs(2745) <= a;
    layer4_outputs(2746) <= not a or b;
    layer4_outputs(2747) <= '0';
    layer4_outputs(2748) <= not (a and b);
    layer4_outputs(2749) <= not a or b;
    layer4_outputs(2750) <= not (a and b);
    layer4_outputs(2751) <= not b;
    layer4_outputs(2752) <= not a;
    layer4_outputs(2753) <= not b;
    layer4_outputs(2754) <= a or b;
    layer4_outputs(2755) <= not b;
    layer4_outputs(2756) <= not a;
    layer4_outputs(2757) <= not a;
    layer4_outputs(2758) <= a;
    layer4_outputs(2759) <= a;
    layer4_outputs(2760) <= a or b;
    layer4_outputs(2761) <= not (a or b);
    layer4_outputs(2762) <= not b or a;
    layer4_outputs(2763) <= not a;
    layer4_outputs(2764) <= not b;
    layer4_outputs(2765) <= not a;
    layer4_outputs(2766) <= b;
    layer4_outputs(2767) <= not (a or b);
    layer4_outputs(2768) <= not (a xor b);
    layer4_outputs(2769) <= a;
    layer4_outputs(2770) <= b and not a;
    layer4_outputs(2771) <= not a;
    layer4_outputs(2772) <= not (a and b);
    layer4_outputs(2773) <= not b or a;
    layer4_outputs(2774) <= a;
    layer4_outputs(2775) <= b and not a;
    layer4_outputs(2776) <= b and not a;
    layer4_outputs(2777) <= not a;
    layer4_outputs(2778) <= a;
    layer4_outputs(2779) <= '0';
    layer4_outputs(2780) <= not b or a;
    layer4_outputs(2781) <= a and b;
    layer4_outputs(2782) <= a xor b;
    layer4_outputs(2783) <= a;
    layer4_outputs(2784) <= a and b;
    layer4_outputs(2785) <= not (a and b);
    layer4_outputs(2786) <= a;
    layer4_outputs(2787) <= not a;
    layer4_outputs(2788) <= not (a xor b);
    layer4_outputs(2789) <= b;
    layer4_outputs(2790) <= not (a xor b);
    layer4_outputs(2791) <= b;
    layer4_outputs(2792) <= not a;
    layer4_outputs(2793) <= a or b;
    layer4_outputs(2794) <= not a;
    layer4_outputs(2795) <= not (a xor b);
    layer4_outputs(2796) <= b;
    layer4_outputs(2797) <= not (a and b);
    layer4_outputs(2798) <= not a or b;
    layer4_outputs(2799) <= not a or b;
    layer4_outputs(2800) <= a and not b;
    layer4_outputs(2801) <= not (a xor b);
    layer4_outputs(2802) <= not b;
    layer4_outputs(2803) <= not a or b;
    layer4_outputs(2804) <= a;
    layer4_outputs(2805) <= not b or a;
    layer4_outputs(2806) <= a xor b;
    layer4_outputs(2807) <= a;
    layer4_outputs(2808) <= not a;
    layer4_outputs(2809) <= not b;
    layer4_outputs(2810) <= a and b;
    layer4_outputs(2811) <= a;
    layer4_outputs(2812) <= not a;
    layer4_outputs(2813) <= b;
    layer4_outputs(2814) <= a or b;
    layer4_outputs(2815) <= not a or b;
    layer4_outputs(2816) <= a xor b;
    layer4_outputs(2817) <= '1';
    layer4_outputs(2818) <= not b or a;
    layer4_outputs(2819) <= not b or a;
    layer4_outputs(2820) <= a and not b;
    layer4_outputs(2821) <= '0';
    layer4_outputs(2822) <= b and not a;
    layer4_outputs(2823) <= not b;
    layer4_outputs(2824) <= not b;
    layer4_outputs(2825) <= '0';
    layer4_outputs(2826) <= a and b;
    layer4_outputs(2827) <= not (a and b);
    layer4_outputs(2828) <= a;
    layer4_outputs(2829) <= not b or a;
    layer4_outputs(2830) <= a;
    layer4_outputs(2831) <= '1';
    layer4_outputs(2832) <= a and not b;
    layer4_outputs(2833) <= a xor b;
    layer4_outputs(2834) <= b;
    layer4_outputs(2835) <= a and not b;
    layer4_outputs(2836) <= a xor b;
    layer4_outputs(2837) <= not (a xor b);
    layer4_outputs(2838) <= not (a or b);
    layer4_outputs(2839) <= not b;
    layer4_outputs(2840) <= not (a xor b);
    layer4_outputs(2841) <= b;
    layer4_outputs(2842) <= not b or a;
    layer4_outputs(2843) <= not a;
    layer4_outputs(2844) <= not (a or b);
    layer4_outputs(2845) <= a;
    layer4_outputs(2846) <= not a;
    layer4_outputs(2847) <= not a;
    layer4_outputs(2848) <= not a;
    layer4_outputs(2849) <= not a;
    layer4_outputs(2850) <= a xor b;
    layer4_outputs(2851) <= b;
    layer4_outputs(2852) <= not a;
    layer4_outputs(2853) <= not a;
    layer4_outputs(2854) <= a xor b;
    layer4_outputs(2855) <= not b;
    layer4_outputs(2856) <= b;
    layer4_outputs(2857) <= not a;
    layer4_outputs(2858) <= not b or a;
    layer4_outputs(2859) <= not (a xor b);
    layer4_outputs(2860) <= not b;
    layer4_outputs(2861) <= not a;
    layer4_outputs(2862) <= b and not a;
    layer4_outputs(2863) <= a and b;
    layer4_outputs(2864) <= not b;
    layer4_outputs(2865) <= not b;
    layer4_outputs(2866) <= a or b;
    layer4_outputs(2867) <= '1';
    layer4_outputs(2868) <= not b;
    layer4_outputs(2869) <= not a;
    layer4_outputs(2870) <= b;
    layer4_outputs(2871) <= not (a and b);
    layer4_outputs(2872) <= '1';
    layer4_outputs(2873) <= a xor b;
    layer4_outputs(2874) <= not b;
    layer4_outputs(2875) <= not b;
    layer4_outputs(2876) <= not a or b;
    layer4_outputs(2877) <= not b;
    layer4_outputs(2878) <= not b or a;
    layer4_outputs(2879) <= not (a xor b);
    layer4_outputs(2880) <= not a;
    layer4_outputs(2881) <= a and not b;
    layer4_outputs(2882) <= a xor b;
    layer4_outputs(2883) <= b;
    layer4_outputs(2884) <= not a;
    layer4_outputs(2885) <= a and not b;
    layer4_outputs(2886) <= b and not a;
    layer4_outputs(2887) <= b;
    layer4_outputs(2888) <= a and not b;
    layer4_outputs(2889) <= a;
    layer4_outputs(2890) <= not (a and b);
    layer4_outputs(2891) <= not a or b;
    layer4_outputs(2892) <= not b or a;
    layer4_outputs(2893) <= not b or a;
    layer4_outputs(2894) <= a;
    layer4_outputs(2895) <= not a;
    layer4_outputs(2896) <= a or b;
    layer4_outputs(2897) <= not a or b;
    layer4_outputs(2898) <= a and not b;
    layer4_outputs(2899) <= not b;
    layer4_outputs(2900) <= not a or b;
    layer4_outputs(2901) <= not a;
    layer4_outputs(2902) <= a;
    layer4_outputs(2903) <= a xor b;
    layer4_outputs(2904) <= a and not b;
    layer4_outputs(2905) <= not (a or b);
    layer4_outputs(2906) <= not (a and b);
    layer4_outputs(2907) <= a or b;
    layer4_outputs(2908) <= not a or b;
    layer4_outputs(2909) <= b and not a;
    layer4_outputs(2910) <= not a;
    layer4_outputs(2911) <= a and not b;
    layer4_outputs(2912) <= a;
    layer4_outputs(2913) <= not b;
    layer4_outputs(2914) <= a xor b;
    layer4_outputs(2915) <= not a;
    layer4_outputs(2916) <= not b;
    layer4_outputs(2917) <= not (a and b);
    layer4_outputs(2918) <= not b;
    layer4_outputs(2919) <= a and not b;
    layer4_outputs(2920) <= a and not b;
    layer4_outputs(2921) <= not a;
    layer4_outputs(2922) <= b and not a;
    layer4_outputs(2923) <= b and not a;
    layer4_outputs(2924) <= a and b;
    layer4_outputs(2925) <= a and b;
    layer4_outputs(2926) <= b;
    layer4_outputs(2927) <= a and b;
    layer4_outputs(2928) <= a and not b;
    layer4_outputs(2929) <= a or b;
    layer4_outputs(2930) <= not a;
    layer4_outputs(2931) <= b and not a;
    layer4_outputs(2932) <= not a;
    layer4_outputs(2933) <= not a;
    layer4_outputs(2934) <= not a;
    layer4_outputs(2935) <= not b or a;
    layer4_outputs(2936) <= a and not b;
    layer4_outputs(2937) <= b and not a;
    layer4_outputs(2938) <= b and not a;
    layer4_outputs(2939) <= a or b;
    layer4_outputs(2940) <= a;
    layer4_outputs(2941) <= not (a xor b);
    layer4_outputs(2942) <= a and not b;
    layer4_outputs(2943) <= not b;
    layer4_outputs(2944) <= a;
    layer4_outputs(2945) <= b;
    layer4_outputs(2946) <= a and not b;
    layer4_outputs(2947) <= a and b;
    layer4_outputs(2948) <= b;
    layer4_outputs(2949) <= b;
    layer4_outputs(2950) <= b and not a;
    layer4_outputs(2951) <= not a;
    layer4_outputs(2952) <= not a;
    layer4_outputs(2953) <= not (a or b);
    layer4_outputs(2954) <= a xor b;
    layer4_outputs(2955) <= a and not b;
    layer4_outputs(2956) <= '1';
    layer4_outputs(2957) <= not a;
    layer4_outputs(2958) <= a;
    layer4_outputs(2959) <= a and not b;
    layer4_outputs(2960) <= a or b;
    layer4_outputs(2961) <= b;
    layer4_outputs(2962) <= a and not b;
    layer4_outputs(2963) <= a xor b;
    layer4_outputs(2964) <= a;
    layer4_outputs(2965) <= b and not a;
    layer4_outputs(2966) <= not b or a;
    layer4_outputs(2967) <= a and b;
    layer4_outputs(2968) <= b;
    layer4_outputs(2969) <= b;
    layer4_outputs(2970) <= not a;
    layer4_outputs(2971) <= b;
    layer4_outputs(2972) <= not b or a;
    layer4_outputs(2973) <= not a;
    layer4_outputs(2974) <= not b;
    layer4_outputs(2975) <= not (a xor b);
    layer4_outputs(2976) <= not (a and b);
    layer4_outputs(2977) <= not (a or b);
    layer4_outputs(2978) <= not (a or b);
    layer4_outputs(2979) <= a or b;
    layer4_outputs(2980) <= b;
    layer4_outputs(2981) <= b and not a;
    layer4_outputs(2982) <= a and b;
    layer4_outputs(2983) <= a xor b;
    layer4_outputs(2984) <= not b or a;
    layer4_outputs(2985) <= not (a or b);
    layer4_outputs(2986) <= a and b;
    layer4_outputs(2987) <= not b;
    layer4_outputs(2988) <= not a or b;
    layer4_outputs(2989) <= not (a and b);
    layer4_outputs(2990) <= not (a xor b);
    layer4_outputs(2991) <= a and not b;
    layer4_outputs(2992) <= b;
    layer4_outputs(2993) <= a and not b;
    layer4_outputs(2994) <= not (a and b);
    layer4_outputs(2995) <= not a or b;
    layer4_outputs(2996) <= not b;
    layer4_outputs(2997) <= not a;
    layer4_outputs(2998) <= a;
    layer4_outputs(2999) <= a;
    layer4_outputs(3000) <= b;
    layer4_outputs(3001) <= a;
    layer4_outputs(3002) <= a xor b;
    layer4_outputs(3003) <= '1';
    layer4_outputs(3004) <= not b or a;
    layer4_outputs(3005) <= not (a or b);
    layer4_outputs(3006) <= a or b;
    layer4_outputs(3007) <= b;
    layer4_outputs(3008) <= not a or b;
    layer4_outputs(3009) <= not b;
    layer4_outputs(3010) <= not b or a;
    layer4_outputs(3011) <= not (a or b);
    layer4_outputs(3012) <= not b;
    layer4_outputs(3013) <= a xor b;
    layer4_outputs(3014) <= not b;
    layer4_outputs(3015) <= not (a or b);
    layer4_outputs(3016) <= b;
    layer4_outputs(3017) <= not (a and b);
    layer4_outputs(3018) <= not (a xor b);
    layer4_outputs(3019) <= not (a xor b);
    layer4_outputs(3020) <= b and not a;
    layer4_outputs(3021) <= not (a or b);
    layer4_outputs(3022) <= b and not a;
    layer4_outputs(3023) <= b;
    layer4_outputs(3024) <= not b;
    layer4_outputs(3025) <= a and not b;
    layer4_outputs(3026) <= a or b;
    layer4_outputs(3027) <= not a;
    layer4_outputs(3028) <= a;
    layer4_outputs(3029) <= not b or a;
    layer4_outputs(3030) <= b and not a;
    layer4_outputs(3031) <= a or b;
    layer4_outputs(3032) <= a;
    layer4_outputs(3033) <= '1';
    layer4_outputs(3034) <= a;
    layer4_outputs(3035) <= not (a and b);
    layer4_outputs(3036) <= a xor b;
    layer4_outputs(3037) <= not a;
    layer4_outputs(3038) <= a;
    layer4_outputs(3039) <= not a;
    layer4_outputs(3040) <= b and not a;
    layer4_outputs(3041) <= b;
    layer4_outputs(3042) <= not (a and b);
    layer4_outputs(3043) <= not a or b;
    layer4_outputs(3044) <= not a;
    layer4_outputs(3045) <= a and not b;
    layer4_outputs(3046) <= not (a and b);
    layer4_outputs(3047) <= b and not a;
    layer4_outputs(3048) <= not (a and b);
    layer4_outputs(3049) <= not a or b;
    layer4_outputs(3050) <= a and not b;
    layer4_outputs(3051) <= a xor b;
    layer4_outputs(3052) <= not a;
    layer4_outputs(3053) <= b and not a;
    layer4_outputs(3054) <= a;
    layer4_outputs(3055) <= a and not b;
    layer4_outputs(3056) <= a and not b;
    layer4_outputs(3057) <= b;
    layer4_outputs(3058) <= not (a and b);
    layer4_outputs(3059) <= not b or a;
    layer4_outputs(3060) <= not b;
    layer4_outputs(3061) <= not b or a;
    layer4_outputs(3062) <= a and b;
    layer4_outputs(3063) <= not a or b;
    layer4_outputs(3064) <= b;
    layer4_outputs(3065) <= b and not a;
    layer4_outputs(3066) <= not (a and b);
    layer4_outputs(3067) <= not b;
    layer4_outputs(3068) <= '0';
    layer4_outputs(3069) <= a and not b;
    layer4_outputs(3070) <= b;
    layer4_outputs(3071) <= not a;
    layer4_outputs(3072) <= not (a xor b);
    layer4_outputs(3073) <= not (a or b);
    layer4_outputs(3074) <= not (a and b);
    layer4_outputs(3075) <= not b;
    layer4_outputs(3076) <= not a;
    layer4_outputs(3077) <= a or b;
    layer4_outputs(3078) <= not b or a;
    layer4_outputs(3079) <= not (a xor b);
    layer4_outputs(3080) <= a xor b;
    layer4_outputs(3081) <= not (a or b);
    layer4_outputs(3082) <= not a or b;
    layer4_outputs(3083) <= not b;
    layer4_outputs(3084) <= not (a or b);
    layer4_outputs(3085) <= not a;
    layer4_outputs(3086) <= not b;
    layer4_outputs(3087) <= not b;
    layer4_outputs(3088) <= not a;
    layer4_outputs(3089) <= a and b;
    layer4_outputs(3090) <= b;
    layer4_outputs(3091) <= not b or a;
    layer4_outputs(3092) <= not b;
    layer4_outputs(3093) <= a;
    layer4_outputs(3094) <= '1';
    layer4_outputs(3095) <= not (a and b);
    layer4_outputs(3096) <= a xor b;
    layer4_outputs(3097) <= not a;
    layer4_outputs(3098) <= not b or a;
    layer4_outputs(3099) <= not b;
    layer4_outputs(3100) <= a and b;
    layer4_outputs(3101) <= not b;
    layer4_outputs(3102) <= a;
    layer4_outputs(3103) <= not (a xor b);
    layer4_outputs(3104) <= not a;
    layer4_outputs(3105) <= not a;
    layer4_outputs(3106) <= not (a xor b);
    layer4_outputs(3107) <= not b or a;
    layer4_outputs(3108) <= b;
    layer4_outputs(3109) <= a or b;
    layer4_outputs(3110) <= not a;
    layer4_outputs(3111) <= not (a and b);
    layer4_outputs(3112) <= not b;
    layer4_outputs(3113) <= not (a xor b);
    layer4_outputs(3114) <= not (a and b);
    layer4_outputs(3115) <= not (a and b);
    layer4_outputs(3116) <= not a;
    layer4_outputs(3117) <= a;
    layer4_outputs(3118) <= not b;
    layer4_outputs(3119) <= '0';
    layer4_outputs(3120) <= '1';
    layer4_outputs(3121) <= not (a xor b);
    layer4_outputs(3122) <= a xor b;
    layer4_outputs(3123) <= not a;
    layer4_outputs(3124) <= not b or a;
    layer4_outputs(3125) <= a or b;
    layer4_outputs(3126) <= not (a xor b);
    layer4_outputs(3127) <= a xor b;
    layer4_outputs(3128) <= b and not a;
    layer4_outputs(3129) <= a and not b;
    layer4_outputs(3130) <= a;
    layer4_outputs(3131) <= not b;
    layer4_outputs(3132) <= '1';
    layer4_outputs(3133) <= not b or a;
    layer4_outputs(3134) <= a xor b;
    layer4_outputs(3135) <= a and not b;
    layer4_outputs(3136) <= not (a or b);
    layer4_outputs(3137) <= a;
    layer4_outputs(3138) <= not (a and b);
    layer4_outputs(3139) <= not (a xor b);
    layer4_outputs(3140) <= not b or a;
    layer4_outputs(3141) <= not a or b;
    layer4_outputs(3142) <= b;
    layer4_outputs(3143) <= not (a xor b);
    layer4_outputs(3144) <= not (a and b);
    layer4_outputs(3145) <= not a or b;
    layer4_outputs(3146) <= not (a or b);
    layer4_outputs(3147) <= not b;
    layer4_outputs(3148) <= '0';
    layer4_outputs(3149) <= not b or a;
    layer4_outputs(3150) <= a and b;
    layer4_outputs(3151) <= not a;
    layer4_outputs(3152) <= b;
    layer4_outputs(3153) <= '1';
    layer4_outputs(3154) <= not (a and b);
    layer4_outputs(3155) <= a;
    layer4_outputs(3156) <= not (a and b);
    layer4_outputs(3157) <= a and not b;
    layer4_outputs(3158) <= a and not b;
    layer4_outputs(3159) <= a;
    layer4_outputs(3160) <= b;
    layer4_outputs(3161) <= a or b;
    layer4_outputs(3162) <= not a;
    layer4_outputs(3163) <= not b or a;
    layer4_outputs(3164) <= not b or a;
    layer4_outputs(3165) <= not b;
    layer4_outputs(3166) <= not a;
    layer4_outputs(3167) <= not b or a;
    layer4_outputs(3168) <= b and not a;
    layer4_outputs(3169) <= a or b;
    layer4_outputs(3170) <= a;
    layer4_outputs(3171) <= not b;
    layer4_outputs(3172) <= '0';
    layer4_outputs(3173) <= not (a xor b);
    layer4_outputs(3174) <= b and not a;
    layer4_outputs(3175) <= '1';
    layer4_outputs(3176) <= b and not a;
    layer4_outputs(3177) <= not b;
    layer4_outputs(3178) <= not (a and b);
    layer4_outputs(3179) <= not a;
    layer4_outputs(3180) <= not a;
    layer4_outputs(3181) <= not a or b;
    layer4_outputs(3182) <= not a;
    layer4_outputs(3183) <= b;
    layer4_outputs(3184) <= not a;
    layer4_outputs(3185) <= not a;
    layer4_outputs(3186) <= not (a and b);
    layer4_outputs(3187) <= '0';
    layer4_outputs(3188) <= b and not a;
    layer4_outputs(3189) <= not b;
    layer4_outputs(3190) <= '1';
    layer4_outputs(3191) <= not (a and b);
    layer4_outputs(3192) <= not (a and b);
    layer4_outputs(3193) <= not (a or b);
    layer4_outputs(3194) <= b;
    layer4_outputs(3195) <= not (a or b);
    layer4_outputs(3196) <= not b;
    layer4_outputs(3197) <= b and not a;
    layer4_outputs(3198) <= not b;
    layer4_outputs(3199) <= not b;
    layer4_outputs(3200) <= a;
    layer4_outputs(3201) <= not (a or b);
    layer4_outputs(3202) <= a;
    layer4_outputs(3203) <= not b or a;
    layer4_outputs(3204) <= a and b;
    layer4_outputs(3205) <= not a;
    layer4_outputs(3206) <= a;
    layer4_outputs(3207) <= not (a or b);
    layer4_outputs(3208) <= a and b;
    layer4_outputs(3209) <= b;
    layer4_outputs(3210) <= not b;
    layer4_outputs(3211) <= a and not b;
    layer4_outputs(3212) <= a;
    layer4_outputs(3213) <= a and not b;
    layer4_outputs(3214) <= a;
    layer4_outputs(3215) <= b and not a;
    layer4_outputs(3216) <= not b;
    layer4_outputs(3217) <= not b or a;
    layer4_outputs(3218) <= not a or b;
    layer4_outputs(3219) <= b;
    layer4_outputs(3220) <= not (a xor b);
    layer4_outputs(3221) <= '1';
    layer4_outputs(3222) <= b and not a;
    layer4_outputs(3223) <= a xor b;
    layer4_outputs(3224) <= not a;
    layer4_outputs(3225) <= a;
    layer4_outputs(3226) <= not (a xor b);
    layer4_outputs(3227) <= a;
    layer4_outputs(3228) <= a;
    layer4_outputs(3229) <= a and not b;
    layer4_outputs(3230) <= b;
    layer4_outputs(3231) <= b and not a;
    layer4_outputs(3232) <= not a;
    layer4_outputs(3233) <= '0';
    layer4_outputs(3234) <= b;
    layer4_outputs(3235) <= '0';
    layer4_outputs(3236) <= not a;
    layer4_outputs(3237) <= a xor b;
    layer4_outputs(3238) <= not (a or b);
    layer4_outputs(3239) <= not a;
    layer4_outputs(3240) <= not (a and b);
    layer4_outputs(3241) <= a xor b;
    layer4_outputs(3242) <= a and not b;
    layer4_outputs(3243) <= not b;
    layer4_outputs(3244) <= not a;
    layer4_outputs(3245) <= a or b;
    layer4_outputs(3246) <= b;
    layer4_outputs(3247) <= b and not a;
    layer4_outputs(3248) <= '1';
    layer4_outputs(3249) <= not a or b;
    layer4_outputs(3250) <= not a;
    layer4_outputs(3251) <= not a;
    layer4_outputs(3252) <= not b;
    layer4_outputs(3253) <= a;
    layer4_outputs(3254) <= not b or a;
    layer4_outputs(3255) <= not a;
    layer4_outputs(3256) <= a or b;
    layer4_outputs(3257) <= not a;
    layer4_outputs(3258) <= a and b;
    layer4_outputs(3259) <= not b;
    layer4_outputs(3260) <= not (a xor b);
    layer4_outputs(3261) <= not (a or b);
    layer4_outputs(3262) <= not (a or b);
    layer4_outputs(3263) <= a;
    layer4_outputs(3264) <= not (a xor b);
    layer4_outputs(3265) <= b and not a;
    layer4_outputs(3266) <= not b;
    layer4_outputs(3267) <= not (a or b);
    layer4_outputs(3268) <= a xor b;
    layer4_outputs(3269) <= not a;
    layer4_outputs(3270) <= a;
    layer4_outputs(3271) <= a xor b;
    layer4_outputs(3272) <= b;
    layer4_outputs(3273) <= a and b;
    layer4_outputs(3274) <= not b;
    layer4_outputs(3275) <= a xor b;
    layer4_outputs(3276) <= not b or a;
    layer4_outputs(3277) <= not a;
    layer4_outputs(3278) <= not b;
    layer4_outputs(3279) <= b;
    layer4_outputs(3280) <= not a;
    layer4_outputs(3281) <= not b or a;
    layer4_outputs(3282) <= a and b;
    layer4_outputs(3283) <= not a;
    layer4_outputs(3284) <= b and not a;
    layer4_outputs(3285) <= not a;
    layer4_outputs(3286) <= a or b;
    layer4_outputs(3287) <= not a;
    layer4_outputs(3288) <= a xor b;
    layer4_outputs(3289) <= not (a xor b);
    layer4_outputs(3290) <= b;
    layer4_outputs(3291) <= not b or a;
    layer4_outputs(3292) <= a;
    layer4_outputs(3293) <= not (a xor b);
    layer4_outputs(3294) <= not a or b;
    layer4_outputs(3295) <= not b or a;
    layer4_outputs(3296) <= a or b;
    layer4_outputs(3297) <= b;
    layer4_outputs(3298) <= a;
    layer4_outputs(3299) <= '1';
    layer4_outputs(3300) <= not (a or b);
    layer4_outputs(3301) <= not a or b;
    layer4_outputs(3302) <= not a;
    layer4_outputs(3303) <= not b;
    layer4_outputs(3304) <= a or b;
    layer4_outputs(3305) <= not (a and b);
    layer4_outputs(3306) <= not a;
    layer4_outputs(3307) <= b and not a;
    layer4_outputs(3308) <= b;
    layer4_outputs(3309) <= b;
    layer4_outputs(3310) <= a;
    layer4_outputs(3311) <= b;
    layer4_outputs(3312) <= a or b;
    layer4_outputs(3313) <= a and not b;
    layer4_outputs(3314) <= b;
    layer4_outputs(3315) <= not (a or b);
    layer4_outputs(3316) <= not a or b;
    layer4_outputs(3317) <= not a or b;
    layer4_outputs(3318) <= not a or b;
    layer4_outputs(3319) <= a xor b;
    layer4_outputs(3320) <= a xor b;
    layer4_outputs(3321) <= a;
    layer4_outputs(3322) <= not b;
    layer4_outputs(3323) <= not a or b;
    layer4_outputs(3324) <= not a;
    layer4_outputs(3325) <= a xor b;
    layer4_outputs(3326) <= a or b;
    layer4_outputs(3327) <= '1';
    layer4_outputs(3328) <= a and b;
    layer4_outputs(3329) <= not a;
    layer4_outputs(3330) <= b;
    layer4_outputs(3331) <= not b;
    layer4_outputs(3332) <= a;
    layer4_outputs(3333) <= a and b;
    layer4_outputs(3334) <= not a;
    layer4_outputs(3335) <= b;
    layer4_outputs(3336) <= a or b;
    layer4_outputs(3337) <= a and b;
    layer4_outputs(3338) <= b;
    layer4_outputs(3339) <= not b or a;
    layer4_outputs(3340) <= a and not b;
    layer4_outputs(3341) <= not b;
    layer4_outputs(3342) <= a;
    layer4_outputs(3343) <= a;
    layer4_outputs(3344) <= a and not b;
    layer4_outputs(3345) <= a;
    layer4_outputs(3346) <= a and b;
    layer4_outputs(3347) <= b;
    layer4_outputs(3348) <= not (a xor b);
    layer4_outputs(3349) <= not b;
    layer4_outputs(3350) <= b;
    layer4_outputs(3351) <= not (a or b);
    layer4_outputs(3352) <= a or b;
    layer4_outputs(3353) <= a and b;
    layer4_outputs(3354) <= not b or a;
    layer4_outputs(3355) <= not a or b;
    layer4_outputs(3356) <= a xor b;
    layer4_outputs(3357) <= a;
    layer4_outputs(3358) <= not (a xor b);
    layer4_outputs(3359) <= a;
    layer4_outputs(3360) <= not (a or b);
    layer4_outputs(3361) <= a;
    layer4_outputs(3362) <= a and b;
    layer4_outputs(3363) <= a and b;
    layer4_outputs(3364) <= not a;
    layer4_outputs(3365) <= a;
    layer4_outputs(3366) <= not a or b;
    layer4_outputs(3367) <= not (a or b);
    layer4_outputs(3368) <= a;
    layer4_outputs(3369) <= a and not b;
    layer4_outputs(3370) <= a or b;
    layer4_outputs(3371) <= not (a or b);
    layer4_outputs(3372) <= not b;
    layer4_outputs(3373) <= not a;
    layer4_outputs(3374) <= not (a xor b);
    layer4_outputs(3375) <= b and not a;
    layer4_outputs(3376) <= not b;
    layer4_outputs(3377) <= not b;
    layer4_outputs(3378) <= a and not b;
    layer4_outputs(3379) <= not b;
    layer4_outputs(3380) <= not a;
    layer4_outputs(3381) <= not a or b;
    layer4_outputs(3382) <= not (a and b);
    layer4_outputs(3383) <= a or b;
    layer4_outputs(3384) <= not b;
    layer4_outputs(3385) <= not a;
    layer4_outputs(3386) <= not a or b;
    layer4_outputs(3387) <= not (a and b);
    layer4_outputs(3388) <= a or b;
    layer4_outputs(3389) <= not a or b;
    layer4_outputs(3390) <= a and b;
    layer4_outputs(3391) <= not a;
    layer4_outputs(3392) <= not a or b;
    layer4_outputs(3393) <= a or b;
    layer4_outputs(3394) <= not a;
    layer4_outputs(3395) <= not a or b;
    layer4_outputs(3396) <= a and not b;
    layer4_outputs(3397) <= a and not b;
    layer4_outputs(3398) <= a or b;
    layer4_outputs(3399) <= a and b;
    layer4_outputs(3400) <= a or b;
    layer4_outputs(3401) <= not b or a;
    layer4_outputs(3402) <= not b or a;
    layer4_outputs(3403) <= b;
    layer4_outputs(3404) <= a or b;
    layer4_outputs(3405) <= '1';
    layer4_outputs(3406) <= not b or a;
    layer4_outputs(3407) <= not b;
    layer4_outputs(3408) <= b;
    layer4_outputs(3409) <= '1';
    layer4_outputs(3410) <= a or b;
    layer4_outputs(3411) <= not a;
    layer4_outputs(3412) <= '0';
    layer4_outputs(3413) <= not a or b;
    layer4_outputs(3414) <= not b;
    layer4_outputs(3415) <= a xor b;
    layer4_outputs(3416) <= not (a or b);
    layer4_outputs(3417) <= a and not b;
    layer4_outputs(3418) <= a;
    layer4_outputs(3419) <= b;
    layer4_outputs(3420) <= not (a xor b);
    layer4_outputs(3421) <= not a;
    layer4_outputs(3422) <= a and b;
    layer4_outputs(3423) <= a;
    layer4_outputs(3424) <= not b;
    layer4_outputs(3425) <= not b;
    layer4_outputs(3426) <= a or b;
    layer4_outputs(3427) <= b;
    layer4_outputs(3428) <= not (a xor b);
    layer4_outputs(3429) <= not b or a;
    layer4_outputs(3430) <= not a or b;
    layer4_outputs(3431) <= not b;
    layer4_outputs(3432) <= not b or a;
    layer4_outputs(3433) <= not b or a;
    layer4_outputs(3434) <= not (a or b);
    layer4_outputs(3435) <= not a;
    layer4_outputs(3436) <= b;
    layer4_outputs(3437) <= b;
    layer4_outputs(3438) <= not b;
    layer4_outputs(3439) <= not (a and b);
    layer4_outputs(3440) <= not a or b;
    layer4_outputs(3441) <= not a or b;
    layer4_outputs(3442) <= not a or b;
    layer4_outputs(3443) <= not b or a;
    layer4_outputs(3444) <= not (a or b);
    layer4_outputs(3445) <= '0';
    layer4_outputs(3446) <= a xor b;
    layer4_outputs(3447) <= a and b;
    layer4_outputs(3448) <= not a;
    layer4_outputs(3449) <= not (a and b);
    layer4_outputs(3450) <= a and b;
    layer4_outputs(3451) <= not b or a;
    layer4_outputs(3452) <= not b or a;
    layer4_outputs(3453) <= b;
    layer4_outputs(3454) <= b;
    layer4_outputs(3455) <= not (a xor b);
    layer4_outputs(3456) <= a;
    layer4_outputs(3457) <= '0';
    layer4_outputs(3458) <= b and not a;
    layer4_outputs(3459) <= a xor b;
    layer4_outputs(3460) <= a and not b;
    layer4_outputs(3461) <= not b or a;
    layer4_outputs(3462) <= a;
    layer4_outputs(3463) <= not b;
    layer4_outputs(3464) <= a;
    layer4_outputs(3465) <= a or b;
    layer4_outputs(3466) <= not (a and b);
    layer4_outputs(3467) <= not (a and b);
    layer4_outputs(3468) <= not b or a;
    layer4_outputs(3469) <= b;
    layer4_outputs(3470) <= b;
    layer4_outputs(3471) <= not b;
    layer4_outputs(3472) <= b and not a;
    layer4_outputs(3473) <= a and not b;
    layer4_outputs(3474) <= not (a xor b);
    layer4_outputs(3475) <= a;
    layer4_outputs(3476) <= not b;
    layer4_outputs(3477) <= a xor b;
    layer4_outputs(3478) <= not b;
    layer4_outputs(3479) <= b and not a;
    layer4_outputs(3480) <= not a or b;
    layer4_outputs(3481) <= not b;
    layer4_outputs(3482) <= a;
    layer4_outputs(3483) <= b;
    layer4_outputs(3484) <= '0';
    layer4_outputs(3485) <= not b or a;
    layer4_outputs(3486) <= not (a or b);
    layer4_outputs(3487) <= b;
    layer4_outputs(3488) <= b and not a;
    layer4_outputs(3489) <= not (a or b);
    layer4_outputs(3490) <= a xor b;
    layer4_outputs(3491) <= not b or a;
    layer4_outputs(3492) <= not b;
    layer4_outputs(3493) <= b;
    layer4_outputs(3494) <= not a or b;
    layer4_outputs(3495) <= a xor b;
    layer4_outputs(3496) <= b and not a;
    layer4_outputs(3497) <= not b;
    layer4_outputs(3498) <= not b;
    layer4_outputs(3499) <= a and not b;
    layer4_outputs(3500) <= a and b;
    layer4_outputs(3501) <= b;
    layer4_outputs(3502) <= not b or a;
    layer4_outputs(3503) <= a;
    layer4_outputs(3504) <= b and not a;
    layer4_outputs(3505) <= b;
    layer4_outputs(3506) <= a;
    layer4_outputs(3507) <= a and not b;
    layer4_outputs(3508) <= b;
    layer4_outputs(3509) <= not a;
    layer4_outputs(3510) <= b and not a;
    layer4_outputs(3511) <= not b or a;
    layer4_outputs(3512) <= not b;
    layer4_outputs(3513) <= not a or b;
    layer4_outputs(3514) <= '1';
    layer4_outputs(3515) <= not a;
    layer4_outputs(3516) <= not (a and b);
    layer4_outputs(3517) <= a;
    layer4_outputs(3518) <= a and not b;
    layer4_outputs(3519) <= not (a or b);
    layer4_outputs(3520) <= a xor b;
    layer4_outputs(3521) <= not b;
    layer4_outputs(3522) <= not a;
    layer4_outputs(3523) <= b;
    layer4_outputs(3524) <= not (a or b);
    layer4_outputs(3525) <= a and not b;
    layer4_outputs(3526) <= not (a and b);
    layer4_outputs(3527) <= not a;
    layer4_outputs(3528) <= not (a and b);
    layer4_outputs(3529) <= a and not b;
    layer4_outputs(3530) <= b and not a;
    layer4_outputs(3531) <= not b;
    layer4_outputs(3532) <= not (a and b);
    layer4_outputs(3533) <= not (a or b);
    layer4_outputs(3534) <= not a;
    layer4_outputs(3535) <= not a;
    layer4_outputs(3536) <= not a;
    layer4_outputs(3537) <= not b;
    layer4_outputs(3538) <= a and b;
    layer4_outputs(3539) <= a;
    layer4_outputs(3540) <= a xor b;
    layer4_outputs(3541) <= a;
    layer4_outputs(3542) <= a;
    layer4_outputs(3543) <= not b;
    layer4_outputs(3544) <= a and b;
    layer4_outputs(3545) <= a and not b;
    layer4_outputs(3546) <= not (a and b);
    layer4_outputs(3547) <= a and not b;
    layer4_outputs(3548) <= not a or b;
    layer4_outputs(3549) <= b;
    layer4_outputs(3550) <= a and b;
    layer4_outputs(3551) <= a and b;
    layer4_outputs(3552) <= not b;
    layer4_outputs(3553) <= not a;
    layer4_outputs(3554) <= not a or b;
    layer4_outputs(3555) <= b;
    layer4_outputs(3556) <= not (a or b);
    layer4_outputs(3557) <= not a;
    layer4_outputs(3558) <= a and not b;
    layer4_outputs(3559) <= not b or a;
    layer4_outputs(3560) <= not a or b;
    layer4_outputs(3561) <= a;
    layer4_outputs(3562) <= not b or a;
    layer4_outputs(3563) <= not a;
    layer4_outputs(3564) <= not (a and b);
    layer4_outputs(3565) <= not a;
    layer4_outputs(3566) <= not a;
    layer4_outputs(3567) <= '1';
    layer4_outputs(3568) <= not (a or b);
    layer4_outputs(3569) <= not a;
    layer4_outputs(3570) <= not a;
    layer4_outputs(3571) <= not (a and b);
    layer4_outputs(3572) <= a xor b;
    layer4_outputs(3573) <= not (a and b);
    layer4_outputs(3574) <= a xor b;
    layer4_outputs(3575) <= '1';
    layer4_outputs(3576) <= not (a or b);
    layer4_outputs(3577) <= not b or a;
    layer4_outputs(3578) <= a or b;
    layer4_outputs(3579) <= not (a and b);
    layer4_outputs(3580) <= not a;
    layer4_outputs(3581) <= a;
    layer4_outputs(3582) <= b and not a;
    layer4_outputs(3583) <= not b;
    layer4_outputs(3584) <= b;
    layer4_outputs(3585) <= a xor b;
    layer4_outputs(3586) <= not b;
    layer4_outputs(3587) <= a;
    layer4_outputs(3588) <= b and not a;
    layer4_outputs(3589) <= a;
    layer4_outputs(3590) <= not b;
    layer4_outputs(3591) <= a xor b;
    layer4_outputs(3592) <= b;
    layer4_outputs(3593) <= not b or a;
    layer4_outputs(3594) <= not b or a;
    layer4_outputs(3595) <= '1';
    layer4_outputs(3596) <= not b;
    layer4_outputs(3597) <= not (a xor b);
    layer4_outputs(3598) <= b;
    layer4_outputs(3599) <= not b;
    layer4_outputs(3600) <= not b or a;
    layer4_outputs(3601) <= not (a or b);
    layer4_outputs(3602) <= a xor b;
    layer4_outputs(3603) <= '1';
    layer4_outputs(3604) <= not (a or b);
    layer4_outputs(3605) <= b and not a;
    layer4_outputs(3606) <= a or b;
    layer4_outputs(3607) <= not (a or b);
    layer4_outputs(3608) <= a xor b;
    layer4_outputs(3609) <= not (a xor b);
    layer4_outputs(3610) <= a;
    layer4_outputs(3611) <= a or b;
    layer4_outputs(3612) <= a and b;
    layer4_outputs(3613) <= not (a and b);
    layer4_outputs(3614) <= not b;
    layer4_outputs(3615) <= not (a xor b);
    layer4_outputs(3616) <= not (a and b);
    layer4_outputs(3617) <= a and not b;
    layer4_outputs(3618) <= not a;
    layer4_outputs(3619) <= not a or b;
    layer4_outputs(3620) <= not (a or b);
    layer4_outputs(3621) <= b;
    layer4_outputs(3622) <= not (a and b);
    layer4_outputs(3623) <= a;
    layer4_outputs(3624) <= not b or a;
    layer4_outputs(3625) <= not (a and b);
    layer4_outputs(3626) <= not a;
    layer4_outputs(3627) <= a xor b;
    layer4_outputs(3628) <= not (a or b);
    layer4_outputs(3629) <= a and b;
    layer4_outputs(3630) <= '0';
    layer4_outputs(3631) <= a or b;
    layer4_outputs(3632) <= not a;
    layer4_outputs(3633) <= '0';
    layer4_outputs(3634) <= not (a xor b);
    layer4_outputs(3635) <= a xor b;
    layer4_outputs(3636) <= not a or b;
    layer4_outputs(3637) <= b;
    layer4_outputs(3638) <= not (a xor b);
    layer4_outputs(3639) <= b and not a;
    layer4_outputs(3640) <= not (a and b);
    layer4_outputs(3641) <= not a;
    layer4_outputs(3642) <= not (a and b);
    layer4_outputs(3643) <= b and not a;
    layer4_outputs(3644) <= b;
    layer4_outputs(3645) <= a and b;
    layer4_outputs(3646) <= b and not a;
    layer4_outputs(3647) <= '0';
    layer4_outputs(3648) <= not (a and b);
    layer4_outputs(3649) <= b and not a;
    layer4_outputs(3650) <= a or b;
    layer4_outputs(3651) <= not a;
    layer4_outputs(3652) <= a xor b;
    layer4_outputs(3653) <= a or b;
    layer4_outputs(3654) <= a and b;
    layer4_outputs(3655) <= a;
    layer4_outputs(3656) <= not b;
    layer4_outputs(3657) <= b;
    layer4_outputs(3658) <= not (a xor b);
    layer4_outputs(3659) <= a and b;
    layer4_outputs(3660) <= not (a or b);
    layer4_outputs(3661) <= '0';
    layer4_outputs(3662) <= not (a and b);
    layer4_outputs(3663) <= not a or b;
    layer4_outputs(3664) <= not (a xor b);
    layer4_outputs(3665) <= a and not b;
    layer4_outputs(3666) <= b and not a;
    layer4_outputs(3667) <= not a;
    layer4_outputs(3668) <= not (a or b);
    layer4_outputs(3669) <= not (a or b);
    layer4_outputs(3670) <= not (a or b);
    layer4_outputs(3671) <= not (a and b);
    layer4_outputs(3672) <= not a or b;
    layer4_outputs(3673) <= b;
    layer4_outputs(3674) <= '1';
    layer4_outputs(3675) <= not b;
    layer4_outputs(3676) <= b and not a;
    layer4_outputs(3677) <= b;
    layer4_outputs(3678) <= not b;
    layer4_outputs(3679) <= b;
    layer4_outputs(3680) <= a;
    layer4_outputs(3681) <= not b;
    layer4_outputs(3682) <= a;
    layer4_outputs(3683) <= b and not a;
    layer4_outputs(3684) <= not (a and b);
    layer4_outputs(3685) <= not b;
    layer4_outputs(3686) <= not b;
    layer4_outputs(3687) <= not b or a;
    layer4_outputs(3688) <= a;
    layer4_outputs(3689) <= a xor b;
    layer4_outputs(3690) <= not a;
    layer4_outputs(3691) <= not (a and b);
    layer4_outputs(3692) <= a;
    layer4_outputs(3693) <= a and b;
    layer4_outputs(3694) <= a and not b;
    layer4_outputs(3695) <= b and not a;
    layer4_outputs(3696) <= not a;
    layer4_outputs(3697) <= b and not a;
    layer4_outputs(3698) <= a;
    layer4_outputs(3699) <= a and b;
    layer4_outputs(3700) <= not b;
    layer4_outputs(3701) <= a;
    layer4_outputs(3702) <= not (a and b);
    layer4_outputs(3703) <= a;
    layer4_outputs(3704) <= not b or a;
    layer4_outputs(3705) <= not (a or b);
    layer4_outputs(3706) <= not (a xor b);
    layer4_outputs(3707) <= b;
    layer4_outputs(3708) <= not a;
    layer4_outputs(3709) <= a;
    layer4_outputs(3710) <= not (a and b);
    layer4_outputs(3711) <= a or b;
    layer4_outputs(3712) <= not a;
    layer4_outputs(3713) <= not (a xor b);
    layer4_outputs(3714) <= b and not a;
    layer4_outputs(3715) <= a;
    layer4_outputs(3716) <= a or b;
    layer4_outputs(3717) <= '0';
    layer4_outputs(3718) <= b;
    layer4_outputs(3719) <= not (a and b);
    layer4_outputs(3720) <= not b or a;
    layer4_outputs(3721) <= b;
    layer4_outputs(3722) <= not a;
    layer4_outputs(3723) <= not b or a;
    layer4_outputs(3724) <= b;
    layer4_outputs(3725) <= a;
    layer4_outputs(3726) <= not b;
    layer4_outputs(3727) <= not (a and b);
    layer4_outputs(3728) <= not b;
    layer4_outputs(3729) <= not b;
    layer4_outputs(3730) <= a;
    layer4_outputs(3731) <= not (a xor b);
    layer4_outputs(3732) <= a or b;
    layer4_outputs(3733) <= b and not a;
    layer4_outputs(3734) <= not a;
    layer4_outputs(3735) <= not b;
    layer4_outputs(3736) <= a;
    layer4_outputs(3737) <= not b or a;
    layer4_outputs(3738) <= b and not a;
    layer4_outputs(3739) <= '1';
    layer4_outputs(3740) <= a and not b;
    layer4_outputs(3741) <= not (a or b);
    layer4_outputs(3742) <= not a or b;
    layer4_outputs(3743) <= a;
    layer4_outputs(3744) <= a or b;
    layer4_outputs(3745) <= a and not b;
    layer4_outputs(3746) <= not b;
    layer4_outputs(3747) <= a;
    layer4_outputs(3748) <= a and not b;
    layer4_outputs(3749) <= b and not a;
    layer4_outputs(3750) <= not (a xor b);
    layer4_outputs(3751) <= not (a xor b);
    layer4_outputs(3752) <= not (a or b);
    layer4_outputs(3753) <= not (a or b);
    layer4_outputs(3754) <= a and b;
    layer4_outputs(3755) <= a or b;
    layer4_outputs(3756) <= a;
    layer4_outputs(3757) <= a xor b;
    layer4_outputs(3758) <= not a;
    layer4_outputs(3759) <= not b or a;
    layer4_outputs(3760) <= a and b;
    layer4_outputs(3761) <= b and not a;
    layer4_outputs(3762) <= not b;
    layer4_outputs(3763) <= '0';
    layer4_outputs(3764) <= a and b;
    layer4_outputs(3765) <= b;
    layer4_outputs(3766) <= a xor b;
    layer4_outputs(3767) <= not b;
    layer4_outputs(3768) <= not b or a;
    layer4_outputs(3769) <= a and b;
    layer4_outputs(3770) <= b;
    layer4_outputs(3771) <= b;
    layer4_outputs(3772) <= a and b;
    layer4_outputs(3773) <= b and not a;
    layer4_outputs(3774) <= not (a and b);
    layer4_outputs(3775) <= a;
    layer4_outputs(3776) <= '0';
    layer4_outputs(3777) <= a or b;
    layer4_outputs(3778) <= not b;
    layer4_outputs(3779) <= not b or a;
    layer4_outputs(3780) <= not b or a;
    layer4_outputs(3781) <= a;
    layer4_outputs(3782) <= b and not a;
    layer4_outputs(3783) <= b;
    layer4_outputs(3784) <= a xor b;
    layer4_outputs(3785) <= b and not a;
    layer4_outputs(3786) <= a xor b;
    layer4_outputs(3787) <= b;
    layer4_outputs(3788) <= not (a and b);
    layer4_outputs(3789) <= not (a xor b);
    layer4_outputs(3790) <= a;
    layer4_outputs(3791) <= not b;
    layer4_outputs(3792) <= not (a xor b);
    layer4_outputs(3793) <= not a;
    layer4_outputs(3794) <= a;
    layer4_outputs(3795) <= not (a and b);
    layer4_outputs(3796) <= not a;
    layer4_outputs(3797) <= not a;
    layer4_outputs(3798) <= not (a xor b);
    layer4_outputs(3799) <= '1';
    layer4_outputs(3800) <= not b or a;
    layer4_outputs(3801) <= a;
    layer4_outputs(3802) <= not b;
    layer4_outputs(3803) <= not (a or b);
    layer4_outputs(3804) <= b and not a;
    layer4_outputs(3805) <= not b;
    layer4_outputs(3806) <= a and not b;
    layer4_outputs(3807) <= a;
    layer4_outputs(3808) <= not b;
    layer4_outputs(3809) <= a;
    layer4_outputs(3810) <= a xor b;
    layer4_outputs(3811) <= a or b;
    layer4_outputs(3812) <= not (a xor b);
    layer4_outputs(3813) <= a;
    layer4_outputs(3814) <= not (a or b);
    layer4_outputs(3815) <= a and not b;
    layer4_outputs(3816) <= a xor b;
    layer4_outputs(3817) <= not b or a;
    layer4_outputs(3818) <= a and b;
    layer4_outputs(3819) <= b;
    layer4_outputs(3820) <= a xor b;
    layer4_outputs(3821) <= not b;
    layer4_outputs(3822) <= a;
    layer4_outputs(3823) <= a or b;
    layer4_outputs(3824) <= not a or b;
    layer4_outputs(3825) <= a or b;
    layer4_outputs(3826) <= a and b;
    layer4_outputs(3827) <= a;
    layer4_outputs(3828) <= b;
    layer4_outputs(3829) <= not b;
    layer4_outputs(3830) <= not b or a;
    layer4_outputs(3831) <= a;
    layer4_outputs(3832) <= a and not b;
    layer4_outputs(3833) <= not (a and b);
    layer4_outputs(3834) <= a or b;
    layer4_outputs(3835) <= b;
    layer4_outputs(3836) <= b and not a;
    layer4_outputs(3837) <= a and not b;
    layer4_outputs(3838) <= not b;
    layer4_outputs(3839) <= not (a or b);
    layer4_outputs(3840) <= not (a xor b);
    layer4_outputs(3841) <= a and not b;
    layer4_outputs(3842) <= b and not a;
    layer4_outputs(3843) <= not b;
    layer4_outputs(3844) <= not (a xor b);
    layer4_outputs(3845) <= not b or a;
    layer4_outputs(3846) <= not (a or b);
    layer4_outputs(3847) <= not (a and b);
    layer4_outputs(3848) <= a and b;
    layer4_outputs(3849) <= not (a xor b);
    layer4_outputs(3850) <= not (a or b);
    layer4_outputs(3851) <= a;
    layer4_outputs(3852) <= b and not a;
    layer4_outputs(3853) <= not (a and b);
    layer4_outputs(3854) <= a and not b;
    layer4_outputs(3855) <= not (a or b);
    layer4_outputs(3856) <= b and not a;
    layer4_outputs(3857) <= a xor b;
    layer4_outputs(3858) <= not b;
    layer4_outputs(3859) <= a;
    layer4_outputs(3860) <= b;
    layer4_outputs(3861) <= a and not b;
    layer4_outputs(3862) <= a and not b;
    layer4_outputs(3863) <= not b;
    layer4_outputs(3864) <= not a;
    layer4_outputs(3865) <= not (a xor b);
    layer4_outputs(3866) <= a xor b;
    layer4_outputs(3867) <= not b or a;
    layer4_outputs(3868) <= a or b;
    layer4_outputs(3869) <= not a or b;
    layer4_outputs(3870) <= not (a or b);
    layer4_outputs(3871) <= not (a or b);
    layer4_outputs(3872) <= not (a and b);
    layer4_outputs(3873) <= not a;
    layer4_outputs(3874) <= not a;
    layer4_outputs(3875) <= a and b;
    layer4_outputs(3876) <= not b;
    layer4_outputs(3877) <= not a;
    layer4_outputs(3878) <= a;
    layer4_outputs(3879) <= a and b;
    layer4_outputs(3880) <= not b;
    layer4_outputs(3881) <= a;
    layer4_outputs(3882) <= a or b;
    layer4_outputs(3883) <= not (a xor b);
    layer4_outputs(3884) <= not a or b;
    layer4_outputs(3885) <= '0';
    layer4_outputs(3886) <= b;
    layer4_outputs(3887) <= a or b;
    layer4_outputs(3888) <= a xor b;
    layer4_outputs(3889) <= a;
    layer4_outputs(3890) <= not (a xor b);
    layer4_outputs(3891) <= not (a and b);
    layer4_outputs(3892) <= not a or b;
    layer4_outputs(3893) <= a;
    layer4_outputs(3894) <= not a;
    layer4_outputs(3895) <= '0';
    layer4_outputs(3896) <= a and not b;
    layer4_outputs(3897) <= not a or b;
    layer4_outputs(3898) <= '0';
    layer4_outputs(3899) <= not (a xor b);
    layer4_outputs(3900) <= a;
    layer4_outputs(3901) <= not a or b;
    layer4_outputs(3902) <= a or b;
    layer4_outputs(3903) <= not (a or b);
    layer4_outputs(3904) <= not (a xor b);
    layer4_outputs(3905) <= b and not a;
    layer4_outputs(3906) <= not (a or b);
    layer4_outputs(3907) <= a or b;
    layer4_outputs(3908) <= not (a or b);
    layer4_outputs(3909) <= not b;
    layer4_outputs(3910) <= not b;
    layer4_outputs(3911) <= a;
    layer4_outputs(3912) <= b;
    layer4_outputs(3913) <= not b;
    layer4_outputs(3914) <= not (a xor b);
    layer4_outputs(3915) <= not a;
    layer4_outputs(3916) <= b;
    layer4_outputs(3917) <= '0';
    layer4_outputs(3918) <= a and b;
    layer4_outputs(3919) <= not b or a;
    layer4_outputs(3920) <= not b or a;
    layer4_outputs(3921) <= not a;
    layer4_outputs(3922) <= not (a or b);
    layer4_outputs(3923) <= a;
    layer4_outputs(3924) <= a or b;
    layer4_outputs(3925) <= a or b;
    layer4_outputs(3926) <= a and not b;
    layer4_outputs(3927) <= b and not a;
    layer4_outputs(3928) <= b;
    layer4_outputs(3929) <= a;
    layer4_outputs(3930) <= a and not b;
    layer4_outputs(3931) <= not a;
    layer4_outputs(3932) <= a or b;
    layer4_outputs(3933) <= not a or b;
    layer4_outputs(3934) <= not b;
    layer4_outputs(3935) <= not a;
    layer4_outputs(3936) <= not b or a;
    layer4_outputs(3937) <= b;
    layer4_outputs(3938) <= not a;
    layer4_outputs(3939) <= not (a or b);
    layer4_outputs(3940) <= not (a or b);
    layer4_outputs(3941) <= b and not a;
    layer4_outputs(3942) <= not a or b;
    layer4_outputs(3943) <= b and not a;
    layer4_outputs(3944) <= not b;
    layer4_outputs(3945) <= a or b;
    layer4_outputs(3946) <= a;
    layer4_outputs(3947) <= not (a or b);
    layer4_outputs(3948) <= a;
    layer4_outputs(3949) <= b;
    layer4_outputs(3950) <= not (a or b);
    layer4_outputs(3951) <= a;
    layer4_outputs(3952) <= b and not a;
    layer4_outputs(3953) <= not b or a;
    layer4_outputs(3954) <= b;
    layer4_outputs(3955) <= not b;
    layer4_outputs(3956) <= not b;
    layer4_outputs(3957) <= a or b;
    layer4_outputs(3958) <= not a or b;
    layer4_outputs(3959) <= not b;
    layer4_outputs(3960) <= not b;
    layer4_outputs(3961) <= not a or b;
    layer4_outputs(3962) <= '1';
    layer4_outputs(3963) <= not a;
    layer4_outputs(3964) <= not (a xor b);
    layer4_outputs(3965) <= not (a or b);
    layer4_outputs(3966) <= not (a or b);
    layer4_outputs(3967) <= not a;
    layer4_outputs(3968) <= a;
    layer4_outputs(3969) <= not b;
    layer4_outputs(3970) <= a or b;
    layer4_outputs(3971) <= not b;
    layer4_outputs(3972) <= a or b;
    layer4_outputs(3973) <= a;
    layer4_outputs(3974) <= not b or a;
    layer4_outputs(3975) <= not b or a;
    layer4_outputs(3976) <= a and b;
    layer4_outputs(3977) <= a;
    layer4_outputs(3978) <= a;
    layer4_outputs(3979) <= a xor b;
    layer4_outputs(3980) <= a and b;
    layer4_outputs(3981) <= a and b;
    layer4_outputs(3982) <= b;
    layer4_outputs(3983) <= a;
    layer4_outputs(3984) <= a;
    layer4_outputs(3985) <= b and not a;
    layer4_outputs(3986) <= b and not a;
    layer4_outputs(3987) <= a or b;
    layer4_outputs(3988) <= b;
    layer4_outputs(3989) <= a;
    layer4_outputs(3990) <= a and b;
    layer4_outputs(3991) <= not (a xor b);
    layer4_outputs(3992) <= a;
    layer4_outputs(3993) <= a or b;
    layer4_outputs(3994) <= not b;
    layer4_outputs(3995) <= a;
    layer4_outputs(3996) <= not a;
    layer4_outputs(3997) <= a and not b;
    layer4_outputs(3998) <= not b;
    layer4_outputs(3999) <= a and not b;
    layer4_outputs(4000) <= not (a xor b);
    layer4_outputs(4001) <= not b;
    layer4_outputs(4002) <= b;
    layer4_outputs(4003) <= b and not a;
    layer4_outputs(4004) <= a and b;
    layer4_outputs(4005) <= b and not a;
    layer4_outputs(4006) <= a;
    layer4_outputs(4007) <= b and not a;
    layer4_outputs(4008) <= '0';
    layer4_outputs(4009) <= not (a and b);
    layer4_outputs(4010) <= not (a and b);
    layer4_outputs(4011) <= not b or a;
    layer4_outputs(4012) <= '1';
    layer4_outputs(4013) <= b;
    layer4_outputs(4014) <= a;
    layer4_outputs(4015) <= not b;
    layer4_outputs(4016) <= '1';
    layer4_outputs(4017) <= not a;
    layer4_outputs(4018) <= b;
    layer4_outputs(4019) <= not b;
    layer4_outputs(4020) <= a xor b;
    layer4_outputs(4021) <= not a;
    layer4_outputs(4022) <= not a;
    layer4_outputs(4023) <= not a or b;
    layer4_outputs(4024) <= not a;
    layer4_outputs(4025) <= not (a and b);
    layer4_outputs(4026) <= not a or b;
    layer4_outputs(4027) <= a;
    layer4_outputs(4028) <= not (a xor b);
    layer4_outputs(4029) <= '0';
    layer4_outputs(4030) <= not b or a;
    layer4_outputs(4031) <= not b;
    layer4_outputs(4032) <= not a;
    layer4_outputs(4033) <= a and b;
    layer4_outputs(4034) <= not b or a;
    layer4_outputs(4035) <= not b;
    layer4_outputs(4036) <= not b;
    layer4_outputs(4037) <= not a;
    layer4_outputs(4038) <= not (a and b);
    layer4_outputs(4039) <= b;
    layer4_outputs(4040) <= a and b;
    layer4_outputs(4041) <= not b;
    layer4_outputs(4042) <= a and not b;
    layer4_outputs(4043) <= a;
    layer4_outputs(4044) <= not b;
    layer4_outputs(4045) <= not b;
    layer4_outputs(4046) <= not b;
    layer4_outputs(4047) <= a;
    layer4_outputs(4048) <= not (a or b);
    layer4_outputs(4049) <= not (a and b);
    layer4_outputs(4050) <= b;
    layer4_outputs(4051) <= not (a or b);
    layer4_outputs(4052) <= not a;
    layer4_outputs(4053) <= not b or a;
    layer4_outputs(4054) <= not b;
    layer4_outputs(4055) <= a;
    layer4_outputs(4056) <= a or b;
    layer4_outputs(4057) <= a and not b;
    layer4_outputs(4058) <= a;
    layer4_outputs(4059) <= not (a and b);
    layer4_outputs(4060) <= not b;
    layer4_outputs(4061) <= '1';
    layer4_outputs(4062) <= not (a or b);
    layer4_outputs(4063) <= not (a or b);
    layer4_outputs(4064) <= '0';
    layer4_outputs(4065) <= not (a xor b);
    layer4_outputs(4066) <= a xor b;
    layer4_outputs(4067) <= b and not a;
    layer4_outputs(4068) <= not (a or b);
    layer4_outputs(4069) <= '1';
    layer4_outputs(4070) <= a and b;
    layer4_outputs(4071) <= a or b;
    layer4_outputs(4072) <= a and b;
    layer4_outputs(4073) <= not a;
    layer4_outputs(4074) <= not b;
    layer4_outputs(4075) <= not a or b;
    layer4_outputs(4076) <= not (a or b);
    layer4_outputs(4077) <= not a or b;
    layer4_outputs(4078) <= not b or a;
    layer4_outputs(4079) <= not (a and b);
    layer4_outputs(4080) <= not (a or b);
    layer4_outputs(4081) <= a and b;
    layer4_outputs(4082) <= a and b;
    layer4_outputs(4083) <= not (a xor b);
    layer4_outputs(4084) <= b;
    layer4_outputs(4085) <= not b;
    layer4_outputs(4086) <= not a or b;
    layer4_outputs(4087) <= not a;
    layer4_outputs(4088) <= not b;
    layer4_outputs(4089) <= not b or a;
    layer4_outputs(4090) <= not (a and b);
    layer4_outputs(4091) <= b and not a;
    layer4_outputs(4092) <= a or b;
    layer4_outputs(4093) <= not a;
    layer4_outputs(4094) <= b;
    layer4_outputs(4095) <= not b;
    layer4_outputs(4096) <= b and not a;
    layer4_outputs(4097) <= b;
    layer4_outputs(4098) <= not (a or b);
    layer4_outputs(4099) <= a;
    layer4_outputs(4100) <= not (a or b);
    layer4_outputs(4101) <= a xor b;
    layer4_outputs(4102) <= '0';
    layer4_outputs(4103) <= not a;
    layer4_outputs(4104) <= not b;
    layer4_outputs(4105) <= not a;
    layer4_outputs(4106) <= a;
    layer4_outputs(4107) <= not b or a;
    layer4_outputs(4108) <= not (a and b);
    layer4_outputs(4109) <= '1';
    layer4_outputs(4110) <= b;
    layer4_outputs(4111) <= not b;
    layer4_outputs(4112) <= a;
    layer4_outputs(4113) <= not (a or b);
    layer4_outputs(4114) <= not b;
    layer4_outputs(4115) <= not a;
    layer4_outputs(4116) <= a and b;
    layer4_outputs(4117) <= not a;
    layer4_outputs(4118) <= not (a or b);
    layer4_outputs(4119) <= not b;
    layer4_outputs(4120) <= b;
    layer4_outputs(4121) <= not a;
    layer4_outputs(4122) <= not a;
    layer4_outputs(4123) <= a xor b;
    layer4_outputs(4124) <= a xor b;
    layer4_outputs(4125) <= not a;
    layer4_outputs(4126) <= b;
    layer4_outputs(4127) <= not (a and b);
    layer4_outputs(4128) <= not (a and b);
    layer4_outputs(4129) <= not (a or b);
    layer4_outputs(4130) <= not a or b;
    layer4_outputs(4131) <= not b or a;
    layer4_outputs(4132) <= a;
    layer4_outputs(4133) <= '1';
    layer4_outputs(4134) <= a or b;
    layer4_outputs(4135) <= a and b;
    layer4_outputs(4136) <= b;
    layer4_outputs(4137) <= a;
    layer4_outputs(4138) <= not (a or b);
    layer4_outputs(4139) <= not a or b;
    layer4_outputs(4140) <= not (a and b);
    layer4_outputs(4141) <= not (a xor b);
    layer4_outputs(4142) <= not (a and b);
    layer4_outputs(4143) <= a xor b;
    layer4_outputs(4144) <= '1';
    layer4_outputs(4145) <= a and b;
    layer4_outputs(4146) <= a xor b;
    layer4_outputs(4147) <= b and not a;
    layer4_outputs(4148) <= not b;
    layer4_outputs(4149) <= not a;
    layer4_outputs(4150) <= b and not a;
    layer4_outputs(4151) <= not (a and b);
    layer4_outputs(4152) <= not a or b;
    layer4_outputs(4153) <= not (a xor b);
    layer4_outputs(4154) <= not a or b;
    layer4_outputs(4155) <= a and not b;
    layer4_outputs(4156) <= a;
    layer4_outputs(4157) <= not a or b;
    layer4_outputs(4158) <= a;
    layer4_outputs(4159) <= a and not b;
    layer4_outputs(4160) <= a;
    layer4_outputs(4161) <= a and b;
    layer4_outputs(4162) <= a;
    layer4_outputs(4163) <= not b;
    layer4_outputs(4164) <= b and not a;
    layer4_outputs(4165) <= a or b;
    layer4_outputs(4166) <= b;
    layer4_outputs(4167) <= a;
    layer4_outputs(4168) <= a and b;
    layer4_outputs(4169) <= not a or b;
    layer4_outputs(4170) <= not (a xor b);
    layer4_outputs(4171) <= b;
    layer4_outputs(4172) <= not a;
    layer4_outputs(4173) <= b and not a;
    layer4_outputs(4174) <= not a or b;
    layer4_outputs(4175) <= not (a or b);
    layer4_outputs(4176) <= b;
    layer4_outputs(4177) <= a or b;
    layer4_outputs(4178) <= not (a and b);
    layer4_outputs(4179) <= b and not a;
    layer4_outputs(4180) <= not (a and b);
    layer4_outputs(4181) <= not b;
    layer4_outputs(4182) <= a or b;
    layer4_outputs(4183) <= not b;
    layer4_outputs(4184) <= b;
    layer4_outputs(4185) <= b;
    layer4_outputs(4186) <= a xor b;
    layer4_outputs(4187) <= not b;
    layer4_outputs(4188) <= not (a or b);
    layer4_outputs(4189) <= a xor b;
    layer4_outputs(4190) <= not (a xor b);
    layer4_outputs(4191) <= not a;
    layer4_outputs(4192) <= b;
    layer4_outputs(4193) <= b;
    layer4_outputs(4194) <= a and not b;
    layer4_outputs(4195) <= '1';
    layer4_outputs(4196) <= b and not a;
    layer4_outputs(4197) <= '0';
    layer4_outputs(4198) <= not b or a;
    layer4_outputs(4199) <= a or b;
    layer4_outputs(4200) <= not (a xor b);
    layer4_outputs(4201) <= b;
    layer4_outputs(4202) <= a;
    layer4_outputs(4203) <= a;
    layer4_outputs(4204) <= not (a and b);
    layer4_outputs(4205) <= not a;
    layer4_outputs(4206) <= b and not a;
    layer4_outputs(4207) <= not a or b;
    layer4_outputs(4208) <= a and b;
    layer4_outputs(4209) <= not b or a;
    layer4_outputs(4210) <= not (a and b);
    layer4_outputs(4211) <= b and not a;
    layer4_outputs(4212) <= b;
    layer4_outputs(4213) <= b;
    layer4_outputs(4214) <= a xor b;
    layer4_outputs(4215) <= b;
    layer4_outputs(4216) <= not a;
    layer4_outputs(4217) <= not a;
    layer4_outputs(4218) <= a;
    layer4_outputs(4219) <= not b;
    layer4_outputs(4220) <= not (a and b);
    layer4_outputs(4221) <= not b or a;
    layer4_outputs(4222) <= a or b;
    layer4_outputs(4223) <= not (a or b);
    layer4_outputs(4224) <= not (a or b);
    layer4_outputs(4225) <= a;
    layer4_outputs(4226) <= not b;
    layer4_outputs(4227) <= a and b;
    layer4_outputs(4228) <= a and not b;
    layer4_outputs(4229) <= '0';
    layer4_outputs(4230) <= b and not a;
    layer4_outputs(4231) <= b;
    layer4_outputs(4232) <= not a or b;
    layer4_outputs(4233) <= not a;
    layer4_outputs(4234) <= a and not b;
    layer4_outputs(4235) <= a and b;
    layer4_outputs(4236) <= not b;
    layer4_outputs(4237) <= not (a and b);
    layer4_outputs(4238) <= b and not a;
    layer4_outputs(4239) <= not (a or b);
    layer4_outputs(4240) <= not (a or b);
    layer4_outputs(4241) <= not (a and b);
    layer4_outputs(4242) <= not (a or b);
    layer4_outputs(4243) <= b;
    layer4_outputs(4244) <= '1';
    layer4_outputs(4245) <= not b or a;
    layer4_outputs(4246) <= not a or b;
    layer4_outputs(4247) <= not b;
    layer4_outputs(4248) <= a xor b;
    layer4_outputs(4249) <= not a or b;
    layer4_outputs(4250) <= a or b;
    layer4_outputs(4251) <= not b or a;
    layer4_outputs(4252) <= not (a xor b);
    layer4_outputs(4253) <= not a;
    layer4_outputs(4254) <= not a or b;
    layer4_outputs(4255) <= a and b;
    layer4_outputs(4256) <= b and not a;
    layer4_outputs(4257) <= not a;
    layer4_outputs(4258) <= b;
    layer4_outputs(4259) <= b;
    layer4_outputs(4260) <= not a;
    layer4_outputs(4261) <= b and not a;
    layer4_outputs(4262) <= a and not b;
    layer4_outputs(4263) <= not b;
    layer4_outputs(4264) <= not a;
    layer4_outputs(4265) <= not b or a;
    layer4_outputs(4266) <= not a;
    layer4_outputs(4267) <= not a;
    layer4_outputs(4268) <= '0';
    layer4_outputs(4269) <= not (a or b);
    layer4_outputs(4270) <= a and not b;
    layer4_outputs(4271) <= not a;
    layer4_outputs(4272) <= not (a and b);
    layer4_outputs(4273) <= not a;
    layer4_outputs(4274) <= not a;
    layer4_outputs(4275) <= b;
    layer4_outputs(4276) <= a;
    layer4_outputs(4277) <= not b;
    layer4_outputs(4278) <= not b or a;
    layer4_outputs(4279) <= not (a xor b);
    layer4_outputs(4280) <= not b;
    layer4_outputs(4281) <= a or b;
    layer4_outputs(4282) <= not b or a;
    layer4_outputs(4283) <= b;
    layer4_outputs(4284) <= not b or a;
    layer4_outputs(4285) <= b;
    layer4_outputs(4286) <= not b;
    layer4_outputs(4287) <= a or b;
    layer4_outputs(4288) <= b;
    layer4_outputs(4289) <= a and not b;
    layer4_outputs(4290) <= not b;
    layer4_outputs(4291) <= a or b;
    layer4_outputs(4292) <= b and not a;
    layer4_outputs(4293) <= not (a or b);
    layer4_outputs(4294) <= b and not a;
    layer4_outputs(4295) <= not a;
    layer4_outputs(4296) <= a;
    layer4_outputs(4297) <= b;
    layer4_outputs(4298) <= not b or a;
    layer4_outputs(4299) <= not b or a;
    layer4_outputs(4300) <= not b or a;
    layer4_outputs(4301) <= not (a and b);
    layer4_outputs(4302) <= not a;
    layer4_outputs(4303) <= not b;
    layer4_outputs(4304) <= not b;
    layer4_outputs(4305) <= not (a or b);
    layer4_outputs(4306) <= not b;
    layer4_outputs(4307) <= not (a xor b);
    layer4_outputs(4308) <= b;
    layer4_outputs(4309) <= not b;
    layer4_outputs(4310) <= not (a and b);
    layer4_outputs(4311) <= not (a or b);
    layer4_outputs(4312) <= b;
    layer4_outputs(4313) <= a and b;
    layer4_outputs(4314) <= b and not a;
    layer4_outputs(4315) <= '0';
    layer4_outputs(4316) <= b;
    layer4_outputs(4317) <= a;
    layer4_outputs(4318) <= not b;
    layer4_outputs(4319) <= a;
    layer4_outputs(4320) <= a;
    layer4_outputs(4321) <= b and not a;
    layer4_outputs(4322) <= a;
    layer4_outputs(4323) <= a or b;
    layer4_outputs(4324) <= a;
    layer4_outputs(4325) <= a or b;
    layer4_outputs(4326) <= not (a and b);
    layer4_outputs(4327) <= b and not a;
    layer4_outputs(4328) <= b;
    layer4_outputs(4329) <= b;
    layer4_outputs(4330) <= not a;
    layer4_outputs(4331) <= not (a xor b);
    layer4_outputs(4332) <= not b or a;
    layer4_outputs(4333) <= not a or b;
    layer4_outputs(4334) <= not b;
    layer4_outputs(4335) <= not (a and b);
    layer4_outputs(4336) <= not a;
    layer4_outputs(4337) <= not (a or b);
    layer4_outputs(4338) <= b;
    layer4_outputs(4339) <= '1';
    layer4_outputs(4340) <= not a;
    layer4_outputs(4341) <= b;
    layer4_outputs(4342) <= not b;
    layer4_outputs(4343) <= b;
    layer4_outputs(4344) <= not b;
    layer4_outputs(4345) <= a;
    layer4_outputs(4346) <= b;
    layer4_outputs(4347) <= not a;
    layer4_outputs(4348) <= a or b;
    layer4_outputs(4349) <= not (a xor b);
    layer4_outputs(4350) <= not (a or b);
    layer4_outputs(4351) <= b;
    layer4_outputs(4352) <= a and b;
    layer4_outputs(4353) <= not a;
    layer4_outputs(4354) <= not a;
    layer4_outputs(4355) <= a;
    layer4_outputs(4356) <= a and not b;
    layer4_outputs(4357) <= not b;
    layer4_outputs(4358) <= b and not a;
    layer4_outputs(4359) <= not a or b;
    layer4_outputs(4360) <= not b;
    layer4_outputs(4361) <= not b or a;
    layer4_outputs(4362) <= not a or b;
    layer4_outputs(4363) <= not a or b;
    layer4_outputs(4364) <= not (a or b);
    layer4_outputs(4365) <= b and not a;
    layer4_outputs(4366) <= not b;
    layer4_outputs(4367) <= a;
    layer4_outputs(4368) <= not a or b;
    layer4_outputs(4369) <= not a;
    layer4_outputs(4370) <= a;
    layer4_outputs(4371) <= a and not b;
    layer4_outputs(4372) <= a and b;
    layer4_outputs(4373) <= not (a xor b);
    layer4_outputs(4374) <= not a or b;
    layer4_outputs(4375) <= not (a xor b);
    layer4_outputs(4376) <= not (a and b);
    layer4_outputs(4377) <= a and not b;
    layer4_outputs(4378) <= b;
    layer4_outputs(4379) <= '1';
    layer4_outputs(4380) <= b;
    layer4_outputs(4381) <= a and not b;
    layer4_outputs(4382) <= a and not b;
    layer4_outputs(4383) <= not (a or b);
    layer4_outputs(4384) <= not a;
    layer4_outputs(4385) <= not a;
    layer4_outputs(4386) <= not (a xor b);
    layer4_outputs(4387) <= a xor b;
    layer4_outputs(4388) <= not a or b;
    layer4_outputs(4389) <= not b;
    layer4_outputs(4390) <= not b;
    layer4_outputs(4391) <= not (a xor b);
    layer4_outputs(4392) <= not (a or b);
    layer4_outputs(4393) <= not (a and b);
    layer4_outputs(4394) <= not b or a;
    layer4_outputs(4395) <= a;
    layer4_outputs(4396) <= b;
    layer4_outputs(4397) <= not b;
    layer4_outputs(4398) <= not a or b;
    layer4_outputs(4399) <= a xor b;
    layer4_outputs(4400) <= a and b;
    layer4_outputs(4401) <= not a;
    layer4_outputs(4402) <= not b;
    layer4_outputs(4403) <= not (a or b);
    layer4_outputs(4404) <= not (a and b);
    layer4_outputs(4405) <= not a;
    layer4_outputs(4406) <= a and not b;
    layer4_outputs(4407) <= a;
    layer4_outputs(4408) <= b and not a;
    layer4_outputs(4409) <= a xor b;
    layer4_outputs(4410) <= b;
    layer4_outputs(4411) <= b;
    layer4_outputs(4412) <= b and not a;
    layer4_outputs(4413) <= a and not b;
    layer4_outputs(4414) <= not a or b;
    layer4_outputs(4415) <= '0';
    layer4_outputs(4416) <= not (a xor b);
    layer4_outputs(4417) <= not b;
    layer4_outputs(4418) <= b;
    layer4_outputs(4419) <= not b;
    layer4_outputs(4420) <= not b or a;
    layer4_outputs(4421) <= not b or a;
    layer4_outputs(4422) <= not (a and b);
    layer4_outputs(4423) <= not (a xor b);
    layer4_outputs(4424) <= not b or a;
    layer4_outputs(4425) <= not (a and b);
    layer4_outputs(4426) <= b;
    layer4_outputs(4427) <= not (a xor b);
    layer4_outputs(4428) <= a or b;
    layer4_outputs(4429) <= not (a xor b);
    layer4_outputs(4430) <= a or b;
    layer4_outputs(4431) <= not a or b;
    layer4_outputs(4432) <= a;
    layer4_outputs(4433) <= a;
    layer4_outputs(4434) <= b;
    layer4_outputs(4435) <= not b or a;
    layer4_outputs(4436) <= a;
    layer4_outputs(4437) <= not a;
    layer4_outputs(4438) <= not a or b;
    layer4_outputs(4439) <= not a;
    layer4_outputs(4440) <= b;
    layer4_outputs(4441) <= a;
    layer4_outputs(4442) <= b;
    layer4_outputs(4443) <= a;
    layer4_outputs(4444) <= a;
    layer4_outputs(4445) <= b;
    layer4_outputs(4446) <= b;
    layer4_outputs(4447) <= a;
    layer4_outputs(4448) <= b;
    layer4_outputs(4449) <= a or b;
    layer4_outputs(4450) <= not b;
    layer4_outputs(4451) <= a;
    layer4_outputs(4452) <= a;
    layer4_outputs(4453) <= a and not b;
    layer4_outputs(4454) <= not a or b;
    layer4_outputs(4455) <= not a;
    layer4_outputs(4456) <= not a;
    layer4_outputs(4457) <= a;
    layer4_outputs(4458) <= not a;
    layer4_outputs(4459) <= b;
    layer4_outputs(4460) <= '0';
    layer4_outputs(4461) <= not a;
    layer4_outputs(4462) <= b;
    layer4_outputs(4463) <= a xor b;
    layer4_outputs(4464) <= b and not a;
    layer4_outputs(4465) <= not (a and b);
    layer4_outputs(4466) <= not b or a;
    layer4_outputs(4467) <= not a;
    layer4_outputs(4468) <= not b;
    layer4_outputs(4469) <= not (a and b);
    layer4_outputs(4470) <= not (a and b);
    layer4_outputs(4471) <= not b;
    layer4_outputs(4472) <= b;
    layer4_outputs(4473) <= not a or b;
    layer4_outputs(4474) <= a and b;
    layer4_outputs(4475) <= not (a and b);
    layer4_outputs(4476) <= a;
    layer4_outputs(4477) <= a and b;
    layer4_outputs(4478) <= not a;
    layer4_outputs(4479) <= a xor b;
    layer4_outputs(4480) <= not a or b;
    layer4_outputs(4481) <= not b or a;
    layer4_outputs(4482) <= not b;
    layer4_outputs(4483) <= not b or a;
    layer4_outputs(4484) <= not (a or b);
    layer4_outputs(4485) <= not a;
    layer4_outputs(4486) <= not (a xor b);
    layer4_outputs(4487) <= b;
    layer4_outputs(4488) <= not b;
    layer4_outputs(4489) <= not a or b;
    layer4_outputs(4490) <= b;
    layer4_outputs(4491) <= b;
    layer4_outputs(4492) <= b;
    layer4_outputs(4493) <= not (a and b);
    layer4_outputs(4494) <= not (a xor b);
    layer4_outputs(4495) <= a;
    layer4_outputs(4496) <= not b or a;
    layer4_outputs(4497) <= a and not b;
    layer4_outputs(4498) <= not a;
    layer4_outputs(4499) <= b;
    layer4_outputs(4500) <= a xor b;
    layer4_outputs(4501) <= b;
    layer4_outputs(4502) <= not a;
    layer4_outputs(4503) <= a and not b;
    layer4_outputs(4504) <= not b;
    layer4_outputs(4505) <= not b;
    layer4_outputs(4506) <= b;
    layer4_outputs(4507) <= not b;
    layer4_outputs(4508) <= a and b;
    layer4_outputs(4509) <= not a or b;
    layer4_outputs(4510) <= not b;
    layer4_outputs(4511) <= a;
    layer4_outputs(4512) <= not a;
    layer4_outputs(4513) <= a and b;
    layer4_outputs(4514) <= not b or a;
    layer4_outputs(4515) <= not b;
    layer4_outputs(4516) <= not b;
    layer4_outputs(4517) <= '0';
    layer4_outputs(4518) <= not a;
    layer4_outputs(4519) <= a;
    layer4_outputs(4520) <= a;
    layer4_outputs(4521) <= not b;
    layer4_outputs(4522) <= not b or a;
    layer4_outputs(4523) <= a and b;
    layer4_outputs(4524) <= not a or b;
    layer4_outputs(4525) <= not a;
    layer4_outputs(4526) <= not (a or b);
    layer4_outputs(4527) <= a and not b;
    layer4_outputs(4528) <= not a or b;
    layer4_outputs(4529) <= b and not a;
    layer4_outputs(4530) <= a or b;
    layer4_outputs(4531) <= a;
    layer4_outputs(4532) <= not b;
    layer4_outputs(4533) <= not b;
    layer4_outputs(4534) <= not a;
    layer4_outputs(4535) <= a;
    layer4_outputs(4536) <= a;
    layer4_outputs(4537) <= a;
    layer4_outputs(4538) <= '0';
    layer4_outputs(4539) <= not a;
    layer4_outputs(4540) <= a and b;
    layer4_outputs(4541) <= a xor b;
    layer4_outputs(4542) <= not b;
    layer4_outputs(4543) <= '0';
    layer4_outputs(4544) <= a and b;
    layer4_outputs(4545) <= b and not a;
    layer4_outputs(4546) <= a and not b;
    layer4_outputs(4547) <= not a;
    layer4_outputs(4548) <= not a;
    layer4_outputs(4549) <= b and not a;
    layer4_outputs(4550) <= not b or a;
    layer4_outputs(4551) <= not (a or b);
    layer4_outputs(4552) <= not b or a;
    layer4_outputs(4553) <= a and b;
    layer4_outputs(4554) <= not a;
    layer4_outputs(4555) <= a or b;
    layer4_outputs(4556) <= a;
    layer4_outputs(4557) <= a and not b;
    layer4_outputs(4558) <= b;
    layer4_outputs(4559) <= not a;
    layer4_outputs(4560) <= not a;
    layer4_outputs(4561) <= a xor b;
    layer4_outputs(4562) <= b;
    layer4_outputs(4563) <= not b or a;
    layer4_outputs(4564) <= not b;
    layer4_outputs(4565) <= not (a and b);
    layer4_outputs(4566) <= not a;
    layer4_outputs(4567) <= a and not b;
    layer4_outputs(4568) <= a;
    layer4_outputs(4569) <= a and b;
    layer4_outputs(4570) <= not a;
    layer4_outputs(4571) <= not b or a;
    layer4_outputs(4572) <= not a;
    layer4_outputs(4573) <= not (a or b);
    layer4_outputs(4574) <= a;
    layer4_outputs(4575) <= a and b;
    layer4_outputs(4576) <= not (a xor b);
    layer4_outputs(4577) <= '1';
    layer4_outputs(4578) <= a;
    layer4_outputs(4579) <= b and not a;
    layer4_outputs(4580) <= not a;
    layer4_outputs(4581) <= b;
    layer4_outputs(4582) <= b and not a;
    layer4_outputs(4583) <= not b;
    layer4_outputs(4584) <= a and b;
    layer4_outputs(4585) <= a;
    layer4_outputs(4586) <= b and not a;
    layer4_outputs(4587) <= b;
    layer4_outputs(4588) <= not b;
    layer4_outputs(4589) <= b and not a;
    layer4_outputs(4590) <= a and b;
    layer4_outputs(4591) <= a xor b;
    layer4_outputs(4592) <= a;
    layer4_outputs(4593) <= not a;
    layer4_outputs(4594) <= not (a xor b);
    layer4_outputs(4595) <= b;
    layer4_outputs(4596) <= b;
    layer4_outputs(4597) <= not (a or b);
    layer4_outputs(4598) <= a or b;
    layer4_outputs(4599) <= a and b;
    layer4_outputs(4600) <= not b;
    layer4_outputs(4601) <= not b;
    layer4_outputs(4602) <= a;
    layer4_outputs(4603) <= a and not b;
    layer4_outputs(4604) <= b;
    layer4_outputs(4605) <= not a;
    layer4_outputs(4606) <= not a or b;
    layer4_outputs(4607) <= not (a or b);
    layer4_outputs(4608) <= not b;
    layer4_outputs(4609) <= not a;
    layer4_outputs(4610) <= a and b;
    layer4_outputs(4611) <= b;
    layer4_outputs(4612) <= not (a or b);
    layer4_outputs(4613) <= a;
    layer4_outputs(4614) <= not (a and b);
    layer4_outputs(4615) <= not b;
    layer4_outputs(4616) <= a and not b;
    layer4_outputs(4617) <= a;
    layer4_outputs(4618) <= not a or b;
    layer4_outputs(4619) <= not (a or b);
    layer4_outputs(4620) <= not a;
    layer4_outputs(4621) <= not a;
    layer4_outputs(4622) <= a and not b;
    layer4_outputs(4623) <= not b;
    layer4_outputs(4624) <= a and not b;
    layer4_outputs(4625) <= not b;
    layer4_outputs(4626) <= b;
    layer4_outputs(4627) <= b;
    layer4_outputs(4628) <= a and not b;
    layer4_outputs(4629) <= a and b;
    layer4_outputs(4630) <= not b or a;
    layer4_outputs(4631) <= b and not a;
    layer4_outputs(4632) <= a and b;
    layer4_outputs(4633) <= not a or b;
    layer4_outputs(4634) <= a xor b;
    layer4_outputs(4635) <= a and not b;
    layer4_outputs(4636) <= a and not b;
    layer4_outputs(4637) <= not b;
    layer4_outputs(4638) <= not b or a;
    layer4_outputs(4639) <= b and not a;
    layer4_outputs(4640) <= not (a and b);
    layer4_outputs(4641) <= not (a and b);
    layer4_outputs(4642) <= not a;
    layer4_outputs(4643) <= b;
    layer4_outputs(4644) <= not a or b;
    layer4_outputs(4645) <= a and b;
    layer4_outputs(4646) <= a and not b;
    layer4_outputs(4647) <= a or b;
    layer4_outputs(4648) <= '1';
    layer4_outputs(4649) <= b and not a;
    layer4_outputs(4650) <= not b or a;
    layer4_outputs(4651) <= not a;
    layer4_outputs(4652) <= a and b;
    layer4_outputs(4653) <= a and b;
    layer4_outputs(4654) <= a;
    layer4_outputs(4655) <= not a;
    layer4_outputs(4656) <= not a or b;
    layer4_outputs(4657) <= b and not a;
    layer4_outputs(4658) <= a;
    layer4_outputs(4659) <= not a or b;
    layer4_outputs(4660) <= a xor b;
    layer4_outputs(4661) <= not (a and b);
    layer4_outputs(4662) <= a;
    layer4_outputs(4663) <= a and not b;
    layer4_outputs(4664) <= not (a and b);
    layer4_outputs(4665) <= a;
    layer4_outputs(4666) <= not b;
    layer4_outputs(4667) <= a and b;
    layer4_outputs(4668) <= not b;
    layer4_outputs(4669) <= not a;
    layer4_outputs(4670) <= not b;
    layer4_outputs(4671) <= a;
    layer4_outputs(4672) <= b;
    layer4_outputs(4673) <= a xor b;
    layer4_outputs(4674) <= a;
    layer4_outputs(4675) <= not (a or b);
    layer4_outputs(4676) <= b;
    layer4_outputs(4677) <= not b;
    layer4_outputs(4678) <= not b;
    layer4_outputs(4679) <= not b or a;
    layer4_outputs(4680) <= a and b;
    layer4_outputs(4681) <= not b;
    layer4_outputs(4682) <= '0';
    layer4_outputs(4683) <= not (a and b);
    layer4_outputs(4684) <= not b or a;
    layer4_outputs(4685) <= not a or b;
    layer4_outputs(4686) <= b;
    layer4_outputs(4687) <= not b or a;
    layer4_outputs(4688) <= not (a xor b);
    layer4_outputs(4689) <= not a;
    layer4_outputs(4690) <= a;
    layer4_outputs(4691) <= not b;
    layer4_outputs(4692) <= a or b;
    layer4_outputs(4693) <= not (a xor b);
    layer4_outputs(4694) <= not a or b;
    layer4_outputs(4695) <= b;
    layer4_outputs(4696) <= not b or a;
    layer4_outputs(4697) <= a;
    layer4_outputs(4698) <= a or b;
    layer4_outputs(4699) <= not a;
    layer4_outputs(4700) <= not (a and b);
    layer4_outputs(4701) <= not b;
    layer4_outputs(4702) <= not b;
    layer4_outputs(4703) <= not (a or b);
    layer4_outputs(4704) <= not (a xor b);
    layer4_outputs(4705) <= not b;
    layer4_outputs(4706) <= not (a and b);
    layer4_outputs(4707) <= a;
    layer4_outputs(4708) <= a and b;
    layer4_outputs(4709) <= a and b;
    layer4_outputs(4710) <= '0';
    layer4_outputs(4711) <= a;
    layer4_outputs(4712) <= a and not b;
    layer4_outputs(4713) <= a or b;
    layer4_outputs(4714) <= a;
    layer4_outputs(4715) <= not b;
    layer4_outputs(4716) <= not (a or b);
    layer4_outputs(4717) <= b and not a;
    layer4_outputs(4718) <= not (a and b);
    layer4_outputs(4719) <= not b;
    layer4_outputs(4720) <= a;
    layer4_outputs(4721) <= not (a and b);
    layer4_outputs(4722) <= a or b;
    layer4_outputs(4723) <= b;
    layer4_outputs(4724) <= a and b;
    layer4_outputs(4725) <= a and not b;
    layer4_outputs(4726) <= a and b;
    layer4_outputs(4727) <= b;
    layer4_outputs(4728) <= not (a and b);
    layer4_outputs(4729) <= a and b;
    layer4_outputs(4730) <= not b or a;
    layer4_outputs(4731) <= not (a and b);
    layer4_outputs(4732) <= a xor b;
    layer4_outputs(4733) <= not b or a;
    layer4_outputs(4734) <= not (a xor b);
    layer4_outputs(4735) <= b;
    layer4_outputs(4736) <= not a or b;
    layer4_outputs(4737) <= a xor b;
    layer4_outputs(4738) <= not (a or b);
    layer4_outputs(4739) <= a or b;
    layer4_outputs(4740) <= not a;
    layer4_outputs(4741) <= a;
    layer4_outputs(4742) <= '1';
    layer4_outputs(4743) <= not (a and b);
    layer4_outputs(4744) <= not a;
    layer4_outputs(4745) <= not a;
    layer4_outputs(4746) <= a;
    layer4_outputs(4747) <= a;
    layer4_outputs(4748) <= a or b;
    layer4_outputs(4749) <= not b or a;
    layer4_outputs(4750) <= not (a xor b);
    layer4_outputs(4751) <= not (a xor b);
    layer4_outputs(4752) <= a or b;
    layer4_outputs(4753) <= not b;
    layer4_outputs(4754) <= not (a or b);
    layer4_outputs(4755) <= not a;
    layer4_outputs(4756) <= not (a xor b);
    layer4_outputs(4757) <= not a or b;
    layer4_outputs(4758) <= not b;
    layer4_outputs(4759) <= a and b;
    layer4_outputs(4760) <= not a or b;
    layer4_outputs(4761) <= a xor b;
    layer4_outputs(4762) <= a or b;
    layer4_outputs(4763) <= b;
    layer4_outputs(4764) <= a and not b;
    layer4_outputs(4765) <= not a;
    layer4_outputs(4766) <= a;
    layer4_outputs(4767) <= not (a xor b);
    layer4_outputs(4768) <= b;
    layer4_outputs(4769) <= not a or b;
    layer4_outputs(4770) <= not (a or b);
    layer4_outputs(4771) <= not a or b;
    layer4_outputs(4772) <= '0';
    layer4_outputs(4773) <= not b or a;
    layer4_outputs(4774) <= a;
    layer4_outputs(4775) <= b;
    layer4_outputs(4776) <= b;
    layer4_outputs(4777) <= not b or a;
    layer4_outputs(4778) <= a and not b;
    layer4_outputs(4779) <= not a;
    layer4_outputs(4780) <= not a or b;
    layer4_outputs(4781) <= b;
    layer4_outputs(4782) <= not b;
    layer4_outputs(4783) <= b;
    layer4_outputs(4784) <= not a;
    layer4_outputs(4785) <= not (a or b);
    layer4_outputs(4786) <= a;
    layer4_outputs(4787) <= b;
    layer4_outputs(4788) <= b;
    layer4_outputs(4789) <= not b;
    layer4_outputs(4790) <= not b or a;
    layer4_outputs(4791) <= not b;
    layer4_outputs(4792) <= not b;
    layer4_outputs(4793) <= a;
    layer4_outputs(4794) <= not (a and b);
    layer4_outputs(4795) <= not b;
    layer4_outputs(4796) <= a and not b;
    layer4_outputs(4797) <= not (a and b);
    layer4_outputs(4798) <= not b;
    layer4_outputs(4799) <= b;
    layer4_outputs(4800) <= not a or b;
    layer4_outputs(4801) <= a and not b;
    layer4_outputs(4802) <= b and not a;
    layer4_outputs(4803) <= a and not b;
    layer4_outputs(4804) <= '1';
    layer4_outputs(4805) <= not a or b;
    layer4_outputs(4806) <= not (a and b);
    layer4_outputs(4807) <= a or b;
    layer4_outputs(4808) <= not a or b;
    layer4_outputs(4809) <= a or b;
    layer4_outputs(4810) <= not a;
    layer4_outputs(4811) <= '0';
    layer4_outputs(4812) <= not a;
    layer4_outputs(4813) <= a and not b;
    layer4_outputs(4814) <= not b;
    layer4_outputs(4815) <= not (a and b);
    layer4_outputs(4816) <= a and b;
    layer4_outputs(4817) <= b;
    layer4_outputs(4818) <= not (a and b);
    layer4_outputs(4819) <= a xor b;
    layer4_outputs(4820) <= a or b;
    layer4_outputs(4821) <= a;
    layer4_outputs(4822) <= a xor b;
    layer4_outputs(4823) <= a and b;
    layer4_outputs(4824) <= '1';
    layer4_outputs(4825) <= not (a xor b);
    layer4_outputs(4826) <= not b or a;
    layer4_outputs(4827) <= not a;
    layer4_outputs(4828) <= not a;
    layer4_outputs(4829) <= not a or b;
    layer4_outputs(4830) <= not a;
    layer4_outputs(4831) <= a;
    layer4_outputs(4832) <= not (a or b);
    layer4_outputs(4833) <= a or b;
    layer4_outputs(4834) <= not a;
    layer4_outputs(4835) <= b;
    layer4_outputs(4836) <= b;
    layer4_outputs(4837) <= b;
    layer4_outputs(4838) <= a and not b;
    layer4_outputs(4839) <= b;
    layer4_outputs(4840) <= not b;
    layer4_outputs(4841) <= a and not b;
    layer4_outputs(4842) <= not a;
    layer4_outputs(4843) <= not (a xor b);
    layer4_outputs(4844) <= not (a and b);
    layer4_outputs(4845) <= a;
    layer4_outputs(4846) <= b;
    layer4_outputs(4847) <= a xor b;
    layer4_outputs(4848) <= a and not b;
    layer4_outputs(4849) <= a;
    layer4_outputs(4850) <= a or b;
    layer4_outputs(4851) <= a;
    layer4_outputs(4852) <= not b or a;
    layer4_outputs(4853) <= a;
    layer4_outputs(4854) <= not b;
    layer4_outputs(4855) <= not a;
    layer4_outputs(4856) <= not (a or b);
    layer4_outputs(4857) <= not (a or b);
    layer4_outputs(4858) <= a or b;
    layer4_outputs(4859) <= b;
    layer4_outputs(4860) <= not b;
    layer4_outputs(4861) <= not (a xor b);
    layer4_outputs(4862) <= not (a and b);
    layer4_outputs(4863) <= not a;
    layer4_outputs(4864) <= a;
    layer4_outputs(4865) <= not a or b;
    layer4_outputs(4866) <= not (a and b);
    layer4_outputs(4867) <= not b;
    layer4_outputs(4868) <= a;
    layer4_outputs(4869) <= not b;
    layer4_outputs(4870) <= a and b;
    layer4_outputs(4871) <= not a;
    layer4_outputs(4872) <= a;
    layer4_outputs(4873) <= a xor b;
    layer4_outputs(4874) <= not a;
    layer4_outputs(4875) <= not b;
    layer4_outputs(4876) <= not (a xor b);
    layer4_outputs(4877) <= a;
    layer4_outputs(4878) <= not a or b;
    layer4_outputs(4879) <= b;
    layer4_outputs(4880) <= not a;
    layer4_outputs(4881) <= b;
    layer4_outputs(4882) <= not (a xor b);
    layer4_outputs(4883) <= a and b;
    layer4_outputs(4884) <= a and not b;
    layer4_outputs(4885) <= not (a and b);
    layer4_outputs(4886) <= not a or b;
    layer4_outputs(4887) <= a and b;
    layer4_outputs(4888) <= b;
    layer4_outputs(4889) <= a;
    layer4_outputs(4890) <= not (a or b);
    layer4_outputs(4891) <= not a;
    layer4_outputs(4892) <= b;
    layer4_outputs(4893) <= '0';
    layer4_outputs(4894) <= b and not a;
    layer4_outputs(4895) <= not a;
    layer4_outputs(4896) <= not b;
    layer4_outputs(4897) <= a;
    layer4_outputs(4898) <= a xor b;
    layer4_outputs(4899) <= not b;
    layer4_outputs(4900) <= a or b;
    layer4_outputs(4901) <= not a;
    layer4_outputs(4902) <= a xor b;
    layer4_outputs(4903) <= b;
    layer4_outputs(4904) <= '1';
    layer4_outputs(4905) <= b and not a;
    layer4_outputs(4906) <= not a;
    layer4_outputs(4907) <= b;
    layer4_outputs(4908) <= b;
    layer4_outputs(4909) <= b;
    layer4_outputs(4910) <= a;
    layer4_outputs(4911) <= a xor b;
    layer4_outputs(4912) <= not b;
    layer4_outputs(4913) <= not a or b;
    layer4_outputs(4914) <= b;
    layer4_outputs(4915) <= not a;
    layer4_outputs(4916) <= a and b;
    layer4_outputs(4917) <= a or b;
    layer4_outputs(4918) <= b;
    layer4_outputs(4919) <= a and not b;
    layer4_outputs(4920) <= not (a or b);
    layer4_outputs(4921) <= b and not a;
    layer4_outputs(4922) <= a and b;
    layer4_outputs(4923) <= not (a or b);
    layer4_outputs(4924) <= '0';
    layer4_outputs(4925) <= not (a and b);
    layer4_outputs(4926) <= not a;
    layer4_outputs(4927) <= not a or b;
    layer4_outputs(4928) <= not b;
    layer4_outputs(4929) <= a and not b;
    layer4_outputs(4930) <= '0';
    layer4_outputs(4931) <= '1';
    layer4_outputs(4932) <= a and b;
    layer4_outputs(4933) <= a or b;
    layer4_outputs(4934) <= b and not a;
    layer4_outputs(4935) <= a xor b;
    layer4_outputs(4936) <= a and not b;
    layer4_outputs(4937) <= a or b;
    layer4_outputs(4938) <= '1';
    layer4_outputs(4939) <= a;
    layer4_outputs(4940) <= not a or b;
    layer4_outputs(4941) <= not a;
    layer4_outputs(4942) <= a and not b;
    layer4_outputs(4943) <= not b;
    layer4_outputs(4944) <= a xor b;
    layer4_outputs(4945) <= a xor b;
    layer4_outputs(4946) <= not b;
    layer4_outputs(4947) <= not a;
    layer4_outputs(4948) <= a xor b;
    layer4_outputs(4949) <= not a or b;
    layer4_outputs(4950) <= a and not b;
    layer4_outputs(4951) <= b;
    layer4_outputs(4952) <= not b;
    layer4_outputs(4953) <= b;
    layer4_outputs(4954) <= a or b;
    layer4_outputs(4955) <= a xor b;
    layer4_outputs(4956) <= not (a xor b);
    layer4_outputs(4957) <= not b;
    layer4_outputs(4958) <= not b;
    layer4_outputs(4959) <= a;
    layer4_outputs(4960) <= not b;
    layer4_outputs(4961) <= a xor b;
    layer4_outputs(4962) <= a;
    layer4_outputs(4963) <= not b or a;
    layer4_outputs(4964) <= not b;
    layer4_outputs(4965) <= a xor b;
    layer4_outputs(4966) <= b;
    layer4_outputs(4967) <= a or b;
    layer4_outputs(4968) <= not a;
    layer4_outputs(4969) <= '0';
    layer4_outputs(4970) <= b;
    layer4_outputs(4971) <= b and not a;
    layer4_outputs(4972) <= not a;
    layer4_outputs(4973) <= a;
    layer4_outputs(4974) <= not a;
    layer4_outputs(4975) <= '1';
    layer4_outputs(4976) <= not (a and b);
    layer4_outputs(4977) <= a and not b;
    layer4_outputs(4978) <= a and not b;
    layer4_outputs(4979) <= not a or b;
    layer4_outputs(4980) <= not (a and b);
    layer4_outputs(4981) <= not b or a;
    layer4_outputs(4982) <= not a;
    layer4_outputs(4983) <= not (a or b);
    layer4_outputs(4984) <= a;
    layer4_outputs(4985) <= a and b;
    layer4_outputs(4986) <= '1';
    layer4_outputs(4987) <= a;
    layer4_outputs(4988) <= not b or a;
    layer4_outputs(4989) <= not a;
    layer4_outputs(4990) <= not (a and b);
    layer4_outputs(4991) <= not a or b;
    layer4_outputs(4992) <= a;
    layer4_outputs(4993) <= not b or a;
    layer4_outputs(4994) <= not (a xor b);
    layer4_outputs(4995) <= not b;
    layer4_outputs(4996) <= a or b;
    layer4_outputs(4997) <= not a;
    layer4_outputs(4998) <= not (a or b);
    layer4_outputs(4999) <= not b;
    layer4_outputs(5000) <= a;
    layer4_outputs(5001) <= b;
    layer4_outputs(5002) <= '1';
    layer4_outputs(5003) <= a xor b;
    layer4_outputs(5004) <= a;
    layer4_outputs(5005) <= not (a and b);
    layer4_outputs(5006) <= not (a or b);
    layer4_outputs(5007) <= not b;
    layer4_outputs(5008) <= a and b;
    layer4_outputs(5009) <= not (a and b);
    layer4_outputs(5010) <= b;
    layer4_outputs(5011) <= b and not a;
    layer4_outputs(5012) <= b;
    layer4_outputs(5013) <= not a or b;
    layer4_outputs(5014) <= not a;
    layer4_outputs(5015) <= not (a or b);
    layer4_outputs(5016) <= a xor b;
    layer4_outputs(5017) <= a;
    layer4_outputs(5018) <= a and b;
    layer4_outputs(5019) <= a or b;
    layer4_outputs(5020) <= '1';
    layer4_outputs(5021) <= '1';
    layer4_outputs(5022) <= not (a or b);
    layer4_outputs(5023) <= not (a and b);
    layer4_outputs(5024) <= not a;
    layer4_outputs(5025) <= a;
    layer4_outputs(5026) <= not b or a;
    layer4_outputs(5027) <= a or b;
    layer4_outputs(5028) <= b and not a;
    layer4_outputs(5029) <= a or b;
    layer4_outputs(5030) <= not (a or b);
    layer4_outputs(5031) <= not b or a;
    layer4_outputs(5032) <= b;
    layer4_outputs(5033) <= not a;
    layer4_outputs(5034) <= not a;
    layer4_outputs(5035) <= not a;
    layer4_outputs(5036) <= a and not b;
    layer4_outputs(5037) <= a and not b;
    layer4_outputs(5038) <= not b;
    layer4_outputs(5039) <= not b or a;
    layer4_outputs(5040) <= not b;
    layer4_outputs(5041) <= b and not a;
    layer4_outputs(5042) <= not b;
    layer4_outputs(5043) <= not (a xor b);
    layer4_outputs(5044) <= a or b;
    layer4_outputs(5045) <= a;
    layer4_outputs(5046) <= not a;
    layer4_outputs(5047) <= not (a or b);
    layer4_outputs(5048) <= not (a xor b);
    layer4_outputs(5049) <= b and not a;
    layer4_outputs(5050) <= b;
    layer4_outputs(5051) <= not b;
    layer4_outputs(5052) <= not b or a;
    layer4_outputs(5053) <= a and b;
    layer4_outputs(5054) <= not b or a;
    layer4_outputs(5055) <= a and not b;
    layer4_outputs(5056) <= b and not a;
    layer4_outputs(5057) <= not b;
    layer4_outputs(5058) <= not a;
    layer4_outputs(5059) <= not b;
    layer4_outputs(5060) <= a;
    layer4_outputs(5061) <= b;
    layer4_outputs(5062) <= a xor b;
    layer4_outputs(5063) <= a;
    layer4_outputs(5064) <= b;
    layer4_outputs(5065) <= not b;
    layer4_outputs(5066) <= not b;
    layer4_outputs(5067) <= a and b;
    layer4_outputs(5068) <= a or b;
    layer4_outputs(5069) <= not b;
    layer4_outputs(5070) <= b and not a;
    layer4_outputs(5071) <= b;
    layer4_outputs(5072) <= not a or b;
    layer4_outputs(5073) <= not (a xor b);
    layer4_outputs(5074) <= b and not a;
    layer4_outputs(5075) <= a or b;
    layer4_outputs(5076) <= b;
    layer4_outputs(5077) <= not (a or b);
    layer4_outputs(5078) <= a and not b;
    layer4_outputs(5079) <= a;
    layer4_outputs(5080) <= a xor b;
    layer4_outputs(5081) <= not b or a;
    layer4_outputs(5082) <= a xor b;
    layer4_outputs(5083) <= b;
    layer4_outputs(5084) <= not a;
    layer4_outputs(5085) <= a;
    layer4_outputs(5086) <= a and not b;
    layer4_outputs(5087) <= not b;
    layer4_outputs(5088) <= not (a or b);
    layer4_outputs(5089) <= a and not b;
    layer4_outputs(5090) <= a;
    layer4_outputs(5091) <= not a or b;
    layer4_outputs(5092) <= a and not b;
    layer4_outputs(5093) <= a;
    layer4_outputs(5094) <= not (a xor b);
    layer4_outputs(5095) <= not a or b;
    layer4_outputs(5096) <= not a or b;
    layer4_outputs(5097) <= not b;
    layer4_outputs(5098) <= a and b;
    layer4_outputs(5099) <= b;
    layer4_outputs(5100) <= a or b;
    layer4_outputs(5101) <= not a;
    layer4_outputs(5102) <= '1';
    layer4_outputs(5103) <= not (a xor b);
    layer4_outputs(5104) <= b;
    layer4_outputs(5105) <= a and not b;
    layer4_outputs(5106) <= not a;
    layer4_outputs(5107) <= a or b;
    layer4_outputs(5108) <= a;
    layer4_outputs(5109) <= not (a xor b);
    layer4_outputs(5110) <= b and not a;
    layer4_outputs(5111) <= not (a or b);
    layer4_outputs(5112) <= not b;
    layer4_outputs(5113) <= '0';
    layer4_outputs(5114) <= not a;
    layer4_outputs(5115) <= not b or a;
    layer4_outputs(5116) <= not a;
    layer4_outputs(5117) <= not (a and b);
    layer4_outputs(5118) <= b;
    layer4_outputs(5119) <= b and not a;
    layer4_outputs(5120) <= a xor b;
    layer4_outputs(5121) <= not b or a;
    layer4_outputs(5122) <= not (a and b);
    layer4_outputs(5123) <= a and b;
    layer4_outputs(5124) <= a;
    layer4_outputs(5125) <= not b;
    layer4_outputs(5126) <= not a;
    layer4_outputs(5127) <= a or b;
    layer4_outputs(5128) <= not (a xor b);
    layer4_outputs(5129) <= '1';
    layer4_outputs(5130) <= '1';
    layer4_outputs(5131) <= a and b;
    layer4_outputs(5132) <= a and not b;
    layer4_outputs(5133) <= a xor b;
    layer4_outputs(5134) <= b;
    layer4_outputs(5135) <= a or b;
    layer4_outputs(5136) <= not b or a;
    layer4_outputs(5137) <= not a;
    layer4_outputs(5138) <= not (a xor b);
    layer4_outputs(5139) <= b and not a;
    layer4_outputs(5140) <= a xor b;
    layer4_outputs(5141) <= not (a or b);
    layer4_outputs(5142) <= b;
    layer4_outputs(5143) <= a and not b;
    layer4_outputs(5144) <= not (a and b);
    layer4_outputs(5145) <= not (a and b);
    layer4_outputs(5146) <= not a;
    layer4_outputs(5147) <= a xor b;
    layer4_outputs(5148) <= '0';
    layer4_outputs(5149) <= b;
    layer4_outputs(5150) <= b and not a;
    layer4_outputs(5151) <= not (a or b);
    layer4_outputs(5152) <= not b or a;
    layer4_outputs(5153) <= '0';
    layer4_outputs(5154) <= a;
    layer4_outputs(5155) <= not b or a;
    layer4_outputs(5156) <= not (a or b);
    layer4_outputs(5157) <= b and not a;
    layer4_outputs(5158) <= not a or b;
    layer4_outputs(5159) <= not b or a;
    layer4_outputs(5160) <= b;
    layer4_outputs(5161) <= not b;
    layer4_outputs(5162) <= a;
    layer4_outputs(5163) <= a or b;
    layer4_outputs(5164) <= not a;
    layer4_outputs(5165) <= a or b;
    layer4_outputs(5166) <= a or b;
    layer4_outputs(5167) <= not (a and b);
    layer4_outputs(5168) <= not (a xor b);
    layer4_outputs(5169) <= not b;
    layer4_outputs(5170) <= not b or a;
    layer4_outputs(5171) <= '0';
    layer4_outputs(5172) <= not (a and b);
    layer4_outputs(5173) <= not b;
    layer4_outputs(5174) <= a;
    layer4_outputs(5175) <= '1';
    layer4_outputs(5176) <= not b;
    layer4_outputs(5177) <= a;
    layer4_outputs(5178) <= not (a xor b);
    layer4_outputs(5179) <= a;
    layer4_outputs(5180) <= a or b;
    layer4_outputs(5181) <= not a;
    layer4_outputs(5182) <= not a;
    layer4_outputs(5183) <= a xor b;
    layer4_outputs(5184) <= b;
    layer4_outputs(5185) <= not a;
    layer4_outputs(5186) <= a;
    layer4_outputs(5187) <= not a;
    layer4_outputs(5188) <= not (a or b);
    layer4_outputs(5189) <= b;
    layer4_outputs(5190) <= a;
    layer4_outputs(5191) <= not (a and b);
    layer4_outputs(5192) <= a and b;
    layer4_outputs(5193) <= a xor b;
    layer4_outputs(5194) <= a;
    layer4_outputs(5195) <= a and b;
    layer4_outputs(5196) <= not a or b;
    layer4_outputs(5197) <= b;
    layer4_outputs(5198) <= not a;
    layer4_outputs(5199) <= a and b;
    layer4_outputs(5200) <= not a;
    layer4_outputs(5201) <= not a;
    layer4_outputs(5202) <= a and b;
    layer4_outputs(5203) <= not (a xor b);
    layer4_outputs(5204) <= not b or a;
    layer4_outputs(5205) <= a and not b;
    layer4_outputs(5206) <= a xor b;
    layer4_outputs(5207) <= b;
    layer4_outputs(5208) <= a xor b;
    layer4_outputs(5209) <= a;
    layer4_outputs(5210) <= not a;
    layer4_outputs(5211) <= not (a and b);
    layer4_outputs(5212) <= not (a xor b);
    layer4_outputs(5213) <= not (a and b);
    layer4_outputs(5214) <= a xor b;
    layer4_outputs(5215) <= not (a and b);
    layer4_outputs(5216) <= b;
    layer4_outputs(5217) <= a;
    layer4_outputs(5218) <= not b or a;
    layer4_outputs(5219) <= b and not a;
    layer4_outputs(5220) <= b;
    layer4_outputs(5221) <= a and not b;
    layer4_outputs(5222) <= b;
    layer4_outputs(5223) <= b;
    layer4_outputs(5224) <= a xor b;
    layer4_outputs(5225) <= a or b;
    layer4_outputs(5226) <= not (a or b);
    layer4_outputs(5227) <= a or b;
    layer4_outputs(5228) <= a xor b;
    layer4_outputs(5229) <= a and not b;
    layer4_outputs(5230) <= b;
    layer4_outputs(5231) <= not a;
    layer4_outputs(5232) <= a and b;
    layer4_outputs(5233) <= a and not b;
    layer4_outputs(5234) <= not b;
    layer4_outputs(5235) <= not (a and b);
    layer4_outputs(5236) <= not (a xor b);
    layer4_outputs(5237) <= b and not a;
    layer4_outputs(5238) <= not (a or b);
    layer4_outputs(5239) <= not a;
    layer4_outputs(5240) <= '0';
    layer4_outputs(5241) <= not (a or b);
    layer4_outputs(5242) <= not b;
    layer4_outputs(5243) <= b;
    layer4_outputs(5244) <= not (a and b);
    layer4_outputs(5245) <= not (a and b);
    layer4_outputs(5246) <= not a;
    layer4_outputs(5247) <= not b;
    layer4_outputs(5248) <= not b;
    layer4_outputs(5249) <= '1';
    layer4_outputs(5250) <= not a;
    layer4_outputs(5251) <= a xor b;
    layer4_outputs(5252) <= b and not a;
    layer4_outputs(5253) <= '1';
    layer4_outputs(5254) <= a;
    layer4_outputs(5255) <= not a;
    layer4_outputs(5256) <= b;
    layer4_outputs(5257) <= not (a or b);
    layer4_outputs(5258) <= not (a and b);
    layer4_outputs(5259) <= not b or a;
    layer4_outputs(5260) <= b;
    layer4_outputs(5261) <= not b;
    layer4_outputs(5262) <= not (a xor b);
    layer4_outputs(5263) <= not a or b;
    layer4_outputs(5264) <= not (a xor b);
    layer4_outputs(5265) <= a or b;
    layer4_outputs(5266) <= b;
    layer4_outputs(5267) <= a and b;
    layer4_outputs(5268) <= a or b;
    layer4_outputs(5269) <= a;
    layer4_outputs(5270) <= not b;
    layer4_outputs(5271) <= b and not a;
    layer4_outputs(5272) <= not a;
    layer4_outputs(5273) <= not a or b;
    layer4_outputs(5274) <= not (a xor b);
    layer4_outputs(5275) <= b;
    layer4_outputs(5276) <= not b or a;
    layer4_outputs(5277) <= not b or a;
    layer4_outputs(5278) <= a xor b;
    layer4_outputs(5279) <= not (a xor b);
    layer4_outputs(5280) <= b and not a;
    layer4_outputs(5281) <= not (a xor b);
    layer4_outputs(5282) <= not (a xor b);
    layer4_outputs(5283) <= b;
    layer4_outputs(5284) <= b and not a;
    layer4_outputs(5285) <= not (a xor b);
    layer4_outputs(5286) <= not b or a;
    layer4_outputs(5287) <= not b or a;
    layer4_outputs(5288) <= not b;
    layer4_outputs(5289) <= a;
    layer4_outputs(5290) <= not b;
    layer4_outputs(5291) <= not (a and b);
    layer4_outputs(5292) <= not a or b;
    layer4_outputs(5293) <= not (a or b);
    layer4_outputs(5294) <= '1';
    layer4_outputs(5295) <= not a;
    layer4_outputs(5296) <= a and b;
    layer4_outputs(5297) <= not b;
    layer4_outputs(5298) <= not a;
    layer4_outputs(5299) <= not a;
    layer4_outputs(5300) <= not b;
    layer4_outputs(5301) <= not (a xor b);
    layer4_outputs(5302) <= a xor b;
    layer4_outputs(5303) <= b and not a;
    layer4_outputs(5304) <= not b;
    layer4_outputs(5305) <= not (a or b);
    layer4_outputs(5306) <= b and not a;
    layer4_outputs(5307) <= b;
    layer4_outputs(5308) <= not (a and b);
    layer4_outputs(5309) <= a xor b;
    layer4_outputs(5310) <= not a;
    layer4_outputs(5311) <= b;
    layer4_outputs(5312) <= not b;
    layer4_outputs(5313) <= not a;
    layer4_outputs(5314) <= not a;
    layer4_outputs(5315) <= not (a or b);
    layer4_outputs(5316) <= not a or b;
    layer4_outputs(5317) <= a and b;
    layer4_outputs(5318) <= b;
    layer4_outputs(5319) <= not (a or b);
    layer4_outputs(5320) <= a;
    layer4_outputs(5321) <= '1';
    layer4_outputs(5322) <= b;
    layer4_outputs(5323) <= b and not a;
    layer4_outputs(5324) <= a xor b;
    layer4_outputs(5325) <= a;
    layer4_outputs(5326) <= b;
    layer4_outputs(5327) <= a and not b;
    layer4_outputs(5328) <= a;
    layer4_outputs(5329) <= not a;
    layer4_outputs(5330) <= b;
    layer4_outputs(5331) <= not a;
    layer4_outputs(5332) <= not (a or b);
    layer4_outputs(5333) <= b;
    layer4_outputs(5334) <= not b;
    layer4_outputs(5335) <= not b or a;
    layer4_outputs(5336) <= not b;
    layer4_outputs(5337) <= not a;
    layer4_outputs(5338) <= not b or a;
    layer4_outputs(5339) <= a xor b;
    layer4_outputs(5340) <= not a;
    layer4_outputs(5341) <= not b or a;
    layer4_outputs(5342) <= b and not a;
    layer4_outputs(5343) <= not (a and b);
    layer4_outputs(5344) <= a and not b;
    layer4_outputs(5345) <= not (a xor b);
    layer4_outputs(5346) <= a;
    layer4_outputs(5347) <= a;
    layer4_outputs(5348) <= not (a and b);
    layer4_outputs(5349) <= a;
    layer4_outputs(5350) <= a and b;
    layer4_outputs(5351) <= b;
    layer4_outputs(5352) <= a xor b;
    layer4_outputs(5353) <= a;
    layer4_outputs(5354) <= not (a and b);
    layer4_outputs(5355) <= not a or b;
    layer4_outputs(5356) <= a;
    layer4_outputs(5357) <= a and b;
    layer4_outputs(5358) <= not a or b;
    layer4_outputs(5359) <= a;
    layer4_outputs(5360) <= not (a and b);
    layer4_outputs(5361) <= a;
    layer4_outputs(5362) <= b and not a;
    layer4_outputs(5363) <= not (a and b);
    layer4_outputs(5364) <= not b;
    layer4_outputs(5365) <= not b;
    layer4_outputs(5366) <= not b;
    layer4_outputs(5367) <= b and not a;
    layer4_outputs(5368) <= b;
    layer4_outputs(5369) <= not b or a;
    layer4_outputs(5370) <= a;
    layer4_outputs(5371) <= not b or a;
    layer4_outputs(5372) <= a or b;
    layer4_outputs(5373) <= not (a or b);
    layer4_outputs(5374) <= not b or a;
    layer4_outputs(5375) <= not b;
    layer4_outputs(5376) <= a and not b;
    layer4_outputs(5377) <= not (a and b);
    layer4_outputs(5378) <= a xor b;
    layer4_outputs(5379) <= not a;
    layer4_outputs(5380) <= not b;
    layer4_outputs(5381) <= not b or a;
    layer4_outputs(5382) <= a;
    layer4_outputs(5383) <= a;
    layer4_outputs(5384) <= a or b;
    layer4_outputs(5385) <= not a or b;
    layer4_outputs(5386) <= not b;
    layer4_outputs(5387) <= not (a or b);
    layer4_outputs(5388) <= a and b;
    layer4_outputs(5389) <= not a;
    layer4_outputs(5390) <= a and b;
    layer4_outputs(5391) <= not a or b;
    layer4_outputs(5392) <= b;
    layer4_outputs(5393) <= not b;
    layer4_outputs(5394) <= not a;
    layer4_outputs(5395) <= a or b;
    layer4_outputs(5396) <= not a;
    layer4_outputs(5397) <= not b or a;
    layer4_outputs(5398) <= a and b;
    layer4_outputs(5399) <= a and b;
    layer4_outputs(5400) <= not b;
    layer4_outputs(5401) <= not (a and b);
    layer4_outputs(5402) <= a;
    layer4_outputs(5403) <= not (a or b);
    layer4_outputs(5404) <= a or b;
    layer4_outputs(5405) <= not (a xor b);
    layer4_outputs(5406) <= b;
    layer4_outputs(5407) <= not (a and b);
    layer4_outputs(5408) <= '1';
    layer4_outputs(5409) <= not (a and b);
    layer4_outputs(5410) <= a;
    layer4_outputs(5411) <= not b or a;
    layer4_outputs(5412) <= a and not b;
    layer4_outputs(5413) <= a and not b;
    layer4_outputs(5414) <= not b;
    layer4_outputs(5415) <= not b;
    layer4_outputs(5416) <= not a;
    layer4_outputs(5417) <= a xor b;
    layer4_outputs(5418) <= b;
    layer4_outputs(5419) <= a and b;
    layer4_outputs(5420) <= a;
    layer4_outputs(5421) <= b;
    layer4_outputs(5422) <= b;
    layer4_outputs(5423) <= not a or b;
    layer4_outputs(5424) <= b and not a;
    layer4_outputs(5425) <= not b or a;
    layer4_outputs(5426) <= a;
    layer4_outputs(5427) <= a;
    layer4_outputs(5428) <= not a or b;
    layer4_outputs(5429) <= a;
    layer4_outputs(5430) <= a and not b;
    layer4_outputs(5431) <= a or b;
    layer4_outputs(5432) <= '1';
    layer4_outputs(5433) <= not b;
    layer4_outputs(5434) <= a or b;
    layer4_outputs(5435) <= a and not b;
    layer4_outputs(5436) <= a;
    layer4_outputs(5437) <= a and b;
    layer4_outputs(5438) <= not a;
    layer4_outputs(5439) <= b and not a;
    layer4_outputs(5440) <= a and b;
    layer4_outputs(5441) <= a xor b;
    layer4_outputs(5442) <= not b or a;
    layer4_outputs(5443) <= a or b;
    layer4_outputs(5444) <= b and not a;
    layer4_outputs(5445) <= b;
    layer4_outputs(5446) <= not a;
    layer4_outputs(5447) <= a;
    layer4_outputs(5448) <= '0';
    layer4_outputs(5449) <= not a;
    layer4_outputs(5450) <= not (a xor b);
    layer4_outputs(5451) <= not b;
    layer4_outputs(5452) <= a;
    layer4_outputs(5453) <= not b;
    layer4_outputs(5454) <= b;
    layer4_outputs(5455) <= a;
    layer4_outputs(5456) <= a and b;
    layer4_outputs(5457) <= not b;
    layer4_outputs(5458) <= not b;
    layer4_outputs(5459) <= not a or b;
    layer4_outputs(5460) <= '0';
    layer4_outputs(5461) <= not b;
    layer4_outputs(5462) <= b;
    layer4_outputs(5463) <= a and b;
    layer4_outputs(5464) <= a;
    layer4_outputs(5465) <= not a;
    layer4_outputs(5466) <= not b;
    layer4_outputs(5467) <= not b;
    layer4_outputs(5468) <= not (a and b);
    layer4_outputs(5469) <= not (a xor b);
    layer4_outputs(5470) <= not (a or b);
    layer4_outputs(5471) <= b;
    layer4_outputs(5472) <= b and not a;
    layer4_outputs(5473) <= not a or b;
    layer4_outputs(5474) <= a xor b;
    layer4_outputs(5475) <= a;
    layer4_outputs(5476) <= a and not b;
    layer4_outputs(5477) <= a xor b;
    layer4_outputs(5478) <= not b;
    layer4_outputs(5479) <= not a;
    layer4_outputs(5480) <= a or b;
    layer4_outputs(5481) <= a;
    layer4_outputs(5482) <= a;
    layer4_outputs(5483) <= not a;
    layer4_outputs(5484) <= not (a and b);
    layer4_outputs(5485) <= not a;
    layer4_outputs(5486) <= a and not b;
    layer4_outputs(5487) <= not a or b;
    layer4_outputs(5488) <= not (a or b);
    layer4_outputs(5489) <= b and not a;
    layer4_outputs(5490) <= a;
    layer4_outputs(5491) <= not b or a;
    layer4_outputs(5492) <= a or b;
    layer4_outputs(5493) <= a;
    layer4_outputs(5494) <= b and not a;
    layer4_outputs(5495) <= b and not a;
    layer4_outputs(5496) <= a;
    layer4_outputs(5497) <= b and not a;
    layer4_outputs(5498) <= not (a and b);
    layer4_outputs(5499) <= a xor b;
    layer4_outputs(5500) <= not a;
    layer4_outputs(5501) <= b and not a;
    layer4_outputs(5502) <= a or b;
    layer4_outputs(5503) <= b;
    layer4_outputs(5504) <= not (a or b);
    layer4_outputs(5505) <= not a or b;
    layer4_outputs(5506) <= a;
    layer4_outputs(5507) <= a and not b;
    layer4_outputs(5508) <= '1';
    layer4_outputs(5509) <= a and b;
    layer4_outputs(5510) <= a and not b;
    layer4_outputs(5511) <= not a;
    layer4_outputs(5512) <= a xor b;
    layer4_outputs(5513) <= '0';
    layer4_outputs(5514) <= b and not a;
    layer4_outputs(5515) <= not b or a;
    layer4_outputs(5516) <= '1';
    layer4_outputs(5517) <= not a or b;
    layer4_outputs(5518) <= not b;
    layer4_outputs(5519) <= a and not b;
    layer4_outputs(5520) <= b;
    layer4_outputs(5521) <= not (a and b);
    layer4_outputs(5522) <= b and not a;
    layer4_outputs(5523) <= not a;
    layer4_outputs(5524) <= a and not b;
    layer4_outputs(5525) <= b;
    layer4_outputs(5526) <= not a;
    layer4_outputs(5527) <= not (a or b);
    layer4_outputs(5528) <= not b or a;
    layer4_outputs(5529) <= not b;
    layer4_outputs(5530) <= a;
    layer4_outputs(5531) <= not b;
    layer4_outputs(5532) <= not (a or b);
    layer4_outputs(5533) <= not (a or b);
    layer4_outputs(5534) <= a;
    layer4_outputs(5535) <= not b;
    layer4_outputs(5536) <= a or b;
    layer4_outputs(5537) <= not (a or b);
    layer4_outputs(5538) <= not (a xor b);
    layer4_outputs(5539) <= not a;
    layer4_outputs(5540) <= not a;
    layer4_outputs(5541) <= a and b;
    layer4_outputs(5542) <= not b;
    layer4_outputs(5543) <= '0';
    layer4_outputs(5544) <= not b;
    layer4_outputs(5545) <= b;
    layer4_outputs(5546) <= not a or b;
    layer4_outputs(5547) <= a and not b;
    layer4_outputs(5548) <= a and not b;
    layer4_outputs(5549) <= a and b;
    layer4_outputs(5550) <= a;
    layer4_outputs(5551) <= not a;
    layer4_outputs(5552) <= a and b;
    layer4_outputs(5553) <= a;
    layer4_outputs(5554) <= a;
    layer4_outputs(5555) <= a or b;
    layer4_outputs(5556) <= not (a and b);
    layer4_outputs(5557) <= not b;
    layer4_outputs(5558) <= a;
    layer4_outputs(5559) <= not (a or b);
    layer4_outputs(5560) <= not (a and b);
    layer4_outputs(5561) <= b;
    layer4_outputs(5562) <= a and b;
    layer4_outputs(5563) <= a;
    layer4_outputs(5564) <= not a;
    layer4_outputs(5565) <= a;
    layer4_outputs(5566) <= a;
    layer4_outputs(5567) <= not a;
    layer4_outputs(5568) <= b;
    layer4_outputs(5569) <= b and not a;
    layer4_outputs(5570) <= b;
    layer4_outputs(5571) <= not (a and b);
    layer4_outputs(5572) <= not b;
    layer4_outputs(5573) <= not b;
    layer4_outputs(5574) <= '1';
    layer4_outputs(5575) <= a xor b;
    layer4_outputs(5576) <= not b;
    layer4_outputs(5577) <= a;
    layer4_outputs(5578) <= b and not a;
    layer4_outputs(5579) <= '1';
    layer4_outputs(5580) <= a;
    layer4_outputs(5581) <= b and not a;
    layer4_outputs(5582) <= a;
    layer4_outputs(5583) <= b and not a;
    layer4_outputs(5584) <= b;
    layer4_outputs(5585) <= not b;
    layer4_outputs(5586) <= not a or b;
    layer4_outputs(5587) <= a;
    layer4_outputs(5588) <= not b or a;
    layer4_outputs(5589) <= b;
    layer4_outputs(5590) <= a;
    layer4_outputs(5591) <= not b;
    layer4_outputs(5592) <= b and not a;
    layer4_outputs(5593) <= a;
    layer4_outputs(5594) <= a and not b;
    layer4_outputs(5595) <= not (a or b);
    layer4_outputs(5596) <= not b or a;
    layer4_outputs(5597) <= not a;
    layer4_outputs(5598) <= not a or b;
    layer4_outputs(5599) <= not (a xor b);
    layer4_outputs(5600) <= not (a and b);
    layer4_outputs(5601) <= a;
    layer4_outputs(5602) <= a and not b;
    layer4_outputs(5603) <= b and not a;
    layer4_outputs(5604) <= '1';
    layer4_outputs(5605) <= b;
    layer4_outputs(5606) <= a or b;
    layer4_outputs(5607) <= '1';
    layer4_outputs(5608) <= a and b;
    layer4_outputs(5609) <= not (a and b);
    layer4_outputs(5610) <= a and b;
    layer4_outputs(5611) <= b and not a;
    layer4_outputs(5612) <= a and b;
    layer4_outputs(5613) <= b;
    layer4_outputs(5614) <= not a;
    layer4_outputs(5615) <= not (a and b);
    layer4_outputs(5616) <= b;
    layer4_outputs(5617) <= not a;
    layer4_outputs(5618) <= b;
    layer4_outputs(5619) <= a;
    layer4_outputs(5620) <= b;
    layer4_outputs(5621) <= not b;
    layer4_outputs(5622) <= a and b;
    layer4_outputs(5623) <= '1';
    layer4_outputs(5624) <= b;
    layer4_outputs(5625) <= a and b;
    layer4_outputs(5626) <= a xor b;
    layer4_outputs(5627) <= a and not b;
    layer4_outputs(5628) <= a;
    layer4_outputs(5629) <= a;
    layer4_outputs(5630) <= not (a or b);
    layer4_outputs(5631) <= not b;
    layer4_outputs(5632) <= b;
    layer4_outputs(5633) <= a xor b;
    layer4_outputs(5634) <= not b;
    layer4_outputs(5635) <= a;
    layer4_outputs(5636) <= b;
    layer4_outputs(5637) <= not b or a;
    layer4_outputs(5638) <= not (a xor b);
    layer4_outputs(5639) <= a or b;
    layer4_outputs(5640) <= a;
    layer4_outputs(5641) <= not a or b;
    layer4_outputs(5642) <= b and not a;
    layer4_outputs(5643) <= not a;
    layer4_outputs(5644) <= a;
    layer4_outputs(5645) <= a and b;
    layer4_outputs(5646) <= a;
    layer4_outputs(5647) <= not a;
    layer4_outputs(5648) <= a;
    layer4_outputs(5649) <= not (a and b);
    layer4_outputs(5650) <= '0';
    layer4_outputs(5651) <= not a;
    layer4_outputs(5652) <= a or b;
    layer4_outputs(5653) <= not a;
    layer4_outputs(5654) <= not a;
    layer4_outputs(5655) <= not a or b;
    layer4_outputs(5656) <= '0';
    layer4_outputs(5657) <= '0';
    layer4_outputs(5658) <= a xor b;
    layer4_outputs(5659) <= b;
    layer4_outputs(5660) <= not b;
    layer4_outputs(5661) <= not b or a;
    layer4_outputs(5662) <= a;
    layer4_outputs(5663) <= not a;
    layer4_outputs(5664) <= b;
    layer4_outputs(5665) <= not (a or b);
    layer4_outputs(5666) <= not (a or b);
    layer4_outputs(5667) <= not a;
    layer4_outputs(5668) <= not (a and b);
    layer4_outputs(5669) <= a;
    layer4_outputs(5670) <= a and b;
    layer4_outputs(5671) <= a and not b;
    layer4_outputs(5672) <= not (a xor b);
    layer4_outputs(5673) <= b and not a;
    layer4_outputs(5674) <= not a or b;
    layer4_outputs(5675) <= not b;
    layer4_outputs(5676) <= a;
    layer4_outputs(5677) <= '1';
    layer4_outputs(5678) <= a and not b;
    layer4_outputs(5679) <= a and not b;
    layer4_outputs(5680) <= not (a xor b);
    layer4_outputs(5681) <= b and not a;
    layer4_outputs(5682) <= not (a or b);
    layer4_outputs(5683) <= a and not b;
    layer4_outputs(5684) <= b;
    layer4_outputs(5685) <= '0';
    layer4_outputs(5686) <= not b;
    layer4_outputs(5687) <= not (a or b);
    layer4_outputs(5688) <= a xor b;
    layer4_outputs(5689) <= not a;
    layer4_outputs(5690) <= not a;
    layer4_outputs(5691) <= b and not a;
    layer4_outputs(5692) <= a;
    layer4_outputs(5693) <= not a;
    layer4_outputs(5694) <= not a;
    layer4_outputs(5695) <= not (a and b);
    layer4_outputs(5696) <= '0';
    layer4_outputs(5697) <= not b or a;
    layer4_outputs(5698) <= a;
    layer4_outputs(5699) <= not b;
    layer4_outputs(5700) <= a and not b;
    layer4_outputs(5701) <= a xor b;
    layer4_outputs(5702) <= not a or b;
    layer4_outputs(5703) <= a or b;
    layer4_outputs(5704) <= not b;
    layer4_outputs(5705) <= not b;
    layer4_outputs(5706) <= a and not b;
    layer4_outputs(5707) <= a;
    layer4_outputs(5708) <= a;
    layer4_outputs(5709) <= a xor b;
    layer4_outputs(5710) <= not a;
    layer4_outputs(5711) <= not b;
    layer4_outputs(5712) <= not a;
    layer4_outputs(5713) <= not a;
    layer4_outputs(5714) <= a;
    layer4_outputs(5715) <= not (a or b);
    layer4_outputs(5716) <= not a;
    layer4_outputs(5717) <= a;
    layer4_outputs(5718) <= not b;
    layer4_outputs(5719) <= not b;
    layer4_outputs(5720) <= not b;
    layer4_outputs(5721) <= a;
    layer4_outputs(5722) <= a and not b;
    layer4_outputs(5723) <= not a or b;
    layer4_outputs(5724) <= not b;
    layer4_outputs(5725) <= not b;
    layer4_outputs(5726) <= not (a or b);
    layer4_outputs(5727) <= b;
    layer4_outputs(5728) <= not (a or b);
    layer4_outputs(5729) <= not b;
    layer4_outputs(5730) <= a and not b;
    layer4_outputs(5731) <= not a;
    layer4_outputs(5732) <= a;
    layer4_outputs(5733) <= not b;
    layer4_outputs(5734) <= not (a xor b);
    layer4_outputs(5735) <= b;
    layer4_outputs(5736) <= b and not a;
    layer4_outputs(5737) <= a;
    layer4_outputs(5738) <= a xor b;
    layer4_outputs(5739) <= not (a and b);
    layer4_outputs(5740) <= a;
    layer4_outputs(5741) <= not a;
    layer4_outputs(5742) <= not b;
    layer4_outputs(5743) <= a;
    layer4_outputs(5744) <= not b or a;
    layer4_outputs(5745) <= not a or b;
    layer4_outputs(5746) <= not a or b;
    layer4_outputs(5747) <= not (a xor b);
    layer4_outputs(5748) <= not b;
    layer4_outputs(5749) <= not a;
    layer4_outputs(5750) <= not (a or b);
    layer4_outputs(5751) <= not (a or b);
    layer4_outputs(5752) <= not (a and b);
    layer4_outputs(5753) <= not b;
    layer4_outputs(5754) <= a xor b;
    layer4_outputs(5755) <= not a;
    layer4_outputs(5756) <= not a or b;
    layer4_outputs(5757) <= not a;
    layer4_outputs(5758) <= a or b;
    layer4_outputs(5759) <= a xor b;
    layer4_outputs(5760) <= b;
    layer4_outputs(5761) <= not (a and b);
    layer4_outputs(5762) <= not (a xor b);
    layer4_outputs(5763) <= not (a xor b);
    layer4_outputs(5764) <= b and not a;
    layer4_outputs(5765) <= not b or a;
    layer4_outputs(5766) <= a xor b;
    layer4_outputs(5767) <= not a;
    layer4_outputs(5768) <= '1';
    layer4_outputs(5769) <= not a or b;
    layer4_outputs(5770) <= a and b;
    layer4_outputs(5771) <= not a;
    layer4_outputs(5772) <= not b;
    layer4_outputs(5773) <= not (a and b);
    layer4_outputs(5774) <= not b or a;
    layer4_outputs(5775) <= a and not b;
    layer4_outputs(5776) <= a and not b;
    layer4_outputs(5777) <= a;
    layer4_outputs(5778) <= b and not a;
    layer4_outputs(5779) <= a and not b;
    layer4_outputs(5780) <= not b;
    layer4_outputs(5781) <= not b or a;
    layer4_outputs(5782) <= a and not b;
    layer4_outputs(5783) <= not b;
    layer4_outputs(5784) <= not b or a;
    layer4_outputs(5785) <= not (a or b);
    layer4_outputs(5786) <= a and b;
    layer4_outputs(5787) <= not b or a;
    layer4_outputs(5788) <= '0';
    layer4_outputs(5789) <= not b;
    layer4_outputs(5790) <= not (a xor b);
    layer4_outputs(5791) <= a and b;
    layer4_outputs(5792) <= not a or b;
    layer4_outputs(5793) <= a and not b;
    layer4_outputs(5794) <= not a;
    layer4_outputs(5795) <= not a or b;
    layer4_outputs(5796) <= a and b;
    layer4_outputs(5797) <= a and not b;
    layer4_outputs(5798) <= '1';
    layer4_outputs(5799) <= not a;
    layer4_outputs(5800) <= a and b;
    layer4_outputs(5801) <= a or b;
    layer4_outputs(5802) <= a and not b;
    layer4_outputs(5803) <= not b or a;
    layer4_outputs(5804) <= not b or a;
    layer4_outputs(5805) <= not a;
    layer4_outputs(5806) <= not a;
    layer4_outputs(5807) <= a and b;
    layer4_outputs(5808) <= '0';
    layer4_outputs(5809) <= a;
    layer4_outputs(5810) <= not b or a;
    layer4_outputs(5811) <= a or b;
    layer4_outputs(5812) <= not b;
    layer4_outputs(5813) <= b;
    layer4_outputs(5814) <= a and b;
    layer4_outputs(5815) <= a xor b;
    layer4_outputs(5816) <= b;
    layer4_outputs(5817) <= a;
    layer4_outputs(5818) <= b;
    layer4_outputs(5819) <= not b;
    layer4_outputs(5820) <= a;
    layer4_outputs(5821) <= not a or b;
    layer4_outputs(5822) <= not b or a;
    layer4_outputs(5823) <= a and not b;
    layer4_outputs(5824) <= not a or b;
    layer4_outputs(5825) <= a or b;
    layer4_outputs(5826) <= a and b;
    layer4_outputs(5827) <= b;
    layer4_outputs(5828) <= a;
    layer4_outputs(5829) <= b;
    layer4_outputs(5830) <= not (a and b);
    layer4_outputs(5831) <= not b or a;
    layer4_outputs(5832) <= not a;
    layer4_outputs(5833) <= not (a xor b);
    layer4_outputs(5834) <= a and b;
    layer4_outputs(5835) <= b and not a;
    layer4_outputs(5836) <= not b;
    layer4_outputs(5837) <= b;
    layer4_outputs(5838) <= not a;
    layer4_outputs(5839) <= not b;
    layer4_outputs(5840) <= a;
    layer4_outputs(5841) <= not b;
    layer4_outputs(5842) <= not (a xor b);
    layer4_outputs(5843) <= not (a xor b);
    layer4_outputs(5844) <= not b;
    layer4_outputs(5845) <= not (a and b);
    layer4_outputs(5846) <= a and b;
    layer4_outputs(5847) <= b;
    layer4_outputs(5848) <= not (a and b);
    layer4_outputs(5849) <= not (a or b);
    layer4_outputs(5850) <= a or b;
    layer4_outputs(5851) <= not a or b;
    layer4_outputs(5852) <= a xor b;
    layer4_outputs(5853) <= not b;
    layer4_outputs(5854) <= a and not b;
    layer4_outputs(5855) <= b;
    layer4_outputs(5856) <= a;
    layer4_outputs(5857) <= b and not a;
    layer4_outputs(5858) <= not (a xor b);
    layer4_outputs(5859) <= not a;
    layer4_outputs(5860) <= a and not b;
    layer4_outputs(5861) <= '1';
    layer4_outputs(5862) <= not (a xor b);
    layer4_outputs(5863) <= b and not a;
    layer4_outputs(5864) <= b and not a;
    layer4_outputs(5865) <= a or b;
    layer4_outputs(5866) <= a xor b;
    layer4_outputs(5867) <= b;
    layer4_outputs(5868) <= b;
    layer4_outputs(5869) <= not (a or b);
    layer4_outputs(5870) <= not (a or b);
    layer4_outputs(5871) <= not (a xor b);
    layer4_outputs(5872) <= not a or b;
    layer4_outputs(5873) <= not (a xor b);
    layer4_outputs(5874) <= not b;
    layer4_outputs(5875) <= a;
    layer4_outputs(5876) <= b;
    layer4_outputs(5877) <= not (a or b);
    layer4_outputs(5878) <= b and not a;
    layer4_outputs(5879) <= a;
    layer4_outputs(5880) <= b;
    layer4_outputs(5881) <= a or b;
    layer4_outputs(5882) <= b and not a;
    layer4_outputs(5883) <= a;
    layer4_outputs(5884) <= not b;
    layer4_outputs(5885) <= a;
    layer4_outputs(5886) <= a or b;
    layer4_outputs(5887) <= not a;
    layer4_outputs(5888) <= not a;
    layer4_outputs(5889) <= b;
    layer4_outputs(5890) <= b;
    layer4_outputs(5891) <= not (a xor b);
    layer4_outputs(5892) <= b and not a;
    layer4_outputs(5893) <= not a or b;
    layer4_outputs(5894) <= a and b;
    layer4_outputs(5895) <= a and not b;
    layer4_outputs(5896) <= '1';
    layer4_outputs(5897) <= a or b;
    layer4_outputs(5898) <= not b;
    layer4_outputs(5899) <= a xor b;
    layer4_outputs(5900) <= a and not b;
    layer4_outputs(5901) <= b and not a;
    layer4_outputs(5902) <= a xor b;
    layer4_outputs(5903) <= not b or a;
    layer4_outputs(5904) <= not b;
    layer4_outputs(5905) <= a;
    layer4_outputs(5906) <= b and not a;
    layer4_outputs(5907) <= b;
    layer4_outputs(5908) <= a and b;
    layer4_outputs(5909) <= a;
    layer4_outputs(5910) <= a or b;
    layer4_outputs(5911) <= b;
    layer4_outputs(5912) <= not (a or b);
    layer4_outputs(5913) <= not a or b;
    layer4_outputs(5914) <= a and not b;
    layer4_outputs(5915) <= a;
    layer4_outputs(5916) <= not (a and b);
    layer4_outputs(5917) <= '0';
    layer4_outputs(5918) <= b;
    layer4_outputs(5919) <= not b;
    layer4_outputs(5920) <= not b;
    layer4_outputs(5921) <= a;
    layer4_outputs(5922) <= not (a xor b);
    layer4_outputs(5923) <= b;
    layer4_outputs(5924) <= not a or b;
    layer4_outputs(5925) <= not a;
    layer4_outputs(5926) <= not a;
    layer4_outputs(5927) <= a xor b;
    layer4_outputs(5928) <= a;
    layer4_outputs(5929) <= not a or b;
    layer4_outputs(5930) <= a or b;
    layer4_outputs(5931) <= b;
    layer4_outputs(5932) <= not a;
    layer4_outputs(5933) <= a;
    layer4_outputs(5934) <= a and b;
    layer4_outputs(5935) <= a or b;
    layer4_outputs(5936) <= b;
    layer4_outputs(5937) <= a;
    layer4_outputs(5938) <= not (a xor b);
    layer4_outputs(5939) <= not (a and b);
    layer4_outputs(5940) <= a and not b;
    layer4_outputs(5941) <= not b;
    layer4_outputs(5942) <= a or b;
    layer4_outputs(5943) <= b;
    layer4_outputs(5944) <= b and not a;
    layer4_outputs(5945) <= '1';
    layer4_outputs(5946) <= not (a xor b);
    layer4_outputs(5947) <= not a or b;
    layer4_outputs(5948) <= not a;
    layer4_outputs(5949) <= not b;
    layer4_outputs(5950) <= not b;
    layer4_outputs(5951) <= b and not a;
    layer4_outputs(5952) <= '0';
    layer4_outputs(5953) <= not b;
    layer4_outputs(5954) <= a;
    layer4_outputs(5955) <= a or b;
    layer4_outputs(5956) <= not (a xor b);
    layer4_outputs(5957) <= not (a and b);
    layer4_outputs(5958) <= b;
    layer4_outputs(5959) <= a xor b;
    layer4_outputs(5960) <= not b;
    layer4_outputs(5961) <= not b or a;
    layer4_outputs(5962) <= not (a or b);
    layer4_outputs(5963) <= a;
    layer4_outputs(5964) <= not a;
    layer4_outputs(5965) <= b and not a;
    layer4_outputs(5966) <= not b;
    layer4_outputs(5967) <= b;
    layer4_outputs(5968) <= not (a xor b);
    layer4_outputs(5969) <= not b;
    layer4_outputs(5970) <= a and not b;
    layer4_outputs(5971) <= a or b;
    layer4_outputs(5972) <= a and not b;
    layer4_outputs(5973) <= not b;
    layer4_outputs(5974) <= not a or b;
    layer4_outputs(5975) <= b and not a;
    layer4_outputs(5976) <= not b;
    layer4_outputs(5977) <= not b;
    layer4_outputs(5978) <= a;
    layer4_outputs(5979) <= b;
    layer4_outputs(5980) <= b;
    layer4_outputs(5981) <= a and b;
    layer4_outputs(5982) <= not (a xor b);
    layer4_outputs(5983) <= not a or b;
    layer4_outputs(5984) <= a;
    layer4_outputs(5985) <= '0';
    layer4_outputs(5986) <= not a;
    layer4_outputs(5987) <= not (a xor b);
    layer4_outputs(5988) <= a and b;
    layer4_outputs(5989) <= b;
    layer4_outputs(5990) <= not a;
    layer4_outputs(5991) <= not a or b;
    layer4_outputs(5992) <= a and not b;
    layer4_outputs(5993) <= a;
    layer4_outputs(5994) <= a and b;
    layer4_outputs(5995) <= b and not a;
    layer4_outputs(5996) <= not (a or b);
    layer4_outputs(5997) <= not (a and b);
    layer4_outputs(5998) <= a;
    layer4_outputs(5999) <= b;
    layer4_outputs(6000) <= '0';
    layer4_outputs(6001) <= a;
    layer4_outputs(6002) <= '1';
    layer4_outputs(6003) <= not (a and b);
    layer4_outputs(6004) <= a;
    layer4_outputs(6005) <= '1';
    layer4_outputs(6006) <= a and b;
    layer4_outputs(6007) <= '0';
    layer4_outputs(6008) <= a;
    layer4_outputs(6009) <= not b;
    layer4_outputs(6010) <= not a;
    layer4_outputs(6011) <= b and not a;
    layer4_outputs(6012) <= a and not b;
    layer4_outputs(6013) <= '0';
    layer4_outputs(6014) <= not a;
    layer4_outputs(6015) <= b;
    layer4_outputs(6016) <= a;
    layer4_outputs(6017) <= a;
    layer4_outputs(6018) <= not a or b;
    layer4_outputs(6019) <= b;
    layer4_outputs(6020) <= b and not a;
    layer4_outputs(6021) <= a and b;
    layer4_outputs(6022) <= not b;
    layer4_outputs(6023) <= a and not b;
    layer4_outputs(6024) <= a xor b;
    layer4_outputs(6025) <= a xor b;
    layer4_outputs(6026) <= not (a or b);
    layer4_outputs(6027) <= not (a and b);
    layer4_outputs(6028) <= '0';
    layer4_outputs(6029) <= a and not b;
    layer4_outputs(6030) <= not (a xor b);
    layer4_outputs(6031) <= b and not a;
    layer4_outputs(6032) <= not (a xor b);
    layer4_outputs(6033) <= not a;
    layer4_outputs(6034) <= b and not a;
    layer4_outputs(6035) <= not b;
    layer4_outputs(6036) <= not b or a;
    layer4_outputs(6037) <= b;
    layer4_outputs(6038) <= a or b;
    layer4_outputs(6039) <= not b;
    layer4_outputs(6040) <= not a;
    layer4_outputs(6041) <= not b or a;
    layer4_outputs(6042) <= a and not b;
    layer4_outputs(6043) <= a and not b;
    layer4_outputs(6044) <= a;
    layer4_outputs(6045) <= a and not b;
    layer4_outputs(6046) <= not b;
    layer4_outputs(6047) <= not b;
    layer4_outputs(6048) <= not a;
    layer4_outputs(6049) <= a xor b;
    layer4_outputs(6050) <= not a or b;
    layer4_outputs(6051) <= not a or b;
    layer4_outputs(6052) <= a;
    layer4_outputs(6053) <= a;
    layer4_outputs(6054) <= not (a and b);
    layer4_outputs(6055) <= not a;
    layer4_outputs(6056) <= b;
    layer4_outputs(6057) <= b;
    layer4_outputs(6058) <= a;
    layer4_outputs(6059) <= not (a xor b);
    layer4_outputs(6060) <= b;
    layer4_outputs(6061) <= a;
    layer4_outputs(6062) <= a or b;
    layer4_outputs(6063) <= not b or a;
    layer4_outputs(6064) <= not b;
    layer4_outputs(6065) <= not a;
    layer4_outputs(6066) <= '0';
    layer4_outputs(6067) <= not b or a;
    layer4_outputs(6068) <= a or b;
    layer4_outputs(6069) <= b and not a;
    layer4_outputs(6070) <= a;
    layer4_outputs(6071) <= a and not b;
    layer4_outputs(6072) <= '1';
    layer4_outputs(6073) <= a or b;
    layer4_outputs(6074) <= not b;
    layer4_outputs(6075) <= a and b;
    layer4_outputs(6076) <= a and b;
    layer4_outputs(6077) <= a xor b;
    layer4_outputs(6078) <= a xor b;
    layer4_outputs(6079) <= b;
    layer4_outputs(6080) <= not a or b;
    layer4_outputs(6081) <= b;
    layer4_outputs(6082) <= not b;
    layer4_outputs(6083) <= '0';
    layer4_outputs(6084) <= a and b;
    layer4_outputs(6085) <= a and b;
    layer4_outputs(6086) <= a;
    layer4_outputs(6087) <= not (a and b);
    layer4_outputs(6088) <= not a or b;
    layer4_outputs(6089) <= not (a or b);
    layer4_outputs(6090) <= a or b;
    layer4_outputs(6091) <= a;
    layer4_outputs(6092) <= a;
    layer4_outputs(6093) <= a;
    layer4_outputs(6094) <= b;
    layer4_outputs(6095) <= a and b;
    layer4_outputs(6096) <= a or b;
    layer4_outputs(6097) <= a;
    layer4_outputs(6098) <= b;
    layer4_outputs(6099) <= not (a or b);
    layer4_outputs(6100) <= not a;
    layer4_outputs(6101) <= a and b;
    layer4_outputs(6102) <= b and not a;
    layer4_outputs(6103) <= a;
    layer4_outputs(6104) <= a;
    layer4_outputs(6105) <= a;
    layer4_outputs(6106) <= not (a xor b);
    layer4_outputs(6107) <= a;
    layer4_outputs(6108) <= b;
    layer4_outputs(6109) <= not a;
    layer4_outputs(6110) <= not a or b;
    layer4_outputs(6111) <= not b;
    layer4_outputs(6112) <= not b or a;
    layer4_outputs(6113) <= b;
    layer4_outputs(6114) <= not a;
    layer4_outputs(6115) <= not (a or b);
    layer4_outputs(6116) <= b;
    layer4_outputs(6117) <= a xor b;
    layer4_outputs(6118) <= b;
    layer4_outputs(6119) <= not (a and b);
    layer4_outputs(6120) <= b and not a;
    layer4_outputs(6121) <= a;
    layer4_outputs(6122) <= not b;
    layer4_outputs(6123) <= a;
    layer4_outputs(6124) <= not b;
    layer4_outputs(6125) <= not a;
    layer4_outputs(6126) <= not a;
    layer4_outputs(6127) <= a xor b;
    layer4_outputs(6128) <= not (a and b);
    layer4_outputs(6129) <= a and not b;
    layer4_outputs(6130) <= not a;
    layer4_outputs(6131) <= not a;
    layer4_outputs(6132) <= not b;
    layer4_outputs(6133) <= a or b;
    layer4_outputs(6134) <= a;
    layer4_outputs(6135) <= a and b;
    layer4_outputs(6136) <= a;
    layer4_outputs(6137) <= not b;
    layer4_outputs(6138) <= not b;
    layer4_outputs(6139) <= a or b;
    layer4_outputs(6140) <= not (a xor b);
    layer4_outputs(6141) <= a;
    layer4_outputs(6142) <= a xor b;
    layer4_outputs(6143) <= a and not b;
    layer4_outputs(6144) <= a or b;
    layer4_outputs(6145) <= not b or a;
    layer4_outputs(6146) <= b;
    layer4_outputs(6147) <= b;
    layer4_outputs(6148) <= a xor b;
    layer4_outputs(6149) <= a xor b;
    layer4_outputs(6150) <= a xor b;
    layer4_outputs(6151) <= not (a and b);
    layer4_outputs(6152) <= not b or a;
    layer4_outputs(6153) <= not a or b;
    layer4_outputs(6154) <= not a;
    layer4_outputs(6155) <= a and not b;
    layer4_outputs(6156) <= a;
    layer4_outputs(6157) <= b;
    layer4_outputs(6158) <= a xor b;
    layer4_outputs(6159) <= not (a xor b);
    layer4_outputs(6160) <= b;
    layer4_outputs(6161) <= a and b;
    layer4_outputs(6162) <= b;
    layer4_outputs(6163) <= a xor b;
    layer4_outputs(6164) <= b;
    layer4_outputs(6165) <= a;
    layer4_outputs(6166) <= not (a or b);
    layer4_outputs(6167) <= b;
    layer4_outputs(6168) <= not (a and b);
    layer4_outputs(6169) <= b and not a;
    layer4_outputs(6170) <= a or b;
    layer4_outputs(6171) <= a;
    layer4_outputs(6172) <= not b or a;
    layer4_outputs(6173) <= b;
    layer4_outputs(6174) <= b;
    layer4_outputs(6175) <= b and not a;
    layer4_outputs(6176) <= b;
    layer4_outputs(6177) <= a;
    layer4_outputs(6178) <= not (a and b);
    layer4_outputs(6179) <= not a or b;
    layer4_outputs(6180) <= a;
    layer4_outputs(6181) <= b;
    layer4_outputs(6182) <= a xor b;
    layer4_outputs(6183) <= not (a or b);
    layer4_outputs(6184) <= not a;
    layer4_outputs(6185) <= not (a and b);
    layer4_outputs(6186) <= not (a and b);
    layer4_outputs(6187) <= a;
    layer4_outputs(6188) <= b;
    layer4_outputs(6189) <= not a;
    layer4_outputs(6190) <= b;
    layer4_outputs(6191) <= a and not b;
    layer4_outputs(6192) <= not a or b;
    layer4_outputs(6193) <= not a or b;
    layer4_outputs(6194) <= not b;
    layer4_outputs(6195) <= a or b;
    layer4_outputs(6196) <= b and not a;
    layer4_outputs(6197) <= not (a or b);
    layer4_outputs(6198) <= not b;
    layer4_outputs(6199) <= a and not b;
    layer4_outputs(6200) <= not (a and b);
    layer4_outputs(6201) <= not (a xor b);
    layer4_outputs(6202) <= not (a and b);
    layer4_outputs(6203) <= a;
    layer4_outputs(6204) <= not a;
    layer4_outputs(6205) <= not b;
    layer4_outputs(6206) <= not a or b;
    layer4_outputs(6207) <= a and b;
    layer4_outputs(6208) <= b;
    layer4_outputs(6209) <= not (a or b);
    layer4_outputs(6210) <= not a;
    layer4_outputs(6211) <= a xor b;
    layer4_outputs(6212) <= b;
    layer4_outputs(6213) <= b;
    layer4_outputs(6214) <= not (a or b);
    layer4_outputs(6215) <= not (a xor b);
    layer4_outputs(6216) <= a;
    layer4_outputs(6217) <= not b;
    layer4_outputs(6218) <= a;
    layer4_outputs(6219) <= b;
    layer4_outputs(6220) <= not b or a;
    layer4_outputs(6221) <= not (a or b);
    layer4_outputs(6222) <= a;
    layer4_outputs(6223) <= a;
    layer4_outputs(6224) <= not b or a;
    layer4_outputs(6225) <= a;
    layer4_outputs(6226) <= not (a and b);
    layer4_outputs(6227) <= not b or a;
    layer4_outputs(6228) <= a;
    layer4_outputs(6229) <= b;
    layer4_outputs(6230) <= not (a and b);
    layer4_outputs(6231) <= not b;
    layer4_outputs(6232) <= a or b;
    layer4_outputs(6233) <= not b;
    layer4_outputs(6234) <= not (a and b);
    layer4_outputs(6235) <= b;
    layer4_outputs(6236) <= not b or a;
    layer4_outputs(6237) <= not b or a;
    layer4_outputs(6238) <= not b;
    layer4_outputs(6239) <= not b or a;
    layer4_outputs(6240) <= b;
    layer4_outputs(6241) <= a or b;
    layer4_outputs(6242) <= a;
    layer4_outputs(6243) <= not (a or b);
    layer4_outputs(6244) <= b;
    layer4_outputs(6245) <= b;
    layer4_outputs(6246) <= b and not a;
    layer4_outputs(6247) <= not b;
    layer4_outputs(6248) <= not (a xor b);
    layer4_outputs(6249) <= a;
    layer4_outputs(6250) <= not a or b;
    layer4_outputs(6251) <= not a;
    layer4_outputs(6252) <= a and b;
    layer4_outputs(6253) <= not b;
    layer4_outputs(6254) <= not (a and b);
    layer4_outputs(6255) <= a;
    layer4_outputs(6256) <= a and not b;
    layer4_outputs(6257) <= not b or a;
    layer4_outputs(6258) <= a and b;
    layer4_outputs(6259) <= a;
    layer4_outputs(6260) <= not b;
    layer4_outputs(6261) <= '0';
    layer4_outputs(6262) <= a xor b;
    layer4_outputs(6263) <= not a or b;
    layer4_outputs(6264) <= not b or a;
    layer4_outputs(6265) <= a or b;
    layer4_outputs(6266) <= not b;
    layer4_outputs(6267) <= not a;
    layer4_outputs(6268) <= not b;
    layer4_outputs(6269) <= not b or a;
    layer4_outputs(6270) <= a;
    layer4_outputs(6271) <= a xor b;
    layer4_outputs(6272) <= not b or a;
    layer4_outputs(6273) <= not a or b;
    layer4_outputs(6274) <= not (a and b);
    layer4_outputs(6275) <= not (a xor b);
    layer4_outputs(6276) <= b and not a;
    layer4_outputs(6277) <= b;
    layer4_outputs(6278) <= not a;
    layer4_outputs(6279) <= b and not a;
    layer4_outputs(6280) <= not (a xor b);
    layer4_outputs(6281) <= b;
    layer4_outputs(6282) <= b;
    layer4_outputs(6283) <= b and not a;
    layer4_outputs(6284) <= b;
    layer4_outputs(6285) <= a and b;
    layer4_outputs(6286) <= '1';
    layer4_outputs(6287) <= a and b;
    layer4_outputs(6288) <= a and not b;
    layer4_outputs(6289) <= not (a and b);
    layer4_outputs(6290) <= '0';
    layer4_outputs(6291) <= a and not b;
    layer4_outputs(6292) <= a xor b;
    layer4_outputs(6293) <= not b;
    layer4_outputs(6294) <= not (a xor b);
    layer4_outputs(6295) <= not b;
    layer4_outputs(6296) <= a and b;
    layer4_outputs(6297) <= a;
    layer4_outputs(6298) <= b and not a;
    layer4_outputs(6299) <= not b or a;
    layer4_outputs(6300) <= not a;
    layer4_outputs(6301) <= not a;
    layer4_outputs(6302) <= not (a and b);
    layer4_outputs(6303) <= not b;
    layer4_outputs(6304) <= b;
    layer4_outputs(6305) <= b and not a;
    layer4_outputs(6306) <= a and b;
    layer4_outputs(6307) <= not (a xor b);
    layer4_outputs(6308) <= not a;
    layer4_outputs(6309) <= a and not b;
    layer4_outputs(6310) <= a or b;
    layer4_outputs(6311) <= not a or b;
    layer4_outputs(6312) <= not b;
    layer4_outputs(6313) <= '1';
    layer4_outputs(6314) <= not (a xor b);
    layer4_outputs(6315) <= a xor b;
    layer4_outputs(6316) <= b;
    layer4_outputs(6317) <= '0';
    layer4_outputs(6318) <= not (a and b);
    layer4_outputs(6319) <= a or b;
    layer4_outputs(6320) <= not a;
    layer4_outputs(6321) <= b;
    layer4_outputs(6322) <= b;
    layer4_outputs(6323) <= a;
    layer4_outputs(6324) <= '0';
    layer4_outputs(6325) <= not (a xor b);
    layer4_outputs(6326) <= a and not b;
    layer4_outputs(6327) <= not b or a;
    layer4_outputs(6328) <= not a;
    layer4_outputs(6329) <= not a;
    layer4_outputs(6330) <= a xor b;
    layer4_outputs(6331) <= not a;
    layer4_outputs(6332) <= not b;
    layer4_outputs(6333) <= not a;
    layer4_outputs(6334) <= not a;
    layer4_outputs(6335) <= not (a or b);
    layer4_outputs(6336) <= not (a or b);
    layer4_outputs(6337) <= a and not b;
    layer4_outputs(6338) <= not a;
    layer4_outputs(6339) <= a xor b;
    layer4_outputs(6340) <= not (a xor b);
    layer4_outputs(6341) <= not (a xor b);
    layer4_outputs(6342) <= not b;
    layer4_outputs(6343) <= a;
    layer4_outputs(6344) <= not a;
    layer4_outputs(6345) <= not (a or b);
    layer4_outputs(6346) <= not (a xor b);
    layer4_outputs(6347) <= not a or b;
    layer4_outputs(6348) <= a and b;
    layer4_outputs(6349) <= a and b;
    layer4_outputs(6350) <= b;
    layer4_outputs(6351) <= b and not a;
    layer4_outputs(6352) <= b;
    layer4_outputs(6353) <= b and not a;
    layer4_outputs(6354) <= not (a or b);
    layer4_outputs(6355) <= '1';
    layer4_outputs(6356) <= not (a and b);
    layer4_outputs(6357) <= b;
    layer4_outputs(6358) <= a xor b;
    layer4_outputs(6359) <= not b;
    layer4_outputs(6360) <= not (a xor b);
    layer4_outputs(6361) <= not a or b;
    layer4_outputs(6362) <= '1';
    layer4_outputs(6363) <= a and not b;
    layer4_outputs(6364) <= not b or a;
    layer4_outputs(6365) <= not (a and b);
    layer4_outputs(6366) <= a xor b;
    layer4_outputs(6367) <= not a;
    layer4_outputs(6368) <= not b;
    layer4_outputs(6369) <= a and b;
    layer4_outputs(6370) <= a and not b;
    layer4_outputs(6371) <= a and not b;
    layer4_outputs(6372) <= a and not b;
    layer4_outputs(6373) <= b;
    layer4_outputs(6374) <= not a;
    layer4_outputs(6375) <= not (a xor b);
    layer4_outputs(6376) <= a and not b;
    layer4_outputs(6377) <= not (a or b);
    layer4_outputs(6378) <= a or b;
    layer4_outputs(6379) <= '0';
    layer4_outputs(6380) <= not (a or b);
    layer4_outputs(6381) <= not a or b;
    layer4_outputs(6382) <= a xor b;
    layer4_outputs(6383) <= not (a xor b);
    layer4_outputs(6384) <= not (a xor b);
    layer4_outputs(6385) <= a or b;
    layer4_outputs(6386) <= not a;
    layer4_outputs(6387) <= not a or b;
    layer4_outputs(6388) <= a and b;
    layer4_outputs(6389) <= a;
    layer4_outputs(6390) <= not b;
    layer4_outputs(6391) <= a and b;
    layer4_outputs(6392) <= b;
    layer4_outputs(6393) <= not a;
    layer4_outputs(6394) <= not a or b;
    layer4_outputs(6395) <= '0';
    layer4_outputs(6396) <= not (a xor b);
    layer4_outputs(6397) <= not a;
    layer4_outputs(6398) <= b;
    layer4_outputs(6399) <= not b or a;
    layer4_outputs(6400) <= a or b;
    layer4_outputs(6401) <= not b;
    layer4_outputs(6402) <= not a or b;
    layer4_outputs(6403) <= not (a xor b);
    layer4_outputs(6404) <= a and not b;
    layer4_outputs(6405) <= not (a xor b);
    layer4_outputs(6406) <= not b or a;
    layer4_outputs(6407) <= not (a or b);
    layer4_outputs(6408) <= not b;
    layer4_outputs(6409) <= not a or b;
    layer4_outputs(6410) <= not (a or b);
    layer4_outputs(6411) <= not a;
    layer4_outputs(6412) <= not a or b;
    layer4_outputs(6413) <= a;
    layer4_outputs(6414) <= b and not a;
    layer4_outputs(6415) <= not a;
    layer4_outputs(6416) <= not (a xor b);
    layer4_outputs(6417) <= a;
    layer4_outputs(6418) <= not (a xor b);
    layer4_outputs(6419) <= a and b;
    layer4_outputs(6420) <= not b or a;
    layer4_outputs(6421) <= b;
    layer4_outputs(6422) <= not (a xor b);
    layer4_outputs(6423) <= a and b;
    layer4_outputs(6424) <= not a;
    layer4_outputs(6425) <= not b;
    layer4_outputs(6426) <= b;
    layer4_outputs(6427) <= not b;
    layer4_outputs(6428) <= not b;
    layer4_outputs(6429) <= not a;
    layer4_outputs(6430) <= b;
    layer4_outputs(6431) <= a and b;
    layer4_outputs(6432) <= b;
    layer4_outputs(6433) <= b and not a;
    layer4_outputs(6434) <= '1';
    layer4_outputs(6435) <= '0';
    layer4_outputs(6436) <= not (a or b);
    layer4_outputs(6437) <= a;
    layer4_outputs(6438) <= not a or b;
    layer4_outputs(6439) <= a and not b;
    layer4_outputs(6440) <= '1';
    layer4_outputs(6441) <= a or b;
    layer4_outputs(6442) <= not b or a;
    layer4_outputs(6443) <= a;
    layer4_outputs(6444) <= b;
    layer4_outputs(6445) <= b;
    layer4_outputs(6446) <= a and not b;
    layer4_outputs(6447) <= not a;
    layer4_outputs(6448) <= b;
    layer4_outputs(6449) <= not (a or b);
    layer4_outputs(6450) <= a or b;
    layer4_outputs(6451) <= a and not b;
    layer4_outputs(6452) <= a;
    layer4_outputs(6453) <= '0';
    layer4_outputs(6454) <= not a or b;
    layer4_outputs(6455) <= not b;
    layer4_outputs(6456) <= a and not b;
    layer4_outputs(6457) <= b;
    layer4_outputs(6458) <= '0';
    layer4_outputs(6459) <= a and b;
    layer4_outputs(6460) <= b and not a;
    layer4_outputs(6461) <= not b;
    layer4_outputs(6462) <= a xor b;
    layer4_outputs(6463) <= not b or a;
    layer4_outputs(6464) <= not (a or b);
    layer4_outputs(6465) <= a;
    layer4_outputs(6466) <= a or b;
    layer4_outputs(6467) <= not b;
    layer4_outputs(6468) <= not b or a;
    layer4_outputs(6469) <= a;
    layer4_outputs(6470) <= not b;
    layer4_outputs(6471) <= not (a xor b);
    layer4_outputs(6472) <= not (a xor b);
    layer4_outputs(6473) <= not b or a;
    layer4_outputs(6474) <= not (a or b);
    layer4_outputs(6475) <= b;
    layer4_outputs(6476) <= a or b;
    layer4_outputs(6477) <= not b;
    layer4_outputs(6478) <= a;
    layer4_outputs(6479) <= a;
    layer4_outputs(6480) <= a;
    layer4_outputs(6481) <= not b;
    layer4_outputs(6482) <= not b or a;
    layer4_outputs(6483) <= a or b;
    layer4_outputs(6484) <= a and b;
    layer4_outputs(6485) <= a;
    layer4_outputs(6486) <= not a;
    layer4_outputs(6487) <= a xor b;
    layer4_outputs(6488) <= not (a or b);
    layer4_outputs(6489) <= b;
    layer4_outputs(6490) <= a;
    layer4_outputs(6491) <= not (a and b);
    layer4_outputs(6492) <= not b;
    layer4_outputs(6493) <= a xor b;
    layer4_outputs(6494) <= not (a xor b);
    layer4_outputs(6495) <= '0';
    layer4_outputs(6496) <= '1';
    layer4_outputs(6497) <= not (a or b);
    layer4_outputs(6498) <= not b or a;
    layer4_outputs(6499) <= not (a xor b);
    layer4_outputs(6500) <= a and not b;
    layer4_outputs(6501) <= not b;
    layer4_outputs(6502) <= b and not a;
    layer4_outputs(6503) <= not a or b;
    layer4_outputs(6504) <= not b;
    layer4_outputs(6505) <= not b;
    layer4_outputs(6506) <= a;
    layer4_outputs(6507) <= not a;
    layer4_outputs(6508) <= b;
    layer4_outputs(6509) <= not a;
    layer4_outputs(6510) <= b;
    layer4_outputs(6511) <= a and b;
    layer4_outputs(6512) <= a;
    layer4_outputs(6513) <= a;
    layer4_outputs(6514) <= not a or b;
    layer4_outputs(6515) <= not a or b;
    layer4_outputs(6516) <= b;
    layer4_outputs(6517) <= not a or b;
    layer4_outputs(6518) <= not b or a;
    layer4_outputs(6519) <= not b;
    layer4_outputs(6520) <= not a or b;
    layer4_outputs(6521) <= a or b;
    layer4_outputs(6522) <= a;
    layer4_outputs(6523) <= not b or a;
    layer4_outputs(6524) <= b and not a;
    layer4_outputs(6525) <= b;
    layer4_outputs(6526) <= a xor b;
    layer4_outputs(6527) <= a and not b;
    layer4_outputs(6528) <= b;
    layer4_outputs(6529) <= a and b;
    layer4_outputs(6530) <= a or b;
    layer4_outputs(6531) <= not a;
    layer4_outputs(6532) <= not a;
    layer4_outputs(6533) <= b;
    layer4_outputs(6534) <= '1';
    layer4_outputs(6535) <= a and b;
    layer4_outputs(6536) <= not b or a;
    layer4_outputs(6537) <= b;
    layer4_outputs(6538) <= b;
    layer4_outputs(6539) <= b and not a;
    layer4_outputs(6540) <= not a;
    layer4_outputs(6541) <= not b;
    layer4_outputs(6542) <= a or b;
    layer4_outputs(6543) <= a xor b;
    layer4_outputs(6544) <= a xor b;
    layer4_outputs(6545) <= not (a or b);
    layer4_outputs(6546) <= a xor b;
    layer4_outputs(6547) <= not (a and b);
    layer4_outputs(6548) <= a and not b;
    layer4_outputs(6549) <= a and b;
    layer4_outputs(6550) <= a;
    layer4_outputs(6551) <= not b;
    layer4_outputs(6552) <= a or b;
    layer4_outputs(6553) <= a and b;
    layer4_outputs(6554) <= '1';
    layer4_outputs(6555) <= a;
    layer4_outputs(6556) <= a and b;
    layer4_outputs(6557) <= a xor b;
    layer4_outputs(6558) <= not (a xor b);
    layer4_outputs(6559) <= not b;
    layer4_outputs(6560) <= a;
    layer4_outputs(6561) <= not a;
    layer4_outputs(6562) <= not a or b;
    layer4_outputs(6563) <= a or b;
    layer4_outputs(6564) <= a and b;
    layer4_outputs(6565) <= b and not a;
    layer4_outputs(6566) <= not (a or b);
    layer4_outputs(6567) <= not a;
    layer4_outputs(6568) <= a and not b;
    layer4_outputs(6569) <= a and b;
    layer4_outputs(6570) <= a and b;
    layer4_outputs(6571) <= not a or b;
    layer4_outputs(6572) <= not (a or b);
    layer4_outputs(6573) <= '1';
    layer4_outputs(6574) <= a xor b;
    layer4_outputs(6575) <= not b;
    layer4_outputs(6576) <= not b or a;
    layer4_outputs(6577) <= a;
    layer4_outputs(6578) <= a xor b;
    layer4_outputs(6579) <= a or b;
    layer4_outputs(6580) <= not b or a;
    layer4_outputs(6581) <= a xor b;
    layer4_outputs(6582) <= b and not a;
    layer4_outputs(6583) <= '1';
    layer4_outputs(6584) <= not b;
    layer4_outputs(6585) <= not (a xor b);
    layer4_outputs(6586) <= a;
    layer4_outputs(6587) <= a xor b;
    layer4_outputs(6588) <= not a;
    layer4_outputs(6589) <= b and not a;
    layer4_outputs(6590) <= not (a or b);
    layer4_outputs(6591) <= not a or b;
    layer4_outputs(6592) <= a and b;
    layer4_outputs(6593) <= a and b;
    layer4_outputs(6594) <= not b;
    layer4_outputs(6595) <= not a or b;
    layer4_outputs(6596) <= a xor b;
    layer4_outputs(6597) <= '1';
    layer4_outputs(6598) <= not (a and b);
    layer4_outputs(6599) <= b;
    layer4_outputs(6600) <= b;
    layer4_outputs(6601) <= not (a and b);
    layer4_outputs(6602) <= not (a xor b);
    layer4_outputs(6603) <= a and not b;
    layer4_outputs(6604) <= a and b;
    layer4_outputs(6605) <= not a or b;
    layer4_outputs(6606) <= not b;
    layer4_outputs(6607) <= not b or a;
    layer4_outputs(6608) <= a or b;
    layer4_outputs(6609) <= a and not b;
    layer4_outputs(6610) <= not (a xor b);
    layer4_outputs(6611) <= not b;
    layer4_outputs(6612) <= a;
    layer4_outputs(6613) <= a and b;
    layer4_outputs(6614) <= not a;
    layer4_outputs(6615) <= not (a xor b);
    layer4_outputs(6616) <= not a;
    layer4_outputs(6617) <= '1';
    layer4_outputs(6618) <= a;
    layer4_outputs(6619) <= a and not b;
    layer4_outputs(6620) <= not b;
    layer4_outputs(6621) <= '1';
    layer4_outputs(6622) <= a and b;
    layer4_outputs(6623) <= not b;
    layer4_outputs(6624) <= '1';
    layer4_outputs(6625) <= a and not b;
    layer4_outputs(6626) <= not (a or b);
    layer4_outputs(6627) <= not a;
    layer4_outputs(6628) <= a or b;
    layer4_outputs(6629) <= a and not b;
    layer4_outputs(6630) <= a or b;
    layer4_outputs(6631) <= a and not b;
    layer4_outputs(6632) <= a;
    layer4_outputs(6633) <= a xor b;
    layer4_outputs(6634) <= not a;
    layer4_outputs(6635) <= a and not b;
    layer4_outputs(6636) <= not a;
    layer4_outputs(6637) <= not a;
    layer4_outputs(6638) <= '1';
    layer4_outputs(6639) <= not b or a;
    layer4_outputs(6640) <= b and not a;
    layer4_outputs(6641) <= a xor b;
    layer4_outputs(6642) <= not a or b;
    layer4_outputs(6643) <= not a;
    layer4_outputs(6644) <= not b or a;
    layer4_outputs(6645) <= '0';
    layer4_outputs(6646) <= b;
    layer4_outputs(6647) <= not a;
    layer4_outputs(6648) <= not a or b;
    layer4_outputs(6649) <= not (a xor b);
    layer4_outputs(6650) <= not a or b;
    layer4_outputs(6651) <= not a;
    layer4_outputs(6652) <= not a;
    layer4_outputs(6653) <= not a;
    layer4_outputs(6654) <= a and not b;
    layer4_outputs(6655) <= a or b;
    layer4_outputs(6656) <= not b;
    layer4_outputs(6657) <= not (a or b);
    layer4_outputs(6658) <= not (a and b);
    layer4_outputs(6659) <= not (a and b);
    layer4_outputs(6660) <= not a;
    layer4_outputs(6661) <= a;
    layer4_outputs(6662) <= b and not a;
    layer4_outputs(6663) <= not (a xor b);
    layer4_outputs(6664) <= not a or b;
    layer4_outputs(6665) <= not b;
    layer4_outputs(6666) <= b;
    layer4_outputs(6667) <= a and not b;
    layer4_outputs(6668) <= not b;
    layer4_outputs(6669) <= not b or a;
    layer4_outputs(6670) <= not (a or b);
    layer4_outputs(6671) <= b;
    layer4_outputs(6672) <= not b;
    layer4_outputs(6673) <= a and not b;
    layer4_outputs(6674) <= a or b;
    layer4_outputs(6675) <= b;
    layer4_outputs(6676) <= b and not a;
    layer4_outputs(6677) <= b;
    layer4_outputs(6678) <= not (a xor b);
    layer4_outputs(6679) <= a;
    layer4_outputs(6680) <= a and not b;
    layer4_outputs(6681) <= not (a or b);
    layer4_outputs(6682) <= b;
    layer4_outputs(6683) <= not (a or b);
    layer4_outputs(6684) <= not b or a;
    layer4_outputs(6685) <= not a or b;
    layer4_outputs(6686) <= not b or a;
    layer4_outputs(6687) <= not a;
    layer4_outputs(6688) <= not b;
    layer4_outputs(6689) <= not (a and b);
    layer4_outputs(6690) <= not b;
    layer4_outputs(6691) <= a or b;
    layer4_outputs(6692) <= not (a xor b);
    layer4_outputs(6693) <= not b;
    layer4_outputs(6694) <= a and b;
    layer4_outputs(6695) <= not b or a;
    layer4_outputs(6696) <= not (a and b);
    layer4_outputs(6697) <= not a;
    layer4_outputs(6698) <= a xor b;
    layer4_outputs(6699) <= not (a xor b);
    layer4_outputs(6700) <= not b;
    layer4_outputs(6701) <= not a or b;
    layer4_outputs(6702) <= not (a or b);
    layer4_outputs(6703) <= b and not a;
    layer4_outputs(6704) <= not a or b;
    layer4_outputs(6705) <= b and not a;
    layer4_outputs(6706) <= not a;
    layer4_outputs(6707) <= not b;
    layer4_outputs(6708) <= not (a or b);
    layer4_outputs(6709) <= a;
    layer4_outputs(6710) <= a and b;
    layer4_outputs(6711) <= not (a xor b);
    layer4_outputs(6712) <= not (a and b);
    layer4_outputs(6713) <= a and not b;
    layer4_outputs(6714) <= a and not b;
    layer4_outputs(6715) <= not b;
    layer4_outputs(6716) <= '1';
    layer4_outputs(6717) <= not a;
    layer4_outputs(6718) <= not a;
    layer4_outputs(6719) <= not b;
    layer4_outputs(6720) <= not a;
    layer4_outputs(6721) <= b;
    layer4_outputs(6722) <= a and not b;
    layer4_outputs(6723) <= not (a or b);
    layer4_outputs(6724) <= not (a or b);
    layer4_outputs(6725) <= not (a and b);
    layer4_outputs(6726) <= a or b;
    layer4_outputs(6727) <= not a or b;
    layer4_outputs(6728) <= not a;
    layer4_outputs(6729) <= a and not b;
    layer4_outputs(6730) <= a;
    layer4_outputs(6731) <= '0';
    layer4_outputs(6732) <= not (a or b);
    layer4_outputs(6733) <= a xor b;
    layer4_outputs(6734) <= not a;
    layer4_outputs(6735) <= not a or b;
    layer4_outputs(6736) <= not a;
    layer4_outputs(6737) <= not (a xor b);
    layer4_outputs(6738) <= not a;
    layer4_outputs(6739) <= not (a and b);
    layer4_outputs(6740) <= not (a xor b);
    layer4_outputs(6741) <= not b;
    layer4_outputs(6742) <= a or b;
    layer4_outputs(6743) <= a and not b;
    layer4_outputs(6744) <= '0';
    layer4_outputs(6745) <= not b;
    layer4_outputs(6746) <= not (a xor b);
    layer4_outputs(6747) <= a;
    layer4_outputs(6748) <= not b;
    layer4_outputs(6749) <= a;
    layer4_outputs(6750) <= '0';
    layer4_outputs(6751) <= a;
    layer4_outputs(6752) <= not a;
    layer4_outputs(6753) <= a;
    layer4_outputs(6754) <= b;
    layer4_outputs(6755) <= b;
    layer4_outputs(6756) <= a and not b;
    layer4_outputs(6757) <= not b;
    layer4_outputs(6758) <= a and not b;
    layer4_outputs(6759) <= b and not a;
    layer4_outputs(6760) <= not b or a;
    layer4_outputs(6761) <= a;
    layer4_outputs(6762) <= not a or b;
    layer4_outputs(6763) <= not (a xor b);
    layer4_outputs(6764) <= not (a or b);
    layer4_outputs(6765) <= not a;
    layer4_outputs(6766) <= not (a and b);
    layer4_outputs(6767) <= not b;
    layer4_outputs(6768) <= b;
    layer4_outputs(6769) <= not (a or b);
    layer4_outputs(6770) <= not (a or b);
    layer4_outputs(6771) <= a and not b;
    layer4_outputs(6772) <= not b;
    layer4_outputs(6773) <= not (a or b);
    layer4_outputs(6774) <= a and not b;
    layer4_outputs(6775) <= b;
    layer4_outputs(6776) <= a and not b;
    layer4_outputs(6777) <= not a;
    layer4_outputs(6778) <= '0';
    layer4_outputs(6779) <= b;
    layer4_outputs(6780) <= not (a and b);
    layer4_outputs(6781) <= b and not a;
    layer4_outputs(6782) <= b and not a;
    layer4_outputs(6783) <= b and not a;
    layer4_outputs(6784) <= a;
    layer4_outputs(6785) <= a and b;
    layer4_outputs(6786) <= not (a and b);
    layer4_outputs(6787) <= b;
    layer4_outputs(6788) <= b and not a;
    layer4_outputs(6789) <= not b;
    layer4_outputs(6790) <= not (a and b);
    layer4_outputs(6791) <= not a;
    layer4_outputs(6792) <= a xor b;
    layer4_outputs(6793) <= not b or a;
    layer4_outputs(6794) <= b and not a;
    layer4_outputs(6795) <= not (a or b);
    layer4_outputs(6796) <= not a;
    layer4_outputs(6797) <= a and not b;
    layer4_outputs(6798) <= a and not b;
    layer4_outputs(6799) <= a and b;
    layer4_outputs(6800) <= a;
    layer4_outputs(6801) <= not b;
    layer4_outputs(6802) <= a and b;
    layer4_outputs(6803) <= a or b;
    layer4_outputs(6804) <= a or b;
    layer4_outputs(6805) <= not a;
    layer4_outputs(6806) <= a and not b;
    layer4_outputs(6807) <= a;
    layer4_outputs(6808) <= not a;
    layer4_outputs(6809) <= not b;
    layer4_outputs(6810) <= a;
    layer4_outputs(6811) <= not (a xor b);
    layer4_outputs(6812) <= not a;
    layer4_outputs(6813) <= not a;
    layer4_outputs(6814) <= a and b;
    layer4_outputs(6815) <= not (a xor b);
    layer4_outputs(6816) <= b and not a;
    layer4_outputs(6817) <= not (a and b);
    layer4_outputs(6818) <= a xor b;
    layer4_outputs(6819) <= not (a and b);
    layer4_outputs(6820) <= a;
    layer4_outputs(6821) <= a;
    layer4_outputs(6822) <= '0';
    layer4_outputs(6823) <= a and b;
    layer4_outputs(6824) <= a xor b;
    layer4_outputs(6825) <= a and b;
    layer4_outputs(6826) <= not a or b;
    layer4_outputs(6827) <= not a or b;
    layer4_outputs(6828) <= not (a or b);
    layer4_outputs(6829) <= b;
    layer4_outputs(6830) <= a xor b;
    layer4_outputs(6831) <= not a or b;
    layer4_outputs(6832) <= not b;
    layer4_outputs(6833) <= not b or a;
    layer4_outputs(6834) <= a;
    layer4_outputs(6835) <= not a;
    layer4_outputs(6836) <= a and not b;
    layer4_outputs(6837) <= b;
    layer4_outputs(6838) <= not (a or b);
    layer4_outputs(6839) <= not (a xor b);
    layer4_outputs(6840) <= not a;
    layer4_outputs(6841) <= not (a or b);
    layer4_outputs(6842) <= not (a xor b);
    layer4_outputs(6843) <= a;
    layer4_outputs(6844) <= not b or a;
    layer4_outputs(6845) <= '0';
    layer4_outputs(6846) <= a or b;
    layer4_outputs(6847) <= b;
    layer4_outputs(6848) <= not (a xor b);
    layer4_outputs(6849) <= a;
    layer4_outputs(6850) <= a;
    layer4_outputs(6851) <= a;
    layer4_outputs(6852) <= not a;
    layer4_outputs(6853) <= not a;
    layer4_outputs(6854) <= b;
    layer4_outputs(6855) <= not b;
    layer4_outputs(6856) <= a or b;
    layer4_outputs(6857) <= a;
    layer4_outputs(6858) <= not b;
    layer4_outputs(6859) <= b;
    layer4_outputs(6860) <= a and not b;
    layer4_outputs(6861) <= b;
    layer4_outputs(6862) <= '0';
    layer4_outputs(6863) <= b and not a;
    layer4_outputs(6864) <= b;
    layer4_outputs(6865) <= b and not a;
    layer4_outputs(6866) <= a and not b;
    layer4_outputs(6867) <= not b;
    layer4_outputs(6868) <= a and b;
    layer4_outputs(6869) <= not b;
    layer4_outputs(6870) <= a and not b;
    layer4_outputs(6871) <= not (a xor b);
    layer4_outputs(6872) <= not a;
    layer4_outputs(6873) <= not a or b;
    layer4_outputs(6874) <= b;
    layer4_outputs(6875) <= a or b;
    layer4_outputs(6876) <= a;
    layer4_outputs(6877) <= not a or b;
    layer4_outputs(6878) <= not a or b;
    layer4_outputs(6879) <= not b;
    layer4_outputs(6880) <= not b;
    layer4_outputs(6881) <= not b or a;
    layer4_outputs(6882) <= b;
    layer4_outputs(6883) <= not a;
    layer4_outputs(6884) <= '0';
    layer4_outputs(6885) <= not a;
    layer4_outputs(6886) <= a xor b;
    layer4_outputs(6887) <= a and b;
    layer4_outputs(6888) <= a;
    layer4_outputs(6889) <= a;
    layer4_outputs(6890) <= not a or b;
    layer4_outputs(6891) <= not (a and b);
    layer4_outputs(6892) <= a;
    layer4_outputs(6893) <= not b;
    layer4_outputs(6894) <= not a;
    layer4_outputs(6895) <= not (a and b);
    layer4_outputs(6896) <= b;
    layer4_outputs(6897) <= not (a or b);
    layer4_outputs(6898) <= not (a xor b);
    layer4_outputs(6899) <= a and not b;
    layer4_outputs(6900) <= not a;
    layer4_outputs(6901) <= a;
    layer4_outputs(6902) <= not b;
    layer4_outputs(6903) <= not b;
    layer4_outputs(6904) <= not b;
    layer4_outputs(6905) <= not a or b;
    layer4_outputs(6906) <= a and b;
    layer4_outputs(6907) <= not b;
    layer4_outputs(6908) <= b;
    layer4_outputs(6909) <= a;
    layer4_outputs(6910) <= a xor b;
    layer4_outputs(6911) <= a;
    layer4_outputs(6912) <= not (a xor b);
    layer4_outputs(6913) <= a xor b;
    layer4_outputs(6914) <= b;
    layer4_outputs(6915) <= a or b;
    layer4_outputs(6916) <= not b;
    layer4_outputs(6917) <= a;
    layer4_outputs(6918) <= not a;
    layer4_outputs(6919) <= not (a xor b);
    layer4_outputs(6920) <= not (a and b);
    layer4_outputs(6921) <= a;
    layer4_outputs(6922) <= a;
    layer4_outputs(6923) <= a;
    layer4_outputs(6924) <= a;
    layer4_outputs(6925) <= '0';
    layer4_outputs(6926) <= not b;
    layer4_outputs(6927) <= not b or a;
    layer4_outputs(6928) <= not a;
    layer4_outputs(6929) <= not a or b;
    layer4_outputs(6930) <= not b;
    layer4_outputs(6931) <= not b;
    layer4_outputs(6932) <= a and not b;
    layer4_outputs(6933) <= a and b;
    layer4_outputs(6934) <= b;
    layer4_outputs(6935) <= b and not a;
    layer4_outputs(6936) <= b;
    layer4_outputs(6937) <= not (a xor b);
    layer4_outputs(6938) <= not (a xor b);
    layer4_outputs(6939) <= not (a and b);
    layer4_outputs(6940) <= a and b;
    layer4_outputs(6941) <= a;
    layer4_outputs(6942) <= not a;
    layer4_outputs(6943) <= b and not a;
    layer4_outputs(6944) <= a and b;
    layer4_outputs(6945) <= not b or a;
    layer4_outputs(6946) <= not a;
    layer4_outputs(6947) <= not b or a;
    layer4_outputs(6948) <= b;
    layer4_outputs(6949) <= not b or a;
    layer4_outputs(6950) <= b;
    layer4_outputs(6951) <= not (a and b);
    layer4_outputs(6952) <= b and not a;
    layer4_outputs(6953) <= b and not a;
    layer4_outputs(6954) <= a;
    layer4_outputs(6955) <= not a or b;
    layer4_outputs(6956) <= a;
    layer4_outputs(6957) <= not a or b;
    layer4_outputs(6958) <= a and b;
    layer4_outputs(6959) <= not a or b;
    layer4_outputs(6960) <= not a;
    layer4_outputs(6961) <= '0';
    layer4_outputs(6962) <= a;
    layer4_outputs(6963) <= a and not b;
    layer4_outputs(6964) <= a;
    layer4_outputs(6965) <= not a;
    layer4_outputs(6966) <= not (a xor b);
    layer4_outputs(6967) <= not (a and b);
    layer4_outputs(6968) <= not (a xor b);
    layer4_outputs(6969) <= a;
    layer4_outputs(6970) <= a and b;
    layer4_outputs(6971) <= not (a and b);
    layer4_outputs(6972) <= not a;
    layer4_outputs(6973) <= '1';
    layer4_outputs(6974) <= b;
    layer4_outputs(6975) <= not (a xor b);
    layer4_outputs(6976) <= '0';
    layer4_outputs(6977) <= not (a or b);
    layer4_outputs(6978) <= a xor b;
    layer4_outputs(6979) <= a;
    layer4_outputs(6980) <= not a;
    layer4_outputs(6981) <= b;
    layer4_outputs(6982) <= not a or b;
    layer4_outputs(6983) <= b and not a;
    layer4_outputs(6984) <= a xor b;
    layer4_outputs(6985) <= not (a xor b);
    layer4_outputs(6986) <= not (a or b);
    layer4_outputs(6987) <= b;
    layer4_outputs(6988) <= not (a or b);
    layer4_outputs(6989) <= not b;
    layer4_outputs(6990) <= a;
    layer4_outputs(6991) <= b;
    layer4_outputs(6992) <= not (a or b);
    layer4_outputs(6993) <= not (a or b);
    layer4_outputs(6994) <= not a;
    layer4_outputs(6995) <= a or b;
    layer4_outputs(6996) <= not b;
    layer4_outputs(6997) <= b;
    layer4_outputs(6998) <= a or b;
    layer4_outputs(6999) <= b;
    layer4_outputs(7000) <= a and b;
    layer4_outputs(7001) <= not a;
    layer4_outputs(7002) <= a or b;
    layer4_outputs(7003) <= not a;
    layer4_outputs(7004) <= not b or a;
    layer4_outputs(7005) <= not (a and b);
    layer4_outputs(7006) <= not b;
    layer4_outputs(7007) <= not a;
    layer4_outputs(7008) <= a;
    layer4_outputs(7009) <= a;
    layer4_outputs(7010) <= a xor b;
    layer4_outputs(7011) <= not (a xor b);
    layer4_outputs(7012) <= b;
    layer4_outputs(7013) <= a and b;
    layer4_outputs(7014) <= '1';
    layer4_outputs(7015) <= not (a and b);
    layer4_outputs(7016) <= not b or a;
    layer4_outputs(7017) <= a and b;
    layer4_outputs(7018) <= a;
    layer4_outputs(7019) <= not a or b;
    layer4_outputs(7020) <= a;
    layer4_outputs(7021) <= a and b;
    layer4_outputs(7022) <= not a;
    layer4_outputs(7023) <= not b or a;
    layer4_outputs(7024) <= a or b;
    layer4_outputs(7025) <= not (a and b);
    layer4_outputs(7026) <= a and b;
    layer4_outputs(7027) <= not a or b;
    layer4_outputs(7028) <= not a;
    layer4_outputs(7029) <= '0';
    layer4_outputs(7030) <= not b;
    layer4_outputs(7031) <= not (a or b);
    layer4_outputs(7032) <= b;
    layer4_outputs(7033) <= not a;
    layer4_outputs(7034) <= '1';
    layer4_outputs(7035) <= a and not b;
    layer4_outputs(7036) <= not a;
    layer4_outputs(7037) <= not (a xor b);
    layer4_outputs(7038) <= a and b;
    layer4_outputs(7039) <= not b or a;
    layer4_outputs(7040) <= not a;
    layer4_outputs(7041) <= a and not b;
    layer4_outputs(7042) <= not b or a;
    layer4_outputs(7043) <= a or b;
    layer4_outputs(7044) <= a and not b;
    layer4_outputs(7045) <= a and b;
    layer4_outputs(7046) <= not a or b;
    layer4_outputs(7047) <= a and b;
    layer4_outputs(7048) <= b;
    layer4_outputs(7049) <= a and b;
    layer4_outputs(7050) <= not (a or b);
    layer4_outputs(7051) <= not b;
    layer4_outputs(7052) <= '0';
    layer4_outputs(7053) <= not b;
    layer4_outputs(7054) <= not a;
    layer4_outputs(7055) <= not b;
    layer4_outputs(7056) <= not a or b;
    layer4_outputs(7057) <= not b or a;
    layer4_outputs(7058) <= not b;
    layer4_outputs(7059) <= not b;
    layer4_outputs(7060) <= not (a xor b);
    layer4_outputs(7061) <= not (a and b);
    layer4_outputs(7062) <= a or b;
    layer4_outputs(7063) <= not a;
    layer4_outputs(7064) <= a;
    layer4_outputs(7065) <= b;
    layer4_outputs(7066) <= not (a and b);
    layer4_outputs(7067) <= a;
    layer4_outputs(7068) <= not a or b;
    layer4_outputs(7069) <= a or b;
    layer4_outputs(7070) <= b;
    layer4_outputs(7071) <= b;
    layer4_outputs(7072) <= not (a or b);
    layer4_outputs(7073) <= b;
    layer4_outputs(7074) <= not (a and b);
    layer4_outputs(7075) <= a;
    layer4_outputs(7076) <= b;
    layer4_outputs(7077) <= a;
    layer4_outputs(7078) <= not (a or b);
    layer4_outputs(7079) <= not (a and b);
    layer4_outputs(7080) <= a xor b;
    layer4_outputs(7081) <= a;
    layer4_outputs(7082) <= a or b;
    layer4_outputs(7083) <= b and not a;
    layer4_outputs(7084) <= not (a or b);
    layer4_outputs(7085) <= not b;
    layer4_outputs(7086) <= not b;
    layer4_outputs(7087) <= a;
    layer4_outputs(7088) <= '0';
    layer4_outputs(7089) <= a;
    layer4_outputs(7090) <= not a or b;
    layer4_outputs(7091) <= not (a or b);
    layer4_outputs(7092) <= b;
    layer4_outputs(7093) <= a or b;
    layer4_outputs(7094) <= not b or a;
    layer4_outputs(7095) <= not (a xor b);
    layer4_outputs(7096) <= b;
    layer4_outputs(7097) <= b;
    layer4_outputs(7098) <= not (a or b);
    layer4_outputs(7099) <= a and not b;
    layer4_outputs(7100) <= a and b;
    layer4_outputs(7101) <= not b or a;
    layer4_outputs(7102) <= '0';
    layer4_outputs(7103) <= not (a or b);
    layer4_outputs(7104) <= a or b;
    layer4_outputs(7105) <= a and not b;
    layer4_outputs(7106) <= a and not b;
    layer4_outputs(7107) <= b;
    layer4_outputs(7108) <= not b;
    layer4_outputs(7109) <= b;
    layer4_outputs(7110) <= a;
    layer4_outputs(7111) <= not (a and b);
    layer4_outputs(7112) <= not a;
    layer4_outputs(7113) <= b;
    layer4_outputs(7114) <= not (a xor b);
    layer4_outputs(7115) <= not (a and b);
    layer4_outputs(7116) <= a and b;
    layer4_outputs(7117) <= not b;
    layer4_outputs(7118) <= a;
    layer4_outputs(7119) <= a xor b;
    layer4_outputs(7120) <= a;
    layer4_outputs(7121) <= a;
    layer4_outputs(7122) <= a and not b;
    layer4_outputs(7123) <= not b or a;
    layer4_outputs(7124) <= not a;
    layer4_outputs(7125) <= a and b;
    layer4_outputs(7126) <= b;
    layer4_outputs(7127) <= a and not b;
    layer4_outputs(7128) <= not (a or b);
    layer4_outputs(7129) <= not a;
    layer4_outputs(7130) <= '0';
    layer4_outputs(7131) <= a and b;
    layer4_outputs(7132) <= b;
    layer4_outputs(7133) <= b;
    layer4_outputs(7134) <= not b;
    layer4_outputs(7135) <= not b or a;
    layer4_outputs(7136) <= a xor b;
    layer4_outputs(7137) <= a or b;
    layer4_outputs(7138) <= a and b;
    layer4_outputs(7139) <= b;
    layer4_outputs(7140) <= a;
    layer4_outputs(7141) <= not (a and b);
    layer4_outputs(7142) <= b and not a;
    layer4_outputs(7143) <= a and b;
    layer4_outputs(7144) <= not a;
    layer4_outputs(7145) <= not (a or b);
    layer4_outputs(7146) <= a and b;
    layer4_outputs(7147) <= a;
    layer4_outputs(7148) <= not (a or b);
    layer4_outputs(7149) <= a and b;
    layer4_outputs(7150) <= not b;
    layer4_outputs(7151) <= not a;
    layer4_outputs(7152) <= not b;
    layer4_outputs(7153) <= a xor b;
    layer4_outputs(7154) <= not a or b;
    layer4_outputs(7155) <= not a;
    layer4_outputs(7156) <= b;
    layer4_outputs(7157) <= a or b;
    layer4_outputs(7158) <= a;
    layer4_outputs(7159) <= '1';
    layer4_outputs(7160) <= not b;
    layer4_outputs(7161) <= b;
    layer4_outputs(7162) <= not b;
    layer4_outputs(7163) <= b;
    layer4_outputs(7164) <= '0';
    layer4_outputs(7165) <= a or b;
    layer4_outputs(7166) <= b;
    layer4_outputs(7167) <= not (a or b);
    layer4_outputs(7168) <= not b;
    layer4_outputs(7169) <= not b;
    layer4_outputs(7170) <= a;
    layer4_outputs(7171) <= b and not a;
    layer4_outputs(7172) <= a;
    layer4_outputs(7173) <= not a;
    layer4_outputs(7174) <= b and not a;
    layer4_outputs(7175) <= not b;
    layer4_outputs(7176) <= a;
    layer4_outputs(7177) <= not (a or b);
    layer4_outputs(7178) <= b;
    layer4_outputs(7179) <= '1';
    layer4_outputs(7180) <= not b or a;
    layer4_outputs(7181) <= not (a and b);
    layer4_outputs(7182) <= not a;
    layer4_outputs(7183) <= a and b;
    layer4_outputs(7184) <= not a;
    layer4_outputs(7185) <= b;
    layer4_outputs(7186) <= a or b;
    layer4_outputs(7187) <= not (a or b);
    layer4_outputs(7188) <= b;
    layer4_outputs(7189) <= b;
    layer4_outputs(7190) <= not b or a;
    layer4_outputs(7191) <= '0';
    layer4_outputs(7192) <= b;
    layer4_outputs(7193) <= not (a or b);
    layer4_outputs(7194) <= not a or b;
    layer4_outputs(7195) <= '1';
    layer4_outputs(7196) <= '0';
    layer4_outputs(7197) <= '1';
    layer4_outputs(7198) <= b;
    layer4_outputs(7199) <= not (a xor b);
    layer4_outputs(7200) <= not a or b;
    layer4_outputs(7201) <= a;
    layer4_outputs(7202) <= not a;
    layer4_outputs(7203) <= b and not a;
    layer4_outputs(7204) <= not b or a;
    layer4_outputs(7205) <= not a;
    layer4_outputs(7206) <= a;
    layer4_outputs(7207) <= not a or b;
    layer4_outputs(7208) <= a and b;
    layer4_outputs(7209) <= not a;
    layer4_outputs(7210) <= not (a xor b);
    layer4_outputs(7211) <= not (a xor b);
    layer4_outputs(7212) <= not a or b;
    layer4_outputs(7213) <= a;
    layer4_outputs(7214) <= b;
    layer4_outputs(7215) <= not b;
    layer4_outputs(7216) <= not (a or b);
    layer4_outputs(7217) <= not a or b;
    layer4_outputs(7218) <= not (a and b);
    layer4_outputs(7219) <= a xor b;
    layer4_outputs(7220) <= a xor b;
    layer4_outputs(7221) <= b;
    layer4_outputs(7222) <= not b;
    layer4_outputs(7223) <= b and not a;
    layer4_outputs(7224) <= a and b;
    layer4_outputs(7225) <= not b or a;
    layer4_outputs(7226) <= a;
    layer4_outputs(7227) <= not b;
    layer4_outputs(7228) <= not a or b;
    layer4_outputs(7229) <= a;
    layer4_outputs(7230) <= b and not a;
    layer4_outputs(7231) <= not b or a;
    layer4_outputs(7232) <= a;
    layer4_outputs(7233) <= not (a or b);
    layer4_outputs(7234) <= not a;
    layer4_outputs(7235) <= not b;
    layer4_outputs(7236) <= not b;
    layer4_outputs(7237) <= b;
    layer4_outputs(7238) <= not b or a;
    layer4_outputs(7239) <= a;
    layer4_outputs(7240) <= not (a or b);
    layer4_outputs(7241) <= a;
    layer4_outputs(7242) <= b and not a;
    layer4_outputs(7243) <= not (a xor b);
    layer4_outputs(7244) <= not (a xor b);
    layer4_outputs(7245) <= not b;
    layer4_outputs(7246) <= b;
    layer4_outputs(7247) <= b;
    layer4_outputs(7248) <= not (a or b);
    layer4_outputs(7249) <= not (a and b);
    layer4_outputs(7250) <= not a;
    layer4_outputs(7251) <= a;
    layer4_outputs(7252) <= not (a xor b);
    layer4_outputs(7253) <= not a;
    layer4_outputs(7254) <= not (a or b);
    layer4_outputs(7255) <= not a or b;
    layer4_outputs(7256) <= not a or b;
    layer4_outputs(7257) <= a and b;
    layer4_outputs(7258) <= b and not a;
    layer4_outputs(7259) <= not a or b;
    layer4_outputs(7260) <= a;
    layer4_outputs(7261) <= not (a or b);
    layer4_outputs(7262) <= a xor b;
    layer4_outputs(7263) <= a or b;
    layer4_outputs(7264) <= a;
    layer4_outputs(7265) <= b;
    layer4_outputs(7266) <= a or b;
    layer4_outputs(7267) <= not (a or b);
    layer4_outputs(7268) <= not b;
    layer4_outputs(7269) <= not b;
    layer4_outputs(7270) <= not a or b;
    layer4_outputs(7271) <= a and not b;
    layer4_outputs(7272) <= a;
    layer4_outputs(7273) <= not a;
    layer4_outputs(7274) <= a and not b;
    layer4_outputs(7275) <= a and not b;
    layer4_outputs(7276) <= not b or a;
    layer4_outputs(7277) <= not a;
    layer4_outputs(7278) <= b;
    layer4_outputs(7279) <= b;
    layer4_outputs(7280) <= '1';
    layer4_outputs(7281) <= not b or a;
    layer4_outputs(7282) <= a xor b;
    layer4_outputs(7283) <= not b or a;
    layer4_outputs(7284) <= '1';
    layer4_outputs(7285) <= not b;
    layer4_outputs(7286) <= a and not b;
    layer4_outputs(7287) <= not a;
    layer4_outputs(7288) <= a or b;
    layer4_outputs(7289) <= not (a xor b);
    layer4_outputs(7290) <= b and not a;
    layer4_outputs(7291) <= not a;
    layer4_outputs(7292) <= not (a and b);
    layer4_outputs(7293) <= a;
    layer4_outputs(7294) <= not (a xor b);
    layer4_outputs(7295) <= not b or a;
    layer4_outputs(7296) <= not (a xor b);
    layer4_outputs(7297) <= b and not a;
    layer4_outputs(7298) <= a xor b;
    layer4_outputs(7299) <= '1';
    layer4_outputs(7300) <= not a;
    layer4_outputs(7301) <= b and not a;
    layer4_outputs(7302) <= a;
    layer4_outputs(7303) <= not b;
    layer4_outputs(7304) <= a and not b;
    layer4_outputs(7305) <= a;
    layer4_outputs(7306) <= not (a and b);
    layer4_outputs(7307) <= a;
    layer4_outputs(7308) <= b and not a;
    layer4_outputs(7309) <= not (a or b);
    layer4_outputs(7310) <= not (a or b);
    layer4_outputs(7311) <= not (a or b);
    layer4_outputs(7312) <= a or b;
    layer4_outputs(7313) <= not b;
    layer4_outputs(7314) <= a;
    layer4_outputs(7315) <= not (a xor b);
    layer4_outputs(7316) <= a;
    layer4_outputs(7317) <= a;
    layer4_outputs(7318) <= a xor b;
    layer4_outputs(7319) <= not a or b;
    layer4_outputs(7320) <= a or b;
    layer4_outputs(7321) <= a;
    layer4_outputs(7322) <= b;
    layer4_outputs(7323) <= a and not b;
    layer4_outputs(7324) <= not a or b;
    layer4_outputs(7325) <= a and not b;
    layer4_outputs(7326) <= a xor b;
    layer4_outputs(7327) <= b;
    layer4_outputs(7328) <= not (a and b);
    layer4_outputs(7329) <= a and not b;
    layer4_outputs(7330) <= b;
    layer4_outputs(7331) <= a and b;
    layer4_outputs(7332) <= a and b;
    layer4_outputs(7333) <= a;
    layer4_outputs(7334) <= b;
    layer4_outputs(7335) <= a or b;
    layer4_outputs(7336) <= a;
    layer4_outputs(7337) <= b;
    layer4_outputs(7338) <= not (a or b);
    layer4_outputs(7339) <= a;
    layer4_outputs(7340) <= '0';
    layer4_outputs(7341) <= a and not b;
    layer4_outputs(7342) <= a and not b;
    layer4_outputs(7343) <= not a;
    layer4_outputs(7344) <= not (a xor b);
    layer4_outputs(7345) <= not (a or b);
    layer4_outputs(7346) <= not a or b;
    layer4_outputs(7347) <= not a or b;
    layer4_outputs(7348) <= not b;
    layer4_outputs(7349) <= not b or a;
    layer4_outputs(7350) <= a and b;
    layer4_outputs(7351) <= not b;
    layer4_outputs(7352) <= not b;
    layer4_outputs(7353) <= '1';
    layer4_outputs(7354) <= b;
    layer4_outputs(7355) <= not b;
    layer4_outputs(7356) <= not a;
    layer4_outputs(7357) <= not (a xor b);
    layer4_outputs(7358) <= not (a xor b);
    layer4_outputs(7359) <= b;
    layer4_outputs(7360) <= a and not b;
    layer4_outputs(7361) <= not a;
    layer4_outputs(7362) <= not (a or b);
    layer4_outputs(7363) <= a or b;
    layer4_outputs(7364) <= a;
    layer4_outputs(7365) <= not a or b;
    layer4_outputs(7366) <= a or b;
    layer4_outputs(7367) <= not (a xor b);
    layer4_outputs(7368) <= b;
    layer4_outputs(7369) <= not (a and b);
    layer4_outputs(7370) <= not a;
    layer4_outputs(7371) <= not a;
    layer4_outputs(7372) <= a and b;
    layer4_outputs(7373) <= a or b;
    layer4_outputs(7374) <= b;
    layer4_outputs(7375) <= a and b;
    layer4_outputs(7376) <= not b;
    layer4_outputs(7377) <= not b;
    layer4_outputs(7378) <= a xor b;
    layer4_outputs(7379) <= b;
    layer4_outputs(7380) <= not (a xor b);
    layer4_outputs(7381) <= a;
    layer4_outputs(7382) <= a and b;
    layer4_outputs(7383) <= not a;
    layer4_outputs(7384) <= a and not b;
    layer4_outputs(7385) <= not a;
    layer4_outputs(7386) <= b;
    layer4_outputs(7387) <= a and not b;
    layer4_outputs(7388) <= not a;
    layer4_outputs(7389) <= not (a and b);
    layer4_outputs(7390) <= a xor b;
    layer4_outputs(7391) <= not a;
    layer4_outputs(7392) <= not b;
    layer4_outputs(7393) <= a xor b;
    layer4_outputs(7394) <= a;
    layer4_outputs(7395) <= b;
    layer4_outputs(7396) <= a xor b;
    layer4_outputs(7397) <= not b;
    layer4_outputs(7398) <= a xor b;
    layer4_outputs(7399) <= not b;
    layer4_outputs(7400) <= not (a and b);
    layer4_outputs(7401) <= not (a or b);
    layer4_outputs(7402) <= not a or b;
    layer4_outputs(7403) <= a;
    layer4_outputs(7404) <= a and not b;
    layer4_outputs(7405) <= not (a xor b);
    layer4_outputs(7406) <= not (a xor b);
    layer4_outputs(7407) <= b and not a;
    layer4_outputs(7408) <= a or b;
    layer4_outputs(7409) <= not (a or b);
    layer4_outputs(7410) <= a;
    layer4_outputs(7411) <= b;
    layer4_outputs(7412) <= a and b;
    layer4_outputs(7413) <= b;
    layer4_outputs(7414) <= b;
    layer4_outputs(7415) <= not b or a;
    layer4_outputs(7416) <= b;
    layer4_outputs(7417) <= not (a or b);
    layer4_outputs(7418) <= a and b;
    layer4_outputs(7419) <= a;
    layer4_outputs(7420) <= a or b;
    layer4_outputs(7421) <= not a;
    layer4_outputs(7422) <= a or b;
    layer4_outputs(7423) <= not b;
    layer4_outputs(7424) <= not (a and b);
    layer4_outputs(7425) <= a and b;
    layer4_outputs(7426) <= not (a and b);
    layer4_outputs(7427) <= not b;
    layer4_outputs(7428) <= not b;
    layer4_outputs(7429) <= a and not b;
    layer4_outputs(7430) <= a;
    layer4_outputs(7431) <= not (a xor b);
    layer4_outputs(7432) <= a;
    layer4_outputs(7433) <= b and not a;
    layer4_outputs(7434) <= b;
    layer4_outputs(7435) <= a xor b;
    layer4_outputs(7436) <= b;
    layer4_outputs(7437) <= not b;
    layer4_outputs(7438) <= a xor b;
    layer4_outputs(7439) <= not a;
    layer4_outputs(7440) <= not b;
    layer4_outputs(7441) <= b;
    layer4_outputs(7442) <= not b;
    layer4_outputs(7443) <= '0';
    layer4_outputs(7444) <= a or b;
    layer4_outputs(7445) <= b;
    layer4_outputs(7446) <= not a or b;
    layer4_outputs(7447) <= not a or b;
    layer4_outputs(7448) <= not b;
    layer4_outputs(7449) <= a;
    layer4_outputs(7450) <= not b or a;
    layer4_outputs(7451) <= not b;
    layer4_outputs(7452) <= not a or b;
    layer4_outputs(7453) <= not (a and b);
    layer4_outputs(7454) <= '1';
    layer4_outputs(7455) <= not (a and b);
    layer4_outputs(7456) <= a;
    layer4_outputs(7457) <= not (a xor b);
    layer4_outputs(7458) <= a and b;
    layer4_outputs(7459) <= b and not a;
    layer4_outputs(7460) <= not a;
    layer4_outputs(7461) <= not (a or b);
    layer4_outputs(7462) <= not b or a;
    layer4_outputs(7463) <= not b;
    layer4_outputs(7464) <= b;
    layer4_outputs(7465) <= a or b;
    layer4_outputs(7466) <= not (a and b);
    layer4_outputs(7467) <= not b;
    layer4_outputs(7468) <= not a;
    layer4_outputs(7469) <= not a;
    layer4_outputs(7470) <= not a;
    layer4_outputs(7471) <= a and b;
    layer4_outputs(7472) <= not a;
    layer4_outputs(7473) <= not b or a;
    layer4_outputs(7474) <= not a or b;
    layer4_outputs(7475) <= b;
    layer4_outputs(7476) <= a or b;
    layer4_outputs(7477) <= a or b;
    layer4_outputs(7478) <= not b;
    layer4_outputs(7479) <= b and not a;
    layer4_outputs(7480) <= a;
    layer4_outputs(7481) <= not (a or b);
    layer4_outputs(7482) <= a and not b;
    layer4_outputs(7483) <= not (a or b);
    layer4_outputs(7484) <= not a;
    layer4_outputs(7485) <= not b;
    layer4_outputs(7486) <= b;
    layer4_outputs(7487) <= a;
    layer4_outputs(7488) <= a and b;
    layer4_outputs(7489) <= a;
    layer4_outputs(7490) <= a or b;
    layer4_outputs(7491) <= not (a or b);
    layer4_outputs(7492) <= a;
    layer4_outputs(7493) <= b and not a;
    layer4_outputs(7494) <= not (a or b);
    layer4_outputs(7495) <= not b;
    layer4_outputs(7496) <= not (a and b);
    layer4_outputs(7497) <= b and not a;
    layer4_outputs(7498) <= a xor b;
    layer4_outputs(7499) <= a and not b;
    layer4_outputs(7500) <= b;
    layer4_outputs(7501) <= b;
    layer4_outputs(7502) <= not a;
    layer4_outputs(7503) <= not a;
    layer4_outputs(7504) <= not b;
    layer4_outputs(7505) <= a and b;
    layer4_outputs(7506) <= b;
    layer4_outputs(7507) <= a;
    layer4_outputs(7508) <= b;
    layer4_outputs(7509) <= a;
    layer4_outputs(7510) <= not (a xor b);
    layer4_outputs(7511) <= a and not b;
    layer4_outputs(7512) <= not b;
    layer4_outputs(7513) <= a or b;
    layer4_outputs(7514) <= not b;
    layer4_outputs(7515) <= b;
    layer4_outputs(7516) <= a and b;
    layer4_outputs(7517) <= a and b;
    layer4_outputs(7518) <= b;
    layer4_outputs(7519) <= '1';
    layer4_outputs(7520) <= b;
    layer4_outputs(7521) <= b;
    layer4_outputs(7522) <= a;
    layer4_outputs(7523) <= not a;
    layer4_outputs(7524) <= not b or a;
    layer4_outputs(7525) <= not a or b;
    layer4_outputs(7526) <= b;
    layer4_outputs(7527) <= b;
    layer4_outputs(7528) <= not (a xor b);
    layer4_outputs(7529) <= '0';
    layer4_outputs(7530) <= a and not b;
    layer4_outputs(7531) <= not a;
    layer4_outputs(7532) <= a or b;
    layer4_outputs(7533) <= not b or a;
    layer4_outputs(7534) <= a and not b;
    layer4_outputs(7535) <= a and not b;
    layer4_outputs(7536) <= not a;
    layer4_outputs(7537) <= not b or a;
    layer4_outputs(7538) <= a;
    layer4_outputs(7539) <= not (a xor b);
    layer4_outputs(7540) <= b;
    layer4_outputs(7541) <= a or b;
    layer4_outputs(7542) <= a xor b;
    layer4_outputs(7543) <= a;
    layer4_outputs(7544) <= not (a or b);
    layer4_outputs(7545) <= not a;
    layer4_outputs(7546) <= not a;
    layer4_outputs(7547) <= not (a or b);
    layer4_outputs(7548) <= b;
    layer4_outputs(7549) <= a xor b;
    layer4_outputs(7550) <= not b;
    layer4_outputs(7551) <= not (a or b);
    layer4_outputs(7552) <= not b;
    layer4_outputs(7553) <= not (a or b);
    layer4_outputs(7554) <= not a;
    layer4_outputs(7555) <= '0';
    layer4_outputs(7556) <= a;
    layer4_outputs(7557) <= a xor b;
    layer4_outputs(7558) <= '0';
    layer4_outputs(7559) <= b;
    layer4_outputs(7560) <= b;
    layer4_outputs(7561) <= a and b;
    layer4_outputs(7562) <= a and not b;
    layer4_outputs(7563) <= not b;
    layer4_outputs(7564) <= b;
    layer4_outputs(7565) <= a and not b;
    layer4_outputs(7566) <= a and not b;
    layer4_outputs(7567) <= not (a or b);
    layer4_outputs(7568) <= not a;
    layer4_outputs(7569) <= not (a and b);
    layer4_outputs(7570) <= not b;
    layer4_outputs(7571) <= not b;
    layer4_outputs(7572) <= a xor b;
    layer4_outputs(7573) <= not b or a;
    layer4_outputs(7574) <= not a;
    layer4_outputs(7575) <= a or b;
    layer4_outputs(7576) <= not b;
    layer4_outputs(7577) <= b;
    layer4_outputs(7578) <= b;
    layer4_outputs(7579) <= not (a or b);
    layer4_outputs(7580) <= a;
    layer4_outputs(7581) <= not b or a;
    layer4_outputs(7582) <= not (a or b);
    layer4_outputs(7583) <= not a;
    layer4_outputs(7584) <= b;
    layer4_outputs(7585) <= b;
    layer4_outputs(7586) <= not (a xor b);
    layer4_outputs(7587) <= a and not b;
    layer4_outputs(7588) <= a;
    layer4_outputs(7589) <= b;
    layer4_outputs(7590) <= not b or a;
    layer4_outputs(7591) <= not (a xor b);
    layer4_outputs(7592) <= '1';
    layer4_outputs(7593) <= a;
    layer4_outputs(7594) <= not b or a;
    layer4_outputs(7595) <= a;
    layer4_outputs(7596) <= not a;
    layer4_outputs(7597) <= a;
    layer4_outputs(7598) <= b;
    layer4_outputs(7599) <= a and b;
    layer4_outputs(7600) <= a;
    layer4_outputs(7601) <= a and b;
    layer4_outputs(7602) <= b and not a;
    layer4_outputs(7603) <= not b or a;
    layer4_outputs(7604) <= a;
    layer4_outputs(7605) <= not (a or b);
    layer4_outputs(7606) <= not a;
    layer4_outputs(7607) <= b;
    layer4_outputs(7608) <= not b;
    layer4_outputs(7609) <= not a;
    layer4_outputs(7610) <= a;
    layer4_outputs(7611) <= not a;
    layer4_outputs(7612) <= not b or a;
    layer4_outputs(7613) <= a and not b;
    layer4_outputs(7614) <= not b;
    layer4_outputs(7615) <= b;
    layer4_outputs(7616) <= a;
    layer4_outputs(7617) <= not (a xor b);
    layer4_outputs(7618) <= not a;
    layer4_outputs(7619) <= not a;
    layer4_outputs(7620) <= not (a or b);
    layer4_outputs(7621) <= '0';
    layer4_outputs(7622) <= a and b;
    layer4_outputs(7623) <= not a;
    layer4_outputs(7624) <= '0';
    layer4_outputs(7625) <= b;
    layer4_outputs(7626) <= not a or b;
    layer4_outputs(7627) <= not a or b;
    layer4_outputs(7628) <= a and b;
    layer4_outputs(7629) <= b;
    layer4_outputs(7630) <= not b;
    layer4_outputs(7631) <= a xor b;
    layer4_outputs(7632) <= not a;
    layer4_outputs(7633) <= a xor b;
    layer4_outputs(7634) <= '0';
    layer4_outputs(7635) <= a;
    layer4_outputs(7636) <= a and b;
    layer4_outputs(7637) <= b;
    layer4_outputs(7638) <= b;
    layer4_outputs(7639) <= not a or b;
    layer4_outputs(7640) <= not a or b;
    layer4_outputs(7641) <= not a or b;
    layer4_outputs(7642) <= a;
    layer4_outputs(7643) <= b;
    layer4_outputs(7644) <= a;
    layer4_outputs(7645) <= b;
    layer4_outputs(7646) <= b;
    layer4_outputs(7647) <= a or b;
    layer4_outputs(7648) <= not a;
    layer4_outputs(7649) <= a;
    layer4_outputs(7650) <= a or b;
    layer4_outputs(7651) <= a and b;
    layer4_outputs(7652) <= a and not b;
    layer4_outputs(7653) <= b;
    layer4_outputs(7654) <= b;
    layer4_outputs(7655) <= not a;
    layer4_outputs(7656) <= not a;
    layer4_outputs(7657) <= not (a xor b);
    layer4_outputs(7658) <= not a;
    layer4_outputs(7659) <= not a;
    layer4_outputs(7660) <= not b or a;
    layer4_outputs(7661) <= not b;
    layer4_outputs(7662) <= a;
    layer4_outputs(7663) <= not b;
    layer4_outputs(7664) <= b and not a;
    layer4_outputs(7665) <= not b;
    layer4_outputs(7666) <= not b;
    layer4_outputs(7667) <= not (a or b);
    layer4_outputs(7668) <= a and not b;
    layer4_outputs(7669) <= a and b;
    layer4_outputs(7670) <= '0';
    layer4_outputs(7671) <= a or b;
    layer4_outputs(7672) <= not b;
    layer4_outputs(7673) <= a;
    layer4_outputs(7674) <= not b or a;
    layer4_outputs(7675) <= a or b;
    layer4_outputs(7676) <= not (a xor b);
    layer4_outputs(7677) <= a and not b;
    layer4_outputs(7678) <= not (a or b);
    layer4_outputs(7679) <= a;
    layer4_outputs(7680) <= not (a or b);
    layer4_outputs(7681) <= not a or b;
    layer4_outputs(7682) <= a and b;
    layer4_outputs(7683) <= a or b;
    layer4_outputs(7684) <= not (a or b);
    layer4_outputs(7685) <= a xor b;
    layer4_outputs(7686) <= not a or b;
    layer4_outputs(7687) <= a and not b;
    layer4_outputs(7688) <= not a;
    layer4_outputs(7689) <= not b;
    layer4_outputs(7690) <= not (a and b);
    layer4_outputs(7691) <= a;
    layer4_outputs(7692) <= b;
    layer4_outputs(7693) <= a or b;
    layer4_outputs(7694) <= a xor b;
    layer4_outputs(7695) <= '1';
    layer4_outputs(7696) <= not b or a;
    layer4_outputs(7697) <= b and not a;
    layer4_outputs(7698) <= '0';
    layer4_outputs(7699) <= not b;
    layer4_outputs(7700) <= not b or a;
    layer4_outputs(7701) <= not a;
    layer4_outputs(7702) <= b and not a;
    layer4_outputs(7703) <= not a;
    layer4_outputs(7704) <= a or b;
    layer4_outputs(7705) <= a;
    layer4_outputs(7706) <= not b or a;
    layer4_outputs(7707) <= a and not b;
    layer4_outputs(7708) <= a;
    layer4_outputs(7709) <= not a;
    layer4_outputs(7710) <= b and not a;
    layer4_outputs(7711) <= '1';
    layer4_outputs(7712) <= a xor b;
    layer4_outputs(7713) <= b;
    layer4_outputs(7714) <= a and not b;
    layer4_outputs(7715) <= not a;
    layer4_outputs(7716) <= not a;
    layer4_outputs(7717) <= not (a xor b);
    layer4_outputs(7718) <= b;
    layer4_outputs(7719) <= not b;
    layer4_outputs(7720) <= not (a and b);
    layer4_outputs(7721) <= not a;
    layer4_outputs(7722) <= a and b;
    layer4_outputs(7723) <= not a;
    layer4_outputs(7724) <= b;
    layer4_outputs(7725) <= '1';
    layer4_outputs(7726) <= not (a xor b);
    layer4_outputs(7727) <= '0';
    layer4_outputs(7728) <= a xor b;
    layer4_outputs(7729) <= b;
    layer4_outputs(7730) <= not b;
    layer4_outputs(7731) <= b;
    layer4_outputs(7732) <= a and not b;
    layer4_outputs(7733) <= not (a xor b);
    layer4_outputs(7734) <= '0';
    layer4_outputs(7735) <= b;
    layer4_outputs(7736) <= a and not b;
    layer4_outputs(7737) <= a and not b;
    layer4_outputs(7738) <= a or b;
    layer4_outputs(7739) <= not a;
    layer4_outputs(7740) <= not (a and b);
    layer4_outputs(7741) <= a and b;
    layer4_outputs(7742) <= a and not b;
    layer4_outputs(7743) <= not a;
    layer4_outputs(7744) <= b and not a;
    layer4_outputs(7745) <= not a;
    layer4_outputs(7746) <= not b;
    layer4_outputs(7747) <= not b;
    layer4_outputs(7748) <= not a;
    layer4_outputs(7749) <= '1';
    layer4_outputs(7750) <= '1';
    layer4_outputs(7751) <= a and not b;
    layer4_outputs(7752) <= '0';
    layer4_outputs(7753) <= not (a and b);
    layer4_outputs(7754) <= a;
    layer4_outputs(7755) <= a or b;
    layer4_outputs(7756) <= a and not b;
    layer4_outputs(7757) <= a;
    layer4_outputs(7758) <= a;
    layer4_outputs(7759) <= not b or a;
    layer4_outputs(7760) <= not (a and b);
    layer4_outputs(7761) <= a or b;
    layer4_outputs(7762) <= b;
    layer4_outputs(7763) <= '1';
    layer4_outputs(7764) <= a and b;
    layer4_outputs(7765) <= a and not b;
    layer4_outputs(7766) <= a and not b;
    layer4_outputs(7767) <= not b;
    layer4_outputs(7768) <= not b or a;
    layer4_outputs(7769) <= b;
    layer4_outputs(7770) <= not (a xor b);
    layer4_outputs(7771) <= not b;
    layer4_outputs(7772) <= b;
    layer4_outputs(7773) <= a;
    layer4_outputs(7774) <= a;
    layer4_outputs(7775) <= not a;
    layer4_outputs(7776) <= not a;
    layer4_outputs(7777) <= b;
    layer4_outputs(7778) <= a and b;
    layer4_outputs(7779) <= b;
    layer4_outputs(7780) <= not b;
    layer4_outputs(7781) <= a;
    layer4_outputs(7782) <= not (a and b);
    layer4_outputs(7783) <= '0';
    layer4_outputs(7784) <= not b;
    layer4_outputs(7785) <= a and b;
    layer4_outputs(7786) <= not b;
    layer4_outputs(7787) <= not a;
    layer4_outputs(7788) <= not (a xor b);
    layer4_outputs(7789) <= b;
    layer4_outputs(7790) <= a and not b;
    layer4_outputs(7791) <= b and not a;
    layer4_outputs(7792) <= not a;
    layer4_outputs(7793) <= b and not a;
    layer4_outputs(7794) <= a xor b;
    layer4_outputs(7795) <= a and not b;
    layer4_outputs(7796) <= a;
    layer4_outputs(7797) <= a or b;
    layer4_outputs(7798) <= a or b;
    layer4_outputs(7799) <= not b or a;
    layer4_outputs(7800) <= b;
    layer4_outputs(7801) <= a;
    layer4_outputs(7802) <= not b;
    layer4_outputs(7803) <= b;
    layer4_outputs(7804) <= not a;
    layer4_outputs(7805) <= a xor b;
    layer4_outputs(7806) <= b and not a;
    layer4_outputs(7807) <= a xor b;
    layer4_outputs(7808) <= b and not a;
    layer4_outputs(7809) <= not b;
    layer4_outputs(7810) <= a or b;
    layer4_outputs(7811) <= '1';
    layer4_outputs(7812) <= a xor b;
    layer4_outputs(7813) <= not a or b;
    layer4_outputs(7814) <= not (a and b);
    layer4_outputs(7815) <= not b;
    layer4_outputs(7816) <= a;
    layer4_outputs(7817) <= b;
    layer4_outputs(7818) <= not (a or b);
    layer4_outputs(7819) <= not b or a;
    layer4_outputs(7820) <= not a;
    layer4_outputs(7821) <= b;
    layer4_outputs(7822) <= not b;
    layer4_outputs(7823) <= a;
    layer4_outputs(7824) <= b;
    layer4_outputs(7825) <= a and not b;
    layer4_outputs(7826) <= not b;
    layer4_outputs(7827) <= not a or b;
    layer4_outputs(7828) <= b;
    layer4_outputs(7829) <= '1';
    layer4_outputs(7830) <= a and b;
    layer4_outputs(7831) <= a;
    layer4_outputs(7832) <= not b;
    layer4_outputs(7833) <= a;
    layer4_outputs(7834) <= not b or a;
    layer4_outputs(7835) <= '0';
    layer4_outputs(7836) <= not b;
    layer4_outputs(7837) <= not a;
    layer4_outputs(7838) <= not b or a;
    layer4_outputs(7839) <= not (a or b);
    layer4_outputs(7840) <= not b or a;
    layer4_outputs(7841) <= not b;
    layer4_outputs(7842) <= a and b;
    layer4_outputs(7843) <= not a;
    layer4_outputs(7844) <= not (a xor b);
    layer4_outputs(7845) <= a or b;
    layer4_outputs(7846) <= a;
    layer4_outputs(7847) <= not a or b;
    layer4_outputs(7848) <= not b or a;
    layer4_outputs(7849) <= not b;
    layer4_outputs(7850) <= not a;
    layer4_outputs(7851) <= not (a xor b);
    layer4_outputs(7852) <= not b;
    layer4_outputs(7853) <= not (a and b);
    layer4_outputs(7854) <= a xor b;
    layer4_outputs(7855) <= b;
    layer4_outputs(7856) <= not (a and b);
    layer4_outputs(7857) <= not a;
    layer4_outputs(7858) <= a;
    layer4_outputs(7859) <= '0';
    layer4_outputs(7860) <= not a;
    layer4_outputs(7861) <= a and b;
    layer4_outputs(7862) <= not (a xor b);
    layer4_outputs(7863) <= a;
    layer4_outputs(7864) <= not b;
    layer4_outputs(7865) <= not (a and b);
    layer4_outputs(7866) <= not a;
    layer4_outputs(7867) <= not a;
    layer4_outputs(7868) <= not a;
    layer4_outputs(7869) <= b;
    layer4_outputs(7870) <= not (a or b);
    layer4_outputs(7871) <= a and b;
    layer4_outputs(7872) <= a;
    layer4_outputs(7873) <= not a or b;
    layer4_outputs(7874) <= not (a xor b);
    layer4_outputs(7875) <= b;
    layer4_outputs(7876) <= a xor b;
    layer4_outputs(7877) <= not a;
    layer4_outputs(7878) <= b;
    layer4_outputs(7879) <= not b or a;
    layer4_outputs(7880) <= not a;
    layer4_outputs(7881) <= not (a or b);
    layer4_outputs(7882) <= not a;
    layer4_outputs(7883) <= not (a and b);
    layer4_outputs(7884) <= not b or a;
    layer4_outputs(7885) <= not a;
    layer4_outputs(7886) <= b;
    layer4_outputs(7887) <= a and not b;
    layer4_outputs(7888) <= not (a xor b);
    layer4_outputs(7889) <= a and not b;
    layer4_outputs(7890) <= b and not a;
    layer4_outputs(7891) <= not b or a;
    layer4_outputs(7892) <= a xor b;
    layer4_outputs(7893) <= not b;
    layer4_outputs(7894) <= a and b;
    layer4_outputs(7895) <= a and not b;
    layer4_outputs(7896) <= b;
    layer4_outputs(7897) <= not a or b;
    layer4_outputs(7898) <= not (a or b);
    layer4_outputs(7899) <= not (a and b);
    layer4_outputs(7900) <= a or b;
    layer4_outputs(7901) <= b and not a;
    layer4_outputs(7902) <= not (a or b);
    layer4_outputs(7903) <= b;
    layer4_outputs(7904) <= not b or a;
    layer4_outputs(7905) <= not (a or b);
    layer4_outputs(7906) <= not b;
    layer4_outputs(7907) <= not b;
    layer4_outputs(7908) <= b;
    layer4_outputs(7909) <= not (a or b);
    layer4_outputs(7910) <= not a or b;
    layer4_outputs(7911) <= a and b;
    layer4_outputs(7912) <= b;
    layer4_outputs(7913) <= a or b;
    layer4_outputs(7914) <= b and not a;
    layer4_outputs(7915) <= b;
    layer4_outputs(7916) <= a;
    layer4_outputs(7917) <= not b or a;
    layer4_outputs(7918) <= a or b;
    layer4_outputs(7919) <= a or b;
    layer4_outputs(7920) <= a and b;
    layer4_outputs(7921) <= '1';
    layer4_outputs(7922) <= not b;
    layer4_outputs(7923) <= '1';
    layer4_outputs(7924) <= not (a and b);
    layer4_outputs(7925) <= not (a or b);
    layer4_outputs(7926) <= a;
    layer4_outputs(7927) <= a or b;
    layer4_outputs(7928) <= b;
    layer4_outputs(7929) <= not a or b;
    layer4_outputs(7930) <= a xor b;
    layer4_outputs(7931) <= a or b;
    layer4_outputs(7932) <= a xor b;
    layer4_outputs(7933) <= not a;
    layer4_outputs(7934) <= b and not a;
    layer4_outputs(7935) <= '1';
    layer4_outputs(7936) <= a;
    layer4_outputs(7937) <= not a;
    layer4_outputs(7938) <= not (a or b);
    layer4_outputs(7939) <= not b or a;
    layer4_outputs(7940) <= a xor b;
    layer4_outputs(7941) <= '0';
    layer4_outputs(7942) <= b;
    layer4_outputs(7943) <= b;
    layer4_outputs(7944) <= not b;
    layer4_outputs(7945) <= a and not b;
    layer4_outputs(7946) <= not a;
    layer4_outputs(7947) <= a;
    layer4_outputs(7948) <= a;
    layer4_outputs(7949) <= a and b;
    layer4_outputs(7950) <= a and b;
    layer4_outputs(7951) <= a xor b;
    layer4_outputs(7952) <= a and b;
    layer4_outputs(7953) <= '0';
    layer4_outputs(7954) <= a and not b;
    layer4_outputs(7955) <= a;
    layer4_outputs(7956) <= b and not a;
    layer4_outputs(7957) <= a or b;
    layer4_outputs(7958) <= a and not b;
    layer4_outputs(7959) <= a xor b;
    layer4_outputs(7960) <= b and not a;
    layer4_outputs(7961) <= a and not b;
    layer4_outputs(7962) <= not a;
    layer4_outputs(7963) <= not (a xor b);
    layer4_outputs(7964) <= not b;
    layer4_outputs(7965) <= not a;
    layer4_outputs(7966) <= b;
    layer4_outputs(7967) <= not b;
    layer4_outputs(7968) <= a or b;
    layer4_outputs(7969) <= not b;
    layer4_outputs(7970) <= not a;
    layer4_outputs(7971) <= not b or a;
    layer4_outputs(7972) <= not a;
    layer4_outputs(7973) <= not (a xor b);
    layer4_outputs(7974) <= not a or b;
    layer4_outputs(7975) <= b;
    layer4_outputs(7976) <= not b or a;
    layer4_outputs(7977) <= '0';
    layer4_outputs(7978) <= a;
    layer4_outputs(7979) <= not a or b;
    layer4_outputs(7980) <= not a;
    layer4_outputs(7981) <= b and not a;
    layer4_outputs(7982) <= a or b;
    layer4_outputs(7983) <= not b;
    layer4_outputs(7984) <= not (a xor b);
    layer4_outputs(7985) <= b and not a;
    layer4_outputs(7986) <= not (a or b);
    layer4_outputs(7987) <= not (a and b);
    layer4_outputs(7988) <= b;
    layer4_outputs(7989) <= a and not b;
    layer4_outputs(7990) <= a xor b;
    layer4_outputs(7991) <= not b;
    layer4_outputs(7992) <= not b;
    layer4_outputs(7993) <= b;
    layer4_outputs(7994) <= not b or a;
    layer4_outputs(7995) <= a or b;
    layer4_outputs(7996) <= not (a and b);
    layer4_outputs(7997) <= b and not a;
    layer4_outputs(7998) <= not b;
    layer4_outputs(7999) <= not b or a;
    layer4_outputs(8000) <= b;
    layer4_outputs(8001) <= a xor b;
    layer4_outputs(8002) <= not b;
    layer4_outputs(8003) <= b and not a;
    layer4_outputs(8004) <= '0';
    layer4_outputs(8005) <= a or b;
    layer4_outputs(8006) <= b and not a;
    layer4_outputs(8007) <= not (a or b);
    layer4_outputs(8008) <= not b;
    layer4_outputs(8009) <= not b;
    layer4_outputs(8010) <= a and not b;
    layer4_outputs(8011) <= not b;
    layer4_outputs(8012) <= not a;
    layer4_outputs(8013) <= a and not b;
    layer4_outputs(8014) <= not a;
    layer4_outputs(8015) <= not a or b;
    layer4_outputs(8016) <= not (a and b);
    layer4_outputs(8017) <= b;
    layer4_outputs(8018) <= not b or a;
    layer4_outputs(8019) <= not a or b;
    layer4_outputs(8020) <= not (a or b);
    layer4_outputs(8021) <= not b;
    layer4_outputs(8022) <= not (a or b);
    layer4_outputs(8023) <= not (a xor b);
    layer4_outputs(8024) <= a;
    layer4_outputs(8025) <= b;
    layer4_outputs(8026) <= a xor b;
    layer4_outputs(8027) <= not b;
    layer4_outputs(8028) <= a xor b;
    layer4_outputs(8029) <= not (a and b);
    layer4_outputs(8030) <= b;
    layer4_outputs(8031) <= '1';
    layer4_outputs(8032) <= not b or a;
    layer4_outputs(8033) <= not b;
    layer4_outputs(8034) <= a;
    layer4_outputs(8035) <= '1';
    layer4_outputs(8036) <= b;
    layer4_outputs(8037) <= a or b;
    layer4_outputs(8038) <= not b or a;
    layer4_outputs(8039) <= not a or b;
    layer4_outputs(8040) <= not (a or b);
    layer4_outputs(8041) <= a and b;
    layer4_outputs(8042) <= not a;
    layer4_outputs(8043) <= '0';
    layer4_outputs(8044) <= not b;
    layer4_outputs(8045) <= not a or b;
    layer4_outputs(8046) <= not a;
    layer4_outputs(8047) <= a or b;
    layer4_outputs(8048) <= '1';
    layer4_outputs(8049) <= not (a and b);
    layer4_outputs(8050) <= a xor b;
    layer4_outputs(8051) <= not b;
    layer4_outputs(8052) <= a and not b;
    layer4_outputs(8053) <= a;
    layer4_outputs(8054) <= not (a or b);
    layer4_outputs(8055) <= a and b;
    layer4_outputs(8056) <= a xor b;
    layer4_outputs(8057) <= a;
    layer4_outputs(8058) <= a and b;
    layer4_outputs(8059) <= b;
    layer4_outputs(8060) <= b;
    layer4_outputs(8061) <= not b;
    layer4_outputs(8062) <= not b or a;
    layer4_outputs(8063) <= not a or b;
    layer4_outputs(8064) <= not b or a;
    layer4_outputs(8065) <= b and not a;
    layer4_outputs(8066) <= not (a and b);
    layer4_outputs(8067) <= not (a or b);
    layer4_outputs(8068) <= not a;
    layer4_outputs(8069) <= not (a or b);
    layer4_outputs(8070) <= not (a or b);
    layer4_outputs(8071) <= a;
    layer4_outputs(8072) <= not a;
    layer4_outputs(8073) <= not a or b;
    layer4_outputs(8074) <= not b or a;
    layer4_outputs(8075) <= '0';
    layer4_outputs(8076) <= a;
    layer4_outputs(8077) <= a or b;
    layer4_outputs(8078) <= not a;
    layer4_outputs(8079) <= b;
    layer4_outputs(8080) <= a;
    layer4_outputs(8081) <= not b or a;
    layer4_outputs(8082) <= not b;
    layer4_outputs(8083) <= b;
    layer4_outputs(8084) <= a xor b;
    layer4_outputs(8085) <= b;
    layer4_outputs(8086) <= not b;
    layer4_outputs(8087) <= not b or a;
    layer4_outputs(8088) <= not a or b;
    layer4_outputs(8089) <= a and b;
    layer4_outputs(8090) <= b and not a;
    layer4_outputs(8091) <= not a;
    layer4_outputs(8092) <= not (a and b);
    layer4_outputs(8093) <= not (a and b);
    layer4_outputs(8094) <= a;
    layer4_outputs(8095) <= not (a or b);
    layer4_outputs(8096) <= not b;
    layer4_outputs(8097) <= a;
    layer4_outputs(8098) <= not a;
    layer4_outputs(8099) <= not a;
    layer4_outputs(8100) <= not b;
    layer4_outputs(8101) <= not (a xor b);
    layer4_outputs(8102) <= b;
    layer4_outputs(8103) <= a xor b;
    layer4_outputs(8104) <= not b;
    layer4_outputs(8105) <= not (a xor b);
    layer4_outputs(8106) <= '0';
    layer4_outputs(8107) <= a;
    layer4_outputs(8108) <= b;
    layer4_outputs(8109) <= '0';
    layer4_outputs(8110) <= '1';
    layer4_outputs(8111) <= a and b;
    layer4_outputs(8112) <= not (a or b);
    layer4_outputs(8113) <= not b or a;
    layer4_outputs(8114) <= a and b;
    layer4_outputs(8115) <= not a;
    layer4_outputs(8116) <= a xor b;
    layer4_outputs(8117) <= not (a and b);
    layer4_outputs(8118) <= not b;
    layer4_outputs(8119) <= not a;
    layer4_outputs(8120) <= not (a and b);
    layer4_outputs(8121) <= not (a or b);
    layer4_outputs(8122) <= not b or a;
    layer4_outputs(8123) <= not a or b;
    layer4_outputs(8124) <= not (a xor b);
    layer4_outputs(8125) <= b;
    layer4_outputs(8126) <= a;
    layer4_outputs(8127) <= not (a and b);
    layer4_outputs(8128) <= not a or b;
    layer4_outputs(8129) <= b;
    layer4_outputs(8130) <= not a or b;
    layer4_outputs(8131) <= a or b;
    layer4_outputs(8132) <= a;
    layer4_outputs(8133) <= a or b;
    layer4_outputs(8134) <= a;
    layer4_outputs(8135) <= b and not a;
    layer4_outputs(8136) <= not a;
    layer4_outputs(8137) <= not a;
    layer4_outputs(8138) <= a and b;
    layer4_outputs(8139) <= not a or b;
    layer4_outputs(8140) <= a and not b;
    layer4_outputs(8141) <= b and not a;
    layer4_outputs(8142) <= b;
    layer4_outputs(8143) <= not b or a;
    layer4_outputs(8144) <= not (a and b);
    layer4_outputs(8145) <= not (a or b);
    layer4_outputs(8146) <= not (a or b);
    layer4_outputs(8147) <= a or b;
    layer4_outputs(8148) <= not b or a;
    layer4_outputs(8149) <= a and b;
    layer4_outputs(8150) <= b;
    layer4_outputs(8151) <= a or b;
    layer4_outputs(8152) <= b and not a;
    layer4_outputs(8153) <= a and not b;
    layer4_outputs(8154) <= b;
    layer4_outputs(8155) <= not (a xor b);
    layer4_outputs(8156) <= not a or b;
    layer4_outputs(8157) <= not a;
    layer4_outputs(8158) <= not b;
    layer4_outputs(8159) <= not a;
    layer4_outputs(8160) <= b;
    layer4_outputs(8161) <= a;
    layer4_outputs(8162) <= b;
    layer4_outputs(8163) <= a and b;
    layer4_outputs(8164) <= a or b;
    layer4_outputs(8165) <= not a;
    layer4_outputs(8166) <= a;
    layer4_outputs(8167) <= a or b;
    layer4_outputs(8168) <= a or b;
    layer4_outputs(8169) <= not a;
    layer4_outputs(8170) <= not (a or b);
    layer4_outputs(8171) <= not (a xor b);
    layer4_outputs(8172) <= b;
    layer4_outputs(8173) <= not a or b;
    layer4_outputs(8174) <= not (a xor b);
    layer4_outputs(8175) <= not b;
    layer4_outputs(8176) <= '1';
    layer4_outputs(8177) <= a;
    layer4_outputs(8178) <= b;
    layer4_outputs(8179) <= b;
    layer4_outputs(8180) <= b and not a;
    layer4_outputs(8181) <= b;
    layer4_outputs(8182) <= a and b;
    layer4_outputs(8183) <= a and not b;
    layer4_outputs(8184) <= a and b;
    layer4_outputs(8185) <= b and not a;
    layer4_outputs(8186) <= not b or a;
    layer4_outputs(8187) <= b and not a;
    layer4_outputs(8188) <= not b;
    layer4_outputs(8189) <= b;
    layer4_outputs(8190) <= not b;
    layer4_outputs(8191) <= a or b;
    layer4_outputs(8192) <= not b;
    layer4_outputs(8193) <= not a or b;
    layer4_outputs(8194) <= not a;
    layer4_outputs(8195) <= a and not b;
    layer4_outputs(8196) <= not a or b;
    layer4_outputs(8197) <= not (a xor b);
    layer4_outputs(8198) <= not a;
    layer4_outputs(8199) <= not (a xor b);
    layer4_outputs(8200) <= a xor b;
    layer4_outputs(8201) <= a;
    layer4_outputs(8202) <= a;
    layer4_outputs(8203) <= not a;
    layer4_outputs(8204) <= not b;
    layer4_outputs(8205) <= not b;
    layer4_outputs(8206) <= not b or a;
    layer4_outputs(8207) <= '1';
    layer4_outputs(8208) <= not b or a;
    layer4_outputs(8209) <= a or b;
    layer4_outputs(8210) <= a;
    layer4_outputs(8211) <= b;
    layer4_outputs(8212) <= a and b;
    layer4_outputs(8213) <= not b or a;
    layer4_outputs(8214) <= not b;
    layer4_outputs(8215) <= not b;
    layer4_outputs(8216) <= a and b;
    layer4_outputs(8217) <= not b;
    layer4_outputs(8218) <= a or b;
    layer4_outputs(8219) <= not a;
    layer4_outputs(8220) <= not b or a;
    layer4_outputs(8221) <= not b;
    layer4_outputs(8222) <= not a;
    layer4_outputs(8223) <= '1';
    layer4_outputs(8224) <= a and not b;
    layer4_outputs(8225) <= not a or b;
    layer4_outputs(8226) <= not a or b;
    layer4_outputs(8227) <= not (a and b);
    layer4_outputs(8228) <= a and not b;
    layer4_outputs(8229) <= not (a or b);
    layer4_outputs(8230) <= not b;
    layer4_outputs(8231) <= a or b;
    layer4_outputs(8232) <= a and not b;
    layer4_outputs(8233) <= b;
    layer4_outputs(8234) <= not b;
    layer4_outputs(8235) <= not a;
    layer4_outputs(8236) <= a;
    layer4_outputs(8237) <= a xor b;
    layer4_outputs(8238) <= a xor b;
    layer4_outputs(8239) <= a;
    layer4_outputs(8240) <= a;
    layer4_outputs(8241) <= not a or b;
    layer4_outputs(8242) <= not b;
    layer4_outputs(8243) <= b;
    layer4_outputs(8244) <= not b;
    layer4_outputs(8245) <= b;
    layer4_outputs(8246) <= not b;
    layer4_outputs(8247) <= a and b;
    layer4_outputs(8248) <= a xor b;
    layer4_outputs(8249) <= '0';
    layer4_outputs(8250) <= not b;
    layer4_outputs(8251) <= not (a or b);
    layer4_outputs(8252) <= not a;
    layer4_outputs(8253) <= not (a and b);
    layer4_outputs(8254) <= b and not a;
    layer4_outputs(8255) <= a and b;
    layer4_outputs(8256) <= a;
    layer4_outputs(8257) <= not (a or b);
    layer4_outputs(8258) <= b;
    layer4_outputs(8259) <= a and b;
    layer4_outputs(8260) <= a xor b;
    layer4_outputs(8261) <= a and b;
    layer4_outputs(8262) <= not b;
    layer4_outputs(8263) <= b;
    layer4_outputs(8264) <= a and b;
    layer4_outputs(8265) <= a or b;
    layer4_outputs(8266) <= not a or b;
    layer4_outputs(8267) <= a and b;
    layer4_outputs(8268) <= a and b;
    layer4_outputs(8269) <= not b;
    layer4_outputs(8270) <= not a or b;
    layer4_outputs(8271) <= a and b;
    layer4_outputs(8272) <= b;
    layer4_outputs(8273) <= not b;
    layer4_outputs(8274) <= b and not a;
    layer4_outputs(8275) <= a and not b;
    layer4_outputs(8276) <= not a or b;
    layer4_outputs(8277) <= a xor b;
    layer4_outputs(8278) <= b;
    layer4_outputs(8279) <= not a;
    layer4_outputs(8280) <= not b or a;
    layer4_outputs(8281) <= '0';
    layer4_outputs(8282) <= not a or b;
    layer4_outputs(8283) <= b;
    layer4_outputs(8284) <= not (a xor b);
    layer4_outputs(8285) <= not b;
    layer4_outputs(8286) <= a and b;
    layer4_outputs(8287) <= not a;
    layer4_outputs(8288) <= a;
    layer4_outputs(8289) <= not b;
    layer4_outputs(8290) <= a;
    layer4_outputs(8291) <= not (a or b);
    layer4_outputs(8292) <= not b;
    layer4_outputs(8293) <= '0';
    layer4_outputs(8294) <= a and b;
    layer4_outputs(8295) <= not a;
    layer4_outputs(8296) <= not b;
    layer4_outputs(8297) <= b and not a;
    layer4_outputs(8298) <= not a or b;
    layer4_outputs(8299) <= not b or a;
    layer4_outputs(8300) <= not b or a;
    layer4_outputs(8301) <= not b;
    layer4_outputs(8302) <= not (a and b);
    layer4_outputs(8303) <= not b;
    layer4_outputs(8304) <= a or b;
    layer4_outputs(8305) <= not b;
    layer4_outputs(8306) <= not a;
    layer4_outputs(8307) <= a xor b;
    layer4_outputs(8308) <= not b;
    layer4_outputs(8309) <= not a;
    layer4_outputs(8310) <= '0';
    layer4_outputs(8311) <= a and b;
    layer4_outputs(8312) <= a and not b;
    layer4_outputs(8313) <= not (a and b);
    layer4_outputs(8314) <= not a;
    layer4_outputs(8315) <= not a;
    layer4_outputs(8316) <= a;
    layer4_outputs(8317) <= b and not a;
    layer4_outputs(8318) <= not a;
    layer4_outputs(8319) <= a or b;
    layer4_outputs(8320) <= not b;
    layer4_outputs(8321) <= a xor b;
    layer4_outputs(8322) <= a;
    layer4_outputs(8323) <= not b or a;
    layer4_outputs(8324) <= a;
    layer4_outputs(8325) <= a;
    layer4_outputs(8326) <= not a;
    layer4_outputs(8327) <= not b;
    layer4_outputs(8328) <= a xor b;
    layer4_outputs(8329) <= b and not a;
    layer4_outputs(8330) <= not a;
    layer4_outputs(8331) <= not (a or b);
    layer4_outputs(8332) <= not (a or b);
    layer4_outputs(8333) <= not a or b;
    layer4_outputs(8334) <= not b or a;
    layer4_outputs(8335) <= not (a or b);
    layer4_outputs(8336) <= a xor b;
    layer4_outputs(8337) <= a or b;
    layer4_outputs(8338) <= a and not b;
    layer4_outputs(8339) <= a xor b;
    layer4_outputs(8340) <= '1';
    layer4_outputs(8341) <= a;
    layer4_outputs(8342) <= b;
    layer4_outputs(8343) <= b and not a;
    layer4_outputs(8344) <= a and b;
    layer4_outputs(8345) <= not b;
    layer4_outputs(8346) <= not b or a;
    layer4_outputs(8347) <= a xor b;
    layer4_outputs(8348) <= a and not b;
    layer4_outputs(8349) <= not b;
    layer4_outputs(8350) <= a;
    layer4_outputs(8351) <= a and not b;
    layer4_outputs(8352) <= a or b;
    layer4_outputs(8353) <= not a;
    layer4_outputs(8354) <= a and b;
    layer4_outputs(8355) <= not b or a;
    layer4_outputs(8356) <= not (a and b);
    layer4_outputs(8357) <= a and not b;
    layer4_outputs(8358) <= a or b;
    layer4_outputs(8359) <= not a or b;
    layer4_outputs(8360) <= a or b;
    layer4_outputs(8361) <= '1';
    layer4_outputs(8362) <= not a or b;
    layer4_outputs(8363) <= not b or a;
    layer4_outputs(8364) <= not (a xor b);
    layer4_outputs(8365) <= not b;
    layer4_outputs(8366) <= b;
    layer4_outputs(8367) <= not b;
    layer4_outputs(8368) <= a xor b;
    layer4_outputs(8369) <= not (a and b);
    layer4_outputs(8370) <= a or b;
    layer4_outputs(8371) <= not (a and b);
    layer4_outputs(8372) <= a xor b;
    layer4_outputs(8373) <= '1';
    layer4_outputs(8374) <= not (a and b);
    layer4_outputs(8375) <= a or b;
    layer4_outputs(8376) <= not b;
    layer4_outputs(8377) <= a or b;
    layer4_outputs(8378) <= not b;
    layer4_outputs(8379) <= a and not b;
    layer4_outputs(8380) <= a or b;
    layer4_outputs(8381) <= not a;
    layer4_outputs(8382) <= not b;
    layer4_outputs(8383) <= b and not a;
    layer4_outputs(8384) <= not a;
    layer4_outputs(8385) <= b and not a;
    layer4_outputs(8386) <= not b;
    layer4_outputs(8387) <= b;
    layer4_outputs(8388) <= not (a or b);
    layer4_outputs(8389) <= a xor b;
    layer4_outputs(8390) <= a xor b;
    layer4_outputs(8391) <= a and not b;
    layer4_outputs(8392) <= not b;
    layer4_outputs(8393) <= a xor b;
    layer4_outputs(8394) <= a or b;
    layer4_outputs(8395) <= not b;
    layer4_outputs(8396) <= a xor b;
    layer4_outputs(8397) <= not b;
    layer4_outputs(8398) <= not (a or b);
    layer4_outputs(8399) <= not a;
    layer4_outputs(8400) <= not b;
    layer4_outputs(8401) <= a and b;
    layer4_outputs(8402) <= not (a xor b);
    layer4_outputs(8403) <= a xor b;
    layer4_outputs(8404) <= a;
    layer4_outputs(8405) <= a and not b;
    layer4_outputs(8406) <= not (a and b);
    layer4_outputs(8407) <= b and not a;
    layer4_outputs(8408) <= not b;
    layer4_outputs(8409) <= not a;
    layer4_outputs(8410) <= not (a and b);
    layer4_outputs(8411) <= a;
    layer4_outputs(8412) <= not b or a;
    layer4_outputs(8413) <= b;
    layer4_outputs(8414) <= a or b;
    layer4_outputs(8415) <= a;
    layer4_outputs(8416) <= a and b;
    layer4_outputs(8417) <= b;
    layer4_outputs(8418) <= not a or b;
    layer4_outputs(8419) <= a xor b;
    layer4_outputs(8420) <= '1';
    layer4_outputs(8421) <= a xor b;
    layer4_outputs(8422) <= a and not b;
    layer4_outputs(8423) <= not (a or b);
    layer4_outputs(8424) <= a and b;
    layer4_outputs(8425) <= not (a or b);
    layer4_outputs(8426) <= a;
    layer4_outputs(8427) <= b and not a;
    layer4_outputs(8428) <= b and not a;
    layer4_outputs(8429) <= not a;
    layer4_outputs(8430) <= b;
    layer4_outputs(8431) <= a;
    layer4_outputs(8432) <= '0';
    layer4_outputs(8433) <= b;
    layer4_outputs(8434) <= b;
    layer4_outputs(8435) <= not (a or b);
    layer4_outputs(8436) <= not (a and b);
    layer4_outputs(8437) <= a and b;
    layer4_outputs(8438) <= not (a xor b);
    layer4_outputs(8439) <= not (a xor b);
    layer4_outputs(8440) <= b;
    layer4_outputs(8441) <= b;
    layer4_outputs(8442) <= a or b;
    layer4_outputs(8443) <= a or b;
    layer4_outputs(8444) <= not a or b;
    layer4_outputs(8445) <= not a;
    layer4_outputs(8446) <= not b or a;
    layer4_outputs(8447) <= not b;
    layer4_outputs(8448) <= a xor b;
    layer4_outputs(8449) <= not b;
    layer4_outputs(8450) <= a and not b;
    layer4_outputs(8451) <= b;
    layer4_outputs(8452) <= not (a xor b);
    layer4_outputs(8453) <= not (a xor b);
    layer4_outputs(8454) <= not b;
    layer4_outputs(8455) <= b;
    layer4_outputs(8456) <= b and not a;
    layer4_outputs(8457) <= b;
    layer4_outputs(8458) <= not b or a;
    layer4_outputs(8459) <= not b;
    layer4_outputs(8460) <= not a;
    layer4_outputs(8461) <= not (a xor b);
    layer4_outputs(8462) <= b and not a;
    layer4_outputs(8463) <= not a or b;
    layer4_outputs(8464) <= not b;
    layer4_outputs(8465) <= b;
    layer4_outputs(8466) <= a;
    layer4_outputs(8467) <= a xor b;
    layer4_outputs(8468) <= b;
    layer4_outputs(8469) <= a or b;
    layer4_outputs(8470) <= a or b;
    layer4_outputs(8471) <= not b or a;
    layer4_outputs(8472) <= '0';
    layer4_outputs(8473) <= not b or a;
    layer4_outputs(8474) <= b and not a;
    layer4_outputs(8475) <= b;
    layer4_outputs(8476) <= a and b;
    layer4_outputs(8477) <= not b;
    layer4_outputs(8478) <= a;
    layer4_outputs(8479) <= not b or a;
    layer4_outputs(8480) <= not a;
    layer4_outputs(8481) <= not a;
    layer4_outputs(8482) <= '0';
    layer4_outputs(8483) <= '1';
    layer4_outputs(8484) <= b and not a;
    layer4_outputs(8485) <= a or b;
    layer4_outputs(8486) <= a or b;
    layer4_outputs(8487) <= b and not a;
    layer4_outputs(8488) <= not (a xor b);
    layer4_outputs(8489) <= not (a or b);
    layer4_outputs(8490) <= not (a and b);
    layer4_outputs(8491) <= a and b;
    layer4_outputs(8492) <= not a;
    layer4_outputs(8493) <= not a;
    layer4_outputs(8494) <= not a;
    layer4_outputs(8495) <= b and not a;
    layer4_outputs(8496) <= not b or a;
    layer4_outputs(8497) <= b and not a;
    layer4_outputs(8498) <= not b;
    layer4_outputs(8499) <= not b;
    layer4_outputs(8500) <= a and b;
    layer4_outputs(8501) <= not a;
    layer4_outputs(8502) <= not a;
    layer4_outputs(8503) <= not b;
    layer4_outputs(8504) <= a;
    layer4_outputs(8505) <= not b;
    layer4_outputs(8506) <= '1';
    layer4_outputs(8507) <= not b;
    layer4_outputs(8508) <= not a or b;
    layer4_outputs(8509) <= a or b;
    layer4_outputs(8510) <= not a;
    layer4_outputs(8511) <= not a;
    layer4_outputs(8512) <= not b;
    layer4_outputs(8513) <= b;
    layer4_outputs(8514) <= not b or a;
    layer4_outputs(8515) <= not b;
    layer4_outputs(8516) <= not a;
    layer4_outputs(8517) <= a xor b;
    layer4_outputs(8518) <= a;
    layer4_outputs(8519) <= b;
    layer4_outputs(8520) <= a and not b;
    layer4_outputs(8521) <= a;
    layer4_outputs(8522) <= not b;
    layer4_outputs(8523) <= not b or a;
    layer4_outputs(8524) <= a;
    layer4_outputs(8525) <= a;
    layer4_outputs(8526) <= a and b;
    layer4_outputs(8527) <= not b;
    layer4_outputs(8528) <= not b or a;
    layer4_outputs(8529) <= a xor b;
    layer4_outputs(8530) <= a;
    layer4_outputs(8531) <= b;
    layer4_outputs(8532) <= not b;
    layer4_outputs(8533) <= b;
    layer4_outputs(8534) <= not b;
    layer4_outputs(8535) <= a;
    layer4_outputs(8536) <= a or b;
    layer4_outputs(8537) <= not b;
    layer4_outputs(8538) <= '0';
    layer4_outputs(8539) <= not (a xor b);
    layer4_outputs(8540) <= not b;
    layer4_outputs(8541) <= not b;
    layer4_outputs(8542) <= a and b;
    layer4_outputs(8543) <= not b;
    layer4_outputs(8544) <= a and b;
    layer4_outputs(8545) <= a and b;
    layer4_outputs(8546) <= a and b;
    layer4_outputs(8547) <= not (a and b);
    layer4_outputs(8548) <= not a;
    layer4_outputs(8549) <= not (a or b);
    layer4_outputs(8550) <= a xor b;
    layer4_outputs(8551) <= a;
    layer4_outputs(8552) <= a and not b;
    layer4_outputs(8553) <= a and not b;
    layer4_outputs(8554) <= a or b;
    layer4_outputs(8555) <= b;
    layer4_outputs(8556) <= not (a or b);
    layer4_outputs(8557) <= not b or a;
    layer4_outputs(8558) <= not a or b;
    layer4_outputs(8559) <= not (a xor b);
    layer4_outputs(8560) <= '1';
    layer4_outputs(8561) <= a or b;
    layer4_outputs(8562) <= a xor b;
    layer4_outputs(8563) <= not b;
    layer4_outputs(8564) <= a and not b;
    layer4_outputs(8565) <= a;
    layer4_outputs(8566) <= not b;
    layer4_outputs(8567) <= not (a and b);
    layer4_outputs(8568) <= a and b;
    layer4_outputs(8569) <= not a;
    layer4_outputs(8570) <= not b;
    layer4_outputs(8571) <= not (a or b);
    layer4_outputs(8572) <= b and not a;
    layer4_outputs(8573) <= a;
    layer4_outputs(8574) <= b;
    layer4_outputs(8575) <= not b;
    layer4_outputs(8576) <= not a;
    layer4_outputs(8577) <= not b or a;
    layer4_outputs(8578) <= a xor b;
    layer4_outputs(8579) <= not (a and b);
    layer4_outputs(8580) <= a;
    layer4_outputs(8581) <= not (a xor b);
    layer4_outputs(8582) <= not (a and b);
    layer4_outputs(8583) <= b;
    layer4_outputs(8584) <= a and b;
    layer4_outputs(8585) <= a or b;
    layer4_outputs(8586) <= b and not a;
    layer4_outputs(8587) <= a xor b;
    layer4_outputs(8588) <= a xor b;
    layer4_outputs(8589) <= a and b;
    layer4_outputs(8590) <= a;
    layer4_outputs(8591) <= not a;
    layer4_outputs(8592) <= b;
    layer4_outputs(8593) <= a or b;
    layer4_outputs(8594) <= a;
    layer4_outputs(8595) <= not (a xor b);
    layer4_outputs(8596) <= b;
    layer4_outputs(8597) <= not a;
    layer4_outputs(8598) <= not a;
    layer4_outputs(8599) <= not b or a;
    layer4_outputs(8600) <= '1';
    layer4_outputs(8601) <= a xor b;
    layer4_outputs(8602) <= b;
    layer4_outputs(8603) <= a and b;
    layer4_outputs(8604) <= not a or b;
    layer4_outputs(8605) <= not a or b;
    layer4_outputs(8606) <= b and not a;
    layer4_outputs(8607) <= a;
    layer4_outputs(8608) <= not b;
    layer4_outputs(8609) <= '0';
    layer4_outputs(8610) <= not b;
    layer4_outputs(8611) <= not (a xor b);
    layer4_outputs(8612) <= not (a xor b);
    layer4_outputs(8613) <= not b;
    layer4_outputs(8614) <= a and b;
    layer4_outputs(8615) <= not (a and b);
    layer4_outputs(8616) <= b;
    layer4_outputs(8617) <= not (a and b);
    layer4_outputs(8618) <= '0';
    layer4_outputs(8619) <= b;
    layer4_outputs(8620) <= a;
    layer4_outputs(8621) <= a and b;
    layer4_outputs(8622) <= b;
    layer4_outputs(8623) <= not a;
    layer4_outputs(8624) <= not b;
    layer4_outputs(8625) <= not a;
    layer4_outputs(8626) <= a xor b;
    layer4_outputs(8627) <= b;
    layer4_outputs(8628) <= not (a xor b);
    layer4_outputs(8629) <= not b;
    layer4_outputs(8630) <= not (a xor b);
    layer4_outputs(8631) <= not b;
    layer4_outputs(8632) <= a;
    layer4_outputs(8633) <= not (a and b);
    layer4_outputs(8634) <= a and not b;
    layer4_outputs(8635) <= a;
    layer4_outputs(8636) <= not (a xor b);
    layer4_outputs(8637) <= a and not b;
    layer4_outputs(8638) <= not a;
    layer4_outputs(8639) <= a or b;
    layer4_outputs(8640) <= not a or b;
    layer4_outputs(8641) <= a and b;
    layer4_outputs(8642) <= a and b;
    layer4_outputs(8643) <= a or b;
    layer4_outputs(8644) <= not (a and b);
    layer4_outputs(8645) <= not b;
    layer4_outputs(8646) <= not b;
    layer4_outputs(8647) <= not b or a;
    layer4_outputs(8648) <= a and not b;
    layer4_outputs(8649) <= not b;
    layer4_outputs(8650) <= not (a or b);
    layer4_outputs(8651) <= not a;
    layer4_outputs(8652) <= not a or b;
    layer4_outputs(8653) <= not b or a;
    layer4_outputs(8654) <= b;
    layer4_outputs(8655) <= not (a or b);
    layer4_outputs(8656) <= not a;
    layer4_outputs(8657) <= not (a or b);
    layer4_outputs(8658) <= a;
    layer4_outputs(8659) <= a and b;
    layer4_outputs(8660) <= not b or a;
    layer4_outputs(8661) <= not b;
    layer4_outputs(8662) <= not a;
    layer4_outputs(8663) <= '0';
    layer4_outputs(8664) <= not b or a;
    layer4_outputs(8665) <= not a;
    layer4_outputs(8666) <= b and not a;
    layer4_outputs(8667) <= b;
    layer4_outputs(8668) <= a and b;
    layer4_outputs(8669) <= b;
    layer4_outputs(8670) <= b and not a;
    layer4_outputs(8671) <= not (a or b);
    layer4_outputs(8672) <= not (a or b);
    layer4_outputs(8673) <= a;
    layer4_outputs(8674) <= not (a or b);
    layer4_outputs(8675) <= not (a or b);
    layer4_outputs(8676) <= not a;
    layer4_outputs(8677) <= '0';
    layer4_outputs(8678) <= '0';
    layer4_outputs(8679) <= not (a xor b);
    layer4_outputs(8680) <= not (a or b);
    layer4_outputs(8681) <= '0';
    layer4_outputs(8682) <= a;
    layer4_outputs(8683) <= not b;
    layer4_outputs(8684) <= not b;
    layer4_outputs(8685) <= not (a or b);
    layer4_outputs(8686) <= a and not b;
    layer4_outputs(8687) <= not b;
    layer4_outputs(8688) <= not a or b;
    layer4_outputs(8689) <= a and b;
    layer4_outputs(8690) <= not b or a;
    layer4_outputs(8691) <= not b or a;
    layer4_outputs(8692) <= a and not b;
    layer4_outputs(8693) <= not a;
    layer4_outputs(8694) <= not (a or b);
    layer4_outputs(8695) <= a;
    layer4_outputs(8696) <= not a or b;
    layer4_outputs(8697) <= a and b;
    layer4_outputs(8698) <= a;
    layer4_outputs(8699) <= a and not b;
    layer4_outputs(8700) <= a;
    layer4_outputs(8701) <= b;
    layer4_outputs(8702) <= a xor b;
    layer4_outputs(8703) <= a xor b;
    layer4_outputs(8704) <= not (a and b);
    layer4_outputs(8705) <= not a;
    layer4_outputs(8706) <= not a or b;
    layer4_outputs(8707) <= b;
    layer4_outputs(8708) <= b;
    layer4_outputs(8709) <= a and b;
    layer4_outputs(8710) <= not (a and b);
    layer4_outputs(8711) <= a;
    layer4_outputs(8712) <= '1';
    layer4_outputs(8713) <= not (a and b);
    layer4_outputs(8714) <= not b;
    layer4_outputs(8715) <= not a or b;
    layer4_outputs(8716) <= b;
    layer4_outputs(8717) <= not b or a;
    layer4_outputs(8718) <= not b;
    layer4_outputs(8719) <= not b;
    layer4_outputs(8720) <= not (a or b);
    layer4_outputs(8721) <= not b or a;
    layer4_outputs(8722) <= b;
    layer4_outputs(8723) <= not a or b;
    layer4_outputs(8724) <= a;
    layer4_outputs(8725) <= not a or b;
    layer4_outputs(8726) <= a xor b;
    layer4_outputs(8727) <= a or b;
    layer4_outputs(8728) <= not (a or b);
    layer4_outputs(8729) <= not a or b;
    layer4_outputs(8730) <= not a;
    layer4_outputs(8731) <= a and not b;
    layer4_outputs(8732) <= a or b;
    layer4_outputs(8733) <= '0';
    layer4_outputs(8734) <= a or b;
    layer4_outputs(8735) <= b;
    layer4_outputs(8736) <= a and not b;
    layer4_outputs(8737) <= a and not b;
    layer4_outputs(8738) <= not a or b;
    layer4_outputs(8739) <= a;
    layer4_outputs(8740) <= '0';
    layer4_outputs(8741) <= a and b;
    layer4_outputs(8742) <= a and not b;
    layer4_outputs(8743) <= b;
    layer4_outputs(8744) <= not (a or b);
    layer4_outputs(8745) <= not b;
    layer4_outputs(8746) <= a;
    layer4_outputs(8747) <= a or b;
    layer4_outputs(8748) <= not (a xor b);
    layer4_outputs(8749) <= '0';
    layer4_outputs(8750) <= a and b;
    layer4_outputs(8751) <= b and not a;
    layer4_outputs(8752) <= not b;
    layer4_outputs(8753) <= a and b;
    layer4_outputs(8754) <= not (a or b);
    layer4_outputs(8755) <= b;
    layer4_outputs(8756) <= not (a xor b);
    layer4_outputs(8757) <= a or b;
    layer4_outputs(8758) <= not (a or b);
    layer4_outputs(8759) <= a xor b;
    layer4_outputs(8760) <= not a;
    layer4_outputs(8761) <= not a;
    layer4_outputs(8762) <= a xor b;
    layer4_outputs(8763) <= not a or b;
    layer4_outputs(8764) <= not b;
    layer4_outputs(8765) <= a and not b;
    layer4_outputs(8766) <= b;
    layer4_outputs(8767) <= not (a and b);
    layer4_outputs(8768) <= not a;
    layer4_outputs(8769) <= not a or b;
    layer4_outputs(8770) <= not a;
    layer4_outputs(8771) <= a;
    layer4_outputs(8772) <= not a or b;
    layer4_outputs(8773) <= not b or a;
    layer4_outputs(8774) <= a and b;
    layer4_outputs(8775) <= b and not a;
    layer4_outputs(8776) <= a and not b;
    layer4_outputs(8777) <= a xor b;
    layer4_outputs(8778) <= b and not a;
    layer4_outputs(8779) <= a or b;
    layer4_outputs(8780) <= b and not a;
    layer4_outputs(8781) <= a;
    layer4_outputs(8782) <= not a or b;
    layer4_outputs(8783) <= not b or a;
    layer4_outputs(8784) <= a and not b;
    layer4_outputs(8785) <= not (a or b);
    layer4_outputs(8786) <= not a;
    layer4_outputs(8787) <= a and b;
    layer4_outputs(8788) <= not a;
    layer4_outputs(8789) <= not (a or b);
    layer4_outputs(8790) <= not a;
    layer4_outputs(8791) <= not a;
    layer4_outputs(8792) <= a and not b;
    layer4_outputs(8793) <= a;
    layer4_outputs(8794) <= not b;
    layer4_outputs(8795) <= not b;
    layer4_outputs(8796) <= not (a and b);
    layer4_outputs(8797) <= b and not a;
    layer4_outputs(8798) <= a;
    layer4_outputs(8799) <= a and not b;
    layer4_outputs(8800) <= not (a and b);
    layer4_outputs(8801) <= a or b;
    layer4_outputs(8802) <= not a;
    layer4_outputs(8803) <= b;
    layer4_outputs(8804) <= not b;
    layer4_outputs(8805) <= '1';
    layer4_outputs(8806) <= b;
    layer4_outputs(8807) <= a and b;
    layer4_outputs(8808) <= not b or a;
    layer4_outputs(8809) <= not (a xor b);
    layer4_outputs(8810) <= b and not a;
    layer4_outputs(8811) <= a and b;
    layer4_outputs(8812) <= '1';
    layer4_outputs(8813) <= not (a or b);
    layer4_outputs(8814) <= not (a or b);
    layer4_outputs(8815) <= a;
    layer4_outputs(8816) <= b;
    layer4_outputs(8817) <= not (a or b);
    layer4_outputs(8818) <= a;
    layer4_outputs(8819) <= a and not b;
    layer4_outputs(8820) <= a and not b;
    layer4_outputs(8821) <= not (a xor b);
    layer4_outputs(8822) <= b;
    layer4_outputs(8823) <= not a or b;
    layer4_outputs(8824) <= a and b;
    layer4_outputs(8825) <= not (a or b);
    layer4_outputs(8826) <= not (a or b);
    layer4_outputs(8827) <= a;
    layer4_outputs(8828) <= not b or a;
    layer4_outputs(8829) <= not a or b;
    layer4_outputs(8830) <= not b or a;
    layer4_outputs(8831) <= a and b;
    layer4_outputs(8832) <= not b;
    layer4_outputs(8833) <= not b;
    layer4_outputs(8834) <= a;
    layer4_outputs(8835) <= not a;
    layer4_outputs(8836) <= not (a and b);
    layer4_outputs(8837) <= a;
    layer4_outputs(8838) <= a;
    layer4_outputs(8839) <= not a;
    layer4_outputs(8840) <= not (a and b);
    layer4_outputs(8841) <= b and not a;
    layer4_outputs(8842) <= not b;
    layer4_outputs(8843) <= not (a and b);
    layer4_outputs(8844) <= not b;
    layer4_outputs(8845) <= a and not b;
    layer4_outputs(8846) <= not a;
    layer4_outputs(8847) <= a and b;
    layer4_outputs(8848) <= not b;
    layer4_outputs(8849) <= a xor b;
    layer4_outputs(8850) <= not b or a;
    layer4_outputs(8851) <= not (a and b);
    layer4_outputs(8852) <= not a;
    layer4_outputs(8853) <= not b;
    layer4_outputs(8854) <= not (a and b);
    layer4_outputs(8855) <= not (a or b);
    layer4_outputs(8856) <= b and not a;
    layer4_outputs(8857) <= a;
    layer4_outputs(8858) <= '0';
    layer4_outputs(8859) <= a and not b;
    layer4_outputs(8860) <= not b;
    layer4_outputs(8861) <= not (a or b);
    layer4_outputs(8862) <= not b;
    layer4_outputs(8863) <= not b or a;
    layer4_outputs(8864) <= b and not a;
    layer4_outputs(8865) <= b;
    layer4_outputs(8866) <= a or b;
    layer4_outputs(8867) <= b;
    layer4_outputs(8868) <= '0';
    layer4_outputs(8869) <= b and not a;
    layer4_outputs(8870) <= not b or a;
    layer4_outputs(8871) <= '0';
    layer4_outputs(8872) <= not b;
    layer4_outputs(8873) <= not a;
    layer4_outputs(8874) <= '0';
    layer4_outputs(8875) <= not a or b;
    layer4_outputs(8876) <= a;
    layer4_outputs(8877) <= b;
    layer4_outputs(8878) <= a and b;
    layer4_outputs(8879) <= not (a or b);
    layer4_outputs(8880) <= not b;
    layer4_outputs(8881) <= not b;
    layer4_outputs(8882) <= b;
    layer4_outputs(8883) <= a or b;
    layer4_outputs(8884) <= not a or b;
    layer4_outputs(8885) <= a;
    layer4_outputs(8886) <= not (a xor b);
    layer4_outputs(8887) <= a and b;
    layer4_outputs(8888) <= b and not a;
    layer4_outputs(8889) <= a and not b;
    layer4_outputs(8890) <= not (a or b);
    layer4_outputs(8891) <= not a;
    layer4_outputs(8892) <= b;
    layer4_outputs(8893) <= not b;
    layer4_outputs(8894) <= not (a or b);
    layer4_outputs(8895) <= '1';
    layer4_outputs(8896) <= a;
    layer4_outputs(8897) <= b;
    layer4_outputs(8898) <= not a;
    layer4_outputs(8899) <= b and not a;
    layer4_outputs(8900) <= not a;
    layer4_outputs(8901) <= b;
    layer4_outputs(8902) <= a and not b;
    layer4_outputs(8903) <= not a or b;
    layer4_outputs(8904) <= a xor b;
    layer4_outputs(8905) <= not b;
    layer4_outputs(8906) <= a and b;
    layer4_outputs(8907) <= b;
    layer4_outputs(8908) <= a xor b;
    layer4_outputs(8909) <= not a;
    layer4_outputs(8910) <= a xor b;
    layer4_outputs(8911) <= not (a xor b);
    layer4_outputs(8912) <= not b;
    layer4_outputs(8913) <= not (a xor b);
    layer4_outputs(8914) <= not a or b;
    layer4_outputs(8915) <= a xor b;
    layer4_outputs(8916) <= not (a and b);
    layer4_outputs(8917) <= not (a or b);
    layer4_outputs(8918) <= not b;
    layer4_outputs(8919) <= b;
    layer4_outputs(8920) <= b and not a;
    layer4_outputs(8921) <= '1';
    layer4_outputs(8922) <= not (a or b);
    layer4_outputs(8923) <= b;
    layer4_outputs(8924) <= a and not b;
    layer4_outputs(8925) <= a and not b;
    layer4_outputs(8926) <= not (a or b);
    layer4_outputs(8927) <= a or b;
    layer4_outputs(8928) <= not b or a;
    layer4_outputs(8929) <= not b;
    layer4_outputs(8930) <= not a;
    layer4_outputs(8931) <= not a or b;
    layer4_outputs(8932) <= a and not b;
    layer4_outputs(8933) <= b;
    layer4_outputs(8934) <= b;
    layer4_outputs(8935) <= b and not a;
    layer4_outputs(8936) <= '1';
    layer4_outputs(8937) <= not a or b;
    layer4_outputs(8938) <= not a or b;
    layer4_outputs(8939) <= a and not b;
    layer4_outputs(8940) <= '1';
    layer4_outputs(8941) <= b;
    layer4_outputs(8942) <= '1';
    layer4_outputs(8943) <= a and b;
    layer4_outputs(8944) <= not b or a;
    layer4_outputs(8945) <= '0';
    layer4_outputs(8946) <= not a;
    layer4_outputs(8947) <= not b or a;
    layer4_outputs(8948) <= not (a xor b);
    layer4_outputs(8949) <= a and not b;
    layer4_outputs(8950) <= a;
    layer4_outputs(8951) <= not a or b;
    layer4_outputs(8952) <= a xor b;
    layer4_outputs(8953) <= a xor b;
    layer4_outputs(8954) <= not b;
    layer4_outputs(8955) <= a;
    layer4_outputs(8956) <= '1';
    layer4_outputs(8957) <= not b;
    layer4_outputs(8958) <= not a;
    layer4_outputs(8959) <= not a or b;
    layer4_outputs(8960) <= a;
    layer4_outputs(8961) <= a and not b;
    layer4_outputs(8962) <= b;
    layer4_outputs(8963) <= not (a or b);
    layer4_outputs(8964) <= a or b;
    layer4_outputs(8965) <= not a;
    layer4_outputs(8966) <= not a;
    layer4_outputs(8967) <= not b or a;
    layer4_outputs(8968) <= not a or b;
    layer4_outputs(8969) <= a and b;
    layer4_outputs(8970) <= not b;
    layer4_outputs(8971) <= a or b;
    layer4_outputs(8972) <= a and not b;
    layer4_outputs(8973) <= not b;
    layer4_outputs(8974) <= not (a or b);
    layer4_outputs(8975) <= b;
    layer4_outputs(8976) <= not a;
    layer4_outputs(8977) <= not a;
    layer4_outputs(8978) <= a;
    layer4_outputs(8979) <= not (a xor b);
    layer4_outputs(8980) <= not b;
    layer4_outputs(8981) <= a and b;
    layer4_outputs(8982) <= a;
    layer4_outputs(8983) <= not a;
    layer4_outputs(8984) <= not (a and b);
    layer4_outputs(8985) <= b;
    layer4_outputs(8986) <= a;
    layer4_outputs(8987) <= not (a and b);
    layer4_outputs(8988) <= not (a xor b);
    layer4_outputs(8989) <= b;
    layer4_outputs(8990) <= not (a xor b);
    layer4_outputs(8991) <= b;
    layer4_outputs(8992) <= a;
    layer4_outputs(8993) <= a;
    layer4_outputs(8994) <= not a or b;
    layer4_outputs(8995) <= not (a or b);
    layer4_outputs(8996) <= not a;
    layer4_outputs(8997) <= not a or b;
    layer4_outputs(8998) <= not b;
    layer4_outputs(8999) <= a or b;
    layer4_outputs(9000) <= not (a or b);
    layer4_outputs(9001) <= b;
    layer4_outputs(9002) <= a;
    layer4_outputs(9003) <= not a or b;
    layer4_outputs(9004) <= not (a or b);
    layer4_outputs(9005) <= b;
    layer4_outputs(9006) <= not (a and b);
    layer4_outputs(9007) <= b and not a;
    layer4_outputs(9008) <= not (a xor b);
    layer4_outputs(9009) <= not b;
    layer4_outputs(9010) <= not b;
    layer4_outputs(9011) <= a xor b;
    layer4_outputs(9012) <= a;
    layer4_outputs(9013) <= not a;
    layer4_outputs(9014) <= a and b;
    layer4_outputs(9015) <= not a or b;
    layer4_outputs(9016) <= not a;
    layer4_outputs(9017) <= not b or a;
    layer4_outputs(9018) <= a;
    layer4_outputs(9019) <= not (a and b);
    layer4_outputs(9020) <= not (a xor b);
    layer4_outputs(9021) <= not b;
    layer4_outputs(9022) <= b and not a;
    layer4_outputs(9023) <= '1';
    layer4_outputs(9024) <= a xor b;
    layer4_outputs(9025) <= not a or b;
    layer4_outputs(9026) <= b and not a;
    layer4_outputs(9027) <= a and b;
    layer4_outputs(9028) <= a or b;
    layer4_outputs(9029) <= not b;
    layer4_outputs(9030) <= '0';
    layer4_outputs(9031) <= a and b;
    layer4_outputs(9032) <= not a;
    layer4_outputs(9033) <= a and not b;
    layer4_outputs(9034) <= not a or b;
    layer4_outputs(9035) <= a or b;
    layer4_outputs(9036) <= not a;
    layer4_outputs(9037) <= b;
    layer4_outputs(9038) <= not a or b;
    layer4_outputs(9039) <= a;
    layer4_outputs(9040) <= not (a and b);
    layer4_outputs(9041) <= not b or a;
    layer4_outputs(9042) <= not (a or b);
    layer4_outputs(9043) <= not b or a;
    layer4_outputs(9044) <= a and b;
    layer4_outputs(9045) <= not b;
    layer4_outputs(9046) <= not (a and b);
    layer4_outputs(9047) <= b and not a;
    layer4_outputs(9048) <= not (a or b);
    layer4_outputs(9049) <= not a;
    layer4_outputs(9050) <= a;
    layer4_outputs(9051) <= a xor b;
    layer4_outputs(9052) <= a and not b;
    layer4_outputs(9053) <= a xor b;
    layer4_outputs(9054) <= a and not b;
    layer4_outputs(9055) <= a;
    layer4_outputs(9056) <= not b or a;
    layer4_outputs(9057) <= '1';
    layer4_outputs(9058) <= not b;
    layer4_outputs(9059) <= a;
    layer4_outputs(9060) <= not a or b;
    layer4_outputs(9061) <= b;
    layer4_outputs(9062) <= not a or b;
    layer4_outputs(9063) <= '0';
    layer4_outputs(9064) <= b;
    layer4_outputs(9065) <= b;
    layer4_outputs(9066) <= b;
    layer4_outputs(9067) <= not a;
    layer4_outputs(9068) <= not (a and b);
    layer4_outputs(9069) <= not b;
    layer4_outputs(9070) <= not b or a;
    layer4_outputs(9071) <= a and not b;
    layer4_outputs(9072) <= not a;
    layer4_outputs(9073) <= not (a and b);
    layer4_outputs(9074) <= a and b;
    layer4_outputs(9075) <= a and b;
    layer4_outputs(9076) <= not b or a;
    layer4_outputs(9077) <= b;
    layer4_outputs(9078) <= not (a or b);
    layer4_outputs(9079) <= a and not b;
    layer4_outputs(9080) <= b;
    layer4_outputs(9081) <= a and b;
    layer4_outputs(9082) <= a;
    layer4_outputs(9083) <= b and not a;
    layer4_outputs(9084) <= not b;
    layer4_outputs(9085) <= '0';
    layer4_outputs(9086) <= a and not b;
    layer4_outputs(9087) <= not b;
    layer4_outputs(9088) <= a;
    layer4_outputs(9089) <= b;
    layer4_outputs(9090) <= not b;
    layer4_outputs(9091) <= not a;
    layer4_outputs(9092) <= not a or b;
    layer4_outputs(9093) <= b;
    layer4_outputs(9094) <= a;
    layer4_outputs(9095) <= a or b;
    layer4_outputs(9096) <= '0';
    layer4_outputs(9097) <= a;
    layer4_outputs(9098) <= not b or a;
    layer4_outputs(9099) <= a and not b;
    layer4_outputs(9100) <= not a;
    layer4_outputs(9101) <= b;
    layer4_outputs(9102) <= b and not a;
    layer4_outputs(9103) <= a or b;
    layer4_outputs(9104) <= a and not b;
    layer4_outputs(9105) <= a;
    layer4_outputs(9106) <= not a;
    layer4_outputs(9107) <= b and not a;
    layer4_outputs(9108) <= not b or a;
    layer4_outputs(9109) <= not (a xor b);
    layer4_outputs(9110) <= a;
    layer4_outputs(9111) <= a and b;
    layer4_outputs(9112) <= not a;
    layer4_outputs(9113) <= b;
    layer4_outputs(9114) <= not b;
    layer4_outputs(9115) <= not a or b;
    layer4_outputs(9116) <= b and not a;
    layer4_outputs(9117) <= '0';
    layer4_outputs(9118) <= not (a or b);
    layer4_outputs(9119) <= not (a xor b);
    layer4_outputs(9120) <= b and not a;
    layer4_outputs(9121) <= not (a or b);
    layer4_outputs(9122) <= not a;
    layer4_outputs(9123) <= '0';
    layer4_outputs(9124) <= a;
    layer4_outputs(9125) <= b;
    layer4_outputs(9126) <= not a or b;
    layer4_outputs(9127) <= b;
    layer4_outputs(9128) <= a;
    layer4_outputs(9129) <= a and not b;
    layer4_outputs(9130) <= not (a or b);
    layer4_outputs(9131) <= a and not b;
    layer4_outputs(9132) <= not b or a;
    layer4_outputs(9133) <= '1';
    layer4_outputs(9134) <= not (a and b);
    layer4_outputs(9135) <= not (a and b);
    layer4_outputs(9136) <= a and not b;
    layer4_outputs(9137) <= b and not a;
    layer4_outputs(9138) <= not b or a;
    layer4_outputs(9139) <= not (a and b);
    layer4_outputs(9140) <= not a;
    layer4_outputs(9141) <= b;
    layer4_outputs(9142) <= a and not b;
    layer4_outputs(9143) <= a or b;
    layer4_outputs(9144) <= b;
    layer4_outputs(9145) <= a;
    layer4_outputs(9146) <= a;
    layer4_outputs(9147) <= not a;
    layer4_outputs(9148) <= a;
    layer4_outputs(9149) <= b;
    layer4_outputs(9150) <= not a;
    layer4_outputs(9151) <= a xor b;
    layer4_outputs(9152) <= b;
    layer4_outputs(9153) <= not (a xor b);
    layer4_outputs(9154) <= b;
    layer4_outputs(9155) <= not b;
    layer4_outputs(9156) <= not b;
    layer4_outputs(9157) <= a;
    layer4_outputs(9158) <= not b;
    layer4_outputs(9159) <= a or b;
    layer4_outputs(9160) <= not a;
    layer4_outputs(9161) <= b and not a;
    layer4_outputs(9162) <= a and b;
    layer4_outputs(9163) <= not b;
    layer4_outputs(9164) <= b and not a;
    layer4_outputs(9165) <= a and not b;
    layer4_outputs(9166) <= b and not a;
    layer4_outputs(9167) <= not (a and b);
    layer4_outputs(9168) <= a and not b;
    layer4_outputs(9169) <= not a;
    layer4_outputs(9170) <= not b;
    layer4_outputs(9171) <= '0';
    layer4_outputs(9172) <= b;
    layer4_outputs(9173) <= not a;
    layer4_outputs(9174) <= not (a xor b);
    layer4_outputs(9175) <= not b;
    layer4_outputs(9176) <= not b;
    layer4_outputs(9177) <= b;
    layer4_outputs(9178) <= a or b;
    layer4_outputs(9179) <= not b;
    layer4_outputs(9180) <= not b;
    layer4_outputs(9181) <= a and not b;
    layer4_outputs(9182) <= a and b;
    layer4_outputs(9183) <= not (a or b);
    layer4_outputs(9184) <= not a;
    layer4_outputs(9185) <= a or b;
    layer4_outputs(9186) <= a and not b;
    layer4_outputs(9187) <= not a;
    layer4_outputs(9188) <= a or b;
    layer4_outputs(9189) <= b;
    layer4_outputs(9190) <= a xor b;
    layer4_outputs(9191) <= not a;
    layer4_outputs(9192) <= not b or a;
    layer4_outputs(9193) <= not (a and b);
    layer4_outputs(9194) <= not (a xor b);
    layer4_outputs(9195) <= not a or b;
    layer4_outputs(9196) <= not b or a;
    layer4_outputs(9197) <= not b;
    layer4_outputs(9198) <= not a;
    layer4_outputs(9199) <= a and not b;
    layer4_outputs(9200) <= a xor b;
    layer4_outputs(9201) <= not (a xor b);
    layer4_outputs(9202) <= not b;
    layer4_outputs(9203) <= not b;
    layer4_outputs(9204) <= a;
    layer4_outputs(9205) <= not (a and b);
    layer4_outputs(9206) <= not (a xor b);
    layer4_outputs(9207) <= not (a or b);
    layer4_outputs(9208) <= a;
    layer4_outputs(9209) <= not a;
    layer4_outputs(9210) <= a xor b;
    layer4_outputs(9211) <= b and not a;
    layer4_outputs(9212) <= b;
    layer4_outputs(9213) <= not b or a;
    layer4_outputs(9214) <= b;
    layer4_outputs(9215) <= not a or b;
    layer4_outputs(9216) <= b;
    layer4_outputs(9217) <= b;
    layer4_outputs(9218) <= not b;
    layer4_outputs(9219) <= a and not b;
    layer4_outputs(9220) <= not a;
    layer4_outputs(9221) <= a and b;
    layer4_outputs(9222) <= a or b;
    layer4_outputs(9223) <= not a;
    layer4_outputs(9224) <= b and not a;
    layer4_outputs(9225) <= not b;
    layer4_outputs(9226) <= not b;
    layer4_outputs(9227) <= a and b;
    layer4_outputs(9228) <= b;
    layer4_outputs(9229) <= not b;
    layer4_outputs(9230) <= not a;
    layer4_outputs(9231) <= a;
    layer4_outputs(9232) <= a and not b;
    layer4_outputs(9233) <= not (a xor b);
    layer4_outputs(9234) <= not (a and b);
    layer4_outputs(9235) <= not b;
    layer4_outputs(9236) <= not (a xor b);
    layer4_outputs(9237) <= a;
    layer4_outputs(9238) <= not a;
    layer4_outputs(9239) <= not a;
    layer4_outputs(9240) <= a;
    layer4_outputs(9241) <= b and not a;
    layer4_outputs(9242) <= '1';
    layer4_outputs(9243) <= not b;
    layer4_outputs(9244) <= '0';
    layer4_outputs(9245) <= a and b;
    layer4_outputs(9246) <= not a;
    layer4_outputs(9247) <= not b;
    layer4_outputs(9248) <= not b;
    layer4_outputs(9249) <= not (a or b);
    layer4_outputs(9250) <= a xor b;
    layer4_outputs(9251) <= not b or a;
    layer4_outputs(9252) <= not b;
    layer4_outputs(9253) <= not a;
    layer4_outputs(9254) <= not (a and b);
    layer4_outputs(9255) <= not a;
    layer4_outputs(9256) <= a and b;
    layer4_outputs(9257) <= not b;
    layer4_outputs(9258) <= not (a xor b);
    layer4_outputs(9259) <= a;
    layer4_outputs(9260) <= not b;
    layer4_outputs(9261) <= a;
    layer4_outputs(9262) <= not b;
    layer4_outputs(9263) <= not a;
    layer4_outputs(9264) <= b;
    layer4_outputs(9265) <= a;
    layer4_outputs(9266) <= b and not a;
    layer4_outputs(9267) <= a and not b;
    layer4_outputs(9268) <= not a;
    layer4_outputs(9269) <= b;
    layer4_outputs(9270) <= not a or b;
    layer4_outputs(9271) <= a and not b;
    layer4_outputs(9272) <= a or b;
    layer4_outputs(9273) <= not a;
    layer4_outputs(9274) <= not a;
    layer4_outputs(9275) <= not a;
    layer4_outputs(9276) <= a and b;
    layer4_outputs(9277) <= not (a and b);
    layer4_outputs(9278) <= not a;
    layer4_outputs(9279) <= '1';
    layer4_outputs(9280) <= not (a and b);
    layer4_outputs(9281) <= not a;
    layer4_outputs(9282) <= b;
    layer4_outputs(9283) <= b;
    layer4_outputs(9284) <= a;
    layer4_outputs(9285) <= a;
    layer4_outputs(9286) <= not b;
    layer4_outputs(9287) <= '0';
    layer4_outputs(9288) <= not a;
    layer4_outputs(9289) <= a and b;
    layer4_outputs(9290) <= a;
    layer4_outputs(9291) <= not a;
    layer4_outputs(9292) <= a;
    layer4_outputs(9293) <= a;
    layer4_outputs(9294) <= b;
    layer4_outputs(9295) <= not (a or b);
    layer4_outputs(9296) <= not b;
    layer4_outputs(9297) <= not (a xor b);
    layer4_outputs(9298) <= not a;
    layer4_outputs(9299) <= not (a and b);
    layer4_outputs(9300) <= a and b;
    layer4_outputs(9301) <= b;
    layer4_outputs(9302) <= not b or a;
    layer4_outputs(9303) <= not a;
    layer4_outputs(9304) <= a;
    layer4_outputs(9305) <= a;
    layer4_outputs(9306) <= a or b;
    layer4_outputs(9307) <= b and not a;
    layer4_outputs(9308) <= a or b;
    layer4_outputs(9309) <= not a;
    layer4_outputs(9310) <= a and not b;
    layer4_outputs(9311) <= not b;
    layer4_outputs(9312) <= b;
    layer4_outputs(9313) <= not b or a;
    layer4_outputs(9314) <= not b;
    layer4_outputs(9315) <= '1';
    layer4_outputs(9316) <= b;
    layer4_outputs(9317) <= not b;
    layer4_outputs(9318) <= not b or a;
    layer4_outputs(9319) <= a and b;
    layer4_outputs(9320) <= '0';
    layer4_outputs(9321) <= a;
    layer4_outputs(9322) <= not a;
    layer4_outputs(9323) <= a and not b;
    layer4_outputs(9324) <= not a or b;
    layer4_outputs(9325) <= a;
    layer4_outputs(9326) <= a and b;
    layer4_outputs(9327) <= not b or a;
    layer4_outputs(9328) <= not (a xor b);
    layer4_outputs(9329) <= b;
    layer4_outputs(9330) <= not a;
    layer4_outputs(9331) <= a xor b;
    layer4_outputs(9332) <= not a;
    layer4_outputs(9333) <= not a;
    layer4_outputs(9334) <= b;
    layer4_outputs(9335) <= a;
    layer4_outputs(9336) <= '1';
    layer4_outputs(9337) <= a;
    layer4_outputs(9338) <= '1';
    layer4_outputs(9339) <= a and not b;
    layer4_outputs(9340) <= not b or a;
    layer4_outputs(9341) <= not (a xor b);
    layer4_outputs(9342) <= not (a or b);
    layer4_outputs(9343) <= not (a or b);
    layer4_outputs(9344) <= not b;
    layer4_outputs(9345) <= a;
    layer4_outputs(9346) <= '1';
    layer4_outputs(9347) <= b and not a;
    layer4_outputs(9348) <= not (a xor b);
    layer4_outputs(9349) <= '1';
    layer4_outputs(9350) <= not a;
    layer4_outputs(9351) <= not a or b;
    layer4_outputs(9352) <= a xor b;
    layer4_outputs(9353) <= a;
    layer4_outputs(9354) <= b;
    layer4_outputs(9355) <= not (a or b);
    layer4_outputs(9356) <= a;
    layer4_outputs(9357) <= a;
    layer4_outputs(9358) <= '1';
    layer4_outputs(9359) <= not b;
    layer4_outputs(9360) <= not a;
    layer4_outputs(9361) <= a or b;
    layer4_outputs(9362) <= b;
    layer4_outputs(9363) <= not (a and b);
    layer4_outputs(9364) <= a;
    layer4_outputs(9365) <= a;
    layer4_outputs(9366) <= not a or b;
    layer4_outputs(9367) <= not a;
    layer4_outputs(9368) <= '1';
    layer4_outputs(9369) <= a xor b;
    layer4_outputs(9370) <= not b or a;
    layer4_outputs(9371) <= not b;
    layer4_outputs(9372) <= not (a and b);
    layer4_outputs(9373) <= not (a or b);
    layer4_outputs(9374) <= not a;
    layer4_outputs(9375) <= not b or a;
    layer4_outputs(9376) <= not b;
    layer4_outputs(9377) <= not a;
    layer4_outputs(9378) <= a or b;
    layer4_outputs(9379) <= a;
    layer4_outputs(9380) <= b;
    layer4_outputs(9381) <= a;
    layer4_outputs(9382) <= not b or a;
    layer4_outputs(9383) <= a and b;
    layer4_outputs(9384) <= not a or b;
    layer4_outputs(9385) <= b;
    layer4_outputs(9386) <= a and b;
    layer4_outputs(9387) <= not a;
    layer4_outputs(9388) <= not (a and b);
    layer4_outputs(9389) <= a;
    layer4_outputs(9390) <= not a;
    layer4_outputs(9391) <= not b;
    layer4_outputs(9392) <= not a;
    layer4_outputs(9393) <= not a or b;
    layer4_outputs(9394) <= not b or a;
    layer4_outputs(9395) <= not b;
    layer4_outputs(9396) <= not b;
    layer4_outputs(9397) <= a xor b;
    layer4_outputs(9398) <= a and not b;
    layer4_outputs(9399) <= a xor b;
    layer4_outputs(9400) <= not a or b;
    layer4_outputs(9401) <= not b;
    layer4_outputs(9402) <= b and not a;
    layer4_outputs(9403) <= not a or b;
    layer4_outputs(9404) <= a and b;
    layer4_outputs(9405) <= not a;
    layer4_outputs(9406) <= b;
    layer4_outputs(9407) <= not a;
    layer4_outputs(9408) <= a and b;
    layer4_outputs(9409) <= b;
    layer4_outputs(9410) <= b and not a;
    layer4_outputs(9411) <= not b;
    layer4_outputs(9412) <= a or b;
    layer4_outputs(9413) <= a;
    layer4_outputs(9414) <= a and b;
    layer4_outputs(9415) <= not b;
    layer4_outputs(9416) <= a;
    layer4_outputs(9417) <= a or b;
    layer4_outputs(9418) <= not a;
    layer4_outputs(9419) <= not b;
    layer4_outputs(9420) <= b;
    layer4_outputs(9421) <= '1';
    layer4_outputs(9422) <= b and not a;
    layer4_outputs(9423) <= not (a and b);
    layer4_outputs(9424) <= not b;
    layer4_outputs(9425) <= a;
    layer4_outputs(9426) <= a and b;
    layer4_outputs(9427) <= b;
    layer4_outputs(9428) <= not (a or b);
    layer4_outputs(9429) <= not (a or b);
    layer4_outputs(9430) <= not b;
    layer4_outputs(9431) <= a or b;
    layer4_outputs(9432) <= b and not a;
    layer4_outputs(9433) <= a;
    layer4_outputs(9434) <= '1';
    layer4_outputs(9435) <= '0';
    layer4_outputs(9436) <= a;
    layer4_outputs(9437) <= a;
    layer4_outputs(9438) <= a or b;
    layer4_outputs(9439) <= not a;
    layer4_outputs(9440) <= b and not a;
    layer4_outputs(9441) <= b;
    layer4_outputs(9442) <= not (a xor b);
    layer4_outputs(9443) <= b and not a;
    layer4_outputs(9444) <= not (a xor b);
    layer4_outputs(9445) <= b;
    layer4_outputs(9446) <= not b;
    layer4_outputs(9447) <= b;
    layer4_outputs(9448) <= not (a xor b);
    layer4_outputs(9449) <= not a;
    layer4_outputs(9450) <= not b;
    layer4_outputs(9451) <= not b;
    layer4_outputs(9452) <= a or b;
    layer4_outputs(9453) <= b;
    layer4_outputs(9454) <= '0';
    layer4_outputs(9455) <= not a or b;
    layer4_outputs(9456) <= b;
    layer4_outputs(9457) <= b;
    layer4_outputs(9458) <= a;
    layer4_outputs(9459) <= not a or b;
    layer4_outputs(9460) <= a and not b;
    layer4_outputs(9461) <= not a;
    layer4_outputs(9462) <= not a;
    layer4_outputs(9463) <= not a;
    layer4_outputs(9464) <= b and not a;
    layer4_outputs(9465) <= a;
    layer4_outputs(9466) <= not a;
    layer4_outputs(9467) <= not a or b;
    layer4_outputs(9468) <= a;
    layer4_outputs(9469) <= b;
    layer4_outputs(9470) <= a;
    layer4_outputs(9471) <= '1';
    layer4_outputs(9472) <= b;
    layer4_outputs(9473) <= not b or a;
    layer4_outputs(9474) <= '1';
    layer4_outputs(9475) <= a;
    layer4_outputs(9476) <= a xor b;
    layer4_outputs(9477) <= not a or b;
    layer4_outputs(9478) <= not b or a;
    layer4_outputs(9479) <= not a or b;
    layer4_outputs(9480) <= not b;
    layer4_outputs(9481) <= not b or a;
    layer4_outputs(9482) <= not a;
    layer4_outputs(9483) <= a and not b;
    layer4_outputs(9484) <= a xor b;
    layer4_outputs(9485) <= not a;
    layer4_outputs(9486) <= not a or b;
    layer4_outputs(9487) <= a and b;
    layer4_outputs(9488) <= a;
    layer4_outputs(9489) <= not (a or b);
    layer4_outputs(9490) <= a;
    layer4_outputs(9491) <= not b or a;
    layer4_outputs(9492) <= a;
    layer4_outputs(9493) <= not b;
    layer4_outputs(9494) <= a;
    layer4_outputs(9495) <= b;
    layer4_outputs(9496) <= b and not a;
    layer4_outputs(9497) <= not b;
    layer4_outputs(9498) <= a and not b;
    layer4_outputs(9499) <= b and not a;
    layer4_outputs(9500) <= b;
    layer4_outputs(9501) <= not a or b;
    layer4_outputs(9502) <= not (a and b);
    layer4_outputs(9503) <= not (a or b);
    layer4_outputs(9504) <= not a;
    layer4_outputs(9505) <= not b or a;
    layer4_outputs(9506) <= a and not b;
    layer4_outputs(9507) <= a or b;
    layer4_outputs(9508) <= a or b;
    layer4_outputs(9509) <= a and b;
    layer4_outputs(9510) <= not b;
    layer4_outputs(9511) <= '0';
    layer4_outputs(9512) <= a and not b;
    layer4_outputs(9513) <= a and b;
    layer4_outputs(9514) <= not b or a;
    layer4_outputs(9515) <= not b or a;
    layer4_outputs(9516) <= b and not a;
    layer4_outputs(9517) <= not (a xor b);
    layer4_outputs(9518) <= not (a and b);
    layer4_outputs(9519) <= b;
    layer4_outputs(9520) <= not (a or b);
    layer4_outputs(9521) <= a;
    layer4_outputs(9522) <= not a;
    layer4_outputs(9523) <= not b;
    layer4_outputs(9524) <= a;
    layer4_outputs(9525) <= a or b;
    layer4_outputs(9526) <= b;
    layer4_outputs(9527) <= b;
    layer4_outputs(9528) <= not (a and b);
    layer4_outputs(9529) <= b and not a;
    layer4_outputs(9530) <= a;
    layer4_outputs(9531) <= a or b;
    layer4_outputs(9532) <= not a;
    layer4_outputs(9533) <= a;
    layer4_outputs(9534) <= not b or a;
    layer4_outputs(9535) <= a and not b;
    layer4_outputs(9536) <= a;
    layer4_outputs(9537) <= not b;
    layer4_outputs(9538) <= a xor b;
    layer4_outputs(9539) <= not (a and b);
    layer4_outputs(9540) <= a;
    layer4_outputs(9541) <= b and not a;
    layer4_outputs(9542) <= a and not b;
    layer4_outputs(9543) <= not b or a;
    layer4_outputs(9544) <= not (a and b);
    layer4_outputs(9545) <= a;
    layer4_outputs(9546) <= a xor b;
    layer4_outputs(9547) <= not b;
    layer4_outputs(9548) <= a;
    layer4_outputs(9549) <= not a;
    layer4_outputs(9550) <= not b or a;
    layer4_outputs(9551) <= not a;
    layer4_outputs(9552) <= not b;
    layer4_outputs(9553) <= a;
    layer4_outputs(9554) <= not (a xor b);
    layer4_outputs(9555) <= a or b;
    layer4_outputs(9556) <= not a;
    layer4_outputs(9557) <= not b or a;
    layer4_outputs(9558) <= a;
    layer4_outputs(9559) <= a and b;
    layer4_outputs(9560) <= not a;
    layer4_outputs(9561) <= a or b;
    layer4_outputs(9562) <= a or b;
    layer4_outputs(9563) <= not (a and b);
    layer4_outputs(9564) <= a and not b;
    layer4_outputs(9565) <= a;
    layer4_outputs(9566) <= not a;
    layer4_outputs(9567) <= a and not b;
    layer4_outputs(9568) <= not b;
    layer4_outputs(9569) <= a and b;
    layer4_outputs(9570) <= b;
    layer4_outputs(9571) <= b and not a;
    layer4_outputs(9572) <= not a;
    layer4_outputs(9573) <= not a;
    layer4_outputs(9574) <= not b;
    layer4_outputs(9575) <= not a or b;
    layer4_outputs(9576) <= not (a and b);
    layer4_outputs(9577) <= not a or b;
    layer4_outputs(9578) <= not a or b;
    layer4_outputs(9579) <= not (a or b);
    layer4_outputs(9580) <= a xor b;
    layer4_outputs(9581) <= b;
    layer4_outputs(9582) <= a and b;
    layer4_outputs(9583) <= b;
    layer4_outputs(9584) <= not a or b;
    layer4_outputs(9585) <= not a;
    layer4_outputs(9586) <= a xor b;
    layer4_outputs(9587) <= not a;
    layer4_outputs(9588) <= a;
    layer4_outputs(9589) <= a;
    layer4_outputs(9590) <= not (a xor b);
    layer4_outputs(9591) <= not (a xor b);
    layer4_outputs(9592) <= b;
    layer4_outputs(9593) <= a;
    layer4_outputs(9594) <= a xor b;
    layer4_outputs(9595) <= not (a xor b);
    layer4_outputs(9596) <= not b or a;
    layer4_outputs(9597) <= a xor b;
    layer4_outputs(9598) <= a and b;
    layer4_outputs(9599) <= not a;
    layer4_outputs(9600) <= a;
    layer4_outputs(9601) <= b and not a;
    layer4_outputs(9602) <= a and b;
    layer4_outputs(9603) <= '1';
    layer4_outputs(9604) <= b and not a;
    layer4_outputs(9605) <= '0';
    layer4_outputs(9606) <= a;
    layer4_outputs(9607) <= a and not b;
    layer4_outputs(9608) <= a;
    layer4_outputs(9609) <= a xor b;
    layer4_outputs(9610) <= b;
    layer4_outputs(9611) <= a and not b;
    layer4_outputs(9612) <= not (a or b);
    layer4_outputs(9613) <= not b or a;
    layer4_outputs(9614) <= not b or a;
    layer4_outputs(9615) <= a;
    layer4_outputs(9616) <= not a;
    layer4_outputs(9617) <= not a;
    layer4_outputs(9618) <= not (a and b);
    layer4_outputs(9619) <= a;
    layer4_outputs(9620) <= not a or b;
    layer4_outputs(9621) <= not a or b;
    layer4_outputs(9622) <= a and b;
    layer4_outputs(9623) <= not a;
    layer4_outputs(9624) <= a and not b;
    layer4_outputs(9625) <= a xor b;
    layer4_outputs(9626) <= a xor b;
    layer4_outputs(9627) <= a or b;
    layer4_outputs(9628) <= not b;
    layer4_outputs(9629) <= not a or b;
    layer4_outputs(9630) <= a or b;
    layer4_outputs(9631) <= a xor b;
    layer4_outputs(9632) <= b;
    layer4_outputs(9633) <= a;
    layer4_outputs(9634) <= not b;
    layer4_outputs(9635) <= not a;
    layer4_outputs(9636) <= a xor b;
    layer4_outputs(9637) <= a and not b;
    layer4_outputs(9638) <= not (a and b);
    layer4_outputs(9639) <= a;
    layer4_outputs(9640) <= not a;
    layer4_outputs(9641) <= '0';
    layer4_outputs(9642) <= not b;
    layer4_outputs(9643) <= a xor b;
    layer4_outputs(9644) <= a;
    layer4_outputs(9645) <= a or b;
    layer4_outputs(9646) <= not a;
    layer4_outputs(9647) <= a and b;
    layer4_outputs(9648) <= not a;
    layer4_outputs(9649) <= not (a and b);
    layer4_outputs(9650) <= not a;
    layer4_outputs(9651) <= not b or a;
    layer4_outputs(9652) <= a;
    layer4_outputs(9653) <= not a;
    layer4_outputs(9654) <= a xor b;
    layer4_outputs(9655) <= a or b;
    layer4_outputs(9656) <= not a;
    layer4_outputs(9657) <= a;
    layer4_outputs(9658) <= b and not a;
    layer4_outputs(9659) <= not b;
    layer4_outputs(9660) <= b and not a;
    layer4_outputs(9661) <= not (a and b);
    layer4_outputs(9662) <= b and not a;
    layer4_outputs(9663) <= a and b;
    layer4_outputs(9664) <= a or b;
    layer4_outputs(9665) <= '0';
    layer4_outputs(9666) <= '0';
    layer4_outputs(9667) <= not (a xor b);
    layer4_outputs(9668) <= b;
    layer4_outputs(9669) <= not (a or b);
    layer4_outputs(9670) <= '1';
    layer4_outputs(9671) <= a;
    layer4_outputs(9672) <= '1';
    layer4_outputs(9673) <= not a;
    layer4_outputs(9674) <= not (a or b);
    layer4_outputs(9675) <= not b or a;
    layer4_outputs(9676) <= not (a and b);
    layer4_outputs(9677) <= not (a or b);
    layer4_outputs(9678) <= a;
    layer4_outputs(9679) <= not b or a;
    layer4_outputs(9680) <= not a or b;
    layer4_outputs(9681) <= not (a or b);
    layer4_outputs(9682) <= not b;
    layer4_outputs(9683) <= a;
    layer4_outputs(9684) <= '1';
    layer4_outputs(9685) <= not b;
    layer4_outputs(9686) <= not b or a;
    layer4_outputs(9687) <= b;
    layer4_outputs(9688) <= '0';
    layer4_outputs(9689) <= not (a or b);
    layer4_outputs(9690) <= a and b;
    layer4_outputs(9691) <= a;
    layer4_outputs(9692) <= a;
    layer4_outputs(9693) <= not a;
    layer4_outputs(9694) <= not (a or b);
    layer4_outputs(9695) <= not b or a;
    layer4_outputs(9696) <= a and not b;
    layer4_outputs(9697) <= b and not a;
    layer4_outputs(9698) <= a;
    layer4_outputs(9699) <= a;
    layer4_outputs(9700) <= not (a or b);
    layer4_outputs(9701) <= a xor b;
    layer4_outputs(9702) <= b and not a;
    layer4_outputs(9703) <= a xor b;
    layer4_outputs(9704) <= not (a and b);
    layer4_outputs(9705) <= not (a and b);
    layer4_outputs(9706) <= not a or b;
    layer4_outputs(9707) <= not (a or b);
    layer4_outputs(9708) <= not a;
    layer4_outputs(9709) <= not b or a;
    layer4_outputs(9710) <= not (a xor b);
    layer4_outputs(9711) <= not b;
    layer4_outputs(9712) <= not b;
    layer4_outputs(9713) <= b and not a;
    layer4_outputs(9714) <= a and b;
    layer4_outputs(9715) <= not (a xor b);
    layer4_outputs(9716) <= a xor b;
    layer4_outputs(9717) <= b and not a;
    layer4_outputs(9718) <= not a or b;
    layer4_outputs(9719) <= a or b;
    layer4_outputs(9720) <= not b or a;
    layer4_outputs(9721) <= not a;
    layer4_outputs(9722) <= not b or a;
    layer4_outputs(9723) <= not a;
    layer4_outputs(9724) <= '0';
    layer4_outputs(9725) <= a and b;
    layer4_outputs(9726) <= '1';
    layer4_outputs(9727) <= b;
    layer4_outputs(9728) <= a or b;
    layer4_outputs(9729) <= not b or a;
    layer4_outputs(9730) <= a and not b;
    layer4_outputs(9731) <= not b or a;
    layer4_outputs(9732) <= not b or a;
    layer4_outputs(9733) <= a;
    layer4_outputs(9734) <= a and b;
    layer4_outputs(9735) <= not (a xor b);
    layer4_outputs(9736) <= a xor b;
    layer4_outputs(9737) <= b;
    layer4_outputs(9738) <= not b;
    layer4_outputs(9739) <= a xor b;
    layer4_outputs(9740) <= not a;
    layer4_outputs(9741) <= not b or a;
    layer4_outputs(9742) <= b and not a;
    layer4_outputs(9743) <= not b;
    layer4_outputs(9744) <= not b;
    layer4_outputs(9745) <= a or b;
    layer4_outputs(9746) <= a xor b;
    layer4_outputs(9747) <= a;
    layer4_outputs(9748) <= a or b;
    layer4_outputs(9749) <= a;
    layer4_outputs(9750) <= a;
    layer4_outputs(9751) <= '1';
    layer4_outputs(9752) <= a and not b;
    layer4_outputs(9753) <= b;
    layer4_outputs(9754) <= not a;
    layer4_outputs(9755) <= not (a or b);
    layer4_outputs(9756) <= '0';
    layer4_outputs(9757) <= b and not a;
    layer4_outputs(9758) <= not b or a;
    layer4_outputs(9759) <= not (a or b);
    layer4_outputs(9760) <= not (a xor b);
    layer4_outputs(9761) <= a and not b;
    layer4_outputs(9762) <= a and b;
    layer4_outputs(9763) <= b;
    layer4_outputs(9764) <= not a or b;
    layer4_outputs(9765) <= not (a or b);
    layer4_outputs(9766) <= not a;
    layer4_outputs(9767) <= not (a xor b);
    layer4_outputs(9768) <= not b;
    layer4_outputs(9769) <= a;
    layer4_outputs(9770) <= a;
    layer4_outputs(9771) <= not b;
    layer4_outputs(9772) <= a;
    layer4_outputs(9773) <= '1';
    layer4_outputs(9774) <= not a or b;
    layer4_outputs(9775) <= a and not b;
    layer4_outputs(9776) <= not (a xor b);
    layer4_outputs(9777) <= a and b;
    layer4_outputs(9778) <= b;
    layer4_outputs(9779) <= a and b;
    layer4_outputs(9780) <= b;
    layer4_outputs(9781) <= not a;
    layer4_outputs(9782) <= not (a and b);
    layer4_outputs(9783) <= '0';
    layer4_outputs(9784) <= a or b;
    layer4_outputs(9785) <= not (a and b);
    layer4_outputs(9786) <= not (a or b);
    layer4_outputs(9787) <= not a;
    layer4_outputs(9788) <= not b or a;
    layer4_outputs(9789) <= not (a xor b);
    layer4_outputs(9790) <= not (a or b);
    layer4_outputs(9791) <= a;
    layer4_outputs(9792) <= a and not b;
    layer4_outputs(9793) <= a;
    layer4_outputs(9794) <= not a;
    layer4_outputs(9795) <= b and not a;
    layer4_outputs(9796) <= b and not a;
    layer4_outputs(9797) <= a;
    layer4_outputs(9798) <= b;
    layer4_outputs(9799) <= not b or a;
    layer4_outputs(9800) <= not b or a;
    layer4_outputs(9801) <= a;
    layer4_outputs(9802) <= a and b;
    layer4_outputs(9803) <= b;
    layer4_outputs(9804) <= not b;
    layer4_outputs(9805) <= a and not b;
    layer4_outputs(9806) <= not a or b;
    layer4_outputs(9807) <= not a or b;
    layer4_outputs(9808) <= b;
    layer4_outputs(9809) <= b and not a;
    layer4_outputs(9810) <= a;
    layer4_outputs(9811) <= not a;
    layer4_outputs(9812) <= b and not a;
    layer4_outputs(9813) <= not (a or b);
    layer4_outputs(9814) <= b;
    layer4_outputs(9815) <= not a;
    layer4_outputs(9816) <= not a or b;
    layer4_outputs(9817) <= a or b;
    layer4_outputs(9818) <= not (a and b);
    layer4_outputs(9819) <= b;
    layer4_outputs(9820) <= a and not b;
    layer4_outputs(9821) <= not b;
    layer4_outputs(9822) <= a or b;
    layer4_outputs(9823) <= a or b;
    layer4_outputs(9824) <= a;
    layer4_outputs(9825) <= a xor b;
    layer4_outputs(9826) <= not b or a;
    layer4_outputs(9827) <= not a or b;
    layer4_outputs(9828) <= not b;
    layer4_outputs(9829) <= a or b;
    layer4_outputs(9830) <= a;
    layer4_outputs(9831) <= not (a or b);
    layer4_outputs(9832) <= not (a and b);
    layer4_outputs(9833) <= a xor b;
    layer4_outputs(9834) <= a;
    layer4_outputs(9835) <= not b;
    layer4_outputs(9836) <= '0';
    layer4_outputs(9837) <= not (a or b);
    layer4_outputs(9838) <= a and not b;
    layer4_outputs(9839) <= a and not b;
    layer4_outputs(9840) <= not (a and b);
    layer4_outputs(9841) <= not b or a;
    layer4_outputs(9842) <= a and b;
    layer4_outputs(9843) <= a and not b;
    layer4_outputs(9844) <= b and not a;
    layer4_outputs(9845) <= a and b;
    layer4_outputs(9846) <= not b;
    layer4_outputs(9847) <= not a;
    layer4_outputs(9848) <= b;
    layer4_outputs(9849) <= not a;
    layer4_outputs(9850) <= a and not b;
    layer4_outputs(9851) <= a and not b;
    layer4_outputs(9852) <= not a;
    layer4_outputs(9853) <= a xor b;
    layer4_outputs(9854) <= a and not b;
    layer4_outputs(9855) <= '0';
    layer4_outputs(9856) <= not b;
    layer4_outputs(9857) <= a or b;
    layer4_outputs(9858) <= b and not a;
    layer4_outputs(9859) <= not b or a;
    layer4_outputs(9860) <= not (a or b);
    layer4_outputs(9861) <= a;
    layer4_outputs(9862) <= not b or a;
    layer4_outputs(9863) <= '1';
    layer4_outputs(9864) <= a;
    layer4_outputs(9865) <= not a;
    layer4_outputs(9866) <= a;
    layer4_outputs(9867) <= a xor b;
    layer4_outputs(9868) <= not (a and b);
    layer4_outputs(9869) <= '0';
    layer4_outputs(9870) <= b;
    layer4_outputs(9871) <= a and not b;
    layer4_outputs(9872) <= not (a or b);
    layer4_outputs(9873) <= a xor b;
    layer4_outputs(9874) <= a;
    layer4_outputs(9875) <= a and b;
    layer4_outputs(9876) <= a xor b;
    layer4_outputs(9877) <= b;
    layer4_outputs(9878) <= a and not b;
    layer4_outputs(9879) <= not a or b;
    layer4_outputs(9880) <= '1';
    layer4_outputs(9881) <= not a or b;
    layer4_outputs(9882) <= not a;
    layer4_outputs(9883) <= a or b;
    layer4_outputs(9884) <= b;
    layer4_outputs(9885) <= a and b;
    layer4_outputs(9886) <= b;
    layer4_outputs(9887) <= a and b;
    layer4_outputs(9888) <= a;
    layer4_outputs(9889) <= a and not b;
    layer4_outputs(9890) <= a or b;
    layer4_outputs(9891) <= a and b;
    layer4_outputs(9892) <= not (a or b);
    layer4_outputs(9893) <= not b;
    layer4_outputs(9894) <= '0';
    layer4_outputs(9895) <= b;
    layer4_outputs(9896) <= not b;
    layer4_outputs(9897) <= b and not a;
    layer4_outputs(9898) <= a;
    layer4_outputs(9899) <= not b;
    layer4_outputs(9900) <= not (a and b);
    layer4_outputs(9901) <= b;
    layer4_outputs(9902) <= a;
    layer4_outputs(9903) <= b;
    layer4_outputs(9904) <= not b;
    layer4_outputs(9905) <= a or b;
    layer4_outputs(9906) <= not (a and b);
    layer4_outputs(9907) <= a;
    layer4_outputs(9908) <= not (a or b);
    layer4_outputs(9909) <= a or b;
    layer4_outputs(9910) <= b;
    layer4_outputs(9911) <= not b;
    layer4_outputs(9912) <= not a or b;
    layer4_outputs(9913) <= a and not b;
    layer4_outputs(9914) <= a;
    layer4_outputs(9915) <= a xor b;
    layer4_outputs(9916) <= a;
    layer4_outputs(9917) <= b;
    layer4_outputs(9918) <= not a;
    layer4_outputs(9919) <= not a;
    layer4_outputs(9920) <= not (a or b);
    layer4_outputs(9921) <= not (a and b);
    layer4_outputs(9922) <= not b or a;
    layer4_outputs(9923) <= b;
    layer4_outputs(9924) <= not (a xor b);
    layer4_outputs(9925) <= not a or b;
    layer4_outputs(9926) <= a and not b;
    layer4_outputs(9927) <= not (a and b);
    layer4_outputs(9928) <= a and not b;
    layer4_outputs(9929) <= a xor b;
    layer4_outputs(9930) <= a and b;
    layer4_outputs(9931) <= b and not a;
    layer4_outputs(9932) <= not b or a;
    layer4_outputs(9933) <= b and not a;
    layer4_outputs(9934) <= not a or b;
    layer4_outputs(9935) <= a;
    layer4_outputs(9936) <= a and not b;
    layer4_outputs(9937) <= b;
    layer4_outputs(9938) <= a;
    layer4_outputs(9939) <= not a;
    layer4_outputs(9940) <= b;
    layer4_outputs(9941) <= not (a and b);
    layer4_outputs(9942) <= a and b;
    layer4_outputs(9943) <= a or b;
    layer4_outputs(9944) <= not b;
    layer4_outputs(9945) <= not (a and b);
    layer4_outputs(9946) <= not a or b;
    layer4_outputs(9947) <= not (a xor b);
    layer4_outputs(9948) <= not a;
    layer4_outputs(9949) <= b and not a;
    layer4_outputs(9950) <= a xor b;
    layer4_outputs(9951) <= a or b;
    layer4_outputs(9952) <= a or b;
    layer4_outputs(9953) <= b;
    layer4_outputs(9954) <= a;
    layer4_outputs(9955) <= not (a xor b);
    layer4_outputs(9956) <= a;
    layer4_outputs(9957) <= a;
    layer4_outputs(9958) <= not (a and b);
    layer4_outputs(9959) <= '1';
    layer4_outputs(9960) <= a and not b;
    layer4_outputs(9961) <= b and not a;
    layer4_outputs(9962) <= not a or b;
    layer4_outputs(9963) <= '1';
    layer4_outputs(9964) <= not a;
    layer4_outputs(9965) <= not (a xor b);
    layer4_outputs(9966) <= a and not b;
    layer4_outputs(9967) <= b;
    layer4_outputs(9968) <= a xor b;
    layer4_outputs(9969) <= not b;
    layer4_outputs(9970) <= not (a or b);
    layer4_outputs(9971) <= b;
    layer4_outputs(9972) <= not b;
    layer4_outputs(9973) <= not b;
    layer4_outputs(9974) <= not (a and b);
    layer4_outputs(9975) <= not (a or b);
    layer4_outputs(9976) <= a and b;
    layer4_outputs(9977) <= b and not a;
    layer4_outputs(9978) <= not b or a;
    layer4_outputs(9979) <= not a;
    layer4_outputs(9980) <= a xor b;
    layer4_outputs(9981) <= a and not b;
    layer4_outputs(9982) <= not a;
    layer4_outputs(9983) <= b;
    layer4_outputs(9984) <= b;
    layer4_outputs(9985) <= '1';
    layer4_outputs(9986) <= not (a and b);
    layer4_outputs(9987) <= a or b;
    layer4_outputs(9988) <= not (a or b);
    layer4_outputs(9989) <= not a;
    layer4_outputs(9990) <= b and not a;
    layer4_outputs(9991) <= b and not a;
    layer4_outputs(9992) <= a and not b;
    layer4_outputs(9993) <= a;
    layer4_outputs(9994) <= not a or b;
    layer4_outputs(9995) <= a;
    layer4_outputs(9996) <= b and not a;
    layer4_outputs(9997) <= not b;
    layer4_outputs(9998) <= not b;
    layer4_outputs(9999) <= a xor b;
    layer4_outputs(10000) <= not a or b;
    layer4_outputs(10001) <= a or b;
    layer4_outputs(10002) <= not (a or b);
    layer4_outputs(10003) <= not a or b;
    layer4_outputs(10004) <= a and b;
    layer4_outputs(10005) <= not a or b;
    layer4_outputs(10006) <= not (a and b);
    layer4_outputs(10007) <= not (a xor b);
    layer4_outputs(10008) <= not a or b;
    layer4_outputs(10009) <= not a or b;
    layer4_outputs(10010) <= a or b;
    layer4_outputs(10011) <= not a or b;
    layer4_outputs(10012) <= not (a and b);
    layer4_outputs(10013) <= b;
    layer4_outputs(10014) <= not a;
    layer4_outputs(10015) <= '0';
    layer4_outputs(10016) <= b and not a;
    layer4_outputs(10017) <= not b;
    layer4_outputs(10018) <= a and b;
    layer4_outputs(10019) <= '1';
    layer4_outputs(10020) <= b;
    layer4_outputs(10021) <= not b or a;
    layer4_outputs(10022) <= not (a or b);
    layer4_outputs(10023) <= b;
    layer4_outputs(10024) <= not b or a;
    layer4_outputs(10025) <= a and not b;
    layer4_outputs(10026) <= b;
    layer4_outputs(10027) <= not b;
    layer4_outputs(10028) <= not a or b;
    layer4_outputs(10029) <= not b;
    layer4_outputs(10030) <= not b;
    layer4_outputs(10031) <= not (a or b);
    layer4_outputs(10032) <= not (a or b);
    layer4_outputs(10033) <= a or b;
    layer4_outputs(10034) <= not a or b;
    layer4_outputs(10035) <= a xor b;
    layer4_outputs(10036) <= not (a or b);
    layer4_outputs(10037) <= a;
    layer4_outputs(10038) <= not a;
    layer4_outputs(10039) <= b;
    layer4_outputs(10040) <= a and b;
    layer4_outputs(10041) <= b and not a;
    layer4_outputs(10042) <= a;
    layer4_outputs(10043) <= not b or a;
    layer4_outputs(10044) <= not b;
    layer4_outputs(10045) <= not b;
    layer4_outputs(10046) <= not a;
    layer4_outputs(10047) <= not (a and b);
    layer4_outputs(10048) <= a and not b;
    layer4_outputs(10049) <= not b;
    layer4_outputs(10050) <= not a;
    layer4_outputs(10051) <= b;
    layer4_outputs(10052) <= a or b;
    layer4_outputs(10053) <= not b;
    layer4_outputs(10054) <= not b;
    layer4_outputs(10055) <= not (a or b);
    layer4_outputs(10056) <= b;
    layer4_outputs(10057) <= b and not a;
    layer4_outputs(10058) <= a and not b;
    layer4_outputs(10059) <= not b;
    layer4_outputs(10060) <= not b;
    layer4_outputs(10061) <= a and b;
    layer4_outputs(10062) <= not b or a;
    layer4_outputs(10063) <= not b;
    layer4_outputs(10064) <= b;
    layer4_outputs(10065) <= not b;
    layer4_outputs(10066) <= b and not a;
    layer4_outputs(10067) <= not a;
    layer4_outputs(10068) <= b;
    layer4_outputs(10069) <= a;
    layer4_outputs(10070) <= a and b;
    layer4_outputs(10071) <= a or b;
    layer4_outputs(10072) <= not a;
    layer4_outputs(10073) <= not (a and b);
    layer4_outputs(10074) <= not a;
    layer4_outputs(10075) <= not b;
    layer4_outputs(10076) <= not b;
    layer4_outputs(10077) <= not a or b;
    layer4_outputs(10078) <= not (a and b);
    layer4_outputs(10079) <= b;
    layer4_outputs(10080) <= '1';
    layer4_outputs(10081) <= not b;
    layer4_outputs(10082) <= a xor b;
    layer4_outputs(10083) <= a;
    layer4_outputs(10084) <= b and not a;
    layer4_outputs(10085) <= b;
    layer4_outputs(10086) <= not a;
    layer4_outputs(10087) <= b;
    layer4_outputs(10088) <= a or b;
    layer4_outputs(10089) <= not b;
    layer4_outputs(10090) <= not a;
    layer4_outputs(10091) <= a;
    layer4_outputs(10092) <= not (a or b);
    layer4_outputs(10093) <= a;
    layer4_outputs(10094) <= not b or a;
    layer4_outputs(10095) <= not a;
    layer4_outputs(10096) <= a and not b;
    layer4_outputs(10097) <= not a or b;
    layer4_outputs(10098) <= a and b;
    layer4_outputs(10099) <= a or b;
    layer4_outputs(10100) <= not a or b;
    layer4_outputs(10101) <= a;
    layer4_outputs(10102) <= '1';
    layer4_outputs(10103) <= not a;
    layer4_outputs(10104) <= a or b;
    layer4_outputs(10105) <= b;
    layer4_outputs(10106) <= not (a and b);
    layer4_outputs(10107) <= not (a or b);
    layer4_outputs(10108) <= '1';
    layer4_outputs(10109) <= a;
    layer4_outputs(10110) <= b;
    layer4_outputs(10111) <= a and not b;
    layer4_outputs(10112) <= a;
    layer4_outputs(10113) <= not a;
    layer4_outputs(10114) <= a xor b;
    layer4_outputs(10115) <= b;
    layer4_outputs(10116) <= not b;
    layer4_outputs(10117) <= not a or b;
    layer4_outputs(10118) <= a or b;
    layer4_outputs(10119) <= a and b;
    layer4_outputs(10120) <= not a;
    layer4_outputs(10121) <= not (a or b);
    layer4_outputs(10122) <= b;
    layer4_outputs(10123) <= not b;
    layer4_outputs(10124) <= not b or a;
    layer4_outputs(10125) <= b;
    layer4_outputs(10126) <= not a;
    layer4_outputs(10127) <= not (a and b);
    layer4_outputs(10128) <= not b;
    layer4_outputs(10129) <= not b or a;
    layer4_outputs(10130) <= a;
    layer4_outputs(10131) <= a xor b;
    layer4_outputs(10132) <= a;
    layer4_outputs(10133) <= a xor b;
    layer4_outputs(10134) <= b;
    layer4_outputs(10135) <= not a;
    layer4_outputs(10136) <= b;
    layer4_outputs(10137) <= a xor b;
    layer4_outputs(10138) <= not a;
    layer4_outputs(10139) <= a and not b;
    layer4_outputs(10140) <= not (a and b);
    layer4_outputs(10141) <= not (a or b);
    layer4_outputs(10142) <= not (a and b);
    layer4_outputs(10143) <= not b;
    layer4_outputs(10144) <= b and not a;
    layer4_outputs(10145) <= not b or a;
    layer4_outputs(10146) <= b;
    layer4_outputs(10147) <= not b;
    layer4_outputs(10148) <= a xor b;
    layer4_outputs(10149) <= a;
    layer4_outputs(10150) <= b and not a;
    layer4_outputs(10151) <= not (a xor b);
    layer4_outputs(10152) <= a and b;
    layer4_outputs(10153) <= a and not b;
    layer4_outputs(10154) <= a and b;
    layer4_outputs(10155) <= not b;
    layer4_outputs(10156) <= a and b;
    layer4_outputs(10157) <= '1';
    layer4_outputs(10158) <= not a or b;
    layer4_outputs(10159) <= not b;
    layer4_outputs(10160) <= a;
    layer4_outputs(10161) <= not a or b;
    layer4_outputs(10162) <= b and not a;
    layer4_outputs(10163) <= not b;
    layer4_outputs(10164) <= a or b;
    layer4_outputs(10165) <= not b;
    layer4_outputs(10166) <= not a or b;
    layer4_outputs(10167) <= not (a and b);
    layer4_outputs(10168) <= b;
    layer4_outputs(10169) <= not a;
    layer4_outputs(10170) <= not b;
    layer4_outputs(10171) <= not b or a;
    layer4_outputs(10172) <= not b;
    layer4_outputs(10173) <= not b or a;
    layer4_outputs(10174) <= not b;
    layer4_outputs(10175) <= a;
    layer4_outputs(10176) <= b;
    layer4_outputs(10177) <= a;
    layer4_outputs(10178) <= a xor b;
    layer4_outputs(10179) <= not a;
    layer4_outputs(10180) <= a and not b;
    layer4_outputs(10181) <= b;
    layer4_outputs(10182) <= b;
    layer4_outputs(10183) <= not a;
    layer4_outputs(10184) <= not (a and b);
    layer4_outputs(10185) <= not (a xor b);
    layer4_outputs(10186) <= not b;
    layer4_outputs(10187) <= not (a xor b);
    layer4_outputs(10188) <= a;
    layer4_outputs(10189) <= a;
    layer4_outputs(10190) <= not b;
    layer4_outputs(10191) <= b;
    layer4_outputs(10192) <= not b;
    layer4_outputs(10193) <= a and not b;
    layer4_outputs(10194) <= not (a xor b);
    layer4_outputs(10195) <= not (a or b);
    layer4_outputs(10196) <= b;
    layer4_outputs(10197) <= a;
    layer4_outputs(10198) <= not a or b;
    layer4_outputs(10199) <= a or b;
    layer4_outputs(10200) <= '1';
    layer4_outputs(10201) <= a xor b;
    layer4_outputs(10202) <= a;
    layer4_outputs(10203) <= b;
    layer4_outputs(10204) <= not a;
    layer4_outputs(10205) <= not (a xor b);
    layer4_outputs(10206) <= not (a xor b);
    layer4_outputs(10207) <= not b or a;
    layer4_outputs(10208) <= a or b;
    layer4_outputs(10209) <= '1';
    layer4_outputs(10210) <= a;
    layer4_outputs(10211) <= a xor b;
    layer4_outputs(10212) <= a and b;
    layer4_outputs(10213) <= a;
    layer4_outputs(10214) <= not a or b;
    layer4_outputs(10215) <= a and not b;
    layer4_outputs(10216) <= a and b;
    layer4_outputs(10217) <= a or b;
    layer4_outputs(10218) <= b and not a;
    layer4_outputs(10219) <= a;
    layer4_outputs(10220) <= a xor b;
    layer4_outputs(10221) <= a or b;
    layer4_outputs(10222) <= a;
    layer4_outputs(10223) <= not (a xor b);
    layer4_outputs(10224) <= a;
    layer4_outputs(10225) <= not b or a;
    layer4_outputs(10226) <= a or b;
    layer4_outputs(10227) <= a;
    layer4_outputs(10228) <= not a or b;
    layer4_outputs(10229) <= a and b;
    layer4_outputs(10230) <= not a;
    layer4_outputs(10231) <= b;
    layer4_outputs(10232) <= not (a xor b);
    layer4_outputs(10233) <= not b or a;
    layer4_outputs(10234) <= not a;
    layer4_outputs(10235) <= not a or b;
    layer4_outputs(10236) <= not b;
    layer4_outputs(10237) <= a and not b;
    layer4_outputs(10238) <= '0';
    layer4_outputs(10239) <= not b;
    layer4_outputs(10240) <= not b;
    layer4_outputs(10241) <= b and not a;
    layer4_outputs(10242) <= not a;
    layer4_outputs(10243) <= not a or b;
    layer4_outputs(10244) <= b and not a;
    layer4_outputs(10245) <= not a;
    layer4_outputs(10246) <= not (a or b);
    layer4_outputs(10247) <= b;
    layer4_outputs(10248) <= a and not b;
    layer4_outputs(10249) <= a;
    layer4_outputs(10250) <= b and not a;
    layer4_outputs(10251) <= a or b;
    layer4_outputs(10252) <= not (a or b);
    layer4_outputs(10253) <= not a;
    layer4_outputs(10254) <= not a or b;
    layer4_outputs(10255) <= b and not a;
    layer4_outputs(10256) <= a;
    layer4_outputs(10257) <= b and not a;
    layer4_outputs(10258) <= not (a and b);
    layer4_outputs(10259) <= not (a and b);
    layer4_outputs(10260) <= b;
    layer4_outputs(10261) <= a and b;
    layer4_outputs(10262) <= a or b;
    layer4_outputs(10263) <= a and not b;
    layer4_outputs(10264) <= a and b;
    layer4_outputs(10265) <= a and not b;
    layer4_outputs(10266) <= not b or a;
    layer4_outputs(10267) <= '1';
    layer4_outputs(10268) <= not b;
    layer4_outputs(10269) <= a;
    layer4_outputs(10270) <= '0';
    layer4_outputs(10271) <= a and b;
    layer4_outputs(10272) <= not b;
    layer4_outputs(10273) <= not a or b;
    layer4_outputs(10274) <= a xor b;
    layer4_outputs(10275) <= not a;
    layer4_outputs(10276) <= not b;
    layer4_outputs(10277) <= a;
    layer4_outputs(10278) <= not a;
    layer4_outputs(10279) <= a;
    layer4_outputs(10280) <= a xor b;
    layer4_outputs(10281) <= a;
    layer4_outputs(10282) <= a xor b;
    layer4_outputs(10283) <= '0';
    layer4_outputs(10284) <= not (a xor b);
    layer4_outputs(10285) <= a;
    layer4_outputs(10286) <= a or b;
    layer4_outputs(10287) <= not b or a;
    layer4_outputs(10288) <= b;
    layer4_outputs(10289) <= a;
    layer4_outputs(10290) <= not b;
    layer4_outputs(10291) <= not a;
    layer4_outputs(10292) <= a;
    layer4_outputs(10293) <= a xor b;
    layer4_outputs(10294) <= a or b;
    layer4_outputs(10295) <= b;
    layer4_outputs(10296) <= a or b;
    layer4_outputs(10297) <= not b;
    layer4_outputs(10298) <= not a;
    layer4_outputs(10299) <= not (a or b);
    layer4_outputs(10300) <= not a;
    layer4_outputs(10301) <= b;
    layer4_outputs(10302) <= not b;
    layer4_outputs(10303) <= not (a and b);
    layer4_outputs(10304) <= b;
    layer4_outputs(10305) <= not b;
    layer4_outputs(10306) <= a;
    layer4_outputs(10307) <= not a or b;
    layer4_outputs(10308) <= a;
    layer4_outputs(10309) <= not b or a;
    layer4_outputs(10310) <= not (a or b);
    layer4_outputs(10311) <= '0';
    layer4_outputs(10312) <= a or b;
    layer4_outputs(10313) <= not (a and b);
    layer4_outputs(10314) <= a and not b;
    layer4_outputs(10315) <= not a or b;
    layer4_outputs(10316) <= not a;
    layer4_outputs(10317) <= not a or b;
    layer4_outputs(10318) <= b and not a;
    layer4_outputs(10319) <= '0';
    layer4_outputs(10320) <= not a or b;
    layer4_outputs(10321) <= b and not a;
    layer4_outputs(10322) <= b;
    layer4_outputs(10323) <= not a or b;
    layer4_outputs(10324) <= b;
    layer4_outputs(10325) <= not (a and b);
    layer4_outputs(10326) <= not b;
    layer4_outputs(10327) <= not (a or b);
    layer4_outputs(10328) <= a and b;
    layer4_outputs(10329) <= b;
    layer4_outputs(10330) <= not (a xor b);
    layer4_outputs(10331) <= not a or b;
    layer4_outputs(10332) <= a and not b;
    layer4_outputs(10333) <= not a;
    layer4_outputs(10334) <= '1';
    layer4_outputs(10335) <= not b;
    layer4_outputs(10336) <= a xor b;
    layer4_outputs(10337) <= not b;
    layer4_outputs(10338) <= not a or b;
    layer4_outputs(10339) <= not a;
    layer4_outputs(10340) <= a or b;
    layer4_outputs(10341) <= not (a and b);
    layer4_outputs(10342) <= not b;
    layer4_outputs(10343) <= a or b;
    layer4_outputs(10344) <= not (a and b);
    layer4_outputs(10345) <= not (a xor b);
    layer4_outputs(10346) <= a and b;
    layer4_outputs(10347) <= not (a and b);
    layer4_outputs(10348) <= a and b;
    layer4_outputs(10349) <= b and not a;
    layer4_outputs(10350) <= a and not b;
    layer4_outputs(10351) <= not (a or b);
    layer4_outputs(10352) <= '1';
    layer4_outputs(10353) <= not b or a;
    layer4_outputs(10354) <= b;
    layer4_outputs(10355) <= a and b;
    layer4_outputs(10356) <= not a or b;
    layer4_outputs(10357) <= not b or a;
    layer4_outputs(10358) <= b;
    layer4_outputs(10359) <= a or b;
    layer4_outputs(10360) <= b;
    layer4_outputs(10361) <= b and not a;
    layer4_outputs(10362) <= not a;
    layer4_outputs(10363) <= a;
    layer4_outputs(10364) <= a and b;
    layer4_outputs(10365) <= a;
    layer4_outputs(10366) <= not b;
    layer4_outputs(10367) <= a;
    layer4_outputs(10368) <= not (a xor b);
    layer4_outputs(10369) <= a;
    layer4_outputs(10370) <= a;
    layer4_outputs(10371) <= b;
    layer4_outputs(10372) <= a and b;
    layer4_outputs(10373) <= not (a and b);
    layer4_outputs(10374) <= not (a and b);
    layer4_outputs(10375) <= a and b;
    layer4_outputs(10376) <= a and not b;
    layer4_outputs(10377) <= not (a or b);
    layer4_outputs(10378) <= a and b;
    layer4_outputs(10379) <= '0';
    layer4_outputs(10380) <= not b;
    layer4_outputs(10381) <= b;
    layer4_outputs(10382) <= a;
    layer4_outputs(10383) <= a and not b;
    layer4_outputs(10384) <= not (a and b);
    layer4_outputs(10385) <= b and not a;
    layer4_outputs(10386) <= a;
    layer4_outputs(10387) <= not b;
    layer4_outputs(10388) <= a;
    layer4_outputs(10389) <= not a or b;
    layer4_outputs(10390) <= a xor b;
    layer4_outputs(10391) <= a;
    layer4_outputs(10392) <= not b;
    layer4_outputs(10393) <= not a;
    layer4_outputs(10394) <= not a;
    layer4_outputs(10395) <= not b or a;
    layer4_outputs(10396) <= not b;
    layer4_outputs(10397) <= not a or b;
    layer4_outputs(10398) <= b and not a;
    layer4_outputs(10399) <= a and b;
    layer4_outputs(10400) <= a or b;
    layer4_outputs(10401) <= '0';
    layer4_outputs(10402) <= not b;
    layer4_outputs(10403) <= b;
    layer4_outputs(10404) <= not b or a;
    layer4_outputs(10405) <= '0';
    layer4_outputs(10406) <= '0';
    layer4_outputs(10407) <= not (a or b);
    layer4_outputs(10408) <= not b;
    layer4_outputs(10409) <= a;
    layer4_outputs(10410) <= not (a and b);
    layer4_outputs(10411) <= a xor b;
    layer4_outputs(10412) <= a and not b;
    layer4_outputs(10413) <= not b or a;
    layer4_outputs(10414) <= '1';
    layer4_outputs(10415) <= b and not a;
    layer4_outputs(10416) <= not a or b;
    layer4_outputs(10417) <= not a;
    layer4_outputs(10418) <= b and not a;
    layer4_outputs(10419) <= not (a or b);
    layer4_outputs(10420) <= not b or a;
    layer4_outputs(10421) <= not (a and b);
    layer4_outputs(10422) <= not a;
    layer4_outputs(10423) <= b;
    layer4_outputs(10424) <= not (a or b);
    layer4_outputs(10425) <= b;
    layer4_outputs(10426) <= not (a xor b);
    layer4_outputs(10427) <= a and b;
    layer4_outputs(10428) <= a xor b;
    layer4_outputs(10429) <= a;
    layer4_outputs(10430) <= not a;
    layer4_outputs(10431) <= a or b;
    layer4_outputs(10432) <= b;
    layer4_outputs(10433) <= '0';
    layer4_outputs(10434) <= not a or b;
    layer4_outputs(10435) <= not b;
    layer4_outputs(10436) <= a and b;
    layer4_outputs(10437) <= not a;
    layer4_outputs(10438) <= a and not b;
    layer4_outputs(10439) <= a;
    layer4_outputs(10440) <= not b;
    layer4_outputs(10441) <= not b;
    layer4_outputs(10442) <= not a;
    layer4_outputs(10443) <= b and not a;
    layer4_outputs(10444) <= b;
    layer4_outputs(10445) <= '0';
    layer4_outputs(10446) <= a xor b;
    layer4_outputs(10447) <= a;
    layer4_outputs(10448) <= a xor b;
    layer4_outputs(10449) <= b and not a;
    layer4_outputs(10450) <= not (a or b);
    layer4_outputs(10451) <= a or b;
    layer4_outputs(10452) <= not b;
    layer4_outputs(10453) <= not b;
    layer4_outputs(10454) <= not a;
    layer4_outputs(10455) <= not a;
    layer4_outputs(10456) <= b;
    layer4_outputs(10457) <= not (a xor b);
    layer4_outputs(10458) <= a xor b;
    layer4_outputs(10459) <= a;
    layer4_outputs(10460) <= a or b;
    layer4_outputs(10461) <= a;
    layer4_outputs(10462) <= not b;
    layer4_outputs(10463) <= not a or b;
    layer4_outputs(10464) <= not a;
    layer4_outputs(10465) <= a and b;
    layer4_outputs(10466) <= b and not a;
    layer4_outputs(10467) <= not b;
    layer4_outputs(10468) <= not a or b;
    layer4_outputs(10469) <= b and not a;
    layer4_outputs(10470) <= '1';
    layer4_outputs(10471) <= b and not a;
    layer4_outputs(10472) <= not (a or b);
    layer4_outputs(10473) <= a;
    layer4_outputs(10474) <= not b or a;
    layer4_outputs(10475) <= a;
    layer4_outputs(10476) <= not (a or b);
    layer4_outputs(10477) <= b;
    layer4_outputs(10478) <= not (a or b);
    layer4_outputs(10479) <= not a;
    layer4_outputs(10480) <= not a;
    layer4_outputs(10481) <= not a;
    layer4_outputs(10482) <= not b;
    layer4_outputs(10483) <= not (a and b);
    layer4_outputs(10484) <= a and b;
    layer4_outputs(10485) <= not (a or b);
    layer4_outputs(10486) <= b;
    layer4_outputs(10487) <= a;
    layer4_outputs(10488) <= not a or b;
    layer4_outputs(10489) <= '0';
    layer4_outputs(10490) <= b and not a;
    layer4_outputs(10491) <= a;
    layer4_outputs(10492) <= b;
    layer4_outputs(10493) <= b;
    layer4_outputs(10494) <= not (a and b);
    layer4_outputs(10495) <= '1';
    layer4_outputs(10496) <= a and not b;
    layer4_outputs(10497) <= not (a and b);
    layer4_outputs(10498) <= b and not a;
    layer4_outputs(10499) <= not a or b;
    layer4_outputs(10500) <= b;
    layer4_outputs(10501) <= not a;
    layer4_outputs(10502) <= a;
    layer4_outputs(10503) <= b;
    layer4_outputs(10504) <= not a or b;
    layer4_outputs(10505) <= b;
    layer4_outputs(10506) <= not (a or b);
    layer4_outputs(10507) <= not (a and b);
    layer4_outputs(10508) <= a xor b;
    layer4_outputs(10509) <= '1';
    layer4_outputs(10510) <= not a;
    layer4_outputs(10511) <= not (a and b);
    layer4_outputs(10512) <= b;
    layer4_outputs(10513) <= not b;
    layer4_outputs(10514) <= a and b;
    layer4_outputs(10515) <= a xor b;
    layer4_outputs(10516) <= b;
    layer4_outputs(10517) <= not b;
    layer4_outputs(10518) <= not b;
    layer4_outputs(10519) <= b;
    layer4_outputs(10520) <= b and not a;
    layer4_outputs(10521) <= not a or b;
    layer4_outputs(10522) <= not (a and b);
    layer4_outputs(10523) <= not b or a;
    layer4_outputs(10524) <= not a;
    layer4_outputs(10525) <= not (a and b);
    layer4_outputs(10526) <= not (a and b);
    layer4_outputs(10527) <= b and not a;
    layer4_outputs(10528) <= not (a or b);
    layer4_outputs(10529) <= not b;
    layer4_outputs(10530) <= a xor b;
    layer4_outputs(10531) <= a;
    layer4_outputs(10532) <= not (a xor b);
    layer4_outputs(10533) <= b;
    layer4_outputs(10534) <= not (a or b);
    layer4_outputs(10535) <= not b or a;
    layer4_outputs(10536) <= not (a or b);
    layer4_outputs(10537) <= a;
    layer4_outputs(10538) <= not a;
    layer4_outputs(10539) <= a;
    layer4_outputs(10540) <= a xor b;
    layer4_outputs(10541) <= a and not b;
    layer4_outputs(10542) <= a and not b;
    layer4_outputs(10543) <= a;
    layer4_outputs(10544) <= not a or b;
    layer4_outputs(10545) <= a and b;
    layer4_outputs(10546) <= not b;
    layer4_outputs(10547) <= not (a or b);
    layer4_outputs(10548) <= a or b;
    layer4_outputs(10549) <= not b;
    layer4_outputs(10550) <= a xor b;
    layer4_outputs(10551) <= not (a xor b);
    layer4_outputs(10552) <= a or b;
    layer4_outputs(10553) <= a xor b;
    layer4_outputs(10554) <= a and not b;
    layer4_outputs(10555) <= b and not a;
    layer4_outputs(10556) <= a;
    layer4_outputs(10557) <= not a;
    layer4_outputs(10558) <= a and b;
    layer4_outputs(10559) <= a and not b;
    layer4_outputs(10560) <= a and not b;
    layer4_outputs(10561) <= not (a or b);
    layer4_outputs(10562) <= not b or a;
    layer4_outputs(10563) <= a and b;
    layer4_outputs(10564) <= not (a or b);
    layer4_outputs(10565) <= not a;
    layer4_outputs(10566) <= a or b;
    layer4_outputs(10567) <= a or b;
    layer4_outputs(10568) <= not a;
    layer4_outputs(10569) <= not a;
    layer4_outputs(10570) <= a;
    layer4_outputs(10571) <= a or b;
    layer4_outputs(10572) <= not b;
    layer4_outputs(10573) <= b;
    layer4_outputs(10574) <= b and not a;
    layer4_outputs(10575) <= not a;
    layer4_outputs(10576) <= a and not b;
    layer4_outputs(10577) <= a or b;
    layer4_outputs(10578) <= not b;
    layer4_outputs(10579) <= not b;
    layer4_outputs(10580) <= a;
    layer4_outputs(10581) <= not b;
    layer4_outputs(10582) <= not a;
    layer4_outputs(10583) <= not (a xor b);
    layer4_outputs(10584) <= a or b;
    layer4_outputs(10585) <= not (a xor b);
    layer4_outputs(10586) <= a;
    layer4_outputs(10587) <= b;
    layer4_outputs(10588) <= not a;
    layer4_outputs(10589) <= not (a and b);
    layer4_outputs(10590) <= b and not a;
    layer4_outputs(10591) <= a or b;
    layer4_outputs(10592) <= a;
    layer4_outputs(10593) <= a and b;
    layer4_outputs(10594) <= not b;
    layer4_outputs(10595) <= a and not b;
    layer4_outputs(10596) <= not a;
    layer4_outputs(10597) <= not b or a;
    layer4_outputs(10598) <= not (a xor b);
    layer4_outputs(10599) <= not b;
    layer4_outputs(10600) <= not b;
    layer4_outputs(10601) <= b;
    layer4_outputs(10602) <= not (a or b);
    layer4_outputs(10603) <= b;
    layer4_outputs(10604) <= not (a or b);
    layer4_outputs(10605) <= not (a and b);
    layer4_outputs(10606) <= a or b;
    layer4_outputs(10607) <= not b;
    layer4_outputs(10608) <= a and b;
    layer4_outputs(10609) <= b;
    layer4_outputs(10610) <= '0';
    layer4_outputs(10611) <= not b;
    layer4_outputs(10612) <= '0';
    layer4_outputs(10613) <= not (a and b);
    layer4_outputs(10614) <= a xor b;
    layer4_outputs(10615) <= not b;
    layer4_outputs(10616) <= a;
    layer4_outputs(10617) <= not a;
    layer4_outputs(10618) <= a xor b;
    layer4_outputs(10619) <= not b;
    layer4_outputs(10620) <= not b;
    layer4_outputs(10621) <= not b;
    layer4_outputs(10622) <= not b;
    layer4_outputs(10623) <= b;
    layer4_outputs(10624) <= not a or b;
    layer4_outputs(10625) <= a;
    layer4_outputs(10626) <= not (a and b);
    layer4_outputs(10627) <= not a;
    layer4_outputs(10628) <= not a;
    layer4_outputs(10629) <= not a;
    layer4_outputs(10630) <= not (a or b);
    layer4_outputs(10631) <= not b;
    layer4_outputs(10632) <= b;
    layer4_outputs(10633) <= not a or b;
    layer4_outputs(10634) <= not b;
    layer4_outputs(10635) <= not b;
    layer4_outputs(10636) <= not b;
    layer4_outputs(10637) <= a and not b;
    layer4_outputs(10638) <= a xor b;
    layer4_outputs(10639) <= not b;
    layer4_outputs(10640) <= not a or b;
    layer4_outputs(10641) <= b;
    layer4_outputs(10642) <= a and b;
    layer4_outputs(10643) <= not (a xor b);
    layer4_outputs(10644) <= b;
    layer4_outputs(10645) <= not a or b;
    layer4_outputs(10646) <= a or b;
    layer4_outputs(10647) <= a;
    layer4_outputs(10648) <= a;
    layer4_outputs(10649) <= not a or b;
    layer4_outputs(10650) <= not a;
    layer4_outputs(10651) <= a xor b;
    layer4_outputs(10652) <= a or b;
    layer4_outputs(10653) <= b;
    layer4_outputs(10654) <= not b;
    layer4_outputs(10655) <= not a;
    layer4_outputs(10656) <= not (a or b);
    layer4_outputs(10657) <= not b;
    layer4_outputs(10658) <= not (a or b);
    layer4_outputs(10659) <= not a;
    layer4_outputs(10660) <= a;
    layer4_outputs(10661) <= a and b;
    layer4_outputs(10662) <= b;
    layer4_outputs(10663) <= not a;
    layer4_outputs(10664) <= a and not b;
    layer4_outputs(10665) <= a xor b;
    layer4_outputs(10666) <= a or b;
    layer4_outputs(10667) <= a;
    layer4_outputs(10668) <= a and b;
    layer4_outputs(10669) <= b and not a;
    layer4_outputs(10670) <= not a;
    layer4_outputs(10671) <= b and not a;
    layer4_outputs(10672) <= not b;
    layer4_outputs(10673) <= not (a or b);
    layer4_outputs(10674) <= '0';
    layer4_outputs(10675) <= not a;
    layer4_outputs(10676) <= not b;
    layer4_outputs(10677) <= a and not b;
    layer4_outputs(10678) <= b;
    layer4_outputs(10679) <= a and b;
    layer4_outputs(10680) <= a;
    layer4_outputs(10681) <= not a or b;
    layer4_outputs(10682) <= not b;
    layer4_outputs(10683) <= b;
    layer4_outputs(10684) <= not a or b;
    layer4_outputs(10685) <= not (a and b);
    layer4_outputs(10686) <= not a or b;
    layer4_outputs(10687) <= '0';
    layer4_outputs(10688) <= a and b;
    layer4_outputs(10689) <= a and b;
    layer4_outputs(10690) <= a and not b;
    layer4_outputs(10691) <= not a;
    layer4_outputs(10692) <= not a;
    layer4_outputs(10693) <= not (a or b);
    layer4_outputs(10694) <= b and not a;
    layer4_outputs(10695) <= not (a xor b);
    layer4_outputs(10696) <= not a;
    layer4_outputs(10697) <= not b;
    layer4_outputs(10698) <= a xor b;
    layer4_outputs(10699) <= not (a xor b);
    layer4_outputs(10700) <= a xor b;
    layer4_outputs(10701) <= not (a and b);
    layer4_outputs(10702) <= a and b;
    layer4_outputs(10703) <= a and not b;
    layer4_outputs(10704) <= not (a and b);
    layer4_outputs(10705) <= a xor b;
    layer4_outputs(10706) <= a or b;
    layer4_outputs(10707) <= not (a or b);
    layer4_outputs(10708) <= '1';
    layer4_outputs(10709) <= not (a xor b);
    layer4_outputs(10710) <= not (a or b);
    layer4_outputs(10711) <= not a;
    layer4_outputs(10712) <= a and not b;
    layer4_outputs(10713) <= a and not b;
    layer4_outputs(10714) <= a or b;
    layer4_outputs(10715) <= not b;
    layer4_outputs(10716) <= not (a and b);
    layer4_outputs(10717) <= not b or a;
    layer4_outputs(10718) <= a;
    layer4_outputs(10719) <= a and not b;
    layer4_outputs(10720) <= not b or a;
    layer4_outputs(10721) <= b;
    layer4_outputs(10722) <= not a;
    layer4_outputs(10723) <= b and not a;
    layer4_outputs(10724) <= not (a or b);
    layer4_outputs(10725) <= not a;
    layer4_outputs(10726) <= not b or a;
    layer4_outputs(10727) <= not a or b;
    layer4_outputs(10728) <= not (a or b);
    layer4_outputs(10729) <= not (a or b);
    layer4_outputs(10730) <= not (a xor b);
    layer4_outputs(10731) <= not (a or b);
    layer4_outputs(10732) <= a xor b;
    layer4_outputs(10733) <= not (a and b);
    layer4_outputs(10734) <= a or b;
    layer4_outputs(10735) <= a xor b;
    layer4_outputs(10736) <= not (a and b);
    layer4_outputs(10737) <= not (a or b);
    layer4_outputs(10738) <= a;
    layer4_outputs(10739) <= a xor b;
    layer4_outputs(10740) <= b;
    layer4_outputs(10741) <= '0';
    layer4_outputs(10742) <= '0';
    layer4_outputs(10743) <= a;
    layer4_outputs(10744) <= not b;
    layer4_outputs(10745) <= not a;
    layer4_outputs(10746) <= b and not a;
    layer4_outputs(10747) <= a xor b;
    layer4_outputs(10748) <= b and not a;
    layer4_outputs(10749) <= a and not b;
    layer4_outputs(10750) <= not (a and b);
    layer4_outputs(10751) <= not (a and b);
    layer4_outputs(10752) <= not (a xor b);
    layer4_outputs(10753) <= a xor b;
    layer4_outputs(10754) <= '0';
    layer4_outputs(10755) <= a or b;
    layer4_outputs(10756) <= a;
    layer4_outputs(10757) <= not a;
    layer4_outputs(10758) <= not a or b;
    layer4_outputs(10759) <= a;
    layer4_outputs(10760) <= b;
    layer4_outputs(10761) <= a or b;
    layer4_outputs(10762) <= not b;
    layer4_outputs(10763) <= not (a xor b);
    layer4_outputs(10764) <= a and not b;
    layer4_outputs(10765) <= not b or a;
    layer4_outputs(10766) <= a and b;
    layer4_outputs(10767) <= b and not a;
    layer4_outputs(10768) <= not b;
    layer4_outputs(10769) <= b;
    layer4_outputs(10770) <= not b;
    layer4_outputs(10771) <= not a or b;
    layer4_outputs(10772) <= not a or b;
    layer4_outputs(10773) <= a;
    layer4_outputs(10774) <= not a;
    layer4_outputs(10775) <= b;
    layer4_outputs(10776) <= not b;
    layer4_outputs(10777) <= not a;
    layer4_outputs(10778) <= not a or b;
    layer4_outputs(10779) <= b and not a;
    layer4_outputs(10780) <= not (a xor b);
    layer4_outputs(10781) <= b and not a;
    layer4_outputs(10782) <= a xor b;
    layer4_outputs(10783) <= not b;
    layer4_outputs(10784) <= b;
    layer4_outputs(10785) <= a and not b;
    layer4_outputs(10786) <= not (a xor b);
    layer4_outputs(10787) <= not a or b;
    layer4_outputs(10788) <= b;
    layer4_outputs(10789) <= not a;
    layer4_outputs(10790) <= a;
    layer4_outputs(10791) <= not (a xor b);
    layer4_outputs(10792) <= a xor b;
    layer4_outputs(10793) <= a and not b;
    layer4_outputs(10794) <= not a;
    layer4_outputs(10795) <= b;
    layer4_outputs(10796) <= not a or b;
    layer4_outputs(10797) <= a;
    layer4_outputs(10798) <= not a;
    layer4_outputs(10799) <= not b;
    layer4_outputs(10800) <= not a;
    layer4_outputs(10801) <= a xor b;
    layer4_outputs(10802) <= a and b;
    layer4_outputs(10803) <= a and b;
    layer4_outputs(10804) <= a or b;
    layer4_outputs(10805) <= a;
    layer4_outputs(10806) <= not a;
    layer4_outputs(10807) <= not (a and b);
    layer4_outputs(10808) <= not (a or b);
    layer4_outputs(10809) <= not a;
    layer4_outputs(10810) <= b;
    layer4_outputs(10811) <= not b;
    layer4_outputs(10812) <= not b;
    layer4_outputs(10813) <= a;
    layer4_outputs(10814) <= not b or a;
    layer4_outputs(10815) <= '0';
    layer4_outputs(10816) <= b;
    layer4_outputs(10817) <= a or b;
    layer4_outputs(10818) <= a;
    layer4_outputs(10819) <= b;
    layer4_outputs(10820) <= not a;
    layer4_outputs(10821) <= a xor b;
    layer4_outputs(10822) <= not a or b;
    layer4_outputs(10823) <= not (a xor b);
    layer4_outputs(10824) <= not b;
    layer4_outputs(10825) <= a;
    layer4_outputs(10826) <= a;
    layer4_outputs(10827) <= not b;
    layer4_outputs(10828) <= not b;
    layer4_outputs(10829) <= a and not b;
    layer4_outputs(10830) <= not b or a;
    layer4_outputs(10831) <= not (a xor b);
    layer4_outputs(10832) <= not b;
    layer4_outputs(10833) <= a xor b;
    layer4_outputs(10834) <= b;
    layer4_outputs(10835) <= not (a and b);
    layer4_outputs(10836) <= a and not b;
    layer4_outputs(10837) <= a and not b;
    layer4_outputs(10838) <= not (a or b);
    layer4_outputs(10839) <= a or b;
    layer4_outputs(10840) <= not a or b;
    layer4_outputs(10841) <= a or b;
    layer4_outputs(10842) <= not (a or b);
    layer4_outputs(10843) <= not a;
    layer4_outputs(10844) <= a;
    layer4_outputs(10845) <= not a;
    layer4_outputs(10846) <= a and not b;
    layer4_outputs(10847) <= not b or a;
    layer4_outputs(10848) <= b;
    layer4_outputs(10849) <= '0';
    layer4_outputs(10850) <= a or b;
    layer4_outputs(10851) <= a or b;
    layer4_outputs(10852) <= not b or a;
    layer4_outputs(10853) <= not a;
    layer4_outputs(10854) <= not b;
    layer4_outputs(10855) <= a and not b;
    layer4_outputs(10856) <= not (a and b);
    layer4_outputs(10857) <= b and not a;
    layer4_outputs(10858) <= a and b;
    layer4_outputs(10859) <= not (a and b);
    layer4_outputs(10860) <= not a;
    layer4_outputs(10861) <= not (a and b);
    layer4_outputs(10862) <= not b;
    layer4_outputs(10863) <= not a;
    layer4_outputs(10864) <= not a;
    layer4_outputs(10865) <= not b;
    layer4_outputs(10866) <= not b or a;
    layer4_outputs(10867) <= '1';
    layer4_outputs(10868) <= '0';
    layer4_outputs(10869) <= a and b;
    layer4_outputs(10870) <= a or b;
    layer4_outputs(10871) <= a and b;
    layer4_outputs(10872) <= not a;
    layer4_outputs(10873) <= a or b;
    layer4_outputs(10874) <= b;
    layer4_outputs(10875) <= not a;
    layer4_outputs(10876) <= not (a xor b);
    layer4_outputs(10877) <= a xor b;
    layer4_outputs(10878) <= a xor b;
    layer4_outputs(10879) <= a xor b;
    layer4_outputs(10880) <= not a or b;
    layer4_outputs(10881) <= a and not b;
    layer4_outputs(10882) <= not b or a;
    layer4_outputs(10883) <= a;
    layer4_outputs(10884) <= a and not b;
    layer4_outputs(10885) <= a and b;
    layer4_outputs(10886) <= b and not a;
    layer4_outputs(10887) <= a and not b;
    layer4_outputs(10888) <= b;
    layer4_outputs(10889) <= not a;
    layer4_outputs(10890) <= not b;
    layer4_outputs(10891) <= a;
    layer4_outputs(10892) <= a xor b;
    layer4_outputs(10893) <= '1';
    layer4_outputs(10894) <= '0';
    layer4_outputs(10895) <= b and not a;
    layer4_outputs(10896) <= not b;
    layer4_outputs(10897) <= not a or b;
    layer4_outputs(10898) <= a and b;
    layer4_outputs(10899) <= not a or b;
    layer4_outputs(10900) <= not b;
    layer4_outputs(10901) <= b;
    layer4_outputs(10902) <= not b or a;
    layer4_outputs(10903) <= a;
    layer4_outputs(10904) <= not b or a;
    layer4_outputs(10905) <= not b;
    layer4_outputs(10906) <= not a or b;
    layer4_outputs(10907) <= '0';
    layer4_outputs(10908) <= a;
    layer4_outputs(10909) <= not b or a;
    layer4_outputs(10910) <= b;
    layer4_outputs(10911) <= a and b;
    layer4_outputs(10912) <= not b;
    layer4_outputs(10913) <= not (a and b);
    layer4_outputs(10914) <= not a or b;
    layer4_outputs(10915) <= b;
    layer4_outputs(10916) <= b;
    layer4_outputs(10917) <= not a or b;
    layer4_outputs(10918) <= b and not a;
    layer4_outputs(10919) <= b;
    layer4_outputs(10920) <= not b;
    layer4_outputs(10921) <= not a;
    layer4_outputs(10922) <= not a;
    layer4_outputs(10923) <= a or b;
    layer4_outputs(10924) <= a;
    layer4_outputs(10925) <= a;
    layer4_outputs(10926) <= not b;
    layer4_outputs(10927) <= '0';
    layer4_outputs(10928) <= b;
    layer4_outputs(10929) <= a xor b;
    layer4_outputs(10930) <= not b or a;
    layer4_outputs(10931) <= a xor b;
    layer4_outputs(10932) <= a;
    layer4_outputs(10933) <= a and b;
    layer4_outputs(10934) <= a and not b;
    layer4_outputs(10935) <= b;
    layer4_outputs(10936) <= a xor b;
    layer4_outputs(10937) <= a and not b;
    layer4_outputs(10938) <= a;
    layer4_outputs(10939) <= not b;
    layer4_outputs(10940) <= not (a and b);
    layer4_outputs(10941) <= a;
    layer4_outputs(10942) <= not b or a;
    layer4_outputs(10943) <= b;
    layer4_outputs(10944) <= b;
    layer4_outputs(10945) <= a;
    layer4_outputs(10946) <= not (a xor b);
    layer4_outputs(10947) <= a;
    layer4_outputs(10948) <= not b;
    layer4_outputs(10949) <= not b or a;
    layer4_outputs(10950) <= not b;
    layer4_outputs(10951) <= a or b;
    layer4_outputs(10952) <= a;
    layer4_outputs(10953) <= '1';
    layer4_outputs(10954) <= a or b;
    layer4_outputs(10955) <= '0';
    layer4_outputs(10956) <= a and b;
    layer4_outputs(10957) <= a;
    layer4_outputs(10958) <= a and b;
    layer4_outputs(10959) <= b;
    layer4_outputs(10960) <= not b;
    layer4_outputs(10961) <= b;
    layer4_outputs(10962) <= not (a or b);
    layer4_outputs(10963) <= a or b;
    layer4_outputs(10964) <= b;
    layer4_outputs(10965) <= not b or a;
    layer4_outputs(10966) <= b;
    layer4_outputs(10967) <= b;
    layer4_outputs(10968) <= not (a or b);
    layer4_outputs(10969) <= a or b;
    layer4_outputs(10970) <= not a;
    layer4_outputs(10971) <= a or b;
    layer4_outputs(10972) <= not b;
    layer4_outputs(10973) <= not a;
    layer4_outputs(10974) <= not b;
    layer4_outputs(10975) <= b;
    layer4_outputs(10976) <= not a;
    layer4_outputs(10977) <= not (a or b);
    layer4_outputs(10978) <= not b;
    layer4_outputs(10979) <= a and not b;
    layer4_outputs(10980) <= a or b;
    layer4_outputs(10981) <= a and not b;
    layer4_outputs(10982) <= not (a or b);
    layer4_outputs(10983) <= not b;
    layer4_outputs(10984) <= not (a xor b);
    layer4_outputs(10985) <= not b or a;
    layer4_outputs(10986) <= b and not a;
    layer4_outputs(10987) <= not b;
    layer4_outputs(10988) <= not b;
    layer4_outputs(10989) <= b;
    layer4_outputs(10990) <= b;
    layer4_outputs(10991) <= b;
    layer4_outputs(10992) <= a;
    layer4_outputs(10993) <= not a or b;
    layer4_outputs(10994) <= not (a xor b);
    layer4_outputs(10995) <= b;
    layer4_outputs(10996) <= b;
    layer4_outputs(10997) <= not a;
    layer4_outputs(10998) <= a;
    layer4_outputs(10999) <= not b;
    layer4_outputs(11000) <= '1';
    layer4_outputs(11001) <= not b;
    layer4_outputs(11002) <= '1';
    layer4_outputs(11003) <= a;
    layer4_outputs(11004) <= not b;
    layer4_outputs(11005) <= a and b;
    layer4_outputs(11006) <= b;
    layer4_outputs(11007) <= a;
    layer4_outputs(11008) <= '0';
    layer4_outputs(11009) <= not (a xor b);
    layer4_outputs(11010) <= a and not b;
    layer4_outputs(11011) <= not a or b;
    layer4_outputs(11012) <= not a;
    layer4_outputs(11013) <= not b or a;
    layer4_outputs(11014) <= a xor b;
    layer4_outputs(11015) <= a;
    layer4_outputs(11016) <= a;
    layer4_outputs(11017) <= a xor b;
    layer4_outputs(11018) <= a;
    layer4_outputs(11019) <= b and not a;
    layer4_outputs(11020) <= b;
    layer4_outputs(11021) <= not a or b;
    layer4_outputs(11022) <= b and not a;
    layer4_outputs(11023) <= not a;
    layer4_outputs(11024) <= a;
    layer4_outputs(11025) <= a and b;
    layer4_outputs(11026) <= b and not a;
    layer4_outputs(11027) <= not (a xor b);
    layer4_outputs(11028) <= b;
    layer4_outputs(11029) <= '0';
    layer4_outputs(11030) <= not a;
    layer4_outputs(11031) <= a;
    layer4_outputs(11032) <= a and not b;
    layer4_outputs(11033) <= b;
    layer4_outputs(11034) <= not b;
    layer4_outputs(11035) <= a;
    layer4_outputs(11036) <= a;
    layer4_outputs(11037) <= not (a and b);
    layer4_outputs(11038) <= a and not b;
    layer4_outputs(11039) <= a xor b;
    layer4_outputs(11040) <= not (a xor b);
    layer4_outputs(11041) <= b;
    layer4_outputs(11042) <= a and not b;
    layer4_outputs(11043) <= not b or a;
    layer4_outputs(11044) <= not (a or b);
    layer4_outputs(11045) <= not (a and b);
    layer4_outputs(11046) <= a;
    layer4_outputs(11047) <= not a;
    layer4_outputs(11048) <= a and b;
    layer4_outputs(11049) <= not (a xor b);
    layer4_outputs(11050) <= a;
    layer4_outputs(11051) <= b and not a;
    layer4_outputs(11052) <= not a;
    layer4_outputs(11053) <= not b;
    layer4_outputs(11054) <= a xor b;
    layer4_outputs(11055) <= not (a xor b);
    layer4_outputs(11056) <= a;
    layer4_outputs(11057) <= not b;
    layer4_outputs(11058) <= b and not a;
    layer4_outputs(11059) <= b;
    layer4_outputs(11060) <= a and not b;
    layer4_outputs(11061) <= a xor b;
    layer4_outputs(11062) <= not a;
    layer4_outputs(11063) <= a or b;
    layer4_outputs(11064) <= a;
    layer4_outputs(11065) <= not b;
    layer4_outputs(11066) <= b;
    layer4_outputs(11067) <= a and not b;
    layer4_outputs(11068) <= a and not b;
    layer4_outputs(11069) <= b and not a;
    layer4_outputs(11070) <= a or b;
    layer4_outputs(11071) <= a and not b;
    layer4_outputs(11072) <= not (a xor b);
    layer4_outputs(11073) <= a and not b;
    layer4_outputs(11074) <= a;
    layer4_outputs(11075) <= not (a and b);
    layer4_outputs(11076) <= a and b;
    layer4_outputs(11077) <= not b;
    layer4_outputs(11078) <= not b or a;
    layer4_outputs(11079) <= not a;
    layer4_outputs(11080) <= not a;
    layer4_outputs(11081) <= b and not a;
    layer4_outputs(11082) <= not b;
    layer4_outputs(11083) <= not (a or b);
    layer4_outputs(11084) <= a and not b;
    layer4_outputs(11085) <= b;
    layer4_outputs(11086) <= b;
    layer4_outputs(11087) <= not (a and b);
    layer4_outputs(11088) <= not b or a;
    layer4_outputs(11089) <= a or b;
    layer4_outputs(11090) <= a xor b;
    layer4_outputs(11091) <= a or b;
    layer4_outputs(11092) <= '0';
    layer4_outputs(11093) <= not a;
    layer4_outputs(11094) <= not b;
    layer4_outputs(11095) <= b;
    layer4_outputs(11096) <= not b or a;
    layer4_outputs(11097) <= not a or b;
    layer4_outputs(11098) <= b;
    layer4_outputs(11099) <= not a;
    layer4_outputs(11100) <= a xor b;
    layer4_outputs(11101) <= not b;
    layer4_outputs(11102) <= a or b;
    layer4_outputs(11103) <= a and b;
    layer4_outputs(11104) <= not b;
    layer4_outputs(11105) <= b and not a;
    layer4_outputs(11106) <= not (a or b);
    layer4_outputs(11107) <= not a or b;
    layer4_outputs(11108) <= not (a or b);
    layer4_outputs(11109) <= not a;
    layer4_outputs(11110) <= not a;
    layer4_outputs(11111) <= '1';
    layer4_outputs(11112) <= a;
    layer4_outputs(11113) <= a;
    layer4_outputs(11114) <= not (a xor b);
    layer4_outputs(11115) <= not a;
    layer4_outputs(11116) <= '0';
    layer4_outputs(11117) <= '0';
    layer4_outputs(11118) <= not (a xor b);
    layer4_outputs(11119) <= a or b;
    layer4_outputs(11120) <= not a;
    layer4_outputs(11121) <= not a or b;
    layer4_outputs(11122) <= a and b;
    layer4_outputs(11123) <= a or b;
    layer4_outputs(11124) <= a xor b;
    layer4_outputs(11125) <= not b;
    layer4_outputs(11126) <= not a;
    layer4_outputs(11127) <= a;
    layer4_outputs(11128) <= a and b;
    layer4_outputs(11129) <= a or b;
    layer4_outputs(11130) <= a xor b;
    layer4_outputs(11131) <= a;
    layer4_outputs(11132) <= not b or a;
    layer4_outputs(11133) <= a;
    layer4_outputs(11134) <= not b;
    layer4_outputs(11135) <= not a or b;
    layer4_outputs(11136) <= not b;
    layer4_outputs(11137) <= a and b;
    layer4_outputs(11138) <= not (a xor b);
    layer4_outputs(11139) <= b and not a;
    layer4_outputs(11140) <= a and not b;
    layer4_outputs(11141) <= not a;
    layer4_outputs(11142) <= not a;
    layer4_outputs(11143) <= b;
    layer4_outputs(11144) <= not b;
    layer4_outputs(11145) <= not (a xor b);
    layer4_outputs(11146) <= b;
    layer4_outputs(11147) <= not (a or b);
    layer4_outputs(11148) <= b;
    layer4_outputs(11149) <= not b or a;
    layer4_outputs(11150) <= b and not a;
    layer4_outputs(11151) <= not a;
    layer4_outputs(11152) <= a;
    layer4_outputs(11153) <= a and not b;
    layer4_outputs(11154) <= not a;
    layer4_outputs(11155) <= a;
    layer4_outputs(11156) <= a and not b;
    layer4_outputs(11157) <= a and b;
    layer4_outputs(11158) <= a;
    layer4_outputs(11159) <= b and not a;
    layer4_outputs(11160) <= not a;
    layer4_outputs(11161) <= a and b;
    layer4_outputs(11162) <= not b or a;
    layer4_outputs(11163) <= not (a or b);
    layer4_outputs(11164) <= b;
    layer4_outputs(11165) <= a and not b;
    layer4_outputs(11166) <= a and b;
    layer4_outputs(11167) <= not (a and b);
    layer4_outputs(11168) <= not a;
    layer4_outputs(11169) <= not (a and b);
    layer4_outputs(11170) <= not (a or b);
    layer4_outputs(11171) <= not (a and b);
    layer4_outputs(11172) <= a;
    layer4_outputs(11173) <= a xor b;
    layer4_outputs(11174) <= a and not b;
    layer4_outputs(11175) <= a;
    layer4_outputs(11176) <= not b;
    layer4_outputs(11177) <= b;
    layer4_outputs(11178) <= b and not a;
    layer4_outputs(11179) <= not a;
    layer4_outputs(11180) <= not (a xor b);
    layer4_outputs(11181) <= not a;
    layer4_outputs(11182) <= '1';
    layer4_outputs(11183) <= b;
    layer4_outputs(11184) <= a;
    layer4_outputs(11185) <= '0';
    layer4_outputs(11186) <= a or b;
    layer4_outputs(11187) <= not b or a;
    layer4_outputs(11188) <= a or b;
    layer4_outputs(11189) <= '1';
    layer4_outputs(11190) <= a xor b;
    layer4_outputs(11191) <= not b;
    layer4_outputs(11192) <= a;
    layer4_outputs(11193) <= b and not a;
    layer4_outputs(11194) <= a xor b;
    layer4_outputs(11195) <= not (a xor b);
    layer4_outputs(11196) <= not b;
    layer4_outputs(11197) <= not (a and b);
    layer4_outputs(11198) <= not b;
    layer4_outputs(11199) <= b and not a;
    layer4_outputs(11200) <= not (a xor b);
    layer4_outputs(11201) <= a and b;
    layer4_outputs(11202) <= not b;
    layer4_outputs(11203) <= a;
    layer4_outputs(11204) <= a and not b;
    layer4_outputs(11205) <= not a;
    layer4_outputs(11206) <= not b or a;
    layer4_outputs(11207) <= not b or a;
    layer4_outputs(11208) <= b;
    layer4_outputs(11209) <= b;
    layer4_outputs(11210) <= b;
    layer4_outputs(11211) <= not a;
    layer4_outputs(11212) <= not (a xor b);
    layer4_outputs(11213) <= not b or a;
    layer4_outputs(11214) <= a;
    layer4_outputs(11215) <= a and b;
    layer4_outputs(11216) <= a;
    layer4_outputs(11217) <= a;
    layer4_outputs(11218) <= a;
    layer4_outputs(11219) <= not a;
    layer4_outputs(11220) <= a xor b;
    layer4_outputs(11221) <= a or b;
    layer4_outputs(11222) <= a or b;
    layer4_outputs(11223) <= not a or b;
    layer4_outputs(11224) <= a;
    layer4_outputs(11225) <= not b;
    layer4_outputs(11226) <= a;
    layer4_outputs(11227) <= a and not b;
    layer4_outputs(11228) <= a and not b;
    layer4_outputs(11229) <= a;
    layer4_outputs(11230) <= not a;
    layer4_outputs(11231) <= a;
    layer4_outputs(11232) <= not a;
    layer4_outputs(11233) <= not a;
    layer4_outputs(11234) <= not a or b;
    layer4_outputs(11235) <= a;
    layer4_outputs(11236) <= b;
    layer4_outputs(11237) <= not b;
    layer4_outputs(11238) <= a and not b;
    layer4_outputs(11239) <= not b or a;
    layer4_outputs(11240) <= not a;
    layer4_outputs(11241) <= not a;
    layer4_outputs(11242) <= not a;
    layer4_outputs(11243) <= a and not b;
    layer4_outputs(11244) <= not b or a;
    layer4_outputs(11245) <= b;
    layer4_outputs(11246) <= b and not a;
    layer4_outputs(11247) <= not b or a;
    layer4_outputs(11248) <= not (a or b);
    layer4_outputs(11249) <= a xor b;
    layer4_outputs(11250) <= not b;
    layer4_outputs(11251) <= a xor b;
    layer4_outputs(11252) <= not b or a;
    layer4_outputs(11253) <= a;
    layer4_outputs(11254) <= b;
    layer4_outputs(11255) <= not b;
    layer4_outputs(11256) <= not a;
    layer4_outputs(11257) <= b and not a;
    layer4_outputs(11258) <= a;
    layer4_outputs(11259) <= not b;
    layer4_outputs(11260) <= a and b;
    layer4_outputs(11261) <= '1';
    layer4_outputs(11262) <= not (a xor b);
    layer4_outputs(11263) <= a or b;
    layer4_outputs(11264) <= b and not a;
    layer4_outputs(11265) <= a xor b;
    layer4_outputs(11266) <= a and not b;
    layer4_outputs(11267) <= not (a and b);
    layer4_outputs(11268) <= not a or b;
    layer4_outputs(11269) <= a or b;
    layer4_outputs(11270) <= not b;
    layer4_outputs(11271) <= not b;
    layer4_outputs(11272) <= not (a or b);
    layer4_outputs(11273) <= a xor b;
    layer4_outputs(11274) <= not a;
    layer4_outputs(11275) <= a or b;
    layer4_outputs(11276) <= not b;
    layer4_outputs(11277) <= not a;
    layer4_outputs(11278) <= not b or a;
    layer4_outputs(11279) <= '1';
    layer4_outputs(11280) <= not (a and b);
    layer4_outputs(11281) <= not (a and b);
    layer4_outputs(11282) <= a or b;
    layer4_outputs(11283) <= not b;
    layer4_outputs(11284) <= a or b;
    layer4_outputs(11285) <= a and b;
    layer4_outputs(11286) <= a and not b;
    layer4_outputs(11287) <= not (a xor b);
    layer4_outputs(11288) <= not (a xor b);
    layer4_outputs(11289) <= not (a or b);
    layer4_outputs(11290) <= not (a xor b);
    layer4_outputs(11291) <= not a;
    layer4_outputs(11292) <= not b;
    layer4_outputs(11293) <= a or b;
    layer4_outputs(11294) <= b and not a;
    layer4_outputs(11295) <= b;
    layer4_outputs(11296) <= not (a or b);
    layer4_outputs(11297) <= a xor b;
    layer4_outputs(11298) <= a or b;
    layer4_outputs(11299) <= a;
    layer4_outputs(11300) <= not b or a;
    layer4_outputs(11301) <= a;
    layer4_outputs(11302) <= not b;
    layer4_outputs(11303) <= not (a or b);
    layer4_outputs(11304) <= not a;
    layer4_outputs(11305) <= not a;
    layer4_outputs(11306) <= b and not a;
    layer4_outputs(11307) <= not b or a;
    layer4_outputs(11308) <= a xor b;
    layer4_outputs(11309) <= a;
    layer4_outputs(11310) <= not (a and b);
    layer4_outputs(11311) <= a and b;
    layer4_outputs(11312) <= a;
    layer4_outputs(11313) <= a xor b;
    layer4_outputs(11314) <= b and not a;
    layer4_outputs(11315) <= not (a xor b);
    layer4_outputs(11316) <= not (a or b);
    layer4_outputs(11317) <= a and b;
    layer4_outputs(11318) <= not b;
    layer4_outputs(11319) <= not a or b;
    layer4_outputs(11320) <= not (a or b);
    layer4_outputs(11321) <= not (a or b);
    layer4_outputs(11322) <= not b;
    layer4_outputs(11323) <= a;
    layer4_outputs(11324) <= a;
    layer4_outputs(11325) <= '0';
    layer4_outputs(11326) <= not (a xor b);
    layer4_outputs(11327) <= a and not b;
    layer4_outputs(11328) <= not b;
    layer4_outputs(11329) <= a and b;
    layer4_outputs(11330) <= a or b;
    layer4_outputs(11331) <= not b;
    layer4_outputs(11332) <= not b;
    layer4_outputs(11333) <= a xor b;
    layer4_outputs(11334) <= not b or a;
    layer4_outputs(11335) <= not a;
    layer4_outputs(11336) <= a or b;
    layer4_outputs(11337) <= not a;
    layer4_outputs(11338) <= a and b;
    layer4_outputs(11339) <= a;
    layer4_outputs(11340) <= a;
    layer4_outputs(11341) <= not (a and b);
    layer4_outputs(11342) <= '1';
    layer4_outputs(11343) <= not b;
    layer4_outputs(11344) <= not (a xor b);
    layer4_outputs(11345) <= not (a and b);
    layer4_outputs(11346) <= not (a and b);
    layer4_outputs(11347) <= a;
    layer4_outputs(11348) <= b and not a;
    layer4_outputs(11349) <= not b;
    layer4_outputs(11350) <= not (a or b);
    layer4_outputs(11351) <= not a;
    layer4_outputs(11352) <= a or b;
    layer4_outputs(11353) <= not a;
    layer4_outputs(11354) <= a or b;
    layer4_outputs(11355) <= a and not b;
    layer4_outputs(11356) <= not b or a;
    layer4_outputs(11357) <= a;
    layer4_outputs(11358) <= a;
    layer4_outputs(11359) <= not a;
    layer4_outputs(11360) <= a;
    layer4_outputs(11361) <= not b or a;
    layer4_outputs(11362) <= not a;
    layer4_outputs(11363) <= b and not a;
    layer4_outputs(11364) <= a;
    layer4_outputs(11365) <= a and b;
    layer4_outputs(11366) <= a and not b;
    layer4_outputs(11367) <= not b;
    layer4_outputs(11368) <= a;
    layer4_outputs(11369) <= a;
    layer4_outputs(11370) <= a or b;
    layer4_outputs(11371) <= a;
    layer4_outputs(11372) <= a;
    layer4_outputs(11373) <= not (a xor b);
    layer4_outputs(11374) <= a or b;
    layer4_outputs(11375) <= not a;
    layer4_outputs(11376) <= a;
    layer4_outputs(11377) <= a;
    layer4_outputs(11378) <= not a or b;
    layer4_outputs(11379) <= b;
    layer4_outputs(11380) <= a and not b;
    layer4_outputs(11381) <= not a or b;
    layer4_outputs(11382) <= b and not a;
    layer4_outputs(11383) <= b;
    layer4_outputs(11384) <= not (a and b);
    layer4_outputs(11385) <= not a;
    layer4_outputs(11386) <= b and not a;
    layer4_outputs(11387) <= not a;
    layer4_outputs(11388) <= a or b;
    layer4_outputs(11389) <= a xor b;
    layer4_outputs(11390) <= a;
    layer4_outputs(11391) <= b;
    layer4_outputs(11392) <= not (a and b);
    layer4_outputs(11393) <= a;
    layer4_outputs(11394) <= a;
    layer4_outputs(11395) <= not a or b;
    layer4_outputs(11396) <= a xor b;
    layer4_outputs(11397) <= '1';
    layer4_outputs(11398) <= not a;
    layer4_outputs(11399) <= not a;
    layer4_outputs(11400) <= not a or b;
    layer4_outputs(11401) <= a;
    layer4_outputs(11402) <= b;
    layer4_outputs(11403) <= not a;
    layer4_outputs(11404) <= a or b;
    layer4_outputs(11405) <= not a;
    layer4_outputs(11406) <= a and not b;
    layer4_outputs(11407) <= b;
    layer4_outputs(11408) <= not b or a;
    layer4_outputs(11409) <= a and b;
    layer4_outputs(11410) <= a and b;
    layer4_outputs(11411) <= not (a or b);
    layer4_outputs(11412) <= not a or b;
    layer4_outputs(11413) <= b;
    layer4_outputs(11414) <= '0';
    layer4_outputs(11415) <= a;
    layer4_outputs(11416) <= a and b;
    layer4_outputs(11417) <= not b;
    layer4_outputs(11418) <= not a;
    layer4_outputs(11419) <= not a;
    layer4_outputs(11420) <= a or b;
    layer4_outputs(11421) <= b;
    layer4_outputs(11422) <= a xor b;
    layer4_outputs(11423) <= not a;
    layer4_outputs(11424) <= a and not b;
    layer4_outputs(11425) <= b;
    layer4_outputs(11426) <= not (a or b);
    layer4_outputs(11427) <= b;
    layer4_outputs(11428) <= b;
    layer4_outputs(11429) <= b;
    layer4_outputs(11430) <= b;
    layer4_outputs(11431) <= a and not b;
    layer4_outputs(11432) <= not b;
    layer4_outputs(11433) <= b;
    layer4_outputs(11434) <= '1';
    layer4_outputs(11435) <= a or b;
    layer4_outputs(11436) <= not (a or b);
    layer4_outputs(11437) <= not (a or b);
    layer4_outputs(11438) <= not b or a;
    layer4_outputs(11439) <= not a;
    layer4_outputs(11440) <= b;
    layer4_outputs(11441) <= a;
    layer4_outputs(11442) <= '0';
    layer4_outputs(11443) <= not b;
    layer4_outputs(11444) <= not (a and b);
    layer4_outputs(11445) <= not a;
    layer4_outputs(11446) <= not b;
    layer4_outputs(11447) <= not (a and b);
    layer4_outputs(11448) <= a;
    layer4_outputs(11449) <= b and not a;
    layer4_outputs(11450) <= a xor b;
    layer4_outputs(11451) <= a and not b;
    layer4_outputs(11452) <= a and b;
    layer4_outputs(11453) <= '1';
    layer4_outputs(11454) <= a and not b;
    layer4_outputs(11455) <= a and b;
    layer4_outputs(11456) <= not (a xor b);
    layer4_outputs(11457) <= not (a and b);
    layer4_outputs(11458) <= not a;
    layer4_outputs(11459) <= '1';
    layer4_outputs(11460) <= b and not a;
    layer4_outputs(11461) <= not b;
    layer4_outputs(11462) <= a and b;
    layer4_outputs(11463) <= not b or a;
    layer4_outputs(11464) <= b;
    layer4_outputs(11465) <= a xor b;
    layer4_outputs(11466) <= not a or b;
    layer4_outputs(11467) <= not b or a;
    layer4_outputs(11468) <= not (a or b);
    layer4_outputs(11469) <= not (a xor b);
    layer4_outputs(11470) <= a;
    layer4_outputs(11471) <= a;
    layer4_outputs(11472) <= not (a and b);
    layer4_outputs(11473) <= '1';
    layer4_outputs(11474) <= not a or b;
    layer4_outputs(11475) <= a xor b;
    layer4_outputs(11476) <= not b or a;
    layer4_outputs(11477) <= b and not a;
    layer4_outputs(11478) <= a and not b;
    layer4_outputs(11479) <= a;
    layer4_outputs(11480) <= a xor b;
    layer4_outputs(11481) <= not (a xor b);
    layer4_outputs(11482) <= not a;
    layer4_outputs(11483) <= a and b;
    layer4_outputs(11484) <= b;
    layer4_outputs(11485) <= not a or b;
    layer4_outputs(11486) <= not a;
    layer4_outputs(11487) <= not b or a;
    layer4_outputs(11488) <= '0';
    layer4_outputs(11489) <= not a;
    layer4_outputs(11490) <= not (a xor b);
    layer4_outputs(11491) <= b;
    layer4_outputs(11492) <= not b;
    layer4_outputs(11493) <= a;
    layer4_outputs(11494) <= not a or b;
    layer4_outputs(11495) <= not (a and b);
    layer4_outputs(11496) <= not b;
    layer4_outputs(11497) <= b;
    layer4_outputs(11498) <= b;
    layer4_outputs(11499) <= b and not a;
    layer4_outputs(11500) <= not (a or b);
    layer4_outputs(11501) <= not b or a;
    layer4_outputs(11502) <= not b or a;
    layer4_outputs(11503) <= not (a or b);
    layer4_outputs(11504) <= a or b;
    layer4_outputs(11505) <= b and not a;
    layer4_outputs(11506) <= a;
    layer4_outputs(11507) <= b;
    layer4_outputs(11508) <= b;
    layer4_outputs(11509) <= not a;
    layer4_outputs(11510) <= not a;
    layer4_outputs(11511) <= '0';
    layer4_outputs(11512) <= a and b;
    layer4_outputs(11513) <= not (a xor b);
    layer4_outputs(11514) <= '0';
    layer4_outputs(11515) <= a or b;
    layer4_outputs(11516) <= a;
    layer4_outputs(11517) <= a or b;
    layer4_outputs(11518) <= not b;
    layer4_outputs(11519) <= not b;
    layer4_outputs(11520) <= b and not a;
    layer4_outputs(11521) <= not a;
    layer4_outputs(11522) <= a or b;
    layer4_outputs(11523) <= b;
    layer4_outputs(11524) <= a xor b;
    layer4_outputs(11525) <= b and not a;
    layer4_outputs(11526) <= a and b;
    layer4_outputs(11527) <= a and not b;
    layer4_outputs(11528) <= not b;
    layer4_outputs(11529) <= b;
    layer4_outputs(11530) <= a;
    layer4_outputs(11531) <= not b;
    layer4_outputs(11532) <= not (a and b);
    layer4_outputs(11533) <= not a;
    layer4_outputs(11534) <= a and not b;
    layer4_outputs(11535) <= not (a xor b);
    layer4_outputs(11536) <= a and b;
    layer4_outputs(11537) <= not (a and b);
    layer4_outputs(11538) <= b;
    layer4_outputs(11539) <= a and b;
    layer4_outputs(11540) <= b;
    layer4_outputs(11541) <= not (a xor b);
    layer4_outputs(11542) <= not a;
    layer4_outputs(11543) <= not b;
    layer4_outputs(11544) <= a or b;
    layer4_outputs(11545) <= b;
    layer4_outputs(11546) <= a or b;
    layer4_outputs(11547) <= not b;
    layer4_outputs(11548) <= a xor b;
    layer4_outputs(11549) <= not a or b;
    layer4_outputs(11550) <= b and not a;
    layer4_outputs(11551) <= not (a and b);
    layer4_outputs(11552) <= '1';
    layer4_outputs(11553) <= not b;
    layer4_outputs(11554) <= not a;
    layer4_outputs(11555) <= not b;
    layer4_outputs(11556) <= b;
    layer4_outputs(11557) <= a;
    layer4_outputs(11558) <= not (a and b);
    layer4_outputs(11559) <= not b;
    layer4_outputs(11560) <= b;
    layer4_outputs(11561) <= not (a or b);
    layer4_outputs(11562) <= b;
    layer4_outputs(11563) <= a and b;
    layer4_outputs(11564) <= not (a and b);
    layer4_outputs(11565) <= not (a xor b);
    layer4_outputs(11566) <= not a or b;
    layer4_outputs(11567) <= not a or b;
    layer4_outputs(11568) <= not b;
    layer4_outputs(11569) <= not (a and b);
    layer4_outputs(11570) <= b and not a;
    layer4_outputs(11571) <= not b;
    layer4_outputs(11572) <= a;
    layer4_outputs(11573) <= a and not b;
    layer4_outputs(11574) <= not b;
    layer4_outputs(11575) <= not (a or b);
    layer4_outputs(11576) <= not (a xor b);
    layer4_outputs(11577) <= not b;
    layer4_outputs(11578) <= not a;
    layer4_outputs(11579) <= b;
    layer4_outputs(11580) <= not b;
    layer4_outputs(11581) <= not a;
    layer4_outputs(11582) <= not (a or b);
    layer4_outputs(11583) <= b;
    layer4_outputs(11584) <= b;
    layer4_outputs(11585) <= not a;
    layer4_outputs(11586) <= not b or a;
    layer4_outputs(11587) <= not (a and b);
    layer4_outputs(11588) <= not a or b;
    layer4_outputs(11589) <= not a;
    layer4_outputs(11590) <= not a;
    layer4_outputs(11591) <= not (a or b);
    layer4_outputs(11592) <= not a or b;
    layer4_outputs(11593) <= a xor b;
    layer4_outputs(11594) <= a;
    layer4_outputs(11595) <= not b or a;
    layer4_outputs(11596) <= b;
    layer4_outputs(11597) <= not (a and b);
    layer4_outputs(11598) <= b;
    layer4_outputs(11599) <= not a;
    layer4_outputs(11600) <= not a or b;
    layer4_outputs(11601) <= not (a or b);
    layer4_outputs(11602) <= a or b;
    layer4_outputs(11603) <= not (a xor b);
    layer4_outputs(11604) <= a and not b;
    layer4_outputs(11605) <= not a or b;
    layer4_outputs(11606) <= b;
    layer4_outputs(11607) <= a and b;
    layer4_outputs(11608) <= not b;
    layer4_outputs(11609) <= b;
    layer4_outputs(11610) <= b;
    layer4_outputs(11611) <= b;
    layer4_outputs(11612) <= not (a and b);
    layer4_outputs(11613) <= a or b;
    layer4_outputs(11614) <= not a or b;
    layer4_outputs(11615) <= not a;
    layer4_outputs(11616) <= a and b;
    layer4_outputs(11617) <= not (a xor b);
    layer4_outputs(11618) <= not a or b;
    layer4_outputs(11619) <= not a;
    layer4_outputs(11620) <= not (a or b);
    layer4_outputs(11621) <= not b;
    layer4_outputs(11622) <= not b;
    layer4_outputs(11623) <= a and not b;
    layer4_outputs(11624) <= not b;
    layer4_outputs(11625) <= not b;
    layer4_outputs(11626) <= not b;
    layer4_outputs(11627) <= not (a or b);
    layer4_outputs(11628) <= not a or b;
    layer4_outputs(11629) <= b;
    layer4_outputs(11630) <= a or b;
    layer4_outputs(11631) <= not b;
    layer4_outputs(11632) <= not (a or b);
    layer4_outputs(11633) <= not a;
    layer4_outputs(11634) <= b;
    layer4_outputs(11635) <= b and not a;
    layer4_outputs(11636) <= a and b;
    layer4_outputs(11637) <= a and not b;
    layer4_outputs(11638) <= a xor b;
    layer4_outputs(11639) <= a or b;
    layer4_outputs(11640) <= not a;
    layer4_outputs(11641) <= a or b;
    layer4_outputs(11642) <= not a;
    layer4_outputs(11643) <= b;
    layer4_outputs(11644) <= not (a and b);
    layer4_outputs(11645) <= '1';
    layer4_outputs(11646) <= b;
    layer4_outputs(11647) <= a xor b;
    layer4_outputs(11648) <= b;
    layer4_outputs(11649) <= b and not a;
    layer4_outputs(11650) <= not a;
    layer4_outputs(11651) <= not a;
    layer4_outputs(11652) <= not b;
    layer4_outputs(11653) <= a;
    layer4_outputs(11654) <= not a;
    layer4_outputs(11655) <= not (a and b);
    layer4_outputs(11656) <= a and b;
    layer4_outputs(11657) <= b;
    layer4_outputs(11658) <= not b;
    layer4_outputs(11659) <= b;
    layer4_outputs(11660) <= not (a xor b);
    layer4_outputs(11661) <= not (a xor b);
    layer4_outputs(11662) <= not (a and b);
    layer4_outputs(11663) <= a and not b;
    layer4_outputs(11664) <= not (a xor b);
    layer4_outputs(11665) <= not b;
    layer4_outputs(11666) <= a xor b;
    layer4_outputs(11667) <= a;
    layer4_outputs(11668) <= a;
    layer4_outputs(11669) <= not (a and b);
    layer4_outputs(11670) <= not a or b;
    layer4_outputs(11671) <= not (a xor b);
    layer4_outputs(11672) <= a and b;
    layer4_outputs(11673) <= a and not b;
    layer4_outputs(11674) <= not (a xor b);
    layer4_outputs(11675) <= a and b;
    layer4_outputs(11676) <= not b;
    layer4_outputs(11677) <= b;
    layer4_outputs(11678) <= '0';
    layer4_outputs(11679) <= a and not b;
    layer4_outputs(11680) <= a or b;
    layer4_outputs(11681) <= not (a and b);
    layer4_outputs(11682) <= a;
    layer4_outputs(11683) <= not b;
    layer4_outputs(11684) <= not a or b;
    layer4_outputs(11685) <= not b or a;
    layer4_outputs(11686) <= a xor b;
    layer4_outputs(11687) <= a xor b;
    layer4_outputs(11688) <= a;
    layer4_outputs(11689) <= b;
    layer4_outputs(11690) <= not b;
    layer4_outputs(11691) <= not b;
    layer4_outputs(11692) <= a;
    layer4_outputs(11693) <= not b;
    layer4_outputs(11694) <= not (a xor b);
    layer4_outputs(11695) <= a and b;
    layer4_outputs(11696) <= b and not a;
    layer4_outputs(11697) <= b;
    layer4_outputs(11698) <= not a or b;
    layer4_outputs(11699) <= a or b;
    layer4_outputs(11700) <= a or b;
    layer4_outputs(11701) <= not a or b;
    layer4_outputs(11702) <= not (a and b);
    layer4_outputs(11703) <= not a;
    layer4_outputs(11704) <= a and not b;
    layer4_outputs(11705) <= b;
    layer4_outputs(11706) <= '1';
    layer4_outputs(11707) <= not b or a;
    layer4_outputs(11708) <= not a;
    layer4_outputs(11709) <= not b;
    layer4_outputs(11710) <= '0';
    layer4_outputs(11711) <= '0';
    layer4_outputs(11712) <= a xor b;
    layer4_outputs(11713) <= not b;
    layer4_outputs(11714) <= b;
    layer4_outputs(11715) <= a;
    layer4_outputs(11716) <= a and not b;
    layer4_outputs(11717) <= not a;
    layer4_outputs(11718) <= not a;
    layer4_outputs(11719) <= a xor b;
    layer4_outputs(11720) <= a and not b;
    layer4_outputs(11721) <= a xor b;
    layer4_outputs(11722) <= not a;
    layer4_outputs(11723) <= not (a or b);
    layer4_outputs(11724) <= b;
    layer4_outputs(11725) <= not a;
    layer4_outputs(11726) <= a;
    layer4_outputs(11727) <= not (a or b);
    layer4_outputs(11728) <= not a;
    layer4_outputs(11729) <= '1';
    layer4_outputs(11730) <= '1';
    layer4_outputs(11731) <= b and not a;
    layer4_outputs(11732) <= not b;
    layer4_outputs(11733) <= '0';
    layer4_outputs(11734) <= a or b;
    layer4_outputs(11735) <= b;
    layer4_outputs(11736) <= a xor b;
    layer4_outputs(11737) <= b;
    layer4_outputs(11738) <= not b or a;
    layer4_outputs(11739) <= a and b;
    layer4_outputs(11740) <= a;
    layer4_outputs(11741) <= not b;
    layer4_outputs(11742) <= not (a or b);
    layer4_outputs(11743) <= not (a xor b);
    layer4_outputs(11744) <= a xor b;
    layer4_outputs(11745) <= a;
    layer4_outputs(11746) <= not a or b;
    layer4_outputs(11747) <= b;
    layer4_outputs(11748) <= not a or b;
    layer4_outputs(11749) <= a and not b;
    layer4_outputs(11750) <= not a or b;
    layer4_outputs(11751) <= '1';
    layer4_outputs(11752) <= not b or a;
    layer4_outputs(11753) <= b and not a;
    layer4_outputs(11754) <= not a;
    layer4_outputs(11755) <= not (a or b);
    layer4_outputs(11756) <= not (a and b);
    layer4_outputs(11757) <= b;
    layer4_outputs(11758) <= a;
    layer4_outputs(11759) <= not a;
    layer4_outputs(11760) <= a;
    layer4_outputs(11761) <= a;
    layer4_outputs(11762) <= not b;
    layer4_outputs(11763) <= a or b;
    layer4_outputs(11764) <= a and not b;
    layer4_outputs(11765) <= b and not a;
    layer4_outputs(11766) <= not (a xor b);
    layer4_outputs(11767) <= not b;
    layer4_outputs(11768) <= not a;
    layer4_outputs(11769) <= not (a xor b);
    layer4_outputs(11770) <= not (a and b);
    layer4_outputs(11771) <= a xor b;
    layer4_outputs(11772) <= not b;
    layer4_outputs(11773) <= not a;
    layer4_outputs(11774) <= not b;
    layer4_outputs(11775) <= b;
    layer4_outputs(11776) <= a and not b;
    layer4_outputs(11777) <= not (a xor b);
    layer4_outputs(11778) <= not b;
    layer4_outputs(11779) <= a;
    layer4_outputs(11780) <= a and b;
    layer4_outputs(11781) <= b;
    layer4_outputs(11782) <= '1';
    layer4_outputs(11783) <= not a;
    layer4_outputs(11784) <= not a;
    layer4_outputs(11785) <= a xor b;
    layer4_outputs(11786) <= b and not a;
    layer4_outputs(11787) <= not a;
    layer4_outputs(11788) <= b;
    layer4_outputs(11789) <= a;
    layer4_outputs(11790) <= b;
    layer4_outputs(11791) <= not (a or b);
    layer4_outputs(11792) <= a xor b;
    layer4_outputs(11793) <= not (a xor b);
    layer4_outputs(11794) <= not a or b;
    layer4_outputs(11795) <= not (a or b);
    layer4_outputs(11796) <= a and b;
    layer4_outputs(11797) <= not (a or b);
    layer4_outputs(11798) <= not a or b;
    layer4_outputs(11799) <= not (a and b);
    layer4_outputs(11800) <= a and not b;
    layer4_outputs(11801) <= '1';
    layer4_outputs(11802) <= not (a and b);
    layer4_outputs(11803) <= a or b;
    layer4_outputs(11804) <= '0';
    layer4_outputs(11805) <= a xor b;
    layer4_outputs(11806) <= a xor b;
    layer4_outputs(11807) <= b;
    layer4_outputs(11808) <= a and b;
    layer4_outputs(11809) <= not b;
    layer4_outputs(11810) <= not (a xor b);
    layer4_outputs(11811) <= not a;
    layer4_outputs(11812) <= not (a xor b);
    layer4_outputs(11813) <= not b;
    layer4_outputs(11814) <= not b;
    layer4_outputs(11815) <= not a;
    layer4_outputs(11816) <= not (a or b);
    layer4_outputs(11817) <= a or b;
    layer4_outputs(11818) <= a;
    layer4_outputs(11819) <= a;
    layer4_outputs(11820) <= not (a or b);
    layer4_outputs(11821) <= b and not a;
    layer4_outputs(11822) <= b and not a;
    layer4_outputs(11823) <= b and not a;
    layer4_outputs(11824) <= a and not b;
    layer4_outputs(11825) <= a xor b;
    layer4_outputs(11826) <= a xor b;
    layer4_outputs(11827) <= '0';
    layer4_outputs(11828) <= not (a and b);
    layer4_outputs(11829) <= not a;
    layer4_outputs(11830) <= a;
    layer4_outputs(11831) <= b;
    layer4_outputs(11832) <= a and not b;
    layer4_outputs(11833) <= not a;
    layer4_outputs(11834) <= a;
    layer4_outputs(11835) <= not b;
    layer4_outputs(11836) <= a;
    layer4_outputs(11837) <= not a or b;
    layer4_outputs(11838) <= not a;
    layer4_outputs(11839) <= a;
    layer4_outputs(11840) <= b and not a;
    layer4_outputs(11841) <= b;
    layer4_outputs(11842) <= not b;
    layer4_outputs(11843) <= not a;
    layer4_outputs(11844) <= not a;
    layer4_outputs(11845) <= b and not a;
    layer4_outputs(11846) <= not a;
    layer4_outputs(11847) <= b and not a;
    layer4_outputs(11848) <= b;
    layer4_outputs(11849) <= a and b;
    layer4_outputs(11850) <= b;
    layer4_outputs(11851) <= not b;
    layer4_outputs(11852) <= not a;
    layer4_outputs(11853) <= a or b;
    layer4_outputs(11854) <= a or b;
    layer4_outputs(11855) <= not a;
    layer4_outputs(11856) <= b;
    layer4_outputs(11857) <= b;
    layer4_outputs(11858) <= not a;
    layer4_outputs(11859) <= b;
    layer4_outputs(11860) <= a and b;
    layer4_outputs(11861) <= not (a and b);
    layer4_outputs(11862) <= not b or a;
    layer4_outputs(11863) <= a and b;
    layer4_outputs(11864) <= a or b;
    layer4_outputs(11865) <= not b;
    layer4_outputs(11866) <= a and b;
    layer4_outputs(11867) <= a;
    layer4_outputs(11868) <= a or b;
    layer4_outputs(11869) <= not a or b;
    layer4_outputs(11870) <= not (a xor b);
    layer4_outputs(11871) <= not (a and b);
    layer4_outputs(11872) <= b and not a;
    layer4_outputs(11873) <= not a;
    layer4_outputs(11874) <= not (a and b);
    layer4_outputs(11875) <= not b or a;
    layer4_outputs(11876) <= b;
    layer4_outputs(11877) <= not a;
    layer4_outputs(11878) <= not (a and b);
    layer4_outputs(11879) <= b and not a;
    layer4_outputs(11880) <= b;
    layer4_outputs(11881) <= b and not a;
    layer4_outputs(11882) <= not (a xor b);
    layer4_outputs(11883) <= not b or a;
    layer4_outputs(11884) <= not a;
    layer4_outputs(11885) <= not (a xor b);
    layer4_outputs(11886) <= not (a and b);
    layer4_outputs(11887) <= not a;
    layer4_outputs(11888) <= not b;
    layer4_outputs(11889) <= not b;
    layer4_outputs(11890) <= b;
    layer4_outputs(11891) <= a;
    layer4_outputs(11892) <= not (a or b);
    layer4_outputs(11893) <= b;
    layer4_outputs(11894) <= a and not b;
    layer4_outputs(11895) <= a and not b;
    layer4_outputs(11896) <= a or b;
    layer4_outputs(11897) <= '1';
    layer4_outputs(11898) <= not (a or b);
    layer4_outputs(11899) <= not a;
    layer4_outputs(11900) <= not (a xor b);
    layer4_outputs(11901) <= not b or a;
    layer4_outputs(11902) <= b and not a;
    layer4_outputs(11903) <= not a;
    layer4_outputs(11904) <= a and b;
    layer4_outputs(11905) <= b;
    layer4_outputs(11906) <= b and not a;
    layer4_outputs(11907) <= not a;
    layer4_outputs(11908) <= not (a and b);
    layer4_outputs(11909) <= b;
    layer4_outputs(11910) <= not b or a;
    layer4_outputs(11911) <= b;
    layer4_outputs(11912) <= not (a or b);
    layer4_outputs(11913) <= a and not b;
    layer4_outputs(11914) <= '1';
    layer4_outputs(11915) <= a xor b;
    layer4_outputs(11916) <= a and not b;
    layer4_outputs(11917) <= b and not a;
    layer4_outputs(11918) <= not (a or b);
    layer4_outputs(11919) <= not a;
    layer4_outputs(11920) <= not (a or b);
    layer4_outputs(11921) <= a;
    layer4_outputs(11922) <= a or b;
    layer4_outputs(11923) <= not a;
    layer4_outputs(11924) <= b;
    layer4_outputs(11925) <= b and not a;
    layer4_outputs(11926) <= not a or b;
    layer4_outputs(11927) <= not a or b;
    layer4_outputs(11928) <= a and b;
    layer4_outputs(11929) <= a or b;
    layer4_outputs(11930) <= not a;
    layer4_outputs(11931) <= not b;
    layer4_outputs(11932) <= a and not b;
    layer4_outputs(11933) <= a or b;
    layer4_outputs(11934) <= not b or a;
    layer4_outputs(11935) <= not a;
    layer4_outputs(11936) <= a;
    layer4_outputs(11937) <= not a;
    layer4_outputs(11938) <= b;
    layer4_outputs(11939) <= a and not b;
    layer4_outputs(11940) <= not a;
    layer4_outputs(11941) <= a and not b;
    layer4_outputs(11942) <= not a or b;
    layer4_outputs(11943) <= not b;
    layer4_outputs(11944) <= a;
    layer4_outputs(11945) <= a and b;
    layer4_outputs(11946) <= b;
    layer4_outputs(11947) <= not (a xor b);
    layer4_outputs(11948) <= not b;
    layer4_outputs(11949) <= not b;
    layer4_outputs(11950) <= not b;
    layer4_outputs(11951) <= '1';
    layer4_outputs(11952) <= '0';
    layer4_outputs(11953) <= not a or b;
    layer4_outputs(11954) <= not a;
    layer4_outputs(11955) <= not b;
    layer4_outputs(11956) <= not (a xor b);
    layer4_outputs(11957) <= a and not b;
    layer4_outputs(11958) <= a and not b;
    layer4_outputs(11959) <= not b;
    layer4_outputs(11960) <= b and not a;
    layer4_outputs(11961) <= a and b;
    layer4_outputs(11962) <= not b or a;
    layer4_outputs(11963) <= not a;
    layer4_outputs(11964) <= not b;
    layer4_outputs(11965) <= not b;
    layer4_outputs(11966) <= a xor b;
    layer4_outputs(11967) <= a xor b;
    layer4_outputs(11968) <= b;
    layer4_outputs(11969) <= b;
    layer4_outputs(11970) <= a;
    layer4_outputs(11971) <= '1';
    layer4_outputs(11972) <= not (a or b);
    layer4_outputs(11973) <= b and not a;
    layer4_outputs(11974) <= not b;
    layer4_outputs(11975) <= a;
    layer4_outputs(11976) <= a and b;
    layer4_outputs(11977) <= a xor b;
    layer4_outputs(11978) <= b;
    layer4_outputs(11979) <= not a;
    layer4_outputs(11980) <= a and b;
    layer4_outputs(11981) <= b and not a;
    layer4_outputs(11982) <= b;
    layer4_outputs(11983) <= not (a xor b);
    layer4_outputs(11984) <= a and not b;
    layer4_outputs(11985) <= not (a and b);
    layer4_outputs(11986) <= not b;
    layer4_outputs(11987) <= '0';
    layer4_outputs(11988) <= not (a and b);
    layer4_outputs(11989) <= a xor b;
    layer4_outputs(11990) <= b;
    layer4_outputs(11991) <= b;
    layer4_outputs(11992) <= not b;
    layer4_outputs(11993) <= not a;
    layer4_outputs(11994) <= not b;
    layer4_outputs(11995) <= not a;
    layer4_outputs(11996) <= b;
    layer4_outputs(11997) <= not b or a;
    layer4_outputs(11998) <= a or b;
    layer4_outputs(11999) <= '0';
    layer4_outputs(12000) <= a;
    layer4_outputs(12001) <= b and not a;
    layer4_outputs(12002) <= not b or a;
    layer4_outputs(12003) <= a and not b;
    layer4_outputs(12004) <= not a;
    layer4_outputs(12005) <= a xor b;
    layer4_outputs(12006) <= not b;
    layer4_outputs(12007) <= not b;
    layer4_outputs(12008) <= not (a and b);
    layer4_outputs(12009) <= b;
    layer4_outputs(12010) <= a or b;
    layer4_outputs(12011) <= not (a or b);
    layer4_outputs(12012) <= not a;
    layer4_outputs(12013) <= a or b;
    layer4_outputs(12014) <= not a;
    layer4_outputs(12015) <= not (a or b);
    layer4_outputs(12016) <= not a;
    layer4_outputs(12017) <= not (a xor b);
    layer4_outputs(12018) <= a xor b;
    layer4_outputs(12019) <= b and not a;
    layer4_outputs(12020) <= not a;
    layer4_outputs(12021) <= a;
    layer4_outputs(12022) <= not (a or b);
    layer4_outputs(12023) <= not a;
    layer4_outputs(12024) <= b;
    layer4_outputs(12025) <= a or b;
    layer4_outputs(12026) <= a or b;
    layer4_outputs(12027) <= b;
    layer4_outputs(12028) <= b;
    layer4_outputs(12029) <= not a;
    layer4_outputs(12030) <= not a;
    layer4_outputs(12031) <= not b or a;
    layer4_outputs(12032) <= b and not a;
    layer4_outputs(12033) <= a or b;
    layer4_outputs(12034) <= not b or a;
    layer4_outputs(12035) <= not a;
    layer4_outputs(12036) <= '0';
    layer4_outputs(12037) <= a and not b;
    layer4_outputs(12038) <= not a;
    layer4_outputs(12039) <= a;
    layer4_outputs(12040) <= not a or b;
    layer4_outputs(12041) <= b;
    layer4_outputs(12042) <= not a;
    layer4_outputs(12043) <= a or b;
    layer4_outputs(12044) <= a;
    layer4_outputs(12045) <= a;
    layer4_outputs(12046) <= a and not b;
    layer4_outputs(12047) <= a and b;
    layer4_outputs(12048) <= not b or a;
    layer4_outputs(12049) <= a or b;
    layer4_outputs(12050) <= a;
    layer4_outputs(12051) <= not (a or b);
    layer4_outputs(12052) <= a or b;
    layer4_outputs(12053) <= not a;
    layer4_outputs(12054) <= not (a or b);
    layer4_outputs(12055) <= not a or b;
    layer4_outputs(12056) <= not (a xor b);
    layer4_outputs(12057) <= a;
    layer4_outputs(12058) <= not a;
    layer4_outputs(12059) <= b;
    layer4_outputs(12060) <= a xor b;
    layer4_outputs(12061) <= not a or b;
    layer4_outputs(12062) <= b and not a;
    layer4_outputs(12063) <= not a;
    layer4_outputs(12064) <= a and b;
    layer4_outputs(12065) <= not a;
    layer4_outputs(12066) <= a and b;
    layer4_outputs(12067) <= a and b;
    layer4_outputs(12068) <= not b;
    layer4_outputs(12069) <= not b or a;
    layer4_outputs(12070) <= not b;
    layer4_outputs(12071) <= '1';
    layer4_outputs(12072) <= '1';
    layer4_outputs(12073) <= a xor b;
    layer4_outputs(12074) <= not b or a;
    layer4_outputs(12075) <= a xor b;
    layer4_outputs(12076) <= not (a xor b);
    layer4_outputs(12077) <= b;
    layer4_outputs(12078) <= a xor b;
    layer4_outputs(12079) <= a or b;
    layer4_outputs(12080) <= not a or b;
    layer4_outputs(12081) <= not (a and b);
    layer4_outputs(12082) <= b;
    layer4_outputs(12083) <= not a or b;
    layer4_outputs(12084) <= b;
    layer4_outputs(12085) <= not b or a;
    layer4_outputs(12086) <= not a;
    layer4_outputs(12087) <= b and not a;
    layer4_outputs(12088) <= a;
    layer4_outputs(12089) <= not a;
    layer4_outputs(12090) <= not a;
    layer4_outputs(12091) <= '0';
    layer4_outputs(12092) <= not b or a;
    layer4_outputs(12093) <= a;
    layer4_outputs(12094) <= a xor b;
    layer4_outputs(12095) <= a and b;
    layer4_outputs(12096) <= not b;
    layer4_outputs(12097) <= b;
    layer4_outputs(12098) <= a and b;
    layer4_outputs(12099) <= a or b;
    layer4_outputs(12100) <= a;
    layer4_outputs(12101) <= not (a or b);
    layer4_outputs(12102) <= a and not b;
    layer4_outputs(12103) <= a and not b;
    layer4_outputs(12104) <= not (a or b);
    layer4_outputs(12105) <= not (a and b);
    layer4_outputs(12106) <= a xor b;
    layer4_outputs(12107) <= '1';
    layer4_outputs(12108) <= a and b;
    layer4_outputs(12109) <= not b or a;
    layer4_outputs(12110) <= not (a or b);
    layer4_outputs(12111) <= not (a xor b);
    layer4_outputs(12112) <= a and not b;
    layer4_outputs(12113) <= not (a and b);
    layer4_outputs(12114) <= not a;
    layer4_outputs(12115) <= a or b;
    layer4_outputs(12116) <= a and b;
    layer4_outputs(12117) <= b and not a;
    layer4_outputs(12118) <= not (a xor b);
    layer4_outputs(12119) <= a and not b;
    layer4_outputs(12120) <= not a;
    layer4_outputs(12121) <= not (a xor b);
    layer4_outputs(12122) <= a xor b;
    layer4_outputs(12123) <= a and not b;
    layer4_outputs(12124) <= b and not a;
    layer4_outputs(12125) <= a and b;
    layer4_outputs(12126) <= not a;
    layer4_outputs(12127) <= a and not b;
    layer4_outputs(12128) <= not b or a;
    layer4_outputs(12129) <= a and not b;
    layer4_outputs(12130) <= not (a or b);
    layer4_outputs(12131) <= not a;
    layer4_outputs(12132) <= b;
    layer4_outputs(12133) <= not a;
    layer4_outputs(12134) <= a or b;
    layer4_outputs(12135) <= not b;
    layer4_outputs(12136) <= not b;
    layer4_outputs(12137) <= '1';
    layer4_outputs(12138) <= a and not b;
    layer4_outputs(12139) <= not b;
    layer4_outputs(12140) <= a and not b;
    layer4_outputs(12141) <= a;
    layer4_outputs(12142) <= a and b;
    layer4_outputs(12143) <= not (a and b);
    layer4_outputs(12144) <= a and not b;
    layer4_outputs(12145) <= not (a or b);
    layer4_outputs(12146) <= not (a xor b);
    layer4_outputs(12147) <= not a;
    layer4_outputs(12148) <= not (a or b);
    layer4_outputs(12149) <= b;
    layer4_outputs(12150) <= not b;
    layer4_outputs(12151) <= not (a or b);
    layer4_outputs(12152) <= not a;
    layer4_outputs(12153) <= b;
    layer4_outputs(12154) <= a and not b;
    layer4_outputs(12155) <= b;
    layer4_outputs(12156) <= not b or a;
    layer4_outputs(12157) <= not b;
    layer4_outputs(12158) <= '0';
    layer4_outputs(12159) <= not (a or b);
    layer4_outputs(12160) <= a;
    layer4_outputs(12161) <= a and not b;
    layer4_outputs(12162) <= not a;
    layer4_outputs(12163) <= a or b;
    layer4_outputs(12164) <= a or b;
    layer4_outputs(12165) <= not (a and b);
    layer4_outputs(12166) <= '0';
    layer4_outputs(12167) <= b;
    layer4_outputs(12168) <= a or b;
    layer4_outputs(12169) <= a or b;
    layer4_outputs(12170) <= a;
    layer4_outputs(12171) <= a;
    layer4_outputs(12172) <= not b or a;
    layer4_outputs(12173) <= b and not a;
    layer4_outputs(12174) <= not a or b;
    layer4_outputs(12175) <= a or b;
    layer4_outputs(12176) <= not a;
    layer4_outputs(12177) <= not b or a;
    layer4_outputs(12178) <= not (a or b);
    layer4_outputs(12179) <= '0';
    layer4_outputs(12180) <= a;
    layer4_outputs(12181) <= not b;
    layer4_outputs(12182) <= b;
    layer4_outputs(12183) <= a or b;
    layer4_outputs(12184) <= a xor b;
    layer4_outputs(12185) <= b;
    layer4_outputs(12186) <= not b or a;
    layer4_outputs(12187) <= a and b;
    layer4_outputs(12188) <= a xor b;
    layer4_outputs(12189) <= not a or b;
    layer4_outputs(12190) <= not (a xor b);
    layer4_outputs(12191) <= not a;
    layer4_outputs(12192) <= not (a and b);
    layer4_outputs(12193) <= a and b;
    layer4_outputs(12194) <= a;
    layer4_outputs(12195) <= not b;
    layer4_outputs(12196) <= a;
    layer4_outputs(12197) <= a;
    layer4_outputs(12198) <= b;
    layer4_outputs(12199) <= b;
    layer4_outputs(12200) <= not (a and b);
    layer4_outputs(12201) <= a and not b;
    layer4_outputs(12202) <= a xor b;
    layer4_outputs(12203) <= not b or a;
    layer4_outputs(12204) <= a xor b;
    layer4_outputs(12205) <= a xor b;
    layer4_outputs(12206) <= b;
    layer4_outputs(12207) <= not (a xor b);
    layer4_outputs(12208) <= a and b;
    layer4_outputs(12209) <= b and not a;
    layer4_outputs(12210) <= b and not a;
    layer4_outputs(12211) <= not b;
    layer4_outputs(12212) <= not a or b;
    layer4_outputs(12213) <= not (a xor b);
    layer4_outputs(12214) <= b;
    layer4_outputs(12215) <= b and not a;
    layer4_outputs(12216) <= b;
    layer4_outputs(12217) <= a or b;
    layer4_outputs(12218) <= a;
    layer4_outputs(12219) <= a and b;
    layer4_outputs(12220) <= not (a xor b);
    layer4_outputs(12221) <= not a or b;
    layer4_outputs(12222) <= not a;
    layer4_outputs(12223) <= not b or a;
    layer4_outputs(12224) <= not (a and b);
    layer4_outputs(12225) <= not (a xor b);
    layer4_outputs(12226) <= not (a and b);
    layer4_outputs(12227) <= a;
    layer4_outputs(12228) <= not a;
    layer4_outputs(12229) <= not a;
    layer4_outputs(12230) <= '1';
    layer4_outputs(12231) <= b;
    layer4_outputs(12232) <= a or b;
    layer4_outputs(12233) <= a xor b;
    layer4_outputs(12234) <= a and not b;
    layer4_outputs(12235) <= not (a xor b);
    layer4_outputs(12236) <= a or b;
    layer4_outputs(12237) <= a;
    layer4_outputs(12238) <= not b;
    layer4_outputs(12239) <= not a;
    layer4_outputs(12240) <= a xor b;
    layer4_outputs(12241) <= a;
    layer4_outputs(12242) <= b and not a;
    layer4_outputs(12243) <= not (a or b);
    layer4_outputs(12244) <= a and b;
    layer4_outputs(12245) <= b;
    layer4_outputs(12246) <= a and not b;
    layer4_outputs(12247) <= a and not b;
    layer4_outputs(12248) <= b;
    layer4_outputs(12249) <= a and b;
    layer4_outputs(12250) <= b and not a;
    layer4_outputs(12251) <= a and b;
    layer4_outputs(12252) <= not b;
    layer4_outputs(12253) <= not (a and b);
    layer4_outputs(12254) <= not (a or b);
    layer4_outputs(12255) <= not a;
    layer4_outputs(12256) <= not (a xor b);
    layer4_outputs(12257) <= not b;
    layer4_outputs(12258) <= not b;
    layer4_outputs(12259) <= not (a or b);
    layer4_outputs(12260) <= a;
    layer4_outputs(12261) <= a or b;
    layer4_outputs(12262) <= b;
    layer4_outputs(12263) <= a;
    layer4_outputs(12264) <= a or b;
    layer4_outputs(12265) <= not (a and b);
    layer4_outputs(12266) <= not b;
    layer4_outputs(12267) <= not b or a;
    layer4_outputs(12268) <= a and b;
    layer4_outputs(12269) <= not b or a;
    layer4_outputs(12270) <= not b;
    layer4_outputs(12271) <= b;
    layer4_outputs(12272) <= not b;
    layer4_outputs(12273) <= b;
    layer4_outputs(12274) <= not b or a;
    layer4_outputs(12275) <= not b or a;
    layer4_outputs(12276) <= not (a or b);
    layer4_outputs(12277) <= not b;
    layer4_outputs(12278) <= a or b;
    layer4_outputs(12279) <= not (a and b);
    layer4_outputs(12280) <= a or b;
    layer4_outputs(12281) <= a and not b;
    layer4_outputs(12282) <= not (a xor b);
    layer4_outputs(12283) <= not b;
    layer4_outputs(12284) <= a;
    layer4_outputs(12285) <= not (a and b);
    layer4_outputs(12286) <= not (a and b);
    layer4_outputs(12287) <= not (a or b);
    layer4_outputs(12288) <= b;
    layer4_outputs(12289) <= a and not b;
    layer4_outputs(12290) <= not a or b;
    layer4_outputs(12291) <= not a;
    layer4_outputs(12292) <= not a or b;
    layer4_outputs(12293) <= not a or b;
    layer4_outputs(12294) <= not b;
    layer4_outputs(12295) <= b;
    layer4_outputs(12296) <= not a or b;
    layer4_outputs(12297) <= not a;
    layer4_outputs(12298) <= a or b;
    layer4_outputs(12299) <= not b;
    layer4_outputs(12300) <= b;
    layer4_outputs(12301) <= b and not a;
    layer4_outputs(12302) <= not a;
    layer4_outputs(12303) <= a or b;
    layer4_outputs(12304) <= not (a xor b);
    layer4_outputs(12305) <= a;
    layer4_outputs(12306) <= b;
    layer4_outputs(12307) <= b and not a;
    layer4_outputs(12308) <= a xor b;
    layer4_outputs(12309) <= a and not b;
    layer4_outputs(12310) <= not a;
    layer4_outputs(12311) <= a and b;
    layer4_outputs(12312) <= a;
    layer4_outputs(12313) <= a;
    layer4_outputs(12314) <= not (a and b);
    layer4_outputs(12315) <= not a or b;
    layer4_outputs(12316) <= a;
    layer4_outputs(12317) <= b;
    layer4_outputs(12318) <= a;
    layer4_outputs(12319) <= not b;
    layer4_outputs(12320) <= '1';
    layer4_outputs(12321) <= not b or a;
    layer4_outputs(12322) <= a;
    layer4_outputs(12323) <= not (a or b);
    layer4_outputs(12324) <= not (a and b);
    layer4_outputs(12325) <= not (a and b);
    layer4_outputs(12326) <= b and not a;
    layer4_outputs(12327) <= a or b;
    layer4_outputs(12328) <= a xor b;
    layer4_outputs(12329) <= a;
    layer4_outputs(12330) <= not b or a;
    layer4_outputs(12331) <= a and not b;
    layer4_outputs(12332) <= a and b;
    layer4_outputs(12333) <= b;
    layer4_outputs(12334) <= b;
    layer4_outputs(12335) <= not b;
    layer4_outputs(12336) <= a xor b;
    layer4_outputs(12337) <= not a or b;
    layer4_outputs(12338) <= not (a or b);
    layer4_outputs(12339) <= not (a and b);
    layer4_outputs(12340) <= a and not b;
    layer4_outputs(12341) <= not (a and b);
    layer4_outputs(12342) <= a and not b;
    layer4_outputs(12343) <= not (a and b);
    layer4_outputs(12344) <= not b;
    layer4_outputs(12345) <= a xor b;
    layer4_outputs(12346) <= not b;
    layer4_outputs(12347) <= not a or b;
    layer4_outputs(12348) <= a and b;
    layer4_outputs(12349) <= not (a or b);
    layer4_outputs(12350) <= not a or b;
    layer4_outputs(12351) <= not (a or b);
    layer4_outputs(12352) <= not a;
    layer4_outputs(12353) <= a and not b;
    layer4_outputs(12354) <= a and b;
    layer4_outputs(12355) <= not (a xor b);
    layer4_outputs(12356) <= a xor b;
    layer4_outputs(12357) <= not a;
    layer4_outputs(12358) <= not a;
    layer4_outputs(12359) <= b;
    layer4_outputs(12360) <= b and not a;
    layer4_outputs(12361) <= a xor b;
    layer4_outputs(12362) <= not (a and b);
    layer4_outputs(12363) <= a xor b;
    layer4_outputs(12364) <= not a;
    layer4_outputs(12365) <= a;
    layer4_outputs(12366) <= not a or b;
    layer4_outputs(12367) <= b and not a;
    layer4_outputs(12368) <= not a or b;
    layer4_outputs(12369) <= not (a and b);
    layer4_outputs(12370) <= '0';
    layer4_outputs(12371) <= b and not a;
    layer4_outputs(12372) <= '0';
    layer4_outputs(12373) <= b;
    layer4_outputs(12374) <= not b or a;
    layer4_outputs(12375) <= not a or b;
    layer4_outputs(12376) <= not b or a;
    layer4_outputs(12377) <= not (a and b);
    layer4_outputs(12378) <= not (a and b);
    layer4_outputs(12379) <= not (a xor b);
    layer4_outputs(12380) <= not b;
    layer4_outputs(12381) <= not a or b;
    layer4_outputs(12382) <= not (a and b);
    layer4_outputs(12383) <= a;
    layer4_outputs(12384) <= a and not b;
    layer4_outputs(12385) <= '0';
    layer4_outputs(12386) <= b and not a;
    layer4_outputs(12387) <= b;
    layer4_outputs(12388) <= not a;
    layer4_outputs(12389) <= not (a and b);
    layer4_outputs(12390) <= '1';
    layer4_outputs(12391) <= not a or b;
    layer4_outputs(12392) <= a and not b;
    layer4_outputs(12393) <= not a or b;
    layer4_outputs(12394) <= not a;
    layer4_outputs(12395) <= not b;
    layer4_outputs(12396) <= not a or b;
    layer4_outputs(12397) <= not b;
    layer4_outputs(12398) <= a or b;
    layer4_outputs(12399) <= a;
    layer4_outputs(12400) <= not (a xor b);
    layer4_outputs(12401) <= a and not b;
    layer4_outputs(12402) <= not (a and b);
    layer4_outputs(12403) <= not b;
    layer4_outputs(12404) <= not a;
    layer4_outputs(12405) <= not a;
    layer4_outputs(12406) <= a xor b;
    layer4_outputs(12407) <= not a or b;
    layer4_outputs(12408) <= a and b;
    layer4_outputs(12409) <= b;
    layer4_outputs(12410) <= a;
    layer4_outputs(12411) <= not (a or b);
    layer4_outputs(12412) <= not b;
    layer4_outputs(12413) <= '0';
    layer4_outputs(12414) <= not b;
    layer4_outputs(12415) <= a;
    layer4_outputs(12416) <= not (a or b);
    layer4_outputs(12417) <= not b;
    layer4_outputs(12418) <= b and not a;
    layer4_outputs(12419) <= a;
    layer4_outputs(12420) <= not a;
    layer4_outputs(12421) <= a;
    layer4_outputs(12422) <= not b;
    layer4_outputs(12423) <= not (a and b);
    layer4_outputs(12424) <= not b;
    layer4_outputs(12425) <= b;
    layer4_outputs(12426) <= b and not a;
    layer4_outputs(12427) <= not b;
    layer4_outputs(12428) <= not a or b;
    layer4_outputs(12429) <= not (a and b);
    layer4_outputs(12430) <= not b or a;
    layer4_outputs(12431) <= b and not a;
    layer4_outputs(12432) <= not b;
    layer4_outputs(12433) <= a;
    layer4_outputs(12434) <= not (a xor b);
    layer4_outputs(12435) <= not (a xor b);
    layer4_outputs(12436) <= not (a or b);
    layer4_outputs(12437) <= a;
    layer4_outputs(12438) <= not a or b;
    layer4_outputs(12439) <= not (a and b);
    layer4_outputs(12440) <= b;
    layer4_outputs(12441) <= not a;
    layer4_outputs(12442) <= b;
    layer4_outputs(12443) <= a and b;
    layer4_outputs(12444) <= not (a or b);
    layer4_outputs(12445) <= not b or a;
    layer4_outputs(12446) <= not a;
    layer4_outputs(12447) <= b;
    layer4_outputs(12448) <= not (a or b);
    layer4_outputs(12449) <= b;
    layer4_outputs(12450) <= a and not b;
    layer4_outputs(12451) <= not b;
    layer4_outputs(12452) <= not b or a;
    layer4_outputs(12453) <= not b;
    layer4_outputs(12454) <= a;
    layer4_outputs(12455) <= not b;
    layer4_outputs(12456) <= not a or b;
    layer4_outputs(12457) <= b and not a;
    layer4_outputs(12458) <= not (a or b);
    layer4_outputs(12459) <= a;
    layer4_outputs(12460) <= not a;
    layer4_outputs(12461) <= b;
    layer4_outputs(12462) <= a and b;
    layer4_outputs(12463) <= a or b;
    layer4_outputs(12464) <= not a;
    layer4_outputs(12465) <= a;
    layer4_outputs(12466) <= not a or b;
    layer4_outputs(12467) <= not b or a;
    layer4_outputs(12468) <= not (a xor b);
    layer4_outputs(12469) <= b and not a;
    layer4_outputs(12470) <= a and not b;
    layer4_outputs(12471) <= not a;
    layer4_outputs(12472) <= '1';
    layer4_outputs(12473) <= not (a or b);
    layer4_outputs(12474) <= a;
    layer4_outputs(12475) <= a;
    layer4_outputs(12476) <= a and not b;
    layer4_outputs(12477) <= not a;
    layer4_outputs(12478) <= a;
    layer4_outputs(12479) <= a;
    layer4_outputs(12480) <= not (a xor b);
    layer4_outputs(12481) <= b;
    layer4_outputs(12482) <= not b;
    layer4_outputs(12483) <= not (a and b);
    layer4_outputs(12484) <= a and not b;
    layer4_outputs(12485) <= b;
    layer4_outputs(12486) <= a and not b;
    layer4_outputs(12487) <= a;
    layer4_outputs(12488) <= not (a or b);
    layer4_outputs(12489) <= b;
    layer4_outputs(12490) <= not a or b;
    layer4_outputs(12491) <= not (a and b);
    layer4_outputs(12492) <= a;
    layer4_outputs(12493) <= not b;
    layer4_outputs(12494) <= '1';
    layer4_outputs(12495) <= not (a or b);
    layer4_outputs(12496) <= not (a or b);
    layer4_outputs(12497) <= a;
    layer4_outputs(12498) <= b;
    layer4_outputs(12499) <= not a;
    layer4_outputs(12500) <= b;
    layer4_outputs(12501) <= not a;
    layer4_outputs(12502) <= not a;
    layer4_outputs(12503) <= b and not a;
    layer4_outputs(12504) <= not b;
    layer4_outputs(12505) <= not (a and b);
    layer4_outputs(12506) <= not a;
    layer4_outputs(12507) <= '0';
    layer4_outputs(12508) <= a;
    layer4_outputs(12509) <= '0';
    layer4_outputs(12510) <= a and not b;
    layer4_outputs(12511) <= not a;
    layer4_outputs(12512) <= a;
    layer4_outputs(12513) <= not b or a;
    layer4_outputs(12514) <= a and not b;
    layer4_outputs(12515) <= not (a xor b);
    layer4_outputs(12516) <= not a;
    layer4_outputs(12517) <= a and not b;
    layer4_outputs(12518) <= b;
    layer4_outputs(12519) <= not a;
    layer4_outputs(12520) <= not (a and b);
    layer4_outputs(12521) <= not b;
    layer4_outputs(12522) <= not a;
    layer4_outputs(12523) <= not a;
    layer4_outputs(12524) <= b;
    layer4_outputs(12525) <= not (a xor b);
    layer4_outputs(12526) <= b and not a;
    layer4_outputs(12527) <= a and b;
    layer4_outputs(12528) <= not a or b;
    layer4_outputs(12529) <= a and b;
    layer4_outputs(12530) <= a and not b;
    layer4_outputs(12531) <= not (a xor b);
    layer4_outputs(12532) <= a;
    layer4_outputs(12533) <= not (a and b);
    layer4_outputs(12534) <= not a;
    layer4_outputs(12535) <= not a;
    layer4_outputs(12536) <= not b;
    layer4_outputs(12537) <= b;
    layer4_outputs(12538) <= not a;
    layer4_outputs(12539) <= a;
    layer4_outputs(12540) <= a;
    layer4_outputs(12541) <= not a;
    layer4_outputs(12542) <= not a;
    layer4_outputs(12543) <= not a;
    layer4_outputs(12544) <= a and b;
    layer4_outputs(12545) <= a;
    layer4_outputs(12546) <= a and not b;
    layer4_outputs(12547) <= a;
    layer4_outputs(12548) <= not (a xor b);
    layer4_outputs(12549) <= not b;
    layer4_outputs(12550) <= '0';
    layer4_outputs(12551) <= not b;
    layer4_outputs(12552) <= not (a xor b);
    layer4_outputs(12553) <= not (a or b);
    layer4_outputs(12554) <= not b or a;
    layer4_outputs(12555) <= a and b;
    layer4_outputs(12556) <= b;
    layer4_outputs(12557) <= a;
    layer4_outputs(12558) <= not a;
    layer4_outputs(12559) <= not b or a;
    layer4_outputs(12560) <= not b;
    layer4_outputs(12561) <= a or b;
    layer4_outputs(12562) <= not a;
    layer4_outputs(12563) <= not a or b;
    layer4_outputs(12564) <= not (a xor b);
    layer4_outputs(12565) <= b;
    layer4_outputs(12566) <= not a or b;
    layer4_outputs(12567) <= not (a and b);
    layer4_outputs(12568) <= not a or b;
    layer4_outputs(12569) <= not (a and b);
    layer4_outputs(12570) <= a and b;
    layer4_outputs(12571) <= a;
    layer4_outputs(12572) <= a and b;
    layer4_outputs(12573) <= not (a or b);
    layer4_outputs(12574) <= a or b;
    layer4_outputs(12575) <= not b or a;
    layer4_outputs(12576) <= not a;
    layer4_outputs(12577) <= a or b;
    layer4_outputs(12578) <= a;
    layer4_outputs(12579) <= not a or b;
    layer4_outputs(12580) <= not (a and b);
    layer4_outputs(12581) <= not b or a;
    layer4_outputs(12582) <= b;
    layer4_outputs(12583) <= not a or b;
    layer4_outputs(12584) <= b;
    layer4_outputs(12585) <= not (a xor b);
    layer4_outputs(12586) <= not a;
    layer4_outputs(12587) <= not (a xor b);
    layer4_outputs(12588) <= b;
    layer4_outputs(12589) <= not (a or b);
    layer4_outputs(12590) <= not (a and b);
    layer4_outputs(12591) <= a and b;
    layer4_outputs(12592) <= not b or a;
    layer4_outputs(12593) <= b and not a;
    layer4_outputs(12594) <= a and not b;
    layer4_outputs(12595) <= not (a and b);
    layer4_outputs(12596) <= not a;
    layer4_outputs(12597) <= b and not a;
    layer4_outputs(12598) <= not b;
    layer4_outputs(12599) <= not a or b;
    layer4_outputs(12600) <= not (a and b);
    layer4_outputs(12601) <= not (a or b);
    layer4_outputs(12602) <= not a or b;
    layer4_outputs(12603) <= not a;
    layer4_outputs(12604) <= a and not b;
    layer4_outputs(12605) <= not a;
    layer4_outputs(12606) <= b and not a;
    layer4_outputs(12607) <= b;
    layer4_outputs(12608) <= not b;
    layer4_outputs(12609) <= not b;
    layer4_outputs(12610) <= not (a and b);
    layer4_outputs(12611) <= b;
    layer4_outputs(12612) <= not a;
    layer4_outputs(12613) <= not a;
    layer4_outputs(12614) <= a xor b;
    layer4_outputs(12615) <= not b;
    layer4_outputs(12616) <= not (a or b);
    layer4_outputs(12617) <= a xor b;
    layer4_outputs(12618) <= a and not b;
    layer4_outputs(12619) <= not b or a;
    layer4_outputs(12620) <= not (a or b);
    layer4_outputs(12621) <= not a or b;
    layer4_outputs(12622) <= not a;
    layer4_outputs(12623) <= b and not a;
    layer4_outputs(12624) <= a and b;
    layer4_outputs(12625) <= a;
    layer4_outputs(12626) <= a;
    layer4_outputs(12627) <= not b or a;
    layer4_outputs(12628) <= a;
    layer4_outputs(12629) <= not b;
    layer4_outputs(12630) <= a;
    layer4_outputs(12631) <= not (a and b);
    layer4_outputs(12632) <= b and not a;
    layer4_outputs(12633) <= not (a or b);
    layer4_outputs(12634) <= a;
    layer4_outputs(12635) <= not b;
    layer4_outputs(12636) <= not (a or b);
    layer4_outputs(12637) <= a xor b;
    layer4_outputs(12638) <= not (a and b);
    layer4_outputs(12639) <= a and b;
    layer4_outputs(12640) <= a and not b;
    layer4_outputs(12641) <= not (a and b);
    layer4_outputs(12642) <= not (a or b);
    layer4_outputs(12643) <= '0';
    layer4_outputs(12644) <= b and not a;
    layer4_outputs(12645) <= not a;
    layer4_outputs(12646) <= a xor b;
    layer4_outputs(12647) <= not a;
    layer4_outputs(12648) <= a and b;
    layer4_outputs(12649) <= b and not a;
    layer4_outputs(12650) <= b;
    layer4_outputs(12651) <= b;
    layer4_outputs(12652) <= not (a and b);
    layer4_outputs(12653) <= not (a xor b);
    layer4_outputs(12654) <= a and b;
    layer4_outputs(12655) <= not b or a;
    layer4_outputs(12656) <= a;
    layer4_outputs(12657) <= a;
    layer4_outputs(12658) <= not b;
    layer4_outputs(12659) <= not (a or b);
    layer4_outputs(12660) <= not b;
    layer4_outputs(12661) <= not a or b;
    layer4_outputs(12662) <= not (a and b);
    layer4_outputs(12663) <= b;
    layer4_outputs(12664) <= a and not b;
    layer4_outputs(12665) <= not a;
    layer4_outputs(12666) <= not (a or b);
    layer4_outputs(12667) <= not (a xor b);
    layer4_outputs(12668) <= a and b;
    layer4_outputs(12669) <= a and b;
    layer4_outputs(12670) <= a;
    layer4_outputs(12671) <= not b;
    layer4_outputs(12672) <= b;
    layer4_outputs(12673) <= a and not b;
    layer4_outputs(12674) <= not b;
    layer4_outputs(12675) <= '1';
    layer4_outputs(12676) <= a xor b;
    layer4_outputs(12677) <= not a;
    layer4_outputs(12678) <= a xor b;
    layer4_outputs(12679) <= b;
    layer4_outputs(12680) <= not (a and b);
    layer4_outputs(12681) <= b;
    layer4_outputs(12682) <= not a or b;
    layer4_outputs(12683) <= not b;
    layer4_outputs(12684) <= not b or a;
    layer4_outputs(12685) <= a and b;
    layer4_outputs(12686) <= not b;
    layer4_outputs(12687) <= not (a xor b);
    layer4_outputs(12688) <= a xor b;
    layer4_outputs(12689) <= a and b;
    layer4_outputs(12690) <= not (a xor b);
    layer4_outputs(12691) <= not (a and b);
    layer4_outputs(12692) <= a and b;
    layer4_outputs(12693) <= not b;
    layer4_outputs(12694) <= b;
    layer4_outputs(12695) <= not b;
    layer4_outputs(12696) <= not a;
    layer4_outputs(12697) <= a and b;
    layer4_outputs(12698) <= not a;
    layer4_outputs(12699) <= a;
    layer4_outputs(12700) <= not a;
    layer4_outputs(12701) <= a xor b;
    layer4_outputs(12702) <= not (a and b);
    layer4_outputs(12703) <= not (a or b);
    layer4_outputs(12704) <= a and not b;
    layer4_outputs(12705) <= not b;
    layer4_outputs(12706) <= not a;
    layer4_outputs(12707) <= not a;
    layer4_outputs(12708) <= a and not b;
    layer4_outputs(12709) <= not b;
    layer4_outputs(12710) <= not a or b;
    layer4_outputs(12711) <= not (a or b);
    layer4_outputs(12712) <= not b or a;
    layer4_outputs(12713) <= not (a and b);
    layer4_outputs(12714) <= a;
    layer4_outputs(12715) <= not a or b;
    layer4_outputs(12716) <= not a or b;
    layer4_outputs(12717) <= not a;
    layer4_outputs(12718) <= b and not a;
    layer4_outputs(12719) <= b and not a;
    layer4_outputs(12720) <= not (a xor b);
    layer4_outputs(12721) <= a and b;
    layer4_outputs(12722) <= b;
    layer4_outputs(12723) <= not a or b;
    layer4_outputs(12724) <= a;
    layer4_outputs(12725) <= not b;
    layer4_outputs(12726) <= not (a and b);
    layer4_outputs(12727) <= a;
    layer4_outputs(12728) <= not b;
    layer4_outputs(12729) <= b;
    layer4_outputs(12730) <= a and b;
    layer4_outputs(12731) <= not a or b;
    layer4_outputs(12732) <= b;
    layer4_outputs(12733) <= not (a and b);
    layer4_outputs(12734) <= not a or b;
    layer4_outputs(12735) <= not a or b;
    layer4_outputs(12736) <= not b or a;
    layer4_outputs(12737) <= not a;
    layer4_outputs(12738) <= a xor b;
    layer4_outputs(12739) <= '0';
    layer4_outputs(12740) <= a;
    layer4_outputs(12741) <= not a;
    layer4_outputs(12742) <= a and b;
    layer4_outputs(12743) <= not (a or b);
    layer4_outputs(12744) <= a xor b;
    layer4_outputs(12745) <= not a;
    layer4_outputs(12746) <= not b;
    layer4_outputs(12747) <= a;
    layer4_outputs(12748) <= b;
    layer4_outputs(12749) <= b;
    layer4_outputs(12750) <= not (a and b);
    layer4_outputs(12751) <= not a;
    layer4_outputs(12752) <= '0';
    layer4_outputs(12753) <= not (a or b);
    layer4_outputs(12754) <= a or b;
    layer4_outputs(12755) <= not (a xor b);
    layer4_outputs(12756) <= b and not a;
    layer4_outputs(12757) <= not b;
    layer4_outputs(12758) <= '0';
    layer4_outputs(12759) <= not (a xor b);
    layer4_outputs(12760) <= a or b;
    layer4_outputs(12761) <= a or b;
    layer4_outputs(12762) <= a;
    layer4_outputs(12763) <= not b;
    layer4_outputs(12764) <= not b;
    layer4_outputs(12765) <= a xor b;
    layer4_outputs(12766) <= a and not b;
    layer4_outputs(12767) <= a xor b;
    layer4_outputs(12768) <= not a;
    layer4_outputs(12769) <= b;
    layer4_outputs(12770) <= b and not a;
    layer4_outputs(12771) <= a;
    layer4_outputs(12772) <= a;
    layer4_outputs(12773) <= a xor b;
    layer4_outputs(12774) <= not b or a;
    layer4_outputs(12775) <= a and not b;
    layer4_outputs(12776) <= a xor b;
    layer4_outputs(12777) <= a and not b;
    layer4_outputs(12778) <= not b or a;
    layer4_outputs(12779) <= b;
    layer4_outputs(12780) <= b;
    layer4_outputs(12781) <= not (a and b);
    layer4_outputs(12782) <= not (a xor b);
    layer4_outputs(12783) <= b and not a;
    layer4_outputs(12784) <= a or b;
    layer4_outputs(12785) <= a and b;
    layer4_outputs(12786) <= not a or b;
    layer4_outputs(12787) <= a;
    layer4_outputs(12788) <= a and not b;
    layer4_outputs(12789) <= not (a or b);
    layer4_outputs(12790) <= a and not b;
    layer4_outputs(12791) <= a xor b;
    layer4_outputs(12792) <= b;
    layer4_outputs(12793) <= not (a or b);
    layer4_outputs(12794) <= not a;
    layer4_outputs(12795) <= b;
    layer4_outputs(12796) <= not (a xor b);
    layer4_outputs(12797) <= b;
    layer4_outputs(12798) <= a;
    layer4_outputs(12799) <= not (a or b);
    layer5_outputs(0) <= a;
    layer5_outputs(1) <= not a or b;
    layer5_outputs(2) <= not b or a;
    layer5_outputs(3) <= not b;
    layer5_outputs(4) <= '1';
    layer5_outputs(5) <= a and b;
    layer5_outputs(6) <= not a;
    layer5_outputs(7) <= not a;
    layer5_outputs(8) <= b;
    layer5_outputs(9) <= a;
    layer5_outputs(10) <= not b;
    layer5_outputs(11) <= not (a and b);
    layer5_outputs(12) <= b;
    layer5_outputs(13) <= b;
    layer5_outputs(14) <= a xor b;
    layer5_outputs(15) <= '0';
    layer5_outputs(16) <= a and b;
    layer5_outputs(17) <= a;
    layer5_outputs(18) <= b;
    layer5_outputs(19) <= not (a xor b);
    layer5_outputs(20) <= not b;
    layer5_outputs(21) <= a;
    layer5_outputs(22) <= not a;
    layer5_outputs(23) <= a and b;
    layer5_outputs(24) <= a and not b;
    layer5_outputs(25) <= b;
    layer5_outputs(26) <= a;
    layer5_outputs(27) <= b and not a;
    layer5_outputs(28) <= a;
    layer5_outputs(29) <= not a or b;
    layer5_outputs(30) <= b;
    layer5_outputs(31) <= not b or a;
    layer5_outputs(32) <= not a;
    layer5_outputs(33) <= not b;
    layer5_outputs(34) <= b;
    layer5_outputs(35) <= not a;
    layer5_outputs(36) <= not a;
    layer5_outputs(37) <= b and not a;
    layer5_outputs(38) <= a and not b;
    layer5_outputs(39) <= not (a and b);
    layer5_outputs(40) <= a or b;
    layer5_outputs(41) <= b;
    layer5_outputs(42) <= a or b;
    layer5_outputs(43) <= b;
    layer5_outputs(44) <= a and not b;
    layer5_outputs(45) <= not a;
    layer5_outputs(46) <= a;
    layer5_outputs(47) <= a and not b;
    layer5_outputs(48) <= a;
    layer5_outputs(49) <= not (a and b);
    layer5_outputs(50) <= a;
    layer5_outputs(51) <= not a;
    layer5_outputs(52) <= not a;
    layer5_outputs(53) <= b and not a;
    layer5_outputs(54) <= not (a xor b);
    layer5_outputs(55) <= not (a and b);
    layer5_outputs(56) <= not (a xor b);
    layer5_outputs(57) <= a;
    layer5_outputs(58) <= not b or a;
    layer5_outputs(59) <= not (a or b);
    layer5_outputs(60) <= not (a and b);
    layer5_outputs(61) <= a;
    layer5_outputs(62) <= a and b;
    layer5_outputs(63) <= a or b;
    layer5_outputs(64) <= a;
    layer5_outputs(65) <= a and not b;
    layer5_outputs(66) <= a xor b;
    layer5_outputs(67) <= b;
    layer5_outputs(68) <= not a;
    layer5_outputs(69) <= a xor b;
    layer5_outputs(70) <= not (a xor b);
    layer5_outputs(71) <= a or b;
    layer5_outputs(72) <= a;
    layer5_outputs(73) <= a xor b;
    layer5_outputs(74) <= b and not a;
    layer5_outputs(75) <= a or b;
    layer5_outputs(76) <= not a;
    layer5_outputs(77) <= not a;
    layer5_outputs(78) <= b and not a;
    layer5_outputs(79) <= not (a and b);
    layer5_outputs(80) <= not a;
    layer5_outputs(81) <= not (a or b);
    layer5_outputs(82) <= not (a xor b);
    layer5_outputs(83) <= a;
    layer5_outputs(84) <= not (a xor b);
    layer5_outputs(85) <= not a;
    layer5_outputs(86) <= not (a xor b);
    layer5_outputs(87) <= a xor b;
    layer5_outputs(88) <= a and not b;
    layer5_outputs(89) <= not a or b;
    layer5_outputs(90) <= not (a xor b);
    layer5_outputs(91) <= not (a xor b);
    layer5_outputs(92) <= '0';
    layer5_outputs(93) <= not a;
    layer5_outputs(94) <= a xor b;
    layer5_outputs(95) <= not a;
    layer5_outputs(96) <= not b;
    layer5_outputs(97) <= not (a and b);
    layer5_outputs(98) <= not a or b;
    layer5_outputs(99) <= not b;
    layer5_outputs(100) <= not b or a;
    layer5_outputs(101) <= b;
    layer5_outputs(102) <= a and b;
    layer5_outputs(103) <= a or b;
    layer5_outputs(104) <= b and not a;
    layer5_outputs(105) <= b;
    layer5_outputs(106) <= b;
    layer5_outputs(107) <= b and not a;
    layer5_outputs(108) <= a;
    layer5_outputs(109) <= b;
    layer5_outputs(110) <= a;
    layer5_outputs(111) <= a;
    layer5_outputs(112) <= a xor b;
    layer5_outputs(113) <= a xor b;
    layer5_outputs(114) <= not b;
    layer5_outputs(115) <= b;
    layer5_outputs(116) <= a;
    layer5_outputs(117) <= b and not a;
    layer5_outputs(118) <= a;
    layer5_outputs(119) <= a;
    layer5_outputs(120) <= not (a xor b);
    layer5_outputs(121) <= a and not b;
    layer5_outputs(122) <= not a or b;
    layer5_outputs(123) <= not a;
    layer5_outputs(124) <= not b;
    layer5_outputs(125) <= a and not b;
    layer5_outputs(126) <= not (a and b);
    layer5_outputs(127) <= a xor b;
    layer5_outputs(128) <= b and not a;
    layer5_outputs(129) <= a and not b;
    layer5_outputs(130) <= b and not a;
    layer5_outputs(131) <= not b;
    layer5_outputs(132) <= not b;
    layer5_outputs(133) <= a;
    layer5_outputs(134) <= b;
    layer5_outputs(135) <= not a or b;
    layer5_outputs(136) <= not a;
    layer5_outputs(137) <= a xor b;
    layer5_outputs(138) <= b and not a;
    layer5_outputs(139) <= not b;
    layer5_outputs(140) <= b;
    layer5_outputs(141) <= a xor b;
    layer5_outputs(142) <= b and not a;
    layer5_outputs(143) <= not b or a;
    layer5_outputs(144) <= b;
    layer5_outputs(145) <= b and not a;
    layer5_outputs(146) <= a xor b;
    layer5_outputs(147) <= b;
    layer5_outputs(148) <= not (a and b);
    layer5_outputs(149) <= a and not b;
    layer5_outputs(150) <= b;
    layer5_outputs(151) <= not a;
    layer5_outputs(152) <= b and not a;
    layer5_outputs(153) <= a;
    layer5_outputs(154) <= not b;
    layer5_outputs(155) <= a;
    layer5_outputs(156) <= b;
    layer5_outputs(157) <= b;
    layer5_outputs(158) <= a;
    layer5_outputs(159) <= a;
    layer5_outputs(160) <= a;
    layer5_outputs(161) <= not b;
    layer5_outputs(162) <= a xor b;
    layer5_outputs(163) <= not b;
    layer5_outputs(164) <= a and b;
    layer5_outputs(165) <= a and b;
    layer5_outputs(166) <= not a;
    layer5_outputs(167) <= not (a and b);
    layer5_outputs(168) <= not b;
    layer5_outputs(169) <= a or b;
    layer5_outputs(170) <= a xor b;
    layer5_outputs(171) <= b;
    layer5_outputs(172) <= not a;
    layer5_outputs(173) <= not (a xor b);
    layer5_outputs(174) <= not a;
    layer5_outputs(175) <= b;
    layer5_outputs(176) <= not a or b;
    layer5_outputs(177) <= a xor b;
    layer5_outputs(178) <= a;
    layer5_outputs(179) <= not b or a;
    layer5_outputs(180) <= not a;
    layer5_outputs(181) <= a and not b;
    layer5_outputs(182) <= not a;
    layer5_outputs(183) <= a and not b;
    layer5_outputs(184) <= not a;
    layer5_outputs(185) <= b;
    layer5_outputs(186) <= b;
    layer5_outputs(187) <= not b;
    layer5_outputs(188) <= not b;
    layer5_outputs(189) <= b and not a;
    layer5_outputs(190) <= a;
    layer5_outputs(191) <= not a or b;
    layer5_outputs(192) <= not a or b;
    layer5_outputs(193) <= a and not b;
    layer5_outputs(194) <= not (a and b);
    layer5_outputs(195) <= not b or a;
    layer5_outputs(196) <= b and not a;
    layer5_outputs(197) <= not b or a;
    layer5_outputs(198) <= '0';
    layer5_outputs(199) <= not a;
    layer5_outputs(200) <= not (a or b);
    layer5_outputs(201) <= not (a and b);
    layer5_outputs(202) <= not a;
    layer5_outputs(203) <= not b or a;
    layer5_outputs(204) <= not b;
    layer5_outputs(205) <= a;
    layer5_outputs(206) <= not b;
    layer5_outputs(207) <= b and not a;
    layer5_outputs(208) <= b and not a;
    layer5_outputs(209) <= not a;
    layer5_outputs(210) <= not b;
    layer5_outputs(211) <= not b;
    layer5_outputs(212) <= b;
    layer5_outputs(213) <= not b;
    layer5_outputs(214) <= a xor b;
    layer5_outputs(215) <= not b or a;
    layer5_outputs(216) <= not (a xor b);
    layer5_outputs(217) <= a xor b;
    layer5_outputs(218) <= not b;
    layer5_outputs(219) <= not b;
    layer5_outputs(220) <= b;
    layer5_outputs(221) <= a;
    layer5_outputs(222) <= not b or a;
    layer5_outputs(223) <= not b;
    layer5_outputs(224) <= a or b;
    layer5_outputs(225) <= not a;
    layer5_outputs(226) <= not b or a;
    layer5_outputs(227) <= not (a xor b);
    layer5_outputs(228) <= a xor b;
    layer5_outputs(229) <= not b or a;
    layer5_outputs(230) <= not (a and b);
    layer5_outputs(231) <= a or b;
    layer5_outputs(232) <= not a;
    layer5_outputs(233) <= a;
    layer5_outputs(234) <= '1';
    layer5_outputs(235) <= b;
    layer5_outputs(236) <= not b or a;
    layer5_outputs(237) <= not b;
    layer5_outputs(238) <= not b or a;
    layer5_outputs(239) <= not b or a;
    layer5_outputs(240) <= not b;
    layer5_outputs(241) <= not b;
    layer5_outputs(242) <= not (a and b);
    layer5_outputs(243) <= a and not b;
    layer5_outputs(244) <= b;
    layer5_outputs(245) <= not a;
    layer5_outputs(246) <= not b;
    layer5_outputs(247) <= b and not a;
    layer5_outputs(248) <= a;
    layer5_outputs(249) <= not a;
    layer5_outputs(250) <= b;
    layer5_outputs(251) <= not (a xor b);
    layer5_outputs(252) <= not a;
    layer5_outputs(253) <= not (a and b);
    layer5_outputs(254) <= not a;
    layer5_outputs(255) <= '1';
    layer5_outputs(256) <= not a;
    layer5_outputs(257) <= not (a and b);
    layer5_outputs(258) <= not b;
    layer5_outputs(259) <= a and b;
    layer5_outputs(260) <= not (a xor b);
    layer5_outputs(261) <= not b;
    layer5_outputs(262) <= not a;
    layer5_outputs(263) <= not b or a;
    layer5_outputs(264) <= b;
    layer5_outputs(265) <= b;
    layer5_outputs(266) <= a and b;
    layer5_outputs(267) <= a;
    layer5_outputs(268) <= not a;
    layer5_outputs(269) <= not b;
    layer5_outputs(270) <= a;
    layer5_outputs(271) <= b and not a;
    layer5_outputs(272) <= a and not b;
    layer5_outputs(273) <= a or b;
    layer5_outputs(274) <= not a or b;
    layer5_outputs(275) <= a;
    layer5_outputs(276) <= a;
    layer5_outputs(277) <= a or b;
    layer5_outputs(278) <= not b or a;
    layer5_outputs(279) <= not (a and b);
    layer5_outputs(280) <= a;
    layer5_outputs(281) <= b and not a;
    layer5_outputs(282) <= not a;
    layer5_outputs(283) <= a and not b;
    layer5_outputs(284) <= not a or b;
    layer5_outputs(285) <= a xor b;
    layer5_outputs(286) <= b;
    layer5_outputs(287) <= not (a xor b);
    layer5_outputs(288) <= a and b;
    layer5_outputs(289) <= not (a xor b);
    layer5_outputs(290) <= a and not b;
    layer5_outputs(291) <= not (a xor b);
    layer5_outputs(292) <= a and not b;
    layer5_outputs(293) <= a;
    layer5_outputs(294) <= b and not a;
    layer5_outputs(295) <= b;
    layer5_outputs(296) <= not b;
    layer5_outputs(297) <= '0';
    layer5_outputs(298) <= not b;
    layer5_outputs(299) <= a;
    layer5_outputs(300) <= a;
    layer5_outputs(301) <= b;
    layer5_outputs(302) <= not (a and b);
    layer5_outputs(303) <= b;
    layer5_outputs(304) <= a and not b;
    layer5_outputs(305) <= not a;
    layer5_outputs(306) <= not (a xor b);
    layer5_outputs(307) <= '1';
    layer5_outputs(308) <= not b;
    layer5_outputs(309) <= not a or b;
    layer5_outputs(310) <= not (a xor b);
    layer5_outputs(311) <= not a;
    layer5_outputs(312) <= a;
    layer5_outputs(313) <= b;
    layer5_outputs(314) <= b;
    layer5_outputs(315) <= a xor b;
    layer5_outputs(316) <= not a or b;
    layer5_outputs(317) <= a and b;
    layer5_outputs(318) <= b and not a;
    layer5_outputs(319) <= not (a xor b);
    layer5_outputs(320) <= not b;
    layer5_outputs(321) <= not a;
    layer5_outputs(322) <= b;
    layer5_outputs(323) <= not b or a;
    layer5_outputs(324) <= not (a xor b);
    layer5_outputs(325) <= a;
    layer5_outputs(326) <= not b;
    layer5_outputs(327) <= b;
    layer5_outputs(328) <= not b;
    layer5_outputs(329) <= not (a and b);
    layer5_outputs(330) <= not b or a;
    layer5_outputs(331) <= not b;
    layer5_outputs(332) <= not a or b;
    layer5_outputs(333) <= b;
    layer5_outputs(334) <= a and not b;
    layer5_outputs(335) <= not b or a;
    layer5_outputs(336) <= '0';
    layer5_outputs(337) <= a;
    layer5_outputs(338) <= not a;
    layer5_outputs(339) <= not a;
    layer5_outputs(340) <= not a;
    layer5_outputs(341) <= a;
    layer5_outputs(342) <= b;
    layer5_outputs(343) <= a;
    layer5_outputs(344) <= a;
    layer5_outputs(345) <= not b;
    layer5_outputs(346) <= a or b;
    layer5_outputs(347) <= b;
    layer5_outputs(348) <= not (a or b);
    layer5_outputs(349) <= not b or a;
    layer5_outputs(350) <= b;
    layer5_outputs(351) <= not a;
    layer5_outputs(352) <= not b;
    layer5_outputs(353) <= not a or b;
    layer5_outputs(354) <= '0';
    layer5_outputs(355) <= not a;
    layer5_outputs(356) <= a or b;
    layer5_outputs(357) <= a;
    layer5_outputs(358) <= b;
    layer5_outputs(359) <= a;
    layer5_outputs(360) <= not a;
    layer5_outputs(361) <= not (a xor b);
    layer5_outputs(362) <= not a;
    layer5_outputs(363) <= not a or b;
    layer5_outputs(364) <= b;
    layer5_outputs(365) <= not a;
    layer5_outputs(366) <= b;
    layer5_outputs(367) <= a and b;
    layer5_outputs(368) <= not a or b;
    layer5_outputs(369) <= not (a xor b);
    layer5_outputs(370) <= not a or b;
    layer5_outputs(371) <= not b;
    layer5_outputs(372) <= b;
    layer5_outputs(373) <= b;
    layer5_outputs(374) <= a and not b;
    layer5_outputs(375) <= not a;
    layer5_outputs(376) <= not a;
    layer5_outputs(377) <= a xor b;
    layer5_outputs(378) <= b and not a;
    layer5_outputs(379) <= a;
    layer5_outputs(380) <= b;
    layer5_outputs(381) <= not a;
    layer5_outputs(382) <= not (a xor b);
    layer5_outputs(383) <= a or b;
    layer5_outputs(384) <= not a;
    layer5_outputs(385) <= not b;
    layer5_outputs(386) <= not (a xor b);
    layer5_outputs(387) <= a and b;
    layer5_outputs(388) <= not a;
    layer5_outputs(389) <= a;
    layer5_outputs(390) <= not b;
    layer5_outputs(391) <= not (a and b);
    layer5_outputs(392) <= a and b;
    layer5_outputs(393) <= not (a and b);
    layer5_outputs(394) <= a;
    layer5_outputs(395) <= b;
    layer5_outputs(396) <= not b or a;
    layer5_outputs(397) <= a and b;
    layer5_outputs(398) <= b and not a;
    layer5_outputs(399) <= b;
    layer5_outputs(400) <= a or b;
    layer5_outputs(401) <= a and b;
    layer5_outputs(402) <= not a or b;
    layer5_outputs(403) <= '1';
    layer5_outputs(404) <= not a;
    layer5_outputs(405) <= not a or b;
    layer5_outputs(406) <= a;
    layer5_outputs(407) <= b;
    layer5_outputs(408) <= b;
    layer5_outputs(409) <= a;
    layer5_outputs(410) <= not a;
    layer5_outputs(411) <= b and not a;
    layer5_outputs(412) <= a and b;
    layer5_outputs(413) <= a and not b;
    layer5_outputs(414) <= a;
    layer5_outputs(415) <= b;
    layer5_outputs(416) <= not a or b;
    layer5_outputs(417) <= a;
    layer5_outputs(418) <= not a;
    layer5_outputs(419) <= a xor b;
    layer5_outputs(420) <= not b;
    layer5_outputs(421) <= not (a xor b);
    layer5_outputs(422) <= not a;
    layer5_outputs(423) <= a;
    layer5_outputs(424) <= a;
    layer5_outputs(425) <= not (a xor b);
    layer5_outputs(426) <= a or b;
    layer5_outputs(427) <= not (a xor b);
    layer5_outputs(428) <= a xor b;
    layer5_outputs(429) <= not (a xor b);
    layer5_outputs(430) <= a or b;
    layer5_outputs(431) <= a xor b;
    layer5_outputs(432) <= not (a xor b);
    layer5_outputs(433) <= a xor b;
    layer5_outputs(434) <= a and not b;
    layer5_outputs(435) <= not (a and b);
    layer5_outputs(436) <= b;
    layer5_outputs(437) <= not (a or b);
    layer5_outputs(438) <= not b;
    layer5_outputs(439) <= not a;
    layer5_outputs(440) <= not a;
    layer5_outputs(441) <= not (a xor b);
    layer5_outputs(442) <= not a;
    layer5_outputs(443) <= not a;
    layer5_outputs(444) <= b;
    layer5_outputs(445) <= b;
    layer5_outputs(446) <= not b;
    layer5_outputs(447) <= not (a and b);
    layer5_outputs(448) <= not (a xor b);
    layer5_outputs(449) <= b;
    layer5_outputs(450) <= a xor b;
    layer5_outputs(451) <= not a or b;
    layer5_outputs(452) <= not (a xor b);
    layer5_outputs(453) <= a;
    layer5_outputs(454) <= not a or b;
    layer5_outputs(455) <= b and not a;
    layer5_outputs(456) <= b;
    layer5_outputs(457) <= not (a xor b);
    layer5_outputs(458) <= not (a xor b);
    layer5_outputs(459) <= not (a xor b);
    layer5_outputs(460) <= a or b;
    layer5_outputs(461) <= not b;
    layer5_outputs(462) <= a and not b;
    layer5_outputs(463) <= not b;
    layer5_outputs(464) <= a xor b;
    layer5_outputs(465) <= not (a or b);
    layer5_outputs(466) <= b;
    layer5_outputs(467) <= not b;
    layer5_outputs(468) <= a xor b;
    layer5_outputs(469) <= b;
    layer5_outputs(470) <= not b or a;
    layer5_outputs(471) <= a;
    layer5_outputs(472) <= not (a and b);
    layer5_outputs(473) <= not (a xor b);
    layer5_outputs(474) <= not b or a;
    layer5_outputs(475) <= not (a xor b);
    layer5_outputs(476) <= not b;
    layer5_outputs(477) <= a and b;
    layer5_outputs(478) <= a xor b;
    layer5_outputs(479) <= a xor b;
    layer5_outputs(480) <= b;
    layer5_outputs(481) <= a and not b;
    layer5_outputs(482) <= not (a xor b);
    layer5_outputs(483) <= not (a or b);
    layer5_outputs(484) <= a xor b;
    layer5_outputs(485) <= not b;
    layer5_outputs(486) <= a and b;
    layer5_outputs(487) <= not b;
    layer5_outputs(488) <= a;
    layer5_outputs(489) <= '0';
    layer5_outputs(490) <= a and not b;
    layer5_outputs(491) <= not a;
    layer5_outputs(492) <= b and not a;
    layer5_outputs(493) <= not (a xor b);
    layer5_outputs(494) <= not a;
    layer5_outputs(495) <= a or b;
    layer5_outputs(496) <= not (a xor b);
    layer5_outputs(497) <= not (a and b);
    layer5_outputs(498) <= '0';
    layer5_outputs(499) <= a xor b;
    layer5_outputs(500) <= not a or b;
    layer5_outputs(501) <= a;
    layer5_outputs(502) <= a xor b;
    layer5_outputs(503) <= b;
    layer5_outputs(504) <= a;
    layer5_outputs(505) <= a and not b;
    layer5_outputs(506) <= not (a or b);
    layer5_outputs(507) <= not (a xor b);
    layer5_outputs(508) <= not a;
    layer5_outputs(509) <= not a;
    layer5_outputs(510) <= b;
    layer5_outputs(511) <= b and not a;
    layer5_outputs(512) <= a and not b;
    layer5_outputs(513) <= not b;
    layer5_outputs(514) <= b;
    layer5_outputs(515) <= b;
    layer5_outputs(516) <= a;
    layer5_outputs(517) <= a;
    layer5_outputs(518) <= not a;
    layer5_outputs(519) <= not b;
    layer5_outputs(520) <= '1';
    layer5_outputs(521) <= not (a or b);
    layer5_outputs(522) <= not a;
    layer5_outputs(523) <= b;
    layer5_outputs(524) <= a;
    layer5_outputs(525) <= a and b;
    layer5_outputs(526) <= a;
    layer5_outputs(527) <= not a;
    layer5_outputs(528) <= not (a xor b);
    layer5_outputs(529) <= not (a or b);
    layer5_outputs(530) <= not (a xor b);
    layer5_outputs(531) <= not (a xor b);
    layer5_outputs(532) <= not b or a;
    layer5_outputs(533) <= a;
    layer5_outputs(534) <= not (a and b);
    layer5_outputs(535) <= b;
    layer5_outputs(536) <= b;
    layer5_outputs(537) <= a and b;
    layer5_outputs(538) <= a or b;
    layer5_outputs(539) <= not (a xor b);
    layer5_outputs(540) <= not (a xor b);
    layer5_outputs(541) <= a;
    layer5_outputs(542) <= not a;
    layer5_outputs(543) <= not (a xor b);
    layer5_outputs(544) <= not a;
    layer5_outputs(545) <= b;
    layer5_outputs(546) <= a and b;
    layer5_outputs(547) <= not a;
    layer5_outputs(548) <= not b;
    layer5_outputs(549) <= a;
    layer5_outputs(550) <= b;
    layer5_outputs(551) <= not b;
    layer5_outputs(552) <= not b;
    layer5_outputs(553) <= a;
    layer5_outputs(554) <= not (a xor b);
    layer5_outputs(555) <= not b or a;
    layer5_outputs(556) <= not b;
    layer5_outputs(557) <= not b;
    layer5_outputs(558) <= b and not a;
    layer5_outputs(559) <= not a;
    layer5_outputs(560) <= a and b;
    layer5_outputs(561) <= not (a and b);
    layer5_outputs(562) <= a;
    layer5_outputs(563) <= not a;
    layer5_outputs(564) <= a and not b;
    layer5_outputs(565) <= a xor b;
    layer5_outputs(566) <= a or b;
    layer5_outputs(567) <= a;
    layer5_outputs(568) <= a xor b;
    layer5_outputs(569) <= not a;
    layer5_outputs(570) <= a;
    layer5_outputs(571) <= not b or a;
    layer5_outputs(572) <= not a;
    layer5_outputs(573) <= not b or a;
    layer5_outputs(574) <= not (a xor b);
    layer5_outputs(575) <= a xor b;
    layer5_outputs(576) <= b and not a;
    layer5_outputs(577) <= not a;
    layer5_outputs(578) <= not a;
    layer5_outputs(579) <= a and b;
    layer5_outputs(580) <= not a;
    layer5_outputs(581) <= not (a xor b);
    layer5_outputs(582) <= a;
    layer5_outputs(583) <= not b;
    layer5_outputs(584) <= not b;
    layer5_outputs(585) <= not (a or b);
    layer5_outputs(586) <= b;
    layer5_outputs(587) <= a;
    layer5_outputs(588) <= a or b;
    layer5_outputs(589) <= not a;
    layer5_outputs(590) <= a and b;
    layer5_outputs(591) <= not a;
    layer5_outputs(592) <= not a;
    layer5_outputs(593) <= a xor b;
    layer5_outputs(594) <= not a;
    layer5_outputs(595) <= not b;
    layer5_outputs(596) <= not (a xor b);
    layer5_outputs(597) <= not a;
    layer5_outputs(598) <= a;
    layer5_outputs(599) <= a or b;
    layer5_outputs(600) <= not a;
    layer5_outputs(601) <= a;
    layer5_outputs(602) <= not b;
    layer5_outputs(603) <= not b;
    layer5_outputs(604) <= not a;
    layer5_outputs(605) <= b;
    layer5_outputs(606) <= not b;
    layer5_outputs(607) <= a;
    layer5_outputs(608) <= not a;
    layer5_outputs(609) <= not b;
    layer5_outputs(610) <= '0';
    layer5_outputs(611) <= not (a or b);
    layer5_outputs(612) <= b and not a;
    layer5_outputs(613) <= a;
    layer5_outputs(614) <= a and not b;
    layer5_outputs(615) <= not (a or b);
    layer5_outputs(616) <= not b;
    layer5_outputs(617) <= a and b;
    layer5_outputs(618) <= a;
    layer5_outputs(619) <= a or b;
    layer5_outputs(620) <= not b;
    layer5_outputs(621) <= not b or a;
    layer5_outputs(622) <= a and not b;
    layer5_outputs(623) <= not (a and b);
    layer5_outputs(624) <= not (a or b);
    layer5_outputs(625) <= a and b;
    layer5_outputs(626) <= a;
    layer5_outputs(627) <= not a;
    layer5_outputs(628) <= not a or b;
    layer5_outputs(629) <= a;
    layer5_outputs(630) <= b;
    layer5_outputs(631) <= not (a and b);
    layer5_outputs(632) <= a and not b;
    layer5_outputs(633) <= b;
    layer5_outputs(634) <= a;
    layer5_outputs(635) <= not a or b;
    layer5_outputs(636) <= a xor b;
    layer5_outputs(637) <= b and not a;
    layer5_outputs(638) <= not (a and b);
    layer5_outputs(639) <= not (a xor b);
    layer5_outputs(640) <= a xor b;
    layer5_outputs(641) <= a and not b;
    layer5_outputs(642) <= not a or b;
    layer5_outputs(643) <= not a;
    layer5_outputs(644) <= not (a and b);
    layer5_outputs(645) <= not (a or b);
    layer5_outputs(646) <= not a;
    layer5_outputs(647) <= not b;
    layer5_outputs(648) <= a;
    layer5_outputs(649) <= not b or a;
    layer5_outputs(650) <= not a or b;
    layer5_outputs(651) <= not (a xor b);
    layer5_outputs(652) <= a and b;
    layer5_outputs(653) <= not b;
    layer5_outputs(654) <= a or b;
    layer5_outputs(655) <= a;
    layer5_outputs(656) <= a;
    layer5_outputs(657) <= b;
    layer5_outputs(658) <= a and b;
    layer5_outputs(659) <= not b or a;
    layer5_outputs(660) <= not (a or b);
    layer5_outputs(661) <= not b;
    layer5_outputs(662) <= not (a or b);
    layer5_outputs(663) <= b;
    layer5_outputs(664) <= a and b;
    layer5_outputs(665) <= a xor b;
    layer5_outputs(666) <= b;
    layer5_outputs(667) <= a;
    layer5_outputs(668) <= a xor b;
    layer5_outputs(669) <= a or b;
    layer5_outputs(670) <= b;
    layer5_outputs(671) <= not b;
    layer5_outputs(672) <= a;
    layer5_outputs(673) <= not (a xor b);
    layer5_outputs(674) <= not a;
    layer5_outputs(675) <= a or b;
    layer5_outputs(676) <= not a or b;
    layer5_outputs(677) <= not b;
    layer5_outputs(678) <= not b or a;
    layer5_outputs(679) <= b;
    layer5_outputs(680) <= a and b;
    layer5_outputs(681) <= not b;
    layer5_outputs(682) <= a and not b;
    layer5_outputs(683) <= a;
    layer5_outputs(684) <= a;
    layer5_outputs(685) <= a or b;
    layer5_outputs(686) <= b;
    layer5_outputs(687) <= not a or b;
    layer5_outputs(688) <= a;
    layer5_outputs(689) <= a and not b;
    layer5_outputs(690) <= a;
    layer5_outputs(691) <= not a;
    layer5_outputs(692) <= a;
    layer5_outputs(693) <= not b;
    layer5_outputs(694) <= a and b;
    layer5_outputs(695) <= not b;
    layer5_outputs(696) <= not (a or b);
    layer5_outputs(697) <= b;
    layer5_outputs(698) <= not a;
    layer5_outputs(699) <= b;
    layer5_outputs(700) <= a;
    layer5_outputs(701) <= a xor b;
    layer5_outputs(702) <= a xor b;
    layer5_outputs(703) <= not b;
    layer5_outputs(704) <= a and not b;
    layer5_outputs(705) <= a and not b;
    layer5_outputs(706) <= not (a xor b);
    layer5_outputs(707) <= not b;
    layer5_outputs(708) <= not b;
    layer5_outputs(709) <= not (a xor b);
    layer5_outputs(710) <= b and not a;
    layer5_outputs(711) <= not b or a;
    layer5_outputs(712) <= not a;
    layer5_outputs(713) <= b and not a;
    layer5_outputs(714) <= b;
    layer5_outputs(715) <= a;
    layer5_outputs(716) <= not b;
    layer5_outputs(717) <= a and b;
    layer5_outputs(718) <= a and not b;
    layer5_outputs(719) <= b;
    layer5_outputs(720) <= not b or a;
    layer5_outputs(721) <= not a or b;
    layer5_outputs(722) <= b;
    layer5_outputs(723) <= not (a xor b);
    layer5_outputs(724) <= '0';
    layer5_outputs(725) <= not b;
    layer5_outputs(726) <= a;
    layer5_outputs(727) <= not a;
    layer5_outputs(728) <= not b;
    layer5_outputs(729) <= b and not a;
    layer5_outputs(730) <= not (a or b);
    layer5_outputs(731) <= not (a xor b);
    layer5_outputs(732) <= not a;
    layer5_outputs(733) <= a;
    layer5_outputs(734) <= b and not a;
    layer5_outputs(735) <= a and b;
    layer5_outputs(736) <= a and not b;
    layer5_outputs(737) <= a;
    layer5_outputs(738) <= a;
    layer5_outputs(739) <= b;
    layer5_outputs(740) <= not b;
    layer5_outputs(741) <= a and b;
    layer5_outputs(742) <= b;
    layer5_outputs(743) <= a or b;
    layer5_outputs(744) <= a and b;
    layer5_outputs(745) <= a and b;
    layer5_outputs(746) <= a;
    layer5_outputs(747) <= not b;
    layer5_outputs(748) <= not a;
    layer5_outputs(749) <= not b;
    layer5_outputs(750) <= b and not a;
    layer5_outputs(751) <= not (a xor b);
    layer5_outputs(752) <= not a;
    layer5_outputs(753) <= not a or b;
    layer5_outputs(754) <= a;
    layer5_outputs(755) <= not a;
    layer5_outputs(756) <= a;
    layer5_outputs(757) <= not a;
    layer5_outputs(758) <= not a;
    layer5_outputs(759) <= not b or a;
    layer5_outputs(760) <= not (a and b);
    layer5_outputs(761) <= not (a or b);
    layer5_outputs(762) <= a;
    layer5_outputs(763) <= a;
    layer5_outputs(764) <= not a;
    layer5_outputs(765) <= not (a xor b);
    layer5_outputs(766) <= not (a xor b);
    layer5_outputs(767) <= '1';
    layer5_outputs(768) <= not (a and b);
    layer5_outputs(769) <= not b;
    layer5_outputs(770) <= not (a or b);
    layer5_outputs(771) <= not (a xor b);
    layer5_outputs(772) <= not b;
    layer5_outputs(773) <= a;
    layer5_outputs(774) <= not b or a;
    layer5_outputs(775) <= not b or a;
    layer5_outputs(776) <= a xor b;
    layer5_outputs(777) <= a xor b;
    layer5_outputs(778) <= b and not a;
    layer5_outputs(779) <= a and b;
    layer5_outputs(780) <= not a;
    layer5_outputs(781) <= a and not b;
    layer5_outputs(782) <= a;
    layer5_outputs(783) <= not a or b;
    layer5_outputs(784) <= not a;
    layer5_outputs(785) <= not a;
    layer5_outputs(786) <= b;
    layer5_outputs(787) <= b and not a;
    layer5_outputs(788) <= a xor b;
    layer5_outputs(789) <= not (a and b);
    layer5_outputs(790) <= not b;
    layer5_outputs(791) <= not b or a;
    layer5_outputs(792) <= not (a or b);
    layer5_outputs(793) <= not (a xor b);
    layer5_outputs(794) <= not b;
    layer5_outputs(795) <= not (a and b);
    layer5_outputs(796) <= b and not a;
    layer5_outputs(797) <= a or b;
    layer5_outputs(798) <= not a;
    layer5_outputs(799) <= not b;
    layer5_outputs(800) <= not (a xor b);
    layer5_outputs(801) <= a xor b;
    layer5_outputs(802) <= not (a or b);
    layer5_outputs(803) <= not a;
    layer5_outputs(804) <= not a;
    layer5_outputs(805) <= not a or b;
    layer5_outputs(806) <= a and b;
    layer5_outputs(807) <= a;
    layer5_outputs(808) <= not (a or b);
    layer5_outputs(809) <= a;
    layer5_outputs(810) <= not b;
    layer5_outputs(811) <= a and b;
    layer5_outputs(812) <= not (a or b);
    layer5_outputs(813) <= a;
    layer5_outputs(814) <= b;
    layer5_outputs(815) <= not a;
    layer5_outputs(816) <= a and not b;
    layer5_outputs(817) <= a or b;
    layer5_outputs(818) <= a and not b;
    layer5_outputs(819) <= b;
    layer5_outputs(820) <= b and not a;
    layer5_outputs(821) <= a or b;
    layer5_outputs(822) <= not b;
    layer5_outputs(823) <= a and b;
    layer5_outputs(824) <= not b;
    layer5_outputs(825) <= a and b;
    layer5_outputs(826) <= not (a and b);
    layer5_outputs(827) <= not a or b;
    layer5_outputs(828) <= not b;
    layer5_outputs(829) <= not a or b;
    layer5_outputs(830) <= not b;
    layer5_outputs(831) <= a xor b;
    layer5_outputs(832) <= a;
    layer5_outputs(833) <= a or b;
    layer5_outputs(834) <= a;
    layer5_outputs(835) <= not (a xor b);
    layer5_outputs(836) <= not b;
    layer5_outputs(837) <= not a;
    layer5_outputs(838) <= b;
    layer5_outputs(839) <= not b;
    layer5_outputs(840) <= not (a or b);
    layer5_outputs(841) <= a xor b;
    layer5_outputs(842) <= not a;
    layer5_outputs(843) <= not a;
    layer5_outputs(844) <= a xor b;
    layer5_outputs(845) <= not a;
    layer5_outputs(846) <= a;
    layer5_outputs(847) <= not (a xor b);
    layer5_outputs(848) <= not a;
    layer5_outputs(849) <= a and not b;
    layer5_outputs(850) <= not a;
    layer5_outputs(851) <= a or b;
    layer5_outputs(852) <= not a or b;
    layer5_outputs(853) <= not b or a;
    layer5_outputs(854) <= '1';
    layer5_outputs(855) <= a or b;
    layer5_outputs(856) <= a xor b;
    layer5_outputs(857) <= a and not b;
    layer5_outputs(858) <= a and b;
    layer5_outputs(859) <= not a;
    layer5_outputs(860) <= not (a and b);
    layer5_outputs(861) <= b;
    layer5_outputs(862) <= not a;
    layer5_outputs(863) <= not b or a;
    layer5_outputs(864) <= not a;
    layer5_outputs(865) <= b;
    layer5_outputs(866) <= not a;
    layer5_outputs(867) <= not a;
    layer5_outputs(868) <= a;
    layer5_outputs(869) <= not b;
    layer5_outputs(870) <= not a or b;
    layer5_outputs(871) <= a;
    layer5_outputs(872) <= not b or a;
    layer5_outputs(873) <= a or b;
    layer5_outputs(874) <= not b;
    layer5_outputs(875) <= a xor b;
    layer5_outputs(876) <= not b;
    layer5_outputs(877) <= not a;
    layer5_outputs(878) <= b;
    layer5_outputs(879) <= a and b;
    layer5_outputs(880) <= a xor b;
    layer5_outputs(881) <= b;
    layer5_outputs(882) <= a xor b;
    layer5_outputs(883) <= not (a and b);
    layer5_outputs(884) <= b and not a;
    layer5_outputs(885) <= a and b;
    layer5_outputs(886) <= a;
    layer5_outputs(887) <= not a;
    layer5_outputs(888) <= not (a or b);
    layer5_outputs(889) <= not b or a;
    layer5_outputs(890) <= a or b;
    layer5_outputs(891) <= a or b;
    layer5_outputs(892) <= a or b;
    layer5_outputs(893) <= '0';
    layer5_outputs(894) <= not b;
    layer5_outputs(895) <= not (a xor b);
    layer5_outputs(896) <= a;
    layer5_outputs(897) <= b and not a;
    layer5_outputs(898) <= a;
    layer5_outputs(899) <= not (a and b);
    layer5_outputs(900) <= not b;
    layer5_outputs(901) <= a and not b;
    layer5_outputs(902) <= not (a and b);
    layer5_outputs(903) <= not (a or b);
    layer5_outputs(904) <= not a or b;
    layer5_outputs(905) <= not (a xor b);
    layer5_outputs(906) <= a and not b;
    layer5_outputs(907) <= a xor b;
    layer5_outputs(908) <= a and b;
    layer5_outputs(909) <= a or b;
    layer5_outputs(910) <= not a or b;
    layer5_outputs(911) <= not b or a;
    layer5_outputs(912) <= a xor b;
    layer5_outputs(913) <= not a or b;
    layer5_outputs(914) <= a xor b;
    layer5_outputs(915) <= a and not b;
    layer5_outputs(916) <= a;
    layer5_outputs(917) <= a and b;
    layer5_outputs(918) <= a or b;
    layer5_outputs(919) <= a and not b;
    layer5_outputs(920) <= b;
    layer5_outputs(921) <= not a;
    layer5_outputs(922) <= not a;
    layer5_outputs(923) <= b;
    layer5_outputs(924) <= not a;
    layer5_outputs(925) <= not b;
    layer5_outputs(926) <= a and b;
    layer5_outputs(927) <= a or b;
    layer5_outputs(928) <= not (a xor b);
    layer5_outputs(929) <= b;
    layer5_outputs(930) <= b;
    layer5_outputs(931) <= a or b;
    layer5_outputs(932) <= not b;
    layer5_outputs(933) <= b;
    layer5_outputs(934) <= '1';
    layer5_outputs(935) <= a xor b;
    layer5_outputs(936) <= a;
    layer5_outputs(937) <= b;
    layer5_outputs(938) <= a;
    layer5_outputs(939) <= not a;
    layer5_outputs(940) <= not b;
    layer5_outputs(941) <= a or b;
    layer5_outputs(942) <= a;
    layer5_outputs(943) <= not a or b;
    layer5_outputs(944) <= b and not a;
    layer5_outputs(945) <= not (a or b);
    layer5_outputs(946) <= not (a and b);
    layer5_outputs(947) <= not b;
    layer5_outputs(948) <= b and not a;
    layer5_outputs(949) <= not (a and b);
    layer5_outputs(950) <= not b;
    layer5_outputs(951) <= b and not a;
    layer5_outputs(952) <= not (a and b);
    layer5_outputs(953) <= not (a and b);
    layer5_outputs(954) <= not b or a;
    layer5_outputs(955) <= not b or a;
    layer5_outputs(956) <= not a;
    layer5_outputs(957) <= a;
    layer5_outputs(958) <= b;
    layer5_outputs(959) <= a and not b;
    layer5_outputs(960) <= a and b;
    layer5_outputs(961) <= not a;
    layer5_outputs(962) <= not b;
    layer5_outputs(963) <= a and not b;
    layer5_outputs(964) <= a;
    layer5_outputs(965) <= a;
    layer5_outputs(966) <= a xor b;
    layer5_outputs(967) <= a;
    layer5_outputs(968) <= a;
    layer5_outputs(969) <= not b;
    layer5_outputs(970) <= not a;
    layer5_outputs(971) <= a and not b;
    layer5_outputs(972) <= a and not b;
    layer5_outputs(973) <= a and not b;
    layer5_outputs(974) <= not (a xor b);
    layer5_outputs(975) <= not b;
    layer5_outputs(976) <= not b;
    layer5_outputs(977) <= not (a xor b);
    layer5_outputs(978) <= a xor b;
    layer5_outputs(979) <= a;
    layer5_outputs(980) <= '0';
    layer5_outputs(981) <= a and b;
    layer5_outputs(982) <= not (a xor b);
    layer5_outputs(983) <= b;
    layer5_outputs(984) <= a and b;
    layer5_outputs(985) <= not (a or b);
    layer5_outputs(986) <= a and not b;
    layer5_outputs(987) <= not a;
    layer5_outputs(988) <= a and not b;
    layer5_outputs(989) <= b;
    layer5_outputs(990) <= not a;
    layer5_outputs(991) <= not b or a;
    layer5_outputs(992) <= a xor b;
    layer5_outputs(993) <= a and b;
    layer5_outputs(994) <= not a;
    layer5_outputs(995) <= b;
    layer5_outputs(996) <= a and not b;
    layer5_outputs(997) <= not (a xor b);
    layer5_outputs(998) <= a and b;
    layer5_outputs(999) <= not a or b;
    layer5_outputs(1000) <= not (a and b);
    layer5_outputs(1001) <= not a or b;
    layer5_outputs(1002) <= not b;
    layer5_outputs(1003) <= not (a and b);
    layer5_outputs(1004) <= a xor b;
    layer5_outputs(1005) <= a or b;
    layer5_outputs(1006) <= a and b;
    layer5_outputs(1007) <= a and not b;
    layer5_outputs(1008) <= not (a or b);
    layer5_outputs(1009) <= not a;
    layer5_outputs(1010) <= not b or a;
    layer5_outputs(1011) <= a xor b;
    layer5_outputs(1012) <= not (a and b);
    layer5_outputs(1013) <= not b;
    layer5_outputs(1014) <= b;
    layer5_outputs(1015) <= b and not a;
    layer5_outputs(1016) <= a and not b;
    layer5_outputs(1017) <= not (a xor b);
    layer5_outputs(1018) <= a xor b;
    layer5_outputs(1019) <= not a;
    layer5_outputs(1020) <= a and not b;
    layer5_outputs(1021) <= not b;
    layer5_outputs(1022) <= a;
    layer5_outputs(1023) <= a xor b;
    layer5_outputs(1024) <= not a;
    layer5_outputs(1025) <= a;
    layer5_outputs(1026) <= a or b;
    layer5_outputs(1027) <= not a;
    layer5_outputs(1028) <= not b;
    layer5_outputs(1029) <= not a or b;
    layer5_outputs(1030) <= not (a and b);
    layer5_outputs(1031) <= b;
    layer5_outputs(1032) <= b and not a;
    layer5_outputs(1033) <= not a;
    layer5_outputs(1034) <= a;
    layer5_outputs(1035) <= a;
    layer5_outputs(1036) <= b and not a;
    layer5_outputs(1037) <= not b;
    layer5_outputs(1038) <= b;
    layer5_outputs(1039) <= not a;
    layer5_outputs(1040) <= b;
    layer5_outputs(1041) <= a or b;
    layer5_outputs(1042) <= b;
    layer5_outputs(1043) <= a or b;
    layer5_outputs(1044) <= a xor b;
    layer5_outputs(1045) <= not a;
    layer5_outputs(1046) <= not (a or b);
    layer5_outputs(1047) <= not b;
    layer5_outputs(1048) <= a;
    layer5_outputs(1049) <= not (a and b);
    layer5_outputs(1050) <= not (a xor b);
    layer5_outputs(1051) <= a;
    layer5_outputs(1052) <= not (a or b);
    layer5_outputs(1053) <= a and not b;
    layer5_outputs(1054) <= not b or a;
    layer5_outputs(1055) <= a;
    layer5_outputs(1056) <= a;
    layer5_outputs(1057) <= '0';
    layer5_outputs(1058) <= not b or a;
    layer5_outputs(1059) <= b;
    layer5_outputs(1060) <= b and not a;
    layer5_outputs(1061) <= a;
    layer5_outputs(1062) <= a or b;
    layer5_outputs(1063) <= not b or a;
    layer5_outputs(1064) <= a and b;
    layer5_outputs(1065) <= b and not a;
    layer5_outputs(1066) <= '1';
    layer5_outputs(1067) <= b;
    layer5_outputs(1068) <= not b or a;
    layer5_outputs(1069) <= not (a or b);
    layer5_outputs(1070) <= not a or b;
    layer5_outputs(1071) <= b;
    layer5_outputs(1072) <= not a;
    layer5_outputs(1073) <= not a;
    layer5_outputs(1074) <= b and not a;
    layer5_outputs(1075) <= a and b;
    layer5_outputs(1076) <= not b;
    layer5_outputs(1077) <= b;
    layer5_outputs(1078) <= not b;
    layer5_outputs(1079) <= not (a xor b);
    layer5_outputs(1080) <= not b;
    layer5_outputs(1081) <= not (a xor b);
    layer5_outputs(1082) <= not a;
    layer5_outputs(1083) <= not (a or b);
    layer5_outputs(1084) <= not b;
    layer5_outputs(1085) <= a;
    layer5_outputs(1086) <= not a;
    layer5_outputs(1087) <= not b;
    layer5_outputs(1088) <= a and b;
    layer5_outputs(1089) <= a;
    layer5_outputs(1090) <= not a;
    layer5_outputs(1091) <= not a;
    layer5_outputs(1092) <= not b;
    layer5_outputs(1093) <= not b;
    layer5_outputs(1094) <= a;
    layer5_outputs(1095) <= not (a and b);
    layer5_outputs(1096) <= not b or a;
    layer5_outputs(1097) <= a or b;
    layer5_outputs(1098) <= not (a or b);
    layer5_outputs(1099) <= a;
    layer5_outputs(1100) <= not a;
    layer5_outputs(1101) <= a and not b;
    layer5_outputs(1102) <= b;
    layer5_outputs(1103) <= b;
    layer5_outputs(1104) <= not b or a;
    layer5_outputs(1105) <= not (a and b);
    layer5_outputs(1106) <= not b;
    layer5_outputs(1107) <= b;
    layer5_outputs(1108) <= not a;
    layer5_outputs(1109) <= a;
    layer5_outputs(1110) <= not (a or b);
    layer5_outputs(1111) <= not a;
    layer5_outputs(1112) <= not a;
    layer5_outputs(1113) <= a;
    layer5_outputs(1114) <= a and not b;
    layer5_outputs(1115) <= not (a or b);
    layer5_outputs(1116) <= a;
    layer5_outputs(1117) <= not (a xor b);
    layer5_outputs(1118) <= not b;
    layer5_outputs(1119) <= not a;
    layer5_outputs(1120) <= a;
    layer5_outputs(1121) <= a;
    layer5_outputs(1122) <= a xor b;
    layer5_outputs(1123) <= not b or a;
    layer5_outputs(1124) <= a;
    layer5_outputs(1125) <= a or b;
    layer5_outputs(1126) <= not b;
    layer5_outputs(1127) <= not b;
    layer5_outputs(1128) <= b;
    layer5_outputs(1129) <= a;
    layer5_outputs(1130) <= a and not b;
    layer5_outputs(1131) <= b and not a;
    layer5_outputs(1132) <= not a;
    layer5_outputs(1133) <= not b;
    layer5_outputs(1134) <= b;
    layer5_outputs(1135) <= a and not b;
    layer5_outputs(1136) <= a;
    layer5_outputs(1137) <= not b or a;
    layer5_outputs(1138) <= not b;
    layer5_outputs(1139) <= a and b;
    layer5_outputs(1140) <= not a;
    layer5_outputs(1141) <= not b or a;
    layer5_outputs(1142) <= not (a or b);
    layer5_outputs(1143) <= b;
    layer5_outputs(1144) <= not (a and b);
    layer5_outputs(1145) <= not a or b;
    layer5_outputs(1146) <= not a or b;
    layer5_outputs(1147) <= a or b;
    layer5_outputs(1148) <= not b;
    layer5_outputs(1149) <= b;
    layer5_outputs(1150) <= not (a or b);
    layer5_outputs(1151) <= not b or a;
    layer5_outputs(1152) <= not a;
    layer5_outputs(1153) <= a or b;
    layer5_outputs(1154) <= not a;
    layer5_outputs(1155) <= b and not a;
    layer5_outputs(1156) <= not (a and b);
    layer5_outputs(1157) <= b and not a;
    layer5_outputs(1158) <= a xor b;
    layer5_outputs(1159) <= a xor b;
    layer5_outputs(1160) <= a xor b;
    layer5_outputs(1161) <= not b;
    layer5_outputs(1162) <= a;
    layer5_outputs(1163) <= a and not b;
    layer5_outputs(1164) <= b;
    layer5_outputs(1165) <= '0';
    layer5_outputs(1166) <= not b;
    layer5_outputs(1167) <= not a or b;
    layer5_outputs(1168) <= not b;
    layer5_outputs(1169) <= not (a or b);
    layer5_outputs(1170) <= a xor b;
    layer5_outputs(1171) <= not (a xor b);
    layer5_outputs(1172) <= not b or a;
    layer5_outputs(1173) <= b and not a;
    layer5_outputs(1174) <= not (a and b);
    layer5_outputs(1175) <= not a;
    layer5_outputs(1176) <= not b or a;
    layer5_outputs(1177) <= not b or a;
    layer5_outputs(1178) <= not (a xor b);
    layer5_outputs(1179) <= a or b;
    layer5_outputs(1180) <= not b;
    layer5_outputs(1181) <= not (a or b);
    layer5_outputs(1182) <= a;
    layer5_outputs(1183) <= a xor b;
    layer5_outputs(1184) <= a xor b;
    layer5_outputs(1185) <= a and not b;
    layer5_outputs(1186) <= b and not a;
    layer5_outputs(1187) <= not b;
    layer5_outputs(1188) <= b;
    layer5_outputs(1189) <= a and b;
    layer5_outputs(1190) <= not (a xor b);
    layer5_outputs(1191) <= not b;
    layer5_outputs(1192) <= a xor b;
    layer5_outputs(1193) <= not (a xor b);
    layer5_outputs(1194) <= a;
    layer5_outputs(1195) <= b;
    layer5_outputs(1196) <= not (a and b);
    layer5_outputs(1197) <= not b;
    layer5_outputs(1198) <= not (a and b);
    layer5_outputs(1199) <= not (a xor b);
    layer5_outputs(1200) <= not b;
    layer5_outputs(1201) <= a;
    layer5_outputs(1202) <= not b or a;
    layer5_outputs(1203) <= a;
    layer5_outputs(1204) <= not a or b;
    layer5_outputs(1205) <= not (a and b);
    layer5_outputs(1206) <= not b or a;
    layer5_outputs(1207) <= not b;
    layer5_outputs(1208) <= a;
    layer5_outputs(1209) <= not b;
    layer5_outputs(1210) <= b;
    layer5_outputs(1211) <= a;
    layer5_outputs(1212) <= a and b;
    layer5_outputs(1213) <= a;
    layer5_outputs(1214) <= not b or a;
    layer5_outputs(1215) <= not a;
    layer5_outputs(1216) <= not a;
    layer5_outputs(1217) <= not b or a;
    layer5_outputs(1218) <= not (a and b);
    layer5_outputs(1219) <= not a;
    layer5_outputs(1220) <= not b or a;
    layer5_outputs(1221) <= b and not a;
    layer5_outputs(1222) <= not (a and b);
    layer5_outputs(1223) <= a or b;
    layer5_outputs(1224) <= not b;
    layer5_outputs(1225) <= not (a or b);
    layer5_outputs(1226) <= not a or b;
    layer5_outputs(1227) <= not (a or b);
    layer5_outputs(1228) <= not (a or b);
    layer5_outputs(1229) <= not a;
    layer5_outputs(1230) <= not (a and b);
    layer5_outputs(1231) <= not a;
    layer5_outputs(1232) <= a;
    layer5_outputs(1233) <= not a;
    layer5_outputs(1234) <= not a or b;
    layer5_outputs(1235) <= a and b;
    layer5_outputs(1236) <= a xor b;
    layer5_outputs(1237) <= b;
    layer5_outputs(1238) <= a;
    layer5_outputs(1239) <= not a or b;
    layer5_outputs(1240) <= not a;
    layer5_outputs(1241) <= not (a xor b);
    layer5_outputs(1242) <= b;
    layer5_outputs(1243) <= not (a xor b);
    layer5_outputs(1244) <= b and not a;
    layer5_outputs(1245) <= a;
    layer5_outputs(1246) <= not (a xor b);
    layer5_outputs(1247) <= not b;
    layer5_outputs(1248) <= not b;
    layer5_outputs(1249) <= b;
    layer5_outputs(1250) <= a and b;
    layer5_outputs(1251) <= b;
    layer5_outputs(1252) <= a;
    layer5_outputs(1253) <= a xor b;
    layer5_outputs(1254) <= b;
    layer5_outputs(1255) <= not (a or b);
    layer5_outputs(1256) <= a;
    layer5_outputs(1257) <= not b or a;
    layer5_outputs(1258) <= not (a xor b);
    layer5_outputs(1259) <= b and not a;
    layer5_outputs(1260) <= a;
    layer5_outputs(1261) <= a or b;
    layer5_outputs(1262) <= not a;
    layer5_outputs(1263) <= not a;
    layer5_outputs(1264) <= b;
    layer5_outputs(1265) <= not b or a;
    layer5_outputs(1266) <= a and not b;
    layer5_outputs(1267) <= a and not b;
    layer5_outputs(1268) <= a;
    layer5_outputs(1269) <= not a;
    layer5_outputs(1270) <= b;
    layer5_outputs(1271) <= a xor b;
    layer5_outputs(1272) <= not b or a;
    layer5_outputs(1273) <= not a;
    layer5_outputs(1274) <= not (a xor b);
    layer5_outputs(1275) <= b and not a;
    layer5_outputs(1276) <= a and b;
    layer5_outputs(1277) <= not b;
    layer5_outputs(1278) <= a;
    layer5_outputs(1279) <= a xor b;
    layer5_outputs(1280) <= a xor b;
    layer5_outputs(1281) <= a xor b;
    layer5_outputs(1282) <= not b;
    layer5_outputs(1283) <= a and b;
    layer5_outputs(1284) <= a;
    layer5_outputs(1285) <= a;
    layer5_outputs(1286) <= a xor b;
    layer5_outputs(1287) <= a xor b;
    layer5_outputs(1288) <= b and not a;
    layer5_outputs(1289) <= not (a or b);
    layer5_outputs(1290) <= not (a xor b);
    layer5_outputs(1291) <= not a or b;
    layer5_outputs(1292) <= a and not b;
    layer5_outputs(1293) <= not b or a;
    layer5_outputs(1294) <= b and not a;
    layer5_outputs(1295) <= not (a or b);
    layer5_outputs(1296) <= b;
    layer5_outputs(1297) <= not (a xor b);
    layer5_outputs(1298) <= not a or b;
    layer5_outputs(1299) <= b;
    layer5_outputs(1300) <= not (a or b);
    layer5_outputs(1301) <= a xor b;
    layer5_outputs(1302) <= b;
    layer5_outputs(1303) <= not a;
    layer5_outputs(1304) <= not a;
    layer5_outputs(1305) <= not (a and b);
    layer5_outputs(1306) <= b and not a;
    layer5_outputs(1307) <= not a;
    layer5_outputs(1308) <= a;
    layer5_outputs(1309) <= a;
    layer5_outputs(1310) <= not a;
    layer5_outputs(1311) <= a xor b;
    layer5_outputs(1312) <= a xor b;
    layer5_outputs(1313) <= not a;
    layer5_outputs(1314) <= a and not b;
    layer5_outputs(1315) <= b;
    layer5_outputs(1316) <= not (a and b);
    layer5_outputs(1317) <= a xor b;
    layer5_outputs(1318) <= not b;
    layer5_outputs(1319) <= not b;
    layer5_outputs(1320) <= not a or b;
    layer5_outputs(1321) <= not b;
    layer5_outputs(1322) <= not a;
    layer5_outputs(1323) <= a;
    layer5_outputs(1324) <= not (a and b);
    layer5_outputs(1325) <= not a;
    layer5_outputs(1326) <= not (a xor b);
    layer5_outputs(1327) <= not (a xor b);
    layer5_outputs(1328) <= not b;
    layer5_outputs(1329) <= not (a xor b);
    layer5_outputs(1330) <= not b;
    layer5_outputs(1331) <= a and b;
    layer5_outputs(1332) <= b and not a;
    layer5_outputs(1333) <= b;
    layer5_outputs(1334) <= not b or a;
    layer5_outputs(1335) <= a or b;
    layer5_outputs(1336) <= not (a or b);
    layer5_outputs(1337) <= not (a xor b);
    layer5_outputs(1338) <= a xor b;
    layer5_outputs(1339) <= a;
    layer5_outputs(1340) <= b;
    layer5_outputs(1341) <= a xor b;
    layer5_outputs(1342) <= not a;
    layer5_outputs(1343) <= a and not b;
    layer5_outputs(1344) <= not b or a;
    layer5_outputs(1345) <= not b;
    layer5_outputs(1346) <= not b;
    layer5_outputs(1347) <= b;
    layer5_outputs(1348) <= a or b;
    layer5_outputs(1349) <= a or b;
    layer5_outputs(1350) <= not b;
    layer5_outputs(1351) <= a;
    layer5_outputs(1352) <= a or b;
    layer5_outputs(1353) <= a;
    layer5_outputs(1354) <= not (a and b);
    layer5_outputs(1355) <= a xor b;
    layer5_outputs(1356) <= not a;
    layer5_outputs(1357) <= not a;
    layer5_outputs(1358) <= not b or a;
    layer5_outputs(1359) <= a;
    layer5_outputs(1360) <= not a;
    layer5_outputs(1361) <= not (a and b);
    layer5_outputs(1362) <= not a;
    layer5_outputs(1363) <= b;
    layer5_outputs(1364) <= not a or b;
    layer5_outputs(1365) <= not (a or b);
    layer5_outputs(1366) <= b and not a;
    layer5_outputs(1367) <= not a;
    layer5_outputs(1368) <= a;
    layer5_outputs(1369) <= a;
    layer5_outputs(1370) <= not (a xor b);
    layer5_outputs(1371) <= b;
    layer5_outputs(1372) <= a or b;
    layer5_outputs(1373) <= not a;
    layer5_outputs(1374) <= b;
    layer5_outputs(1375) <= a xor b;
    layer5_outputs(1376) <= not (a and b);
    layer5_outputs(1377) <= not (a and b);
    layer5_outputs(1378) <= not (a and b);
    layer5_outputs(1379) <= a;
    layer5_outputs(1380) <= b;
    layer5_outputs(1381) <= not b or a;
    layer5_outputs(1382) <= b;
    layer5_outputs(1383) <= not a or b;
    layer5_outputs(1384) <= not (a and b);
    layer5_outputs(1385) <= b and not a;
    layer5_outputs(1386) <= '1';
    layer5_outputs(1387) <= not a;
    layer5_outputs(1388) <= not b or a;
    layer5_outputs(1389) <= a;
    layer5_outputs(1390) <= a;
    layer5_outputs(1391) <= a;
    layer5_outputs(1392) <= a or b;
    layer5_outputs(1393) <= not (a and b);
    layer5_outputs(1394) <= not b;
    layer5_outputs(1395) <= not (a xor b);
    layer5_outputs(1396) <= b;
    layer5_outputs(1397) <= not b;
    layer5_outputs(1398) <= a xor b;
    layer5_outputs(1399) <= a and not b;
    layer5_outputs(1400) <= not a;
    layer5_outputs(1401) <= not (a xor b);
    layer5_outputs(1402) <= not a;
    layer5_outputs(1403) <= not a;
    layer5_outputs(1404) <= not a;
    layer5_outputs(1405) <= a and b;
    layer5_outputs(1406) <= b and not a;
    layer5_outputs(1407) <= a and not b;
    layer5_outputs(1408) <= not a;
    layer5_outputs(1409) <= not b or a;
    layer5_outputs(1410) <= a and b;
    layer5_outputs(1411) <= not b or a;
    layer5_outputs(1412) <= a and b;
    layer5_outputs(1413) <= a and not b;
    layer5_outputs(1414) <= a;
    layer5_outputs(1415) <= a and not b;
    layer5_outputs(1416) <= not a;
    layer5_outputs(1417) <= not (a and b);
    layer5_outputs(1418) <= a;
    layer5_outputs(1419) <= not (a xor b);
    layer5_outputs(1420) <= not (a xor b);
    layer5_outputs(1421) <= a xor b;
    layer5_outputs(1422) <= not (a xor b);
    layer5_outputs(1423) <= not a;
    layer5_outputs(1424) <= a or b;
    layer5_outputs(1425) <= b;
    layer5_outputs(1426) <= not b or a;
    layer5_outputs(1427) <= not b or a;
    layer5_outputs(1428) <= not b;
    layer5_outputs(1429) <= not b;
    layer5_outputs(1430) <= '0';
    layer5_outputs(1431) <= not a or b;
    layer5_outputs(1432) <= a xor b;
    layer5_outputs(1433) <= not a;
    layer5_outputs(1434) <= not (a xor b);
    layer5_outputs(1435) <= not a;
    layer5_outputs(1436) <= not a;
    layer5_outputs(1437) <= a;
    layer5_outputs(1438) <= not a or b;
    layer5_outputs(1439) <= not a;
    layer5_outputs(1440) <= not a;
    layer5_outputs(1441) <= a or b;
    layer5_outputs(1442) <= b;
    layer5_outputs(1443) <= not b;
    layer5_outputs(1444) <= not a;
    layer5_outputs(1445) <= not a;
    layer5_outputs(1446) <= '1';
    layer5_outputs(1447) <= a xor b;
    layer5_outputs(1448) <= not b;
    layer5_outputs(1449) <= not (a xor b);
    layer5_outputs(1450) <= not a;
    layer5_outputs(1451) <= a;
    layer5_outputs(1452) <= b;
    layer5_outputs(1453) <= a;
    layer5_outputs(1454) <= a and b;
    layer5_outputs(1455) <= a;
    layer5_outputs(1456) <= not (a xor b);
    layer5_outputs(1457) <= b;
    layer5_outputs(1458) <= not a;
    layer5_outputs(1459) <= a or b;
    layer5_outputs(1460) <= not b;
    layer5_outputs(1461) <= not b or a;
    layer5_outputs(1462) <= a;
    layer5_outputs(1463) <= not a;
    layer5_outputs(1464) <= a or b;
    layer5_outputs(1465) <= not (a and b);
    layer5_outputs(1466) <= not b;
    layer5_outputs(1467) <= not b;
    layer5_outputs(1468) <= b;
    layer5_outputs(1469) <= a and not b;
    layer5_outputs(1470) <= a xor b;
    layer5_outputs(1471) <= a;
    layer5_outputs(1472) <= a;
    layer5_outputs(1473) <= a;
    layer5_outputs(1474) <= a;
    layer5_outputs(1475) <= not a or b;
    layer5_outputs(1476) <= not b;
    layer5_outputs(1477) <= not b;
    layer5_outputs(1478) <= not (a or b);
    layer5_outputs(1479) <= not (a and b);
    layer5_outputs(1480) <= not a;
    layer5_outputs(1481) <= b;
    layer5_outputs(1482) <= a xor b;
    layer5_outputs(1483) <= not (a or b);
    layer5_outputs(1484) <= a and not b;
    layer5_outputs(1485) <= a;
    layer5_outputs(1486) <= a xor b;
    layer5_outputs(1487) <= not a;
    layer5_outputs(1488) <= a and b;
    layer5_outputs(1489) <= not b;
    layer5_outputs(1490) <= not b;
    layer5_outputs(1491) <= a and b;
    layer5_outputs(1492) <= not b or a;
    layer5_outputs(1493) <= not (a xor b);
    layer5_outputs(1494) <= not (a or b);
    layer5_outputs(1495) <= b and not a;
    layer5_outputs(1496) <= a;
    layer5_outputs(1497) <= not a or b;
    layer5_outputs(1498) <= not (a and b);
    layer5_outputs(1499) <= not a;
    layer5_outputs(1500) <= a xor b;
    layer5_outputs(1501) <= a and b;
    layer5_outputs(1502) <= b;
    layer5_outputs(1503) <= not a or b;
    layer5_outputs(1504) <= b;
    layer5_outputs(1505) <= a and b;
    layer5_outputs(1506) <= a or b;
    layer5_outputs(1507) <= a;
    layer5_outputs(1508) <= not (a xor b);
    layer5_outputs(1509) <= not (a xor b);
    layer5_outputs(1510) <= not a;
    layer5_outputs(1511) <= not b;
    layer5_outputs(1512) <= b and not a;
    layer5_outputs(1513) <= not a;
    layer5_outputs(1514) <= not (a or b);
    layer5_outputs(1515) <= not b;
    layer5_outputs(1516) <= b;
    layer5_outputs(1517) <= not a;
    layer5_outputs(1518) <= a;
    layer5_outputs(1519) <= b;
    layer5_outputs(1520) <= not b;
    layer5_outputs(1521) <= a and not b;
    layer5_outputs(1522) <= b;
    layer5_outputs(1523) <= b and not a;
    layer5_outputs(1524) <= not b;
    layer5_outputs(1525) <= a or b;
    layer5_outputs(1526) <= not b or a;
    layer5_outputs(1527) <= a;
    layer5_outputs(1528) <= not (a and b);
    layer5_outputs(1529) <= not a or b;
    layer5_outputs(1530) <= not (a xor b);
    layer5_outputs(1531) <= a and b;
    layer5_outputs(1532) <= a and b;
    layer5_outputs(1533) <= not a;
    layer5_outputs(1534) <= a;
    layer5_outputs(1535) <= not b;
    layer5_outputs(1536) <= not b;
    layer5_outputs(1537) <= not b or a;
    layer5_outputs(1538) <= a;
    layer5_outputs(1539) <= '0';
    layer5_outputs(1540) <= a or b;
    layer5_outputs(1541) <= not b;
    layer5_outputs(1542) <= b;
    layer5_outputs(1543) <= not b;
    layer5_outputs(1544) <= b;
    layer5_outputs(1545) <= not a;
    layer5_outputs(1546) <= not b;
    layer5_outputs(1547) <= a and not b;
    layer5_outputs(1548) <= not b;
    layer5_outputs(1549) <= a;
    layer5_outputs(1550) <= a and not b;
    layer5_outputs(1551) <= not (a or b);
    layer5_outputs(1552) <= a and not b;
    layer5_outputs(1553) <= not (a xor b);
    layer5_outputs(1554) <= a and b;
    layer5_outputs(1555) <= a xor b;
    layer5_outputs(1556) <= not a;
    layer5_outputs(1557) <= a and not b;
    layer5_outputs(1558) <= not (a xor b);
    layer5_outputs(1559) <= b;
    layer5_outputs(1560) <= not a or b;
    layer5_outputs(1561) <= a or b;
    layer5_outputs(1562) <= not a or b;
    layer5_outputs(1563) <= a xor b;
    layer5_outputs(1564) <= a or b;
    layer5_outputs(1565) <= not (a xor b);
    layer5_outputs(1566) <= not a;
    layer5_outputs(1567) <= a xor b;
    layer5_outputs(1568) <= not b or a;
    layer5_outputs(1569) <= a xor b;
    layer5_outputs(1570) <= '1';
    layer5_outputs(1571) <= '1';
    layer5_outputs(1572) <= not (a and b);
    layer5_outputs(1573) <= not b;
    layer5_outputs(1574) <= a;
    layer5_outputs(1575) <= not a;
    layer5_outputs(1576) <= a xor b;
    layer5_outputs(1577) <= a or b;
    layer5_outputs(1578) <= not (a xor b);
    layer5_outputs(1579) <= not a;
    layer5_outputs(1580) <= not a or b;
    layer5_outputs(1581) <= not b;
    layer5_outputs(1582) <= not a;
    layer5_outputs(1583) <= a and not b;
    layer5_outputs(1584) <= a and not b;
    layer5_outputs(1585) <= not a or b;
    layer5_outputs(1586) <= a and not b;
    layer5_outputs(1587) <= a xor b;
    layer5_outputs(1588) <= a;
    layer5_outputs(1589) <= not b;
    layer5_outputs(1590) <= not a;
    layer5_outputs(1591) <= b;
    layer5_outputs(1592) <= a and not b;
    layer5_outputs(1593) <= b and not a;
    layer5_outputs(1594) <= not a;
    layer5_outputs(1595) <= not b;
    layer5_outputs(1596) <= a xor b;
    layer5_outputs(1597) <= b and not a;
    layer5_outputs(1598) <= a and b;
    layer5_outputs(1599) <= not b;
    layer5_outputs(1600) <= a or b;
    layer5_outputs(1601) <= b;
    layer5_outputs(1602) <= '0';
    layer5_outputs(1603) <= a;
    layer5_outputs(1604) <= not a or b;
    layer5_outputs(1605) <= not b or a;
    layer5_outputs(1606) <= not a;
    layer5_outputs(1607) <= b;
    layer5_outputs(1608) <= b;
    layer5_outputs(1609) <= a or b;
    layer5_outputs(1610) <= b;
    layer5_outputs(1611) <= not (a and b);
    layer5_outputs(1612) <= b;
    layer5_outputs(1613) <= not (a xor b);
    layer5_outputs(1614) <= not (a xor b);
    layer5_outputs(1615) <= not (a xor b);
    layer5_outputs(1616) <= b;
    layer5_outputs(1617) <= not b;
    layer5_outputs(1618) <= a xor b;
    layer5_outputs(1619) <= b;
    layer5_outputs(1620) <= not a or b;
    layer5_outputs(1621) <= a;
    layer5_outputs(1622) <= a and b;
    layer5_outputs(1623) <= not (a xor b);
    layer5_outputs(1624) <= a and b;
    layer5_outputs(1625) <= b and not a;
    layer5_outputs(1626) <= not (a xor b);
    layer5_outputs(1627) <= not b;
    layer5_outputs(1628) <= a;
    layer5_outputs(1629) <= not (a or b);
    layer5_outputs(1630) <= a;
    layer5_outputs(1631) <= a;
    layer5_outputs(1632) <= not (a xor b);
    layer5_outputs(1633) <= not b;
    layer5_outputs(1634) <= not a;
    layer5_outputs(1635) <= a xor b;
    layer5_outputs(1636) <= a xor b;
    layer5_outputs(1637) <= a xor b;
    layer5_outputs(1638) <= not a;
    layer5_outputs(1639) <= not (a xor b);
    layer5_outputs(1640) <= not (a or b);
    layer5_outputs(1641) <= not (a and b);
    layer5_outputs(1642) <= not a;
    layer5_outputs(1643) <= not (a and b);
    layer5_outputs(1644) <= not a;
    layer5_outputs(1645) <= not a;
    layer5_outputs(1646) <= not a or b;
    layer5_outputs(1647) <= not a;
    layer5_outputs(1648) <= not (a xor b);
    layer5_outputs(1649) <= a or b;
    layer5_outputs(1650) <= not (a xor b);
    layer5_outputs(1651) <= a or b;
    layer5_outputs(1652) <= not (a and b);
    layer5_outputs(1653) <= b;
    layer5_outputs(1654) <= b and not a;
    layer5_outputs(1655) <= not b;
    layer5_outputs(1656) <= not a;
    layer5_outputs(1657) <= b;
    layer5_outputs(1658) <= a and b;
    layer5_outputs(1659) <= not b;
    layer5_outputs(1660) <= not (a and b);
    layer5_outputs(1661) <= a xor b;
    layer5_outputs(1662) <= a xor b;
    layer5_outputs(1663) <= b and not a;
    layer5_outputs(1664) <= a;
    layer5_outputs(1665) <= not (a or b);
    layer5_outputs(1666) <= not a;
    layer5_outputs(1667) <= b;
    layer5_outputs(1668) <= not b or a;
    layer5_outputs(1669) <= not (a and b);
    layer5_outputs(1670) <= a or b;
    layer5_outputs(1671) <= a;
    layer5_outputs(1672) <= b;
    layer5_outputs(1673) <= a and b;
    layer5_outputs(1674) <= a and not b;
    layer5_outputs(1675) <= b;
    layer5_outputs(1676) <= a and not b;
    layer5_outputs(1677) <= a;
    layer5_outputs(1678) <= '0';
    layer5_outputs(1679) <= a;
    layer5_outputs(1680) <= a or b;
    layer5_outputs(1681) <= not b;
    layer5_outputs(1682) <= not (a and b);
    layer5_outputs(1683) <= not (a xor b);
    layer5_outputs(1684) <= not a;
    layer5_outputs(1685) <= not a;
    layer5_outputs(1686) <= a and not b;
    layer5_outputs(1687) <= a and not b;
    layer5_outputs(1688) <= a xor b;
    layer5_outputs(1689) <= a;
    layer5_outputs(1690) <= a xor b;
    layer5_outputs(1691) <= not a or b;
    layer5_outputs(1692) <= a and not b;
    layer5_outputs(1693) <= a;
    layer5_outputs(1694) <= not (a xor b);
    layer5_outputs(1695) <= a;
    layer5_outputs(1696) <= a xor b;
    layer5_outputs(1697) <= not a;
    layer5_outputs(1698) <= a and not b;
    layer5_outputs(1699) <= not b;
    layer5_outputs(1700) <= b;
    layer5_outputs(1701) <= a or b;
    layer5_outputs(1702) <= a xor b;
    layer5_outputs(1703) <= a xor b;
    layer5_outputs(1704) <= a xor b;
    layer5_outputs(1705) <= a and b;
    layer5_outputs(1706) <= not a or b;
    layer5_outputs(1707) <= not (a and b);
    layer5_outputs(1708) <= not b;
    layer5_outputs(1709) <= not (a or b);
    layer5_outputs(1710) <= a;
    layer5_outputs(1711) <= not b;
    layer5_outputs(1712) <= b and not a;
    layer5_outputs(1713) <= not b;
    layer5_outputs(1714) <= not a;
    layer5_outputs(1715) <= not (a xor b);
    layer5_outputs(1716) <= not (a or b);
    layer5_outputs(1717) <= b;
    layer5_outputs(1718) <= not (a or b);
    layer5_outputs(1719) <= a;
    layer5_outputs(1720) <= not (a xor b);
    layer5_outputs(1721) <= a and not b;
    layer5_outputs(1722) <= not (a and b);
    layer5_outputs(1723) <= not a;
    layer5_outputs(1724) <= a or b;
    layer5_outputs(1725) <= not (a xor b);
    layer5_outputs(1726) <= a or b;
    layer5_outputs(1727) <= b;
    layer5_outputs(1728) <= not (a xor b);
    layer5_outputs(1729) <= not b or a;
    layer5_outputs(1730) <= a;
    layer5_outputs(1731) <= b;
    layer5_outputs(1732) <= b;
    layer5_outputs(1733) <= not a;
    layer5_outputs(1734) <= not b;
    layer5_outputs(1735) <= not b;
    layer5_outputs(1736) <= not (a or b);
    layer5_outputs(1737) <= a and b;
    layer5_outputs(1738) <= not (a xor b);
    layer5_outputs(1739) <= a and b;
    layer5_outputs(1740) <= a;
    layer5_outputs(1741) <= not a or b;
    layer5_outputs(1742) <= '1';
    layer5_outputs(1743) <= a;
    layer5_outputs(1744) <= not (a or b);
    layer5_outputs(1745) <= b;
    layer5_outputs(1746) <= not b;
    layer5_outputs(1747) <= not b;
    layer5_outputs(1748) <= a;
    layer5_outputs(1749) <= a;
    layer5_outputs(1750) <= not a;
    layer5_outputs(1751) <= b;
    layer5_outputs(1752) <= not (a xor b);
    layer5_outputs(1753) <= a and b;
    layer5_outputs(1754) <= not a;
    layer5_outputs(1755) <= not b;
    layer5_outputs(1756) <= a and b;
    layer5_outputs(1757) <= a or b;
    layer5_outputs(1758) <= b;
    layer5_outputs(1759) <= a or b;
    layer5_outputs(1760) <= not (a or b);
    layer5_outputs(1761) <= a or b;
    layer5_outputs(1762) <= not (a xor b);
    layer5_outputs(1763) <= a;
    layer5_outputs(1764) <= not (a xor b);
    layer5_outputs(1765) <= not a;
    layer5_outputs(1766) <= not b;
    layer5_outputs(1767) <= a xor b;
    layer5_outputs(1768) <= not a;
    layer5_outputs(1769) <= a;
    layer5_outputs(1770) <= not b or a;
    layer5_outputs(1771) <= a;
    layer5_outputs(1772) <= not (a and b);
    layer5_outputs(1773) <= b;
    layer5_outputs(1774) <= a;
    layer5_outputs(1775) <= a or b;
    layer5_outputs(1776) <= b;
    layer5_outputs(1777) <= b;
    layer5_outputs(1778) <= b and not a;
    layer5_outputs(1779) <= a and not b;
    layer5_outputs(1780) <= a and b;
    layer5_outputs(1781) <= a and b;
    layer5_outputs(1782) <= a or b;
    layer5_outputs(1783) <= a and not b;
    layer5_outputs(1784) <= not (a xor b);
    layer5_outputs(1785) <= not b;
    layer5_outputs(1786) <= a and b;
    layer5_outputs(1787) <= not b;
    layer5_outputs(1788) <= a and b;
    layer5_outputs(1789) <= b;
    layer5_outputs(1790) <= a or b;
    layer5_outputs(1791) <= a;
    layer5_outputs(1792) <= a and not b;
    layer5_outputs(1793) <= a;
    layer5_outputs(1794) <= not b;
    layer5_outputs(1795) <= not (a and b);
    layer5_outputs(1796) <= a xor b;
    layer5_outputs(1797) <= not (a and b);
    layer5_outputs(1798) <= not b or a;
    layer5_outputs(1799) <= not a;
    layer5_outputs(1800) <= '0';
    layer5_outputs(1801) <= a;
    layer5_outputs(1802) <= not b;
    layer5_outputs(1803) <= not (a or b);
    layer5_outputs(1804) <= not (a and b);
    layer5_outputs(1805) <= a;
    layer5_outputs(1806) <= b;
    layer5_outputs(1807) <= not b;
    layer5_outputs(1808) <= b and not a;
    layer5_outputs(1809) <= a and b;
    layer5_outputs(1810) <= b;
    layer5_outputs(1811) <= not a or b;
    layer5_outputs(1812) <= a;
    layer5_outputs(1813) <= b;
    layer5_outputs(1814) <= a and b;
    layer5_outputs(1815) <= not b;
    layer5_outputs(1816) <= a;
    layer5_outputs(1817) <= not b;
    layer5_outputs(1818) <= not a;
    layer5_outputs(1819) <= a and not b;
    layer5_outputs(1820) <= a and not b;
    layer5_outputs(1821) <= b;
    layer5_outputs(1822) <= not a or b;
    layer5_outputs(1823) <= not a;
    layer5_outputs(1824) <= not a;
    layer5_outputs(1825) <= b;
    layer5_outputs(1826) <= not b;
    layer5_outputs(1827) <= a;
    layer5_outputs(1828) <= not (a and b);
    layer5_outputs(1829) <= a and not b;
    layer5_outputs(1830) <= a;
    layer5_outputs(1831) <= a;
    layer5_outputs(1832) <= not a;
    layer5_outputs(1833) <= a;
    layer5_outputs(1834) <= a or b;
    layer5_outputs(1835) <= not b;
    layer5_outputs(1836) <= b and not a;
    layer5_outputs(1837) <= not a or b;
    layer5_outputs(1838) <= a or b;
    layer5_outputs(1839) <= not a or b;
    layer5_outputs(1840) <= not (a and b);
    layer5_outputs(1841) <= not a;
    layer5_outputs(1842) <= not a;
    layer5_outputs(1843) <= not b;
    layer5_outputs(1844) <= a;
    layer5_outputs(1845) <= b;
    layer5_outputs(1846) <= b;
    layer5_outputs(1847) <= not b;
    layer5_outputs(1848) <= not b or a;
    layer5_outputs(1849) <= not b or a;
    layer5_outputs(1850) <= a xor b;
    layer5_outputs(1851) <= a;
    layer5_outputs(1852) <= a or b;
    layer5_outputs(1853) <= not a;
    layer5_outputs(1854) <= not b or a;
    layer5_outputs(1855) <= b and not a;
    layer5_outputs(1856) <= not (a xor b);
    layer5_outputs(1857) <= a and b;
    layer5_outputs(1858) <= not a;
    layer5_outputs(1859) <= a;
    layer5_outputs(1860) <= a xor b;
    layer5_outputs(1861) <= not (a xor b);
    layer5_outputs(1862) <= a and b;
    layer5_outputs(1863) <= not (a xor b);
    layer5_outputs(1864) <= a xor b;
    layer5_outputs(1865) <= not (a xor b);
    layer5_outputs(1866) <= not b or a;
    layer5_outputs(1867) <= not b or a;
    layer5_outputs(1868) <= '1';
    layer5_outputs(1869) <= a;
    layer5_outputs(1870) <= not a;
    layer5_outputs(1871) <= b;
    layer5_outputs(1872) <= a;
    layer5_outputs(1873) <= a;
    layer5_outputs(1874) <= not b;
    layer5_outputs(1875) <= a or b;
    layer5_outputs(1876) <= b;
    layer5_outputs(1877) <= a xor b;
    layer5_outputs(1878) <= not a;
    layer5_outputs(1879) <= not b;
    layer5_outputs(1880) <= b and not a;
    layer5_outputs(1881) <= a and not b;
    layer5_outputs(1882) <= not b;
    layer5_outputs(1883) <= a xor b;
    layer5_outputs(1884) <= a or b;
    layer5_outputs(1885) <= not a;
    layer5_outputs(1886) <= not (a or b);
    layer5_outputs(1887) <= not (a or b);
    layer5_outputs(1888) <= b;
    layer5_outputs(1889) <= not b;
    layer5_outputs(1890) <= a;
    layer5_outputs(1891) <= not (a xor b);
    layer5_outputs(1892) <= b;
    layer5_outputs(1893) <= a and not b;
    layer5_outputs(1894) <= not b;
    layer5_outputs(1895) <= not a;
    layer5_outputs(1896) <= not (a or b);
    layer5_outputs(1897) <= not a;
    layer5_outputs(1898) <= not b or a;
    layer5_outputs(1899) <= not (a xor b);
    layer5_outputs(1900) <= not (a or b);
    layer5_outputs(1901) <= a and not b;
    layer5_outputs(1902) <= a or b;
    layer5_outputs(1903) <= a or b;
    layer5_outputs(1904) <= not (a and b);
    layer5_outputs(1905) <= a and b;
    layer5_outputs(1906) <= not (a or b);
    layer5_outputs(1907) <= not a;
    layer5_outputs(1908) <= not b or a;
    layer5_outputs(1909) <= b;
    layer5_outputs(1910) <= b and not a;
    layer5_outputs(1911) <= b and not a;
    layer5_outputs(1912) <= b;
    layer5_outputs(1913) <= a xor b;
    layer5_outputs(1914) <= not a;
    layer5_outputs(1915) <= not (a and b);
    layer5_outputs(1916) <= not b;
    layer5_outputs(1917) <= not (a xor b);
    layer5_outputs(1918) <= not a or b;
    layer5_outputs(1919) <= b;
    layer5_outputs(1920) <= a or b;
    layer5_outputs(1921) <= a xor b;
    layer5_outputs(1922) <= not b;
    layer5_outputs(1923) <= not a;
    layer5_outputs(1924) <= a and b;
    layer5_outputs(1925) <= not (a or b);
    layer5_outputs(1926) <= not (a xor b);
    layer5_outputs(1927) <= not b;
    layer5_outputs(1928) <= not a;
    layer5_outputs(1929) <= not (a and b);
    layer5_outputs(1930) <= not b or a;
    layer5_outputs(1931) <= not a;
    layer5_outputs(1932) <= not a;
    layer5_outputs(1933) <= not (a and b);
    layer5_outputs(1934) <= not b or a;
    layer5_outputs(1935) <= not a or b;
    layer5_outputs(1936) <= not b;
    layer5_outputs(1937) <= a;
    layer5_outputs(1938) <= b;
    layer5_outputs(1939) <= not b;
    layer5_outputs(1940) <= not (a or b);
    layer5_outputs(1941) <= not a or b;
    layer5_outputs(1942) <= b;
    layer5_outputs(1943) <= b and not a;
    layer5_outputs(1944) <= a or b;
    layer5_outputs(1945) <= not b;
    layer5_outputs(1946) <= b and not a;
    layer5_outputs(1947) <= not b;
    layer5_outputs(1948) <= a;
    layer5_outputs(1949) <= b;
    layer5_outputs(1950) <= not b or a;
    layer5_outputs(1951) <= not b or a;
    layer5_outputs(1952) <= not (a xor b);
    layer5_outputs(1953) <= not b;
    layer5_outputs(1954) <= a and not b;
    layer5_outputs(1955) <= b;
    layer5_outputs(1956) <= b and not a;
    layer5_outputs(1957) <= a;
    layer5_outputs(1958) <= not (a xor b);
    layer5_outputs(1959) <= not (a xor b);
    layer5_outputs(1960) <= not (a xor b);
    layer5_outputs(1961) <= a and b;
    layer5_outputs(1962) <= b;
    layer5_outputs(1963) <= not a;
    layer5_outputs(1964) <= a;
    layer5_outputs(1965) <= b;
    layer5_outputs(1966) <= a or b;
    layer5_outputs(1967) <= a and b;
    layer5_outputs(1968) <= '0';
    layer5_outputs(1969) <= not b or a;
    layer5_outputs(1970) <= a;
    layer5_outputs(1971) <= a and not b;
    layer5_outputs(1972) <= not (a xor b);
    layer5_outputs(1973) <= not (a and b);
    layer5_outputs(1974) <= not a;
    layer5_outputs(1975) <= not b;
    layer5_outputs(1976) <= a and not b;
    layer5_outputs(1977) <= not b or a;
    layer5_outputs(1978) <= a;
    layer5_outputs(1979) <= a;
    layer5_outputs(1980) <= a or b;
    layer5_outputs(1981) <= a and b;
    layer5_outputs(1982) <= not b;
    layer5_outputs(1983) <= not a;
    layer5_outputs(1984) <= a;
    layer5_outputs(1985) <= not b;
    layer5_outputs(1986) <= not b;
    layer5_outputs(1987) <= b;
    layer5_outputs(1988) <= b;
    layer5_outputs(1989) <= b;
    layer5_outputs(1990) <= '1';
    layer5_outputs(1991) <= a and not b;
    layer5_outputs(1992) <= a and not b;
    layer5_outputs(1993) <= a;
    layer5_outputs(1994) <= not b;
    layer5_outputs(1995) <= not (a and b);
    layer5_outputs(1996) <= not a;
    layer5_outputs(1997) <= a and not b;
    layer5_outputs(1998) <= not (a or b);
    layer5_outputs(1999) <= not (a and b);
    layer5_outputs(2000) <= not a or b;
    layer5_outputs(2001) <= a;
    layer5_outputs(2002) <= a and b;
    layer5_outputs(2003) <= a or b;
    layer5_outputs(2004) <= a;
    layer5_outputs(2005) <= a or b;
    layer5_outputs(2006) <= b and not a;
    layer5_outputs(2007) <= b;
    layer5_outputs(2008) <= not (a xor b);
    layer5_outputs(2009) <= b;
    layer5_outputs(2010) <= a and not b;
    layer5_outputs(2011) <= a;
    layer5_outputs(2012) <= a xor b;
    layer5_outputs(2013) <= a;
    layer5_outputs(2014) <= '0';
    layer5_outputs(2015) <= not (a and b);
    layer5_outputs(2016) <= a;
    layer5_outputs(2017) <= b and not a;
    layer5_outputs(2018) <= b;
    layer5_outputs(2019) <= not (a or b);
    layer5_outputs(2020) <= a;
    layer5_outputs(2021) <= a and b;
    layer5_outputs(2022) <= '1';
    layer5_outputs(2023) <= not (a xor b);
    layer5_outputs(2024) <= not b;
    layer5_outputs(2025) <= b;
    layer5_outputs(2026) <= a or b;
    layer5_outputs(2027) <= not a or b;
    layer5_outputs(2028) <= not b;
    layer5_outputs(2029) <= a xor b;
    layer5_outputs(2030) <= b and not a;
    layer5_outputs(2031) <= not b;
    layer5_outputs(2032) <= not a;
    layer5_outputs(2033) <= not a;
    layer5_outputs(2034) <= a;
    layer5_outputs(2035) <= not (a xor b);
    layer5_outputs(2036) <= b;
    layer5_outputs(2037) <= not (a xor b);
    layer5_outputs(2038) <= a or b;
    layer5_outputs(2039) <= b and not a;
    layer5_outputs(2040) <= a or b;
    layer5_outputs(2041) <= a;
    layer5_outputs(2042) <= a and not b;
    layer5_outputs(2043) <= b;
    layer5_outputs(2044) <= not a;
    layer5_outputs(2045) <= a;
    layer5_outputs(2046) <= not b;
    layer5_outputs(2047) <= b;
    layer5_outputs(2048) <= a;
    layer5_outputs(2049) <= not (a or b);
    layer5_outputs(2050) <= not b;
    layer5_outputs(2051) <= b and not a;
    layer5_outputs(2052) <= a or b;
    layer5_outputs(2053) <= a and b;
    layer5_outputs(2054) <= not b or a;
    layer5_outputs(2055) <= a xor b;
    layer5_outputs(2056) <= not b;
    layer5_outputs(2057) <= not b;
    layer5_outputs(2058) <= not (a and b);
    layer5_outputs(2059) <= not b;
    layer5_outputs(2060) <= not a;
    layer5_outputs(2061) <= b;
    layer5_outputs(2062) <= not a or b;
    layer5_outputs(2063) <= a xor b;
    layer5_outputs(2064) <= not b;
    layer5_outputs(2065) <= a;
    layer5_outputs(2066) <= a;
    layer5_outputs(2067) <= not b or a;
    layer5_outputs(2068) <= not b or a;
    layer5_outputs(2069) <= not (a and b);
    layer5_outputs(2070) <= not b;
    layer5_outputs(2071) <= not (a xor b);
    layer5_outputs(2072) <= b and not a;
    layer5_outputs(2073) <= not a;
    layer5_outputs(2074) <= not (a or b);
    layer5_outputs(2075) <= a xor b;
    layer5_outputs(2076) <= not b or a;
    layer5_outputs(2077) <= a;
    layer5_outputs(2078) <= not (a and b);
    layer5_outputs(2079) <= a;
    layer5_outputs(2080) <= not (a and b);
    layer5_outputs(2081) <= not b;
    layer5_outputs(2082) <= a xor b;
    layer5_outputs(2083) <= a xor b;
    layer5_outputs(2084) <= b and not a;
    layer5_outputs(2085) <= not b;
    layer5_outputs(2086) <= not a;
    layer5_outputs(2087) <= b;
    layer5_outputs(2088) <= b;
    layer5_outputs(2089) <= not a;
    layer5_outputs(2090) <= not a;
    layer5_outputs(2091) <= '0';
    layer5_outputs(2092) <= not b or a;
    layer5_outputs(2093) <= not (a and b);
    layer5_outputs(2094) <= a xor b;
    layer5_outputs(2095) <= b and not a;
    layer5_outputs(2096) <= a;
    layer5_outputs(2097) <= a;
    layer5_outputs(2098) <= b and not a;
    layer5_outputs(2099) <= not a or b;
    layer5_outputs(2100) <= not (a xor b);
    layer5_outputs(2101) <= not b;
    layer5_outputs(2102) <= b;
    layer5_outputs(2103) <= b;
    layer5_outputs(2104) <= a;
    layer5_outputs(2105) <= b;
    layer5_outputs(2106) <= a;
    layer5_outputs(2107) <= not (a and b);
    layer5_outputs(2108) <= '0';
    layer5_outputs(2109) <= a;
    layer5_outputs(2110) <= b;
    layer5_outputs(2111) <= a and not b;
    layer5_outputs(2112) <= not (a or b);
    layer5_outputs(2113) <= a;
    layer5_outputs(2114) <= b;
    layer5_outputs(2115) <= a;
    layer5_outputs(2116) <= b and not a;
    layer5_outputs(2117) <= not a or b;
    layer5_outputs(2118) <= not b;
    layer5_outputs(2119) <= a xor b;
    layer5_outputs(2120) <= not a;
    layer5_outputs(2121) <= not (a xor b);
    layer5_outputs(2122) <= not b;
    layer5_outputs(2123) <= not (a or b);
    layer5_outputs(2124) <= a;
    layer5_outputs(2125) <= not b;
    layer5_outputs(2126) <= a xor b;
    layer5_outputs(2127) <= not b or a;
    layer5_outputs(2128) <= not b or a;
    layer5_outputs(2129) <= not b;
    layer5_outputs(2130) <= not b or a;
    layer5_outputs(2131) <= not b;
    layer5_outputs(2132) <= b;
    layer5_outputs(2133) <= a;
    layer5_outputs(2134) <= b and not a;
    layer5_outputs(2135) <= not (a xor b);
    layer5_outputs(2136) <= not (a xor b);
    layer5_outputs(2137) <= a;
    layer5_outputs(2138) <= a xor b;
    layer5_outputs(2139) <= not (a xor b);
    layer5_outputs(2140) <= not a or b;
    layer5_outputs(2141) <= a and not b;
    layer5_outputs(2142) <= b and not a;
    layer5_outputs(2143) <= a;
    layer5_outputs(2144) <= a and b;
    layer5_outputs(2145) <= not (a or b);
    layer5_outputs(2146) <= a and b;
    layer5_outputs(2147) <= not b;
    layer5_outputs(2148) <= a or b;
    layer5_outputs(2149) <= a xor b;
    layer5_outputs(2150) <= not b;
    layer5_outputs(2151) <= b;
    layer5_outputs(2152) <= a or b;
    layer5_outputs(2153) <= not a;
    layer5_outputs(2154) <= a and b;
    layer5_outputs(2155) <= not a;
    layer5_outputs(2156) <= b;
    layer5_outputs(2157) <= not a;
    layer5_outputs(2158) <= not (a or b);
    layer5_outputs(2159) <= b;
    layer5_outputs(2160) <= a;
    layer5_outputs(2161) <= not b;
    layer5_outputs(2162) <= not a;
    layer5_outputs(2163) <= not b;
    layer5_outputs(2164) <= not b;
    layer5_outputs(2165) <= not b or a;
    layer5_outputs(2166) <= '0';
    layer5_outputs(2167) <= not b;
    layer5_outputs(2168) <= a;
    layer5_outputs(2169) <= not b or a;
    layer5_outputs(2170) <= b;
    layer5_outputs(2171) <= not a or b;
    layer5_outputs(2172) <= a;
    layer5_outputs(2173) <= not a;
    layer5_outputs(2174) <= a or b;
    layer5_outputs(2175) <= a xor b;
    layer5_outputs(2176) <= a;
    layer5_outputs(2177) <= not (a xor b);
    layer5_outputs(2178) <= not b or a;
    layer5_outputs(2179) <= not b;
    layer5_outputs(2180) <= not (a xor b);
    layer5_outputs(2181) <= not (a xor b);
    layer5_outputs(2182) <= not b;
    layer5_outputs(2183) <= a xor b;
    layer5_outputs(2184) <= b;
    layer5_outputs(2185) <= not b;
    layer5_outputs(2186) <= not (a xor b);
    layer5_outputs(2187) <= not (a and b);
    layer5_outputs(2188) <= b;
    layer5_outputs(2189) <= not a;
    layer5_outputs(2190) <= not b;
    layer5_outputs(2191) <= not (a and b);
    layer5_outputs(2192) <= not b;
    layer5_outputs(2193) <= not a or b;
    layer5_outputs(2194) <= not b;
    layer5_outputs(2195) <= not b;
    layer5_outputs(2196) <= not (a and b);
    layer5_outputs(2197) <= b;
    layer5_outputs(2198) <= a;
    layer5_outputs(2199) <= not a;
    layer5_outputs(2200) <= a;
    layer5_outputs(2201) <= a xor b;
    layer5_outputs(2202) <= not a;
    layer5_outputs(2203) <= not b;
    layer5_outputs(2204) <= not a or b;
    layer5_outputs(2205) <= a and b;
    layer5_outputs(2206) <= b;
    layer5_outputs(2207) <= not a;
    layer5_outputs(2208) <= a and b;
    layer5_outputs(2209) <= not b or a;
    layer5_outputs(2210) <= not b or a;
    layer5_outputs(2211) <= a xor b;
    layer5_outputs(2212) <= a or b;
    layer5_outputs(2213) <= a xor b;
    layer5_outputs(2214) <= not (a and b);
    layer5_outputs(2215) <= a xor b;
    layer5_outputs(2216) <= not (a xor b);
    layer5_outputs(2217) <= not (a xor b);
    layer5_outputs(2218) <= a xor b;
    layer5_outputs(2219) <= b;
    layer5_outputs(2220) <= b;
    layer5_outputs(2221) <= not a or b;
    layer5_outputs(2222) <= a;
    layer5_outputs(2223) <= not (a and b);
    layer5_outputs(2224) <= not (a xor b);
    layer5_outputs(2225) <= b and not a;
    layer5_outputs(2226) <= b and not a;
    layer5_outputs(2227) <= not (a or b);
    layer5_outputs(2228) <= not b;
    layer5_outputs(2229) <= a;
    layer5_outputs(2230) <= b;
    layer5_outputs(2231) <= not (a and b);
    layer5_outputs(2232) <= not b;
    layer5_outputs(2233) <= not (a and b);
    layer5_outputs(2234) <= a and not b;
    layer5_outputs(2235) <= b;
    layer5_outputs(2236) <= b;
    layer5_outputs(2237) <= not (a xor b);
    layer5_outputs(2238) <= not (a or b);
    layer5_outputs(2239) <= a or b;
    layer5_outputs(2240) <= not a;
    layer5_outputs(2241) <= b;
    layer5_outputs(2242) <= a or b;
    layer5_outputs(2243) <= a or b;
    layer5_outputs(2244) <= not a;
    layer5_outputs(2245) <= '1';
    layer5_outputs(2246) <= b;
    layer5_outputs(2247) <= b;
    layer5_outputs(2248) <= a xor b;
    layer5_outputs(2249) <= b and not a;
    layer5_outputs(2250) <= not b;
    layer5_outputs(2251) <= not (a or b);
    layer5_outputs(2252) <= a or b;
    layer5_outputs(2253) <= a xor b;
    layer5_outputs(2254) <= a;
    layer5_outputs(2255) <= a;
    layer5_outputs(2256) <= b;
    layer5_outputs(2257) <= '1';
    layer5_outputs(2258) <= b and not a;
    layer5_outputs(2259) <= not b;
    layer5_outputs(2260) <= a xor b;
    layer5_outputs(2261) <= not b;
    layer5_outputs(2262) <= not b;
    layer5_outputs(2263) <= not (a and b);
    layer5_outputs(2264) <= b and not a;
    layer5_outputs(2265) <= not a;
    layer5_outputs(2266) <= b and not a;
    layer5_outputs(2267) <= not b;
    layer5_outputs(2268) <= not a;
    layer5_outputs(2269) <= a and b;
    layer5_outputs(2270) <= a and b;
    layer5_outputs(2271) <= not (a xor b);
    layer5_outputs(2272) <= '0';
    layer5_outputs(2273) <= b;
    layer5_outputs(2274) <= b;
    layer5_outputs(2275) <= b and not a;
    layer5_outputs(2276) <= b;
    layer5_outputs(2277) <= b;
    layer5_outputs(2278) <= not b;
    layer5_outputs(2279) <= not b;
    layer5_outputs(2280) <= a xor b;
    layer5_outputs(2281) <= not a or b;
    layer5_outputs(2282) <= not (a and b);
    layer5_outputs(2283) <= not b;
    layer5_outputs(2284) <= not (a or b);
    layer5_outputs(2285) <= not a;
    layer5_outputs(2286) <= not (a xor b);
    layer5_outputs(2287) <= not b;
    layer5_outputs(2288) <= not (a and b);
    layer5_outputs(2289) <= not b or a;
    layer5_outputs(2290) <= not a or b;
    layer5_outputs(2291) <= not a;
    layer5_outputs(2292) <= not (a and b);
    layer5_outputs(2293) <= b;
    layer5_outputs(2294) <= a or b;
    layer5_outputs(2295) <= not (a xor b);
    layer5_outputs(2296) <= not a or b;
    layer5_outputs(2297) <= not a;
    layer5_outputs(2298) <= a xor b;
    layer5_outputs(2299) <= b;
    layer5_outputs(2300) <= a and b;
    layer5_outputs(2301) <= not (a or b);
    layer5_outputs(2302) <= a and b;
    layer5_outputs(2303) <= not a or b;
    layer5_outputs(2304) <= not (a xor b);
    layer5_outputs(2305) <= a;
    layer5_outputs(2306) <= not (a or b);
    layer5_outputs(2307) <= a and b;
    layer5_outputs(2308) <= not (a and b);
    layer5_outputs(2309) <= b;
    layer5_outputs(2310) <= not b;
    layer5_outputs(2311) <= not a;
    layer5_outputs(2312) <= a and not b;
    layer5_outputs(2313) <= b and not a;
    layer5_outputs(2314) <= a and b;
    layer5_outputs(2315) <= not (a xor b);
    layer5_outputs(2316) <= not b;
    layer5_outputs(2317) <= a;
    layer5_outputs(2318) <= not a or b;
    layer5_outputs(2319) <= a xor b;
    layer5_outputs(2320) <= not a;
    layer5_outputs(2321) <= b;
    layer5_outputs(2322) <= b;
    layer5_outputs(2323) <= a and not b;
    layer5_outputs(2324) <= a and not b;
    layer5_outputs(2325) <= not b or a;
    layer5_outputs(2326) <= not a or b;
    layer5_outputs(2327) <= a;
    layer5_outputs(2328) <= not b;
    layer5_outputs(2329) <= not a or b;
    layer5_outputs(2330) <= b and not a;
    layer5_outputs(2331) <= b;
    layer5_outputs(2332) <= not b;
    layer5_outputs(2333) <= not a;
    layer5_outputs(2334) <= a and b;
    layer5_outputs(2335) <= not a;
    layer5_outputs(2336) <= b;
    layer5_outputs(2337) <= not a or b;
    layer5_outputs(2338) <= b and not a;
    layer5_outputs(2339) <= not (a xor b);
    layer5_outputs(2340) <= not a or b;
    layer5_outputs(2341) <= a;
    layer5_outputs(2342) <= a or b;
    layer5_outputs(2343) <= a;
    layer5_outputs(2344) <= not (a and b);
    layer5_outputs(2345) <= a xor b;
    layer5_outputs(2346) <= not b;
    layer5_outputs(2347) <= not (a and b);
    layer5_outputs(2348) <= b;
    layer5_outputs(2349) <= not (a xor b);
    layer5_outputs(2350) <= not b;
    layer5_outputs(2351) <= a;
    layer5_outputs(2352) <= not (a and b);
    layer5_outputs(2353) <= not b;
    layer5_outputs(2354) <= a xor b;
    layer5_outputs(2355) <= not (a xor b);
    layer5_outputs(2356) <= not (a and b);
    layer5_outputs(2357) <= a xor b;
    layer5_outputs(2358) <= a and b;
    layer5_outputs(2359) <= not a or b;
    layer5_outputs(2360) <= not b or a;
    layer5_outputs(2361) <= not (a xor b);
    layer5_outputs(2362) <= b;
    layer5_outputs(2363) <= a or b;
    layer5_outputs(2364) <= not a;
    layer5_outputs(2365) <= a;
    layer5_outputs(2366) <= not a;
    layer5_outputs(2367) <= a;
    layer5_outputs(2368) <= '0';
    layer5_outputs(2369) <= not a;
    layer5_outputs(2370) <= not a;
    layer5_outputs(2371) <= '0';
    layer5_outputs(2372) <= b;
    layer5_outputs(2373) <= a or b;
    layer5_outputs(2374) <= a xor b;
    layer5_outputs(2375) <= a xor b;
    layer5_outputs(2376) <= a xor b;
    layer5_outputs(2377) <= not (a and b);
    layer5_outputs(2378) <= not a;
    layer5_outputs(2379) <= not (a xor b);
    layer5_outputs(2380) <= not b or a;
    layer5_outputs(2381) <= not a;
    layer5_outputs(2382) <= not b;
    layer5_outputs(2383) <= a;
    layer5_outputs(2384) <= not a;
    layer5_outputs(2385) <= not b or a;
    layer5_outputs(2386) <= not b;
    layer5_outputs(2387) <= a;
    layer5_outputs(2388) <= not b;
    layer5_outputs(2389) <= a xor b;
    layer5_outputs(2390) <= a xor b;
    layer5_outputs(2391) <= a xor b;
    layer5_outputs(2392) <= a;
    layer5_outputs(2393) <= not b;
    layer5_outputs(2394) <= not b or a;
    layer5_outputs(2395) <= b;
    layer5_outputs(2396) <= not (a xor b);
    layer5_outputs(2397) <= not b;
    layer5_outputs(2398) <= a or b;
    layer5_outputs(2399) <= a;
    layer5_outputs(2400) <= not b;
    layer5_outputs(2401) <= a xor b;
    layer5_outputs(2402) <= a;
    layer5_outputs(2403) <= not b;
    layer5_outputs(2404) <= not (a or b);
    layer5_outputs(2405) <= not (a or b);
    layer5_outputs(2406) <= not (a or b);
    layer5_outputs(2407) <= b;
    layer5_outputs(2408) <= a xor b;
    layer5_outputs(2409) <= not (a or b);
    layer5_outputs(2410) <= not (a xor b);
    layer5_outputs(2411) <= not b;
    layer5_outputs(2412) <= a xor b;
    layer5_outputs(2413) <= not (a and b);
    layer5_outputs(2414) <= b and not a;
    layer5_outputs(2415) <= not b;
    layer5_outputs(2416) <= a;
    layer5_outputs(2417) <= not b;
    layer5_outputs(2418) <= not (a xor b);
    layer5_outputs(2419) <= not a or b;
    layer5_outputs(2420) <= a xor b;
    layer5_outputs(2421) <= not a or b;
    layer5_outputs(2422) <= not b or a;
    layer5_outputs(2423) <= a and not b;
    layer5_outputs(2424) <= a and not b;
    layer5_outputs(2425) <= b;
    layer5_outputs(2426) <= a;
    layer5_outputs(2427) <= a;
    layer5_outputs(2428) <= a and b;
    layer5_outputs(2429) <= '0';
    layer5_outputs(2430) <= a xor b;
    layer5_outputs(2431) <= not a;
    layer5_outputs(2432) <= not b;
    layer5_outputs(2433) <= not b or a;
    layer5_outputs(2434) <= a;
    layer5_outputs(2435) <= not (a and b);
    layer5_outputs(2436) <= b;
    layer5_outputs(2437) <= not a;
    layer5_outputs(2438) <= b;
    layer5_outputs(2439) <= not b or a;
    layer5_outputs(2440) <= not (a and b);
    layer5_outputs(2441) <= not a;
    layer5_outputs(2442) <= a;
    layer5_outputs(2443) <= not a;
    layer5_outputs(2444) <= a;
    layer5_outputs(2445) <= a or b;
    layer5_outputs(2446) <= a and b;
    layer5_outputs(2447) <= not b;
    layer5_outputs(2448) <= a xor b;
    layer5_outputs(2449) <= not a or b;
    layer5_outputs(2450) <= not a;
    layer5_outputs(2451) <= not (a or b);
    layer5_outputs(2452) <= not (a xor b);
    layer5_outputs(2453) <= b;
    layer5_outputs(2454) <= b and not a;
    layer5_outputs(2455) <= a;
    layer5_outputs(2456) <= not (a or b);
    layer5_outputs(2457) <= a;
    layer5_outputs(2458) <= not a;
    layer5_outputs(2459) <= b;
    layer5_outputs(2460) <= b and not a;
    layer5_outputs(2461) <= not (a xor b);
    layer5_outputs(2462) <= not (a xor b);
    layer5_outputs(2463) <= not a or b;
    layer5_outputs(2464) <= a;
    layer5_outputs(2465) <= not (a or b);
    layer5_outputs(2466) <= a;
    layer5_outputs(2467) <= not a;
    layer5_outputs(2468) <= a and b;
    layer5_outputs(2469) <= b;
    layer5_outputs(2470) <= not a;
    layer5_outputs(2471) <= not b;
    layer5_outputs(2472) <= not b or a;
    layer5_outputs(2473) <= not (a xor b);
    layer5_outputs(2474) <= not b;
    layer5_outputs(2475) <= not (a xor b);
    layer5_outputs(2476) <= a or b;
    layer5_outputs(2477) <= a and b;
    layer5_outputs(2478) <= not a;
    layer5_outputs(2479) <= a and not b;
    layer5_outputs(2480) <= a;
    layer5_outputs(2481) <= not b or a;
    layer5_outputs(2482) <= not b;
    layer5_outputs(2483) <= not b;
    layer5_outputs(2484) <= a or b;
    layer5_outputs(2485) <= not a or b;
    layer5_outputs(2486) <= not a;
    layer5_outputs(2487) <= b;
    layer5_outputs(2488) <= not b;
    layer5_outputs(2489) <= not (a xor b);
    layer5_outputs(2490) <= a and b;
    layer5_outputs(2491) <= a;
    layer5_outputs(2492) <= not a;
    layer5_outputs(2493) <= not b;
    layer5_outputs(2494) <= a and b;
    layer5_outputs(2495) <= b;
    layer5_outputs(2496) <= not b;
    layer5_outputs(2497) <= not b;
    layer5_outputs(2498) <= a xor b;
    layer5_outputs(2499) <= b;
    layer5_outputs(2500) <= b;
    layer5_outputs(2501) <= a;
    layer5_outputs(2502) <= not a;
    layer5_outputs(2503) <= b;
    layer5_outputs(2504) <= not a;
    layer5_outputs(2505) <= not b;
    layer5_outputs(2506) <= a and not b;
    layer5_outputs(2507) <= not (a or b);
    layer5_outputs(2508) <= b and not a;
    layer5_outputs(2509) <= not b;
    layer5_outputs(2510) <= a;
    layer5_outputs(2511) <= b and not a;
    layer5_outputs(2512) <= b and not a;
    layer5_outputs(2513) <= not a;
    layer5_outputs(2514) <= a;
    layer5_outputs(2515) <= not (a and b);
    layer5_outputs(2516) <= not a;
    layer5_outputs(2517) <= not b;
    layer5_outputs(2518) <= b;
    layer5_outputs(2519) <= not (a or b);
    layer5_outputs(2520) <= not a;
    layer5_outputs(2521) <= not a or b;
    layer5_outputs(2522) <= not a;
    layer5_outputs(2523) <= not (a xor b);
    layer5_outputs(2524) <= a;
    layer5_outputs(2525) <= not b;
    layer5_outputs(2526) <= a and b;
    layer5_outputs(2527) <= b;
    layer5_outputs(2528) <= a xor b;
    layer5_outputs(2529) <= not a;
    layer5_outputs(2530) <= not b;
    layer5_outputs(2531) <= b;
    layer5_outputs(2532) <= not a;
    layer5_outputs(2533) <= a;
    layer5_outputs(2534) <= not a;
    layer5_outputs(2535) <= not b;
    layer5_outputs(2536) <= a;
    layer5_outputs(2537) <= b;
    layer5_outputs(2538) <= not b or a;
    layer5_outputs(2539) <= a and b;
    layer5_outputs(2540) <= not (a or b);
    layer5_outputs(2541) <= a or b;
    layer5_outputs(2542) <= a or b;
    layer5_outputs(2543) <= not (a or b);
    layer5_outputs(2544) <= a or b;
    layer5_outputs(2545) <= not b;
    layer5_outputs(2546) <= b;
    layer5_outputs(2547) <= a xor b;
    layer5_outputs(2548) <= not (a xor b);
    layer5_outputs(2549) <= a xor b;
    layer5_outputs(2550) <= b;
    layer5_outputs(2551) <= a;
    layer5_outputs(2552) <= a xor b;
    layer5_outputs(2553) <= not (a and b);
    layer5_outputs(2554) <= b;
    layer5_outputs(2555) <= b;
    layer5_outputs(2556) <= not a;
    layer5_outputs(2557) <= not b;
    layer5_outputs(2558) <= not a or b;
    layer5_outputs(2559) <= b;
    layer5_outputs(2560) <= b;
    layer5_outputs(2561) <= a xor b;
    layer5_outputs(2562) <= not a or b;
    layer5_outputs(2563) <= a and not b;
    layer5_outputs(2564) <= a and b;
    layer5_outputs(2565) <= not b or a;
    layer5_outputs(2566) <= not a;
    layer5_outputs(2567) <= b and not a;
    layer5_outputs(2568) <= a;
    layer5_outputs(2569) <= not (a and b);
    layer5_outputs(2570) <= a;
    layer5_outputs(2571) <= '1';
    layer5_outputs(2572) <= not b;
    layer5_outputs(2573) <= a xor b;
    layer5_outputs(2574) <= b;
    layer5_outputs(2575) <= '0';
    layer5_outputs(2576) <= not b;
    layer5_outputs(2577) <= not a;
    layer5_outputs(2578) <= not a;
    layer5_outputs(2579) <= not b;
    layer5_outputs(2580) <= not b;
    layer5_outputs(2581) <= not a;
    layer5_outputs(2582) <= b;
    layer5_outputs(2583) <= not b or a;
    layer5_outputs(2584) <= a;
    layer5_outputs(2585) <= a;
    layer5_outputs(2586) <= not (a or b);
    layer5_outputs(2587) <= not (a or b);
    layer5_outputs(2588) <= not b;
    layer5_outputs(2589) <= not (a or b);
    layer5_outputs(2590) <= a xor b;
    layer5_outputs(2591) <= not a;
    layer5_outputs(2592) <= a xor b;
    layer5_outputs(2593) <= not b;
    layer5_outputs(2594) <= not b or a;
    layer5_outputs(2595) <= a or b;
    layer5_outputs(2596) <= not b;
    layer5_outputs(2597) <= a xor b;
    layer5_outputs(2598) <= a and b;
    layer5_outputs(2599) <= a or b;
    layer5_outputs(2600) <= a;
    layer5_outputs(2601) <= '1';
    layer5_outputs(2602) <= a and b;
    layer5_outputs(2603) <= not (a or b);
    layer5_outputs(2604) <= not (a xor b);
    layer5_outputs(2605) <= a;
    layer5_outputs(2606) <= a and b;
    layer5_outputs(2607) <= a and not b;
    layer5_outputs(2608) <= not b;
    layer5_outputs(2609) <= not a;
    layer5_outputs(2610) <= a;
    layer5_outputs(2611) <= a;
    layer5_outputs(2612) <= a;
    layer5_outputs(2613) <= b and not a;
    layer5_outputs(2614) <= not b;
    layer5_outputs(2615) <= a and not b;
    layer5_outputs(2616) <= a or b;
    layer5_outputs(2617) <= not (a or b);
    layer5_outputs(2618) <= a xor b;
    layer5_outputs(2619) <= not b;
    layer5_outputs(2620) <= a;
    layer5_outputs(2621) <= a xor b;
    layer5_outputs(2622) <= not (a xor b);
    layer5_outputs(2623) <= b;
    layer5_outputs(2624) <= a or b;
    layer5_outputs(2625) <= not b;
    layer5_outputs(2626) <= a;
    layer5_outputs(2627) <= not (a xor b);
    layer5_outputs(2628) <= not b;
    layer5_outputs(2629) <= not (a and b);
    layer5_outputs(2630) <= a xor b;
    layer5_outputs(2631) <= '1';
    layer5_outputs(2632) <= b;
    layer5_outputs(2633) <= a and not b;
    layer5_outputs(2634) <= a;
    layer5_outputs(2635) <= not b or a;
    layer5_outputs(2636) <= b;
    layer5_outputs(2637) <= not b or a;
    layer5_outputs(2638) <= b;
    layer5_outputs(2639) <= a and b;
    layer5_outputs(2640) <= not a;
    layer5_outputs(2641) <= not (a xor b);
    layer5_outputs(2642) <= a;
    layer5_outputs(2643) <= not (a and b);
    layer5_outputs(2644) <= not b;
    layer5_outputs(2645) <= b and not a;
    layer5_outputs(2646) <= a;
    layer5_outputs(2647) <= b;
    layer5_outputs(2648) <= not a;
    layer5_outputs(2649) <= b;
    layer5_outputs(2650) <= not b;
    layer5_outputs(2651) <= a or b;
    layer5_outputs(2652) <= not a or b;
    layer5_outputs(2653) <= a and not b;
    layer5_outputs(2654) <= a;
    layer5_outputs(2655) <= not (a and b);
    layer5_outputs(2656) <= not (a or b);
    layer5_outputs(2657) <= not b or a;
    layer5_outputs(2658) <= not a;
    layer5_outputs(2659) <= a and not b;
    layer5_outputs(2660) <= not b;
    layer5_outputs(2661) <= a;
    layer5_outputs(2662) <= b;
    layer5_outputs(2663) <= b;
    layer5_outputs(2664) <= a;
    layer5_outputs(2665) <= not a or b;
    layer5_outputs(2666) <= a;
    layer5_outputs(2667) <= a;
    layer5_outputs(2668) <= a;
    layer5_outputs(2669) <= not b;
    layer5_outputs(2670) <= a;
    layer5_outputs(2671) <= not b;
    layer5_outputs(2672) <= '1';
    layer5_outputs(2673) <= not (a and b);
    layer5_outputs(2674) <= '0';
    layer5_outputs(2675) <= not (a xor b);
    layer5_outputs(2676) <= b and not a;
    layer5_outputs(2677) <= '1';
    layer5_outputs(2678) <= not a;
    layer5_outputs(2679) <= a and b;
    layer5_outputs(2680) <= b and not a;
    layer5_outputs(2681) <= not b;
    layer5_outputs(2682) <= not (a and b);
    layer5_outputs(2683) <= not (a and b);
    layer5_outputs(2684) <= b;
    layer5_outputs(2685) <= not a or b;
    layer5_outputs(2686) <= b;
    layer5_outputs(2687) <= not b;
    layer5_outputs(2688) <= not b;
    layer5_outputs(2689) <= not a;
    layer5_outputs(2690) <= not b;
    layer5_outputs(2691) <= not a;
    layer5_outputs(2692) <= not a or b;
    layer5_outputs(2693) <= not a;
    layer5_outputs(2694) <= a and not b;
    layer5_outputs(2695) <= a and not b;
    layer5_outputs(2696) <= not (a xor b);
    layer5_outputs(2697) <= b;
    layer5_outputs(2698) <= a;
    layer5_outputs(2699) <= not (a or b);
    layer5_outputs(2700) <= b;
    layer5_outputs(2701) <= a xor b;
    layer5_outputs(2702) <= a;
    layer5_outputs(2703) <= a and not b;
    layer5_outputs(2704) <= not (a or b);
    layer5_outputs(2705) <= not (a or b);
    layer5_outputs(2706) <= not a or b;
    layer5_outputs(2707) <= not b;
    layer5_outputs(2708) <= not b;
    layer5_outputs(2709) <= not a;
    layer5_outputs(2710) <= a;
    layer5_outputs(2711) <= not (a xor b);
    layer5_outputs(2712) <= not b;
    layer5_outputs(2713) <= b;
    layer5_outputs(2714) <= a and b;
    layer5_outputs(2715) <= not a;
    layer5_outputs(2716) <= not a;
    layer5_outputs(2717) <= a xor b;
    layer5_outputs(2718) <= a xor b;
    layer5_outputs(2719) <= a and b;
    layer5_outputs(2720) <= b;
    layer5_outputs(2721) <= a and not b;
    layer5_outputs(2722) <= not b or a;
    layer5_outputs(2723) <= b;
    layer5_outputs(2724) <= not (a and b);
    layer5_outputs(2725) <= a and b;
    layer5_outputs(2726) <= not b;
    layer5_outputs(2727) <= a;
    layer5_outputs(2728) <= not a;
    layer5_outputs(2729) <= not (a xor b);
    layer5_outputs(2730) <= not b;
    layer5_outputs(2731) <= a;
    layer5_outputs(2732) <= a or b;
    layer5_outputs(2733) <= a;
    layer5_outputs(2734) <= not b;
    layer5_outputs(2735) <= b;
    layer5_outputs(2736) <= b and not a;
    layer5_outputs(2737) <= a xor b;
    layer5_outputs(2738) <= a and not b;
    layer5_outputs(2739) <= a;
    layer5_outputs(2740) <= not b;
    layer5_outputs(2741) <= a and not b;
    layer5_outputs(2742) <= b;
    layer5_outputs(2743) <= not (a or b);
    layer5_outputs(2744) <= a;
    layer5_outputs(2745) <= a;
    layer5_outputs(2746) <= not b;
    layer5_outputs(2747) <= not b;
    layer5_outputs(2748) <= b;
    layer5_outputs(2749) <= a;
    layer5_outputs(2750) <= a or b;
    layer5_outputs(2751) <= a;
    layer5_outputs(2752) <= b and not a;
    layer5_outputs(2753) <= not a;
    layer5_outputs(2754) <= not a or b;
    layer5_outputs(2755) <= not a;
    layer5_outputs(2756) <= b and not a;
    layer5_outputs(2757) <= b;
    layer5_outputs(2758) <= a;
    layer5_outputs(2759) <= b;
    layer5_outputs(2760) <= not b;
    layer5_outputs(2761) <= '0';
    layer5_outputs(2762) <= a xor b;
    layer5_outputs(2763) <= a and not b;
    layer5_outputs(2764) <= not b;
    layer5_outputs(2765) <= not a or b;
    layer5_outputs(2766) <= a and not b;
    layer5_outputs(2767) <= not a;
    layer5_outputs(2768) <= a xor b;
    layer5_outputs(2769) <= a;
    layer5_outputs(2770) <= a;
    layer5_outputs(2771) <= a;
    layer5_outputs(2772) <= a and b;
    layer5_outputs(2773) <= not b;
    layer5_outputs(2774) <= not (a or b);
    layer5_outputs(2775) <= not (a or b);
    layer5_outputs(2776) <= not a or b;
    layer5_outputs(2777) <= not b;
    layer5_outputs(2778) <= not (a xor b);
    layer5_outputs(2779) <= a xor b;
    layer5_outputs(2780) <= b;
    layer5_outputs(2781) <= a xor b;
    layer5_outputs(2782) <= not b;
    layer5_outputs(2783) <= a;
    layer5_outputs(2784) <= a and not b;
    layer5_outputs(2785) <= a and not b;
    layer5_outputs(2786) <= a or b;
    layer5_outputs(2787) <= a;
    layer5_outputs(2788) <= not b or a;
    layer5_outputs(2789) <= not b;
    layer5_outputs(2790) <= b;
    layer5_outputs(2791) <= b;
    layer5_outputs(2792) <= not a;
    layer5_outputs(2793) <= not (a and b);
    layer5_outputs(2794) <= a xor b;
    layer5_outputs(2795) <= not (a and b);
    layer5_outputs(2796) <= not (a and b);
    layer5_outputs(2797) <= a or b;
    layer5_outputs(2798) <= not b or a;
    layer5_outputs(2799) <= a;
    layer5_outputs(2800) <= not a;
    layer5_outputs(2801) <= not a;
    layer5_outputs(2802) <= not (a xor b);
    layer5_outputs(2803) <= a;
    layer5_outputs(2804) <= not a or b;
    layer5_outputs(2805) <= a;
    layer5_outputs(2806) <= b;
    layer5_outputs(2807) <= b;
    layer5_outputs(2808) <= b;
    layer5_outputs(2809) <= a;
    layer5_outputs(2810) <= a;
    layer5_outputs(2811) <= b;
    layer5_outputs(2812) <= '1';
    layer5_outputs(2813) <= b;
    layer5_outputs(2814) <= b;
    layer5_outputs(2815) <= b;
    layer5_outputs(2816) <= not a or b;
    layer5_outputs(2817) <= b;
    layer5_outputs(2818) <= not a;
    layer5_outputs(2819) <= a or b;
    layer5_outputs(2820) <= a xor b;
    layer5_outputs(2821) <= a;
    layer5_outputs(2822) <= not (a xor b);
    layer5_outputs(2823) <= a and b;
    layer5_outputs(2824) <= a xor b;
    layer5_outputs(2825) <= a;
    layer5_outputs(2826) <= not a;
    layer5_outputs(2827) <= b;
    layer5_outputs(2828) <= a xor b;
    layer5_outputs(2829) <= a;
    layer5_outputs(2830) <= b and not a;
    layer5_outputs(2831) <= not b;
    layer5_outputs(2832) <= not b;
    layer5_outputs(2833) <= not a;
    layer5_outputs(2834) <= not b or a;
    layer5_outputs(2835) <= a or b;
    layer5_outputs(2836) <= a and b;
    layer5_outputs(2837) <= a;
    layer5_outputs(2838) <= not b;
    layer5_outputs(2839) <= not a;
    layer5_outputs(2840) <= b;
    layer5_outputs(2841) <= a;
    layer5_outputs(2842) <= b and not a;
    layer5_outputs(2843) <= a xor b;
    layer5_outputs(2844) <= a and not b;
    layer5_outputs(2845) <= a and not b;
    layer5_outputs(2846) <= a;
    layer5_outputs(2847) <= not a or b;
    layer5_outputs(2848) <= b;
    layer5_outputs(2849) <= a;
    layer5_outputs(2850) <= not a;
    layer5_outputs(2851) <= b;
    layer5_outputs(2852) <= a xor b;
    layer5_outputs(2853) <= not a;
    layer5_outputs(2854) <= b;
    layer5_outputs(2855) <= b;
    layer5_outputs(2856) <= b;
    layer5_outputs(2857) <= a xor b;
    layer5_outputs(2858) <= not b or a;
    layer5_outputs(2859) <= a and b;
    layer5_outputs(2860) <= not b or a;
    layer5_outputs(2861) <= b and not a;
    layer5_outputs(2862) <= not b or a;
    layer5_outputs(2863) <= not a;
    layer5_outputs(2864) <= not b;
    layer5_outputs(2865) <= not a or b;
    layer5_outputs(2866) <= not b;
    layer5_outputs(2867) <= a and not b;
    layer5_outputs(2868) <= not (a xor b);
    layer5_outputs(2869) <= not a;
    layer5_outputs(2870) <= b;
    layer5_outputs(2871) <= a;
    layer5_outputs(2872) <= not b;
    layer5_outputs(2873) <= not a;
    layer5_outputs(2874) <= b;
    layer5_outputs(2875) <= a xor b;
    layer5_outputs(2876) <= not (a xor b);
    layer5_outputs(2877) <= b and not a;
    layer5_outputs(2878) <= a and not b;
    layer5_outputs(2879) <= '1';
    layer5_outputs(2880) <= not b;
    layer5_outputs(2881) <= a;
    layer5_outputs(2882) <= not a;
    layer5_outputs(2883) <= a;
    layer5_outputs(2884) <= not a;
    layer5_outputs(2885) <= not b;
    layer5_outputs(2886) <= not b or a;
    layer5_outputs(2887) <= not b or a;
    layer5_outputs(2888) <= a and b;
    layer5_outputs(2889) <= not a;
    layer5_outputs(2890) <= not (a xor b);
    layer5_outputs(2891) <= a or b;
    layer5_outputs(2892) <= not b or a;
    layer5_outputs(2893) <= not a;
    layer5_outputs(2894) <= not (a and b);
    layer5_outputs(2895) <= not (a and b);
    layer5_outputs(2896) <= b;
    layer5_outputs(2897) <= b;
    layer5_outputs(2898) <= a and not b;
    layer5_outputs(2899) <= a or b;
    layer5_outputs(2900) <= not (a and b);
    layer5_outputs(2901) <= not a;
    layer5_outputs(2902) <= a;
    layer5_outputs(2903) <= not (a or b);
    layer5_outputs(2904) <= b;
    layer5_outputs(2905) <= not a;
    layer5_outputs(2906) <= b;
    layer5_outputs(2907) <= not (a and b);
    layer5_outputs(2908) <= not b;
    layer5_outputs(2909) <= a;
    layer5_outputs(2910) <= '0';
    layer5_outputs(2911) <= not a;
    layer5_outputs(2912) <= b;
    layer5_outputs(2913) <= not (a xor b);
    layer5_outputs(2914) <= a;
    layer5_outputs(2915) <= a;
    layer5_outputs(2916) <= a or b;
    layer5_outputs(2917) <= not (a or b);
    layer5_outputs(2918) <= a and not b;
    layer5_outputs(2919) <= a;
    layer5_outputs(2920) <= not (a xor b);
    layer5_outputs(2921) <= a and not b;
    layer5_outputs(2922) <= not b or a;
    layer5_outputs(2923) <= b;
    layer5_outputs(2924) <= not a or b;
    layer5_outputs(2925) <= not a;
    layer5_outputs(2926) <= a or b;
    layer5_outputs(2927) <= a xor b;
    layer5_outputs(2928) <= a and not b;
    layer5_outputs(2929) <= not (a xor b);
    layer5_outputs(2930) <= a xor b;
    layer5_outputs(2931) <= b;
    layer5_outputs(2932) <= not b;
    layer5_outputs(2933) <= a;
    layer5_outputs(2934) <= a xor b;
    layer5_outputs(2935) <= not b;
    layer5_outputs(2936) <= b;
    layer5_outputs(2937) <= not (a or b);
    layer5_outputs(2938) <= a or b;
    layer5_outputs(2939) <= b;
    layer5_outputs(2940) <= not (a or b);
    layer5_outputs(2941) <= not (a xor b);
    layer5_outputs(2942) <= '0';
    layer5_outputs(2943) <= not b;
    layer5_outputs(2944) <= a or b;
    layer5_outputs(2945) <= b;
    layer5_outputs(2946) <= a and not b;
    layer5_outputs(2947) <= a and b;
    layer5_outputs(2948) <= a and b;
    layer5_outputs(2949) <= a;
    layer5_outputs(2950) <= a;
    layer5_outputs(2951) <= b and not a;
    layer5_outputs(2952) <= not b;
    layer5_outputs(2953) <= a xor b;
    layer5_outputs(2954) <= a;
    layer5_outputs(2955) <= not a;
    layer5_outputs(2956) <= b;
    layer5_outputs(2957) <= not a;
    layer5_outputs(2958) <= a;
    layer5_outputs(2959) <= b and not a;
    layer5_outputs(2960) <= a and not b;
    layer5_outputs(2961) <= a;
    layer5_outputs(2962) <= not a;
    layer5_outputs(2963) <= not b or a;
    layer5_outputs(2964) <= not (a xor b);
    layer5_outputs(2965) <= not a;
    layer5_outputs(2966) <= not b;
    layer5_outputs(2967) <= a xor b;
    layer5_outputs(2968) <= b and not a;
    layer5_outputs(2969) <= not (a and b);
    layer5_outputs(2970) <= not (a xor b);
    layer5_outputs(2971) <= not b or a;
    layer5_outputs(2972) <= a and b;
    layer5_outputs(2973) <= not (a and b);
    layer5_outputs(2974) <= a or b;
    layer5_outputs(2975) <= a;
    layer5_outputs(2976) <= not (a xor b);
    layer5_outputs(2977) <= b;
    layer5_outputs(2978) <= a and b;
    layer5_outputs(2979) <= not (a or b);
    layer5_outputs(2980) <= not b or a;
    layer5_outputs(2981) <= not (a or b);
    layer5_outputs(2982) <= not (a or b);
    layer5_outputs(2983) <= not (a and b);
    layer5_outputs(2984) <= b;
    layer5_outputs(2985) <= b;
    layer5_outputs(2986) <= not a or b;
    layer5_outputs(2987) <= b;
    layer5_outputs(2988) <= not a or b;
    layer5_outputs(2989) <= not (a and b);
    layer5_outputs(2990) <= a xor b;
    layer5_outputs(2991) <= a and b;
    layer5_outputs(2992) <= a and not b;
    layer5_outputs(2993) <= not b or a;
    layer5_outputs(2994) <= b;
    layer5_outputs(2995) <= not b or a;
    layer5_outputs(2996) <= a xor b;
    layer5_outputs(2997) <= not b;
    layer5_outputs(2998) <= b;
    layer5_outputs(2999) <= not (a xor b);
    layer5_outputs(3000) <= b;
    layer5_outputs(3001) <= not b;
    layer5_outputs(3002) <= not (a or b);
    layer5_outputs(3003) <= b;
    layer5_outputs(3004) <= a and not b;
    layer5_outputs(3005) <= not a or b;
    layer5_outputs(3006) <= b;
    layer5_outputs(3007) <= not b;
    layer5_outputs(3008) <= not (a and b);
    layer5_outputs(3009) <= b;
    layer5_outputs(3010) <= b;
    layer5_outputs(3011) <= not b;
    layer5_outputs(3012) <= not (a xor b);
    layer5_outputs(3013) <= not (a and b);
    layer5_outputs(3014) <= not b or a;
    layer5_outputs(3015) <= not (a xor b);
    layer5_outputs(3016) <= not a or b;
    layer5_outputs(3017) <= a;
    layer5_outputs(3018) <= a;
    layer5_outputs(3019) <= a or b;
    layer5_outputs(3020) <= not a;
    layer5_outputs(3021) <= not (a or b);
    layer5_outputs(3022) <= not b;
    layer5_outputs(3023) <= not a;
    layer5_outputs(3024) <= a and not b;
    layer5_outputs(3025) <= a or b;
    layer5_outputs(3026) <= b;
    layer5_outputs(3027) <= not a or b;
    layer5_outputs(3028) <= a or b;
    layer5_outputs(3029) <= b;
    layer5_outputs(3030) <= a;
    layer5_outputs(3031) <= b;
    layer5_outputs(3032) <= not (a and b);
    layer5_outputs(3033) <= b;
    layer5_outputs(3034) <= not (a or b);
    layer5_outputs(3035) <= a;
    layer5_outputs(3036) <= b;
    layer5_outputs(3037) <= not (a xor b);
    layer5_outputs(3038) <= not (a xor b);
    layer5_outputs(3039) <= not a;
    layer5_outputs(3040) <= a xor b;
    layer5_outputs(3041) <= not a;
    layer5_outputs(3042) <= b and not a;
    layer5_outputs(3043) <= not (a or b);
    layer5_outputs(3044) <= b;
    layer5_outputs(3045) <= not a;
    layer5_outputs(3046) <= not a;
    layer5_outputs(3047) <= not (a or b);
    layer5_outputs(3048) <= not (a xor b);
    layer5_outputs(3049) <= not a;
    layer5_outputs(3050) <= not a;
    layer5_outputs(3051) <= not a;
    layer5_outputs(3052) <= a and not b;
    layer5_outputs(3053) <= not a;
    layer5_outputs(3054) <= not (a and b);
    layer5_outputs(3055) <= a;
    layer5_outputs(3056) <= a xor b;
    layer5_outputs(3057) <= a xor b;
    layer5_outputs(3058) <= a;
    layer5_outputs(3059) <= not (a xor b);
    layer5_outputs(3060) <= b and not a;
    layer5_outputs(3061) <= a or b;
    layer5_outputs(3062) <= b;
    layer5_outputs(3063) <= not b or a;
    layer5_outputs(3064) <= not a;
    layer5_outputs(3065) <= a;
    layer5_outputs(3066) <= not a or b;
    layer5_outputs(3067) <= b;
    layer5_outputs(3068) <= not a;
    layer5_outputs(3069) <= not (a and b);
    layer5_outputs(3070) <= a and not b;
    layer5_outputs(3071) <= not b;
    layer5_outputs(3072) <= not b or a;
    layer5_outputs(3073) <= b and not a;
    layer5_outputs(3074) <= a;
    layer5_outputs(3075) <= not a;
    layer5_outputs(3076) <= a or b;
    layer5_outputs(3077) <= b and not a;
    layer5_outputs(3078) <= not (a or b);
    layer5_outputs(3079) <= a xor b;
    layer5_outputs(3080) <= b;
    layer5_outputs(3081) <= not (a xor b);
    layer5_outputs(3082) <= b;
    layer5_outputs(3083) <= not (a and b);
    layer5_outputs(3084) <= a xor b;
    layer5_outputs(3085) <= a;
    layer5_outputs(3086) <= not a;
    layer5_outputs(3087) <= b and not a;
    layer5_outputs(3088) <= not (a xor b);
    layer5_outputs(3089) <= not (a xor b);
    layer5_outputs(3090) <= not b or a;
    layer5_outputs(3091) <= not (a xor b);
    layer5_outputs(3092) <= not (a and b);
    layer5_outputs(3093) <= not a or b;
    layer5_outputs(3094) <= b;
    layer5_outputs(3095) <= a or b;
    layer5_outputs(3096) <= b;
    layer5_outputs(3097) <= not a;
    layer5_outputs(3098) <= not (a xor b);
    layer5_outputs(3099) <= a and not b;
    layer5_outputs(3100) <= not (a and b);
    layer5_outputs(3101) <= a xor b;
    layer5_outputs(3102) <= a and not b;
    layer5_outputs(3103) <= not b;
    layer5_outputs(3104) <= a;
    layer5_outputs(3105) <= '0';
    layer5_outputs(3106) <= a;
    layer5_outputs(3107) <= a;
    layer5_outputs(3108) <= a and b;
    layer5_outputs(3109) <= '0';
    layer5_outputs(3110) <= not a or b;
    layer5_outputs(3111) <= not (a or b);
    layer5_outputs(3112) <= a or b;
    layer5_outputs(3113) <= a xor b;
    layer5_outputs(3114) <= not b;
    layer5_outputs(3115) <= a;
    layer5_outputs(3116) <= b;
    layer5_outputs(3117) <= a;
    layer5_outputs(3118) <= a and not b;
    layer5_outputs(3119) <= a;
    layer5_outputs(3120) <= a xor b;
    layer5_outputs(3121) <= not a;
    layer5_outputs(3122) <= not a;
    layer5_outputs(3123) <= a;
    layer5_outputs(3124) <= a and b;
    layer5_outputs(3125) <= a xor b;
    layer5_outputs(3126) <= not a;
    layer5_outputs(3127) <= not (a or b);
    layer5_outputs(3128) <= not (a xor b);
    layer5_outputs(3129) <= not (a xor b);
    layer5_outputs(3130) <= not b;
    layer5_outputs(3131) <= not a or b;
    layer5_outputs(3132) <= not b;
    layer5_outputs(3133) <= not b;
    layer5_outputs(3134) <= a and b;
    layer5_outputs(3135) <= not a;
    layer5_outputs(3136) <= a and b;
    layer5_outputs(3137) <= a or b;
    layer5_outputs(3138) <= not (a and b);
    layer5_outputs(3139) <= not b or a;
    layer5_outputs(3140) <= a and not b;
    layer5_outputs(3141) <= b;
    layer5_outputs(3142) <= a xor b;
    layer5_outputs(3143) <= a;
    layer5_outputs(3144) <= a or b;
    layer5_outputs(3145) <= not b or a;
    layer5_outputs(3146) <= not b;
    layer5_outputs(3147) <= '1';
    layer5_outputs(3148) <= b;
    layer5_outputs(3149) <= b;
    layer5_outputs(3150) <= a;
    layer5_outputs(3151) <= not a;
    layer5_outputs(3152) <= a or b;
    layer5_outputs(3153) <= not a;
    layer5_outputs(3154) <= b;
    layer5_outputs(3155) <= not (a and b);
    layer5_outputs(3156) <= a and b;
    layer5_outputs(3157) <= not b;
    layer5_outputs(3158) <= not (a and b);
    layer5_outputs(3159) <= not b or a;
    layer5_outputs(3160) <= a;
    layer5_outputs(3161) <= a;
    layer5_outputs(3162) <= not a or b;
    layer5_outputs(3163) <= b;
    layer5_outputs(3164) <= not (a xor b);
    layer5_outputs(3165) <= b;
    layer5_outputs(3166) <= not a;
    layer5_outputs(3167) <= not b;
    layer5_outputs(3168) <= not (a and b);
    layer5_outputs(3169) <= b and not a;
    layer5_outputs(3170) <= not a;
    layer5_outputs(3171) <= a;
    layer5_outputs(3172) <= not (a or b);
    layer5_outputs(3173) <= not (a and b);
    layer5_outputs(3174) <= not b;
    layer5_outputs(3175) <= not a;
    layer5_outputs(3176) <= a xor b;
    layer5_outputs(3177) <= not a;
    layer5_outputs(3178) <= a;
    layer5_outputs(3179) <= '0';
    layer5_outputs(3180) <= a or b;
    layer5_outputs(3181) <= not (a and b);
    layer5_outputs(3182) <= not a;
    layer5_outputs(3183) <= b;
    layer5_outputs(3184) <= not a;
    layer5_outputs(3185) <= '1';
    layer5_outputs(3186) <= b;
    layer5_outputs(3187) <= a;
    layer5_outputs(3188) <= a;
    layer5_outputs(3189) <= not (a or b);
    layer5_outputs(3190) <= not b;
    layer5_outputs(3191) <= a xor b;
    layer5_outputs(3192) <= not a;
    layer5_outputs(3193) <= a;
    layer5_outputs(3194) <= a and b;
    layer5_outputs(3195) <= not b;
    layer5_outputs(3196) <= a and not b;
    layer5_outputs(3197) <= not (a or b);
    layer5_outputs(3198) <= not b or a;
    layer5_outputs(3199) <= not a;
    layer5_outputs(3200) <= not a;
    layer5_outputs(3201) <= a xor b;
    layer5_outputs(3202) <= not a;
    layer5_outputs(3203) <= not b;
    layer5_outputs(3204) <= b;
    layer5_outputs(3205) <= not b;
    layer5_outputs(3206) <= b;
    layer5_outputs(3207) <= a and not b;
    layer5_outputs(3208) <= not (a and b);
    layer5_outputs(3209) <= a;
    layer5_outputs(3210) <= not (a or b);
    layer5_outputs(3211) <= not b or a;
    layer5_outputs(3212) <= not b;
    layer5_outputs(3213) <= not b;
    layer5_outputs(3214) <= not b or a;
    layer5_outputs(3215) <= a or b;
    layer5_outputs(3216) <= not a or b;
    layer5_outputs(3217) <= not a;
    layer5_outputs(3218) <= b;
    layer5_outputs(3219) <= not b;
    layer5_outputs(3220) <= not b or a;
    layer5_outputs(3221) <= not b;
    layer5_outputs(3222) <= '0';
    layer5_outputs(3223) <= not a;
    layer5_outputs(3224) <= b;
    layer5_outputs(3225) <= not b;
    layer5_outputs(3226) <= a and b;
    layer5_outputs(3227) <= a and b;
    layer5_outputs(3228) <= not b;
    layer5_outputs(3229) <= b;
    layer5_outputs(3230) <= not a;
    layer5_outputs(3231) <= b and not a;
    layer5_outputs(3232) <= not (a or b);
    layer5_outputs(3233) <= '0';
    layer5_outputs(3234) <= not b;
    layer5_outputs(3235) <= not a or b;
    layer5_outputs(3236) <= not (a and b);
    layer5_outputs(3237) <= b;
    layer5_outputs(3238) <= a xor b;
    layer5_outputs(3239) <= not (a xor b);
    layer5_outputs(3240) <= not (a and b);
    layer5_outputs(3241) <= b;
    layer5_outputs(3242) <= a;
    layer5_outputs(3243) <= not (a and b);
    layer5_outputs(3244) <= not a;
    layer5_outputs(3245) <= not (a and b);
    layer5_outputs(3246) <= not (a and b);
    layer5_outputs(3247) <= b;
    layer5_outputs(3248) <= not a;
    layer5_outputs(3249) <= not a or b;
    layer5_outputs(3250) <= a;
    layer5_outputs(3251) <= not (a xor b);
    layer5_outputs(3252) <= a and not b;
    layer5_outputs(3253) <= '0';
    layer5_outputs(3254) <= b;
    layer5_outputs(3255) <= not (a xor b);
    layer5_outputs(3256) <= not a;
    layer5_outputs(3257) <= not b;
    layer5_outputs(3258) <= not a;
    layer5_outputs(3259) <= a and not b;
    layer5_outputs(3260) <= b;
    layer5_outputs(3261) <= not a or b;
    layer5_outputs(3262) <= not a or b;
    layer5_outputs(3263) <= a and b;
    layer5_outputs(3264) <= not (a and b);
    layer5_outputs(3265) <= a;
    layer5_outputs(3266) <= not a;
    layer5_outputs(3267) <= a or b;
    layer5_outputs(3268) <= b and not a;
    layer5_outputs(3269) <= not a;
    layer5_outputs(3270) <= b;
    layer5_outputs(3271) <= not a;
    layer5_outputs(3272) <= not a;
    layer5_outputs(3273) <= not b;
    layer5_outputs(3274) <= not a or b;
    layer5_outputs(3275) <= a and not b;
    layer5_outputs(3276) <= not (a and b);
    layer5_outputs(3277) <= not (a or b);
    layer5_outputs(3278) <= not b;
    layer5_outputs(3279) <= not b;
    layer5_outputs(3280) <= b;
    layer5_outputs(3281) <= not (a or b);
    layer5_outputs(3282) <= not (a and b);
    layer5_outputs(3283) <= not (a xor b);
    layer5_outputs(3284) <= not a;
    layer5_outputs(3285) <= a;
    layer5_outputs(3286) <= not a or b;
    layer5_outputs(3287) <= not (a or b);
    layer5_outputs(3288) <= b;
    layer5_outputs(3289) <= a or b;
    layer5_outputs(3290) <= not (a and b);
    layer5_outputs(3291) <= not a;
    layer5_outputs(3292) <= not b;
    layer5_outputs(3293) <= not b;
    layer5_outputs(3294) <= a xor b;
    layer5_outputs(3295) <= not a;
    layer5_outputs(3296) <= not (a and b);
    layer5_outputs(3297) <= a;
    layer5_outputs(3298) <= not (a or b);
    layer5_outputs(3299) <= not b;
    layer5_outputs(3300) <= a;
    layer5_outputs(3301) <= not a;
    layer5_outputs(3302) <= not (a or b);
    layer5_outputs(3303) <= a and not b;
    layer5_outputs(3304) <= not (a xor b);
    layer5_outputs(3305) <= a xor b;
    layer5_outputs(3306) <= b and not a;
    layer5_outputs(3307) <= not (a xor b);
    layer5_outputs(3308) <= not a;
    layer5_outputs(3309) <= not (a and b);
    layer5_outputs(3310) <= b;
    layer5_outputs(3311) <= not a;
    layer5_outputs(3312) <= a xor b;
    layer5_outputs(3313) <= a xor b;
    layer5_outputs(3314) <= a and b;
    layer5_outputs(3315) <= b;
    layer5_outputs(3316) <= a xor b;
    layer5_outputs(3317) <= not b or a;
    layer5_outputs(3318) <= not (a and b);
    layer5_outputs(3319) <= a or b;
    layer5_outputs(3320) <= b;
    layer5_outputs(3321) <= a and b;
    layer5_outputs(3322) <= not a;
    layer5_outputs(3323) <= not b or a;
    layer5_outputs(3324) <= not b;
    layer5_outputs(3325) <= b;
    layer5_outputs(3326) <= not a or b;
    layer5_outputs(3327) <= not (a and b);
    layer5_outputs(3328) <= not b;
    layer5_outputs(3329) <= a;
    layer5_outputs(3330) <= not b;
    layer5_outputs(3331) <= b;
    layer5_outputs(3332) <= not a;
    layer5_outputs(3333) <= a;
    layer5_outputs(3334) <= b;
    layer5_outputs(3335) <= a;
    layer5_outputs(3336) <= a;
    layer5_outputs(3337) <= a or b;
    layer5_outputs(3338) <= not (a or b);
    layer5_outputs(3339) <= not a or b;
    layer5_outputs(3340) <= a and not b;
    layer5_outputs(3341) <= not b;
    layer5_outputs(3342) <= a and b;
    layer5_outputs(3343) <= not a;
    layer5_outputs(3344) <= a;
    layer5_outputs(3345) <= b;
    layer5_outputs(3346) <= a and b;
    layer5_outputs(3347) <= a or b;
    layer5_outputs(3348) <= not a;
    layer5_outputs(3349) <= not b;
    layer5_outputs(3350) <= '0';
    layer5_outputs(3351) <= not a or b;
    layer5_outputs(3352) <= not (a xor b);
    layer5_outputs(3353) <= a;
    layer5_outputs(3354) <= not (a and b);
    layer5_outputs(3355) <= a xor b;
    layer5_outputs(3356) <= not (a or b);
    layer5_outputs(3357) <= not (a or b);
    layer5_outputs(3358) <= b;
    layer5_outputs(3359) <= a;
    layer5_outputs(3360) <= not (a xor b);
    layer5_outputs(3361) <= not b;
    layer5_outputs(3362) <= b;
    layer5_outputs(3363) <= not b;
    layer5_outputs(3364) <= a or b;
    layer5_outputs(3365) <= b;
    layer5_outputs(3366) <= a;
    layer5_outputs(3367) <= a;
    layer5_outputs(3368) <= not a;
    layer5_outputs(3369) <= a xor b;
    layer5_outputs(3370) <= a or b;
    layer5_outputs(3371) <= a;
    layer5_outputs(3372) <= a;
    layer5_outputs(3373) <= not (a xor b);
    layer5_outputs(3374) <= not (a and b);
    layer5_outputs(3375) <= a or b;
    layer5_outputs(3376) <= a;
    layer5_outputs(3377) <= not b;
    layer5_outputs(3378) <= a xor b;
    layer5_outputs(3379) <= not b;
    layer5_outputs(3380) <= not (a xor b);
    layer5_outputs(3381) <= not b;
    layer5_outputs(3382) <= a;
    layer5_outputs(3383) <= not (a or b);
    layer5_outputs(3384) <= b and not a;
    layer5_outputs(3385) <= not b or a;
    layer5_outputs(3386) <= a;
    layer5_outputs(3387) <= not b;
    layer5_outputs(3388) <= a or b;
    layer5_outputs(3389) <= a;
    layer5_outputs(3390) <= a and not b;
    layer5_outputs(3391) <= a;
    layer5_outputs(3392) <= a and b;
    layer5_outputs(3393) <= a or b;
    layer5_outputs(3394) <= not b or a;
    layer5_outputs(3395) <= a;
    layer5_outputs(3396) <= not a;
    layer5_outputs(3397) <= a;
    layer5_outputs(3398) <= not (a and b);
    layer5_outputs(3399) <= not a;
    layer5_outputs(3400) <= b;
    layer5_outputs(3401) <= not (a xor b);
    layer5_outputs(3402) <= b and not a;
    layer5_outputs(3403) <= a or b;
    layer5_outputs(3404) <= not a;
    layer5_outputs(3405) <= not b;
    layer5_outputs(3406) <= not a;
    layer5_outputs(3407) <= a;
    layer5_outputs(3408) <= a;
    layer5_outputs(3409) <= b;
    layer5_outputs(3410) <= b and not a;
    layer5_outputs(3411) <= b;
    layer5_outputs(3412) <= a and b;
    layer5_outputs(3413) <= not b;
    layer5_outputs(3414) <= b and not a;
    layer5_outputs(3415) <= a;
    layer5_outputs(3416) <= b;
    layer5_outputs(3417) <= b;
    layer5_outputs(3418) <= a;
    layer5_outputs(3419) <= not (a xor b);
    layer5_outputs(3420) <= not a;
    layer5_outputs(3421) <= a xor b;
    layer5_outputs(3422) <= not a;
    layer5_outputs(3423) <= not b;
    layer5_outputs(3424) <= not (a xor b);
    layer5_outputs(3425) <= a xor b;
    layer5_outputs(3426) <= b and not a;
    layer5_outputs(3427) <= b;
    layer5_outputs(3428) <= b;
    layer5_outputs(3429) <= a or b;
    layer5_outputs(3430) <= b;
    layer5_outputs(3431) <= a and not b;
    layer5_outputs(3432) <= a xor b;
    layer5_outputs(3433) <= b;
    layer5_outputs(3434) <= '0';
    layer5_outputs(3435) <= not b or a;
    layer5_outputs(3436) <= a;
    layer5_outputs(3437) <= a;
    layer5_outputs(3438) <= a xor b;
    layer5_outputs(3439) <= not (a xor b);
    layer5_outputs(3440) <= b;
    layer5_outputs(3441) <= not b or a;
    layer5_outputs(3442) <= not a;
    layer5_outputs(3443) <= a and not b;
    layer5_outputs(3444) <= b;
    layer5_outputs(3445) <= '0';
    layer5_outputs(3446) <= a or b;
    layer5_outputs(3447) <= not b;
    layer5_outputs(3448) <= '0';
    layer5_outputs(3449) <= not (a xor b);
    layer5_outputs(3450) <= not b;
    layer5_outputs(3451) <= not a or b;
    layer5_outputs(3452) <= a xor b;
    layer5_outputs(3453) <= b;
    layer5_outputs(3454) <= b and not a;
    layer5_outputs(3455) <= a xor b;
    layer5_outputs(3456) <= a or b;
    layer5_outputs(3457) <= not (a xor b);
    layer5_outputs(3458) <= b;
    layer5_outputs(3459) <= a xor b;
    layer5_outputs(3460) <= not b;
    layer5_outputs(3461) <= not a;
    layer5_outputs(3462) <= not (a xor b);
    layer5_outputs(3463) <= a;
    layer5_outputs(3464) <= not (a xor b);
    layer5_outputs(3465) <= a;
    layer5_outputs(3466) <= not a or b;
    layer5_outputs(3467) <= not a;
    layer5_outputs(3468) <= a xor b;
    layer5_outputs(3469) <= b;
    layer5_outputs(3470) <= a and b;
    layer5_outputs(3471) <= '1';
    layer5_outputs(3472) <= b;
    layer5_outputs(3473) <= a;
    layer5_outputs(3474) <= not b;
    layer5_outputs(3475) <= not b;
    layer5_outputs(3476) <= '1';
    layer5_outputs(3477) <= a and not b;
    layer5_outputs(3478) <= a and b;
    layer5_outputs(3479) <= not a or b;
    layer5_outputs(3480) <= a and b;
    layer5_outputs(3481) <= a xor b;
    layer5_outputs(3482) <= not b;
    layer5_outputs(3483) <= not a;
    layer5_outputs(3484) <= not b;
    layer5_outputs(3485) <= b and not a;
    layer5_outputs(3486) <= not (a and b);
    layer5_outputs(3487) <= not (a or b);
    layer5_outputs(3488) <= a;
    layer5_outputs(3489) <= not (a and b);
    layer5_outputs(3490) <= not (a or b);
    layer5_outputs(3491) <= not (a and b);
    layer5_outputs(3492) <= b;
    layer5_outputs(3493) <= b;
    layer5_outputs(3494) <= not a or b;
    layer5_outputs(3495) <= not (a or b);
    layer5_outputs(3496) <= a or b;
    layer5_outputs(3497) <= a;
    layer5_outputs(3498) <= not a;
    layer5_outputs(3499) <= not (a xor b);
    layer5_outputs(3500) <= not b;
    layer5_outputs(3501) <= not (a xor b);
    layer5_outputs(3502) <= a and b;
    layer5_outputs(3503) <= a and b;
    layer5_outputs(3504) <= a;
    layer5_outputs(3505) <= '0';
    layer5_outputs(3506) <= not (a or b);
    layer5_outputs(3507) <= '1';
    layer5_outputs(3508) <= not (a xor b);
    layer5_outputs(3509) <= b and not a;
    layer5_outputs(3510) <= not (a or b);
    layer5_outputs(3511) <= b;
    layer5_outputs(3512) <= b;
    layer5_outputs(3513) <= not (a xor b);
    layer5_outputs(3514) <= not b;
    layer5_outputs(3515) <= not (a and b);
    layer5_outputs(3516) <= b and not a;
    layer5_outputs(3517) <= not b;
    layer5_outputs(3518) <= a;
    layer5_outputs(3519) <= not a or b;
    layer5_outputs(3520) <= not (a and b);
    layer5_outputs(3521) <= not (a xor b);
    layer5_outputs(3522) <= a xor b;
    layer5_outputs(3523) <= not b;
    layer5_outputs(3524) <= b and not a;
    layer5_outputs(3525) <= b;
    layer5_outputs(3526) <= a;
    layer5_outputs(3527) <= a;
    layer5_outputs(3528) <= a;
    layer5_outputs(3529) <= a xor b;
    layer5_outputs(3530) <= a;
    layer5_outputs(3531) <= not b;
    layer5_outputs(3532) <= b;
    layer5_outputs(3533) <= not (a or b);
    layer5_outputs(3534) <= not b;
    layer5_outputs(3535) <= not a;
    layer5_outputs(3536) <= a xor b;
    layer5_outputs(3537) <= b;
    layer5_outputs(3538) <= not a;
    layer5_outputs(3539) <= not a;
    layer5_outputs(3540) <= not b;
    layer5_outputs(3541) <= not a;
    layer5_outputs(3542) <= not b;
    layer5_outputs(3543) <= not a or b;
    layer5_outputs(3544) <= b;
    layer5_outputs(3545) <= b;
    layer5_outputs(3546) <= not b or a;
    layer5_outputs(3547) <= not a;
    layer5_outputs(3548) <= a and b;
    layer5_outputs(3549) <= '1';
    layer5_outputs(3550) <= not (a xor b);
    layer5_outputs(3551) <= not b or a;
    layer5_outputs(3552) <= not b or a;
    layer5_outputs(3553) <= not b;
    layer5_outputs(3554) <= b;
    layer5_outputs(3555) <= not (a or b);
    layer5_outputs(3556) <= a and b;
    layer5_outputs(3557) <= a and b;
    layer5_outputs(3558) <= a xor b;
    layer5_outputs(3559) <= a and b;
    layer5_outputs(3560) <= a and not b;
    layer5_outputs(3561) <= b;
    layer5_outputs(3562) <= b;
    layer5_outputs(3563) <= b and not a;
    layer5_outputs(3564) <= not b;
    layer5_outputs(3565) <= b and not a;
    layer5_outputs(3566) <= '0';
    layer5_outputs(3567) <= a;
    layer5_outputs(3568) <= b;
    layer5_outputs(3569) <= a or b;
    layer5_outputs(3570) <= not a;
    layer5_outputs(3571) <= not a;
    layer5_outputs(3572) <= not (a and b);
    layer5_outputs(3573) <= not b;
    layer5_outputs(3574) <= not b or a;
    layer5_outputs(3575) <= not b or a;
    layer5_outputs(3576) <= a;
    layer5_outputs(3577) <= a and not b;
    layer5_outputs(3578) <= a or b;
    layer5_outputs(3579) <= not b;
    layer5_outputs(3580) <= not b;
    layer5_outputs(3581) <= b;
    layer5_outputs(3582) <= not (a xor b);
    layer5_outputs(3583) <= not a;
    layer5_outputs(3584) <= not a or b;
    layer5_outputs(3585) <= not a;
    layer5_outputs(3586) <= b;
    layer5_outputs(3587) <= not b;
    layer5_outputs(3588) <= b;
    layer5_outputs(3589) <= not (a and b);
    layer5_outputs(3590) <= a and b;
    layer5_outputs(3591) <= not b or a;
    layer5_outputs(3592) <= not b;
    layer5_outputs(3593) <= a or b;
    layer5_outputs(3594) <= b and not a;
    layer5_outputs(3595) <= not a;
    layer5_outputs(3596) <= not (a or b);
    layer5_outputs(3597) <= a;
    layer5_outputs(3598) <= not a;
    layer5_outputs(3599) <= b;
    layer5_outputs(3600) <= not b or a;
    layer5_outputs(3601) <= b and not a;
    layer5_outputs(3602) <= a xor b;
    layer5_outputs(3603) <= not a;
    layer5_outputs(3604) <= not (a xor b);
    layer5_outputs(3605) <= b and not a;
    layer5_outputs(3606) <= not (a or b);
    layer5_outputs(3607) <= not (a xor b);
    layer5_outputs(3608) <= '1';
    layer5_outputs(3609) <= not b;
    layer5_outputs(3610) <= a and b;
    layer5_outputs(3611) <= a or b;
    layer5_outputs(3612) <= b and not a;
    layer5_outputs(3613) <= not b;
    layer5_outputs(3614) <= b;
    layer5_outputs(3615) <= a or b;
    layer5_outputs(3616) <= not a or b;
    layer5_outputs(3617) <= a;
    layer5_outputs(3618) <= b;
    layer5_outputs(3619) <= not a;
    layer5_outputs(3620) <= not (a xor b);
    layer5_outputs(3621) <= not b or a;
    layer5_outputs(3622) <= a or b;
    layer5_outputs(3623) <= b;
    layer5_outputs(3624) <= a;
    layer5_outputs(3625) <= a xor b;
    layer5_outputs(3626) <= b;
    layer5_outputs(3627) <= not b;
    layer5_outputs(3628) <= a or b;
    layer5_outputs(3629) <= not (a or b);
    layer5_outputs(3630) <= '1';
    layer5_outputs(3631) <= a;
    layer5_outputs(3632) <= a;
    layer5_outputs(3633) <= a;
    layer5_outputs(3634) <= not b;
    layer5_outputs(3635) <= '0';
    layer5_outputs(3636) <= '1';
    layer5_outputs(3637) <= b and not a;
    layer5_outputs(3638) <= not b;
    layer5_outputs(3639) <= not b;
    layer5_outputs(3640) <= a and not b;
    layer5_outputs(3641) <= not b or a;
    layer5_outputs(3642) <= not (a or b);
    layer5_outputs(3643) <= b;
    layer5_outputs(3644) <= not (a and b);
    layer5_outputs(3645) <= not b;
    layer5_outputs(3646) <= not (a xor b);
    layer5_outputs(3647) <= not (a and b);
    layer5_outputs(3648) <= a;
    layer5_outputs(3649) <= b;
    layer5_outputs(3650) <= a and not b;
    layer5_outputs(3651) <= not (a xor b);
    layer5_outputs(3652) <= not (a and b);
    layer5_outputs(3653) <= not (a or b);
    layer5_outputs(3654) <= a xor b;
    layer5_outputs(3655) <= not (a and b);
    layer5_outputs(3656) <= a and b;
    layer5_outputs(3657) <= not (a or b);
    layer5_outputs(3658) <= a or b;
    layer5_outputs(3659) <= a;
    layer5_outputs(3660) <= a;
    layer5_outputs(3661) <= not b;
    layer5_outputs(3662) <= a;
    layer5_outputs(3663) <= b;
    layer5_outputs(3664) <= not a or b;
    layer5_outputs(3665) <= not a or b;
    layer5_outputs(3666) <= a xor b;
    layer5_outputs(3667) <= not a;
    layer5_outputs(3668) <= not b;
    layer5_outputs(3669) <= a;
    layer5_outputs(3670) <= b;
    layer5_outputs(3671) <= b and not a;
    layer5_outputs(3672) <= a and b;
    layer5_outputs(3673) <= a;
    layer5_outputs(3674) <= not b;
    layer5_outputs(3675) <= not (a xor b);
    layer5_outputs(3676) <= not b;
    layer5_outputs(3677) <= a;
    layer5_outputs(3678) <= not (a xor b);
    layer5_outputs(3679) <= not (a and b);
    layer5_outputs(3680) <= a or b;
    layer5_outputs(3681) <= not b or a;
    layer5_outputs(3682) <= '0';
    layer5_outputs(3683) <= a xor b;
    layer5_outputs(3684) <= a;
    layer5_outputs(3685) <= not a;
    layer5_outputs(3686) <= a;
    layer5_outputs(3687) <= b;
    layer5_outputs(3688) <= not a;
    layer5_outputs(3689) <= not (a xor b);
    layer5_outputs(3690) <= not (a and b);
    layer5_outputs(3691) <= a xor b;
    layer5_outputs(3692) <= not b;
    layer5_outputs(3693) <= not (a xor b);
    layer5_outputs(3694) <= a and not b;
    layer5_outputs(3695) <= a xor b;
    layer5_outputs(3696) <= a and not b;
    layer5_outputs(3697) <= not a;
    layer5_outputs(3698) <= a;
    layer5_outputs(3699) <= b;
    layer5_outputs(3700) <= a;
    layer5_outputs(3701) <= not b;
    layer5_outputs(3702) <= not (a and b);
    layer5_outputs(3703) <= not a;
    layer5_outputs(3704) <= a;
    layer5_outputs(3705) <= a xor b;
    layer5_outputs(3706) <= a;
    layer5_outputs(3707) <= not b;
    layer5_outputs(3708) <= b and not a;
    layer5_outputs(3709) <= not b;
    layer5_outputs(3710) <= not a;
    layer5_outputs(3711) <= not (a and b);
    layer5_outputs(3712) <= not (a or b);
    layer5_outputs(3713) <= not (a xor b);
    layer5_outputs(3714) <= not (a and b);
    layer5_outputs(3715) <= not a;
    layer5_outputs(3716) <= not b or a;
    layer5_outputs(3717) <= b and not a;
    layer5_outputs(3718) <= not b;
    layer5_outputs(3719) <= a or b;
    layer5_outputs(3720) <= not b;
    layer5_outputs(3721) <= not b;
    layer5_outputs(3722) <= a and not b;
    layer5_outputs(3723) <= a;
    layer5_outputs(3724) <= not (a xor b);
    layer5_outputs(3725) <= not a;
    layer5_outputs(3726) <= not (a and b);
    layer5_outputs(3727) <= a xor b;
    layer5_outputs(3728) <= b and not a;
    layer5_outputs(3729) <= not a;
    layer5_outputs(3730) <= a and not b;
    layer5_outputs(3731) <= a xor b;
    layer5_outputs(3732) <= not (a xor b);
    layer5_outputs(3733) <= not a;
    layer5_outputs(3734) <= not b or a;
    layer5_outputs(3735) <= not a;
    layer5_outputs(3736) <= b;
    layer5_outputs(3737) <= not (a xor b);
    layer5_outputs(3738) <= not a;
    layer5_outputs(3739) <= a or b;
    layer5_outputs(3740) <= not a;
    layer5_outputs(3741) <= a and not b;
    layer5_outputs(3742) <= not a;
    layer5_outputs(3743) <= not (a and b);
    layer5_outputs(3744) <= not (a or b);
    layer5_outputs(3745) <= a;
    layer5_outputs(3746) <= not b or a;
    layer5_outputs(3747) <= a or b;
    layer5_outputs(3748) <= a or b;
    layer5_outputs(3749) <= not a or b;
    layer5_outputs(3750) <= not a;
    layer5_outputs(3751) <= a and not b;
    layer5_outputs(3752) <= a and not b;
    layer5_outputs(3753) <= '0';
    layer5_outputs(3754) <= not b;
    layer5_outputs(3755) <= b;
    layer5_outputs(3756) <= not b;
    layer5_outputs(3757) <= a xor b;
    layer5_outputs(3758) <= a;
    layer5_outputs(3759) <= a and not b;
    layer5_outputs(3760) <= not b;
    layer5_outputs(3761) <= a;
    layer5_outputs(3762) <= not a;
    layer5_outputs(3763) <= b and not a;
    layer5_outputs(3764) <= not b;
    layer5_outputs(3765) <= not (a and b);
    layer5_outputs(3766) <= not b;
    layer5_outputs(3767) <= not b or a;
    layer5_outputs(3768) <= a or b;
    layer5_outputs(3769) <= not a;
    layer5_outputs(3770) <= a;
    layer5_outputs(3771) <= b and not a;
    layer5_outputs(3772) <= not a or b;
    layer5_outputs(3773) <= a xor b;
    layer5_outputs(3774) <= not b;
    layer5_outputs(3775) <= a;
    layer5_outputs(3776) <= not b;
    layer5_outputs(3777) <= a xor b;
    layer5_outputs(3778) <= a;
    layer5_outputs(3779) <= a and not b;
    layer5_outputs(3780) <= a;
    layer5_outputs(3781) <= not (a xor b);
    layer5_outputs(3782) <= not b;
    layer5_outputs(3783) <= a or b;
    layer5_outputs(3784) <= a xor b;
    layer5_outputs(3785) <= a;
    layer5_outputs(3786) <= b and not a;
    layer5_outputs(3787) <= not a;
    layer5_outputs(3788) <= a xor b;
    layer5_outputs(3789) <= not b or a;
    layer5_outputs(3790) <= not b or a;
    layer5_outputs(3791) <= a;
    layer5_outputs(3792) <= not b or a;
    layer5_outputs(3793) <= not a;
    layer5_outputs(3794) <= not b;
    layer5_outputs(3795) <= not (a or b);
    layer5_outputs(3796) <= not b or a;
    layer5_outputs(3797) <= not (a xor b);
    layer5_outputs(3798) <= not b;
    layer5_outputs(3799) <= not (a xor b);
    layer5_outputs(3800) <= not a;
    layer5_outputs(3801) <= a and b;
    layer5_outputs(3802) <= a and not b;
    layer5_outputs(3803) <= not b;
    layer5_outputs(3804) <= not (a or b);
    layer5_outputs(3805) <= not a;
    layer5_outputs(3806) <= b and not a;
    layer5_outputs(3807) <= not b or a;
    layer5_outputs(3808) <= not b;
    layer5_outputs(3809) <= b;
    layer5_outputs(3810) <= not b or a;
    layer5_outputs(3811) <= not (a or b);
    layer5_outputs(3812) <= not b;
    layer5_outputs(3813) <= not (a or b);
    layer5_outputs(3814) <= b;
    layer5_outputs(3815) <= a or b;
    layer5_outputs(3816) <= a;
    layer5_outputs(3817) <= not (a or b);
    layer5_outputs(3818) <= a;
    layer5_outputs(3819) <= not b or a;
    layer5_outputs(3820) <= a;
    layer5_outputs(3821) <= a xor b;
    layer5_outputs(3822) <= not a;
    layer5_outputs(3823) <= a and b;
    layer5_outputs(3824) <= not a or b;
    layer5_outputs(3825) <= not (a xor b);
    layer5_outputs(3826) <= not b;
    layer5_outputs(3827) <= not b or a;
    layer5_outputs(3828) <= b;
    layer5_outputs(3829) <= a and b;
    layer5_outputs(3830) <= a or b;
    layer5_outputs(3831) <= not a;
    layer5_outputs(3832) <= not (a and b);
    layer5_outputs(3833) <= not (a or b);
    layer5_outputs(3834) <= b;
    layer5_outputs(3835) <= '1';
    layer5_outputs(3836) <= not a or b;
    layer5_outputs(3837) <= not a or b;
    layer5_outputs(3838) <= a or b;
    layer5_outputs(3839) <= not a;
    layer5_outputs(3840) <= not (a xor b);
    layer5_outputs(3841) <= not (a or b);
    layer5_outputs(3842) <= not (a or b);
    layer5_outputs(3843) <= b and not a;
    layer5_outputs(3844) <= not (a or b);
    layer5_outputs(3845) <= b and not a;
    layer5_outputs(3846) <= b and not a;
    layer5_outputs(3847) <= a;
    layer5_outputs(3848) <= a and not b;
    layer5_outputs(3849) <= not (a and b);
    layer5_outputs(3850) <= a;
    layer5_outputs(3851) <= not (a or b);
    layer5_outputs(3852) <= not (a and b);
    layer5_outputs(3853) <= not a;
    layer5_outputs(3854) <= a and b;
    layer5_outputs(3855) <= not b;
    layer5_outputs(3856) <= not b;
    layer5_outputs(3857) <= a xor b;
    layer5_outputs(3858) <= a xor b;
    layer5_outputs(3859) <= a;
    layer5_outputs(3860) <= not a;
    layer5_outputs(3861) <= not b;
    layer5_outputs(3862) <= a and not b;
    layer5_outputs(3863) <= not a or b;
    layer5_outputs(3864) <= b and not a;
    layer5_outputs(3865) <= not b;
    layer5_outputs(3866) <= not b;
    layer5_outputs(3867) <= not (a or b);
    layer5_outputs(3868) <= not b;
    layer5_outputs(3869) <= not b or a;
    layer5_outputs(3870) <= not (a or b);
    layer5_outputs(3871) <= a and not b;
    layer5_outputs(3872) <= not a;
    layer5_outputs(3873) <= not (a xor b);
    layer5_outputs(3874) <= not b;
    layer5_outputs(3875) <= not b or a;
    layer5_outputs(3876) <= not a;
    layer5_outputs(3877) <= not a;
    layer5_outputs(3878) <= not (a xor b);
    layer5_outputs(3879) <= not b;
    layer5_outputs(3880) <= not b;
    layer5_outputs(3881) <= a;
    layer5_outputs(3882) <= a xor b;
    layer5_outputs(3883) <= a or b;
    layer5_outputs(3884) <= a and not b;
    layer5_outputs(3885) <= b;
    layer5_outputs(3886) <= not b or a;
    layer5_outputs(3887) <= not a;
    layer5_outputs(3888) <= not a;
    layer5_outputs(3889) <= '1';
    layer5_outputs(3890) <= b;
    layer5_outputs(3891) <= b and not a;
    layer5_outputs(3892) <= b;
    layer5_outputs(3893) <= a;
    layer5_outputs(3894) <= a and not b;
    layer5_outputs(3895) <= not (a xor b);
    layer5_outputs(3896) <= not (a and b);
    layer5_outputs(3897) <= not b;
    layer5_outputs(3898) <= a and not b;
    layer5_outputs(3899) <= b;
    layer5_outputs(3900) <= not a;
    layer5_outputs(3901) <= b and not a;
    layer5_outputs(3902) <= a;
    layer5_outputs(3903) <= b;
    layer5_outputs(3904) <= not (a and b);
    layer5_outputs(3905) <= a xor b;
    layer5_outputs(3906) <= '1';
    layer5_outputs(3907) <= b and not a;
    layer5_outputs(3908) <= not (a xor b);
    layer5_outputs(3909) <= not b or a;
    layer5_outputs(3910) <= not a;
    layer5_outputs(3911) <= a and b;
    layer5_outputs(3912) <= a xor b;
    layer5_outputs(3913) <= a;
    layer5_outputs(3914) <= a xor b;
    layer5_outputs(3915) <= b;
    layer5_outputs(3916) <= b;
    layer5_outputs(3917) <= a or b;
    layer5_outputs(3918) <= not a or b;
    layer5_outputs(3919) <= a and b;
    layer5_outputs(3920) <= a and b;
    layer5_outputs(3921) <= not a or b;
    layer5_outputs(3922) <= not b;
    layer5_outputs(3923) <= not a or b;
    layer5_outputs(3924) <= a xor b;
    layer5_outputs(3925) <= not (a xor b);
    layer5_outputs(3926) <= b;
    layer5_outputs(3927) <= not b;
    layer5_outputs(3928) <= b;
    layer5_outputs(3929) <= b;
    layer5_outputs(3930) <= not (a xor b);
    layer5_outputs(3931) <= not a or b;
    layer5_outputs(3932) <= a;
    layer5_outputs(3933) <= a or b;
    layer5_outputs(3934) <= a xor b;
    layer5_outputs(3935) <= not a;
    layer5_outputs(3936) <= a or b;
    layer5_outputs(3937) <= not (a and b);
    layer5_outputs(3938) <= b and not a;
    layer5_outputs(3939) <= a and b;
    layer5_outputs(3940) <= a;
    layer5_outputs(3941) <= a xor b;
    layer5_outputs(3942) <= not (a xor b);
    layer5_outputs(3943) <= a and not b;
    layer5_outputs(3944) <= not (a or b);
    layer5_outputs(3945) <= b;
    layer5_outputs(3946) <= not b;
    layer5_outputs(3947) <= a;
    layer5_outputs(3948) <= a;
    layer5_outputs(3949) <= a and b;
    layer5_outputs(3950) <= a and not b;
    layer5_outputs(3951) <= b;
    layer5_outputs(3952) <= not b;
    layer5_outputs(3953) <= not b or a;
    layer5_outputs(3954) <= not (a or b);
    layer5_outputs(3955) <= b;
    layer5_outputs(3956) <= a and b;
    layer5_outputs(3957) <= not b;
    layer5_outputs(3958) <= b;
    layer5_outputs(3959) <= not a;
    layer5_outputs(3960) <= not a;
    layer5_outputs(3961) <= not b;
    layer5_outputs(3962) <= not (a xor b);
    layer5_outputs(3963) <= a;
    layer5_outputs(3964) <= b;
    layer5_outputs(3965) <= not (a or b);
    layer5_outputs(3966) <= not (a and b);
    layer5_outputs(3967) <= a;
    layer5_outputs(3968) <= not (a xor b);
    layer5_outputs(3969) <= not b;
    layer5_outputs(3970) <= a or b;
    layer5_outputs(3971) <= not b;
    layer5_outputs(3972) <= not b;
    layer5_outputs(3973) <= a;
    layer5_outputs(3974) <= a;
    layer5_outputs(3975) <= a;
    layer5_outputs(3976) <= a;
    layer5_outputs(3977) <= a;
    layer5_outputs(3978) <= a or b;
    layer5_outputs(3979) <= b;
    layer5_outputs(3980) <= not (a or b);
    layer5_outputs(3981) <= not (a and b);
    layer5_outputs(3982) <= b;
    layer5_outputs(3983) <= not b;
    layer5_outputs(3984) <= b;
    layer5_outputs(3985) <= not a;
    layer5_outputs(3986) <= b;
    layer5_outputs(3987) <= not a or b;
    layer5_outputs(3988) <= a or b;
    layer5_outputs(3989) <= not (a and b);
    layer5_outputs(3990) <= not b;
    layer5_outputs(3991) <= a and not b;
    layer5_outputs(3992) <= a xor b;
    layer5_outputs(3993) <= a and not b;
    layer5_outputs(3994) <= not b;
    layer5_outputs(3995) <= not a;
    layer5_outputs(3996) <= a and b;
    layer5_outputs(3997) <= b;
    layer5_outputs(3998) <= a and b;
    layer5_outputs(3999) <= not (a and b);
    layer5_outputs(4000) <= not a;
    layer5_outputs(4001) <= b;
    layer5_outputs(4002) <= b and not a;
    layer5_outputs(4003) <= not b;
    layer5_outputs(4004) <= b;
    layer5_outputs(4005) <= not b;
    layer5_outputs(4006) <= not a;
    layer5_outputs(4007) <= a;
    layer5_outputs(4008) <= a;
    layer5_outputs(4009) <= not b;
    layer5_outputs(4010) <= not a or b;
    layer5_outputs(4011) <= not b or a;
    layer5_outputs(4012) <= b;
    layer5_outputs(4013) <= not b;
    layer5_outputs(4014) <= b;
    layer5_outputs(4015) <= not a or b;
    layer5_outputs(4016) <= not (a xor b);
    layer5_outputs(4017) <= a or b;
    layer5_outputs(4018) <= not (a xor b);
    layer5_outputs(4019) <= not b;
    layer5_outputs(4020) <= a xor b;
    layer5_outputs(4021) <= b;
    layer5_outputs(4022) <= a;
    layer5_outputs(4023) <= not b or a;
    layer5_outputs(4024) <= b;
    layer5_outputs(4025) <= not (a xor b);
    layer5_outputs(4026) <= b and not a;
    layer5_outputs(4027) <= a and not b;
    layer5_outputs(4028) <= a or b;
    layer5_outputs(4029) <= a;
    layer5_outputs(4030) <= not (a or b);
    layer5_outputs(4031) <= not (a xor b);
    layer5_outputs(4032) <= not a or b;
    layer5_outputs(4033) <= not (a or b);
    layer5_outputs(4034) <= b;
    layer5_outputs(4035) <= b;
    layer5_outputs(4036) <= a xor b;
    layer5_outputs(4037) <= not b;
    layer5_outputs(4038) <= not (a or b);
    layer5_outputs(4039) <= b;
    layer5_outputs(4040) <= not (a xor b);
    layer5_outputs(4041) <= a xor b;
    layer5_outputs(4042) <= a or b;
    layer5_outputs(4043) <= not b;
    layer5_outputs(4044) <= not b;
    layer5_outputs(4045) <= a or b;
    layer5_outputs(4046) <= a xor b;
    layer5_outputs(4047) <= b;
    layer5_outputs(4048) <= a or b;
    layer5_outputs(4049) <= not a;
    layer5_outputs(4050) <= a;
    layer5_outputs(4051) <= a;
    layer5_outputs(4052) <= b;
    layer5_outputs(4053) <= not a;
    layer5_outputs(4054) <= a and b;
    layer5_outputs(4055) <= not (a or b);
    layer5_outputs(4056) <= b;
    layer5_outputs(4057) <= not b;
    layer5_outputs(4058) <= a;
    layer5_outputs(4059) <= a xor b;
    layer5_outputs(4060) <= not b;
    layer5_outputs(4061) <= a;
    layer5_outputs(4062) <= not (a and b);
    layer5_outputs(4063) <= not b;
    layer5_outputs(4064) <= a and not b;
    layer5_outputs(4065) <= not (a or b);
    layer5_outputs(4066) <= b;
    layer5_outputs(4067) <= not (a or b);
    layer5_outputs(4068) <= not a or b;
    layer5_outputs(4069) <= a or b;
    layer5_outputs(4070) <= b;
    layer5_outputs(4071) <= a;
    layer5_outputs(4072) <= not (a xor b);
    layer5_outputs(4073) <= a or b;
    layer5_outputs(4074) <= not (a or b);
    layer5_outputs(4075) <= b;
    layer5_outputs(4076) <= not a or b;
    layer5_outputs(4077) <= not b;
    layer5_outputs(4078) <= b;
    layer5_outputs(4079) <= a or b;
    layer5_outputs(4080) <= a and b;
    layer5_outputs(4081) <= a xor b;
    layer5_outputs(4082) <= '0';
    layer5_outputs(4083) <= not (a or b);
    layer5_outputs(4084) <= a;
    layer5_outputs(4085) <= a and not b;
    layer5_outputs(4086) <= not a;
    layer5_outputs(4087) <= '1';
    layer5_outputs(4088) <= a;
    layer5_outputs(4089) <= not b or a;
    layer5_outputs(4090) <= not (a or b);
    layer5_outputs(4091) <= a and not b;
    layer5_outputs(4092) <= not b;
    layer5_outputs(4093) <= not (a xor b);
    layer5_outputs(4094) <= not a or b;
    layer5_outputs(4095) <= not (a and b);
    layer5_outputs(4096) <= not b;
    layer5_outputs(4097) <= not (a or b);
    layer5_outputs(4098) <= not (a xor b);
    layer5_outputs(4099) <= not (a and b);
    layer5_outputs(4100) <= a or b;
    layer5_outputs(4101) <= not a or b;
    layer5_outputs(4102) <= not (a xor b);
    layer5_outputs(4103) <= b;
    layer5_outputs(4104) <= a and not b;
    layer5_outputs(4105) <= a;
    layer5_outputs(4106) <= not b or a;
    layer5_outputs(4107) <= not b;
    layer5_outputs(4108) <= not a or b;
    layer5_outputs(4109) <= a;
    layer5_outputs(4110) <= b;
    layer5_outputs(4111) <= a or b;
    layer5_outputs(4112) <= b and not a;
    layer5_outputs(4113) <= not (a xor b);
    layer5_outputs(4114) <= a and b;
    layer5_outputs(4115) <= a;
    layer5_outputs(4116) <= a xor b;
    layer5_outputs(4117) <= a;
    layer5_outputs(4118) <= not b or a;
    layer5_outputs(4119) <= a and b;
    layer5_outputs(4120) <= '1';
    layer5_outputs(4121) <= not b or a;
    layer5_outputs(4122) <= not a;
    layer5_outputs(4123) <= a and b;
    layer5_outputs(4124) <= a;
    layer5_outputs(4125) <= not a;
    layer5_outputs(4126) <= not b or a;
    layer5_outputs(4127) <= a;
    layer5_outputs(4128) <= not a;
    layer5_outputs(4129) <= not a;
    layer5_outputs(4130) <= b and not a;
    layer5_outputs(4131) <= not (a and b);
    layer5_outputs(4132) <= a;
    layer5_outputs(4133) <= not (a or b);
    layer5_outputs(4134) <= not b;
    layer5_outputs(4135) <= a and not b;
    layer5_outputs(4136) <= not (a or b);
    layer5_outputs(4137) <= not (a xor b);
    layer5_outputs(4138) <= b;
    layer5_outputs(4139) <= b;
    layer5_outputs(4140) <= a xor b;
    layer5_outputs(4141) <= a or b;
    layer5_outputs(4142) <= b;
    layer5_outputs(4143) <= a;
    layer5_outputs(4144) <= b;
    layer5_outputs(4145) <= not b;
    layer5_outputs(4146) <= '0';
    layer5_outputs(4147) <= not b or a;
    layer5_outputs(4148) <= not (a xor b);
    layer5_outputs(4149) <= not b or a;
    layer5_outputs(4150) <= not (a xor b);
    layer5_outputs(4151) <= not (a and b);
    layer5_outputs(4152) <= not a;
    layer5_outputs(4153) <= not a;
    layer5_outputs(4154) <= not b or a;
    layer5_outputs(4155) <= a;
    layer5_outputs(4156) <= a and not b;
    layer5_outputs(4157) <= a and not b;
    layer5_outputs(4158) <= a;
    layer5_outputs(4159) <= not b;
    layer5_outputs(4160) <= not (a and b);
    layer5_outputs(4161) <= a;
    layer5_outputs(4162) <= not a;
    layer5_outputs(4163) <= not (a xor b);
    layer5_outputs(4164) <= not b or a;
    layer5_outputs(4165) <= b and not a;
    layer5_outputs(4166) <= a xor b;
    layer5_outputs(4167) <= a and b;
    layer5_outputs(4168) <= not b;
    layer5_outputs(4169) <= not b or a;
    layer5_outputs(4170) <= b and not a;
    layer5_outputs(4171) <= b;
    layer5_outputs(4172) <= not (a xor b);
    layer5_outputs(4173) <= a and not b;
    layer5_outputs(4174) <= a or b;
    layer5_outputs(4175) <= b;
    layer5_outputs(4176) <= b;
    layer5_outputs(4177) <= not b or a;
    layer5_outputs(4178) <= not a;
    layer5_outputs(4179) <= not (a xor b);
    layer5_outputs(4180) <= not (a xor b);
    layer5_outputs(4181) <= not (a and b);
    layer5_outputs(4182) <= not (a and b);
    layer5_outputs(4183) <= b and not a;
    layer5_outputs(4184) <= a xor b;
    layer5_outputs(4185) <= a or b;
    layer5_outputs(4186) <= a xor b;
    layer5_outputs(4187) <= a and b;
    layer5_outputs(4188) <= not b;
    layer5_outputs(4189) <= b;
    layer5_outputs(4190) <= not a;
    layer5_outputs(4191) <= a xor b;
    layer5_outputs(4192) <= not a or b;
    layer5_outputs(4193) <= not b or a;
    layer5_outputs(4194) <= b;
    layer5_outputs(4195) <= not a;
    layer5_outputs(4196) <= a and not b;
    layer5_outputs(4197) <= a and b;
    layer5_outputs(4198) <= not (a xor b);
    layer5_outputs(4199) <= b;
    layer5_outputs(4200) <= a;
    layer5_outputs(4201) <= '1';
    layer5_outputs(4202) <= not (a or b);
    layer5_outputs(4203) <= not a;
    layer5_outputs(4204) <= b;
    layer5_outputs(4205) <= not b;
    layer5_outputs(4206) <= not a or b;
    layer5_outputs(4207) <= not b;
    layer5_outputs(4208) <= not b;
    layer5_outputs(4209) <= not a;
    layer5_outputs(4210) <= b;
    layer5_outputs(4211) <= not (a xor b);
    layer5_outputs(4212) <= a or b;
    layer5_outputs(4213) <= b;
    layer5_outputs(4214) <= a or b;
    layer5_outputs(4215) <= a or b;
    layer5_outputs(4216) <= b;
    layer5_outputs(4217) <= b;
    layer5_outputs(4218) <= not a;
    layer5_outputs(4219) <= a;
    layer5_outputs(4220) <= '1';
    layer5_outputs(4221) <= not a;
    layer5_outputs(4222) <= not a or b;
    layer5_outputs(4223) <= not b or a;
    layer5_outputs(4224) <= not a;
    layer5_outputs(4225) <= not b;
    layer5_outputs(4226) <= a and b;
    layer5_outputs(4227) <= not b;
    layer5_outputs(4228) <= not a or b;
    layer5_outputs(4229) <= not (a xor b);
    layer5_outputs(4230) <= a xor b;
    layer5_outputs(4231) <= a xor b;
    layer5_outputs(4232) <= a xor b;
    layer5_outputs(4233) <= not a;
    layer5_outputs(4234) <= a and b;
    layer5_outputs(4235) <= b and not a;
    layer5_outputs(4236) <= b;
    layer5_outputs(4237) <= not a or b;
    layer5_outputs(4238) <= a and not b;
    layer5_outputs(4239) <= b and not a;
    layer5_outputs(4240) <= b;
    layer5_outputs(4241) <= not a;
    layer5_outputs(4242) <= a;
    layer5_outputs(4243) <= b and not a;
    layer5_outputs(4244) <= b;
    layer5_outputs(4245) <= a and not b;
    layer5_outputs(4246) <= a or b;
    layer5_outputs(4247) <= not (a xor b);
    layer5_outputs(4248) <= not b;
    layer5_outputs(4249) <= not (a xor b);
    layer5_outputs(4250) <= a and not b;
    layer5_outputs(4251) <= a;
    layer5_outputs(4252) <= a xor b;
    layer5_outputs(4253) <= not a or b;
    layer5_outputs(4254) <= a and not b;
    layer5_outputs(4255) <= not b;
    layer5_outputs(4256) <= not (a xor b);
    layer5_outputs(4257) <= not b;
    layer5_outputs(4258) <= not b;
    layer5_outputs(4259) <= b;
    layer5_outputs(4260) <= a and b;
    layer5_outputs(4261) <= not b;
    layer5_outputs(4262) <= '1';
    layer5_outputs(4263) <= not (a and b);
    layer5_outputs(4264) <= b and not a;
    layer5_outputs(4265) <= b;
    layer5_outputs(4266) <= not (a xor b);
    layer5_outputs(4267) <= not a;
    layer5_outputs(4268) <= not a;
    layer5_outputs(4269) <= a;
    layer5_outputs(4270) <= not b;
    layer5_outputs(4271) <= not b;
    layer5_outputs(4272) <= not b;
    layer5_outputs(4273) <= not (a or b);
    layer5_outputs(4274) <= not a;
    layer5_outputs(4275) <= not b or a;
    layer5_outputs(4276) <= not (a and b);
    layer5_outputs(4277) <= b and not a;
    layer5_outputs(4278) <= not a or b;
    layer5_outputs(4279) <= not b;
    layer5_outputs(4280) <= not (a xor b);
    layer5_outputs(4281) <= not b;
    layer5_outputs(4282) <= a xor b;
    layer5_outputs(4283) <= a;
    layer5_outputs(4284) <= a and not b;
    layer5_outputs(4285) <= not b;
    layer5_outputs(4286) <= not b or a;
    layer5_outputs(4287) <= a xor b;
    layer5_outputs(4288) <= b;
    layer5_outputs(4289) <= '0';
    layer5_outputs(4290) <= not (a xor b);
    layer5_outputs(4291) <= not b;
    layer5_outputs(4292) <= b;
    layer5_outputs(4293) <= not a;
    layer5_outputs(4294) <= b;
    layer5_outputs(4295) <= not a;
    layer5_outputs(4296) <= a;
    layer5_outputs(4297) <= b and not a;
    layer5_outputs(4298) <= '1';
    layer5_outputs(4299) <= b and not a;
    layer5_outputs(4300) <= a xor b;
    layer5_outputs(4301) <= a and not b;
    layer5_outputs(4302) <= not b or a;
    layer5_outputs(4303) <= a;
    layer5_outputs(4304) <= a;
    layer5_outputs(4305) <= not (a and b);
    layer5_outputs(4306) <= b;
    layer5_outputs(4307) <= a or b;
    layer5_outputs(4308) <= b;
    layer5_outputs(4309) <= not (a xor b);
    layer5_outputs(4310) <= a;
    layer5_outputs(4311) <= b and not a;
    layer5_outputs(4312) <= a and b;
    layer5_outputs(4313) <= a;
    layer5_outputs(4314) <= not (a or b);
    layer5_outputs(4315) <= a;
    layer5_outputs(4316) <= a and not b;
    layer5_outputs(4317) <= not b;
    layer5_outputs(4318) <= a;
    layer5_outputs(4319) <= not b;
    layer5_outputs(4320) <= b and not a;
    layer5_outputs(4321) <= a;
    layer5_outputs(4322) <= not b or a;
    layer5_outputs(4323) <= b and not a;
    layer5_outputs(4324) <= a xor b;
    layer5_outputs(4325) <= not b;
    layer5_outputs(4326) <= not (a or b);
    layer5_outputs(4327) <= a and not b;
    layer5_outputs(4328) <= a;
    layer5_outputs(4329) <= not b;
    layer5_outputs(4330) <= not a;
    layer5_outputs(4331) <= b and not a;
    layer5_outputs(4332) <= a;
    layer5_outputs(4333) <= not a or b;
    layer5_outputs(4334) <= not b;
    layer5_outputs(4335) <= a and b;
    layer5_outputs(4336) <= not b;
    layer5_outputs(4337) <= a;
    layer5_outputs(4338) <= a;
    layer5_outputs(4339) <= not a or b;
    layer5_outputs(4340) <= '0';
    layer5_outputs(4341) <= a;
    layer5_outputs(4342) <= a and b;
    layer5_outputs(4343) <= not a;
    layer5_outputs(4344) <= a and b;
    layer5_outputs(4345) <= b;
    layer5_outputs(4346) <= not (a and b);
    layer5_outputs(4347) <= b and not a;
    layer5_outputs(4348) <= b;
    layer5_outputs(4349) <= b;
    layer5_outputs(4350) <= not b or a;
    layer5_outputs(4351) <= a xor b;
    layer5_outputs(4352) <= not b;
    layer5_outputs(4353) <= a and b;
    layer5_outputs(4354) <= a;
    layer5_outputs(4355) <= a or b;
    layer5_outputs(4356) <= not (a and b);
    layer5_outputs(4357) <= a xor b;
    layer5_outputs(4358) <= not a;
    layer5_outputs(4359) <= a;
    layer5_outputs(4360) <= a and b;
    layer5_outputs(4361) <= not (a and b);
    layer5_outputs(4362) <= not (a or b);
    layer5_outputs(4363) <= not a or b;
    layer5_outputs(4364) <= not b or a;
    layer5_outputs(4365) <= b;
    layer5_outputs(4366) <= not (a xor b);
    layer5_outputs(4367) <= a xor b;
    layer5_outputs(4368) <= a or b;
    layer5_outputs(4369) <= not a;
    layer5_outputs(4370) <= b;
    layer5_outputs(4371) <= b and not a;
    layer5_outputs(4372) <= b;
    layer5_outputs(4373) <= b and not a;
    layer5_outputs(4374) <= not b;
    layer5_outputs(4375) <= not b or a;
    layer5_outputs(4376) <= not a;
    layer5_outputs(4377) <= a xor b;
    layer5_outputs(4378) <= not a;
    layer5_outputs(4379) <= b;
    layer5_outputs(4380) <= not b;
    layer5_outputs(4381) <= '0';
    layer5_outputs(4382) <= not b or a;
    layer5_outputs(4383) <= a and not b;
    layer5_outputs(4384) <= not a;
    layer5_outputs(4385) <= b;
    layer5_outputs(4386) <= not (a xor b);
    layer5_outputs(4387) <= a;
    layer5_outputs(4388) <= b and not a;
    layer5_outputs(4389) <= not b or a;
    layer5_outputs(4390) <= b;
    layer5_outputs(4391) <= a and not b;
    layer5_outputs(4392) <= not b;
    layer5_outputs(4393) <= not (a and b);
    layer5_outputs(4394) <= not b or a;
    layer5_outputs(4395) <= b;
    layer5_outputs(4396) <= not b;
    layer5_outputs(4397) <= b;
    layer5_outputs(4398) <= not (a xor b);
    layer5_outputs(4399) <= a and not b;
    layer5_outputs(4400) <= not (a and b);
    layer5_outputs(4401) <= not a;
    layer5_outputs(4402) <= not a;
    layer5_outputs(4403) <= a and b;
    layer5_outputs(4404) <= a;
    layer5_outputs(4405) <= not b;
    layer5_outputs(4406) <= not b or a;
    layer5_outputs(4407) <= not b or a;
    layer5_outputs(4408) <= not (a and b);
    layer5_outputs(4409) <= not a;
    layer5_outputs(4410) <= not (a xor b);
    layer5_outputs(4411) <= not a or b;
    layer5_outputs(4412) <= not a;
    layer5_outputs(4413) <= a;
    layer5_outputs(4414) <= a;
    layer5_outputs(4415) <= a xor b;
    layer5_outputs(4416) <= a;
    layer5_outputs(4417) <= not b or a;
    layer5_outputs(4418) <= not a or b;
    layer5_outputs(4419) <= not (a or b);
    layer5_outputs(4420) <= a or b;
    layer5_outputs(4421) <= not a;
    layer5_outputs(4422) <= not a or b;
    layer5_outputs(4423) <= not a;
    layer5_outputs(4424) <= b;
    layer5_outputs(4425) <= b;
    layer5_outputs(4426) <= a xor b;
    layer5_outputs(4427) <= a or b;
    layer5_outputs(4428) <= a and b;
    layer5_outputs(4429) <= not b;
    layer5_outputs(4430) <= not (a xor b);
    layer5_outputs(4431) <= a;
    layer5_outputs(4432) <= '0';
    layer5_outputs(4433) <= a;
    layer5_outputs(4434) <= not a;
    layer5_outputs(4435) <= not b or a;
    layer5_outputs(4436) <= a xor b;
    layer5_outputs(4437) <= not (a or b);
    layer5_outputs(4438) <= a xor b;
    layer5_outputs(4439) <= b;
    layer5_outputs(4440) <= a;
    layer5_outputs(4441) <= a and not b;
    layer5_outputs(4442) <= not (a and b);
    layer5_outputs(4443) <= a and not b;
    layer5_outputs(4444) <= '0';
    layer5_outputs(4445) <= not a;
    layer5_outputs(4446) <= a xor b;
    layer5_outputs(4447) <= not a or b;
    layer5_outputs(4448) <= not b;
    layer5_outputs(4449) <= a and b;
    layer5_outputs(4450) <= not (a or b);
    layer5_outputs(4451) <= not b;
    layer5_outputs(4452) <= not a;
    layer5_outputs(4453) <= not a;
    layer5_outputs(4454) <= a xor b;
    layer5_outputs(4455) <= not b or a;
    layer5_outputs(4456) <= not b;
    layer5_outputs(4457) <= not b;
    layer5_outputs(4458) <= not b;
    layer5_outputs(4459) <= b;
    layer5_outputs(4460) <= a and not b;
    layer5_outputs(4461) <= not (a and b);
    layer5_outputs(4462) <= a or b;
    layer5_outputs(4463) <= not b or a;
    layer5_outputs(4464) <= a or b;
    layer5_outputs(4465) <= not a;
    layer5_outputs(4466) <= not a;
    layer5_outputs(4467) <= a and b;
    layer5_outputs(4468) <= not (a xor b);
    layer5_outputs(4469) <= a or b;
    layer5_outputs(4470) <= b and not a;
    layer5_outputs(4471) <= not a;
    layer5_outputs(4472) <= not b;
    layer5_outputs(4473) <= not (a and b);
    layer5_outputs(4474) <= not b;
    layer5_outputs(4475) <= a xor b;
    layer5_outputs(4476) <= b and not a;
    layer5_outputs(4477) <= not b or a;
    layer5_outputs(4478) <= not b;
    layer5_outputs(4479) <= not a or b;
    layer5_outputs(4480) <= not (a or b);
    layer5_outputs(4481) <= not b;
    layer5_outputs(4482) <= b;
    layer5_outputs(4483) <= a xor b;
    layer5_outputs(4484) <= a;
    layer5_outputs(4485) <= not (a xor b);
    layer5_outputs(4486) <= not a or b;
    layer5_outputs(4487) <= b;
    layer5_outputs(4488) <= a and not b;
    layer5_outputs(4489) <= not a;
    layer5_outputs(4490) <= b and not a;
    layer5_outputs(4491) <= b;
    layer5_outputs(4492) <= not b or a;
    layer5_outputs(4493) <= b;
    layer5_outputs(4494) <= b;
    layer5_outputs(4495) <= not b;
    layer5_outputs(4496) <= not (a or b);
    layer5_outputs(4497) <= '0';
    layer5_outputs(4498) <= not a;
    layer5_outputs(4499) <= a;
    layer5_outputs(4500) <= not (a or b);
    layer5_outputs(4501) <= a or b;
    layer5_outputs(4502) <= b;
    layer5_outputs(4503) <= a and not b;
    layer5_outputs(4504) <= a;
    layer5_outputs(4505) <= not b;
    layer5_outputs(4506) <= not a;
    layer5_outputs(4507) <= not a;
    layer5_outputs(4508) <= b;
    layer5_outputs(4509) <= a;
    layer5_outputs(4510) <= not b or a;
    layer5_outputs(4511) <= not a or b;
    layer5_outputs(4512) <= b;
    layer5_outputs(4513) <= a or b;
    layer5_outputs(4514) <= a or b;
    layer5_outputs(4515) <= not (a and b);
    layer5_outputs(4516) <= b;
    layer5_outputs(4517) <= not a;
    layer5_outputs(4518) <= not (a and b);
    layer5_outputs(4519) <= not (a xor b);
    layer5_outputs(4520) <= b;
    layer5_outputs(4521) <= not b or a;
    layer5_outputs(4522) <= a;
    layer5_outputs(4523) <= not a;
    layer5_outputs(4524) <= not (a xor b);
    layer5_outputs(4525) <= a xor b;
    layer5_outputs(4526) <= a or b;
    layer5_outputs(4527) <= a xor b;
    layer5_outputs(4528) <= not (a xor b);
    layer5_outputs(4529) <= b;
    layer5_outputs(4530) <= b and not a;
    layer5_outputs(4531) <= a;
    layer5_outputs(4532) <= a and not b;
    layer5_outputs(4533) <= a;
    layer5_outputs(4534) <= not a;
    layer5_outputs(4535) <= a;
    layer5_outputs(4536) <= a or b;
    layer5_outputs(4537) <= not b;
    layer5_outputs(4538) <= a and not b;
    layer5_outputs(4539) <= a;
    layer5_outputs(4540) <= not (a xor b);
    layer5_outputs(4541) <= b;
    layer5_outputs(4542) <= not b or a;
    layer5_outputs(4543) <= a xor b;
    layer5_outputs(4544) <= b;
    layer5_outputs(4545) <= b;
    layer5_outputs(4546) <= not b;
    layer5_outputs(4547) <= a or b;
    layer5_outputs(4548) <= not b or a;
    layer5_outputs(4549) <= a and not b;
    layer5_outputs(4550) <= a;
    layer5_outputs(4551) <= a and b;
    layer5_outputs(4552) <= not b or a;
    layer5_outputs(4553) <= a;
    layer5_outputs(4554) <= not b;
    layer5_outputs(4555) <= not (a xor b);
    layer5_outputs(4556) <= not (a xor b);
    layer5_outputs(4557) <= a;
    layer5_outputs(4558) <= a xor b;
    layer5_outputs(4559) <= a or b;
    layer5_outputs(4560) <= not b;
    layer5_outputs(4561) <= b;
    layer5_outputs(4562) <= b and not a;
    layer5_outputs(4563) <= a or b;
    layer5_outputs(4564) <= not (a or b);
    layer5_outputs(4565) <= not a;
    layer5_outputs(4566) <= not (a and b);
    layer5_outputs(4567) <= not (a or b);
    layer5_outputs(4568) <= not a;
    layer5_outputs(4569) <= not a or b;
    layer5_outputs(4570) <= not (a or b);
    layer5_outputs(4571) <= a xor b;
    layer5_outputs(4572) <= not (a xor b);
    layer5_outputs(4573) <= not a;
    layer5_outputs(4574) <= not a;
    layer5_outputs(4575) <= a or b;
    layer5_outputs(4576) <= a or b;
    layer5_outputs(4577) <= a;
    layer5_outputs(4578) <= not (a xor b);
    layer5_outputs(4579) <= not (a xor b);
    layer5_outputs(4580) <= b;
    layer5_outputs(4581) <= not (a and b);
    layer5_outputs(4582) <= not a or b;
    layer5_outputs(4583) <= not a or b;
    layer5_outputs(4584) <= not (a xor b);
    layer5_outputs(4585) <= a and b;
    layer5_outputs(4586) <= b;
    layer5_outputs(4587) <= not b or a;
    layer5_outputs(4588) <= not a;
    layer5_outputs(4589) <= b and not a;
    layer5_outputs(4590) <= not b;
    layer5_outputs(4591) <= not b;
    layer5_outputs(4592) <= a and not b;
    layer5_outputs(4593) <= not b;
    layer5_outputs(4594) <= not b or a;
    layer5_outputs(4595) <= b;
    layer5_outputs(4596) <= not (a xor b);
    layer5_outputs(4597) <= not (a and b);
    layer5_outputs(4598) <= not (a xor b);
    layer5_outputs(4599) <= a xor b;
    layer5_outputs(4600) <= not (a or b);
    layer5_outputs(4601) <= not b;
    layer5_outputs(4602) <= not (a xor b);
    layer5_outputs(4603) <= not a or b;
    layer5_outputs(4604) <= not (a and b);
    layer5_outputs(4605) <= not a;
    layer5_outputs(4606) <= a or b;
    layer5_outputs(4607) <= not (a xor b);
    layer5_outputs(4608) <= not a;
    layer5_outputs(4609) <= not a;
    layer5_outputs(4610) <= b;
    layer5_outputs(4611) <= a;
    layer5_outputs(4612) <= not b;
    layer5_outputs(4613) <= not (a xor b);
    layer5_outputs(4614) <= not (a xor b);
    layer5_outputs(4615) <= not b or a;
    layer5_outputs(4616) <= a xor b;
    layer5_outputs(4617) <= a;
    layer5_outputs(4618) <= a or b;
    layer5_outputs(4619) <= not (a or b);
    layer5_outputs(4620) <= not (a and b);
    layer5_outputs(4621) <= a xor b;
    layer5_outputs(4622) <= a and b;
    layer5_outputs(4623) <= a and b;
    layer5_outputs(4624) <= a;
    layer5_outputs(4625) <= not a;
    layer5_outputs(4626) <= a and b;
    layer5_outputs(4627) <= not b or a;
    layer5_outputs(4628) <= not (a and b);
    layer5_outputs(4629) <= not (a xor b);
    layer5_outputs(4630) <= a xor b;
    layer5_outputs(4631) <= a;
    layer5_outputs(4632) <= not b or a;
    layer5_outputs(4633) <= not (a or b);
    layer5_outputs(4634) <= not a;
    layer5_outputs(4635) <= not b;
    layer5_outputs(4636) <= not a or b;
    layer5_outputs(4637) <= not a;
    layer5_outputs(4638) <= not b;
    layer5_outputs(4639) <= not (a and b);
    layer5_outputs(4640) <= not b;
    layer5_outputs(4641) <= not a or b;
    layer5_outputs(4642) <= a;
    layer5_outputs(4643) <= a and b;
    layer5_outputs(4644) <= b;
    layer5_outputs(4645) <= not a;
    layer5_outputs(4646) <= a;
    layer5_outputs(4647) <= a xor b;
    layer5_outputs(4648) <= a xor b;
    layer5_outputs(4649) <= not (a xor b);
    layer5_outputs(4650) <= not (a xor b);
    layer5_outputs(4651) <= not (a or b);
    layer5_outputs(4652) <= a or b;
    layer5_outputs(4653) <= a xor b;
    layer5_outputs(4654) <= '1';
    layer5_outputs(4655) <= not b;
    layer5_outputs(4656) <= not (a and b);
    layer5_outputs(4657) <= a;
    layer5_outputs(4658) <= a and b;
    layer5_outputs(4659) <= not a;
    layer5_outputs(4660) <= a or b;
    layer5_outputs(4661) <= not b;
    layer5_outputs(4662) <= not (a or b);
    layer5_outputs(4663) <= b and not a;
    layer5_outputs(4664) <= not (a xor b);
    layer5_outputs(4665) <= not a;
    layer5_outputs(4666) <= not a;
    layer5_outputs(4667) <= a and not b;
    layer5_outputs(4668) <= b;
    layer5_outputs(4669) <= not a;
    layer5_outputs(4670) <= a;
    layer5_outputs(4671) <= not a or b;
    layer5_outputs(4672) <= a and b;
    layer5_outputs(4673) <= b;
    layer5_outputs(4674) <= not a or b;
    layer5_outputs(4675) <= not b;
    layer5_outputs(4676) <= not (a and b);
    layer5_outputs(4677) <= b;
    layer5_outputs(4678) <= a;
    layer5_outputs(4679) <= not (a and b);
    layer5_outputs(4680) <= not b;
    layer5_outputs(4681) <= b;
    layer5_outputs(4682) <= not b;
    layer5_outputs(4683) <= not (a or b);
    layer5_outputs(4684) <= '0';
    layer5_outputs(4685) <= not b;
    layer5_outputs(4686) <= b;
    layer5_outputs(4687) <= a;
    layer5_outputs(4688) <= a and not b;
    layer5_outputs(4689) <= a and not b;
    layer5_outputs(4690) <= a and not b;
    layer5_outputs(4691) <= a;
    layer5_outputs(4692) <= not (a xor b);
    layer5_outputs(4693) <= a xor b;
    layer5_outputs(4694) <= not b;
    layer5_outputs(4695) <= not (a and b);
    layer5_outputs(4696) <= not (a xor b);
    layer5_outputs(4697) <= a xor b;
    layer5_outputs(4698) <= not (a or b);
    layer5_outputs(4699) <= b;
    layer5_outputs(4700) <= a or b;
    layer5_outputs(4701) <= not b;
    layer5_outputs(4702) <= a;
    layer5_outputs(4703) <= not b;
    layer5_outputs(4704) <= a and not b;
    layer5_outputs(4705) <= not b or a;
    layer5_outputs(4706) <= not (a xor b);
    layer5_outputs(4707) <= a and not b;
    layer5_outputs(4708) <= b;
    layer5_outputs(4709) <= not b or a;
    layer5_outputs(4710) <= b;
    layer5_outputs(4711) <= not (a and b);
    layer5_outputs(4712) <= b;
    layer5_outputs(4713) <= a;
    layer5_outputs(4714) <= b and not a;
    layer5_outputs(4715) <= b;
    layer5_outputs(4716) <= '0';
    layer5_outputs(4717) <= '1';
    layer5_outputs(4718) <= b;
    layer5_outputs(4719) <= not b or a;
    layer5_outputs(4720) <= b;
    layer5_outputs(4721) <= not b;
    layer5_outputs(4722) <= b;
    layer5_outputs(4723) <= not b or a;
    layer5_outputs(4724) <= a and not b;
    layer5_outputs(4725) <= b and not a;
    layer5_outputs(4726) <= a;
    layer5_outputs(4727) <= a and b;
    layer5_outputs(4728) <= not a;
    layer5_outputs(4729) <= not (a xor b);
    layer5_outputs(4730) <= a;
    layer5_outputs(4731) <= '0';
    layer5_outputs(4732) <= not (a and b);
    layer5_outputs(4733) <= not (a or b);
    layer5_outputs(4734) <= a;
    layer5_outputs(4735) <= not b or a;
    layer5_outputs(4736) <= not (a and b);
    layer5_outputs(4737) <= not a;
    layer5_outputs(4738) <= b;
    layer5_outputs(4739) <= not a;
    layer5_outputs(4740) <= a and not b;
    layer5_outputs(4741) <= not (a xor b);
    layer5_outputs(4742) <= a;
    layer5_outputs(4743) <= b and not a;
    layer5_outputs(4744) <= a and b;
    layer5_outputs(4745) <= not a;
    layer5_outputs(4746) <= not a or b;
    layer5_outputs(4747) <= not a or b;
    layer5_outputs(4748) <= a and b;
    layer5_outputs(4749) <= not (a or b);
    layer5_outputs(4750) <= not b;
    layer5_outputs(4751) <= b;
    layer5_outputs(4752) <= a and not b;
    layer5_outputs(4753) <= not a;
    layer5_outputs(4754) <= '1';
    layer5_outputs(4755) <= b;
    layer5_outputs(4756) <= not (a xor b);
    layer5_outputs(4757) <= not (a and b);
    layer5_outputs(4758) <= not (a xor b);
    layer5_outputs(4759) <= not a;
    layer5_outputs(4760) <= not a;
    layer5_outputs(4761) <= a and b;
    layer5_outputs(4762) <= a;
    layer5_outputs(4763) <= not b or a;
    layer5_outputs(4764) <= not (a xor b);
    layer5_outputs(4765) <= not b or a;
    layer5_outputs(4766) <= not a or b;
    layer5_outputs(4767) <= not b or a;
    layer5_outputs(4768) <= a;
    layer5_outputs(4769) <= b;
    layer5_outputs(4770) <= not (a xor b);
    layer5_outputs(4771) <= a xor b;
    layer5_outputs(4772) <= a xor b;
    layer5_outputs(4773) <= not (a and b);
    layer5_outputs(4774) <= a;
    layer5_outputs(4775) <= a;
    layer5_outputs(4776) <= not a or b;
    layer5_outputs(4777) <= '1';
    layer5_outputs(4778) <= b and not a;
    layer5_outputs(4779) <= not b;
    layer5_outputs(4780) <= a xor b;
    layer5_outputs(4781) <= not a;
    layer5_outputs(4782) <= not b;
    layer5_outputs(4783) <= not b or a;
    layer5_outputs(4784) <= not (a and b);
    layer5_outputs(4785) <= a;
    layer5_outputs(4786) <= not (a and b);
    layer5_outputs(4787) <= a and b;
    layer5_outputs(4788) <= not b;
    layer5_outputs(4789) <= not a;
    layer5_outputs(4790) <= a xor b;
    layer5_outputs(4791) <= a;
    layer5_outputs(4792) <= a;
    layer5_outputs(4793) <= not a;
    layer5_outputs(4794) <= not a;
    layer5_outputs(4795) <= a and not b;
    layer5_outputs(4796) <= a xor b;
    layer5_outputs(4797) <= b;
    layer5_outputs(4798) <= a or b;
    layer5_outputs(4799) <= not b;
    layer5_outputs(4800) <= not a or b;
    layer5_outputs(4801) <= a and not b;
    layer5_outputs(4802) <= b;
    layer5_outputs(4803) <= a;
    layer5_outputs(4804) <= not a;
    layer5_outputs(4805) <= a;
    layer5_outputs(4806) <= a;
    layer5_outputs(4807) <= not (a and b);
    layer5_outputs(4808) <= not (a and b);
    layer5_outputs(4809) <= b;
    layer5_outputs(4810) <= not (a and b);
    layer5_outputs(4811) <= not (a xor b);
    layer5_outputs(4812) <= b;
    layer5_outputs(4813) <= b;
    layer5_outputs(4814) <= b and not a;
    layer5_outputs(4815) <= not a;
    layer5_outputs(4816) <= a;
    layer5_outputs(4817) <= b;
    layer5_outputs(4818) <= not b;
    layer5_outputs(4819) <= not a;
    layer5_outputs(4820) <= not a;
    layer5_outputs(4821) <= a and b;
    layer5_outputs(4822) <= a;
    layer5_outputs(4823) <= not b or a;
    layer5_outputs(4824) <= not b;
    layer5_outputs(4825) <= a and b;
    layer5_outputs(4826) <= not (a xor b);
    layer5_outputs(4827) <= not (a and b);
    layer5_outputs(4828) <= a or b;
    layer5_outputs(4829) <= a or b;
    layer5_outputs(4830) <= not b;
    layer5_outputs(4831) <= a;
    layer5_outputs(4832) <= not (a xor b);
    layer5_outputs(4833) <= not b or a;
    layer5_outputs(4834) <= not (a and b);
    layer5_outputs(4835) <= '1';
    layer5_outputs(4836) <= b;
    layer5_outputs(4837) <= not a or b;
    layer5_outputs(4838) <= a and not b;
    layer5_outputs(4839) <= b;
    layer5_outputs(4840) <= not (a or b);
    layer5_outputs(4841) <= not (a xor b);
    layer5_outputs(4842) <= not (a xor b);
    layer5_outputs(4843) <= not (a or b);
    layer5_outputs(4844) <= not a;
    layer5_outputs(4845) <= a xor b;
    layer5_outputs(4846) <= not a;
    layer5_outputs(4847) <= a and b;
    layer5_outputs(4848) <= not b;
    layer5_outputs(4849) <= b;
    layer5_outputs(4850) <= not a or b;
    layer5_outputs(4851) <= a xor b;
    layer5_outputs(4852) <= b;
    layer5_outputs(4853) <= a;
    layer5_outputs(4854) <= a;
    layer5_outputs(4855) <= not b;
    layer5_outputs(4856) <= a;
    layer5_outputs(4857) <= a;
    layer5_outputs(4858) <= a or b;
    layer5_outputs(4859) <= b and not a;
    layer5_outputs(4860) <= b and not a;
    layer5_outputs(4861) <= not (a and b);
    layer5_outputs(4862) <= not a;
    layer5_outputs(4863) <= not (a and b);
    layer5_outputs(4864) <= b;
    layer5_outputs(4865) <= not a;
    layer5_outputs(4866) <= b;
    layer5_outputs(4867) <= a;
    layer5_outputs(4868) <= a;
    layer5_outputs(4869) <= not b;
    layer5_outputs(4870) <= not (a xor b);
    layer5_outputs(4871) <= a and b;
    layer5_outputs(4872) <= a and b;
    layer5_outputs(4873) <= not b;
    layer5_outputs(4874) <= b;
    layer5_outputs(4875) <= a and b;
    layer5_outputs(4876) <= not (a and b);
    layer5_outputs(4877) <= not (a and b);
    layer5_outputs(4878) <= b;
    layer5_outputs(4879) <= not a or b;
    layer5_outputs(4880) <= not a;
    layer5_outputs(4881) <= b;
    layer5_outputs(4882) <= not b;
    layer5_outputs(4883) <= a or b;
    layer5_outputs(4884) <= not (a and b);
    layer5_outputs(4885) <= a;
    layer5_outputs(4886) <= b;
    layer5_outputs(4887) <= a;
    layer5_outputs(4888) <= not (a xor b);
    layer5_outputs(4889) <= a;
    layer5_outputs(4890) <= b;
    layer5_outputs(4891) <= not (a and b);
    layer5_outputs(4892) <= a xor b;
    layer5_outputs(4893) <= b and not a;
    layer5_outputs(4894) <= b;
    layer5_outputs(4895) <= a;
    layer5_outputs(4896) <= a xor b;
    layer5_outputs(4897) <= not b;
    layer5_outputs(4898) <= '1';
    layer5_outputs(4899) <= not a or b;
    layer5_outputs(4900) <= not (a xor b);
    layer5_outputs(4901) <= not a or b;
    layer5_outputs(4902) <= not b or a;
    layer5_outputs(4903) <= a xor b;
    layer5_outputs(4904) <= a and b;
    layer5_outputs(4905) <= a xor b;
    layer5_outputs(4906) <= not b;
    layer5_outputs(4907) <= not a or b;
    layer5_outputs(4908) <= a;
    layer5_outputs(4909) <= not a;
    layer5_outputs(4910) <= not a;
    layer5_outputs(4911) <= not (a and b);
    layer5_outputs(4912) <= a or b;
    layer5_outputs(4913) <= b;
    layer5_outputs(4914) <= not b or a;
    layer5_outputs(4915) <= b;
    layer5_outputs(4916) <= not a;
    layer5_outputs(4917) <= not (a or b);
    layer5_outputs(4918) <= a and not b;
    layer5_outputs(4919) <= not (a and b);
    layer5_outputs(4920) <= b;
    layer5_outputs(4921) <= not (a or b);
    layer5_outputs(4922) <= b and not a;
    layer5_outputs(4923) <= not a;
    layer5_outputs(4924) <= not (a and b);
    layer5_outputs(4925) <= b and not a;
    layer5_outputs(4926) <= a and b;
    layer5_outputs(4927) <= a and b;
    layer5_outputs(4928) <= a or b;
    layer5_outputs(4929) <= not a;
    layer5_outputs(4930) <= not b;
    layer5_outputs(4931) <= a;
    layer5_outputs(4932) <= not b;
    layer5_outputs(4933) <= not b;
    layer5_outputs(4934) <= a and b;
    layer5_outputs(4935) <= not b;
    layer5_outputs(4936) <= a;
    layer5_outputs(4937) <= a xor b;
    layer5_outputs(4938) <= not (a and b);
    layer5_outputs(4939) <= b and not a;
    layer5_outputs(4940) <= not a;
    layer5_outputs(4941) <= not b;
    layer5_outputs(4942) <= not b;
    layer5_outputs(4943) <= a xor b;
    layer5_outputs(4944) <= not b or a;
    layer5_outputs(4945) <= not a or b;
    layer5_outputs(4946) <= '0';
    layer5_outputs(4947) <= '1';
    layer5_outputs(4948) <= a xor b;
    layer5_outputs(4949) <= not (a xor b);
    layer5_outputs(4950) <= b;
    layer5_outputs(4951) <= a or b;
    layer5_outputs(4952) <= not b;
    layer5_outputs(4953) <= not b;
    layer5_outputs(4954) <= b;
    layer5_outputs(4955) <= not a or b;
    layer5_outputs(4956) <= '1';
    layer5_outputs(4957) <= not a or b;
    layer5_outputs(4958) <= not b;
    layer5_outputs(4959) <= a or b;
    layer5_outputs(4960) <= not a;
    layer5_outputs(4961) <= a or b;
    layer5_outputs(4962) <= not b or a;
    layer5_outputs(4963) <= not (a xor b);
    layer5_outputs(4964) <= a and b;
    layer5_outputs(4965) <= b;
    layer5_outputs(4966) <= a and not b;
    layer5_outputs(4967) <= not b or a;
    layer5_outputs(4968) <= not b;
    layer5_outputs(4969) <= not a;
    layer5_outputs(4970) <= a and b;
    layer5_outputs(4971) <= not (a or b);
    layer5_outputs(4972) <= b and not a;
    layer5_outputs(4973) <= b;
    layer5_outputs(4974) <= a and b;
    layer5_outputs(4975) <= not a or b;
    layer5_outputs(4976) <= a and b;
    layer5_outputs(4977) <= not (a xor b);
    layer5_outputs(4978) <= a;
    layer5_outputs(4979) <= a xor b;
    layer5_outputs(4980) <= a;
    layer5_outputs(4981) <= not (a or b);
    layer5_outputs(4982) <= not (a xor b);
    layer5_outputs(4983) <= not b;
    layer5_outputs(4984) <= not (a or b);
    layer5_outputs(4985) <= not a;
    layer5_outputs(4986) <= a and b;
    layer5_outputs(4987) <= b;
    layer5_outputs(4988) <= a;
    layer5_outputs(4989) <= a and b;
    layer5_outputs(4990) <= b;
    layer5_outputs(4991) <= b and not a;
    layer5_outputs(4992) <= not (a and b);
    layer5_outputs(4993) <= not b;
    layer5_outputs(4994) <= a;
    layer5_outputs(4995) <= a xor b;
    layer5_outputs(4996) <= a;
    layer5_outputs(4997) <= not a;
    layer5_outputs(4998) <= b and not a;
    layer5_outputs(4999) <= a;
    layer5_outputs(5000) <= not (a or b);
    layer5_outputs(5001) <= a and not b;
    layer5_outputs(5002) <= a or b;
    layer5_outputs(5003) <= a xor b;
    layer5_outputs(5004) <= not (a and b);
    layer5_outputs(5005) <= not b;
    layer5_outputs(5006) <= a xor b;
    layer5_outputs(5007) <= not a;
    layer5_outputs(5008) <= not (a xor b);
    layer5_outputs(5009) <= not b or a;
    layer5_outputs(5010) <= a and b;
    layer5_outputs(5011) <= not (a xor b);
    layer5_outputs(5012) <= a;
    layer5_outputs(5013) <= not a;
    layer5_outputs(5014) <= not (a or b);
    layer5_outputs(5015) <= not a;
    layer5_outputs(5016) <= not b;
    layer5_outputs(5017) <= a or b;
    layer5_outputs(5018) <= a;
    layer5_outputs(5019) <= not (a xor b);
    layer5_outputs(5020) <= a and b;
    layer5_outputs(5021) <= not (a and b);
    layer5_outputs(5022) <= b and not a;
    layer5_outputs(5023) <= a xor b;
    layer5_outputs(5024) <= a;
    layer5_outputs(5025) <= not a or b;
    layer5_outputs(5026) <= not b;
    layer5_outputs(5027) <= '0';
    layer5_outputs(5028) <= b;
    layer5_outputs(5029) <= a;
    layer5_outputs(5030) <= a or b;
    layer5_outputs(5031) <= not b;
    layer5_outputs(5032) <= not a;
    layer5_outputs(5033) <= a;
    layer5_outputs(5034) <= '0';
    layer5_outputs(5035) <= not a;
    layer5_outputs(5036) <= a;
    layer5_outputs(5037) <= a;
    layer5_outputs(5038) <= not b;
    layer5_outputs(5039) <= not b;
    layer5_outputs(5040) <= not b;
    layer5_outputs(5041) <= not b;
    layer5_outputs(5042) <= a and b;
    layer5_outputs(5043) <= not (a and b);
    layer5_outputs(5044) <= b;
    layer5_outputs(5045) <= not (a xor b);
    layer5_outputs(5046) <= b and not a;
    layer5_outputs(5047) <= not a;
    layer5_outputs(5048) <= a;
    layer5_outputs(5049) <= not (a xor b);
    layer5_outputs(5050) <= not a;
    layer5_outputs(5051) <= a;
    layer5_outputs(5052) <= b and not a;
    layer5_outputs(5053) <= not b;
    layer5_outputs(5054) <= b;
    layer5_outputs(5055) <= not b;
    layer5_outputs(5056) <= not (a or b);
    layer5_outputs(5057) <= a;
    layer5_outputs(5058) <= not a or b;
    layer5_outputs(5059) <= a or b;
    layer5_outputs(5060) <= b;
    layer5_outputs(5061) <= a;
    layer5_outputs(5062) <= a or b;
    layer5_outputs(5063) <= b;
    layer5_outputs(5064) <= b;
    layer5_outputs(5065) <= a and not b;
    layer5_outputs(5066) <= not a;
    layer5_outputs(5067) <= b;
    layer5_outputs(5068) <= not (a and b);
    layer5_outputs(5069) <= not (a or b);
    layer5_outputs(5070) <= not a;
    layer5_outputs(5071) <= not b;
    layer5_outputs(5072) <= not b or a;
    layer5_outputs(5073) <= a and not b;
    layer5_outputs(5074) <= a and b;
    layer5_outputs(5075) <= not (a and b);
    layer5_outputs(5076) <= b;
    layer5_outputs(5077) <= not a;
    layer5_outputs(5078) <= a;
    layer5_outputs(5079) <= not a;
    layer5_outputs(5080) <= not a;
    layer5_outputs(5081) <= b;
    layer5_outputs(5082) <= not a;
    layer5_outputs(5083) <= not b;
    layer5_outputs(5084) <= a and not b;
    layer5_outputs(5085) <= a and b;
    layer5_outputs(5086) <= not b or a;
    layer5_outputs(5087) <= a xor b;
    layer5_outputs(5088) <= not b;
    layer5_outputs(5089) <= a xor b;
    layer5_outputs(5090) <= not a;
    layer5_outputs(5091) <= not a;
    layer5_outputs(5092) <= a and not b;
    layer5_outputs(5093) <= not (a or b);
    layer5_outputs(5094) <= a;
    layer5_outputs(5095) <= a xor b;
    layer5_outputs(5096) <= a or b;
    layer5_outputs(5097) <= not a;
    layer5_outputs(5098) <= b and not a;
    layer5_outputs(5099) <= not (a xor b);
    layer5_outputs(5100) <= b;
    layer5_outputs(5101) <= not b;
    layer5_outputs(5102) <= a or b;
    layer5_outputs(5103) <= a xor b;
    layer5_outputs(5104) <= b and not a;
    layer5_outputs(5105) <= not (a xor b);
    layer5_outputs(5106) <= not a;
    layer5_outputs(5107) <= not b;
    layer5_outputs(5108) <= not (a xor b);
    layer5_outputs(5109) <= not (a or b);
    layer5_outputs(5110) <= not (a xor b);
    layer5_outputs(5111) <= a or b;
    layer5_outputs(5112) <= a xor b;
    layer5_outputs(5113) <= not (a xor b);
    layer5_outputs(5114) <= a;
    layer5_outputs(5115) <= not b or a;
    layer5_outputs(5116) <= b;
    layer5_outputs(5117) <= not a or b;
    layer5_outputs(5118) <= a and b;
    layer5_outputs(5119) <= a and not b;
    layer5_outputs(5120) <= a and b;
    layer5_outputs(5121) <= not a;
    layer5_outputs(5122) <= b and not a;
    layer5_outputs(5123) <= not (a and b);
    layer5_outputs(5124) <= not b or a;
    layer5_outputs(5125) <= not a;
    layer5_outputs(5126) <= a or b;
    layer5_outputs(5127) <= not a;
    layer5_outputs(5128) <= not a;
    layer5_outputs(5129) <= a and not b;
    layer5_outputs(5130) <= not (a xor b);
    layer5_outputs(5131) <= not (a xor b);
    layer5_outputs(5132) <= a;
    layer5_outputs(5133) <= not a or b;
    layer5_outputs(5134) <= not (a xor b);
    layer5_outputs(5135) <= not b;
    layer5_outputs(5136) <= not b;
    layer5_outputs(5137) <= not b;
    layer5_outputs(5138) <= a and b;
    layer5_outputs(5139) <= not a;
    layer5_outputs(5140) <= b;
    layer5_outputs(5141) <= a;
    layer5_outputs(5142) <= a and b;
    layer5_outputs(5143) <= b and not a;
    layer5_outputs(5144) <= b and not a;
    layer5_outputs(5145) <= a and not b;
    layer5_outputs(5146) <= not (a or b);
    layer5_outputs(5147) <= not b;
    layer5_outputs(5148) <= not (a or b);
    layer5_outputs(5149) <= b;
    layer5_outputs(5150) <= a;
    layer5_outputs(5151) <= b and not a;
    layer5_outputs(5152) <= not (a or b);
    layer5_outputs(5153) <= a and not b;
    layer5_outputs(5154) <= b;
    layer5_outputs(5155) <= b and not a;
    layer5_outputs(5156) <= a xor b;
    layer5_outputs(5157) <= '1';
    layer5_outputs(5158) <= not (a or b);
    layer5_outputs(5159) <= a;
    layer5_outputs(5160) <= not b;
    layer5_outputs(5161) <= not (a or b);
    layer5_outputs(5162) <= not (a and b);
    layer5_outputs(5163) <= not b;
    layer5_outputs(5164) <= not b or a;
    layer5_outputs(5165) <= not b or a;
    layer5_outputs(5166) <= a and b;
    layer5_outputs(5167) <= not a;
    layer5_outputs(5168) <= b and not a;
    layer5_outputs(5169) <= not a or b;
    layer5_outputs(5170) <= a and not b;
    layer5_outputs(5171) <= not a or b;
    layer5_outputs(5172) <= a xor b;
    layer5_outputs(5173) <= not b;
    layer5_outputs(5174) <= a or b;
    layer5_outputs(5175) <= not b or a;
    layer5_outputs(5176) <= not b or a;
    layer5_outputs(5177) <= not a or b;
    layer5_outputs(5178) <= a;
    layer5_outputs(5179) <= not (a xor b);
    layer5_outputs(5180) <= b and not a;
    layer5_outputs(5181) <= not a;
    layer5_outputs(5182) <= a xor b;
    layer5_outputs(5183) <= a or b;
    layer5_outputs(5184) <= not (a or b);
    layer5_outputs(5185) <= a;
    layer5_outputs(5186) <= not b or a;
    layer5_outputs(5187) <= not b or a;
    layer5_outputs(5188) <= not (a xor b);
    layer5_outputs(5189) <= a;
    layer5_outputs(5190) <= not a or b;
    layer5_outputs(5191) <= a;
    layer5_outputs(5192) <= a xor b;
    layer5_outputs(5193) <= a xor b;
    layer5_outputs(5194) <= b;
    layer5_outputs(5195) <= not a or b;
    layer5_outputs(5196) <= not (a xor b);
    layer5_outputs(5197) <= not a;
    layer5_outputs(5198) <= a xor b;
    layer5_outputs(5199) <= a or b;
    layer5_outputs(5200) <= not (a or b);
    layer5_outputs(5201) <= a;
    layer5_outputs(5202) <= not b or a;
    layer5_outputs(5203) <= '0';
    layer5_outputs(5204) <= not a;
    layer5_outputs(5205) <= a and not b;
    layer5_outputs(5206) <= not (a xor b);
    layer5_outputs(5207) <= not (a and b);
    layer5_outputs(5208) <= not a or b;
    layer5_outputs(5209) <= not (a xor b);
    layer5_outputs(5210) <= not (a xor b);
    layer5_outputs(5211) <= not b;
    layer5_outputs(5212) <= a;
    layer5_outputs(5213) <= a and not b;
    layer5_outputs(5214) <= not b or a;
    layer5_outputs(5215) <= b;
    layer5_outputs(5216) <= not a;
    layer5_outputs(5217) <= a;
    layer5_outputs(5218) <= b;
    layer5_outputs(5219) <= b;
    layer5_outputs(5220) <= b;
    layer5_outputs(5221) <= a or b;
    layer5_outputs(5222) <= not b;
    layer5_outputs(5223) <= b;
    layer5_outputs(5224) <= not a;
    layer5_outputs(5225) <= b and not a;
    layer5_outputs(5226) <= not a or b;
    layer5_outputs(5227) <= a;
    layer5_outputs(5228) <= not (a or b);
    layer5_outputs(5229) <= a or b;
    layer5_outputs(5230) <= not a;
    layer5_outputs(5231) <= not b or a;
    layer5_outputs(5232) <= not (a xor b);
    layer5_outputs(5233) <= a and not b;
    layer5_outputs(5234) <= a xor b;
    layer5_outputs(5235) <= not b;
    layer5_outputs(5236) <= b and not a;
    layer5_outputs(5237) <= b;
    layer5_outputs(5238) <= not b or a;
    layer5_outputs(5239) <= not a;
    layer5_outputs(5240) <= not a;
    layer5_outputs(5241) <= a xor b;
    layer5_outputs(5242) <= b and not a;
    layer5_outputs(5243) <= not (a xor b);
    layer5_outputs(5244) <= a;
    layer5_outputs(5245) <= a or b;
    layer5_outputs(5246) <= a and b;
    layer5_outputs(5247) <= not b;
    layer5_outputs(5248) <= not a;
    layer5_outputs(5249) <= not (a and b);
    layer5_outputs(5250) <= a and not b;
    layer5_outputs(5251) <= a;
    layer5_outputs(5252) <= not (a or b);
    layer5_outputs(5253) <= a or b;
    layer5_outputs(5254) <= not (a xor b);
    layer5_outputs(5255) <= not a;
    layer5_outputs(5256) <= not b or a;
    layer5_outputs(5257) <= not (a xor b);
    layer5_outputs(5258) <= not (a or b);
    layer5_outputs(5259) <= a;
    layer5_outputs(5260) <= not a;
    layer5_outputs(5261) <= not b;
    layer5_outputs(5262) <= a or b;
    layer5_outputs(5263) <= b;
    layer5_outputs(5264) <= a xor b;
    layer5_outputs(5265) <= a;
    layer5_outputs(5266) <= b;
    layer5_outputs(5267) <= not (a xor b);
    layer5_outputs(5268) <= a xor b;
    layer5_outputs(5269) <= not (a xor b);
    layer5_outputs(5270) <= not b;
    layer5_outputs(5271) <= not a or b;
    layer5_outputs(5272) <= a and b;
    layer5_outputs(5273) <= not b or a;
    layer5_outputs(5274) <= b;
    layer5_outputs(5275) <= not b;
    layer5_outputs(5276) <= a;
    layer5_outputs(5277) <= not a;
    layer5_outputs(5278) <= a;
    layer5_outputs(5279) <= '1';
    layer5_outputs(5280) <= not (a xor b);
    layer5_outputs(5281) <= '1';
    layer5_outputs(5282) <= not b;
    layer5_outputs(5283) <= not b;
    layer5_outputs(5284) <= not a;
    layer5_outputs(5285) <= not (a xor b);
    layer5_outputs(5286) <= not a;
    layer5_outputs(5287) <= '0';
    layer5_outputs(5288) <= '1';
    layer5_outputs(5289) <= a and not b;
    layer5_outputs(5290) <= not (a or b);
    layer5_outputs(5291) <= a and not b;
    layer5_outputs(5292) <= a and b;
    layer5_outputs(5293) <= a xor b;
    layer5_outputs(5294) <= b;
    layer5_outputs(5295) <= a xor b;
    layer5_outputs(5296) <= a and b;
    layer5_outputs(5297) <= b;
    layer5_outputs(5298) <= not a;
    layer5_outputs(5299) <= not b;
    layer5_outputs(5300) <= b and not a;
    layer5_outputs(5301) <= not b;
    layer5_outputs(5302) <= b and not a;
    layer5_outputs(5303) <= b;
    layer5_outputs(5304) <= b;
    layer5_outputs(5305) <= not b or a;
    layer5_outputs(5306) <= not b or a;
    layer5_outputs(5307) <= a;
    layer5_outputs(5308) <= a and not b;
    layer5_outputs(5309) <= '0';
    layer5_outputs(5310) <= a xor b;
    layer5_outputs(5311) <= a;
    layer5_outputs(5312) <= a;
    layer5_outputs(5313) <= a and not b;
    layer5_outputs(5314) <= a or b;
    layer5_outputs(5315) <= b and not a;
    layer5_outputs(5316) <= b;
    layer5_outputs(5317) <= not b;
    layer5_outputs(5318) <= not b;
    layer5_outputs(5319) <= a or b;
    layer5_outputs(5320) <= not b;
    layer5_outputs(5321) <= a;
    layer5_outputs(5322) <= a;
    layer5_outputs(5323) <= a;
    layer5_outputs(5324) <= b;
    layer5_outputs(5325) <= b;
    layer5_outputs(5326) <= not (a xor b);
    layer5_outputs(5327) <= a and b;
    layer5_outputs(5328) <= not (a or b);
    layer5_outputs(5329) <= a xor b;
    layer5_outputs(5330) <= not (a xor b);
    layer5_outputs(5331) <= a;
    layer5_outputs(5332) <= a and b;
    layer5_outputs(5333) <= a;
    layer5_outputs(5334) <= '0';
    layer5_outputs(5335) <= a;
    layer5_outputs(5336) <= a or b;
    layer5_outputs(5337) <= a xor b;
    layer5_outputs(5338) <= not (a and b);
    layer5_outputs(5339) <= not (a xor b);
    layer5_outputs(5340) <= a xor b;
    layer5_outputs(5341) <= b;
    layer5_outputs(5342) <= a or b;
    layer5_outputs(5343) <= not a or b;
    layer5_outputs(5344) <= a and not b;
    layer5_outputs(5345) <= a;
    layer5_outputs(5346) <= not (a xor b);
    layer5_outputs(5347) <= a and not b;
    layer5_outputs(5348) <= not (a xor b);
    layer5_outputs(5349) <= a and not b;
    layer5_outputs(5350) <= not a;
    layer5_outputs(5351) <= not (a and b);
    layer5_outputs(5352) <= a;
    layer5_outputs(5353) <= a;
    layer5_outputs(5354) <= not (a xor b);
    layer5_outputs(5355) <= a xor b;
    layer5_outputs(5356) <= b;
    layer5_outputs(5357) <= b and not a;
    layer5_outputs(5358) <= not a;
    layer5_outputs(5359) <= b;
    layer5_outputs(5360) <= not b or a;
    layer5_outputs(5361) <= not b;
    layer5_outputs(5362) <= a;
    layer5_outputs(5363) <= not a or b;
    layer5_outputs(5364) <= not (a xor b);
    layer5_outputs(5365) <= not b or a;
    layer5_outputs(5366) <= not b;
    layer5_outputs(5367) <= not a;
    layer5_outputs(5368) <= not a or b;
    layer5_outputs(5369) <= not a;
    layer5_outputs(5370) <= not (a and b);
    layer5_outputs(5371) <= a;
    layer5_outputs(5372) <= a;
    layer5_outputs(5373) <= a;
    layer5_outputs(5374) <= not a;
    layer5_outputs(5375) <= b and not a;
    layer5_outputs(5376) <= a and not b;
    layer5_outputs(5377) <= not b;
    layer5_outputs(5378) <= a xor b;
    layer5_outputs(5379) <= not a or b;
    layer5_outputs(5380) <= b;
    layer5_outputs(5381) <= a;
    layer5_outputs(5382) <= not a;
    layer5_outputs(5383) <= not b or a;
    layer5_outputs(5384) <= a;
    layer5_outputs(5385) <= b;
    layer5_outputs(5386) <= a and not b;
    layer5_outputs(5387) <= a xor b;
    layer5_outputs(5388) <= a;
    layer5_outputs(5389) <= a;
    layer5_outputs(5390) <= b;
    layer5_outputs(5391) <= not a;
    layer5_outputs(5392) <= a;
    layer5_outputs(5393) <= not a;
    layer5_outputs(5394) <= '1';
    layer5_outputs(5395) <= a and not b;
    layer5_outputs(5396) <= not a;
    layer5_outputs(5397) <= '0';
    layer5_outputs(5398) <= a or b;
    layer5_outputs(5399) <= not b;
    layer5_outputs(5400) <= not a;
    layer5_outputs(5401) <= not b;
    layer5_outputs(5402) <= not b;
    layer5_outputs(5403) <= b;
    layer5_outputs(5404) <= not a;
    layer5_outputs(5405) <= not (a or b);
    layer5_outputs(5406) <= '0';
    layer5_outputs(5407) <= not b;
    layer5_outputs(5408) <= not a;
    layer5_outputs(5409) <= a and b;
    layer5_outputs(5410) <= a;
    layer5_outputs(5411) <= not b;
    layer5_outputs(5412) <= not b;
    layer5_outputs(5413) <= not (a xor b);
    layer5_outputs(5414) <= not (a xor b);
    layer5_outputs(5415) <= a;
    layer5_outputs(5416) <= not b or a;
    layer5_outputs(5417) <= not (a xor b);
    layer5_outputs(5418) <= a;
    layer5_outputs(5419) <= not a;
    layer5_outputs(5420) <= not b or a;
    layer5_outputs(5421) <= a and b;
    layer5_outputs(5422) <= a xor b;
    layer5_outputs(5423) <= not b or a;
    layer5_outputs(5424) <= b;
    layer5_outputs(5425) <= not a or b;
    layer5_outputs(5426) <= '0';
    layer5_outputs(5427) <= b and not a;
    layer5_outputs(5428) <= not (a or b);
    layer5_outputs(5429) <= b and not a;
    layer5_outputs(5430) <= a and not b;
    layer5_outputs(5431) <= a;
    layer5_outputs(5432) <= a and not b;
    layer5_outputs(5433) <= a and b;
    layer5_outputs(5434) <= not (a and b);
    layer5_outputs(5435) <= a and b;
    layer5_outputs(5436) <= not a;
    layer5_outputs(5437) <= not (a xor b);
    layer5_outputs(5438) <= not a or b;
    layer5_outputs(5439) <= a;
    layer5_outputs(5440) <= a;
    layer5_outputs(5441) <= a xor b;
    layer5_outputs(5442) <= a and not b;
    layer5_outputs(5443) <= a;
    layer5_outputs(5444) <= a xor b;
    layer5_outputs(5445) <= b and not a;
    layer5_outputs(5446) <= b;
    layer5_outputs(5447) <= a;
    layer5_outputs(5448) <= a and b;
    layer5_outputs(5449) <= b;
    layer5_outputs(5450) <= a;
    layer5_outputs(5451) <= not b;
    layer5_outputs(5452) <= not b;
    layer5_outputs(5453) <= not a;
    layer5_outputs(5454) <= a xor b;
    layer5_outputs(5455) <= a;
    layer5_outputs(5456) <= not a or b;
    layer5_outputs(5457) <= not (a and b);
    layer5_outputs(5458) <= not (a xor b);
    layer5_outputs(5459) <= a xor b;
    layer5_outputs(5460) <= '0';
    layer5_outputs(5461) <= b and not a;
    layer5_outputs(5462) <= not b;
    layer5_outputs(5463) <= not a;
    layer5_outputs(5464) <= not (a xor b);
    layer5_outputs(5465) <= b;
    layer5_outputs(5466) <= a;
    layer5_outputs(5467) <= a or b;
    layer5_outputs(5468) <= not a;
    layer5_outputs(5469) <= not a or b;
    layer5_outputs(5470) <= not (a and b);
    layer5_outputs(5471) <= a or b;
    layer5_outputs(5472) <= not a;
    layer5_outputs(5473) <= a;
    layer5_outputs(5474) <= not a;
    layer5_outputs(5475) <= a or b;
    layer5_outputs(5476) <= not a;
    layer5_outputs(5477) <= not a;
    layer5_outputs(5478) <= not (a or b);
    layer5_outputs(5479) <= a;
    layer5_outputs(5480) <= not (a or b);
    layer5_outputs(5481) <= a xor b;
    layer5_outputs(5482) <= b and not a;
    layer5_outputs(5483) <= b;
    layer5_outputs(5484) <= not b;
    layer5_outputs(5485) <= a xor b;
    layer5_outputs(5486) <= b;
    layer5_outputs(5487) <= a and not b;
    layer5_outputs(5488) <= not (a or b);
    layer5_outputs(5489) <= b;
    layer5_outputs(5490) <= not a;
    layer5_outputs(5491) <= not b or a;
    layer5_outputs(5492) <= not b or a;
    layer5_outputs(5493) <= not a;
    layer5_outputs(5494) <= a xor b;
    layer5_outputs(5495) <= not b;
    layer5_outputs(5496) <= a and b;
    layer5_outputs(5497) <= not (a or b);
    layer5_outputs(5498) <= a xor b;
    layer5_outputs(5499) <= not a;
    layer5_outputs(5500) <= not (a and b);
    layer5_outputs(5501) <= a xor b;
    layer5_outputs(5502) <= a xor b;
    layer5_outputs(5503) <= b;
    layer5_outputs(5504) <= not a or b;
    layer5_outputs(5505) <= not (a or b);
    layer5_outputs(5506) <= a xor b;
    layer5_outputs(5507) <= not (a or b);
    layer5_outputs(5508) <= not a;
    layer5_outputs(5509) <= b and not a;
    layer5_outputs(5510) <= b;
    layer5_outputs(5511) <= not a;
    layer5_outputs(5512) <= a and b;
    layer5_outputs(5513) <= not (a and b);
    layer5_outputs(5514) <= not a;
    layer5_outputs(5515) <= a;
    layer5_outputs(5516) <= a and b;
    layer5_outputs(5517) <= b;
    layer5_outputs(5518) <= a and not b;
    layer5_outputs(5519) <= not a or b;
    layer5_outputs(5520) <= not (a and b);
    layer5_outputs(5521) <= a or b;
    layer5_outputs(5522) <= not a;
    layer5_outputs(5523) <= a or b;
    layer5_outputs(5524) <= not a or b;
    layer5_outputs(5525) <= a;
    layer5_outputs(5526) <= not b;
    layer5_outputs(5527) <= not b;
    layer5_outputs(5528) <= not b or a;
    layer5_outputs(5529) <= not b or a;
    layer5_outputs(5530) <= a;
    layer5_outputs(5531) <= a and b;
    layer5_outputs(5532) <= b;
    layer5_outputs(5533) <= not a;
    layer5_outputs(5534) <= not (a or b);
    layer5_outputs(5535) <= a;
    layer5_outputs(5536) <= not (a and b);
    layer5_outputs(5537) <= a xor b;
    layer5_outputs(5538) <= not a;
    layer5_outputs(5539) <= b;
    layer5_outputs(5540) <= not a;
    layer5_outputs(5541) <= b;
    layer5_outputs(5542) <= not b;
    layer5_outputs(5543) <= not (a and b);
    layer5_outputs(5544) <= b;
    layer5_outputs(5545) <= not a;
    layer5_outputs(5546) <= not (a and b);
    layer5_outputs(5547) <= a;
    layer5_outputs(5548) <= a;
    layer5_outputs(5549) <= not a;
    layer5_outputs(5550) <= a;
    layer5_outputs(5551) <= a or b;
    layer5_outputs(5552) <= b;
    layer5_outputs(5553) <= b and not a;
    layer5_outputs(5554) <= a xor b;
    layer5_outputs(5555) <= a or b;
    layer5_outputs(5556) <= a xor b;
    layer5_outputs(5557) <= not a;
    layer5_outputs(5558) <= a;
    layer5_outputs(5559) <= not b;
    layer5_outputs(5560) <= a;
    layer5_outputs(5561) <= a xor b;
    layer5_outputs(5562) <= a and b;
    layer5_outputs(5563) <= not b or a;
    layer5_outputs(5564) <= a;
    layer5_outputs(5565) <= a xor b;
    layer5_outputs(5566) <= '1';
    layer5_outputs(5567) <= not a;
    layer5_outputs(5568) <= not (a xor b);
    layer5_outputs(5569) <= not a;
    layer5_outputs(5570) <= not (a or b);
    layer5_outputs(5571) <= a xor b;
    layer5_outputs(5572) <= not (a and b);
    layer5_outputs(5573) <= not b;
    layer5_outputs(5574) <= not (a and b);
    layer5_outputs(5575) <= a and not b;
    layer5_outputs(5576) <= a xor b;
    layer5_outputs(5577) <= not a;
    layer5_outputs(5578) <= not (a or b);
    layer5_outputs(5579) <= not a or b;
    layer5_outputs(5580) <= not b or a;
    layer5_outputs(5581) <= a and b;
    layer5_outputs(5582) <= not a or b;
    layer5_outputs(5583) <= a xor b;
    layer5_outputs(5584) <= not b;
    layer5_outputs(5585) <= b;
    layer5_outputs(5586) <= not b;
    layer5_outputs(5587) <= not (a xor b);
    layer5_outputs(5588) <= a or b;
    layer5_outputs(5589) <= not (a and b);
    layer5_outputs(5590) <= not a;
    layer5_outputs(5591) <= not (a xor b);
    layer5_outputs(5592) <= a or b;
    layer5_outputs(5593) <= b;
    layer5_outputs(5594) <= not b or a;
    layer5_outputs(5595) <= not a or b;
    layer5_outputs(5596) <= b and not a;
    layer5_outputs(5597) <= not b or a;
    layer5_outputs(5598) <= a;
    layer5_outputs(5599) <= not b or a;
    layer5_outputs(5600) <= not b or a;
    layer5_outputs(5601) <= not a or b;
    layer5_outputs(5602) <= not b;
    layer5_outputs(5603) <= not b;
    layer5_outputs(5604) <= not a or b;
    layer5_outputs(5605) <= b and not a;
    layer5_outputs(5606) <= a;
    layer5_outputs(5607) <= not a;
    layer5_outputs(5608) <= a and not b;
    layer5_outputs(5609) <= not a;
    layer5_outputs(5610) <= not b;
    layer5_outputs(5611) <= not a;
    layer5_outputs(5612) <= not a or b;
    layer5_outputs(5613) <= not (a and b);
    layer5_outputs(5614) <= b and not a;
    layer5_outputs(5615) <= not (a or b);
    layer5_outputs(5616) <= a;
    layer5_outputs(5617) <= a and b;
    layer5_outputs(5618) <= b;
    layer5_outputs(5619) <= not (a and b);
    layer5_outputs(5620) <= a;
    layer5_outputs(5621) <= b;
    layer5_outputs(5622) <= a and b;
    layer5_outputs(5623) <= b;
    layer5_outputs(5624) <= a and b;
    layer5_outputs(5625) <= b and not a;
    layer5_outputs(5626) <= a and b;
    layer5_outputs(5627) <= not (a xor b);
    layer5_outputs(5628) <= not a or b;
    layer5_outputs(5629) <= not b;
    layer5_outputs(5630) <= b;
    layer5_outputs(5631) <= a xor b;
    layer5_outputs(5632) <= a xor b;
    layer5_outputs(5633) <= not a;
    layer5_outputs(5634) <= not a or b;
    layer5_outputs(5635) <= b and not a;
    layer5_outputs(5636) <= b;
    layer5_outputs(5637) <= not (a xor b);
    layer5_outputs(5638) <= not b;
    layer5_outputs(5639) <= not b or a;
    layer5_outputs(5640) <= not (a and b);
    layer5_outputs(5641) <= not (a and b);
    layer5_outputs(5642) <= not b;
    layer5_outputs(5643) <= a and b;
    layer5_outputs(5644) <= not (a xor b);
    layer5_outputs(5645) <= not (a and b);
    layer5_outputs(5646) <= b;
    layer5_outputs(5647) <= a xor b;
    layer5_outputs(5648) <= not (a or b);
    layer5_outputs(5649) <= not a;
    layer5_outputs(5650) <= a;
    layer5_outputs(5651) <= a;
    layer5_outputs(5652) <= a and b;
    layer5_outputs(5653) <= not b;
    layer5_outputs(5654) <= a;
    layer5_outputs(5655) <= a xor b;
    layer5_outputs(5656) <= not a;
    layer5_outputs(5657) <= a xor b;
    layer5_outputs(5658) <= not (a or b);
    layer5_outputs(5659) <= not (a and b);
    layer5_outputs(5660) <= not b;
    layer5_outputs(5661) <= b;
    layer5_outputs(5662) <= not b;
    layer5_outputs(5663) <= a or b;
    layer5_outputs(5664) <= b and not a;
    layer5_outputs(5665) <= a and b;
    layer5_outputs(5666) <= a;
    layer5_outputs(5667) <= not a or b;
    layer5_outputs(5668) <= a;
    layer5_outputs(5669) <= not a;
    layer5_outputs(5670) <= a or b;
    layer5_outputs(5671) <= a;
    layer5_outputs(5672) <= not b;
    layer5_outputs(5673) <= a xor b;
    layer5_outputs(5674) <= not b;
    layer5_outputs(5675) <= a;
    layer5_outputs(5676) <= not a;
    layer5_outputs(5677) <= a;
    layer5_outputs(5678) <= '1';
    layer5_outputs(5679) <= not (a xor b);
    layer5_outputs(5680) <= b;
    layer5_outputs(5681) <= a;
    layer5_outputs(5682) <= a;
    layer5_outputs(5683) <= a or b;
    layer5_outputs(5684) <= not b;
    layer5_outputs(5685) <= not b;
    layer5_outputs(5686) <= a and b;
    layer5_outputs(5687) <= b;
    layer5_outputs(5688) <= a;
    layer5_outputs(5689) <= not a;
    layer5_outputs(5690) <= not a or b;
    layer5_outputs(5691) <= not b;
    layer5_outputs(5692) <= a;
    layer5_outputs(5693) <= not (a xor b);
    layer5_outputs(5694) <= not (a xor b);
    layer5_outputs(5695) <= a or b;
    layer5_outputs(5696) <= b;
    layer5_outputs(5697) <= b and not a;
    layer5_outputs(5698) <= a;
    layer5_outputs(5699) <= not a or b;
    layer5_outputs(5700) <= not (a xor b);
    layer5_outputs(5701) <= a or b;
    layer5_outputs(5702) <= b;
    layer5_outputs(5703) <= a and b;
    layer5_outputs(5704) <= not b;
    layer5_outputs(5705) <= a xor b;
    layer5_outputs(5706) <= b and not a;
    layer5_outputs(5707) <= a and not b;
    layer5_outputs(5708) <= b and not a;
    layer5_outputs(5709) <= not (a xor b);
    layer5_outputs(5710) <= a;
    layer5_outputs(5711) <= not (a xor b);
    layer5_outputs(5712) <= '0';
    layer5_outputs(5713) <= '1';
    layer5_outputs(5714) <= not a;
    layer5_outputs(5715) <= not b;
    layer5_outputs(5716) <= not (a or b);
    layer5_outputs(5717) <= a;
    layer5_outputs(5718) <= not b;
    layer5_outputs(5719) <= a xor b;
    layer5_outputs(5720) <= not (a xor b);
    layer5_outputs(5721) <= not b or a;
    layer5_outputs(5722) <= not (a xor b);
    layer5_outputs(5723) <= b;
    layer5_outputs(5724) <= a or b;
    layer5_outputs(5725) <= a xor b;
    layer5_outputs(5726) <= not (a or b);
    layer5_outputs(5727) <= a;
    layer5_outputs(5728) <= a and not b;
    layer5_outputs(5729) <= b;
    layer5_outputs(5730) <= not a;
    layer5_outputs(5731) <= not b;
    layer5_outputs(5732) <= a or b;
    layer5_outputs(5733) <= not (a and b);
    layer5_outputs(5734) <= not a;
    layer5_outputs(5735) <= b;
    layer5_outputs(5736) <= not (a and b);
    layer5_outputs(5737) <= not (a xor b);
    layer5_outputs(5738) <= b and not a;
    layer5_outputs(5739) <= not a;
    layer5_outputs(5740) <= a or b;
    layer5_outputs(5741) <= not (a or b);
    layer5_outputs(5742) <= not b or a;
    layer5_outputs(5743) <= not a;
    layer5_outputs(5744) <= a and not b;
    layer5_outputs(5745) <= not b;
    layer5_outputs(5746) <= not a;
    layer5_outputs(5747) <= not (a or b);
    layer5_outputs(5748) <= a;
    layer5_outputs(5749) <= not (a xor b);
    layer5_outputs(5750) <= not a or b;
    layer5_outputs(5751) <= b;
    layer5_outputs(5752) <= b;
    layer5_outputs(5753) <= not b;
    layer5_outputs(5754) <= a;
    layer5_outputs(5755) <= not b or a;
    layer5_outputs(5756) <= a;
    layer5_outputs(5757) <= b and not a;
    layer5_outputs(5758) <= a;
    layer5_outputs(5759) <= not a or b;
    layer5_outputs(5760) <= not (a and b);
    layer5_outputs(5761) <= a xor b;
    layer5_outputs(5762) <= a and not b;
    layer5_outputs(5763) <= a and b;
    layer5_outputs(5764) <= b and not a;
    layer5_outputs(5765) <= a and b;
    layer5_outputs(5766) <= not b;
    layer5_outputs(5767) <= not a or b;
    layer5_outputs(5768) <= not a or b;
    layer5_outputs(5769) <= not b or a;
    layer5_outputs(5770) <= b;
    layer5_outputs(5771) <= not (a xor b);
    layer5_outputs(5772) <= not a or b;
    layer5_outputs(5773) <= not a;
    layer5_outputs(5774) <= not b;
    layer5_outputs(5775) <= a and b;
    layer5_outputs(5776) <= a and b;
    layer5_outputs(5777) <= not b;
    layer5_outputs(5778) <= not b;
    layer5_outputs(5779) <= not b;
    layer5_outputs(5780) <= a;
    layer5_outputs(5781) <= b;
    layer5_outputs(5782) <= a;
    layer5_outputs(5783) <= not a;
    layer5_outputs(5784) <= a and b;
    layer5_outputs(5785) <= not a or b;
    layer5_outputs(5786) <= not a;
    layer5_outputs(5787) <= b;
    layer5_outputs(5788) <= not b or a;
    layer5_outputs(5789) <= not a;
    layer5_outputs(5790) <= a;
    layer5_outputs(5791) <= not a;
    layer5_outputs(5792) <= a;
    layer5_outputs(5793) <= not b or a;
    layer5_outputs(5794) <= b;
    layer5_outputs(5795) <= not a;
    layer5_outputs(5796) <= a xor b;
    layer5_outputs(5797) <= not b;
    layer5_outputs(5798) <= not (a xor b);
    layer5_outputs(5799) <= not a;
    layer5_outputs(5800) <= b and not a;
    layer5_outputs(5801) <= a;
    layer5_outputs(5802) <= a or b;
    layer5_outputs(5803) <= not a;
    layer5_outputs(5804) <= not b;
    layer5_outputs(5805) <= a and not b;
    layer5_outputs(5806) <= b;
    layer5_outputs(5807) <= not a;
    layer5_outputs(5808) <= a and not b;
    layer5_outputs(5809) <= not a;
    layer5_outputs(5810) <= not a or b;
    layer5_outputs(5811) <= not a;
    layer5_outputs(5812) <= '1';
    layer5_outputs(5813) <= not (a or b);
    layer5_outputs(5814) <= not a;
    layer5_outputs(5815) <= not a;
    layer5_outputs(5816) <= b and not a;
    layer5_outputs(5817) <= a and b;
    layer5_outputs(5818) <= not a;
    layer5_outputs(5819) <= a or b;
    layer5_outputs(5820) <= b;
    layer5_outputs(5821) <= a;
    layer5_outputs(5822) <= a xor b;
    layer5_outputs(5823) <= b;
    layer5_outputs(5824) <= a and b;
    layer5_outputs(5825) <= b;
    layer5_outputs(5826) <= '1';
    layer5_outputs(5827) <= not (a or b);
    layer5_outputs(5828) <= not a;
    layer5_outputs(5829) <= not (a xor b);
    layer5_outputs(5830) <= not a or b;
    layer5_outputs(5831) <= not b;
    layer5_outputs(5832) <= not a;
    layer5_outputs(5833) <= a;
    layer5_outputs(5834) <= not b;
    layer5_outputs(5835) <= '0';
    layer5_outputs(5836) <= a;
    layer5_outputs(5837) <= not b or a;
    layer5_outputs(5838) <= '1';
    layer5_outputs(5839) <= b and not a;
    layer5_outputs(5840) <= not a;
    layer5_outputs(5841) <= b and not a;
    layer5_outputs(5842) <= a and not b;
    layer5_outputs(5843) <= not b or a;
    layer5_outputs(5844) <= b;
    layer5_outputs(5845) <= b;
    layer5_outputs(5846) <= not a;
    layer5_outputs(5847) <= not a;
    layer5_outputs(5848) <= a and not b;
    layer5_outputs(5849) <= not a or b;
    layer5_outputs(5850) <= not a;
    layer5_outputs(5851) <= b;
    layer5_outputs(5852) <= not a;
    layer5_outputs(5853) <= a;
    layer5_outputs(5854) <= not b;
    layer5_outputs(5855) <= not b;
    layer5_outputs(5856) <= not a;
    layer5_outputs(5857) <= not a;
    layer5_outputs(5858) <= a or b;
    layer5_outputs(5859) <= not (a xor b);
    layer5_outputs(5860) <= not b or a;
    layer5_outputs(5861) <= b;
    layer5_outputs(5862) <= a and not b;
    layer5_outputs(5863) <= a and not b;
    layer5_outputs(5864) <= a and not b;
    layer5_outputs(5865) <= not a or b;
    layer5_outputs(5866) <= not b or a;
    layer5_outputs(5867) <= not b;
    layer5_outputs(5868) <= a and b;
    layer5_outputs(5869) <= a;
    layer5_outputs(5870) <= a and not b;
    layer5_outputs(5871) <= not b;
    layer5_outputs(5872) <= not (a xor b);
    layer5_outputs(5873) <= b;
    layer5_outputs(5874) <= b;
    layer5_outputs(5875) <= a xor b;
    layer5_outputs(5876) <= b;
    layer5_outputs(5877) <= not (a or b);
    layer5_outputs(5878) <= a and not b;
    layer5_outputs(5879) <= a;
    layer5_outputs(5880) <= b;
    layer5_outputs(5881) <= a;
    layer5_outputs(5882) <= not a or b;
    layer5_outputs(5883) <= a and b;
    layer5_outputs(5884) <= a and not b;
    layer5_outputs(5885) <= a;
    layer5_outputs(5886) <= not b;
    layer5_outputs(5887) <= b and not a;
    layer5_outputs(5888) <= a and b;
    layer5_outputs(5889) <= not b or a;
    layer5_outputs(5890) <= not a;
    layer5_outputs(5891) <= not a or b;
    layer5_outputs(5892) <= not a;
    layer5_outputs(5893) <= b and not a;
    layer5_outputs(5894) <= not b;
    layer5_outputs(5895) <= a;
    layer5_outputs(5896) <= a xor b;
    layer5_outputs(5897) <= not a or b;
    layer5_outputs(5898) <= b;
    layer5_outputs(5899) <= a and not b;
    layer5_outputs(5900) <= not b or a;
    layer5_outputs(5901) <= b;
    layer5_outputs(5902) <= not a;
    layer5_outputs(5903) <= not a or b;
    layer5_outputs(5904) <= b;
    layer5_outputs(5905) <= not (a and b);
    layer5_outputs(5906) <= not (a or b);
    layer5_outputs(5907) <= a and b;
    layer5_outputs(5908) <= not b;
    layer5_outputs(5909) <= b;
    layer5_outputs(5910) <= not a or b;
    layer5_outputs(5911) <= a;
    layer5_outputs(5912) <= not a;
    layer5_outputs(5913) <= not b;
    layer5_outputs(5914) <= b;
    layer5_outputs(5915) <= not a;
    layer5_outputs(5916) <= not (a or b);
    layer5_outputs(5917) <= not (a xor b);
    layer5_outputs(5918) <= not (a or b);
    layer5_outputs(5919) <= not b;
    layer5_outputs(5920) <= a xor b;
    layer5_outputs(5921) <= b;
    layer5_outputs(5922) <= '1';
    layer5_outputs(5923) <= not a or b;
    layer5_outputs(5924) <= b and not a;
    layer5_outputs(5925) <= b and not a;
    layer5_outputs(5926) <= not b;
    layer5_outputs(5927) <= not b or a;
    layer5_outputs(5928) <= b;
    layer5_outputs(5929) <= not a;
    layer5_outputs(5930) <= not a;
    layer5_outputs(5931) <= b and not a;
    layer5_outputs(5932) <= b;
    layer5_outputs(5933) <= not b;
    layer5_outputs(5934) <= not b;
    layer5_outputs(5935) <= not b;
    layer5_outputs(5936) <= not a;
    layer5_outputs(5937) <= a and b;
    layer5_outputs(5938) <= not b;
    layer5_outputs(5939) <= not (a or b);
    layer5_outputs(5940) <= b and not a;
    layer5_outputs(5941) <= a and b;
    layer5_outputs(5942) <= a and b;
    layer5_outputs(5943) <= not a or b;
    layer5_outputs(5944) <= not b;
    layer5_outputs(5945) <= not a or b;
    layer5_outputs(5946) <= b and not a;
    layer5_outputs(5947) <= a xor b;
    layer5_outputs(5948) <= a or b;
    layer5_outputs(5949) <= not a;
    layer5_outputs(5950) <= a and b;
    layer5_outputs(5951) <= b;
    layer5_outputs(5952) <= '1';
    layer5_outputs(5953) <= not (a xor b);
    layer5_outputs(5954) <= a or b;
    layer5_outputs(5955) <= '0';
    layer5_outputs(5956) <= not b;
    layer5_outputs(5957) <= not a or b;
    layer5_outputs(5958) <= a;
    layer5_outputs(5959) <= a xor b;
    layer5_outputs(5960) <= not (a xor b);
    layer5_outputs(5961) <= not b or a;
    layer5_outputs(5962) <= b;
    layer5_outputs(5963) <= a and not b;
    layer5_outputs(5964) <= not a;
    layer5_outputs(5965) <= not a or b;
    layer5_outputs(5966) <= not a;
    layer5_outputs(5967) <= b;
    layer5_outputs(5968) <= not (a xor b);
    layer5_outputs(5969) <= not b;
    layer5_outputs(5970) <= not b;
    layer5_outputs(5971) <= b;
    layer5_outputs(5972) <= b;
    layer5_outputs(5973) <= a and not b;
    layer5_outputs(5974) <= a xor b;
    layer5_outputs(5975) <= not a or b;
    layer5_outputs(5976) <= not b or a;
    layer5_outputs(5977) <= not (a and b);
    layer5_outputs(5978) <= not a;
    layer5_outputs(5979) <= b;
    layer5_outputs(5980) <= a xor b;
    layer5_outputs(5981) <= a and not b;
    layer5_outputs(5982) <= not (a and b);
    layer5_outputs(5983) <= not (a or b);
    layer5_outputs(5984) <= b;
    layer5_outputs(5985) <= not (a or b);
    layer5_outputs(5986) <= b;
    layer5_outputs(5987) <= b;
    layer5_outputs(5988) <= b;
    layer5_outputs(5989) <= not b;
    layer5_outputs(5990) <= not (a or b);
    layer5_outputs(5991) <= not a or b;
    layer5_outputs(5992) <= a;
    layer5_outputs(5993) <= a;
    layer5_outputs(5994) <= not b;
    layer5_outputs(5995) <= not b;
    layer5_outputs(5996) <= not b;
    layer5_outputs(5997) <= a and b;
    layer5_outputs(5998) <= not a;
    layer5_outputs(5999) <= a or b;
    layer5_outputs(6000) <= not a;
    layer5_outputs(6001) <= not (a xor b);
    layer5_outputs(6002) <= not b;
    layer5_outputs(6003) <= not b or a;
    layer5_outputs(6004) <= a;
    layer5_outputs(6005) <= a;
    layer5_outputs(6006) <= a;
    layer5_outputs(6007) <= not (a and b);
    layer5_outputs(6008) <= b;
    layer5_outputs(6009) <= not (a and b);
    layer5_outputs(6010) <= a and b;
    layer5_outputs(6011) <= not a;
    layer5_outputs(6012) <= b;
    layer5_outputs(6013) <= a;
    layer5_outputs(6014) <= b;
    layer5_outputs(6015) <= a;
    layer5_outputs(6016) <= a and b;
    layer5_outputs(6017) <= not a;
    layer5_outputs(6018) <= a xor b;
    layer5_outputs(6019) <= not a;
    layer5_outputs(6020) <= not (a and b);
    layer5_outputs(6021) <= not (a xor b);
    layer5_outputs(6022) <= a xor b;
    layer5_outputs(6023) <= b and not a;
    layer5_outputs(6024) <= a xor b;
    layer5_outputs(6025) <= b;
    layer5_outputs(6026) <= not a;
    layer5_outputs(6027) <= not b or a;
    layer5_outputs(6028) <= not (a xor b);
    layer5_outputs(6029) <= not (a or b);
    layer5_outputs(6030) <= not a or b;
    layer5_outputs(6031) <= not a;
    layer5_outputs(6032) <= not a or b;
    layer5_outputs(6033) <= not (a and b);
    layer5_outputs(6034) <= a xor b;
    layer5_outputs(6035) <= not a;
    layer5_outputs(6036) <= b;
    layer5_outputs(6037) <= '1';
    layer5_outputs(6038) <= a and not b;
    layer5_outputs(6039) <= a;
    layer5_outputs(6040) <= b;
    layer5_outputs(6041) <= not a;
    layer5_outputs(6042) <= a;
    layer5_outputs(6043) <= not a;
    layer5_outputs(6044) <= a;
    layer5_outputs(6045) <= not a or b;
    layer5_outputs(6046) <= a xor b;
    layer5_outputs(6047) <= a xor b;
    layer5_outputs(6048) <= a and b;
    layer5_outputs(6049) <= not b;
    layer5_outputs(6050) <= '1';
    layer5_outputs(6051) <= not a;
    layer5_outputs(6052) <= not a;
    layer5_outputs(6053) <= a;
    layer5_outputs(6054) <= a and b;
    layer5_outputs(6055) <= '1';
    layer5_outputs(6056) <= a;
    layer5_outputs(6057) <= a or b;
    layer5_outputs(6058) <= not b;
    layer5_outputs(6059) <= b and not a;
    layer5_outputs(6060) <= a xor b;
    layer5_outputs(6061) <= a and not b;
    layer5_outputs(6062) <= not a;
    layer5_outputs(6063) <= b;
    layer5_outputs(6064) <= b and not a;
    layer5_outputs(6065) <= b and not a;
    layer5_outputs(6066) <= not (a or b);
    layer5_outputs(6067) <= not b or a;
    layer5_outputs(6068) <= a xor b;
    layer5_outputs(6069) <= a and not b;
    layer5_outputs(6070) <= not a or b;
    layer5_outputs(6071) <= a and b;
    layer5_outputs(6072) <= a and not b;
    layer5_outputs(6073) <= a or b;
    layer5_outputs(6074) <= a and b;
    layer5_outputs(6075) <= a;
    layer5_outputs(6076) <= a xor b;
    layer5_outputs(6077) <= b and not a;
    layer5_outputs(6078) <= not b;
    layer5_outputs(6079) <= not a;
    layer5_outputs(6080) <= not a or b;
    layer5_outputs(6081) <= b;
    layer5_outputs(6082) <= b;
    layer5_outputs(6083) <= b and not a;
    layer5_outputs(6084) <= b;
    layer5_outputs(6085) <= '0';
    layer5_outputs(6086) <= b and not a;
    layer5_outputs(6087) <= not b;
    layer5_outputs(6088) <= not (a and b);
    layer5_outputs(6089) <= not (a xor b);
    layer5_outputs(6090) <= a;
    layer5_outputs(6091) <= not b;
    layer5_outputs(6092) <= not a;
    layer5_outputs(6093) <= not a;
    layer5_outputs(6094) <= a;
    layer5_outputs(6095) <= not (a xor b);
    layer5_outputs(6096) <= a;
    layer5_outputs(6097) <= a xor b;
    layer5_outputs(6098) <= not a or b;
    layer5_outputs(6099) <= a and b;
    layer5_outputs(6100) <= not a;
    layer5_outputs(6101) <= not b;
    layer5_outputs(6102) <= b and not a;
    layer5_outputs(6103) <= a;
    layer5_outputs(6104) <= not b;
    layer5_outputs(6105) <= a and b;
    layer5_outputs(6106) <= a;
    layer5_outputs(6107) <= a or b;
    layer5_outputs(6108) <= a xor b;
    layer5_outputs(6109) <= not b;
    layer5_outputs(6110) <= a or b;
    layer5_outputs(6111) <= a and not b;
    layer5_outputs(6112) <= '0';
    layer5_outputs(6113) <= not b;
    layer5_outputs(6114) <= a and not b;
    layer5_outputs(6115) <= a xor b;
    layer5_outputs(6116) <= a and not b;
    layer5_outputs(6117) <= b and not a;
    layer5_outputs(6118) <= a or b;
    layer5_outputs(6119) <= not b or a;
    layer5_outputs(6120) <= a and not b;
    layer5_outputs(6121) <= b;
    layer5_outputs(6122) <= not a;
    layer5_outputs(6123) <= a;
    layer5_outputs(6124) <= not b;
    layer5_outputs(6125) <= not a;
    layer5_outputs(6126) <= not a;
    layer5_outputs(6127) <= a xor b;
    layer5_outputs(6128) <= not (a or b);
    layer5_outputs(6129) <= not (a and b);
    layer5_outputs(6130) <= b;
    layer5_outputs(6131) <= b and not a;
    layer5_outputs(6132) <= a;
    layer5_outputs(6133) <= not (a and b);
    layer5_outputs(6134) <= a;
    layer5_outputs(6135) <= not b;
    layer5_outputs(6136) <= not a;
    layer5_outputs(6137) <= a or b;
    layer5_outputs(6138) <= b and not a;
    layer5_outputs(6139) <= not a;
    layer5_outputs(6140) <= not a;
    layer5_outputs(6141) <= a;
    layer5_outputs(6142) <= '0';
    layer5_outputs(6143) <= b and not a;
    layer5_outputs(6144) <= not a;
    layer5_outputs(6145) <= a or b;
    layer5_outputs(6146) <= a;
    layer5_outputs(6147) <= a and b;
    layer5_outputs(6148) <= not a or b;
    layer5_outputs(6149) <= b;
    layer5_outputs(6150) <= a xor b;
    layer5_outputs(6151) <= not a or b;
    layer5_outputs(6152) <= not (a or b);
    layer5_outputs(6153) <= a and b;
    layer5_outputs(6154) <= a;
    layer5_outputs(6155) <= a xor b;
    layer5_outputs(6156) <= a;
    layer5_outputs(6157) <= not a or b;
    layer5_outputs(6158) <= not b or a;
    layer5_outputs(6159) <= not a;
    layer5_outputs(6160) <= a or b;
    layer5_outputs(6161) <= b;
    layer5_outputs(6162) <= a;
    layer5_outputs(6163) <= not a;
    layer5_outputs(6164) <= b;
    layer5_outputs(6165) <= not (a xor b);
    layer5_outputs(6166) <= not b or a;
    layer5_outputs(6167) <= not b;
    layer5_outputs(6168) <= not a or b;
    layer5_outputs(6169) <= '0';
    layer5_outputs(6170) <= not b;
    layer5_outputs(6171) <= not (a and b);
    layer5_outputs(6172) <= not a;
    layer5_outputs(6173) <= not b;
    layer5_outputs(6174) <= not a or b;
    layer5_outputs(6175) <= a xor b;
    layer5_outputs(6176) <= not b or a;
    layer5_outputs(6177) <= not b;
    layer5_outputs(6178) <= b;
    layer5_outputs(6179) <= b;
    layer5_outputs(6180) <= not (a xor b);
    layer5_outputs(6181) <= b and not a;
    layer5_outputs(6182) <= a or b;
    layer5_outputs(6183) <= not a;
    layer5_outputs(6184) <= a and b;
    layer5_outputs(6185) <= a and not b;
    layer5_outputs(6186) <= a;
    layer5_outputs(6187) <= b;
    layer5_outputs(6188) <= b;
    layer5_outputs(6189) <= not a;
    layer5_outputs(6190) <= b and not a;
    layer5_outputs(6191) <= a xor b;
    layer5_outputs(6192) <= not (a and b);
    layer5_outputs(6193) <= not a or b;
    layer5_outputs(6194) <= not a;
    layer5_outputs(6195) <= a;
    layer5_outputs(6196) <= not (a xor b);
    layer5_outputs(6197) <= not (a and b);
    layer5_outputs(6198) <= not a;
    layer5_outputs(6199) <= not a;
    layer5_outputs(6200) <= not (a or b);
    layer5_outputs(6201) <= b;
    layer5_outputs(6202) <= not b;
    layer5_outputs(6203) <= not b;
    layer5_outputs(6204) <= a xor b;
    layer5_outputs(6205) <= not b;
    layer5_outputs(6206) <= not b;
    layer5_outputs(6207) <= b;
    layer5_outputs(6208) <= a and b;
    layer5_outputs(6209) <= not a;
    layer5_outputs(6210) <= not b;
    layer5_outputs(6211) <= a and b;
    layer5_outputs(6212) <= not b or a;
    layer5_outputs(6213) <= a xor b;
    layer5_outputs(6214) <= not b;
    layer5_outputs(6215) <= a xor b;
    layer5_outputs(6216) <= a xor b;
    layer5_outputs(6217) <= not a;
    layer5_outputs(6218) <= b;
    layer5_outputs(6219) <= a xor b;
    layer5_outputs(6220) <= a or b;
    layer5_outputs(6221) <= not (a and b);
    layer5_outputs(6222) <= '0';
    layer5_outputs(6223) <= a xor b;
    layer5_outputs(6224) <= not (a xor b);
    layer5_outputs(6225) <= b;
    layer5_outputs(6226) <= '0';
    layer5_outputs(6227) <= not (a xor b);
    layer5_outputs(6228) <= a or b;
    layer5_outputs(6229) <= not b or a;
    layer5_outputs(6230) <= not b;
    layer5_outputs(6231) <= a;
    layer5_outputs(6232) <= a;
    layer5_outputs(6233) <= b;
    layer5_outputs(6234) <= not b or a;
    layer5_outputs(6235) <= a and b;
    layer5_outputs(6236) <= not (a or b);
    layer5_outputs(6237) <= b;
    layer5_outputs(6238) <= not b;
    layer5_outputs(6239) <= a xor b;
    layer5_outputs(6240) <= not b;
    layer5_outputs(6241) <= not b or a;
    layer5_outputs(6242) <= b;
    layer5_outputs(6243) <= a xor b;
    layer5_outputs(6244) <= not b;
    layer5_outputs(6245) <= b and not a;
    layer5_outputs(6246) <= a and b;
    layer5_outputs(6247) <= not a or b;
    layer5_outputs(6248) <= a xor b;
    layer5_outputs(6249) <= not a;
    layer5_outputs(6250) <= not b or a;
    layer5_outputs(6251) <= not (a xor b);
    layer5_outputs(6252) <= not b;
    layer5_outputs(6253) <= a or b;
    layer5_outputs(6254) <= not b;
    layer5_outputs(6255) <= a;
    layer5_outputs(6256) <= a;
    layer5_outputs(6257) <= a and b;
    layer5_outputs(6258) <= not b or a;
    layer5_outputs(6259) <= a or b;
    layer5_outputs(6260) <= a xor b;
    layer5_outputs(6261) <= not b;
    layer5_outputs(6262) <= not a;
    layer5_outputs(6263) <= a xor b;
    layer5_outputs(6264) <= not (a or b);
    layer5_outputs(6265) <= a and not b;
    layer5_outputs(6266) <= a;
    layer5_outputs(6267) <= not (a and b);
    layer5_outputs(6268) <= b;
    layer5_outputs(6269) <= a xor b;
    layer5_outputs(6270) <= not (a xor b);
    layer5_outputs(6271) <= not b or a;
    layer5_outputs(6272) <= '1';
    layer5_outputs(6273) <= a and b;
    layer5_outputs(6274) <= a;
    layer5_outputs(6275) <= not b;
    layer5_outputs(6276) <= not (a xor b);
    layer5_outputs(6277) <= not a;
    layer5_outputs(6278) <= a and not b;
    layer5_outputs(6279) <= not b;
    layer5_outputs(6280) <= b;
    layer5_outputs(6281) <= not b;
    layer5_outputs(6282) <= a or b;
    layer5_outputs(6283) <= not (a or b);
    layer5_outputs(6284) <= a;
    layer5_outputs(6285) <= a or b;
    layer5_outputs(6286) <= not a or b;
    layer5_outputs(6287) <= not a or b;
    layer5_outputs(6288) <= not a;
    layer5_outputs(6289) <= '0';
    layer5_outputs(6290) <= a and not b;
    layer5_outputs(6291) <= not a or b;
    layer5_outputs(6292) <= a xor b;
    layer5_outputs(6293) <= not (a xor b);
    layer5_outputs(6294) <= b;
    layer5_outputs(6295) <= not b or a;
    layer5_outputs(6296) <= b and not a;
    layer5_outputs(6297) <= not (a and b);
    layer5_outputs(6298) <= not a;
    layer5_outputs(6299) <= a and b;
    layer5_outputs(6300) <= a;
    layer5_outputs(6301) <= not a;
    layer5_outputs(6302) <= not b;
    layer5_outputs(6303) <= a;
    layer5_outputs(6304) <= '0';
    layer5_outputs(6305) <= not (a xor b);
    layer5_outputs(6306) <= a and not b;
    layer5_outputs(6307) <= a;
    layer5_outputs(6308) <= not a;
    layer5_outputs(6309) <= not (a and b);
    layer5_outputs(6310) <= not a;
    layer5_outputs(6311) <= a;
    layer5_outputs(6312) <= not a or b;
    layer5_outputs(6313) <= b;
    layer5_outputs(6314) <= a or b;
    layer5_outputs(6315) <= not a;
    layer5_outputs(6316) <= not a;
    layer5_outputs(6317) <= not b;
    layer5_outputs(6318) <= not a or b;
    layer5_outputs(6319) <= not b;
    layer5_outputs(6320) <= not b;
    layer5_outputs(6321) <= not a;
    layer5_outputs(6322) <= not a;
    layer5_outputs(6323) <= a;
    layer5_outputs(6324) <= not b;
    layer5_outputs(6325) <= a or b;
    layer5_outputs(6326) <= a and not b;
    layer5_outputs(6327) <= a;
    layer5_outputs(6328) <= a xor b;
    layer5_outputs(6329) <= a;
    layer5_outputs(6330) <= not a;
    layer5_outputs(6331) <= not (a and b);
    layer5_outputs(6332) <= not a or b;
    layer5_outputs(6333) <= not (a xor b);
    layer5_outputs(6334) <= b and not a;
    layer5_outputs(6335) <= not b or a;
    layer5_outputs(6336) <= not (a xor b);
    layer5_outputs(6337) <= b;
    layer5_outputs(6338) <= a and b;
    layer5_outputs(6339) <= not (a and b);
    layer5_outputs(6340) <= not (a or b);
    layer5_outputs(6341) <= a and not b;
    layer5_outputs(6342) <= not a;
    layer5_outputs(6343) <= b;
    layer5_outputs(6344) <= not a or b;
    layer5_outputs(6345) <= not a or b;
    layer5_outputs(6346) <= not (a or b);
    layer5_outputs(6347) <= a and b;
    layer5_outputs(6348) <= a and not b;
    layer5_outputs(6349) <= not b;
    layer5_outputs(6350) <= not (a xor b);
    layer5_outputs(6351) <= not b or a;
    layer5_outputs(6352) <= a xor b;
    layer5_outputs(6353) <= a;
    layer5_outputs(6354) <= not a or b;
    layer5_outputs(6355) <= a;
    layer5_outputs(6356) <= not a;
    layer5_outputs(6357) <= a and b;
    layer5_outputs(6358) <= not (a or b);
    layer5_outputs(6359) <= a;
    layer5_outputs(6360) <= b;
    layer5_outputs(6361) <= not b or a;
    layer5_outputs(6362) <= a;
    layer5_outputs(6363) <= not a or b;
    layer5_outputs(6364) <= not a;
    layer5_outputs(6365) <= not a;
    layer5_outputs(6366) <= a or b;
    layer5_outputs(6367) <= not b;
    layer5_outputs(6368) <= not b;
    layer5_outputs(6369) <= not a;
    layer5_outputs(6370) <= not a;
    layer5_outputs(6371) <= not b;
    layer5_outputs(6372) <= '1';
    layer5_outputs(6373) <= not (a and b);
    layer5_outputs(6374) <= not a or b;
    layer5_outputs(6375) <= b;
    layer5_outputs(6376) <= not (a xor b);
    layer5_outputs(6377) <= b and not a;
    layer5_outputs(6378) <= not (a or b);
    layer5_outputs(6379) <= not (a xor b);
    layer5_outputs(6380) <= a;
    layer5_outputs(6381) <= not b;
    layer5_outputs(6382) <= a and b;
    layer5_outputs(6383) <= not (a and b);
    layer5_outputs(6384) <= not b or a;
    layer5_outputs(6385) <= not a or b;
    layer5_outputs(6386) <= a and not b;
    layer5_outputs(6387) <= not b;
    layer5_outputs(6388) <= not a or b;
    layer5_outputs(6389) <= not b or a;
    layer5_outputs(6390) <= a and b;
    layer5_outputs(6391) <= a and b;
    layer5_outputs(6392) <= not (a and b);
    layer5_outputs(6393) <= not a;
    layer5_outputs(6394) <= b;
    layer5_outputs(6395) <= not b;
    layer5_outputs(6396) <= a or b;
    layer5_outputs(6397) <= not b;
    layer5_outputs(6398) <= a;
    layer5_outputs(6399) <= not a or b;
    layer5_outputs(6400) <= not (a or b);
    layer5_outputs(6401) <= not (a and b);
    layer5_outputs(6402) <= b;
    layer5_outputs(6403) <= not b;
    layer5_outputs(6404) <= a and not b;
    layer5_outputs(6405) <= not b;
    layer5_outputs(6406) <= not (a xor b);
    layer5_outputs(6407) <= a xor b;
    layer5_outputs(6408) <= not (a or b);
    layer5_outputs(6409) <= a or b;
    layer5_outputs(6410) <= not b;
    layer5_outputs(6411) <= a and b;
    layer5_outputs(6412) <= a and not b;
    layer5_outputs(6413) <= not a;
    layer5_outputs(6414) <= a and b;
    layer5_outputs(6415) <= not b;
    layer5_outputs(6416) <= a and b;
    layer5_outputs(6417) <= not a;
    layer5_outputs(6418) <= a;
    layer5_outputs(6419) <= not b;
    layer5_outputs(6420) <= not (a xor b);
    layer5_outputs(6421) <= a;
    layer5_outputs(6422) <= a;
    layer5_outputs(6423) <= a and b;
    layer5_outputs(6424) <= b;
    layer5_outputs(6425) <= not b or a;
    layer5_outputs(6426) <= a xor b;
    layer5_outputs(6427) <= a xor b;
    layer5_outputs(6428) <= a;
    layer5_outputs(6429) <= not a or b;
    layer5_outputs(6430) <= not (a xor b);
    layer5_outputs(6431) <= b and not a;
    layer5_outputs(6432) <= b and not a;
    layer5_outputs(6433) <= a;
    layer5_outputs(6434) <= not (a or b);
    layer5_outputs(6435) <= b;
    layer5_outputs(6436) <= a and b;
    layer5_outputs(6437) <= not b;
    layer5_outputs(6438) <= b;
    layer5_outputs(6439) <= b;
    layer5_outputs(6440) <= not b;
    layer5_outputs(6441) <= not (a and b);
    layer5_outputs(6442) <= b and not a;
    layer5_outputs(6443) <= '1';
    layer5_outputs(6444) <= a;
    layer5_outputs(6445) <= a and not b;
    layer5_outputs(6446) <= not b;
    layer5_outputs(6447) <= a and not b;
    layer5_outputs(6448) <= a;
    layer5_outputs(6449) <= not (a xor b);
    layer5_outputs(6450) <= not a or b;
    layer5_outputs(6451) <= a and b;
    layer5_outputs(6452) <= b;
    layer5_outputs(6453) <= b;
    layer5_outputs(6454) <= not b or a;
    layer5_outputs(6455) <= '1';
    layer5_outputs(6456) <= a;
    layer5_outputs(6457) <= a or b;
    layer5_outputs(6458) <= not b;
    layer5_outputs(6459) <= not (a or b);
    layer5_outputs(6460) <= not (a and b);
    layer5_outputs(6461) <= a;
    layer5_outputs(6462) <= a or b;
    layer5_outputs(6463) <= not b;
    layer5_outputs(6464) <= not b;
    layer5_outputs(6465) <= not b or a;
    layer5_outputs(6466) <= b and not a;
    layer5_outputs(6467) <= not a;
    layer5_outputs(6468) <= not b or a;
    layer5_outputs(6469) <= b;
    layer5_outputs(6470) <= a xor b;
    layer5_outputs(6471) <= not (a and b);
    layer5_outputs(6472) <= not a;
    layer5_outputs(6473) <= not b;
    layer5_outputs(6474) <= not b;
    layer5_outputs(6475) <= not (a and b);
    layer5_outputs(6476) <= a;
    layer5_outputs(6477) <= not a;
    layer5_outputs(6478) <= a xor b;
    layer5_outputs(6479) <= not b;
    layer5_outputs(6480) <= not b or a;
    layer5_outputs(6481) <= a;
    layer5_outputs(6482) <= not b;
    layer5_outputs(6483) <= not b;
    layer5_outputs(6484) <= a and not b;
    layer5_outputs(6485) <= not (a xor b);
    layer5_outputs(6486) <= a;
    layer5_outputs(6487) <= a or b;
    layer5_outputs(6488) <= not a;
    layer5_outputs(6489) <= not a or b;
    layer5_outputs(6490) <= not a;
    layer5_outputs(6491) <= a;
    layer5_outputs(6492) <= not a;
    layer5_outputs(6493) <= not (a or b);
    layer5_outputs(6494) <= b;
    layer5_outputs(6495) <= not b;
    layer5_outputs(6496) <= not (a xor b);
    layer5_outputs(6497) <= b and not a;
    layer5_outputs(6498) <= a or b;
    layer5_outputs(6499) <= a;
    layer5_outputs(6500) <= a;
    layer5_outputs(6501) <= a and b;
    layer5_outputs(6502) <= not (a or b);
    layer5_outputs(6503) <= not a;
    layer5_outputs(6504) <= not (a xor b);
    layer5_outputs(6505) <= a xor b;
    layer5_outputs(6506) <= b;
    layer5_outputs(6507) <= a;
    layer5_outputs(6508) <= not (a or b);
    layer5_outputs(6509) <= not b or a;
    layer5_outputs(6510) <= not a;
    layer5_outputs(6511) <= b;
    layer5_outputs(6512) <= a;
    layer5_outputs(6513) <= not b;
    layer5_outputs(6514) <= '0';
    layer5_outputs(6515) <= not a;
    layer5_outputs(6516) <= not a or b;
    layer5_outputs(6517) <= b;
    layer5_outputs(6518) <= b;
    layer5_outputs(6519) <= a and b;
    layer5_outputs(6520) <= not a;
    layer5_outputs(6521) <= not (a or b);
    layer5_outputs(6522) <= a and b;
    layer5_outputs(6523) <= a xor b;
    layer5_outputs(6524) <= b;
    layer5_outputs(6525) <= b and not a;
    layer5_outputs(6526) <= not a or b;
    layer5_outputs(6527) <= not (a xor b);
    layer5_outputs(6528) <= a;
    layer5_outputs(6529) <= not (a xor b);
    layer5_outputs(6530) <= not b;
    layer5_outputs(6531) <= a;
    layer5_outputs(6532) <= a and not b;
    layer5_outputs(6533) <= not (a xor b);
    layer5_outputs(6534) <= a xor b;
    layer5_outputs(6535) <= not b or a;
    layer5_outputs(6536) <= b;
    layer5_outputs(6537) <= b and not a;
    layer5_outputs(6538) <= not (a xor b);
    layer5_outputs(6539) <= a;
    layer5_outputs(6540) <= a;
    layer5_outputs(6541) <= a;
    layer5_outputs(6542) <= not a;
    layer5_outputs(6543) <= a;
    layer5_outputs(6544) <= a and b;
    layer5_outputs(6545) <= a;
    layer5_outputs(6546) <= a;
    layer5_outputs(6547) <= a xor b;
    layer5_outputs(6548) <= not a;
    layer5_outputs(6549) <= not (a xor b);
    layer5_outputs(6550) <= not (a xor b);
    layer5_outputs(6551) <= not (a and b);
    layer5_outputs(6552) <= b;
    layer5_outputs(6553) <= a and not b;
    layer5_outputs(6554) <= a and b;
    layer5_outputs(6555) <= not a;
    layer5_outputs(6556) <= a;
    layer5_outputs(6557) <= not b;
    layer5_outputs(6558) <= a;
    layer5_outputs(6559) <= not b or a;
    layer5_outputs(6560) <= not a;
    layer5_outputs(6561) <= not (a or b);
    layer5_outputs(6562) <= not (a xor b);
    layer5_outputs(6563) <= b;
    layer5_outputs(6564) <= a xor b;
    layer5_outputs(6565) <= not a or b;
    layer5_outputs(6566) <= not b or a;
    layer5_outputs(6567) <= a and b;
    layer5_outputs(6568) <= b and not a;
    layer5_outputs(6569) <= not (a xor b);
    layer5_outputs(6570) <= not b or a;
    layer5_outputs(6571) <= not b or a;
    layer5_outputs(6572) <= b and not a;
    layer5_outputs(6573) <= b and not a;
    layer5_outputs(6574) <= b;
    layer5_outputs(6575) <= b and not a;
    layer5_outputs(6576) <= not b;
    layer5_outputs(6577) <= not b or a;
    layer5_outputs(6578) <= not b;
    layer5_outputs(6579) <= not b;
    layer5_outputs(6580) <= not a;
    layer5_outputs(6581) <= not a;
    layer5_outputs(6582) <= a;
    layer5_outputs(6583) <= not (a and b);
    layer5_outputs(6584) <= b and not a;
    layer5_outputs(6585) <= not (a and b);
    layer5_outputs(6586) <= not b or a;
    layer5_outputs(6587) <= not a or b;
    layer5_outputs(6588) <= not (a xor b);
    layer5_outputs(6589) <= not a or b;
    layer5_outputs(6590) <= not b or a;
    layer5_outputs(6591) <= not b;
    layer5_outputs(6592) <= not a;
    layer5_outputs(6593) <= not b or a;
    layer5_outputs(6594) <= a xor b;
    layer5_outputs(6595) <= not (a xor b);
    layer5_outputs(6596) <= a xor b;
    layer5_outputs(6597) <= not b or a;
    layer5_outputs(6598) <= a or b;
    layer5_outputs(6599) <= not b;
    layer5_outputs(6600) <= not (a or b);
    layer5_outputs(6601) <= not a;
    layer5_outputs(6602) <= b and not a;
    layer5_outputs(6603) <= '1';
    layer5_outputs(6604) <= not a;
    layer5_outputs(6605) <= b;
    layer5_outputs(6606) <= b;
    layer5_outputs(6607) <= not a or b;
    layer5_outputs(6608) <= b;
    layer5_outputs(6609) <= a or b;
    layer5_outputs(6610) <= b;
    layer5_outputs(6611) <= not (a xor b);
    layer5_outputs(6612) <= not b or a;
    layer5_outputs(6613) <= a;
    layer5_outputs(6614) <= not a;
    layer5_outputs(6615) <= a;
    layer5_outputs(6616) <= not (a or b);
    layer5_outputs(6617) <= b;
    layer5_outputs(6618) <= b;
    layer5_outputs(6619) <= b and not a;
    layer5_outputs(6620) <= not b or a;
    layer5_outputs(6621) <= '0';
    layer5_outputs(6622) <= a;
    layer5_outputs(6623) <= not a;
    layer5_outputs(6624) <= not a;
    layer5_outputs(6625) <= not b;
    layer5_outputs(6626) <= a and not b;
    layer5_outputs(6627) <= b;
    layer5_outputs(6628) <= not (a or b);
    layer5_outputs(6629) <= a;
    layer5_outputs(6630) <= not b or a;
    layer5_outputs(6631) <= b and not a;
    layer5_outputs(6632) <= a or b;
    layer5_outputs(6633) <= not (a or b);
    layer5_outputs(6634) <= not a;
    layer5_outputs(6635) <= a;
    layer5_outputs(6636) <= not a or b;
    layer5_outputs(6637) <= a and b;
    layer5_outputs(6638) <= b;
    layer5_outputs(6639) <= not b or a;
    layer5_outputs(6640) <= not a;
    layer5_outputs(6641) <= not b or a;
    layer5_outputs(6642) <= a or b;
    layer5_outputs(6643) <= a or b;
    layer5_outputs(6644) <= a;
    layer5_outputs(6645) <= not (a and b);
    layer5_outputs(6646) <= not a or b;
    layer5_outputs(6647) <= a and b;
    layer5_outputs(6648) <= a and not b;
    layer5_outputs(6649) <= a and b;
    layer5_outputs(6650) <= not b or a;
    layer5_outputs(6651) <= not a or b;
    layer5_outputs(6652) <= b;
    layer5_outputs(6653) <= not b;
    layer5_outputs(6654) <= b;
    layer5_outputs(6655) <= not (a xor b);
    layer5_outputs(6656) <= not b;
    layer5_outputs(6657) <= not a;
    layer5_outputs(6658) <= a and not b;
    layer5_outputs(6659) <= not b;
    layer5_outputs(6660) <= b and not a;
    layer5_outputs(6661) <= not a;
    layer5_outputs(6662) <= a xor b;
    layer5_outputs(6663) <= a;
    layer5_outputs(6664) <= b;
    layer5_outputs(6665) <= not (a or b);
    layer5_outputs(6666) <= not b;
    layer5_outputs(6667) <= a and not b;
    layer5_outputs(6668) <= not (a or b);
    layer5_outputs(6669) <= not a;
    layer5_outputs(6670) <= b;
    layer5_outputs(6671) <= a;
    layer5_outputs(6672) <= not (a or b);
    layer5_outputs(6673) <= not b;
    layer5_outputs(6674) <= b;
    layer5_outputs(6675) <= b;
    layer5_outputs(6676) <= not a;
    layer5_outputs(6677) <= a and b;
    layer5_outputs(6678) <= '1';
    layer5_outputs(6679) <= not a;
    layer5_outputs(6680) <= b;
    layer5_outputs(6681) <= a xor b;
    layer5_outputs(6682) <= not (a xor b);
    layer5_outputs(6683) <= a;
    layer5_outputs(6684) <= not b or a;
    layer5_outputs(6685) <= b;
    layer5_outputs(6686) <= a and not b;
    layer5_outputs(6687) <= a and not b;
    layer5_outputs(6688) <= not (a xor b);
    layer5_outputs(6689) <= not b or a;
    layer5_outputs(6690) <= not b;
    layer5_outputs(6691) <= not (a and b);
    layer5_outputs(6692) <= a;
    layer5_outputs(6693) <= not a;
    layer5_outputs(6694) <= not a;
    layer5_outputs(6695) <= not b or a;
    layer5_outputs(6696) <= not b;
    layer5_outputs(6697) <= a and not b;
    layer5_outputs(6698) <= b;
    layer5_outputs(6699) <= not b;
    layer5_outputs(6700) <= not a;
    layer5_outputs(6701) <= a xor b;
    layer5_outputs(6702) <= not (a xor b);
    layer5_outputs(6703) <= a and not b;
    layer5_outputs(6704) <= not a;
    layer5_outputs(6705) <= not (a xor b);
    layer5_outputs(6706) <= not b or a;
    layer5_outputs(6707) <= b;
    layer5_outputs(6708) <= a;
    layer5_outputs(6709) <= a;
    layer5_outputs(6710) <= not b;
    layer5_outputs(6711) <= not (a xor b);
    layer5_outputs(6712) <= not a;
    layer5_outputs(6713) <= not a or b;
    layer5_outputs(6714) <= not a;
    layer5_outputs(6715) <= not (a xor b);
    layer5_outputs(6716) <= not a;
    layer5_outputs(6717) <= not b;
    layer5_outputs(6718) <= a;
    layer5_outputs(6719) <= a and not b;
    layer5_outputs(6720) <= a xor b;
    layer5_outputs(6721) <= not b;
    layer5_outputs(6722) <= not (a and b);
    layer5_outputs(6723) <= a and b;
    layer5_outputs(6724) <= not b or a;
    layer5_outputs(6725) <= not a;
    layer5_outputs(6726) <= a xor b;
    layer5_outputs(6727) <= not b;
    layer5_outputs(6728) <= a;
    layer5_outputs(6729) <= not a or b;
    layer5_outputs(6730) <= not (a xor b);
    layer5_outputs(6731) <= not (a xor b);
    layer5_outputs(6732) <= b;
    layer5_outputs(6733) <= a xor b;
    layer5_outputs(6734) <= not b;
    layer5_outputs(6735) <= not (a and b);
    layer5_outputs(6736) <= a and not b;
    layer5_outputs(6737) <= a xor b;
    layer5_outputs(6738) <= a and b;
    layer5_outputs(6739) <= not (a or b);
    layer5_outputs(6740) <= a;
    layer5_outputs(6741) <= not (a and b);
    layer5_outputs(6742) <= a and not b;
    layer5_outputs(6743) <= not (a and b);
    layer5_outputs(6744) <= not a;
    layer5_outputs(6745) <= not a;
    layer5_outputs(6746) <= not a or b;
    layer5_outputs(6747) <= a xor b;
    layer5_outputs(6748) <= '0';
    layer5_outputs(6749) <= not b;
    layer5_outputs(6750) <= a xor b;
    layer5_outputs(6751) <= a;
    layer5_outputs(6752) <= not a;
    layer5_outputs(6753) <= a;
    layer5_outputs(6754) <= not a;
    layer5_outputs(6755) <= b;
    layer5_outputs(6756) <= b;
    layer5_outputs(6757) <= a xor b;
    layer5_outputs(6758) <= a xor b;
    layer5_outputs(6759) <= not a;
    layer5_outputs(6760) <= not (a and b);
    layer5_outputs(6761) <= b;
    layer5_outputs(6762) <= a and not b;
    layer5_outputs(6763) <= a xor b;
    layer5_outputs(6764) <= b;
    layer5_outputs(6765) <= b;
    layer5_outputs(6766) <= not (a xor b);
    layer5_outputs(6767) <= not a;
    layer5_outputs(6768) <= not a;
    layer5_outputs(6769) <= a and not b;
    layer5_outputs(6770) <= not b;
    layer5_outputs(6771) <= not (a and b);
    layer5_outputs(6772) <= a;
    layer5_outputs(6773) <= not b;
    layer5_outputs(6774) <= not (a or b);
    layer5_outputs(6775) <= b;
    layer5_outputs(6776) <= a or b;
    layer5_outputs(6777) <= not a;
    layer5_outputs(6778) <= a or b;
    layer5_outputs(6779) <= '0';
    layer5_outputs(6780) <= not (a xor b);
    layer5_outputs(6781) <= not b;
    layer5_outputs(6782) <= b;
    layer5_outputs(6783) <= not b;
    layer5_outputs(6784) <= not a;
    layer5_outputs(6785) <= a and not b;
    layer5_outputs(6786) <= not a or b;
    layer5_outputs(6787) <= a;
    layer5_outputs(6788) <= a xor b;
    layer5_outputs(6789) <= b and not a;
    layer5_outputs(6790) <= not (a and b);
    layer5_outputs(6791) <= a or b;
    layer5_outputs(6792) <= not (a xor b);
    layer5_outputs(6793) <= not a;
    layer5_outputs(6794) <= not b or a;
    layer5_outputs(6795) <= a xor b;
    layer5_outputs(6796) <= a and not b;
    layer5_outputs(6797) <= not a;
    layer5_outputs(6798) <= b;
    layer5_outputs(6799) <= not (a xor b);
    layer5_outputs(6800) <= not (a xor b);
    layer5_outputs(6801) <= not a;
    layer5_outputs(6802) <= not a or b;
    layer5_outputs(6803) <= not b or a;
    layer5_outputs(6804) <= not a;
    layer5_outputs(6805) <= not (a xor b);
    layer5_outputs(6806) <= not b;
    layer5_outputs(6807) <= not (a xor b);
    layer5_outputs(6808) <= not a;
    layer5_outputs(6809) <= b;
    layer5_outputs(6810) <= b;
    layer5_outputs(6811) <= not (a and b);
    layer5_outputs(6812) <= not a;
    layer5_outputs(6813) <= a or b;
    layer5_outputs(6814) <= not (a and b);
    layer5_outputs(6815) <= not a;
    layer5_outputs(6816) <= a and not b;
    layer5_outputs(6817) <= a;
    layer5_outputs(6818) <= b;
    layer5_outputs(6819) <= not b;
    layer5_outputs(6820) <= a and not b;
    layer5_outputs(6821) <= b;
    layer5_outputs(6822) <= a or b;
    layer5_outputs(6823) <= not b;
    layer5_outputs(6824) <= b and not a;
    layer5_outputs(6825) <= b and not a;
    layer5_outputs(6826) <= not b or a;
    layer5_outputs(6827) <= b;
    layer5_outputs(6828) <= a and b;
    layer5_outputs(6829) <= a;
    layer5_outputs(6830) <= not (a xor b);
    layer5_outputs(6831) <= not b;
    layer5_outputs(6832) <= not b or a;
    layer5_outputs(6833) <= a and b;
    layer5_outputs(6834) <= not (a and b);
    layer5_outputs(6835) <= a;
    layer5_outputs(6836) <= a;
    layer5_outputs(6837) <= not (a or b);
    layer5_outputs(6838) <= not b or a;
    layer5_outputs(6839) <= b and not a;
    layer5_outputs(6840) <= not a;
    layer5_outputs(6841) <= not b or a;
    layer5_outputs(6842) <= not (a or b);
    layer5_outputs(6843) <= a or b;
    layer5_outputs(6844) <= a xor b;
    layer5_outputs(6845) <= a and not b;
    layer5_outputs(6846) <= a and not b;
    layer5_outputs(6847) <= not b or a;
    layer5_outputs(6848) <= not a;
    layer5_outputs(6849) <= a xor b;
    layer5_outputs(6850) <= not b;
    layer5_outputs(6851) <= a;
    layer5_outputs(6852) <= not a;
    layer5_outputs(6853) <= not a;
    layer5_outputs(6854) <= a;
    layer5_outputs(6855) <= not b;
    layer5_outputs(6856) <= b and not a;
    layer5_outputs(6857) <= not a;
    layer5_outputs(6858) <= a;
    layer5_outputs(6859) <= not b;
    layer5_outputs(6860) <= not (a or b);
    layer5_outputs(6861) <= not (a and b);
    layer5_outputs(6862) <= not (a xor b);
    layer5_outputs(6863) <= a xor b;
    layer5_outputs(6864) <= not (a or b);
    layer5_outputs(6865) <= not a or b;
    layer5_outputs(6866) <= not a;
    layer5_outputs(6867) <= a or b;
    layer5_outputs(6868) <= not (a xor b);
    layer5_outputs(6869) <= b and not a;
    layer5_outputs(6870) <= a xor b;
    layer5_outputs(6871) <= not b or a;
    layer5_outputs(6872) <= a xor b;
    layer5_outputs(6873) <= a;
    layer5_outputs(6874) <= not a;
    layer5_outputs(6875) <= b;
    layer5_outputs(6876) <= not (a xor b);
    layer5_outputs(6877) <= not (a or b);
    layer5_outputs(6878) <= not b or a;
    layer5_outputs(6879) <= a;
    layer5_outputs(6880) <= not a;
    layer5_outputs(6881) <= not (a xor b);
    layer5_outputs(6882) <= a xor b;
    layer5_outputs(6883) <= not (a and b);
    layer5_outputs(6884) <= not b;
    layer5_outputs(6885) <= a or b;
    layer5_outputs(6886) <= b and not a;
    layer5_outputs(6887) <= not a or b;
    layer5_outputs(6888) <= not (a xor b);
    layer5_outputs(6889) <= not b;
    layer5_outputs(6890) <= not b;
    layer5_outputs(6891) <= not (a or b);
    layer5_outputs(6892) <= not a;
    layer5_outputs(6893) <= not (a and b);
    layer5_outputs(6894) <= a;
    layer5_outputs(6895) <= not a or b;
    layer5_outputs(6896) <= not (a and b);
    layer5_outputs(6897) <= b;
    layer5_outputs(6898) <= b;
    layer5_outputs(6899) <= a or b;
    layer5_outputs(6900) <= a and b;
    layer5_outputs(6901) <= not a;
    layer5_outputs(6902) <= a;
    layer5_outputs(6903) <= '1';
    layer5_outputs(6904) <= b;
    layer5_outputs(6905) <= not b;
    layer5_outputs(6906) <= b;
    layer5_outputs(6907) <= b and not a;
    layer5_outputs(6908) <= '0';
    layer5_outputs(6909) <= a or b;
    layer5_outputs(6910) <= not a;
    layer5_outputs(6911) <= not (a xor b);
    layer5_outputs(6912) <= a or b;
    layer5_outputs(6913) <= a and not b;
    layer5_outputs(6914) <= not (a xor b);
    layer5_outputs(6915) <= a;
    layer5_outputs(6916) <= not b;
    layer5_outputs(6917) <= a xor b;
    layer5_outputs(6918) <= not a;
    layer5_outputs(6919) <= a;
    layer5_outputs(6920) <= not b;
    layer5_outputs(6921) <= not (a xor b);
    layer5_outputs(6922) <= a;
    layer5_outputs(6923) <= not (a or b);
    layer5_outputs(6924) <= a and not b;
    layer5_outputs(6925) <= a xor b;
    layer5_outputs(6926) <= not a or b;
    layer5_outputs(6927) <= a and not b;
    layer5_outputs(6928) <= not a;
    layer5_outputs(6929) <= not b;
    layer5_outputs(6930) <= not (a or b);
    layer5_outputs(6931) <= a;
    layer5_outputs(6932) <= not a or b;
    layer5_outputs(6933) <= not (a or b);
    layer5_outputs(6934) <= not a;
    layer5_outputs(6935) <= a or b;
    layer5_outputs(6936) <= a xor b;
    layer5_outputs(6937) <= a and not b;
    layer5_outputs(6938) <= a and b;
    layer5_outputs(6939) <= not a;
    layer5_outputs(6940) <= b;
    layer5_outputs(6941) <= not (a and b);
    layer5_outputs(6942) <= b;
    layer5_outputs(6943) <= not b or a;
    layer5_outputs(6944) <= b;
    layer5_outputs(6945) <= a;
    layer5_outputs(6946) <= a;
    layer5_outputs(6947) <= a;
    layer5_outputs(6948) <= b;
    layer5_outputs(6949) <= not (a xor b);
    layer5_outputs(6950) <= a or b;
    layer5_outputs(6951) <= a xor b;
    layer5_outputs(6952) <= a;
    layer5_outputs(6953) <= not a;
    layer5_outputs(6954) <= b;
    layer5_outputs(6955) <= not a;
    layer5_outputs(6956) <= a;
    layer5_outputs(6957) <= a;
    layer5_outputs(6958) <= not (a xor b);
    layer5_outputs(6959) <= b and not a;
    layer5_outputs(6960) <= a and b;
    layer5_outputs(6961) <= b;
    layer5_outputs(6962) <= a and not b;
    layer5_outputs(6963) <= a xor b;
    layer5_outputs(6964) <= b;
    layer5_outputs(6965) <= a and b;
    layer5_outputs(6966) <= a and not b;
    layer5_outputs(6967) <= a;
    layer5_outputs(6968) <= not b;
    layer5_outputs(6969) <= not (a xor b);
    layer5_outputs(6970) <= b;
    layer5_outputs(6971) <= a and not b;
    layer5_outputs(6972) <= '0';
    layer5_outputs(6973) <= not a;
    layer5_outputs(6974) <= '0';
    layer5_outputs(6975) <= not (a or b);
    layer5_outputs(6976) <= a and b;
    layer5_outputs(6977) <= a;
    layer5_outputs(6978) <= a and not b;
    layer5_outputs(6979) <= not (a xor b);
    layer5_outputs(6980) <= b;
    layer5_outputs(6981) <= not (a or b);
    layer5_outputs(6982) <= not b;
    layer5_outputs(6983) <= a or b;
    layer5_outputs(6984) <= not a or b;
    layer5_outputs(6985) <= not (a and b);
    layer5_outputs(6986) <= a or b;
    layer5_outputs(6987) <= a;
    layer5_outputs(6988) <= not (a xor b);
    layer5_outputs(6989) <= a;
    layer5_outputs(6990) <= not b;
    layer5_outputs(6991) <= b;
    layer5_outputs(6992) <= not b or a;
    layer5_outputs(6993) <= not a or b;
    layer5_outputs(6994) <= not (a or b);
    layer5_outputs(6995) <= a and not b;
    layer5_outputs(6996) <= not (a or b);
    layer5_outputs(6997) <= b;
    layer5_outputs(6998) <= a and b;
    layer5_outputs(6999) <= not a;
    layer5_outputs(7000) <= a or b;
    layer5_outputs(7001) <= not (a and b);
    layer5_outputs(7002) <= b and not a;
    layer5_outputs(7003) <= not (a and b);
    layer5_outputs(7004) <= not (a xor b);
    layer5_outputs(7005) <= b and not a;
    layer5_outputs(7006) <= not a or b;
    layer5_outputs(7007) <= not a;
    layer5_outputs(7008) <= not a;
    layer5_outputs(7009) <= b;
    layer5_outputs(7010) <= a and b;
    layer5_outputs(7011) <= not a;
    layer5_outputs(7012) <= not b or a;
    layer5_outputs(7013) <= not a;
    layer5_outputs(7014) <= not (a or b);
    layer5_outputs(7015) <= not a;
    layer5_outputs(7016) <= not b;
    layer5_outputs(7017) <= a;
    layer5_outputs(7018) <= not a;
    layer5_outputs(7019) <= a and b;
    layer5_outputs(7020) <= a xor b;
    layer5_outputs(7021) <= a xor b;
    layer5_outputs(7022) <= '1';
    layer5_outputs(7023) <= a or b;
    layer5_outputs(7024) <= a and not b;
    layer5_outputs(7025) <= not (a xor b);
    layer5_outputs(7026) <= a and b;
    layer5_outputs(7027) <= a;
    layer5_outputs(7028) <= a and b;
    layer5_outputs(7029) <= a xor b;
    layer5_outputs(7030) <= not (a and b);
    layer5_outputs(7031) <= b;
    layer5_outputs(7032) <= a;
    layer5_outputs(7033) <= not a;
    layer5_outputs(7034) <= a;
    layer5_outputs(7035) <= b and not a;
    layer5_outputs(7036) <= a or b;
    layer5_outputs(7037) <= b;
    layer5_outputs(7038) <= not (a xor b);
    layer5_outputs(7039) <= not (a xor b);
    layer5_outputs(7040) <= not a;
    layer5_outputs(7041) <= a;
    layer5_outputs(7042) <= a or b;
    layer5_outputs(7043) <= not a or b;
    layer5_outputs(7044) <= not b or a;
    layer5_outputs(7045) <= not a;
    layer5_outputs(7046) <= not b;
    layer5_outputs(7047) <= b;
    layer5_outputs(7048) <= a and b;
    layer5_outputs(7049) <= a;
    layer5_outputs(7050) <= not a;
    layer5_outputs(7051) <= a and not b;
    layer5_outputs(7052) <= a xor b;
    layer5_outputs(7053) <= not (a xor b);
    layer5_outputs(7054) <= a or b;
    layer5_outputs(7055) <= a xor b;
    layer5_outputs(7056) <= not a;
    layer5_outputs(7057) <= not (a and b);
    layer5_outputs(7058) <= a xor b;
    layer5_outputs(7059) <= not b;
    layer5_outputs(7060) <= not b;
    layer5_outputs(7061) <= not a;
    layer5_outputs(7062) <= a;
    layer5_outputs(7063) <= a and not b;
    layer5_outputs(7064) <= a and b;
    layer5_outputs(7065) <= b and not a;
    layer5_outputs(7066) <= a and not b;
    layer5_outputs(7067) <= a and b;
    layer5_outputs(7068) <= not (a xor b);
    layer5_outputs(7069) <= not a or b;
    layer5_outputs(7070) <= a and b;
    layer5_outputs(7071) <= a;
    layer5_outputs(7072) <= not b;
    layer5_outputs(7073) <= a and not b;
    layer5_outputs(7074) <= not a or b;
    layer5_outputs(7075) <= not (a and b);
    layer5_outputs(7076) <= not a;
    layer5_outputs(7077) <= not (a or b);
    layer5_outputs(7078) <= not a or b;
    layer5_outputs(7079) <= a or b;
    layer5_outputs(7080) <= b;
    layer5_outputs(7081) <= not b;
    layer5_outputs(7082) <= a and not b;
    layer5_outputs(7083) <= a and b;
    layer5_outputs(7084) <= not b;
    layer5_outputs(7085) <= b;
    layer5_outputs(7086) <= b;
    layer5_outputs(7087) <= not b;
    layer5_outputs(7088) <= not b or a;
    layer5_outputs(7089) <= a;
    layer5_outputs(7090) <= b;
    layer5_outputs(7091) <= '1';
    layer5_outputs(7092) <= a xor b;
    layer5_outputs(7093) <= a xor b;
    layer5_outputs(7094) <= a;
    layer5_outputs(7095) <= not (a xor b);
    layer5_outputs(7096) <= b and not a;
    layer5_outputs(7097) <= not (a or b);
    layer5_outputs(7098) <= not (a and b);
    layer5_outputs(7099) <= not b;
    layer5_outputs(7100) <= b and not a;
    layer5_outputs(7101) <= b;
    layer5_outputs(7102) <= a;
    layer5_outputs(7103) <= not a or b;
    layer5_outputs(7104) <= a xor b;
    layer5_outputs(7105) <= not a;
    layer5_outputs(7106) <= not a;
    layer5_outputs(7107) <= a and b;
    layer5_outputs(7108) <= not a;
    layer5_outputs(7109) <= not a or b;
    layer5_outputs(7110) <= not b;
    layer5_outputs(7111) <= not b;
    layer5_outputs(7112) <= not a;
    layer5_outputs(7113) <= a or b;
    layer5_outputs(7114) <= b;
    layer5_outputs(7115) <= not a;
    layer5_outputs(7116) <= not a;
    layer5_outputs(7117) <= a;
    layer5_outputs(7118) <= a xor b;
    layer5_outputs(7119) <= a xor b;
    layer5_outputs(7120) <= not a or b;
    layer5_outputs(7121) <= not b;
    layer5_outputs(7122) <= not (a xor b);
    layer5_outputs(7123) <= not (a and b);
    layer5_outputs(7124) <= b;
    layer5_outputs(7125) <= a and not b;
    layer5_outputs(7126) <= b and not a;
    layer5_outputs(7127) <= not a or b;
    layer5_outputs(7128) <= not b or a;
    layer5_outputs(7129) <= not b or a;
    layer5_outputs(7130) <= not a;
    layer5_outputs(7131) <= not b or a;
    layer5_outputs(7132) <= b and not a;
    layer5_outputs(7133) <= a;
    layer5_outputs(7134) <= a;
    layer5_outputs(7135) <= not (a xor b);
    layer5_outputs(7136) <= a;
    layer5_outputs(7137) <= not (a xor b);
    layer5_outputs(7138) <= not b;
    layer5_outputs(7139) <= not a;
    layer5_outputs(7140) <= '0';
    layer5_outputs(7141) <= a;
    layer5_outputs(7142) <= b;
    layer5_outputs(7143) <= a or b;
    layer5_outputs(7144) <= not (a xor b);
    layer5_outputs(7145) <= not a;
    layer5_outputs(7146) <= not b;
    layer5_outputs(7147) <= not a;
    layer5_outputs(7148) <= not a or b;
    layer5_outputs(7149) <= not b;
    layer5_outputs(7150) <= not (a and b);
    layer5_outputs(7151) <= b;
    layer5_outputs(7152) <= b;
    layer5_outputs(7153) <= b;
    layer5_outputs(7154) <= a;
    layer5_outputs(7155) <= not (a or b);
    layer5_outputs(7156) <= not b;
    layer5_outputs(7157) <= not a;
    layer5_outputs(7158) <= a and not b;
    layer5_outputs(7159) <= a and b;
    layer5_outputs(7160) <= not b or a;
    layer5_outputs(7161) <= b;
    layer5_outputs(7162) <= b;
    layer5_outputs(7163) <= a;
    layer5_outputs(7164) <= a and not b;
    layer5_outputs(7165) <= not b or a;
    layer5_outputs(7166) <= a xor b;
    layer5_outputs(7167) <= b;
    layer5_outputs(7168) <= '1';
    layer5_outputs(7169) <= b;
    layer5_outputs(7170) <= not (a and b);
    layer5_outputs(7171) <= a and not b;
    layer5_outputs(7172) <= not a;
    layer5_outputs(7173) <= b and not a;
    layer5_outputs(7174) <= a;
    layer5_outputs(7175) <= not (a or b);
    layer5_outputs(7176) <= not a or b;
    layer5_outputs(7177) <= not b;
    layer5_outputs(7178) <= b and not a;
    layer5_outputs(7179) <= not a;
    layer5_outputs(7180) <= b and not a;
    layer5_outputs(7181) <= b;
    layer5_outputs(7182) <= not a or b;
    layer5_outputs(7183) <= not (a xor b);
    layer5_outputs(7184) <= a;
    layer5_outputs(7185) <= a xor b;
    layer5_outputs(7186) <= b and not a;
    layer5_outputs(7187) <= b;
    layer5_outputs(7188) <= b;
    layer5_outputs(7189) <= not b or a;
    layer5_outputs(7190) <= not a;
    layer5_outputs(7191) <= b;
    layer5_outputs(7192) <= a;
    layer5_outputs(7193) <= not a or b;
    layer5_outputs(7194) <= not (a and b);
    layer5_outputs(7195) <= a xor b;
    layer5_outputs(7196) <= a and not b;
    layer5_outputs(7197) <= a;
    layer5_outputs(7198) <= a and b;
    layer5_outputs(7199) <= b;
    layer5_outputs(7200) <= a;
    layer5_outputs(7201) <= not b;
    layer5_outputs(7202) <= b and not a;
    layer5_outputs(7203) <= not a;
    layer5_outputs(7204) <= not b;
    layer5_outputs(7205) <= not (a xor b);
    layer5_outputs(7206) <= not b;
    layer5_outputs(7207) <= b;
    layer5_outputs(7208) <= not b;
    layer5_outputs(7209) <= b;
    layer5_outputs(7210) <= a and not b;
    layer5_outputs(7211) <= not (a or b);
    layer5_outputs(7212) <= not (a xor b);
    layer5_outputs(7213) <= not b or a;
    layer5_outputs(7214) <= not (a and b);
    layer5_outputs(7215) <= a and not b;
    layer5_outputs(7216) <= not (a xor b);
    layer5_outputs(7217) <= b;
    layer5_outputs(7218) <= not b;
    layer5_outputs(7219) <= a or b;
    layer5_outputs(7220) <= a and b;
    layer5_outputs(7221) <= a;
    layer5_outputs(7222) <= a;
    layer5_outputs(7223) <= a and b;
    layer5_outputs(7224) <= not b or a;
    layer5_outputs(7225) <= a xor b;
    layer5_outputs(7226) <= not b or a;
    layer5_outputs(7227) <= a and b;
    layer5_outputs(7228) <= not a;
    layer5_outputs(7229) <= not (a xor b);
    layer5_outputs(7230) <= not b or a;
    layer5_outputs(7231) <= b;
    layer5_outputs(7232) <= a or b;
    layer5_outputs(7233) <= a and not b;
    layer5_outputs(7234) <= not a;
    layer5_outputs(7235) <= not b;
    layer5_outputs(7236) <= not a;
    layer5_outputs(7237) <= not (a xor b);
    layer5_outputs(7238) <= not b or a;
    layer5_outputs(7239) <= b and not a;
    layer5_outputs(7240) <= a or b;
    layer5_outputs(7241) <= not b or a;
    layer5_outputs(7242) <= not a;
    layer5_outputs(7243) <= b and not a;
    layer5_outputs(7244) <= b;
    layer5_outputs(7245) <= not a or b;
    layer5_outputs(7246) <= a xor b;
    layer5_outputs(7247) <= not a;
    layer5_outputs(7248) <= not b;
    layer5_outputs(7249) <= not b or a;
    layer5_outputs(7250) <= a and not b;
    layer5_outputs(7251) <= not (a or b);
    layer5_outputs(7252) <= b;
    layer5_outputs(7253) <= not a or b;
    layer5_outputs(7254) <= a xor b;
    layer5_outputs(7255) <= not (a and b);
    layer5_outputs(7256) <= a and b;
    layer5_outputs(7257) <= not (a xor b);
    layer5_outputs(7258) <= not (a xor b);
    layer5_outputs(7259) <= not a or b;
    layer5_outputs(7260) <= a xor b;
    layer5_outputs(7261) <= not a or b;
    layer5_outputs(7262) <= b;
    layer5_outputs(7263) <= not b or a;
    layer5_outputs(7264) <= not a;
    layer5_outputs(7265) <= a;
    layer5_outputs(7266) <= not (a and b);
    layer5_outputs(7267) <= a xor b;
    layer5_outputs(7268) <= a;
    layer5_outputs(7269) <= a xor b;
    layer5_outputs(7270) <= a xor b;
    layer5_outputs(7271) <= not (a xor b);
    layer5_outputs(7272) <= a;
    layer5_outputs(7273) <= a or b;
    layer5_outputs(7274) <= a and not b;
    layer5_outputs(7275) <= a and not b;
    layer5_outputs(7276) <= not (a or b);
    layer5_outputs(7277) <= not (a and b);
    layer5_outputs(7278) <= not a or b;
    layer5_outputs(7279) <= not b;
    layer5_outputs(7280) <= not (a and b);
    layer5_outputs(7281) <= not (a and b);
    layer5_outputs(7282) <= not b or a;
    layer5_outputs(7283) <= a;
    layer5_outputs(7284) <= b;
    layer5_outputs(7285) <= a;
    layer5_outputs(7286) <= not (a or b);
    layer5_outputs(7287) <= a xor b;
    layer5_outputs(7288) <= not (a or b);
    layer5_outputs(7289) <= b and not a;
    layer5_outputs(7290) <= not (a xor b);
    layer5_outputs(7291) <= not (a xor b);
    layer5_outputs(7292) <= not a;
    layer5_outputs(7293) <= not a or b;
    layer5_outputs(7294) <= not a or b;
    layer5_outputs(7295) <= not a;
    layer5_outputs(7296) <= not b or a;
    layer5_outputs(7297) <= a xor b;
    layer5_outputs(7298) <= a;
    layer5_outputs(7299) <= not b;
    layer5_outputs(7300) <= not b or a;
    layer5_outputs(7301) <= b;
    layer5_outputs(7302) <= not b;
    layer5_outputs(7303) <= not (a xor b);
    layer5_outputs(7304) <= not a;
    layer5_outputs(7305) <= not (a xor b);
    layer5_outputs(7306) <= not a;
    layer5_outputs(7307) <= a or b;
    layer5_outputs(7308) <= a or b;
    layer5_outputs(7309) <= b;
    layer5_outputs(7310) <= a or b;
    layer5_outputs(7311) <= not b;
    layer5_outputs(7312) <= not (a or b);
    layer5_outputs(7313) <= not a;
    layer5_outputs(7314) <= b and not a;
    layer5_outputs(7315) <= not a or b;
    layer5_outputs(7316) <= a or b;
    layer5_outputs(7317) <= not (a and b);
    layer5_outputs(7318) <= b;
    layer5_outputs(7319) <= a;
    layer5_outputs(7320) <= a;
    layer5_outputs(7321) <= b;
    layer5_outputs(7322) <= b and not a;
    layer5_outputs(7323) <= not b;
    layer5_outputs(7324) <= not (a or b);
    layer5_outputs(7325) <= b;
    layer5_outputs(7326) <= not (a or b);
    layer5_outputs(7327) <= not a;
    layer5_outputs(7328) <= not b or a;
    layer5_outputs(7329) <= b;
    layer5_outputs(7330) <= '1';
    layer5_outputs(7331) <= a and b;
    layer5_outputs(7332) <= a xor b;
    layer5_outputs(7333) <= a;
    layer5_outputs(7334) <= not (a xor b);
    layer5_outputs(7335) <= b and not a;
    layer5_outputs(7336) <= not a;
    layer5_outputs(7337) <= not (a xor b);
    layer5_outputs(7338) <= not a;
    layer5_outputs(7339) <= not b;
    layer5_outputs(7340) <= b;
    layer5_outputs(7341) <= a and b;
    layer5_outputs(7342) <= not b;
    layer5_outputs(7343) <= a;
    layer5_outputs(7344) <= b;
    layer5_outputs(7345) <= b;
    layer5_outputs(7346) <= not a;
    layer5_outputs(7347) <= a or b;
    layer5_outputs(7348) <= not a;
    layer5_outputs(7349) <= not b or a;
    layer5_outputs(7350) <= not (a or b);
    layer5_outputs(7351) <= a and b;
    layer5_outputs(7352) <= not (a xor b);
    layer5_outputs(7353) <= b;
    layer5_outputs(7354) <= not (a xor b);
    layer5_outputs(7355) <= a xor b;
    layer5_outputs(7356) <= not (a xor b);
    layer5_outputs(7357) <= a;
    layer5_outputs(7358) <= b;
    layer5_outputs(7359) <= b;
    layer5_outputs(7360) <= '0';
    layer5_outputs(7361) <= not a or b;
    layer5_outputs(7362) <= a;
    layer5_outputs(7363) <= b;
    layer5_outputs(7364) <= b;
    layer5_outputs(7365) <= a;
    layer5_outputs(7366) <= not (a or b);
    layer5_outputs(7367) <= a;
    layer5_outputs(7368) <= not b;
    layer5_outputs(7369) <= '1';
    layer5_outputs(7370) <= not (a and b);
    layer5_outputs(7371) <= not (a xor b);
    layer5_outputs(7372) <= not (a xor b);
    layer5_outputs(7373) <= not a or b;
    layer5_outputs(7374) <= not b or a;
    layer5_outputs(7375) <= not a;
    layer5_outputs(7376) <= not (a or b);
    layer5_outputs(7377) <= not b;
    layer5_outputs(7378) <= a and b;
    layer5_outputs(7379) <= not (a xor b);
    layer5_outputs(7380) <= '0';
    layer5_outputs(7381) <= not b;
    layer5_outputs(7382) <= b;
    layer5_outputs(7383) <= b;
    layer5_outputs(7384) <= not (a and b);
    layer5_outputs(7385) <= a;
    layer5_outputs(7386) <= not a or b;
    layer5_outputs(7387) <= a xor b;
    layer5_outputs(7388) <= '0';
    layer5_outputs(7389) <= not b;
    layer5_outputs(7390) <= b;
    layer5_outputs(7391) <= not a or b;
    layer5_outputs(7392) <= not b;
    layer5_outputs(7393) <= not (a or b);
    layer5_outputs(7394) <= not a or b;
    layer5_outputs(7395) <= a;
    layer5_outputs(7396) <= a;
    layer5_outputs(7397) <= not a or b;
    layer5_outputs(7398) <= not b or a;
    layer5_outputs(7399) <= not (a xor b);
    layer5_outputs(7400) <= not b;
    layer5_outputs(7401) <= a and not b;
    layer5_outputs(7402) <= a or b;
    layer5_outputs(7403) <= a and not b;
    layer5_outputs(7404) <= b;
    layer5_outputs(7405) <= a;
    layer5_outputs(7406) <= b;
    layer5_outputs(7407) <= a;
    layer5_outputs(7408) <= not (a xor b);
    layer5_outputs(7409) <= not b or a;
    layer5_outputs(7410) <= not (a and b);
    layer5_outputs(7411) <= not b;
    layer5_outputs(7412) <= a or b;
    layer5_outputs(7413) <= '1';
    layer5_outputs(7414) <= not b;
    layer5_outputs(7415) <= b and not a;
    layer5_outputs(7416) <= not a or b;
    layer5_outputs(7417) <= not (a xor b);
    layer5_outputs(7418) <= a;
    layer5_outputs(7419) <= '1';
    layer5_outputs(7420) <= not (a or b);
    layer5_outputs(7421) <= not a or b;
    layer5_outputs(7422) <= not a or b;
    layer5_outputs(7423) <= a and not b;
    layer5_outputs(7424) <= a and not b;
    layer5_outputs(7425) <= not b;
    layer5_outputs(7426) <= a;
    layer5_outputs(7427) <= not a or b;
    layer5_outputs(7428) <= not a or b;
    layer5_outputs(7429) <= not b;
    layer5_outputs(7430) <= b and not a;
    layer5_outputs(7431) <= a xor b;
    layer5_outputs(7432) <= a and not b;
    layer5_outputs(7433) <= not (a or b);
    layer5_outputs(7434) <= a and not b;
    layer5_outputs(7435) <= a;
    layer5_outputs(7436) <= not b;
    layer5_outputs(7437) <= not (a xor b);
    layer5_outputs(7438) <= not b;
    layer5_outputs(7439) <= a;
    layer5_outputs(7440) <= not a;
    layer5_outputs(7441) <= a xor b;
    layer5_outputs(7442) <= not b or a;
    layer5_outputs(7443) <= not a;
    layer5_outputs(7444) <= not b;
    layer5_outputs(7445) <= not a;
    layer5_outputs(7446) <= a;
    layer5_outputs(7447) <= b;
    layer5_outputs(7448) <= not a;
    layer5_outputs(7449) <= not a;
    layer5_outputs(7450) <= a;
    layer5_outputs(7451) <= b and not a;
    layer5_outputs(7452) <= a;
    layer5_outputs(7453) <= a and b;
    layer5_outputs(7454) <= not (a or b);
    layer5_outputs(7455) <= not a or b;
    layer5_outputs(7456) <= a;
    layer5_outputs(7457) <= a;
    layer5_outputs(7458) <= a and b;
    layer5_outputs(7459) <= not a or b;
    layer5_outputs(7460) <= b and not a;
    layer5_outputs(7461) <= not (a xor b);
    layer5_outputs(7462) <= not a or b;
    layer5_outputs(7463) <= not a;
    layer5_outputs(7464) <= not (a or b);
    layer5_outputs(7465) <= b and not a;
    layer5_outputs(7466) <= a and not b;
    layer5_outputs(7467) <= not a;
    layer5_outputs(7468) <= a and b;
    layer5_outputs(7469) <= not b or a;
    layer5_outputs(7470) <= a xor b;
    layer5_outputs(7471) <= not b;
    layer5_outputs(7472) <= a xor b;
    layer5_outputs(7473) <= not a;
    layer5_outputs(7474) <= b;
    layer5_outputs(7475) <= not b;
    layer5_outputs(7476) <= a;
    layer5_outputs(7477) <= not a;
    layer5_outputs(7478) <= a;
    layer5_outputs(7479) <= b;
    layer5_outputs(7480) <= not (a or b);
    layer5_outputs(7481) <= not a;
    layer5_outputs(7482) <= not a;
    layer5_outputs(7483) <= a and b;
    layer5_outputs(7484) <= not b;
    layer5_outputs(7485) <= not b or a;
    layer5_outputs(7486) <= not b;
    layer5_outputs(7487) <= not (a xor b);
    layer5_outputs(7488) <= not a or b;
    layer5_outputs(7489) <= not (a and b);
    layer5_outputs(7490) <= a and not b;
    layer5_outputs(7491) <= a and not b;
    layer5_outputs(7492) <= a;
    layer5_outputs(7493) <= not b;
    layer5_outputs(7494) <= not (a or b);
    layer5_outputs(7495) <= not (a or b);
    layer5_outputs(7496) <= a xor b;
    layer5_outputs(7497) <= not a;
    layer5_outputs(7498) <= not (a and b);
    layer5_outputs(7499) <= b and not a;
    layer5_outputs(7500) <= a;
    layer5_outputs(7501) <= not a or b;
    layer5_outputs(7502) <= not (a or b);
    layer5_outputs(7503) <= not (a or b);
    layer5_outputs(7504) <= not b;
    layer5_outputs(7505) <= b and not a;
    layer5_outputs(7506) <= b;
    layer5_outputs(7507) <= b and not a;
    layer5_outputs(7508) <= a xor b;
    layer5_outputs(7509) <= b;
    layer5_outputs(7510) <= a;
    layer5_outputs(7511) <= not b;
    layer5_outputs(7512) <= b;
    layer5_outputs(7513) <= not (a xor b);
    layer5_outputs(7514) <= a or b;
    layer5_outputs(7515) <= b;
    layer5_outputs(7516) <= a;
    layer5_outputs(7517) <= not b;
    layer5_outputs(7518) <= not (a or b);
    layer5_outputs(7519) <= not b;
    layer5_outputs(7520) <= not b or a;
    layer5_outputs(7521) <= not a;
    layer5_outputs(7522) <= not (a or b);
    layer5_outputs(7523) <= b;
    layer5_outputs(7524) <= not a;
    layer5_outputs(7525) <= a;
    layer5_outputs(7526) <= not b;
    layer5_outputs(7527) <= a;
    layer5_outputs(7528) <= a;
    layer5_outputs(7529) <= not a or b;
    layer5_outputs(7530) <= not a;
    layer5_outputs(7531) <= b;
    layer5_outputs(7532) <= not b or a;
    layer5_outputs(7533) <= not b;
    layer5_outputs(7534) <= a and b;
    layer5_outputs(7535) <= b and not a;
    layer5_outputs(7536) <= a or b;
    layer5_outputs(7537) <= not (a xor b);
    layer5_outputs(7538) <= b;
    layer5_outputs(7539) <= a;
    layer5_outputs(7540) <= a xor b;
    layer5_outputs(7541) <= b;
    layer5_outputs(7542) <= b;
    layer5_outputs(7543) <= not b or a;
    layer5_outputs(7544) <= not a;
    layer5_outputs(7545) <= a;
    layer5_outputs(7546) <= not (a xor b);
    layer5_outputs(7547) <= not (a and b);
    layer5_outputs(7548) <= a and not b;
    layer5_outputs(7549) <= not b or a;
    layer5_outputs(7550) <= a and not b;
    layer5_outputs(7551) <= b;
    layer5_outputs(7552) <= a and b;
    layer5_outputs(7553) <= not a;
    layer5_outputs(7554) <= not a;
    layer5_outputs(7555) <= not a;
    layer5_outputs(7556) <= a or b;
    layer5_outputs(7557) <= '0';
    layer5_outputs(7558) <= a xor b;
    layer5_outputs(7559) <= not (a and b);
    layer5_outputs(7560) <= not a;
    layer5_outputs(7561) <= b;
    layer5_outputs(7562) <= not b;
    layer5_outputs(7563) <= b;
    layer5_outputs(7564) <= not (a and b);
    layer5_outputs(7565) <= b;
    layer5_outputs(7566) <= not a;
    layer5_outputs(7567) <= b and not a;
    layer5_outputs(7568) <= not b or a;
    layer5_outputs(7569) <= b and not a;
    layer5_outputs(7570) <= a or b;
    layer5_outputs(7571) <= b;
    layer5_outputs(7572) <= not a or b;
    layer5_outputs(7573) <= a or b;
    layer5_outputs(7574) <= '0';
    layer5_outputs(7575) <= not (a and b);
    layer5_outputs(7576) <= not (a or b);
    layer5_outputs(7577) <= not a;
    layer5_outputs(7578) <= b and not a;
    layer5_outputs(7579) <= a xor b;
    layer5_outputs(7580) <= not a;
    layer5_outputs(7581) <= not b or a;
    layer5_outputs(7582) <= not a;
    layer5_outputs(7583) <= not a or b;
    layer5_outputs(7584) <= a xor b;
    layer5_outputs(7585) <= not (a and b);
    layer5_outputs(7586) <= a and b;
    layer5_outputs(7587) <= a xor b;
    layer5_outputs(7588) <= a and b;
    layer5_outputs(7589) <= not b;
    layer5_outputs(7590) <= not b;
    layer5_outputs(7591) <= a or b;
    layer5_outputs(7592) <= not a;
    layer5_outputs(7593) <= a and b;
    layer5_outputs(7594) <= b;
    layer5_outputs(7595) <= a or b;
    layer5_outputs(7596) <= not b;
    layer5_outputs(7597) <= not a;
    layer5_outputs(7598) <= not (a xor b);
    layer5_outputs(7599) <= b;
    layer5_outputs(7600) <= a and not b;
    layer5_outputs(7601) <= a and not b;
    layer5_outputs(7602) <= a and not b;
    layer5_outputs(7603) <= a and not b;
    layer5_outputs(7604) <= a;
    layer5_outputs(7605) <= a or b;
    layer5_outputs(7606) <= not a;
    layer5_outputs(7607) <= b;
    layer5_outputs(7608) <= a or b;
    layer5_outputs(7609) <= not (a or b);
    layer5_outputs(7610) <= not b or a;
    layer5_outputs(7611) <= not a or b;
    layer5_outputs(7612) <= not b;
    layer5_outputs(7613) <= a or b;
    layer5_outputs(7614) <= b and not a;
    layer5_outputs(7615) <= not b;
    layer5_outputs(7616) <= a;
    layer5_outputs(7617) <= a and not b;
    layer5_outputs(7618) <= a and b;
    layer5_outputs(7619) <= not (a or b);
    layer5_outputs(7620) <= a or b;
    layer5_outputs(7621) <= not a;
    layer5_outputs(7622) <= not b;
    layer5_outputs(7623) <= a and b;
    layer5_outputs(7624) <= a or b;
    layer5_outputs(7625) <= a;
    layer5_outputs(7626) <= a and b;
    layer5_outputs(7627) <= a and b;
    layer5_outputs(7628) <= '1';
    layer5_outputs(7629) <= not a;
    layer5_outputs(7630) <= not a;
    layer5_outputs(7631) <= not a;
    layer5_outputs(7632) <= not (a xor b);
    layer5_outputs(7633) <= not a;
    layer5_outputs(7634) <= not a;
    layer5_outputs(7635) <= not a or b;
    layer5_outputs(7636) <= not b;
    layer5_outputs(7637) <= a;
    layer5_outputs(7638) <= not a or b;
    layer5_outputs(7639) <= not b;
    layer5_outputs(7640) <= a xor b;
    layer5_outputs(7641) <= b and not a;
    layer5_outputs(7642) <= not (a and b);
    layer5_outputs(7643) <= not b;
    layer5_outputs(7644) <= not (a and b);
    layer5_outputs(7645) <= not (a and b);
    layer5_outputs(7646) <= not (a or b);
    layer5_outputs(7647) <= a;
    layer5_outputs(7648) <= b and not a;
    layer5_outputs(7649) <= a;
    layer5_outputs(7650) <= not a;
    layer5_outputs(7651) <= a;
    layer5_outputs(7652) <= b;
    layer5_outputs(7653) <= not (a and b);
    layer5_outputs(7654) <= '1';
    layer5_outputs(7655) <= b;
    layer5_outputs(7656) <= b and not a;
    layer5_outputs(7657) <= a and not b;
    layer5_outputs(7658) <= a;
    layer5_outputs(7659) <= not (a xor b);
    layer5_outputs(7660) <= not (a and b);
    layer5_outputs(7661) <= b and not a;
    layer5_outputs(7662) <= b and not a;
    layer5_outputs(7663) <= not b;
    layer5_outputs(7664) <= b;
    layer5_outputs(7665) <= not b;
    layer5_outputs(7666) <= not b;
    layer5_outputs(7667) <= b;
    layer5_outputs(7668) <= not (a or b);
    layer5_outputs(7669) <= not (a xor b);
    layer5_outputs(7670) <= not a or b;
    layer5_outputs(7671) <= b and not a;
    layer5_outputs(7672) <= a and b;
    layer5_outputs(7673) <= not a or b;
    layer5_outputs(7674) <= b and not a;
    layer5_outputs(7675) <= not a;
    layer5_outputs(7676) <= b and not a;
    layer5_outputs(7677) <= a xor b;
    layer5_outputs(7678) <= a and not b;
    layer5_outputs(7679) <= not (a and b);
    layer5_outputs(7680) <= a;
    layer5_outputs(7681) <= a;
    layer5_outputs(7682) <= not (a xor b);
    layer5_outputs(7683) <= not a or b;
    layer5_outputs(7684) <= b;
    layer5_outputs(7685) <= not b;
    layer5_outputs(7686) <= a;
    layer5_outputs(7687) <= a or b;
    layer5_outputs(7688) <= b;
    layer5_outputs(7689) <= a;
    layer5_outputs(7690) <= b;
    layer5_outputs(7691) <= not b;
    layer5_outputs(7692) <= a xor b;
    layer5_outputs(7693) <= b;
    layer5_outputs(7694) <= a;
    layer5_outputs(7695) <= b and not a;
    layer5_outputs(7696) <= not b;
    layer5_outputs(7697) <= a xor b;
    layer5_outputs(7698) <= a and not b;
    layer5_outputs(7699) <= not b;
    layer5_outputs(7700) <= b;
    layer5_outputs(7701) <= not a;
    layer5_outputs(7702) <= b and not a;
    layer5_outputs(7703) <= not (a or b);
    layer5_outputs(7704) <= not (a and b);
    layer5_outputs(7705) <= not b;
    layer5_outputs(7706) <= not b;
    layer5_outputs(7707) <= not a;
    layer5_outputs(7708) <= b;
    layer5_outputs(7709) <= a;
    layer5_outputs(7710) <= a xor b;
    layer5_outputs(7711) <= not b or a;
    layer5_outputs(7712) <= not b;
    layer5_outputs(7713) <= a or b;
    layer5_outputs(7714) <= a xor b;
    layer5_outputs(7715) <= not a;
    layer5_outputs(7716) <= b;
    layer5_outputs(7717) <= b and not a;
    layer5_outputs(7718) <= not (a and b);
    layer5_outputs(7719) <= b;
    layer5_outputs(7720) <= not b or a;
    layer5_outputs(7721) <= a xor b;
    layer5_outputs(7722) <= b;
    layer5_outputs(7723) <= not a or b;
    layer5_outputs(7724) <= not b;
    layer5_outputs(7725) <= not a;
    layer5_outputs(7726) <= not b or a;
    layer5_outputs(7727) <= a and not b;
    layer5_outputs(7728) <= not (a and b);
    layer5_outputs(7729) <= not b;
    layer5_outputs(7730) <= a or b;
    layer5_outputs(7731) <= a xor b;
    layer5_outputs(7732) <= not a;
    layer5_outputs(7733) <= '0';
    layer5_outputs(7734) <= b;
    layer5_outputs(7735) <= not a;
    layer5_outputs(7736) <= a or b;
    layer5_outputs(7737) <= '0';
    layer5_outputs(7738) <= not (a and b);
    layer5_outputs(7739) <= a xor b;
    layer5_outputs(7740) <= not a;
    layer5_outputs(7741) <= a xor b;
    layer5_outputs(7742) <= b;
    layer5_outputs(7743) <= a;
    layer5_outputs(7744) <= a and b;
    layer5_outputs(7745) <= not a or b;
    layer5_outputs(7746) <= not b;
    layer5_outputs(7747) <= not a;
    layer5_outputs(7748) <= not a;
    layer5_outputs(7749) <= not a;
    layer5_outputs(7750) <= not a;
    layer5_outputs(7751) <= a;
    layer5_outputs(7752) <= a or b;
    layer5_outputs(7753) <= not (a or b);
    layer5_outputs(7754) <= b;
    layer5_outputs(7755) <= a;
    layer5_outputs(7756) <= not (a and b);
    layer5_outputs(7757) <= a;
    layer5_outputs(7758) <= not b;
    layer5_outputs(7759) <= not (a xor b);
    layer5_outputs(7760) <= not b;
    layer5_outputs(7761) <= not b or a;
    layer5_outputs(7762) <= '0';
    layer5_outputs(7763) <= b;
    layer5_outputs(7764) <= a or b;
    layer5_outputs(7765) <= b;
    layer5_outputs(7766) <= b;
    layer5_outputs(7767) <= a or b;
    layer5_outputs(7768) <= b;
    layer5_outputs(7769) <= b and not a;
    layer5_outputs(7770) <= a;
    layer5_outputs(7771) <= not b;
    layer5_outputs(7772) <= not b;
    layer5_outputs(7773) <= a;
    layer5_outputs(7774) <= a;
    layer5_outputs(7775) <= b and not a;
    layer5_outputs(7776) <= a or b;
    layer5_outputs(7777) <= a and b;
    layer5_outputs(7778) <= not (a or b);
    layer5_outputs(7779) <= a;
    layer5_outputs(7780) <= not b;
    layer5_outputs(7781) <= not b;
    layer5_outputs(7782) <= not b;
    layer5_outputs(7783) <= not a or b;
    layer5_outputs(7784) <= not (a or b);
    layer5_outputs(7785) <= not b;
    layer5_outputs(7786) <= b;
    layer5_outputs(7787) <= not b;
    layer5_outputs(7788) <= not a;
    layer5_outputs(7789) <= not a;
    layer5_outputs(7790) <= not (a or b);
    layer5_outputs(7791) <= a;
    layer5_outputs(7792) <= b;
    layer5_outputs(7793) <= not (a xor b);
    layer5_outputs(7794) <= not (a or b);
    layer5_outputs(7795) <= not a;
    layer5_outputs(7796) <= b;
    layer5_outputs(7797) <= a or b;
    layer5_outputs(7798) <= not (a or b);
    layer5_outputs(7799) <= b;
    layer5_outputs(7800) <= not b or a;
    layer5_outputs(7801) <= a xor b;
    layer5_outputs(7802) <= '1';
    layer5_outputs(7803) <= a;
    layer5_outputs(7804) <= not (a xor b);
    layer5_outputs(7805) <= not b or a;
    layer5_outputs(7806) <= b;
    layer5_outputs(7807) <= not (a or b);
    layer5_outputs(7808) <= a;
    layer5_outputs(7809) <= a xor b;
    layer5_outputs(7810) <= b;
    layer5_outputs(7811) <= not a;
    layer5_outputs(7812) <= not a;
    layer5_outputs(7813) <= a or b;
    layer5_outputs(7814) <= b;
    layer5_outputs(7815) <= b;
    layer5_outputs(7816) <= not (a xor b);
    layer5_outputs(7817) <= not b or a;
    layer5_outputs(7818) <= not (a xor b);
    layer5_outputs(7819) <= a and not b;
    layer5_outputs(7820) <= b;
    layer5_outputs(7821) <= not a;
    layer5_outputs(7822) <= a xor b;
    layer5_outputs(7823) <= a and not b;
    layer5_outputs(7824) <= a;
    layer5_outputs(7825) <= not a or b;
    layer5_outputs(7826) <= not b or a;
    layer5_outputs(7827) <= b;
    layer5_outputs(7828) <= not a;
    layer5_outputs(7829) <= b;
    layer5_outputs(7830) <= b;
    layer5_outputs(7831) <= not (a and b);
    layer5_outputs(7832) <= b;
    layer5_outputs(7833) <= not (a or b);
    layer5_outputs(7834) <= not a or b;
    layer5_outputs(7835) <= not b or a;
    layer5_outputs(7836) <= not a;
    layer5_outputs(7837) <= not (a xor b);
    layer5_outputs(7838) <= a xor b;
    layer5_outputs(7839) <= a;
    layer5_outputs(7840) <= not a;
    layer5_outputs(7841) <= not a;
    layer5_outputs(7842) <= not a;
    layer5_outputs(7843) <= b;
    layer5_outputs(7844) <= not a;
    layer5_outputs(7845) <= not a;
    layer5_outputs(7846) <= not (a xor b);
    layer5_outputs(7847) <= not a;
    layer5_outputs(7848) <= a;
    layer5_outputs(7849) <= b;
    layer5_outputs(7850) <= not a;
    layer5_outputs(7851) <= '0';
    layer5_outputs(7852) <= b and not a;
    layer5_outputs(7853) <= a;
    layer5_outputs(7854) <= not (a xor b);
    layer5_outputs(7855) <= a and b;
    layer5_outputs(7856) <= b;
    layer5_outputs(7857) <= not a;
    layer5_outputs(7858) <= not (a or b);
    layer5_outputs(7859) <= not a or b;
    layer5_outputs(7860) <= a;
    layer5_outputs(7861) <= b;
    layer5_outputs(7862) <= not b;
    layer5_outputs(7863) <= a xor b;
    layer5_outputs(7864) <= '0';
    layer5_outputs(7865) <= a;
    layer5_outputs(7866) <= a or b;
    layer5_outputs(7867) <= a and not b;
    layer5_outputs(7868) <= b and not a;
    layer5_outputs(7869) <= not a or b;
    layer5_outputs(7870) <= not b or a;
    layer5_outputs(7871) <= b;
    layer5_outputs(7872) <= not a;
    layer5_outputs(7873) <= b;
    layer5_outputs(7874) <= not b or a;
    layer5_outputs(7875) <= not (a and b);
    layer5_outputs(7876) <= not (a or b);
    layer5_outputs(7877) <= not a;
    layer5_outputs(7878) <= b;
    layer5_outputs(7879) <= not b or a;
    layer5_outputs(7880) <= a xor b;
    layer5_outputs(7881) <= a xor b;
    layer5_outputs(7882) <= a and b;
    layer5_outputs(7883) <= not a;
    layer5_outputs(7884) <= not (a or b);
    layer5_outputs(7885) <= not a;
    layer5_outputs(7886) <= not a;
    layer5_outputs(7887) <= not a;
    layer5_outputs(7888) <= b;
    layer5_outputs(7889) <= not (a xor b);
    layer5_outputs(7890) <= b;
    layer5_outputs(7891) <= not b or a;
    layer5_outputs(7892) <= not b;
    layer5_outputs(7893) <= b;
    layer5_outputs(7894) <= not b;
    layer5_outputs(7895) <= not a;
    layer5_outputs(7896) <= not (a xor b);
    layer5_outputs(7897) <= a;
    layer5_outputs(7898) <= a;
    layer5_outputs(7899) <= b and not a;
    layer5_outputs(7900) <= not (a and b);
    layer5_outputs(7901) <= b;
    layer5_outputs(7902) <= a xor b;
    layer5_outputs(7903) <= not (a and b);
    layer5_outputs(7904) <= a xor b;
    layer5_outputs(7905) <= b and not a;
    layer5_outputs(7906) <= a;
    layer5_outputs(7907) <= not a;
    layer5_outputs(7908) <= a or b;
    layer5_outputs(7909) <= not b;
    layer5_outputs(7910) <= a xor b;
    layer5_outputs(7911) <= not a;
    layer5_outputs(7912) <= not (a xor b);
    layer5_outputs(7913) <= not (a xor b);
    layer5_outputs(7914) <= '1';
    layer5_outputs(7915) <= not a;
    layer5_outputs(7916) <= a;
    layer5_outputs(7917) <= a or b;
    layer5_outputs(7918) <= a xor b;
    layer5_outputs(7919) <= a;
    layer5_outputs(7920) <= a xor b;
    layer5_outputs(7921) <= b;
    layer5_outputs(7922) <= b;
    layer5_outputs(7923) <= not (a or b);
    layer5_outputs(7924) <= not a;
    layer5_outputs(7925) <= not a;
    layer5_outputs(7926) <= a;
    layer5_outputs(7927) <= not b or a;
    layer5_outputs(7928) <= not (a xor b);
    layer5_outputs(7929) <= a xor b;
    layer5_outputs(7930) <= not (a xor b);
    layer5_outputs(7931) <= not (a or b);
    layer5_outputs(7932) <= not a;
    layer5_outputs(7933) <= '0';
    layer5_outputs(7934) <= b and not a;
    layer5_outputs(7935) <= not a;
    layer5_outputs(7936) <= not (a and b);
    layer5_outputs(7937) <= a xor b;
    layer5_outputs(7938) <= not b or a;
    layer5_outputs(7939) <= a or b;
    layer5_outputs(7940) <= not (a or b);
    layer5_outputs(7941) <= not (a or b);
    layer5_outputs(7942) <= b;
    layer5_outputs(7943) <= not a or b;
    layer5_outputs(7944) <= a and not b;
    layer5_outputs(7945) <= a and b;
    layer5_outputs(7946) <= a;
    layer5_outputs(7947) <= not b or a;
    layer5_outputs(7948) <= not (a xor b);
    layer5_outputs(7949) <= not b;
    layer5_outputs(7950) <= not (a or b);
    layer5_outputs(7951) <= a and b;
    layer5_outputs(7952) <= a xor b;
    layer5_outputs(7953) <= '1';
    layer5_outputs(7954) <= a;
    layer5_outputs(7955) <= not (a and b);
    layer5_outputs(7956) <= a;
    layer5_outputs(7957) <= a and b;
    layer5_outputs(7958) <= not a;
    layer5_outputs(7959) <= not (a or b);
    layer5_outputs(7960) <= a and not b;
    layer5_outputs(7961) <= a;
    layer5_outputs(7962) <= a;
    layer5_outputs(7963) <= not (a or b);
    layer5_outputs(7964) <= a;
    layer5_outputs(7965) <= not a;
    layer5_outputs(7966) <= not (a or b);
    layer5_outputs(7967) <= a xor b;
    layer5_outputs(7968) <= not b;
    layer5_outputs(7969) <= not b;
    layer5_outputs(7970) <= a and not b;
    layer5_outputs(7971) <= b;
    layer5_outputs(7972) <= a;
    layer5_outputs(7973) <= b and not a;
    layer5_outputs(7974) <= b and not a;
    layer5_outputs(7975) <= not (a and b);
    layer5_outputs(7976) <= not a;
    layer5_outputs(7977) <= not b;
    layer5_outputs(7978) <= not b or a;
    layer5_outputs(7979) <= not (a xor b);
    layer5_outputs(7980) <= b and not a;
    layer5_outputs(7981) <= a;
    layer5_outputs(7982) <= not b;
    layer5_outputs(7983) <= a;
    layer5_outputs(7984) <= not (a or b);
    layer5_outputs(7985) <= not a;
    layer5_outputs(7986) <= a and not b;
    layer5_outputs(7987) <= not b or a;
    layer5_outputs(7988) <= a and b;
    layer5_outputs(7989) <= not (a xor b);
    layer5_outputs(7990) <= a or b;
    layer5_outputs(7991) <= b;
    layer5_outputs(7992) <= not (a or b);
    layer5_outputs(7993) <= b;
    layer5_outputs(7994) <= not b;
    layer5_outputs(7995) <= a;
    layer5_outputs(7996) <= a;
    layer5_outputs(7997) <= a;
    layer5_outputs(7998) <= b and not a;
    layer5_outputs(7999) <= a and not b;
    layer5_outputs(8000) <= a;
    layer5_outputs(8001) <= not b;
    layer5_outputs(8002) <= not b;
    layer5_outputs(8003) <= not (a and b);
    layer5_outputs(8004) <= b and not a;
    layer5_outputs(8005) <= not a;
    layer5_outputs(8006) <= a and not b;
    layer5_outputs(8007) <= a and not b;
    layer5_outputs(8008) <= a xor b;
    layer5_outputs(8009) <= b and not a;
    layer5_outputs(8010) <= a and b;
    layer5_outputs(8011) <= a xor b;
    layer5_outputs(8012) <= not b;
    layer5_outputs(8013) <= not a;
    layer5_outputs(8014) <= not (a xor b);
    layer5_outputs(8015) <= a xor b;
    layer5_outputs(8016) <= not a or b;
    layer5_outputs(8017) <= not b;
    layer5_outputs(8018) <= not (a or b);
    layer5_outputs(8019) <= b and not a;
    layer5_outputs(8020) <= not a or b;
    layer5_outputs(8021) <= not a or b;
    layer5_outputs(8022) <= a and not b;
    layer5_outputs(8023) <= a and not b;
    layer5_outputs(8024) <= not (a xor b);
    layer5_outputs(8025) <= a;
    layer5_outputs(8026) <= b and not a;
    layer5_outputs(8027) <= not b;
    layer5_outputs(8028) <= b and not a;
    layer5_outputs(8029) <= a or b;
    layer5_outputs(8030) <= a;
    layer5_outputs(8031) <= not (a xor b);
    layer5_outputs(8032) <= not b or a;
    layer5_outputs(8033) <= a xor b;
    layer5_outputs(8034) <= not (a xor b);
    layer5_outputs(8035) <= not b;
    layer5_outputs(8036) <= a;
    layer5_outputs(8037) <= b and not a;
    layer5_outputs(8038) <= a xor b;
    layer5_outputs(8039) <= not (a and b);
    layer5_outputs(8040) <= a and not b;
    layer5_outputs(8041) <= not b;
    layer5_outputs(8042) <= a and not b;
    layer5_outputs(8043) <= a xor b;
    layer5_outputs(8044) <= a;
    layer5_outputs(8045) <= a or b;
    layer5_outputs(8046) <= a xor b;
    layer5_outputs(8047) <= not a or b;
    layer5_outputs(8048) <= a and not b;
    layer5_outputs(8049) <= a or b;
    layer5_outputs(8050) <= not (a and b);
    layer5_outputs(8051) <= b and not a;
    layer5_outputs(8052) <= not a or b;
    layer5_outputs(8053) <= b and not a;
    layer5_outputs(8054) <= a;
    layer5_outputs(8055) <= not b;
    layer5_outputs(8056) <= not a;
    layer5_outputs(8057) <= not a;
    layer5_outputs(8058) <= not b or a;
    layer5_outputs(8059) <= not (a xor b);
    layer5_outputs(8060) <= not b;
    layer5_outputs(8061) <= a and not b;
    layer5_outputs(8062) <= not (a or b);
    layer5_outputs(8063) <= not b;
    layer5_outputs(8064) <= not a;
    layer5_outputs(8065) <= a and not b;
    layer5_outputs(8066) <= b;
    layer5_outputs(8067) <= not (a xor b);
    layer5_outputs(8068) <= not a;
    layer5_outputs(8069) <= a xor b;
    layer5_outputs(8070) <= not a;
    layer5_outputs(8071) <= not b or a;
    layer5_outputs(8072) <= b;
    layer5_outputs(8073) <= not a;
    layer5_outputs(8074) <= not (a xor b);
    layer5_outputs(8075) <= a or b;
    layer5_outputs(8076) <= a and not b;
    layer5_outputs(8077) <= not b;
    layer5_outputs(8078) <= b;
    layer5_outputs(8079) <= not a;
    layer5_outputs(8080) <= not (a xor b);
    layer5_outputs(8081) <= a xor b;
    layer5_outputs(8082) <= a;
    layer5_outputs(8083) <= not (a or b);
    layer5_outputs(8084) <= '0';
    layer5_outputs(8085) <= not b;
    layer5_outputs(8086) <= b;
    layer5_outputs(8087) <= not (a xor b);
    layer5_outputs(8088) <= not (a or b);
    layer5_outputs(8089) <= a and b;
    layer5_outputs(8090) <= b;
    layer5_outputs(8091) <= not b;
    layer5_outputs(8092) <= not b;
    layer5_outputs(8093) <= not a or b;
    layer5_outputs(8094) <= not (a or b);
    layer5_outputs(8095) <= b;
    layer5_outputs(8096) <= not b;
    layer5_outputs(8097) <= not (a and b);
    layer5_outputs(8098) <= not a;
    layer5_outputs(8099) <= '0';
    layer5_outputs(8100) <= a;
    layer5_outputs(8101) <= a;
    layer5_outputs(8102) <= b;
    layer5_outputs(8103) <= not a;
    layer5_outputs(8104) <= not b;
    layer5_outputs(8105) <= not a;
    layer5_outputs(8106) <= not b;
    layer5_outputs(8107) <= a and not b;
    layer5_outputs(8108) <= a and b;
    layer5_outputs(8109) <= not (a or b);
    layer5_outputs(8110) <= a;
    layer5_outputs(8111) <= not (a and b);
    layer5_outputs(8112) <= not a;
    layer5_outputs(8113) <= a;
    layer5_outputs(8114) <= b;
    layer5_outputs(8115) <= b;
    layer5_outputs(8116) <= not b or a;
    layer5_outputs(8117) <= a and b;
    layer5_outputs(8118) <= not b;
    layer5_outputs(8119) <= a or b;
    layer5_outputs(8120) <= a or b;
    layer5_outputs(8121) <= b;
    layer5_outputs(8122) <= b and not a;
    layer5_outputs(8123) <= not a;
    layer5_outputs(8124) <= a;
    layer5_outputs(8125) <= not a;
    layer5_outputs(8126) <= b;
    layer5_outputs(8127) <= b;
    layer5_outputs(8128) <= b;
    layer5_outputs(8129) <= a and b;
    layer5_outputs(8130) <= not (a xor b);
    layer5_outputs(8131) <= a xor b;
    layer5_outputs(8132) <= a xor b;
    layer5_outputs(8133) <= not b;
    layer5_outputs(8134) <= a;
    layer5_outputs(8135) <= a;
    layer5_outputs(8136) <= not a;
    layer5_outputs(8137) <= a;
    layer5_outputs(8138) <= not (a and b);
    layer5_outputs(8139) <= a xor b;
    layer5_outputs(8140) <= a and not b;
    layer5_outputs(8141) <= not a;
    layer5_outputs(8142) <= not a;
    layer5_outputs(8143) <= not (a and b);
    layer5_outputs(8144) <= a and b;
    layer5_outputs(8145) <= a;
    layer5_outputs(8146) <= not (a and b);
    layer5_outputs(8147) <= not (a xor b);
    layer5_outputs(8148) <= not a;
    layer5_outputs(8149) <= a;
    layer5_outputs(8150) <= a or b;
    layer5_outputs(8151) <= not a;
    layer5_outputs(8152) <= not b or a;
    layer5_outputs(8153) <= a or b;
    layer5_outputs(8154) <= not b;
    layer5_outputs(8155) <= a or b;
    layer5_outputs(8156) <= not (a and b);
    layer5_outputs(8157) <= a xor b;
    layer5_outputs(8158) <= not (a xor b);
    layer5_outputs(8159) <= b and not a;
    layer5_outputs(8160) <= not b;
    layer5_outputs(8161) <= a or b;
    layer5_outputs(8162) <= not a;
    layer5_outputs(8163) <= not a;
    layer5_outputs(8164) <= b;
    layer5_outputs(8165) <= not b;
    layer5_outputs(8166) <= a xor b;
    layer5_outputs(8167) <= not (a xor b);
    layer5_outputs(8168) <= b;
    layer5_outputs(8169) <= not (a xor b);
    layer5_outputs(8170) <= not b;
    layer5_outputs(8171) <= not b;
    layer5_outputs(8172) <= b;
    layer5_outputs(8173) <= not b;
    layer5_outputs(8174) <= a xor b;
    layer5_outputs(8175) <= a or b;
    layer5_outputs(8176) <= not a;
    layer5_outputs(8177) <= a and b;
    layer5_outputs(8178) <= not b;
    layer5_outputs(8179) <= a and not b;
    layer5_outputs(8180) <= not b or a;
    layer5_outputs(8181) <= a;
    layer5_outputs(8182) <= a and not b;
    layer5_outputs(8183) <= a and not b;
    layer5_outputs(8184) <= not b or a;
    layer5_outputs(8185) <= a;
    layer5_outputs(8186) <= not a or b;
    layer5_outputs(8187) <= a xor b;
    layer5_outputs(8188) <= not (a and b);
    layer5_outputs(8189) <= a xor b;
    layer5_outputs(8190) <= a;
    layer5_outputs(8191) <= a or b;
    layer5_outputs(8192) <= a xor b;
    layer5_outputs(8193) <= b and not a;
    layer5_outputs(8194) <= not (a xor b);
    layer5_outputs(8195) <= '1';
    layer5_outputs(8196) <= a or b;
    layer5_outputs(8197) <= not b;
    layer5_outputs(8198) <= b;
    layer5_outputs(8199) <= not a;
    layer5_outputs(8200) <= b;
    layer5_outputs(8201) <= not (a and b);
    layer5_outputs(8202) <= b;
    layer5_outputs(8203) <= b;
    layer5_outputs(8204) <= not b;
    layer5_outputs(8205) <= b and not a;
    layer5_outputs(8206) <= b;
    layer5_outputs(8207) <= '0';
    layer5_outputs(8208) <= b;
    layer5_outputs(8209) <= not a;
    layer5_outputs(8210) <= not b;
    layer5_outputs(8211) <= a;
    layer5_outputs(8212) <= a;
    layer5_outputs(8213) <= not a;
    layer5_outputs(8214) <= b and not a;
    layer5_outputs(8215) <= a;
    layer5_outputs(8216) <= not b;
    layer5_outputs(8217) <= not b or a;
    layer5_outputs(8218) <= b;
    layer5_outputs(8219) <= not (a xor b);
    layer5_outputs(8220) <= a;
    layer5_outputs(8221) <= a xor b;
    layer5_outputs(8222) <= not a;
    layer5_outputs(8223) <= not (a and b);
    layer5_outputs(8224) <= a;
    layer5_outputs(8225) <= b and not a;
    layer5_outputs(8226) <= a;
    layer5_outputs(8227) <= not (a and b);
    layer5_outputs(8228) <= not b;
    layer5_outputs(8229) <= a;
    layer5_outputs(8230) <= a or b;
    layer5_outputs(8231) <= not a;
    layer5_outputs(8232) <= not b or a;
    layer5_outputs(8233) <= not a;
    layer5_outputs(8234) <= a xor b;
    layer5_outputs(8235) <= b;
    layer5_outputs(8236) <= not b;
    layer5_outputs(8237) <= not a;
    layer5_outputs(8238) <= a;
    layer5_outputs(8239) <= not b;
    layer5_outputs(8240) <= '0';
    layer5_outputs(8241) <= a and not b;
    layer5_outputs(8242) <= not b;
    layer5_outputs(8243) <= a;
    layer5_outputs(8244) <= not a;
    layer5_outputs(8245) <= b and not a;
    layer5_outputs(8246) <= not b;
    layer5_outputs(8247) <= not b or a;
    layer5_outputs(8248) <= not b;
    layer5_outputs(8249) <= a;
    layer5_outputs(8250) <= not a;
    layer5_outputs(8251) <= a;
    layer5_outputs(8252) <= not (a and b);
    layer5_outputs(8253) <= not a;
    layer5_outputs(8254) <= not (a or b);
    layer5_outputs(8255) <= not (a or b);
    layer5_outputs(8256) <= '0';
    layer5_outputs(8257) <= a and not b;
    layer5_outputs(8258) <= not a;
    layer5_outputs(8259) <= not a or b;
    layer5_outputs(8260) <= not b;
    layer5_outputs(8261) <= not (a xor b);
    layer5_outputs(8262) <= not b or a;
    layer5_outputs(8263) <= '1';
    layer5_outputs(8264) <= not (a xor b);
    layer5_outputs(8265) <= a and b;
    layer5_outputs(8266) <= not a or b;
    layer5_outputs(8267) <= not a;
    layer5_outputs(8268) <= not (a and b);
    layer5_outputs(8269) <= a and b;
    layer5_outputs(8270) <= not a;
    layer5_outputs(8271) <= not a or b;
    layer5_outputs(8272) <= a xor b;
    layer5_outputs(8273) <= not (a and b);
    layer5_outputs(8274) <= not a;
    layer5_outputs(8275) <= not a;
    layer5_outputs(8276) <= a xor b;
    layer5_outputs(8277) <= not b;
    layer5_outputs(8278) <= a and not b;
    layer5_outputs(8279) <= a;
    layer5_outputs(8280) <= not a or b;
    layer5_outputs(8281) <= not b;
    layer5_outputs(8282) <= not a;
    layer5_outputs(8283) <= not b;
    layer5_outputs(8284) <= not b;
    layer5_outputs(8285) <= not a;
    layer5_outputs(8286) <= not b;
    layer5_outputs(8287) <= b and not a;
    layer5_outputs(8288) <= not a;
    layer5_outputs(8289) <= '0';
    layer5_outputs(8290) <= a;
    layer5_outputs(8291) <= not b or a;
    layer5_outputs(8292) <= not a or b;
    layer5_outputs(8293) <= a and b;
    layer5_outputs(8294) <= a and b;
    layer5_outputs(8295) <= b and not a;
    layer5_outputs(8296) <= not b;
    layer5_outputs(8297) <= not a;
    layer5_outputs(8298) <= not b or a;
    layer5_outputs(8299) <= a xor b;
    layer5_outputs(8300) <= not (a xor b);
    layer5_outputs(8301) <= a;
    layer5_outputs(8302) <= a and not b;
    layer5_outputs(8303) <= a xor b;
    layer5_outputs(8304) <= not a;
    layer5_outputs(8305) <= b;
    layer5_outputs(8306) <= a and b;
    layer5_outputs(8307) <= a;
    layer5_outputs(8308) <= a;
    layer5_outputs(8309) <= not (a and b);
    layer5_outputs(8310) <= a and not b;
    layer5_outputs(8311) <= a;
    layer5_outputs(8312) <= b;
    layer5_outputs(8313) <= not b;
    layer5_outputs(8314) <= not b or a;
    layer5_outputs(8315) <= not a;
    layer5_outputs(8316) <= not a;
    layer5_outputs(8317) <= a and b;
    layer5_outputs(8318) <= not (a xor b);
    layer5_outputs(8319) <= not a;
    layer5_outputs(8320) <= not (a xor b);
    layer5_outputs(8321) <= a xor b;
    layer5_outputs(8322) <= not (a xor b);
    layer5_outputs(8323) <= a or b;
    layer5_outputs(8324) <= not b;
    layer5_outputs(8325) <= a xor b;
    layer5_outputs(8326) <= not (a or b);
    layer5_outputs(8327) <= a xor b;
    layer5_outputs(8328) <= b;
    layer5_outputs(8329) <= a and b;
    layer5_outputs(8330) <= b;
    layer5_outputs(8331) <= not a or b;
    layer5_outputs(8332) <= a or b;
    layer5_outputs(8333) <= not b;
    layer5_outputs(8334) <= b;
    layer5_outputs(8335) <= a or b;
    layer5_outputs(8336) <= a;
    layer5_outputs(8337) <= not (a xor b);
    layer5_outputs(8338) <= a or b;
    layer5_outputs(8339) <= not b or a;
    layer5_outputs(8340) <= a and b;
    layer5_outputs(8341) <= a;
    layer5_outputs(8342) <= a xor b;
    layer5_outputs(8343) <= b;
    layer5_outputs(8344) <= not (a xor b);
    layer5_outputs(8345) <= a;
    layer5_outputs(8346) <= '1';
    layer5_outputs(8347) <= not a or b;
    layer5_outputs(8348) <= a;
    layer5_outputs(8349) <= not b or a;
    layer5_outputs(8350) <= not a;
    layer5_outputs(8351) <= not (a and b);
    layer5_outputs(8352) <= not b or a;
    layer5_outputs(8353) <= not a or b;
    layer5_outputs(8354) <= a xor b;
    layer5_outputs(8355) <= a xor b;
    layer5_outputs(8356) <= a or b;
    layer5_outputs(8357) <= b;
    layer5_outputs(8358) <= not b or a;
    layer5_outputs(8359) <= not a;
    layer5_outputs(8360) <= not (a xor b);
    layer5_outputs(8361) <= '1';
    layer5_outputs(8362) <= a and not b;
    layer5_outputs(8363) <= not a or b;
    layer5_outputs(8364) <= a or b;
    layer5_outputs(8365) <= a and b;
    layer5_outputs(8366) <= a and not b;
    layer5_outputs(8367) <= not (a or b);
    layer5_outputs(8368) <= '1';
    layer5_outputs(8369) <= not (a or b);
    layer5_outputs(8370) <= not b or a;
    layer5_outputs(8371) <= b and not a;
    layer5_outputs(8372) <= not b;
    layer5_outputs(8373) <= a;
    layer5_outputs(8374) <= not a;
    layer5_outputs(8375) <= not (a xor b);
    layer5_outputs(8376) <= not (a and b);
    layer5_outputs(8377) <= b and not a;
    layer5_outputs(8378) <= not (a xor b);
    layer5_outputs(8379) <= not a;
    layer5_outputs(8380) <= a;
    layer5_outputs(8381) <= b;
    layer5_outputs(8382) <= a and b;
    layer5_outputs(8383) <= not (a xor b);
    layer5_outputs(8384) <= b;
    layer5_outputs(8385) <= b and not a;
    layer5_outputs(8386) <= '1';
    layer5_outputs(8387) <= a;
    layer5_outputs(8388) <= not (a and b);
    layer5_outputs(8389) <= b;
    layer5_outputs(8390) <= not (a and b);
    layer5_outputs(8391) <= a;
    layer5_outputs(8392) <= not b;
    layer5_outputs(8393) <= a;
    layer5_outputs(8394) <= b;
    layer5_outputs(8395) <= a xor b;
    layer5_outputs(8396) <= '1';
    layer5_outputs(8397) <= not b;
    layer5_outputs(8398) <= a xor b;
    layer5_outputs(8399) <= not a;
    layer5_outputs(8400) <= b;
    layer5_outputs(8401) <= not (a and b);
    layer5_outputs(8402) <= a xor b;
    layer5_outputs(8403) <= a xor b;
    layer5_outputs(8404) <= b;
    layer5_outputs(8405) <= a or b;
    layer5_outputs(8406) <= a and b;
    layer5_outputs(8407) <= a;
    layer5_outputs(8408) <= a xor b;
    layer5_outputs(8409) <= not a;
    layer5_outputs(8410) <= b and not a;
    layer5_outputs(8411) <= not (a and b);
    layer5_outputs(8412) <= not a or b;
    layer5_outputs(8413) <= '0';
    layer5_outputs(8414) <= b;
    layer5_outputs(8415) <= a xor b;
    layer5_outputs(8416) <= a;
    layer5_outputs(8417) <= a and b;
    layer5_outputs(8418) <= not b or a;
    layer5_outputs(8419) <= a;
    layer5_outputs(8420) <= not b or a;
    layer5_outputs(8421) <= '1';
    layer5_outputs(8422) <= a;
    layer5_outputs(8423) <= '0';
    layer5_outputs(8424) <= not b;
    layer5_outputs(8425) <= not b or a;
    layer5_outputs(8426) <= a and b;
    layer5_outputs(8427) <= not a or b;
    layer5_outputs(8428) <= b and not a;
    layer5_outputs(8429) <= not a;
    layer5_outputs(8430) <= b;
    layer5_outputs(8431) <= '1';
    layer5_outputs(8432) <= a;
    layer5_outputs(8433) <= b;
    layer5_outputs(8434) <= a xor b;
    layer5_outputs(8435) <= not a;
    layer5_outputs(8436) <= a and b;
    layer5_outputs(8437) <= b;
    layer5_outputs(8438) <= a;
    layer5_outputs(8439) <= not a or b;
    layer5_outputs(8440) <= not a;
    layer5_outputs(8441) <= not b or a;
    layer5_outputs(8442) <= b and not a;
    layer5_outputs(8443) <= b;
    layer5_outputs(8444) <= a or b;
    layer5_outputs(8445) <= not b or a;
    layer5_outputs(8446) <= a;
    layer5_outputs(8447) <= a;
    layer5_outputs(8448) <= b;
    layer5_outputs(8449) <= not (a or b);
    layer5_outputs(8450) <= not b or a;
    layer5_outputs(8451) <= not b;
    layer5_outputs(8452) <= not a;
    layer5_outputs(8453) <= a;
    layer5_outputs(8454) <= not (a xor b);
    layer5_outputs(8455) <= a or b;
    layer5_outputs(8456) <= not (a or b);
    layer5_outputs(8457) <= b;
    layer5_outputs(8458) <= a;
    layer5_outputs(8459) <= not a;
    layer5_outputs(8460) <= not b;
    layer5_outputs(8461) <= a and b;
    layer5_outputs(8462) <= a or b;
    layer5_outputs(8463) <= a;
    layer5_outputs(8464) <= b;
    layer5_outputs(8465) <= a and b;
    layer5_outputs(8466) <= a and not b;
    layer5_outputs(8467) <= a and b;
    layer5_outputs(8468) <= not (a or b);
    layer5_outputs(8469) <= b;
    layer5_outputs(8470) <= not (a xor b);
    layer5_outputs(8471) <= a;
    layer5_outputs(8472) <= a;
    layer5_outputs(8473) <= a or b;
    layer5_outputs(8474) <= not a or b;
    layer5_outputs(8475) <= not b or a;
    layer5_outputs(8476) <= not b or a;
    layer5_outputs(8477) <= b;
    layer5_outputs(8478) <= a and b;
    layer5_outputs(8479) <= not (a or b);
    layer5_outputs(8480) <= not (a or b);
    layer5_outputs(8481) <= not (a xor b);
    layer5_outputs(8482) <= not b;
    layer5_outputs(8483) <= not a or b;
    layer5_outputs(8484) <= a and b;
    layer5_outputs(8485) <= a;
    layer5_outputs(8486) <= a or b;
    layer5_outputs(8487) <= b and not a;
    layer5_outputs(8488) <= b;
    layer5_outputs(8489) <= a and not b;
    layer5_outputs(8490) <= not (a and b);
    layer5_outputs(8491) <= a xor b;
    layer5_outputs(8492) <= a;
    layer5_outputs(8493) <= not (a xor b);
    layer5_outputs(8494) <= not b;
    layer5_outputs(8495) <= b;
    layer5_outputs(8496) <= not (a xor b);
    layer5_outputs(8497) <= not a;
    layer5_outputs(8498) <= b and not a;
    layer5_outputs(8499) <= not (a xor b);
    layer5_outputs(8500) <= a and b;
    layer5_outputs(8501) <= b and not a;
    layer5_outputs(8502) <= a xor b;
    layer5_outputs(8503) <= not (a or b);
    layer5_outputs(8504) <= not b;
    layer5_outputs(8505) <= '0';
    layer5_outputs(8506) <= not b;
    layer5_outputs(8507) <= not a;
    layer5_outputs(8508) <= not a or b;
    layer5_outputs(8509) <= not (a or b);
    layer5_outputs(8510) <= not (a xor b);
    layer5_outputs(8511) <= not b or a;
    layer5_outputs(8512) <= not a or b;
    layer5_outputs(8513) <= a;
    layer5_outputs(8514) <= not a;
    layer5_outputs(8515) <= a xor b;
    layer5_outputs(8516) <= b;
    layer5_outputs(8517) <= b and not a;
    layer5_outputs(8518) <= not b or a;
    layer5_outputs(8519) <= a and not b;
    layer5_outputs(8520) <= not b;
    layer5_outputs(8521) <= not (a xor b);
    layer5_outputs(8522) <= a and not b;
    layer5_outputs(8523) <= a;
    layer5_outputs(8524) <= not (a xor b);
    layer5_outputs(8525) <= not a;
    layer5_outputs(8526) <= a;
    layer5_outputs(8527) <= not (a or b);
    layer5_outputs(8528) <= a and not b;
    layer5_outputs(8529) <= a and not b;
    layer5_outputs(8530) <= b and not a;
    layer5_outputs(8531) <= not a;
    layer5_outputs(8532) <= a xor b;
    layer5_outputs(8533) <= not (a and b);
    layer5_outputs(8534) <= not (a xor b);
    layer5_outputs(8535) <= not b;
    layer5_outputs(8536) <= not a or b;
    layer5_outputs(8537) <= not (a xor b);
    layer5_outputs(8538) <= a;
    layer5_outputs(8539) <= not b;
    layer5_outputs(8540) <= a;
    layer5_outputs(8541) <= a xor b;
    layer5_outputs(8542) <= not b or a;
    layer5_outputs(8543) <= not b;
    layer5_outputs(8544) <= a and not b;
    layer5_outputs(8545) <= not a;
    layer5_outputs(8546) <= a xor b;
    layer5_outputs(8547) <= not b;
    layer5_outputs(8548) <= b and not a;
    layer5_outputs(8549) <= a xor b;
    layer5_outputs(8550) <= b;
    layer5_outputs(8551) <= not (a and b);
    layer5_outputs(8552) <= not b;
    layer5_outputs(8553) <= not a or b;
    layer5_outputs(8554) <= a xor b;
    layer5_outputs(8555) <= not b;
    layer5_outputs(8556) <= a xor b;
    layer5_outputs(8557) <= a or b;
    layer5_outputs(8558) <= not (a xor b);
    layer5_outputs(8559) <= b;
    layer5_outputs(8560) <= a or b;
    layer5_outputs(8561) <= not (a or b);
    layer5_outputs(8562) <= a and b;
    layer5_outputs(8563) <= '0';
    layer5_outputs(8564) <= not b or a;
    layer5_outputs(8565) <= not (a and b);
    layer5_outputs(8566) <= not a or b;
    layer5_outputs(8567) <= not b;
    layer5_outputs(8568) <= not (a xor b);
    layer5_outputs(8569) <= a and not b;
    layer5_outputs(8570) <= b;
    layer5_outputs(8571) <= a;
    layer5_outputs(8572) <= a or b;
    layer5_outputs(8573) <= '0';
    layer5_outputs(8574) <= a and not b;
    layer5_outputs(8575) <= b;
    layer5_outputs(8576) <= not (a xor b);
    layer5_outputs(8577) <= not (a xor b);
    layer5_outputs(8578) <= a xor b;
    layer5_outputs(8579) <= a;
    layer5_outputs(8580) <= a xor b;
    layer5_outputs(8581) <= a or b;
    layer5_outputs(8582) <= not a;
    layer5_outputs(8583) <= a xor b;
    layer5_outputs(8584) <= not b;
    layer5_outputs(8585) <= not b;
    layer5_outputs(8586) <= not a;
    layer5_outputs(8587) <= not (a xor b);
    layer5_outputs(8588) <= not (a xor b);
    layer5_outputs(8589) <= a and b;
    layer5_outputs(8590) <= not (a and b);
    layer5_outputs(8591) <= not b or a;
    layer5_outputs(8592) <= not a;
    layer5_outputs(8593) <= a or b;
    layer5_outputs(8594) <= not b;
    layer5_outputs(8595) <= a;
    layer5_outputs(8596) <= not b;
    layer5_outputs(8597) <= not b;
    layer5_outputs(8598) <= b;
    layer5_outputs(8599) <= a;
    layer5_outputs(8600) <= b and not a;
    layer5_outputs(8601) <= not a or b;
    layer5_outputs(8602) <= not a or b;
    layer5_outputs(8603) <= a and not b;
    layer5_outputs(8604) <= not (a and b);
    layer5_outputs(8605) <= not b;
    layer5_outputs(8606) <= not a;
    layer5_outputs(8607) <= not (a xor b);
    layer5_outputs(8608) <= a and not b;
    layer5_outputs(8609) <= a xor b;
    layer5_outputs(8610) <= a and b;
    layer5_outputs(8611) <= b and not a;
    layer5_outputs(8612) <= b and not a;
    layer5_outputs(8613) <= b;
    layer5_outputs(8614) <= b;
    layer5_outputs(8615) <= b and not a;
    layer5_outputs(8616) <= a xor b;
    layer5_outputs(8617) <= not a;
    layer5_outputs(8618) <= b;
    layer5_outputs(8619) <= not a;
    layer5_outputs(8620) <= a and b;
    layer5_outputs(8621) <= a xor b;
    layer5_outputs(8622) <= not b;
    layer5_outputs(8623) <= b and not a;
    layer5_outputs(8624) <= not b;
    layer5_outputs(8625) <= a and b;
    layer5_outputs(8626) <= not a or b;
    layer5_outputs(8627) <= not b or a;
    layer5_outputs(8628) <= b;
    layer5_outputs(8629) <= not a or b;
    layer5_outputs(8630) <= not a or b;
    layer5_outputs(8631) <= a;
    layer5_outputs(8632) <= b;
    layer5_outputs(8633) <= a xor b;
    layer5_outputs(8634) <= not b;
    layer5_outputs(8635) <= not b or a;
    layer5_outputs(8636) <= a;
    layer5_outputs(8637) <= a xor b;
    layer5_outputs(8638) <= not (a and b);
    layer5_outputs(8639) <= not (a or b);
    layer5_outputs(8640) <= a or b;
    layer5_outputs(8641) <= not b;
    layer5_outputs(8642) <= b and not a;
    layer5_outputs(8643) <= a;
    layer5_outputs(8644) <= not b;
    layer5_outputs(8645) <= not a;
    layer5_outputs(8646) <= not a;
    layer5_outputs(8647) <= b;
    layer5_outputs(8648) <= not (a xor b);
    layer5_outputs(8649) <= a;
    layer5_outputs(8650) <= not (a xor b);
    layer5_outputs(8651) <= a;
    layer5_outputs(8652) <= not (a xor b);
    layer5_outputs(8653) <= a xor b;
    layer5_outputs(8654) <= a;
    layer5_outputs(8655) <= b;
    layer5_outputs(8656) <= a;
    layer5_outputs(8657) <= b and not a;
    layer5_outputs(8658) <= a and b;
    layer5_outputs(8659) <= b;
    layer5_outputs(8660) <= not (a and b);
    layer5_outputs(8661) <= a and not b;
    layer5_outputs(8662) <= not a or b;
    layer5_outputs(8663) <= a;
    layer5_outputs(8664) <= not a;
    layer5_outputs(8665) <= '1';
    layer5_outputs(8666) <= a and b;
    layer5_outputs(8667) <= not (a and b);
    layer5_outputs(8668) <= not a or b;
    layer5_outputs(8669) <= not (a and b);
    layer5_outputs(8670) <= a;
    layer5_outputs(8671) <= a or b;
    layer5_outputs(8672) <= not b;
    layer5_outputs(8673) <= a or b;
    layer5_outputs(8674) <= not (a or b);
    layer5_outputs(8675) <= a or b;
    layer5_outputs(8676) <= a xor b;
    layer5_outputs(8677) <= b;
    layer5_outputs(8678) <= a;
    layer5_outputs(8679) <= a;
    layer5_outputs(8680) <= not b;
    layer5_outputs(8681) <= not a or b;
    layer5_outputs(8682) <= not b or a;
    layer5_outputs(8683) <= a xor b;
    layer5_outputs(8684) <= not a or b;
    layer5_outputs(8685) <= a;
    layer5_outputs(8686) <= a xor b;
    layer5_outputs(8687) <= not b;
    layer5_outputs(8688) <= a and not b;
    layer5_outputs(8689) <= a;
    layer5_outputs(8690) <= not (a and b);
    layer5_outputs(8691) <= a or b;
    layer5_outputs(8692) <= not a;
    layer5_outputs(8693) <= not a or b;
    layer5_outputs(8694) <= a;
    layer5_outputs(8695) <= b;
    layer5_outputs(8696) <= b;
    layer5_outputs(8697) <= a or b;
    layer5_outputs(8698) <= a and not b;
    layer5_outputs(8699) <= b;
    layer5_outputs(8700) <= b;
    layer5_outputs(8701) <= b and not a;
    layer5_outputs(8702) <= not a;
    layer5_outputs(8703) <= not (a xor b);
    layer5_outputs(8704) <= b;
    layer5_outputs(8705) <= not a;
    layer5_outputs(8706) <= b;
    layer5_outputs(8707) <= not (a xor b);
    layer5_outputs(8708) <= not b;
    layer5_outputs(8709) <= a xor b;
    layer5_outputs(8710) <= not b;
    layer5_outputs(8711) <= not a;
    layer5_outputs(8712) <= a;
    layer5_outputs(8713) <= a xor b;
    layer5_outputs(8714) <= b;
    layer5_outputs(8715) <= a;
    layer5_outputs(8716) <= not a;
    layer5_outputs(8717) <= not a;
    layer5_outputs(8718) <= a and not b;
    layer5_outputs(8719) <= not b;
    layer5_outputs(8720) <= not (a or b);
    layer5_outputs(8721) <= b;
    layer5_outputs(8722) <= a xor b;
    layer5_outputs(8723) <= not b or a;
    layer5_outputs(8724) <= a;
    layer5_outputs(8725) <= a or b;
    layer5_outputs(8726) <= not (a or b);
    layer5_outputs(8727) <= a xor b;
    layer5_outputs(8728) <= not (a and b);
    layer5_outputs(8729) <= a;
    layer5_outputs(8730) <= a;
    layer5_outputs(8731) <= not a;
    layer5_outputs(8732) <= a xor b;
    layer5_outputs(8733) <= a;
    layer5_outputs(8734) <= a and b;
    layer5_outputs(8735) <= b;
    layer5_outputs(8736) <= not a;
    layer5_outputs(8737) <= a and b;
    layer5_outputs(8738) <= not b;
    layer5_outputs(8739) <= not (a xor b);
    layer5_outputs(8740) <= a;
    layer5_outputs(8741) <= a;
    layer5_outputs(8742) <= b;
    layer5_outputs(8743) <= '0';
    layer5_outputs(8744) <= a xor b;
    layer5_outputs(8745) <= a;
    layer5_outputs(8746) <= a;
    layer5_outputs(8747) <= not b;
    layer5_outputs(8748) <= not b or a;
    layer5_outputs(8749) <= b;
    layer5_outputs(8750) <= a;
    layer5_outputs(8751) <= b and not a;
    layer5_outputs(8752) <= not (a or b);
    layer5_outputs(8753) <= not (a and b);
    layer5_outputs(8754) <= a and b;
    layer5_outputs(8755) <= a;
    layer5_outputs(8756) <= not a or b;
    layer5_outputs(8757) <= a;
    layer5_outputs(8758) <= b;
    layer5_outputs(8759) <= not (a xor b);
    layer5_outputs(8760) <= a or b;
    layer5_outputs(8761) <= not b or a;
    layer5_outputs(8762) <= a;
    layer5_outputs(8763) <= not b;
    layer5_outputs(8764) <= not b;
    layer5_outputs(8765) <= not b;
    layer5_outputs(8766) <= a or b;
    layer5_outputs(8767) <= not (a or b);
    layer5_outputs(8768) <= not a;
    layer5_outputs(8769) <= a and not b;
    layer5_outputs(8770) <= b;
    layer5_outputs(8771) <= not (a xor b);
    layer5_outputs(8772) <= not b or a;
    layer5_outputs(8773) <= b;
    layer5_outputs(8774) <= a and b;
    layer5_outputs(8775) <= a and not b;
    layer5_outputs(8776) <= b and not a;
    layer5_outputs(8777) <= not (a xor b);
    layer5_outputs(8778) <= a and not b;
    layer5_outputs(8779) <= b;
    layer5_outputs(8780) <= b and not a;
    layer5_outputs(8781) <= not (a xor b);
    layer5_outputs(8782) <= '0';
    layer5_outputs(8783) <= a;
    layer5_outputs(8784) <= not (a xor b);
    layer5_outputs(8785) <= not (a and b);
    layer5_outputs(8786) <= not (a and b);
    layer5_outputs(8787) <= not a or b;
    layer5_outputs(8788) <= not a or b;
    layer5_outputs(8789) <= not (a and b);
    layer5_outputs(8790) <= not a or b;
    layer5_outputs(8791) <= a;
    layer5_outputs(8792) <= a xor b;
    layer5_outputs(8793) <= a;
    layer5_outputs(8794) <= not b or a;
    layer5_outputs(8795) <= not (a and b);
    layer5_outputs(8796) <= not (a and b);
    layer5_outputs(8797) <= not (a or b);
    layer5_outputs(8798) <= '0';
    layer5_outputs(8799) <= not a or b;
    layer5_outputs(8800) <= a;
    layer5_outputs(8801) <= '1';
    layer5_outputs(8802) <= a;
    layer5_outputs(8803) <= a and b;
    layer5_outputs(8804) <= a;
    layer5_outputs(8805) <= a;
    layer5_outputs(8806) <= not (a or b);
    layer5_outputs(8807) <= not a;
    layer5_outputs(8808) <= not a;
    layer5_outputs(8809) <= not (a xor b);
    layer5_outputs(8810) <= '0';
    layer5_outputs(8811) <= a;
    layer5_outputs(8812) <= not b;
    layer5_outputs(8813) <= a xor b;
    layer5_outputs(8814) <= b;
    layer5_outputs(8815) <= not a;
    layer5_outputs(8816) <= a and b;
    layer5_outputs(8817) <= not b;
    layer5_outputs(8818) <= not (a and b);
    layer5_outputs(8819) <= not (a or b);
    layer5_outputs(8820) <= not b or a;
    layer5_outputs(8821) <= not a;
    layer5_outputs(8822) <= a and not b;
    layer5_outputs(8823) <= a;
    layer5_outputs(8824) <= not a or b;
    layer5_outputs(8825) <= a and not b;
    layer5_outputs(8826) <= not b or a;
    layer5_outputs(8827) <= not (a and b);
    layer5_outputs(8828) <= a;
    layer5_outputs(8829) <= a and b;
    layer5_outputs(8830) <= not b;
    layer5_outputs(8831) <= a or b;
    layer5_outputs(8832) <= a and b;
    layer5_outputs(8833) <= not b;
    layer5_outputs(8834) <= a and not b;
    layer5_outputs(8835) <= a;
    layer5_outputs(8836) <= not (a xor b);
    layer5_outputs(8837) <= a;
    layer5_outputs(8838) <= a;
    layer5_outputs(8839) <= a;
    layer5_outputs(8840) <= a;
    layer5_outputs(8841) <= not b;
    layer5_outputs(8842) <= a or b;
    layer5_outputs(8843) <= a;
    layer5_outputs(8844) <= b;
    layer5_outputs(8845) <= b;
    layer5_outputs(8846) <= not b;
    layer5_outputs(8847) <= a xor b;
    layer5_outputs(8848) <= not (a and b);
    layer5_outputs(8849) <= a;
    layer5_outputs(8850) <= b;
    layer5_outputs(8851) <= not (a or b);
    layer5_outputs(8852) <= not a;
    layer5_outputs(8853) <= b;
    layer5_outputs(8854) <= b and not a;
    layer5_outputs(8855) <= a and b;
    layer5_outputs(8856) <= not (a xor b);
    layer5_outputs(8857) <= not a;
    layer5_outputs(8858) <= a and b;
    layer5_outputs(8859) <= not (a xor b);
    layer5_outputs(8860) <= a;
    layer5_outputs(8861) <= b;
    layer5_outputs(8862) <= a;
    layer5_outputs(8863) <= not (a xor b);
    layer5_outputs(8864) <= not a;
    layer5_outputs(8865) <= not a;
    layer5_outputs(8866) <= b;
    layer5_outputs(8867) <= not b;
    layer5_outputs(8868) <= a xor b;
    layer5_outputs(8869) <= not a;
    layer5_outputs(8870) <= a;
    layer5_outputs(8871) <= not (a or b);
    layer5_outputs(8872) <= a and b;
    layer5_outputs(8873) <= not a or b;
    layer5_outputs(8874) <= b;
    layer5_outputs(8875) <= a or b;
    layer5_outputs(8876) <= a;
    layer5_outputs(8877) <= a and b;
    layer5_outputs(8878) <= b;
    layer5_outputs(8879) <= b and not a;
    layer5_outputs(8880) <= a or b;
    layer5_outputs(8881) <= b;
    layer5_outputs(8882) <= not (a xor b);
    layer5_outputs(8883) <= a;
    layer5_outputs(8884) <= b;
    layer5_outputs(8885) <= b;
    layer5_outputs(8886) <= not a;
    layer5_outputs(8887) <= not b;
    layer5_outputs(8888) <= a and not b;
    layer5_outputs(8889) <= not (a and b);
    layer5_outputs(8890) <= '0';
    layer5_outputs(8891) <= b;
    layer5_outputs(8892) <= not a;
    layer5_outputs(8893) <= b and not a;
    layer5_outputs(8894) <= not b;
    layer5_outputs(8895) <= not a;
    layer5_outputs(8896) <= a;
    layer5_outputs(8897) <= a;
    layer5_outputs(8898) <= not a or b;
    layer5_outputs(8899) <= not b;
    layer5_outputs(8900) <= not (a and b);
    layer5_outputs(8901) <= a and b;
    layer5_outputs(8902) <= not a;
    layer5_outputs(8903) <= a or b;
    layer5_outputs(8904) <= a or b;
    layer5_outputs(8905) <= not (a xor b);
    layer5_outputs(8906) <= a;
    layer5_outputs(8907) <= not (a xor b);
    layer5_outputs(8908) <= '1';
    layer5_outputs(8909) <= a;
    layer5_outputs(8910) <= a xor b;
    layer5_outputs(8911) <= not a;
    layer5_outputs(8912) <= a or b;
    layer5_outputs(8913) <= not a;
    layer5_outputs(8914) <= not (a or b);
    layer5_outputs(8915) <= a;
    layer5_outputs(8916) <= a or b;
    layer5_outputs(8917) <= b and not a;
    layer5_outputs(8918) <= a;
    layer5_outputs(8919) <= a;
    layer5_outputs(8920) <= not (a or b);
    layer5_outputs(8921) <= not b;
    layer5_outputs(8922) <= b;
    layer5_outputs(8923) <= a;
    layer5_outputs(8924) <= not b;
    layer5_outputs(8925) <= not b;
    layer5_outputs(8926) <= a xor b;
    layer5_outputs(8927) <= a;
    layer5_outputs(8928) <= b and not a;
    layer5_outputs(8929) <= not (a xor b);
    layer5_outputs(8930) <= not (a xor b);
    layer5_outputs(8931) <= a and not b;
    layer5_outputs(8932) <= b and not a;
    layer5_outputs(8933) <= b;
    layer5_outputs(8934) <= a and not b;
    layer5_outputs(8935) <= a;
    layer5_outputs(8936) <= not b or a;
    layer5_outputs(8937) <= a or b;
    layer5_outputs(8938) <= a;
    layer5_outputs(8939) <= a or b;
    layer5_outputs(8940) <= a xor b;
    layer5_outputs(8941) <= not a;
    layer5_outputs(8942) <= a or b;
    layer5_outputs(8943) <= not (a and b);
    layer5_outputs(8944) <= not (a and b);
    layer5_outputs(8945) <= a and b;
    layer5_outputs(8946) <= not b;
    layer5_outputs(8947) <= a or b;
    layer5_outputs(8948) <= not (a xor b);
    layer5_outputs(8949) <= a xor b;
    layer5_outputs(8950) <= not a;
    layer5_outputs(8951) <= not b or a;
    layer5_outputs(8952) <= not b;
    layer5_outputs(8953) <= not a or b;
    layer5_outputs(8954) <= not (a or b);
    layer5_outputs(8955) <= b;
    layer5_outputs(8956) <= not (a and b);
    layer5_outputs(8957) <= not a;
    layer5_outputs(8958) <= not a;
    layer5_outputs(8959) <= b and not a;
    layer5_outputs(8960) <= a or b;
    layer5_outputs(8961) <= not (a xor b);
    layer5_outputs(8962) <= a;
    layer5_outputs(8963) <= a and not b;
    layer5_outputs(8964) <= not b or a;
    layer5_outputs(8965) <= not (a and b);
    layer5_outputs(8966) <= not a;
    layer5_outputs(8967) <= a or b;
    layer5_outputs(8968) <= a xor b;
    layer5_outputs(8969) <= not (a xor b);
    layer5_outputs(8970) <= not (a xor b);
    layer5_outputs(8971) <= a;
    layer5_outputs(8972) <= not (a xor b);
    layer5_outputs(8973) <= a and b;
    layer5_outputs(8974) <= a and not b;
    layer5_outputs(8975) <= a xor b;
    layer5_outputs(8976) <= not b;
    layer5_outputs(8977) <= not b;
    layer5_outputs(8978) <= a;
    layer5_outputs(8979) <= not a or b;
    layer5_outputs(8980) <= b;
    layer5_outputs(8981) <= not a;
    layer5_outputs(8982) <= a or b;
    layer5_outputs(8983) <= b and not a;
    layer5_outputs(8984) <= not b or a;
    layer5_outputs(8985) <= b and not a;
    layer5_outputs(8986) <= b;
    layer5_outputs(8987) <= a;
    layer5_outputs(8988) <= not b;
    layer5_outputs(8989) <= b;
    layer5_outputs(8990) <= not a or b;
    layer5_outputs(8991) <= a;
    layer5_outputs(8992) <= a;
    layer5_outputs(8993) <= b;
    layer5_outputs(8994) <= not (a xor b);
    layer5_outputs(8995) <= b;
    layer5_outputs(8996) <= a and b;
    layer5_outputs(8997) <= not (a and b);
    layer5_outputs(8998) <= b;
    layer5_outputs(8999) <= not b;
    layer5_outputs(9000) <= not (a and b);
    layer5_outputs(9001) <= not (a xor b);
    layer5_outputs(9002) <= not a;
    layer5_outputs(9003) <= not b;
    layer5_outputs(9004) <= not b;
    layer5_outputs(9005) <= a and not b;
    layer5_outputs(9006) <= not b;
    layer5_outputs(9007) <= a;
    layer5_outputs(9008) <= a;
    layer5_outputs(9009) <= not b;
    layer5_outputs(9010) <= not a or b;
    layer5_outputs(9011) <= a or b;
    layer5_outputs(9012) <= b;
    layer5_outputs(9013) <= b;
    layer5_outputs(9014) <= b;
    layer5_outputs(9015) <= b;
    layer5_outputs(9016) <= not (a xor b);
    layer5_outputs(9017) <= a or b;
    layer5_outputs(9018) <= not (a and b);
    layer5_outputs(9019) <= a and b;
    layer5_outputs(9020) <= not a or b;
    layer5_outputs(9021) <= not a or b;
    layer5_outputs(9022) <= not (a xor b);
    layer5_outputs(9023) <= a;
    layer5_outputs(9024) <= a;
    layer5_outputs(9025) <= not a;
    layer5_outputs(9026) <= a and b;
    layer5_outputs(9027) <= not a;
    layer5_outputs(9028) <= a xor b;
    layer5_outputs(9029) <= a;
    layer5_outputs(9030) <= a or b;
    layer5_outputs(9031) <= a and not b;
    layer5_outputs(9032) <= b and not a;
    layer5_outputs(9033) <= not (a xor b);
    layer5_outputs(9034) <= a and b;
    layer5_outputs(9035) <= a and b;
    layer5_outputs(9036) <= b;
    layer5_outputs(9037) <= a;
    layer5_outputs(9038) <= not b;
    layer5_outputs(9039) <= not (a xor b);
    layer5_outputs(9040) <= not b;
    layer5_outputs(9041) <= a;
    layer5_outputs(9042) <= not (a xor b);
    layer5_outputs(9043) <= not a;
    layer5_outputs(9044) <= b and not a;
    layer5_outputs(9045) <= not a;
    layer5_outputs(9046) <= not b or a;
    layer5_outputs(9047) <= a;
    layer5_outputs(9048) <= not b;
    layer5_outputs(9049) <= not b;
    layer5_outputs(9050) <= not a or b;
    layer5_outputs(9051) <= not b;
    layer5_outputs(9052) <= b and not a;
    layer5_outputs(9053) <= b;
    layer5_outputs(9054) <= not b;
    layer5_outputs(9055) <= not (a or b);
    layer5_outputs(9056) <= not b;
    layer5_outputs(9057) <= not a;
    layer5_outputs(9058) <= not b;
    layer5_outputs(9059) <= not a;
    layer5_outputs(9060) <= a xor b;
    layer5_outputs(9061) <= not (a or b);
    layer5_outputs(9062) <= a;
    layer5_outputs(9063) <= not (a or b);
    layer5_outputs(9064) <= not (a and b);
    layer5_outputs(9065) <= a or b;
    layer5_outputs(9066) <= not b;
    layer5_outputs(9067) <= not (a and b);
    layer5_outputs(9068) <= a xor b;
    layer5_outputs(9069) <= not a or b;
    layer5_outputs(9070) <= not (a and b);
    layer5_outputs(9071) <= not b or a;
    layer5_outputs(9072) <= b;
    layer5_outputs(9073) <= not a;
    layer5_outputs(9074) <= not a;
    layer5_outputs(9075) <= a and not b;
    layer5_outputs(9076) <= not (a or b);
    layer5_outputs(9077) <= not a;
    layer5_outputs(9078) <= not b;
    layer5_outputs(9079) <= not a or b;
    layer5_outputs(9080) <= b;
    layer5_outputs(9081) <= b;
    layer5_outputs(9082) <= not b or a;
    layer5_outputs(9083) <= a xor b;
    layer5_outputs(9084) <= not a;
    layer5_outputs(9085) <= not (a or b);
    layer5_outputs(9086) <= not (a and b);
    layer5_outputs(9087) <= a xor b;
    layer5_outputs(9088) <= not a;
    layer5_outputs(9089) <= a;
    layer5_outputs(9090) <= not b;
    layer5_outputs(9091) <= a xor b;
    layer5_outputs(9092) <= not a;
    layer5_outputs(9093) <= b;
    layer5_outputs(9094) <= a or b;
    layer5_outputs(9095) <= not a;
    layer5_outputs(9096) <= a;
    layer5_outputs(9097) <= b;
    layer5_outputs(9098) <= not (a or b);
    layer5_outputs(9099) <= a;
    layer5_outputs(9100) <= not (a and b);
    layer5_outputs(9101) <= a or b;
    layer5_outputs(9102) <= b and not a;
    layer5_outputs(9103) <= a xor b;
    layer5_outputs(9104) <= a and b;
    layer5_outputs(9105) <= a or b;
    layer5_outputs(9106) <= not (a and b);
    layer5_outputs(9107) <= b and not a;
    layer5_outputs(9108) <= a and b;
    layer5_outputs(9109) <= not b;
    layer5_outputs(9110) <= not b;
    layer5_outputs(9111) <= not b or a;
    layer5_outputs(9112) <= not a or b;
    layer5_outputs(9113) <= a;
    layer5_outputs(9114) <= not (a xor b);
    layer5_outputs(9115) <= not b or a;
    layer5_outputs(9116) <= a and b;
    layer5_outputs(9117) <= a and not b;
    layer5_outputs(9118) <= not (a and b);
    layer5_outputs(9119) <= not a;
    layer5_outputs(9120) <= a;
    layer5_outputs(9121) <= a and b;
    layer5_outputs(9122) <= b;
    layer5_outputs(9123) <= a and not b;
    layer5_outputs(9124) <= '0';
    layer5_outputs(9125) <= a or b;
    layer5_outputs(9126) <= a;
    layer5_outputs(9127) <= a xor b;
    layer5_outputs(9128) <= '1';
    layer5_outputs(9129) <= not a;
    layer5_outputs(9130) <= not a;
    layer5_outputs(9131) <= '0';
    layer5_outputs(9132) <= a xor b;
    layer5_outputs(9133) <= not b or a;
    layer5_outputs(9134) <= not (a xor b);
    layer5_outputs(9135) <= b and not a;
    layer5_outputs(9136) <= a;
    layer5_outputs(9137) <= a;
    layer5_outputs(9138) <= a xor b;
    layer5_outputs(9139) <= b;
    layer5_outputs(9140) <= b;
    layer5_outputs(9141) <= not b or a;
    layer5_outputs(9142) <= not (a xor b);
    layer5_outputs(9143) <= a and b;
    layer5_outputs(9144) <= not (a xor b);
    layer5_outputs(9145) <= not b or a;
    layer5_outputs(9146) <= a and not b;
    layer5_outputs(9147) <= not (a or b);
    layer5_outputs(9148) <= a;
    layer5_outputs(9149) <= not b;
    layer5_outputs(9150) <= b and not a;
    layer5_outputs(9151) <= not (a or b);
    layer5_outputs(9152) <= not a or b;
    layer5_outputs(9153) <= '1';
    layer5_outputs(9154) <= b;
    layer5_outputs(9155) <= not b;
    layer5_outputs(9156) <= not b or a;
    layer5_outputs(9157) <= a and not b;
    layer5_outputs(9158) <= a or b;
    layer5_outputs(9159) <= a or b;
    layer5_outputs(9160) <= not b;
    layer5_outputs(9161) <= not (a and b);
    layer5_outputs(9162) <= a xor b;
    layer5_outputs(9163) <= not (a or b);
    layer5_outputs(9164) <= not b;
    layer5_outputs(9165) <= not (a and b);
    layer5_outputs(9166) <= not (a or b);
    layer5_outputs(9167) <= b and not a;
    layer5_outputs(9168) <= a;
    layer5_outputs(9169) <= not a;
    layer5_outputs(9170) <= b and not a;
    layer5_outputs(9171) <= a;
    layer5_outputs(9172) <= not b;
    layer5_outputs(9173) <= not b;
    layer5_outputs(9174) <= b;
    layer5_outputs(9175) <= '1';
    layer5_outputs(9176) <= a and not b;
    layer5_outputs(9177) <= b;
    layer5_outputs(9178) <= b;
    layer5_outputs(9179) <= not (a or b);
    layer5_outputs(9180) <= a xor b;
    layer5_outputs(9181) <= not a or b;
    layer5_outputs(9182) <= a or b;
    layer5_outputs(9183) <= not (a and b);
    layer5_outputs(9184) <= a xor b;
    layer5_outputs(9185) <= not a;
    layer5_outputs(9186) <= not a;
    layer5_outputs(9187) <= a;
    layer5_outputs(9188) <= a;
    layer5_outputs(9189) <= a or b;
    layer5_outputs(9190) <= a;
    layer5_outputs(9191) <= a xor b;
    layer5_outputs(9192) <= not a or b;
    layer5_outputs(9193) <= not (a or b);
    layer5_outputs(9194) <= not a;
    layer5_outputs(9195) <= not b;
    layer5_outputs(9196) <= not a or b;
    layer5_outputs(9197) <= not (a and b);
    layer5_outputs(9198) <= b;
    layer5_outputs(9199) <= not a or b;
    layer5_outputs(9200) <= not a;
    layer5_outputs(9201) <= not (a and b);
    layer5_outputs(9202) <= a and not b;
    layer5_outputs(9203) <= not b or a;
    layer5_outputs(9204) <= not b;
    layer5_outputs(9205) <= a and not b;
    layer5_outputs(9206) <= a and not b;
    layer5_outputs(9207) <= b;
    layer5_outputs(9208) <= '0';
    layer5_outputs(9209) <= not b or a;
    layer5_outputs(9210) <= not b;
    layer5_outputs(9211) <= a and not b;
    layer5_outputs(9212) <= not a or b;
    layer5_outputs(9213) <= not (a or b);
    layer5_outputs(9214) <= not b;
    layer5_outputs(9215) <= not a;
    layer5_outputs(9216) <= b;
    layer5_outputs(9217) <= a;
    layer5_outputs(9218) <= not a;
    layer5_outputs(9219) <= not a;
    layer5_outputs(9220) <= not (a and b);
    layer5_outputs(9221) <= a xor b;
    layer5_outputs(9222) <= a and not b;
    layer5_outputs(9223) <= not (a xor b);
    layer5_outputs(9224) <= not b or a;
    layer5_outputs(9225) <= not (a xor b);
    layer5_outputs(9226) <= a and not b;
    layer5_outputs(9227) <= not b;
    layer5_outputs(9228) <= not a;
    layer5_outputs(9229) <= not b;
    layer5_outputs(9230) <= a;
    layer5_outputs(9231) <= '0';
    layer5_outputs(9232) <= b;
    layer5_outputs(9233) <= b;
    layer5_outputs(9234) <= not a or b;
    layer5_outputs(9235) <= not b;
    layer5_outputs(9236) <= not a;
    layer5_outputs(9237) <= a or b;
    layer5_outputs(9238) <= not (a xor b);
    layer5_outputs(9239) <= not (a xor b);
    layer5_outputs(9240) <= a and b;
    layer5_outputs(9241) <= not b;
    layer5_outputs(9242) <= not b or a;
    layer5_outputs(9243) <= a;
    layer5_outputs(9244) <= not (a and b);
    layer5_outputs(9245) <= not b;
    layer5_outputs(9246) <= not (a or b);
    layer5_outputs(9247) <= not (a xor b);
    layer5_outputs(9248) <= b;
    layer5_outputs(9249) <= not b;
    layer5_outputs(9250) <= not (a and b);
    layer5_outputs(9251) <= a and b;
    layer5_outputs(9252) <= a and not b;
    layer5_outputs(9253) <= a;
    layer5_outputs(9254) <= a or b;
    layer5_outputs(9255) <= b;
    layer5_outputs(9256) <= not b;
    layer5_outputs(9257) <= not b or a;
    layer5_outputs(9258) <= not a;
    layer5_outputs(9259) <= a xor b;
    layer5_outputs(9260) <= not b;
    layer5_outputs(9261) <= not (a and b);
    layer5_outputs(9262) <= not b;
    layer5_outputs(9263) <= not (a or b);
    layer5_outputs(9264) <= not b or a;
    layer5_outputs(9265) <= not a;
    layer5_outputs(9266) <= a xor b;
    layer5_outputs(9267) <= not (a and b);
    layer5_outputs(9268) <= '0';
    layer5_outputs(9269) <= '0';
    layer5_outputs(9270) <= a;
    layer5_outputs(9271) <= not a;
    layer5_outputs(9272) <= b and not a;
    layer5_outputs(9273) <= a;
    layer5_outputs(9274) <= '0';
    layer5_outputs(9275) <= a;
    layer5_outputs(9276) <= a or b;
    layer5_outputs(9277) <= b and not a;
    layer5_outputs(9278) <= a or b;
    layer5_outputs(9279) <= a;
    layer5_outputs(9280) <= a and not b;
    layer5_outputs(9281) <= not (a xor b);
    layer5_outputs(9282) <= not (a or b);
    layer5_outputs(9283) <= not a or b;
    layer5_outputs(9284) <= b;
    layer5_outputs(9285) <= a xor b;
    layer5_outputs(9286) <= not a;
    layer5_outputs(9287) <= not a;
    layer5_outputs(9288) <= not (a xor b);
    layer5_outputs(9289) <= not b;
    layer5_outputs(9290) <= b and not a;
    layer5_outputs(9291) <= not a;
    layer5_outputs(9292) <= b;
    layer5_outputs(9293) <= a;
    layer5_outputs(9294) <= '0';
    layer5_outputs(9295) <= not b or a;
    layer5_outputs(9296) <= a xor b;
    layer5_outputs(9297) <= a xor b;
    layer5_outputs(9298) <= a;
    layer5_outputs(9299) <= not (a or b);
    layer5_outputs(9300) <= b;
    layer5_outputs(9301) <= not (a xor b);
    layer5_outputs(9302) <= not b;
    layer5_outputs(9303) <= not b;
    layer5_outputs(9304) <= a or b;
    layer5_outputs(9305) <= not b or a;
    layer5_outputs(9306) <= not b or a;
    layer5_outputs(9307) <= a;
    layer5_outputs(9308) <= b and not a;
    layer5_outputs(9309) <= not (a or b);
    layer5_outputs(9310) <= not (a and b);
    layer5_outputs(9311) <= not b;
    layer5_outputs(9312) <= not (a xor b);
    layer5_outputs(9313) <= b and not a;
    layer5_outputs(9314) <= not (a and b);
    layer5_outputs(9315) <= not (a xor b);
    layer5_outputs(9316) <= not b;
    layer5_outputs(9317) <= b;
    layer5_outputs(9318) <= not b;
    layer5_outputs(9319) <= a or b;
    layer5_outputs(9320) <= b;
    layer5_outputs(9321) <= not a or b;
    layer5_outputs(9322) <= a;
    layer5_outputs(9323) <= a xor b;
    layer5_outputs(9324) <= not (a xor b);
    layer5_outputs(9325) <= a;
    layer5_outputs(9326) <= not b;
    layer5_outputs(9327) <= a;
    layer5_outputs(9328) <= not b;
    layer5_outputs(9329) <= a or b;
    layer5_outputs(9330) <= not b or a;
    layer5_outputs(9331) <= not (a and b);
    layer5_outputs(9332) <= a;
    layer5_outputs(9333) <= not (a xor b);
    layer5_outputs(9334) <= a;
    layer5_outputs(9335) <= b;
    layer5_outputs(9336) <= not b;
    layer5_outputs(9337) <= a;
    layer5_outputs(9338) <= not a;
    layer5_outputs(9339) <= not b or a;
    layer5_outputs(9340) <= not b;
    layer5_outputs(9341) <= not a or b;
    layer5_outputs(9342) <= not (a and b);
    layer5_outputs(9343) <= not a;
    layer5_outputs(9344) <= not (a xor b);
    layer5_outputs(9345) <= a;
    layer5_outputs(9346) <= a or b;
    layer5_outputs(9347) <= b and not a;
    layer5_outputs(9348) <= a and not b;
    layer5_outputs(9349) <= b;
    layer5_outputs(9350) <= a xor b;
    layer5_outputs(9351) <= a;
    layer5_outputs(9352) <= b;
    layer5_outputs(9353) <= not a;
    layer5_outputs(9354) <= b;
    layer5_outputs(9355) <= a and b;
    layer5_outputs(9356) <= a;
    layer5_outputs(9357) <= b and not a;
    layer5_outputs(9358) <= not a;
    layer5_outputs(9359) <= not b or a;
    layer5_outputs(9360) <= a;
    layer5_outputs(9361) <= '1';
    layer5_outputs(9362) <= b and not a;
    layer5_outputs(9363) <= b;
    layer5_outputs(9364) <= b;
    layer5_outputs(9365) <= not a;
    layer5_outputs(9366) <= not (a or b);
    layer5_outputs(9367) <= not a;
    layer5_outputs(9368) <= not (a xor b);
    layer5_outputs(9369) <= b;
    layer5_outputs(9370) <= not a or b;
    layer5_outputs(9371) <= b;
    layer5_outputs(9372) <= a and not b;
    layer5_outputs(9373) <= a;
    layer5_outputs(9374) <= a;
    layer5_outputs(9375) <= b and not a;
    layer5_outputs(9376) <= a and b;
    layer5_outputs(9377) <= not (a and b);
    layer5_outputs(9378) <= not (a and b);
    layer5_outputs(9379) <= b and not a;
    layer5_outputs(9380) <= a and not b;
    layer5_outputs(9381) <= b;
    layer5_outputs(9382) <= '0';
    layer5_outputs(9383) <= a;
    layer5_outputs(9384) <= b;
    layer5_outputs(9385) <= not b;
    layer5_outputs(9386) <= a or b;
    layer5_outputs(9387) <= not a;
    layer5_outputs(9388) <= not (a xor b);
    layer5_outputs(9389) <= not b;
    layer5_outputs(9390) <= not (a and b);
    layer5_outputs(9391) <= not (a and b);
    layer5_outputs(9392) <= not (a xor b);
    layer5_outputs(9393) <= not a or b;
    layer5_outputs(9394) <= not b or a;
    layer5_outputs(9395) <= a and not b;
    layer5_outputs(9396) <= not a;
    layer5_outputs(9397) <= not (a xor b);
    layer5_outputs(9398) <= a;
    layer5_outputs(9399) <= not (a and b);
    layer5_outputs(9400) <= b;
    layer5_outputs(9401) <= b and not a;
    layer5_outputs(9402) <= not b;
    layer5_outputs(9403) <= not (a or b);
    layer5_outputs(9404) <= not (a or b);
    layer5_outputs(9405) <= a;
    layer5_outputs(9406) <= not (a and b);
    layer5_outputs(9407) <= a and b;
    layer5_outputs(9408) <= a xor b;
    layer5_outputs(9409) <= not a;
    layer5_outputs(9410) <= a and not b;
    layer5_outputs(9411) <= '0';
    layer5_outputs(9412) <= a;
    layer5_outputs(9413) <= not (a or b);
    layer5_outputs(9414) <= a;
    layer5_outputs(9415) <= b and not a;
    layer5_outputs(9416) <= not b;
    layer5_outputs(9417) <= a;
    layer5_outputs(9418) <= not (a or b);
    layer5_outputs(9419) <= not b;
    layer5_outputs(9420) <= a or b;
    layer5_outputs(9421) <= not (a xor b);
    layer5_outputs(9422) <= b;
    layer5_outputs(9423) <= a and not b;
    layer5_outputs(9424) <= b;
    layer5_outputs(9425) <= not a;
    layer5_outputs(9426) <= b and not a;
    layer5_outputs(9427) <= not a;
    layer5_outputs(9428) <= not (a or b);
    layer5_outputs(9429) <= '0';
    layer5_outputs(9430) <= a and b;
    layer5_outputs(9431) <= not a;
    layer5_outputs(9432) <= not a;
    layer5_outputs(9433) <= b and not a;
    layer5_outputs(9434) <= not a;
    layer5_outputs(9435) <= not b or a;
    layer5_outputs(9436) <= b;
    layer5_outputs(9437) <= not b or a;
    layer5_outputs(9438) <= not a;
    layer5_outputs(9439) <= not a or b;
    layer5_outputs(9440) <= not b;
    layer5_outputs(9441) <= not b;
    layer5_outputs(9442) <= not a;
    layer5_outputs(9443) <= b and not a;
    layer5_outputs(9444) <= not (a and b);
    layer5_outputs(9445) <= not b;
    layer5_outputs(9446) <= a;
    layer5_outputs(9447) <= a and b;
    layer5_outputs(9448) <= not (a and b);
    layer5_outputs(9449) <= not a or b;
    layer5_outputs(9450) <= not b or a;
    layer5_outputs(9451) <= b;
    layer5_outputs(9452) <= a and not b;
    layer5_outputs(9453) <= not a;
    layer5_outputs(9454) <= a and not b;
    layer5_outputs(9455) <= not b;
    layer5_outputs(9456) <= a;
    layer5_outputs(9457) <= a xor b;
    layer5_outputs(9458) <= b;
    layer5_outputs(9459) <= not b;
    layer5_outputs(9460) <= a and b;
    layer5_outputs(9461) <= a and b;
    layer5_outputs(9462) <= a or b;
    layer5_outputs(9463) <= not b;
    layer5_outputs(9464) <= b;
    layer5_outputs(9465) <= a xor b;
    layer5_outputs(9466) <= a;
    layer5_outputs(9467) <= a xor b;
    layer5_outputs(9468) <= not a;
    layer5_outputs(9469) <= not (a or b);
    layer5_outputs(9470) <= not b;
    layer5_outputs(9471) <= a;
    layer5_outputs(9472) <= a;
    layer5_outputs(9473) <= b and not a;
    layer5_outputs(9474) <= not (a xor b);
    layer5_outputs(9475) <= not (a and b);
    layer5_outputs(9476) <= not a;
    layer5_outputs(9477) <= not a or b;
    layer5_outputs(9478) <= a xor b;
    layer5_outputs(9479) <= a;
    layer5_outputs(9480) <= not a;
    layer5_outputs(9481) <= not b;
    layer5_outputs(9482) <= a or b;
    layer5_outputs(9483) <= a;
    layer5_outputs(9484) <= not (a xor b);
    layer5_outputs(9485) <= a;
    layer5_outputs(9486) <= a and not b;
    layer5_outputs(9487) <= not b;
    layer5_outputs(9488) <= b;
    layer5_outputs(9489) <= a xor b;
    layer5_outputs(9490) <= not a;
    layer5_outputs(9491) <= not b or a;
    layer5_outputs(9492) <= not b or a;
    layer5_outputs(9493) <= not a;
    layer5_outputs(9494) <= not a;
    layer5_outputs(9495) <= not (a xor b);
    layer5_outputs(9496) <= b;
    layer5_outputs(9497) <= b;
    layer5_outputs(9498) <= a xor b;
    layer5_outputs(9499) <= not (a xor b);
    layer5_outputs(9500) <= not b;
    layer5_outputs(9501) <= not b or a;
    layer5_outputs(9502) <= not a;
    layer5_outputs(9503) <= a and b;
    layer5_outputs(9504) <= not a;
    layer5_outputs(9505) <= a;
    layer5_outputs(9506) <= a xor b;
    layer5_outputs(9507) <= a;
    layer5_outputs(9508) <= b;
    layer5_outputs(9509) <= not b or a;
    layer5_outputs(9510) <= not (a or b);
    layer5_outputs(9511) <= not a;
    layer5_outputs(9512) <= not (a and b);
    layer5_outputs(9513) <= not (a and b);
    layer5_outputs(9514) <= a;
    layer5_outputs(9515) <= not (a or b);
    layer5_outputs(9516) <= not a or b;
    layer5_outputs(9517) <= a xor b;
    layer5_outputs(9518) <= b;
    layer5_outputs(9519) <= not b;
    layer5_outputs(9520) <= not b;
    layer5_outputs(9521) <= not b;
    layer5_outputs(9522) <= a;
    layer5_outputs(9523) <= a or b;
    layer5_outputs(9524) <= not (a or b);
    layer5_outputs(9525) <= not b or a;
    layer5_outputs(9526) <= b;
    layer5_outputs(9527) <= a or b;
    layer5_outputs(9528) <= not b;
    layer5_outputs(9529) <= not (a or b);
    layer5_outputs(9530) <= a;
    layer5_outputs(9531) <= not b;
    layer5_outputs(9532) <= a;
    layer5_outputs(9533) <= a and b;
    layer5_outputs(9534) <= b;
    layer5_outputs(9535) <= b and not a;
    layer5_outputs(9536) <= not b;
    layer5_outputs(9537) <= a;
    layer5_outputs(9538) <= a xor b;
    layer5_outputs(9539) <= a xor b;
    layer5_outputs(9540) <= a xor b;
    layer5_outputs(9541) <= not (a and b);
    layer5_outputs(9542) <= not (a xor b);
    layer5_outputs(9543) <= not a;
    layer5_outputs(9544) <= b;
    layer5_outputs(9545) <= b;
    layer5_outputs(9546) <= not a;
    layer5_outputs(9547) <= not (a or b);
    layer5_outputs(9548) <= not (a and b);
    layer5_outputs(9549) <= not (a xor b);
    layer5_outputs(9550) <= not (a or b);
    layer5_outputs(9551) <= b;
    layer5_outputs(9552) <= not a;
    layer5_outputs(9553) <= b;
    layer5_outputs(9554) <= b;
    layer5_outputs(9555) <= b and not a;
    layer5_outputs(9556) <= a or b;
    layer5_outputs(9557) <= a xor b;
    layer5_outputs(9558) <= '1';
    layer5_outputs(9559) <= not a;
    layer5_outputs(9560) <= not a or b;
    layer5_outputs(9561) <= not b or a;
    layer5_outputs(9562) <= a xor b;
    layer5_outputs(9563) <= a;
    layer5_outputs(9564) <= not a;
    layer5_outputs(9565) <= a and not b;
    layer5_outputs(9566) <= '0';
    layer5_outputs(9567) <= a;
    layer5_outputs(9568) <= a and not b;
    layer5_outputs(9569) <= a;
    layer5_outputs(9570) <= a or b;
    layer5_outputs(9571) <= b;
    layer5_outputs(9572) <= '1';
    layer5_outputs(9573) <= a xor b;
    layer5_outputs(9574) <= not a or b;
    layer5_outputs(9575) <= not a or b;
    layer5_outputs(9576) <= a;
    layer5_outputs(9577) <= not a;
    layer5_outputs(9578) <= not a;
    layer5_outputs(9579) <= a xor b;
    layer5_outputs(9580) <= a;
    layer5_outputs(9581) <= not b or a;
    layer5_outputs(9582) <= not a;
    layer5_outputs(9583) <= not b or a;
    layer5_outputs(9584) <= not (a or b);
    layer5_outputs(9585) <= a xor b;
    layer5_outputs(9586) <= a;
    layer5_outputs(9587) <= not (a or b);
    layer5_outputs(9588) <= a;
    layer5_outputs(9589) <= a or b;
    layer5_outputs(9590) <= b;
    layer5_outputs(9591) <= not (a xor b);
    layer5_outputs(9592) <= not (a xor b);
    layer5_outputs(9593) <= b;
    layer5_outputs(9594) <= not b;
    layer5_outputs(9595) <= a;
    layer5_outputs(9596) <= not b or a;
    layer5_outputs(9597) <= not b;
    layer5_outputs(9598) <= not b;
    layer5_outputs(9599) <= not (a or b);
    layer5_outputs(9600) <= not (a and b);
    layer5_outputs(9601) <= not a;
    layer5_outputs(9602) <= a;
    layer5_outputs(9603) <= not b or a;
    layer5_outputs(9604) <= a or b;
    layer5_outputs(9605) <= not a;
    layer5_outputs(9606) <= a;
    layer5_outputs(9607) <= not a or b;
    layer5_outputs(9608) <= not a;
    layer5_outputs(9609) <= a;
    layer5_outputs(9610) <= a and b;
    layer5_outputs(9611) <= a;
    layer5_outputs(9612) <= a;
    layer5_outputs(9613) <= not (a xor b);
    layer5_outputs(9614) <= not a;
    layer5_outputs(9615) <= a and b;
    layer5_outputs(9616) <= not a;
    layer5_outputs(9617) <= b and not a;
    layer5_outputs(9618) <= a and b;
    layer5_outputs(9619) <= a or b;
    layer5_outputs(9620) <= b;
    layer5_outputs(9621) <= not a;
    layer5_outputs(9622) <= not a;
    layer5_outputs(9623) <= '0';
    layer5_outputs(9624) <= '0';
    layer5_outputs(9625) <= b;
    layer5_outputs(9626) <= '1';
    layer5_outputs(9627) <= b;
    layer5_outputs(9628) <= a xor b;
    layer5_outputs(9629) <= not b;
    layer5_outputs(9630) <= not (a or b);
    layer5_outputs(9631) <= a and not b;
    layer5_outputs(9632) <= not b;
    layer5_outputs(9633) <= not b or a;
    layer5_outputs(9634) <= a;
    layer5_outputs(9635) <= not a;
    layer5_outputs(9636) <= a and b;
    layer5_outputs(9637) <= a;
    layer5_outputs(9638) <= a xor b;
    layer5_outputs(9639) <= not (a xor b);
    layer5_outputs(9640) <= not b;
    layer5_outputs(9641) <= a or b;
    layer5_outputs(9642) <= not a;
    layer5_outputs(9643) <= a and not b;
    layer5_outputs(9644) <= a;
    layer5_outputs(9645) <= not a;
    layer5_outputs(9646) <= b and not a;
    layer5_outputs(9647) <= a and b;
    layer5_outputs(9648) <= b;
    layer5_outputs(9649) <= not (a and b);
    layer5_outputs(9650) <= not b;
    layer5_outputs(9651) <= b;
    layer5_outputs(9652) <= a or b;
    layer5_outputs(9653) <= not (a or b);
    layer5_outputs(9654) <= b;
    layer5_outputs(9655) <= b;
    layer5_outputs(9656) <= a xor b;
    layer5_outputs(9657) <= not (a or b);
    layer5_outputs(9658) <= not (a and b);
    layer5_outputs(9659) <= a and b;
    layer5_outputs(9660) <= not a;
    layer5_outputs(9661) <= not a;
    layer5_outputs(9662) <= not b;
    layer5_outputs(9663) <= a and b;
    layer5_outputs(9664) <= not b;
    layer5_outputs(9665) <= not b;
    layer5_outputs(9666) <= not (a and b);
    layer5_outputs(9667) <= not a;
    layer5_outputs(9668) <= b;
    layer5_outputs(9669) <= not b;
    layer5_outputs(9670) <= not (a xor b);
    layer5_outputs(9671) <= '1';
    layer5_outputs(9672) <= '1';
    layer5_outputs(9673) <= not b;
    layer5_outputs(9674) <= a;
    layer5_outputs(9675) <= b and not a;
    layer5_outputs(9676) <= not b;
    layer5_outputs(9677) <= a or b;
    layer5_outputs(9678) <= not (a or b);
    layer5_outputs(9679) <= a;
    layer5_outputs(9680) <= b;
    layer5_outputs(9681) <= not a;
    layer5_outputs(9682) <= not (a and b);
    layer5_outputs(9683) <= b;
    layer5_outputs(9684) <= b;
    layer5_outputs(9685) <= a or b;
    layer5_outputs(9686) <= not b or a;
    layer5_outputs(9687) <= not b;
    layer5_outputs(9688) <= a;
    layer5_outputs(9689) <= not b;
    layer5_outputs(9690) <= a or b;
    layer5_outputs(9691) <= not a or b;
    layer5_outputs(9692) <= not a;
    layer5_outputs(9693) <= a;
    layer5_outputs(9694) <= not b;
    layer5_outputs(9695) <= not b;
    layer5_outputs(9696) <= not a;
    layer5_outputs(9697) <= a;
    layer5_outputs(9698) <= not a or b;
    layer5_outputs(9699) <= not b or a;
    layer5_outputs(9700) <= a and b;
    layer5_outputs(9701) <= not a;
    layer5_outputs(9702) <= not a or b;
    layer5_outputs(9703) <= a and b;
    layer5_outputs(9704) <= not b;
    layer5_outputs(9705) <= not b or a;
    layer5_outputs(9706) <= not (a and b);
    layer5_outputs(9707) <= not a;
    layer5_outputs(9708) <= not b or a;
    layer5_outputs(9709) <= not a;
    layer5_outputs(9710) <= not b or a;
    layer5_outputs(9711) <= a xor b;
    layer5_outputs(9712) <= a and not b;
    layer5_outputs(9713) <= not b;
    layer5_outputs(9714) <= a xor b;
    layer5_outputs(9715) <= b and not a;
    layer5_outputs(9716) <= a;
    layer5_outputs(9717) <= a;
    layer5_outputs(9718) <= a and not b;
    layer5_outputs(9719) <= not (a and b);
    layer5_outputs(9720) <= b;
    layer5_outputs(9721) <= a and not b;
    layer5_outputs(9722) <= not b or a;
    layer5_outputs(9723) <= not a;
    layer5_outputs(9724) <= a xor b;
    layer5_outputs(9725) <= not a;
    layer5_outputs(9726) <= not a;
    layer5_outputs(9727) <= a and b;
    layer5_outputs(9728) <= not b;
    layer5_outputs(9729) <= not (a xor b);
    layer5_outputs(9730) <= b;
    layer5_outputs(9731) <= not a;
    layer5_outputs(9732) <= not a or b;
    layer5_outputs(9733) <= b;
    layer5_outputs(9734) <= not (a and b);
    layer5_outputs(9735) <= not b;
    layer5_outputs(9736) <= a xor b;
    layer5_outputs(9737) <= not (a xor b);
    layer5_outputs(9738) <= a and b;
    layer5_outputs(9739) <= a or b;
    layer5_outputs(9740) <= not b or a;
    layer5_outputs(9741) <= not a;
    layer5_outputs(9742) <= not a or b;
    layer5_outputs(9743) <= not a;
    layer5_outputs(9744) <= not b;
    layer5_outputs(9745) <= not (a and b);
    layer5_outputs(9746) <= not (a or b);
    layer5_outputs(9747) <= not a;
    layer5_outputs(9748) <= not (a xor b);
    layer5_outputs(9749) <= a xor b;
    layer5_outputs(9750) <= not b;
    layer5_outputs(9751) <= not a;
    layer5_outputs(9752) <= a or b;
    layer5_outputs(9753) <= not (a xor b);
    layer5_outputs(9754) <= a;
    layer5_outputs(9755) <= not b;
    layer5_outputs(9756) <= b;
    layer5_outputs(9757) <= not a;
    layer5_outputs(9758) <= a;
    layer5_outputs(9759) <= not b;
    layer5_outputs(9760) <= b;
    layer5_outputs(9761) <= not b;
    layer5_outputs(9762) <= not b or a;
    layer5_outputs(9763) <= not b;
    layer5_outputs(9764) <= b;
    layer5_outputs(9765) <= not b;
    layer5_outputs(9766) <= not b or a;
    layer5_outputs(9767) <= a;
    layer5_outputs(9768) <= not (a and b);
    layer5_outputs(9769) <= a;
    layer5_outputs(9770) <= '1';
    layer5_outputs(9771) <= b and not a;
    layer5_outputs(9772) <= b and not a;
    layer5_outputs(9773) <= not a or b;
    layer5_outputs(9774) <= a;
    layer5_outputs(9775) <= not (a xor b);
    layer5_outputs(9776) <= b and not a;
    layer5_outputs(9777) <= not b or a;
    layer5_outputs(9778) <= not (a and b);
    layer5_outputs(9779) <= not b;
    layer5_outputs(9780) <= a;
    layer5_outputs(9781) <= not a;
    layer5_outputs(9782) <= b;
    layer5_outputs(9783) <= b;
    layer5_outputs(9784) <= not a or b;
    layer5_outputs(9785) <= not (a or b);
    layer5_outputs(9786) <= not (a or b);
    layer5_outputs(9787) <= a or b;
    layer5_outputs(9788) <= a and b;
    layer5_outputs(9789) <= not a or b;
    layer5_outputs(9790) <= a;
    layer5_outputs(9791) <= not b;
    layer5_outputs(9792) <= not b;
    layer5_outputs(9793) <= not b;
    layer5_outputs(9794) <= '1';
    layer5_outputs(9795) <= a;
    layer5_outputs(9796) <= not (a and b);
    layer5_outputs(9797) <= a and not b;
    layer5_outputs(9798) <= a;
    layer5_outputs(9799) <= b;
    layer5_outputs(9800) <= not (a xor b);
    layer5_outputs(9801) <= not (a or b);
    layer5_outputs(9802) <= a xor b;
    layer5_outputs(9803) <= a and not b;
    layer5_outputs(9804) <= b;
    layer5_outputs(9805) <= b;
    layer5_outputs(9806) <= a and not b;
    layer5_outputs(9807) <= a;
    layer5_outputs(9808) <= a xor b;
    layer5_outputs(9809) <= b;
    layer5_outputs(9810) <= not b;
    layer5_outputs(9811) <= not (a and b);
    layer5_outputs(9812) <= a or b;
    layer5_outputs(9813) <= a and b;
    layer5_outputs(9814) <= a;
    layer5_outputs(9815) <= b and not a;
    layer5_outputs(9816) <= not a;
    layer5_outputs(9817) <= '1';
    layer5_outputs(9818) <= not a or b;
    layer5_outputs(9819) <= not (a xor b);
    layer5_outputs(9820) <= b;
    layer5_outputs(9821) <= a and b;
    layer5_outputs(9822) <= not a;
    layer5_outputs(9823) <= not a;
    layer5_outputs(9824) <= b;
    layer5_outputs(9825) <= not b or a;
    layer5_outputs(9826) <= a or b;
    layer5_outputs(9827) <= a and b;
    layer5_outputs(9828) <= a or b;
    layer5_outputs(9829) <= not (a or b);
    layer5_outputs(9830) <= a or b;
    layer5_outputs(9831) <= not b;
    layer5_outputs(9832) <= not b;
    layer5_outputs(9833) <= b and not a;
    layer5_outputs(9834) <= a xor b;
    layer5_outputs(9835) <= a;
    layer5_outputs(9836) <= b;
    layer5_outputs(9837) <= b;
    layer5_outputs(9838) <= b;
    layer5_outputs(9839) <= not (a xor b);
    layer5_outputs(9840) <= a xor b;
    layer5_outputs(9841) <= not (a xor b);
    layer5_outputs(9842) <= not (a xor b);
    layer5_outputs(9843) <= not (a xor b);
    layer5_outputs(9844) <= b and not a;
    layer5_outputs(9845) <= a xor b;
    layer5_outputs(9846) <= b;
    layer5_outputs(9847) <= b and not a;
    layer5_outputs(9848) <= b and not a;
    layer5_outputs(9849) <= not b or a;
    layer5_outputs(9850) <= a and b;
    layer5_outputs(9851) <= a or b;
    layer5_outputs(9852) <= b;
    layer5_outputs(9853) <= a xor b;
    layer5_outputs(9854) <= not (a or b);
    layer5_outputs(9855) <= b;
    layer5_outputs(9856) <= not a or b;
    layer5_outputs(9857) <= b;
    layer5_outputs(9858) <= not a;
    layer5_outputs(9859) <= a;
    layer5_outputs(9860) <= not (a or b);
    layer5_outputs(9861) <= not (a xor b);
    layer5_outputs(9862) <= not (a or b);
    layer5_outputs(9863) <= b;
    layer5_outputs(9864) <= a or b;
    layer5_outputs(9865) <= not a;
    layer5_outputs(9866) <= a and b;
    layer5_outputs(9867) <= not a or b;
    layer5_outputs(9868) <= not b;
    layer5_outputs(9869) <= not (a xor b);
    layer5_outputs(9870) <= b;
    layer5_outputs(9871) <= not (a xor b);
    layer5_outputs(9872) <= b;
    layer5_outputs(9873) <= not b;
    layer5_outputs(9874) <= a;
    layer5_outputs(9875) <= a xor b;
    layer5_outputs(9876) <= a or b;
    layer5_outputs(9877) <= a;
    layer5_outputs(9878) <= not (a and b);
    layer5_outputs(9879) <= a xor b;
    layer5_outputs(9880) <= not (a or b);
    layer5_outputs(9881) <= a and not b;
    layer5_outputs(9882) <= '1';
    layer5_outputs(9883) <= a and b;
    layer5_outputs(9884) <= a xor b;
    layer5_outputs(9885) <= a xor b;
    layer5_outputs(9886) <= a;
    layer5_outputs(9887) <= a;
    layer5_outputs(9888) <= a or b;
    layer5_outputs(9889) <= '1';
    layer5_outputs(9890) <= a xor b;
    layer5_outputs(9891) <= not a;
    layer5_outputs(9892) <= not (a and b);
    layer5_outputs(9893) <= '0';
    layer5_outputs(9894) <= a and b;
    layer5_outputs(9895) <= not (a and b);
    layer5_outputs(9896) <= not (a or b);
    layer5_outputs(9897) <= a xor b;
    layer5_outputs(9898) <= not (a and b);
    layer5_outputs(9899) <= a and b;
    layer5_outputs(9900) <= a;
    layer5_outputs(9901) <= b;
    layer5_outputs(9902) <= b;
    layer5_outputs(9903) <= not a or b;
    layer5_outputs(9904) <= a or b;
    layer5_outputs(9905) <= a or b;
    layer5_outputs(9906) <= not a;
    layer5_outputs(9907) <= '1';
    layer5_outputs(9908) <= b;
    layer5_outputs(9909) <= not a or b;
    layer5_outputs(9910) <= a xor b;
    layer5_outputs(9911) <= a or b;
    layer5_outputs(9912) <= not b;
    layer5_outputs(9913) <= not b or a;
    layer5_outputs(9914) <= a and b;
    layer5_outputs(9915) <= a xor b;
    layer5_outputs(9916) <= a xor b;
    layer5_outputs(9917) <= b;
    layer5_outputs(9918) <= b;
    layer5_outputs(9919) <= b;
    layer5_outputs(9920) <= not (a xor b);
    layer5_outputs(9921) <= not (a and b);
    layer5_outputs(9922) <= b;
    layer5_outputs(9923) <= b and not a;
    layer5_outputs(9924) <= b;
    layer5_outputs(9925) <= not a;
    layer5_outputs(9926) <= a xor b;
    layer5_outputs(9927) <= not (a or b);
    layer5_outputs(9928) <= not a;
    layer5_outputs(9929) <= not a or b;
    layer5_outputs(9930) <= a and b;
    layer5_outputs(9931) <= a or b;
    layer5_outputs(9932) <= not (a and b);
    layer5_outputs(9933) <= not a or b;
    layer5_outputs(9934) <= a xor b;
    layer5_outputs(9935) <= a xor b;
    layer5_outputs(9936) <= a and b;
    layer5_outputs(9937) <= a;
    layer5_outputs(9938) <= a and b;
    layer5_outputs(9939) <= a and not b;
    layer5_outputs(9940) <= not b;
    layer5_outputs(9941) <= b;
    layer5_outputs(9942) <= b;
    layer5_outputs(9943) <= not (a and b);
    layer5_outputs(9944) <= not a;
    layer5_outputs(9945) <= not a;
    layer5_outputs(9946) <= a or b;
    layer5_outputs(9947) <= not b;
    layer5_outputs(9948) <= a;
    layer5_outputs(9949) <= not b or a;
    layer5_outputs(9950) <= a or b;
    layer5_outputs(9951) <= not (a and b);
    layer5_outputs(9952) <= not a;
    layer5_outputs(9953) <= a and not b;
    layer5_outputs(9954) <= not a;
    layer5_outputs(9955) <= not a;
    layer5_outputs(9956) <= b;
    layer5_outputs(9957) <= a and b;
    layer5_outputs(9958) <= not a;
    layer5_outputs(9959) <= not (a xor b);
    layer5_outputs(9960) <= b and not a;
    layer5_outputs(9961) <= not b or a;
    layer5_outputs(9962) <= not (a and b);
    layer5_outputs(9963) <= not (a or b);
    layer5_outputs(9964) <= not (a or b);
    layer5_outputs(9965) <= a xor b;
    layer5_outputs(9966) <= b;
    layer5_outputs(9967) <= b and not a;
    layer5_outputs(9968) <= a and b;
    layer5_outputs(9969) <= a;
    layer5_outputs(9970) <= not b;
    layer5_outputs(9971) <= not a;
    layer5_outputs(9972) <= a xor b;
    layer5_outputs(9973) <= not (a xor b);
    layer5_outputs(9974) <= b;
    layer5_outputs(9975) <= b;
    layer5_outputs(9976) <= b;
    layer5_outputs(9977) <= not a;
    layer5_outputs(9978) <= b and not a;
    layer5_outputs(9979) <= not a;
    layer5_outputs(9980) <= not b;
    layer5_outputs(9981) <= a;
    layer5_outputs(9982) <= not b;
    layer5_outputs(9983) <= b;
    layer5_outputs(9984) <= a;
    layer5_outputs(9985) <= '0';
    layer5_outputs(9986) <= a and b;
    layer5_outputs(9987) <= b;
    layer5_outputs(9988) <= b and not a;
    layer5_outputs(9989) <= a;
    layer5_outputs(9990) <= a and b;
    layer5_outputs(9991) <= b;
    layer5_outputs(9992) <= a;
    layer5_outputs(9993) <= b and not a;
    layer5_outputs(9994) <= '0';
    layer5_outputs(9995) <= not (a xor b);
    layer5_outputs(9996) <= a or b;
    layer5_outputs(9997) <= a;
    layer5_outputs(9998) <= not b;
    layer5_outputs(9999) <= b and not a;
    layer5_outputs(10000) <= not (a xor b);
    layer5_outputs(10001) <= not a;
    layer5_outputs(10002) <= not a;
    layer5_outputs(10003) <= a or b;
    layer5_outputs(10004) <= not a;
    layer5_outputs(10005) <= a;
    layer5_outputs(10006) <= not b;
    layer5_outputs(10007) <= not a;
    layer5_outputs(10008) <= not a or b;
    layer5_outputs(10009) <= not a or b;
    layer5_outputs(10010) <= b;
    layer5_outputs(10011) <= a xor b;
    layer5_outputs(10012) <= a or b;
    layer5_outputs(10013) <= a;
    layer5_outputs(10014) <= not b;
    layer5_outputs(10015) <= not b or a;
    layer5_outputs(10016) <= a xor b;
    layer5_outputs(10017) <= a;
    layer5_outputs(10018) <= a and b;
    layer5_outputs(10019) <= a and b;
    layer5_outputs(10020) <= a xor b;
    layer5_outputs(10021) <= a xor b;
    layer5_outputs(10022) <= a;
    layer5_outputs(10023) <= not b or a;
    layer5_outputs(10024) <= not b;
    layer5_outputs(10025) <= not b or a;
    layer5_outputs(10026) <= a and not b;
    layer5_outputs(10027) <= not (a and b);
    layer5_outputs(10028) <= a or b;
    layer5_outputs(10029) <= b;
    layer5_outputs(10030) <= b and not a;
    layer5_outputs(10031) <= not (a xor b);
    layer5_outputs(10032) <= a;
    layer5_outputs(10033) <= not (a or b);
    layer5_outputs(10034) <= a xor b;
    layer5_outputs(10035) <= a and not b;
    layer5_outputs(10036) <= a;
    layer5_outputs(10037) <= b;
    layer5_outputs(10038) <= not b;
    layer5_outputs(10039) <= not (a or b);
    layer5_outputs(10040) <= not a;
    layer5_outputs(10041) <= b and not a;
    layer5_outputs(10042) <= not b;
    layer5_outputs(10043) <= not b;
    layer5_outputs(10044) <= not (a or b);
    layer5_outputs(10045) <= not (a and b);
    layer5_outputs(10046) <= a;
    layer5_outputs(10047) <= not (a and b);
    layer5_outputs(10048) <= a and b;
    layer5_outputs(10049) <= b;
    layer5_outputs(10050) <= a or b;
    layer5_outputs(10051) <= b and not a;
    layer5_outputs(10052) <= not b;
    layer5_outputs(10053) <= not b;
    layer5_outputs(10054) <= not b;
    layer5_outputs(10055) <= not a;
    layer5_outputs(10056) <= a;
    layer5_outputs(10057) <= not b;
    layer5_outputs(10058) <= b;
    layer5_outputs(10059) <= not (a xor b);
    layer5_outputs(10060) <= not a;
    layer5_outputs(10061) <= a;
    layer5_outputs(10062) <= not a;
    layer5_outputs(10063) <= not b;
    layer5_outputs(10064) <= a and not b;
    layer5_outputs(10065) <= a and not b;
    layer5_outputs(10066) <= not b or a;
    layer5_outputs(10067) <= not (a and b);
    layer5_outputs(10068) <= b and not a;
    layer5_outputs(10069) <= not a or b;
    layer5_outputs(10070) <= b;
    layer5_outputs(10071) <= a xor b;
    layer5_outputs(10072) <= b and not a;
    layer5_outputs(10073) <= a;
    layer5_outputs(10074) <= a xor b;
    layer5_outputs(10075) <= not (a or b);
    layer5_outputs(10076) <= a or b;
    layer5_outputs(10077) <= not b;
    layer5_outputs(10078) <= a and not b;
    layer5_outputs(10079) <= a;
    layer5_outputs(10080) <= not (a xor b);
    layer5_outputs(10081) <= a;
    layer5_outputs(10082) <= not (a xor b);
    layer5_outputs(10083) <= '0';
    layer5_outputs(10084) <= a xor b;
    layer5_outputs(10085) <= not a;
    layer5_outputs(10086) <= not a;
    layer5_outputs(10087) <= not (a and b);
    layer5_outputs(10088) <= b;
    layer5_outputs(10089) <= a xor b;
    layer5_outputs(10090) <= a and b;
    layer5_outputs(10091) <= a and not b;
    layer5_outputs(10092) <= not b or a;
    layer5_outputs(10093) <= not a;
    layer5_outputs(10094) <= a;
    layer5_outputs(10095) <= not (a and b);
    layer5_outputs(10096) <= a and not b;
    layer5_outputs(10097) <= a xor b;
    layer5_outputs(10098) <= not b;
    layer5_outputs(10099) <= a and not b;
    layer5_outputs(10100) <= not (a and b);
    layer5_outputs(10101) <= not (a and b);
    layer5_outputs(10102) <= b and not a;
    layer5_outputs(10103) <= a and not b;
    layer5_outputs(10104) <= b;
    layer5_outputs(10105) <= b;
    layer5_outputs(10106) <= '0';
    layer5_outputs(10107) <= b and not a;
    layer5_outputs(10108) <= b;
    layer5_outputs(10109) <= b and not a;
    layer5_outputs(10110) <= not a;
    layer5_outputs(10111) <= a;
    layer5_outputs(10112) <= not a;
    layer5_outputs(10113) <= not (a xor b);
    layer5_outputs(10114) <= not a;
    layer5_outputs(10115) <= not a;
    layer5_outputs(10116) <= not b;
    layer5_outputs(10117) <= not (a or b);
    layer5_outputs(10118) <= b;
    layer5_outputs(10119) <= not a;
    layer5_outputs(10120) <= not a or b;
    layer5_outputs(10121) <= a or b;
    layer5_outputs(10122) <= not (a and b);
    layer5_outputs(10123) <= a;
    layer5_outputs(10124) <= not b;
    layer5_outputs(10125) <= a;
    layer5_outputs(10126) <= a;
    layer5_outputs(10127) <= a xor b;
    layer5_outputs(10128) <= '1';
    layer5_outputs(10129) <= not (a or b);
    layer5_outputs(10130) <= a;
    layer5_outputs(10131) <= a;
    layer5_outputs(10132) <= a xor b;
    layer5_outputs(10133) <= b;
    layer5_outputs(10134) <= not (a or b);
    layer5_outputs(10135) <= a;
    layer5_outputs(10136) <= a and not b;
    layer5_outputs(10137) <= not a;
    layer5_outputs(10138) <= b;
    layer5_outputs(10139) <= not b;
    layer5_outputs(10140) <= not a or b;
    layer5_outputs(10141) <= b;
    layer5_outputs(10142) <= a;
    layer5_outputs(10143) <= b;
    layer5_outputs(10144) <= not (a xor b);
    layer5_outputs(10145) <= not (a and b);
    layer5_outputs(10146) <= a or b;
    layer5_outputs(10147) <= not (a xor b);
    layer5_outputs(10148) <= not b;
    layer5_outputs(10149) <= b;
    layer5_outputs(10150) <= a;
    layer5_outputs(10151) <= a or b;
    layer5_outputs(10152) <= b;
    layer5_outputs(10153) <= not b or a;
    layer5_outputs(10154) <= a;
    layer5_outputs(10155) <= not a or b;
    layer5_outputs(10156) <= not b;
    layer5_outputs(10157) <= not b or a;
    layer5_outputs(10158) <= a or b;
    layer5_outputs(10159) <= not a or b;
    layer5_outputs(10160) <= a and b;
    layer5_outputs(10161) <= not b;
    layer5_outputs(10162) <= not (a or b);
    layer5_outputs(10163) <= not (a xor b);
    layer5_outputs(10164) <= b;
    layer5_outputs(10165) <= not a or b;
    layer5_outputs(10166) <= b;
    layer5_outputs(10167) <= b;
    layer5_outputs(10168) <= not a;
    layer5_outputs(10169) <= not a;
    layer5_outputs(10170) <= a or b;
    layer5_outputs(10171) <= a;
    layer5_outputs(10172) <= a xor b;
    layer5_outputs(10173) <= not a;
    layer5_outputs(10174) <= a xor b;
    layer5_outputs(10175) <= b and not a;
    layer5_outputs(10176) <= a;
    layer5_outputs(10177) <= not (a or b);
    layer5_outputs(10178) <= not (a and b);
    layer5_outputs(10179) <= not a;
    layer5_outputs(10180) <= not b;
    layer5_outputs(10181) <= a xor b;
    layer5_outputs(10182) <= a;
    layer5_outputs(10183) <= b;
    layer5_outputs(10184) <= a;
    layer5_outputs(10185) <= b;
    layer5_outputs(10186) <= b;
    layer5_outputs(10187) <= not (a and b);
    layer5_outputs(10188) <= not a or b;
    layer5_outputs(10189) <= b;
    layer5_outputs(10190) <= a or b;
    layer5_outputs(10191) <= a or b;
    layer5_outputs(10192) <= not b;
    layer5_outputs(10193) <= not (a or b);
    layer5_outputs(10194) <= a;
    layer5_outputs(10195) <= not (a xor b);
    layer5_outputs(10196) <= a;
    layer5_outputs(10197) <= b;
    layer5_outputs(10198) <= not a or b;
    layer5_outputs(10199) <= a;
    layer5_outputs(10200) <= a xor b;
    layer5_outputs(10201) <= not (a or b);
    layer5_outputs(10202) <= b;
    layer5_outputs(10203) <= not (a and b);
    layer5_outputs(10204) <= a and not b;
    layer5_outputs(10205) <= not b;
    layer5_outputs(10206) <= not b;
    layer5_outputs(10207) <= a and b;
    layer5_outputs(10208) <= a and b;
    layer5_outputs(10209) <= a and not b;
    layer5_outputs(10210) <= not a;
    layer5_outputs(10211) <= a;
    layer5_outputs(10212) <= not a;
    layer5_outputs(10213) <= not (a or b);
    layer5_outputs(10214) <= not a;
    layer5_outputs(10215) <= a;
    layer5_outputs(10216) <= a and not b;
    layer5_outputs(10217) <= a or b;
    layer5_outputs(10218) <= not (a xor b);
    layer5_outputs(10219) <= b;
    layer5_outputs(10220) <= not a;
    layer5_outputs(10221) <= a;
    layer5_outputs(10222) <= not a;
    layer5_outputs(10223) <= not a;
    layer5_outputs(10224) <= not (a or b);
    layer5_outputs(10225) <= not (a and b);
    layer5_outputs(10226) <= a;
    layer5_outputs(10227) <= not b or a;
    layer5_outputs(10228) <= b and not a;
    layer5_outputs(10229) <= not (a or b);
    layer5_outputs(10230) <= b;
    layer5_outputs(10231) <= a and b;
    layer5_outputs(10232) <= b;
    layer5_outputs(10233) <= not a;
    layer5_outputs(10234) <= b;
    layer5_outputs(10235) <= a;
    layer5_outputs(10236) <= not a;
    layer5_outputs(10237) <= not b;
    layer5_outputs(10238) <= not (a or b);
    layer5_outputs(10239) <= a and not b;
    layer5_outputs(10240) <= not (a or b);
    layer5_outputs(10241) <= not a;
    layer5_outputs(10242) <= not b or a;
    layer5_outputs(10243) <= b;
    layer5_outputs(10244) <= not b;
    layer5_outputs(10245) <= a;
    layer5_outputs(10246) <= b;
    layer5_outputs(10247) <= not a;
    layer5_outputs(10248) <= a;
    layer5_outputs(10249) <= not b;
    layer5_outputs(10250) <= b;
    layer5_outputs(10251) <= b and not a;
    layer5_outputs(10252) <= not b or a;
    layer5_outputs(10253) <= a xor b;
    layer5_outputs(10254) <= a or b;
    layer5_outputs(10255) <= not b or a;
    layer5_outputs(10256) <= not a;
    layer5_outputs(10257) <= not (a and b);
    layer5_outputs(10258) <= a;
    layer5_outputs(10259) <= b;
    layer5_outputs(10260) <= a or b;
    layer5_outputs(10261) <= not a;
    layer5_outputs(10262) <= a xor b;
    layer5_outputs(10263) <= not (a and b);
    layer5_outputs(10264) <= a and not b;
    layer5_outputs(10265) <= not b;
    layer5_outputs(10266) <= not a or b;
    layer5_outputs(10267) <= not (a xor b);
    layer5_outputs(10268) <= not a;
    layer5_outputs(10269) <= b;
    layer5_outputs(10270) <= a and not b;
    layer5_outputs(10271) <= not a;
    layer5_outputs(10272) <= b;
    layer5_outputs(10273) <= a;
    layer5_outputs(10274) <= not b or a;
    layer5_outputs(10275) <= not a;
    layer5_outputs(10276) <= a;
    layer5_outputs(10277) <= not b;
    layer5_outputs(10278) <= not b or a;
    layer5_outputs(10279) <= a xor b;
    layer5_outputs(10280) <= not (a or b);
    layer5_outputs(10281) <= b and not a;
    layer5_outputs(10282) <= not (a and b);
    layer5_outputs(10283) <= not (a xor b);
    layer5_outputs(10284) <= not a or b;
    layer5_outputs(10285) <= a and b;
    layer5_outputs(10286) <= a and b;
    layer5_outputs(10287) <= not (a and b);
    layer5_outputs(10288) <= not (a xor b);
    layer5_outputs(10289) <= b and not a;
    layer5_outputs(10290) <= a;
    layer5_outputs(10291) <= not b;
    layer5_outputs(10292) <= not (a and b);
    layer5_outputs(10293) <= a;
    layer5_outputs(10294) <= not (a or b);
    layer5_outputs(10295) <= a and b;
    layer5_outputs(10296) <= b;
    layer5_outputs(10297) <= b;
    layer5_outputs(10298) <= b and not a;
    layer5_outputs(10299) <= b;
    layer5_outputs(10300) <= b;
    layer5_outputs(10301) <= not a;
    layer5_outputs(10302) <= not (a xor b);
    layer5_outputs(10303) <= not a or b;
    layer5_outputs(10304) <= b and not a;
    layer5_outputs(10305) <= not a;
    layer5_outputs(10306) <= not b;
    layer5_outputs(10307) <= a;
    layer5_outputs(10308) <= b and not a;
    layer5_outputs(10309) <= not b or a;
    layer5_outputs(10310) <= not (a or b);
    layer5_outputs(10311) <= not (a or b);
    layer5_outputs(10312) <= b;
    layer5_outputs(10313) <= not a;
    layer5_outputs(10314) <= a;
    layer5_outputs(10315) <= not b or a;
    layer5_outputs(10316) <= not a;
    layer5_outputs(10317) <= not a or b;
    layer5_outputs(10318) <= a xor b;
    layer5_outputs(10319) <= a or b;
    layer5_outputs(10320) <= not (a or b);
    layer5_outputs(10321) <= a xor b;
    layer5_outputs(10322) <= a xor b;
    layer5_outputs(10323) <= not (a xor b);
    layer5_outputs(10324) <= a and b;
    layer5_outputs(10325) <= a and not b;
    layer5_outputs(10326) <= a and not b;
    layer5_outputs(10327) <= not a;
    layer5_outputs(10328) <= a and b;
    layer5_outputs(10329) <= not b or a;
    layer5_outputs(10330) <= a and b;
    layer5_outputs(10331) <= not a;
    layer5_outputs(10332) <= not (a or b);
    layer5_outputs(10333) <= a xor b;
    layer5_outputs(10334) <= a or b;
    layer5_outputs(10335) <= not a;
    layer5_outputs(10336) <= not (a and b);
    layer5_outputs(10337) <= a and not b;
    layer5_outputs(10338) <= not a or b;
    layer5_outputs(10339) <= not a;
    layer5_outputs(10340) <= not (a or b);
    layer5_outputs(10341) <= a and b;
    layer5_outputs(10342) <= not (a xor b);
    layer5_outputs(10343) <= not (a xor b);
    layer5_outputs(10344) <= not (a or b);
    layer5_outputs(10345) <= not (a xor b);
    layer5_outputs(10346) <= not b;
    layer5_outputs(10347) <= a and not b;
    layer5_outputs(10348) <= not b or a;
    layer5_outputs(10349) <= not a;
    layer5_outputs(10350) <= not b;
    layer5_outputs(10351) <= not (a or b);
    layer5_outputs(10352) <= not b;
    layer5_outputs(10353) <= a;
    layer5_outputs(10354) <= not b or a;
    layer5_outputs(10355) <= a and not b;
    layer5_outputs(10356) <= a;
    layer5_outputs(10357) <= not (a xor b);
    layer5_outputs(10358) <= not (a xor b);
    layer5_outputs(10359) <= b;
    layer5_outputs(10360) <= a or b;
    layer5_outputs(10361) <= b and not a;
    layer5_outputs(10362) <= a and not b;
    layer5_outputs(10363) <= not (a or b);
    layer5_outputs(10364) <= not a;
    layer5_outputs(10365) <= not b;
    layer5_outputs(10366) <= a and not b;
    layer5_outputs(10367) <= b;
    layer5_outputs(10368) <= not b or a;
    layer5_outputs(10369) <= not b or a;
    layer5_outputs(10370) <= b;
    layer5_outputs(10371) <= a xor b;
    layer5_outputs(10372) <= a;
    layer5_outputs(10373) <= not b;
    layer5_outputs(10374) <= a and not b;
    layer5_outputs(10375) <= not (a and b);
    layer5_outputs(10376) <= not (a and b);
    layer5_outputs(10377) <= a xor b;
    layer5_outputs(10378) <= not (a or b);
    layer5_outputs(10379) <= not a or b;
    layer5_outputs(10380) <= not (a or b);
    layer5_outputs(10381) <= not (a xor b);
    layer5_outputs(10382) <= a;
    layer5_outputs(10383) <= not b;
    layer5_outputs(10384) <= b and not a;
    layer5_outputs(10385) <= not b;
    layer5_outputs(10386) <= not (a or b);
    layer5_outputs(10387) <= not a;
    layer5_outputs(10388) <= not b;
    layer5_outputs(10389) <= b;
    layer5_outputs(10390) <= b and not a;
    layer5_outputs(10391) <= not (a and b);
    layer5_outputs(10392) <= b;
    layer5_outputs(10393) <= a and b;
    layer5_outputs(10394) <= not a or b;
    layer5_outputs(10395) <= not a or b;
    layer5_outputs(10396) <= not (a xor b);
    layer5_outputs(10397) <= a xor b;
    layer5_outputs(10398) <= b;
    layer5_outputs(10399) <= not (a or b);
    layer5_outputs(10400) <= not (a xor b);
    layer5_outputs(10401) <= not b;
    layer5_outputs(10402) <= a and b;
    layer5_outputs(10403) <= not a;
    layer5_outputs(10404) <= not b;
    layer5_outputs(10405) <= not b;
    layer5_outputs(10406) <= not b or a;
    layer5_outputs(10407) <= not (a xor b);
    layer5_outputs(10408) <= not (a and b);
    layer5_outputs(10409) <= b;
    layer5_outputs(10410) <= not a;
    layer5_outputs(10411) <= a;
    layer5_outputs(10412) <= a xor b;
    layer5_outputs(10413) <= a xor b;
    layer5_outputs(10414) <= not (a or b);
    layer5_outputs(10415) <= a and not b;
    layer5_outputs(10416) <= a;
    layer5_outputs(10417) <= a xor b;
    layer5_outputs(10418) <= a and b;
    layer5_outputs(10419) <= not b;
    layer5_outputs(10420) <= not a;
    layer5_outputs(10421) <= a or b;
    layer5_outputs(10422) <= not (a and b);
    layer5_outputs(10423) <= b;
    layer5_outputs(10424) <= not b or a;
    layer5_outputs(10425) <= b;
    layer5_outputs(10426) <= not a;
    layer5_outputs(10427) <= not b;
    layer5_outputs(10428) <= not (a xor b);
    layer5_outputs(10429) <= a;
    layer5_outputs(10430) <= not a;
    layer5_outputs(10431) <= b;
    layer5_outputs(10432) <= a xor b;
    layer5_outputs(10433) <= a and b;
    layer5_outputs(10434) <= not b;
    layer5_outputs(10435) <= b and not a;
    layer5_outputs(10436) <= b;
    layer5_outputs(10437) <= a xor b;
    layer5_outputs(10438) <= a and b;
    layer5_outputs(10439) <= a;
    layer5_outputs(10440) <= not a;
    layer5_outputs(10441) <= b and not a;
    layer5_outputs(10442) <= a xor b;
    layer5_outputs(10443) <= a;
    layer5_outputs(10444) <= not a;
    layer5_outputs(10445) <= not (a or b);
    layer5_outputs(10446) <= a and not b;
    layer5_outputs(10447) <= not a;
    layer5_outputs(10448) <= a xor b;
    layer5_outputs(10449) <= not a or b;
    layer5_outputs(10450) <= not a or b;
    layer5_outputs(10451) <= a;
    layer5_outputs(10452) <= a and not b;
    layer5_outputs(10453) <= not (a xor b);
    layer5_outputs(10454) <= a and b;
    layer5_outputs(10455) <= not (a and b);
    layer5_outputs(10456) <= a or b;
    layer5_outputs(10457) <= a and not b;
    layer5_outputs(10458) <= not b;
    layer5_outputs(10459) <= a or b;
    layer5_outputs(10460) <= a and b;
    layer5_outputs(10461) <= not a or b;
    layer5_outputs(10462) <= not b or a;
    layer5_outputs(10463) <= b and not a;
    layer5_outputs(10464) <= not a;
    layer5_outputs(10465) <= not a;
    layer5_outputs(10466) <= not b;
    layer5_outputs(10467) <= not a;
    layer5_outputs(10468) <= not b or a;
    layer5_outputs(10469) <= not b or a;
    layer5_outputs(10470) <= not b or a;
    layer5_outputs(10471) <= a;
    layer5_outputs(10472) <= not a;
    layer5_outputs(10473) <= a;
    layer5_outputs(10474) <= not (a xor b);
    layer5_outputs(10475) <= a;
    layer5_outputs(10476) <= a xor b;
    layer5_outputs(10477) <= a xor b;
    layer5_outputs(10478) <= a;
    layer5_outputs(10479) <= b;
    layer5_outputs(10480) <= a xor b;
    layer5_outputs(10481) <= not (a and b);
    layer5_outputs(10482) <= not a;
    layer5_outputs(10483) <= b and not a;
    layer5_outputs(10484) <= b and not a;
    layer5_outputs(10485) <= b;
    layer5_outputs(10486) <= a;
    layer5_outputs(10487) <= b;
    layer5_outputs(10488) <= not (a or b);
    layer5_outputs(10489) <= not (a or b);
    layer5_outputs(10490) <= a;
    layer5_outputs(10491) <= a and b;
    layer5_outputs(10492) <= not a;
    layer5_outputs(10493) <= not b;
    layer5_outputs(10494) <= a;
    layer5_outputs(10495) <= b;
    layer5_outputs(10496) <= b and not a;
    layer5_outputs(10497) <= not b;
    layer5_outputs(10498) <= not b;
    layer5_outputs(10499) <= not b or a;
    layer5_outputs(10500) <= a or b;
    layer5_outputs(10501) <= not a;
    layer5_outputs(10502) <= a;
    layer5_outputs(10503) <= not a;
    layer5_outputs(10504) <= not (a xor b);
    layer5_outputs(10505) <= a and b;
    layer5_outputs(10506) <= a;
    layer5_outputs(10507) <= b;
    layer5_outputs(10508) <= not a;
    layer5_outputs(10509) <= a or b;
    layer5_outputs(10510) <= not (a xor b);
    layer5_outputs(10511) <= a;
    layer5_outputs(10512) <= not (a or b);
    layer5_outputs(10513) <= not b;
    layer5_outputs(10514) <= a and b;
    layer5_outputs(10515) <= b;
    layer5_outputs(10516) <= not b;
    layer5_outputs(10517) <= b;
    layer5_outputs(10518) <= b and not a;
    layer5_outputs(10519) <= a;
    layer5_outputs(10520) <= not (a or b);
    layer5_outputs(10521) <= a and b;
    layer5_outputs(10522) <= not b;
    layer5_outputs(10523) <= not b;
    layer5_outputs(10524) <= not (a or b);
    layer5_outputs(10525) <= not b or a;
    layer5_outputs(10526) <= a and b;
    layer5_outputs(10527) <= a xor b;
    layer5_outputs(10528) <= a or b;
    layer5_outputs(10529) <= not a;
    layer5_outputs(10530) <= '0';
    layer5_outputs(10531) <= a;
    layer5_outputs(10532) <= not b;
    layer5_outputs(10533) <= a;
    layer5_outputs(10534) <= not b;
    layer5_outputs(10535) <= not a or b;
    layer5_outputs(10536) <= a;
    layer5_outputs(10537) <= a and b;
    layer5_outputs(10538) <= not a;
    layer5_outputs(10539) <= b;
    layer5_outputs(10540) <= '1';
    layer5_outputs(10541) <= not b or a;
    layer5_outputs(10542) <= a;
    layer5_outputs(10543) <= a xor b;
    layer5_outputs(10544) <= not (a xor b);
    layer5_outputs(10545) <= a;
    layer5_outputs(10546) <= not (a xor b);
    layer5_outputs(10547) <= not a;
    layer5_outputs(10548) <= b and not a;
    layer5_outputs(10549) <= a;
    layer5_outputs(10550) <= a xor b;
    layer5_outputs(10551) <= not a or b;
    layer5_outputs(10552) <= not (a xor b);
    layer5_outputs(10553) <= not b or a;
    layer5_outputs(10554) <= b;
    layer5_outputs(10555) <= not a;
    layer5_outputs(10556) <= b;
    layer5_outputs(10557) <= b and not a;
    layer5_outputs(10558) <= a or b;
    layer5_outputs(10559) <= b;
    layer5_outputs(10560) <= b and not a;
    layer5_outputs(10561) <= not (a xor b);
    layer5_outputs(10562) <= a;
    layer5_outputs(10563) <= not a;
    layer5_outputs(10564) <= a and not b;
    layer5_outputs(10565) <= not a;
    layer5_outputs(10566) <= a or b;
    layer5_outputs(10567) <= b;
    layer5_outputs(10568) <= b and not a;
    layer5_outputs(10569) <= not b;
    layer5_outputs(10570) <= not a;
    layer5_outputs(10571) <= not b or a;
    layer5_outputs(10572) <= a;
    layer5_outputs(10573) <= not (a xor b);
    layer5_outputs(10574) <= not b;
    layer5_outputs(10575) <= not a;
    layer5_outputs(10576) <= b and not a;
    layer5_outputs(10577) <= not (a and b);
    layer5_outputs(10578) <= b;
    layer5_outputs(10579) <= a;
    layer5_outputs(10580) <= b and not a;
    layer5_outputs(10581) <= not a;
    layer5_outputs(10582) <= not (a xor b);
    layer5_outputs(10583) <= a;
    layer5_outputs(10584) <= a;
    layer5_outputs(10585) <= not (a or b);
    layer5_outputs(10586) <= not a or b;
    layer5_outputs(10587) <= a xor b;
    layer5_outputs(10588) <= not a;
    layer5_outputs(10589) <= b;
    layer5_outputs(10590) <= not a;
    layer5_outputs(10591) <= '0';
    layer5_outputs(10592) <= not a;
    layer5_outputs(10593) <= not a;
    layer5_outputs(10594) <= not a or b;
    layer5_outputs(10595) <= a;
    layer5_outputs(10596) <= not (a or b);
    layer5_outputs(10597) <= b;
    layer5_outputs(10598) <= not (a xor b);
    layer5_outputs(10599) <= a or b;
    layer5_outputs(10600) <= not b or a;
    layer5_outputs(10601) <= a and not b;
    layer5_outputs(10602) <= a;
    layer5_outputs(10603) <= a;
    layer5_outputs(10604) <= not a;
    layer5_outputs(10605) <= a;
    layer5_outputs(10606) <= not b;
    layer5_outputs(10607) <= not b or a;
    layer5_outputs(10608) <= not a;
    layer5_outputs(10609) <= a and b;
    layer5_outputs(10610) <= not (a xor b);
    layer5_outputs(10611) <= a xor b;
    layer5_outputs(10612) <= not b;
    layer5_outputs(10613) <= a;
    layer5_outputs(10614) <= a;
    layer5_outputs(10615) <= not (a and b);
    layer5_outputs(10616) <= a and not b;
    layer5_outputs(10617) <= not (a xor b);
    layer5_outputs(10618) <= a and b;
    layer5_outputs(10619) <= a and not b;
    layer5_outputs(10620) <= not a;
    layer5_outputs(10621) <= not b;
    layer5_outputs(10622) <= a xor b;
    layer5_outputs(10623) <= a and b;
    layer5_outputs(10624) <= not b;
    layer5_outputs(10625) <= not a;
    layer5_outputs(10626) <= not a;
    layer5_outputs(10627) <= a and b;
    layer5_outputs(10628) <= not a;
    layer5_outputs(10629) <= a and not b;
    layer5_outputs(10630) <= not b or a;
    layer5_outputs(10631) <= not a;
    layer5_outputs(10632) <= '1';
    layer5_outputs(10633) <= not (a or b);
    layer5_outputs(10634) <= not b;
    layer5_outputs(10635) <= not (a xor b);
    layer5_outputs(10636) <= a and not b;
    layer5_outputs(10637) <= a xor b;
    layer5_outputs(10638) <= not a;
    layer5_outputs(10639) <= b;
    layer5_outputs(10640) <= not a or b;
    layer5_outputs(10641) <= not (a xor b);
    layer5_outputs(10642) <= a and b;
    layer5_outputs(10643) <= not b;
    layer5_outputs(10644) <= not a;
    layer5_outputs(10645) <= not a;
    layer5_outputs(10646) <= not (a and b);
    layer5_outputs(10647) <= b and not a;
    layer5_outputs(10648) <= not b or a;
    layer5_outputs(10649) <= a;
    layer5_outputs(10650) <= b and not a;
    layer5_outputs(10651) <= not (a and b);
    layer5_outputs(10652) <= not a;
    layer5_outputs(10653) <= not b;
    layer5_outputs(10654) <= a;
    layer5_outputs(10655) <= '0';
    layer5_outputs(10656) <= not b;
    layer5_outputs(10657) <= b and not a;
    layer5_outputs(10658) <= a;
    layer5_outputs(10659) <= a;
    layer5_outputs(10660) <= b;
    layer5_outputs(10661) <= not a;
    layer5_outputs(10662) <= not (a xor b);
    layer5_outputs(10663) <= not (a and b);
    layer5_outputs(10664) <= not a;
    layer5_outputs(10665) <= not a;
    layer5_outputs(10666) <= not a;
    layer5_outputs(10667) <= not (a xor b);
    layer5_outputs(10668) <= b and not a;
    layer5_outputs(10669) <= a;
    layer5_outputs(10670) <= a and b;
    layer5_outputs(10671) <= a or b;
    layer5_outputs(10672) <= a xor b;
    layer5_outputs(10673) <= not b;
    layer5_outputs(10674) <= not (a xor b);
    layer5_outputs(10675) <= not a or b;
    layer5_outputs(10676) <= b and not a;
    layer5_outputs(10677) <= not b;
    layer5_outputs(10678) <= a or b;
    layer5_outputs(10679) <= not b or a;
    layer5_outputs(10680) <= not b or a;
    layer5_outputs(10681) <= '0';
    layer5_outputs(10682) <= not (a or b);
    layer5_outputs(10683) <= not a;
    layer5_outputs(10684) <= b and not a;
    layer5_outputs(10685) <= '1';
    layer5_outputs(10686) <= not b;
    layer5_outputs(10687) <= a and not b;
    layer5_outputs(10688) <= not b or a;
    layer5_outputs(10689) <= not (a and b);
    layer5_outputs(10690) <= not (a xor b);
    layer5_outputs(10691) <= not a or b;
    layer5_outputs(10692) <= a or b;
    layer5_outputs(10693) <= a xor b;
    layer5_outputs(10694) <= not b or a;
    layer5_outputs(10695) <= a and b;
    layer5_outputs(10696) <= b;
    layer5_outputs(10697) <= a or b;
    layer5_outputs(10698) <= a;
    layer5_outputs(10699) <= a or b;
    layer5_outputs(10700) <= not (a xor b);
    layer5_outputs(10701) <= not (a and b);
    layer5_outputs(10702) <= a and not b;
    layer5_outputs(10703) <= b;
    layer5_outputs(10704) <= not a;
    layer5_outputs(10705) <= a;
    layer5_outputs(10706) <= a xor b;
    layer5_outputs(10707) <= not b;
    layer5_outputs(10708) <= not (a or b);
    layer5_outputs(10709) <= a or b;
    layer5_outputs(10710) <= not a;
    layer5_outputs(10711) <= not (a xor b);
    layer5_outputs(10712) <= a xor b;
    layer5_outputs(10713) <= '0';
    layer5_outputs(10714) <= not a or b;
    layer5_outputs(10715) <= not (a and b);
    layer5_outputs(10716) <= b;
    layer5_outputs(10717) <= not (a xor b);
    layer5_outputs(10718) <= a and b;
    layer5_outputs(10719) <= not a;
    layer5_outputs(10720) <= not (a or b);
    layer5_outputs(10721) <= a and b;
    layer5_outputs(10722) <= not a;
    layer5_outputs(10723) <= not b;
    layer5_outputs(10724) <= not b or a;
    layer5_outputs(10725) <= not (a xor b);
    layer5_outputs(10726) <= a;
    layer5_outputs(10727) <= not (a xor b);
    layer5_outputs(10728) <= b;
    layer5_outputs(10729) <= not a or b;
    layer5_outputs(10730) <= not (a and b);
    layer5_outputs(10731) <= a and b;
    layer5_outputs(10732) <= not b;
    layer5_outputs(10733) <= not a;
    layer5_outputs(10734) <= not a;
    layer5_outputs(10735) <= b and not a;
    layer5_outputs(10736) <= a;
    layer5_outputs(10737) <= '0';
    layer5_outputs(10738) <= not b or a;
    layer5_outputs(10739) <= not (a xor b);
    layer5_outputs(10740) <= not b;
    layer5_outputs(10741) <= b and not a;
    layer5_outputs(10742) <= b;
    layer5_outputs(10743) <= not b;
    layer5_outputs(10744) <= a xor b;
    layer5_outputs(10745) <= a xor b;
    layer5_outputs(10746) <= a and b;
    layer5_outputs(10747) <= a;
    layer5_outputs(10748) <= a xor b;
    layer5_outputs(10749) <= a;
    layer5_outputs(10750) <= not (a or b);
    layer5_outputs(10751) <= not b;
    layer5_outputs(10752) <= not b;
    layer5_outputs(10753) <= b;
    layer5_outputs(10754) <= not a;
    layer5_outputs(10755) <= a;
    layer5_outputs(10756) <= a and not b;
    layer5_outputs(10757) <= not b;
    layer5_outputs(10758) <= not (a or b);
    layer5_outputs(10759) <= not (a and b);
    layer5_outputs(10760) <= not (a and b);
    layer5_outputs(10761) <= not b or a;
    layer5_outputs(10762) <= not a;
    layer5_outputs(10763) <= not a;
    layer5_outputs(10764) <= not a;
    layer5_outputs(10765) <= not a;
    layer5_outputs(10766) <= a or b;
    layer5_outputs(10767) <= not (a or b);
    layer5_outputs(10768) <= a xor b;
    layer5_outputs(10769) <= not (a or b);
    layer5_outputs(10770) <= b;
    layer5_outputs(10771) <= a;
    layer5_outputs(10772) <= not b;
    layer5_outputs(10773) <= not a or b;
    layer5_outputs(10774) <= a or b;
    layer5_outputs(10775) <= not a;
    layer5_outputs(10776) <= b;
    layer5_outputs(10777) <= a;
    layer5_outputs(10778) <= not a or b;
    layer5_outputs(10779) <= b;
    layer5_outputs(10780) <= b;
    layer5_outputs(10781) <= a;
    layer5_outputs(10782) <= a;
    layer5_outputs(10783) <= a xor b;
    layer5_outputs(10784) <= a xor b;
    layer5_outputs(10785) <= a or b;
    layer5_outputs(10786) <= not (a and b);
    layer5_outputs(10787) <= not a or b;
    layer5_outputs(10788) <= not (a xor b);
    layer5_outputs(10789) <= not a;
    layer5_outputs(10790) <= b;
    layer5_outputs(10791) <= not a;
    layer5_outputs(10792) <= not (a or b);
    layer5_outputs(10793) <= not a;
    layer5_outputs(10794) <= a or b;
    layer5_outputs(10795) <= not a;
    layer5_outputs(10796) <= a or b;
    layer5_outputs(10797) <= b;
    layer5_outputs(10798) <= not a or b;
    layer5_outputs(10799) <= not a;
    layer5_outputs(10800) <= not a;
    layer5_outputs(10801) <= not b;
    layer5_outputs(10802) <= not b or a;
    layer5_outputs(10803) <= not a;
    layer5_outputs(10804) <= not a;
    layer5_outputs(10805) <= not (a or b);
    layer5_outputs(10806) <= b;
    layer5_outputs(10807) <= not b or a;
    layer5_outputs(10808) <= a xor b;
    layer5_outputs(10809) <= not b;
    layer5_outputs(10810) <= a;
    layer5_outputs(10811) <= a or b;
    layer5_outputs(10812) <= a and not b;
    layer5_outputs(10813) <= b;
    layer5_outputs(10814) <= not (a or b);
    layer5_outputs(10815) <= a or b;
    layer5_outputs(10816) <= '0';
    layer5_outputs(10817) <= not a;
    layer5_outputs(10818) <= a and not b;
    layer5_outputs(10819) <= a;
    layer5_outputs(10820) <= not b;
    layer5_outputs(10821) <= not b or a;
    layer5_outputs(10822) <= not a;
    layer5_outputs(10823) <= '0';
    layer5_outputs(10824) <= a and b;
    layer5_outputs(10825) <= b and not a;
    layer5_outputs(10826) <= a xor b;
    layer5_outputs(10827) <= b and not a;
    layer5_outputs(10828) <= a xor b;
    layer5_outputs(10829) <= a;
    layer5_outputs(10830) <= b;
    layer5_outputs(10831) <= not b;
    layer5_outputs(10832) <= not a;
    layer5_outputs(10833) <= a;
    layer5_outputs(10834) <= a and not b;
    layer5_outputs(10835) <= a xor b;
    layer5_outputs(10836) <= not b;
    layer5_outputs(10837) <= b;
    layer5_outputs(10838) <= a;
    layer5_outputs(10839) <= not a or b;
    layer5_outputs(10840) <= a;
    layer5_outputs(10841) <= not (a or b);
    layer5_outputs(10842) <= not a;
    layer5_outputs(10843) <= not a;
    layer5_outputs(10844) <= not (a and b);
    layer5_outputs(10845) <= not b or a;
    layer5_outputs(10846) <= not b or a;
    layer5_outputs(10847) <= not (a or b);
    layer5_outputs(10848) <= b and not a;
    layer5_outputs(10849) <= b and not a;
    layer5_outputs(10850) <= not a or b;
    layer5_outputs(10851) <= a;
    layer5_outputs(10852) <= a;
    layer5_outputs(10853) <= b and not a;
    layer5_outputs(10854) <= a and not b;
    layer5_outputs(10855) <= not b;
    layer5_outputs(10856) <= a or b;
    layer5_outputs(10857) <= not (a and b);
    layer5_outputs(10858) <= not b;
    layer5_outputs(10859) <= not (a xor b);
    layer5_outputs(10860) <= not a;
    layer5_outputs(10861) <= a;
    layer5_outputs(10862) <= not a;
    layer5_outputs(10863) <= a;
    layer5_outputs(10864) <= not (a or b);
    layer5_outputs(10865) <= '0';
    layer5_outputs(10866) <= not (a xor b);
    layer5_outputs(10867) <= b;
    layer5_outputs(10868) <= not a;
    layer5_outputs(10869) <= not a;
    layer5_outputs(10870) <= not b;
    layer5_outputs(10871) <= not a or b;
    layer5_outputs(10872) <= not b;
    layer5_outputs(10873) <= a and not b;
    layer5_outputs(10874) <= not b or a;
    layer5_outputs(10875) <= b;
    layer5_outputs(10876) <= not a;
    layer5_outputs(10877) <= b;
    layer5_outputs(10878) <= a xor b;
    layer5_outputs(10879) <= a xor b;
    layer5_outputs(10880) <= '0';
    layer5_outputs(10881) <= b and not a;
    layer5_outputs(10882) <= a;
    layer5_outputs(10883) <= not a;
    layer5_outputs(10884) <= a and not b;
    layer5_outputs(10885) <= not (a or b);
    layer5_outputs(10886) <= not a;
    layer5_outputs(10887) <= b and not a;
    layer5_outputs(10888) <= '0';
    layer5_outputs(10889) <= not a;
    layer5_outputs(10890) <= b and not a;
    layer5_outputs(10891) <= b and not a;
    layer5_outputs(10892) <= a or b;
    layer5_outputs(10893) <= not (a xor b);
    layer5_outputs(10894) <= not a;
    layer5_outputs(10895) <= b and not a;
    layer5_outputs(10896) <= a xor b;
    layer5_outputs(10897) <= a or b;
    layer5_outputs(10898) <= not a;
    layer5_outputs(10899) <= not b or a;
    layer5_outputs(10900) <= not b;
    layer5_outputs(10901) <= a;
    layer5_outputs(10902) <= b and not a;
    layer5_outputs(10903) <= not a;
    layer5_outputs(10904) <= a;
    layer5_outputs(10905) <= not b or a;
    layer5_outputs(10906) <= b;
    layer5_outputs(10907) <= a;
    layer5_outputs(10908) <= a;
    layer5_outputs(10909) <= not (a or b);
    layer5_outputs(10910) <= a xor b;
    layer5_outputs(10911) <= not (a xor b);
    layer5_outputs(10912) <= a and not b;
    layer5_outputs(10913) <= a or b;
    layer5_outputs(10914) <= not (a xor b);
    layer5_outputs(10915) <= not (a and b);
    layer5_outputs(10916) <= not b or a;
    layer5_outputs(10917) <= not (a or b);
    layer5_outputs(10918) <= a and not b;
    layer5_outputs(10919) <= not (a or b);
    layer5_outputs(10920) <= not b or a;
    layer5_outputs(10921) <= not a or b;
    layer5_outputs(10922) <= b;
    layer5_outputs(10923) <= not a;
    layer5_outputs(10924) <= not a or b;
    layer5_outputs(10925) <= not a;
    layer5_outputs(10926) <= not a;
    layer5_outputs(10927) <= not (a or b);
    layer5_outputs(10928) <= not b;
    layer5_outputs(10929) <= not (a xor b);
    layer5_outputs(10930) <= not b or a;
    layer5_outputs(10931) <= not a;
    layer5_outputs(10932) <= a or b;
    layer5_outputs(10933) <= not b;
    layer5_outputs(10934) <= not a;
    layer5_outputs(10935) <= not (a or b);
    layer5_outputs(10936) <= b;
    layer5_outputs(10937) <= b and not a;
    layer5_outputs(10938) <= b;
    layer5_outputs(10939) <= a and b;
    layer5_outputs(10940) <= a or b;
    layer5_outputs(10941) <= not a;
    layer5_outputs(10942) <= a xor b;
    layer5_outputs(10943) <= not a;
    layer5_outputs(10944) <= not b;
    layer5_outputs(10945) <= b;
    layer5_outputs(10946) <= a;
    layer5_outputs(10947) <= not a or b;
    layer5_outputs(10948) <= not a;
    layer5_outputs(10949) <= not a;
    layer5_outputs(10950) <= '1';
    layer5_outputs(10951) <= not a or b;
    layer5_outputs(10952) <= not b;
    layer5_outputs(10953) <= not (a xor b);
    layer5_outputs(10954) <= not b or a;
    layer5_outputs(10955) <= not (a xor b);
    layer5_outputs(10956) <= not (a or b);
    layer5_outputs(10957) <= a and not b;
    layer5_outputs(10958) <= not b;
    layer5_outputs(10959) <= not a;
    layer5_outputs(10960) <= not b;
    layer5_outputs(10961) <= b;
    layer5_outputs(10962) <= a xor b;
    layer5_outputs(10963) <= not a;
    layer5_outputs(10964) <= a xor b;
    layer5_outputs(10965) <= not (a or b);
    layer5_outputs(10966) <= a and not b;
    layer5_outputs(10967) <= not b;
    layer5_outputs(10968) <= not b;
    layer5_outputs(10969) <= b;
    layer5_outputs(10970) <= not b or a;
    layer5_outputs(10971) <= not (a xor b);
    layer5_outputs(10972) <= a xor b;
    layer5_outputs(10973) <= not b;
    layer5_outputs(10974) <= a and not b;
    layer5_outputs(10975) <= a xor b;
    layer5_outputs(10976) <= not (a and b);
    layer5_outputs(10977) <= a;
    layer5_outputs(10978) <= not a or b;
    layer5_outputs(10979) <= not b;
    layer5_outputs(10980) <= a and b;
    layer5_outputs(10981) <= b;
    layer5_outputs(10982) <= not a;
    layer5_outputs(10983) <= not b;
    layer5_outputs(10984) <= '1';
    layer5_outputs(10985) <= a xor b;
    layer5_outputs(10986) <= not a or b;
    layer5_outputs(10987) <= a and b;
    layer5_outputs(10988) <= not (a xor b);
    layer5_outputs(10989) <= not (a or b);
    layer5_outputs(10990) <= not a or b;
    layer5_outputs(10991) <= a xor b;
    layer5_outputs(10992) <= a or b;
    layer5_outputs(10993) <= a and b;
    layer5_outputs(10994) <= a or b;
    layer5_outputs(10995) <= b;
    layer5_outputs(10996) <= b;
    layer5_outputs(10997) <= a and b;
    layer5_outputs(10998) <= a and not b;
    layer5_outputs(10999) <= not a;
    layer5_outputs(11000) <= not a;
    layer5_outputs(11001) <= not b;
    layer5_outputs(11002) <= not (a and b);
    layer5_outputs(11003) <= not b or a;
    layer5_outputs(11004) <= b;
    layer5_outputs(11005) <= not a or b;
    layer5_outputs(11006) <= a and b;
    layer5_outputs(11007) <= not b;
    layer5_outputs(11008) <= not b or a;
    layer5_outputs(11009) <= not (a xor b);
    layer5_outputs(11010) <= not b;
    layer5_outputs(11011) <= not a;
    layer5_outputs(11012) <= b and not a;
    layer5_outputs(11013) <= not b or a;
    layer5_outputs(11014) <= b;
    layer5_outputs(11015) <= a and b;
    layer5_outputs(11016) <= a and b;
    layer5_outputs(11017) <= not (a xor b);
    layer5_outputs(11018) <= not (a xor b);
    layer5_outputs(11019) <= not b;
    layer5_outputs(11020) <= a or b;
    layer5_outputs(11021) <= not b;
    layer5_outputs(11022) <= not a or b;
    layer5_outputs(11023) <= not a or b;
    layer5_outputs(11024) <= a xor b;
    layer5_outputs(11025) <= a or b;
    layer5_outputs(11026) <= not (a and b);
    layer5_outputs(11027) <= b;
    layer5_outputs(11028) <= a or b;
    layer5_outputs(11029) <= not (a and b);
    layer5_outputs(11030) <= not a;
    layer5_outputs(11031) <= not (a xor b);
    layer5_outputs(11032) <= not b or a;
    layer5_outputs(11033) <= not (a and b);
    layer5_outputs(11034) <= not a or b;
    layer5_outputs(11035) <= not a or b;
    layer5_outputs(11036) <= not (a or b);
    layer5_outputs(11037) <= not b;
    layer5_outputs(11038) <= not b;
    layer5_outputs(11039) <= not (a xor b);
    layer5_outputs(11040) <= b;
    layer5_outputs(11041) <= not a;
    layer5_outputs(11042) <= not (a and b);
    layer5_outputs(11043) <= a and b;
    layer5_outputs(11044) <= a or b;
    layer5_outputs(11045) <= a;
    layer5_outputs(11046) <= a;
    layer5_outputs(11047) <= b;
    layer5_outputs(11048) <= not a or b;
    layer5_outputs(11049) <= not a;
    layer5_outputs(11050) <= not (a xor b);
    layer5_outputs(11051) <= b and not a;
    layer5_outputs(11052) <= not (a xor b);
    layer5_outputs(11053) <= not b;
    layer5_outputs(11054) <= not (a or b);
    layer5_outputs(11055) <= a xor b;
    layer5_outputs(11056) <= a xor b;
    layer5_outputs(11057) <= b;
    layer5_outputs(11058) <= not a;
    layer5_outputs(11059) <= not a;
    layer5_outputs(11060) <= a xor b;
    layer5_outputs(11061) <= b and not a;
    layer5_outputs(11062) <= not (a xor b);
    layer5_outputs(11063) <= not a or b;
    layer5_outputs(11064) <= not a;
    layer5_outputs(11065) <= a xor b;
    layer5_outputs(11066) <= not (a xor b);
    layer5_outputs(11067) <= b and not a;
    layer5_outputs(11068) <= b and not a;
    layer5_outputs(11069) <= not a or b;
    layer5_outputs(11070) <= a xor b;
    layer5_outputs(11071) <= a xor b;
    layer5_outputs(11072) <= a and not b;
    layer5_outputs(11073) <= b and not a;
    layer5_outputs(11074) <= a or b;
    layer5_outputs(11075) <= a and b;
    layer5_outputs(11076) <= b;
    layer5_outputs(11077) <= a and b;
    layer5_outputs(11078) <= not a;
    layer5_outputs(11079) <= a;
    layer5_outputs(11080) <= not (a or b);
    layer5_outputs(11081) <= a;
    layer5_outputs(11082) <= not b;
    layer5_outputs(11083) <= a;
    layer5_outputs(11084) <= not (a and b);
    layer5_outputs(11085) <= not b;
    layer5_outputs(11086) <= b;
    layer5_outputs(11087) <= a xor b;
    layer5_outputs(11088) <= not a or b;
    layer5_outputs(11089) <= not (a xor b);
    layer5_outputs(11090) <= a or b;
    layer5_outputs(11091) <= '0';
    layer5_outputs(11092) <= not (a xor b);
    layer5_outputs(11093) <= a xor b;
    layer5_outputs(11094) <= b and not a;
    layer5_outputs(11095) <= a or b;
    layer5_outputs(11096) <= a;
    layer5_outputs(11097) <= a and b;
    layer5_outputs(11098) <= b and not a;
    layer5_outputs(11099) <= not b;
    layer5_outputs(11100) <= not (a or b);
    layer5_outputs(11101) <= not (a and b);
    layer5_outputs(11102) <= a;
    layer5_outputs(11103) <= not (a xor b);
    layer5_outputs(11104) <= a or b;
    layer5_outputs(11105) <= not b or a;
    layer5_outputs(11106) <= not b or a;
    layer5_outputs(11107) <= not (a xor b);
    layer5_outputs(11108) <= not (a xor b);
    layer5_outputs(11109) <= a;
    layer5_outputs(11110) <= not (a or b);
    layer5_outputs(11111) <= b;
    layer5_outputs(11112) <= a xor b;
    layer5_outputs(11113) <= not b or a;
    layer5_outputs(11114) <= a xor b;
    layer5_outputs(11115) <= not (a or b);
    layer5_outputs(11116) <= a and b;
    layer5_outputs(11117) <= a and not b;
    layer5_outputs(11118) <= not b;
    layer5_outputs(11119) <= not b;
    layer5_outputs(11120) <= a xor b;
    layer5_outputs(11121) <= not (a and b);
    layer5_outputs(11122) <= a xor b;
    layer5_outputs(11123) <= a and not b;
    layer5_outputs(11124) <= not b;
    layer5_outputs(11125) <= b;
    layer5_outputs(11126) <= '0';
    layer5_outputs(11127) <= b;
    layer5_outputs(11128) <= a and b;
    layer5_outputs(11129) <= '1';
    layer5_outputs(11130) <= a and b;
    layer5_outputs(11131) <= a xor b;
    layer5_outputs(11132) <= b and not a;
    layer5_outputs(11133) <= not a;
    layer5_outputs(11134) <= b and not a;
    layer5_outputs(11135) <= not a;
    layer5_outputs(11136) <= not b;
    layer5_outputs(11137) <= b;
    layer5_outputs(11138) <= not b;
    layer5_outputs(11139) <= not b;
    layer5_outputs(11140) <= b;
    layer5_outputs(11141) <= not b;
    layer5_outputs(11142) <= a xor b;
    layer5_outputs(11143) <= b;
    layer5_outputs(11144) <= b;
    layer5_outputs(11145) <= not a;
    layer5_outputs(11146) <= not b;
    layer5_outputs(11147) <= a;
    layer5_outputs(11148) <= not (a and b);
    layer5_outputs(11149) <= not a;
    layer5_outputs(11150) <= a;
    layer5_outputs(11151) <= b;
    layer5_outputs(11152) <= b;
    layer5_outputs(11153) <= a and b;
    layer5_outputs(11154) <= a and not b;
    layer5_outputs(11155) <= a and not b;
    layer5_outputs(11156) <= a and not b;
    layer5_outputs(11157) <= a and not b;
    layer5_outputs(11158) <= not (a or b);
    layer5_outputs(11159) <= a or b;
    layer5_outputs(11160) <= not a;
    layer5_outputs(11161) <= not (a or b);
    layer5_outputs(11162) <= not b or a;
    layer5_outputs(11163) <= '0';
    layer5_outputs(11164) <= a or b;
    layer5_outputs(11165) <= not a;
    layer5_outputs(11166) <= a or b;
    layer5_outputs(11167) <= not (a xor b);
    layer5_outputs(11168) <= a xor b;
    layer5_outputs(11169) <= not (a or b);
    layer5_outputs(11170) <= not (a xor b);
    layer5_outputs(11171) <= not (a or b);
    layer5_outputs(11172) <= not (a or b);
    layer5_outputs(11173) <= not b;
    layer5_outputs(11174) <= a;
    layer5_outputs(11175) <= not (a and b);
    layer5_outputs(11176) <= a;
    layer5_outputs(11177) <= not (a xor b);
    layer5_outputs(11178) <= not b or a;
    layer5_outputs(11179) <= b;
    layer5_outputs(11180) <= not a;
    layer5_outputs(11181) <= not a;
    layer5_outputs(11182) <= a and b;
    layer5_outputs(11183) <= not (a and b);
    layer5_outputs(11184) <= a xor b;
    layer5_outputs(11185) <= a and not b;
    layer5_outputs(11186) <= a xor b;
    layer5_outputs(11187) <= not a;
    layer5_outputs(11188) <= b;
    layer5_outputs(11189) <= a;
    layer5_outputs(11190) <= not a;
    layer5_outputs(11191) <= b and not a;
    layer5_outputs(11192) <= not (a and b);
    layer5_outputs(11193) <= not b or a;
    layer5_outputs(11194) <= a and not b;
    layer5_outputs(11195) <= not b;
    layer5_outputs(11196) <= not a;
    layer5_outputs(11197) <= a xor b;
    layer5_outputs(11198) <= not b;
    layer5_outputs(11199) <= a and not b;
    layer5_outputs(11200) <= not b;
    layer5_outputs(11201) <= not (a xor b);
    layer5_outputs(11202) <= not (a or b);
    layer5_outputs(11203) <= not (a and b);
    layer5_outputs(11204) <= b;
    layer5_outputs(11205) <= not (a or b);
    layer5_outputs(11206) <= not (a xor b);
    layer5_outputs(11207) <= a;
    layer5_outputs(11208) <= not (a xor b);
    layer5_outputs(11209) <= not (a xor b);
    layer5_outputs(11210) <= b and not a;
    layer5_outputs(11211) <= b;
    layer5_outputs(11212) <= a;
    layer5_outputs(11213) <= a;
    layer5_outputs(11214) <= not a;
    layer5_outputs(11215) <= a xor b;
    layer5_outputs(11216) <= not b;
    layer5_outputs(11217) <= b;
    layer5_outputs(11218) <= a xor b;
    layer5_outputs(11219) <= a;
    layer5_outputs(11220) <= not a or b;
    layer5_outputs(11221) <= not a;
    layer5_outputs(11222) <= not (a and b);
    layer5_outputs(11223) <= not b;
    layer5_outputs(11224) <= b;
    layer5_outputs(11225) <= a or b;
    layer5_outputs(11226) <= b;
    layer5_outputs(11227) <= not a or b;
    layer5_outputs(11228) <= not (a or b);
    layer5_outputs(11229) <= a or b;
    layer5_outputs(11230) <= a;
    layer5_outputs(11231) <= b and not a;
    layer5_outputs(11232) <= not a;
    layer5_outputs(11233) <= a;
    layer5_outputs(11234) <= not (a and b);
    layer5_outputs(11235) <= not a;
    layer5_outputs(11236) <= not a;
    layer5_outputs(11237) <= not a or b;
    layer5_outputs(11238) <= b;
    layer5_outputs(11239) <= not a or b;
    layer5_outputs(11240) <= not b or a;
    layer5_outputs(11241) <= b;
    layer5_outputs(11242) <= a or b;
    layer5_outputs(11243) <= not b;
    layer5_outputs(11244) <= not (a and b);
    layer5_outputs(11245) <= not (a xor b);
    layer5_outputs(11246) <= a and b;
    layer5_outputs(11247) <= a or b;
    layer5_outputs(11248) <= not b;
    layer5_outputs(11249) <= a;
    layer5_outputs(11250) <= a xor b;
    layer5_outputs(11251) <= not (a and b);
    layer5_outputs(11252) <= not b;
    layer5_outputs(11253) <= a xor b;
    layer5_outputs(11254) <= not b;
    layer5_outputs(11255) <= not (a xor b);
    layer5_outputs(11256) <= not b;
    layer5_outputs(11257) <= b;
    layer5_outputs(11258) <= not a;
    layer5_outputs(11259) <= not (a xor b);
    layer5_outputs(11260) <= a xor b;
    layer5_outputs(11261) <= a and b;
    layer5_outputs(11262) <= b;
    layer5_outputs(11263) <= b;
    layer5_outputs(11264) <= b;
    layer5_outputs(11265) <= not (a or b);
    layer5_outputs(11266) <= a or b;
    layer5_outputs(11267) <= not (a and b);
    layer5_outputs(11268) <= not (a xor b);
    layer5_outputs(11269) <= not b or a;
    layer5_outputs(11270) <= not (a and b);
    layer5_outputs(11271) <= a and b;
    layer5_outputs(11272) <= b;
    layer5_outputs(11273) <= not (a xor b);
    layer5_outputs(11274) <= b and not a;
    layer5_outputs(11275) <= a xor b;
    layer5_outputs(11276) <= not b;
    layer5_outputs(11277) <= not a;
    layer5_outputs(11278) <= b;
    layer5_outputs(11279) <= b and not a;
    layer5_outputs(11280) <= b;
    layer5_outputs(11281) <= a and b;
    layer5_outputs(11282) <= b;
    layer5_outputs(11283) <= not b;
    layer5_outputs(11284) <= not a;
    layer5_outputs(11285) <= not (a or b);
    layer5_outputs(11286) <= not b or a;
    layer5_outputs(11287) <= not a;
    layer5_outputs(11288) <= not b;
    layer5_outputs(11289) <= a or b;
    layer5_outputs(11290) <= a and not b;
    layer5_outputs(11291) <= a xor b;
    layer5_outputs(11292) <= a;
    layer5_outputs(11293) <= not a;
    layer5_outputs(11294) <= not b;
    layer5_outputs(11295) <= not (a or b);
    layer5_outputs(11296) <= not (a or b);
    layer5_outputs(11297) <= a xor b;
    layer5_outputs(11298) <= b;
    layer5_outputs(11299) <= a and not b;
    layer5_outputs(11300) <= not b or a;
    layer5_outputs(11301) <= not a;
    layer5_outputs(11302) <= a and b;
    layer5_outputs(11303) <= '0';
    layer5_outputs(11304) <= not a;
    layer5_outputs(11305) <= b and not a;
    layer5_outputs(11306) <= a or b;
    layer5_outputs(11307) <= not b or a;
    layer5_outputs(11308) <= a xor b;
    layer5_outputs(11309) <= not a;
    layer5_outputs(11310) <= not (a and b);
    layer5_outputs(11311) <= not b;
    layer5_outputs(11312) <= b and not a;
    layer5_outputs(11313) <= a;
    layer5_outputs(11314) <= not (a xor b);
    layer5_outputs(11315) <= not b or a;
    layer5_outputs(11316) <= a or b;
    layer5_outputs(11317) <= not a or b;
    layer5_outputs(11318) <= not b or a;
    layer5_outputs(11319) <= a;
    layer5_outputs(11320) <= not b;
    layer5_outputs(11321) <= not b or a;
    layer5_outputs(11322) <= not (a and b);
    layer5_outputs(11323) <= a or b;
    layer5_outputs(11324) <= not b or a;
    layer5_outputs(11325) <= b and not a;
    layer5_outputs(11326) <= a and b;
    layer5_outputs(11327) <= a xor b;
    layer5_outputs(11328) <= a or b;
    layer5_outputs(11329) <= not (a or b);
    layer5_outputs(11330) <= not b;
    layer5_outputs(11331) <= not a;
    layer5_outputs(11332) <= a and not b;
    layer5_outputs(11333) <= not (a or b);
    layer5_outputs(11334) <= not b;
    layer5_outputs(11335) <= not a;
    layer5_outputs(11336) <= not (a xor b);
    layer5_outputs(11337) <= a;
    layer5_outputs(11338) <= a and not b;
    layer5_outputs(11339) <= not b or a;
    layer5_outputs(11340) <= not (a or b);
    layer5_outputs(11341) <= not (a xor b);
    layer5_outputs(11342) <= a or b;
    layer5_outputs(11343) <= not b;
    layer5_outputs(11344) <= not b or a;
    layer5_outputs(11345) <= not b;
    layer5_outputs(11346) <= not b;
    layer5_outputs(11347) <= not (a and b);
    layer5_outputs(11348) <= a;
    layer5_outputs(11349) <= b;
    layer5_outputs(11350) <= a and b;
    layer5_outputs(11351) <= not b or a;
    layer5_outputs(11352) <= not a;
    layer5_outputs(11353) <= a;
    layer5_outputs(11354) <= a;
    layer5_outputs(11355) <= not (a or b);
    layer5_outputs(11356) <= a and not b;
    layer5_outputs(11357) <= not (a or b);
    layer5_outputs(11358) <= not a or b;
    layer5_outputs(11359) <= b and not a;
    layer5_outputs(11360) <= not b;
    layer5_outputs(11361) <= a;
    layer5_outputs(11362) <= not a;
    layer5_outputs(11363) <= not b;
    layer5_outputs(11364) <= not b;
    layer5_outputs(11365) <= not b;
    layer5_outputs(11366) <= not b;
    layer5_outputs(11367) <= b;
    layer5_outputs(11368) <= b;
    layer5_outputs(11369) <= a;
    layer5_outputs(11370) <= a;
    layer5_outputs(11371) <= not a;
    layer5_outputs(11372) <= b;
    layer5_outputs(11373) <= not (a xor b);
    layer5_outputs(11374) <= b;
    layer5_outputs(11375) <= b and not a;
    layer5_outputs(11376) <= a;
    layer5_outputs(11377) <= not a or b;
    layer5_outputs(11378) <= not a;
    layer5_outputs(11379) <= not b or a;
    layer5_outputs(11380) <= not (a and b);
    layer5_outputs(11381) <= not (a xor b);
    layer5_outputs(11382) <= '1';
    layer5_outputs(11383) <= not b;
    layer5_outputs(11384) <= b;
    layer5_outputs(11385) <= not a;
    layer5_outputs(11386) <= not (a xor b);
    layer5_outputs(11387) <= not b;
    layer5_outputs(11388) <= not a;
    layer5_outputs(11389) <= not a;
    layer5_outputs(11390) <= a and b;
    layer5_outputs(11391) <= not a;
    layer5_outputs(11392) <= b;
    layer5_outputs(11393) <= not a;
    layer5_outputs(11394) <= a;
    layer5_outputs(11395) <= not b or a;
    layer5_outputs(11396) <= not b or a;
    layer5_outputs(11397) <= not (a and b);
    layer5_outputs(11398) <= a or b;
    layer5_outputs(11399) <= a or b;
    layer5_outputs(11400) <= not (a or b);
    layer5_outputs(11401) <= a and not b;
    layer5_outputs(11402) <= not (a or b);
    layer5_outputs(11403) <= a xor b;
    layer5_outputs(11404) <= not b or a;
    layer5_outputs(11405) <= a xor b;
    layer5_outputs(11406) <= b;
    layer5_outputs(11407) <= a or b;
    layer5_outputs(11408) <= b;
    layer5_outputs(11409) <= a and b;
    layer5_outputs(11410) <= not b or a;
    layer5_outputs(11411) <= a;
    layer5_outputs(11412) <= not a;
    layer5_outputs(11413) <= a;
    layer5_outputs(11414) <= a xor b;
    layer5_outputs(11415) <= a and b;
    layer5_outputs(11416) <= b;
    layer5_outputs(11417) <= not a or b;
    layer5_outputs(11418) <= not b;
    layer5_outputs(11419) <= b;
    layer5_outputs(11420) <= b;
    layer5_outputs(11421) <= a xor b;
    layer5_outputs(11422) <= a xor b;
    layer5_outputs(11423) <= not a;
    layer5_outputs(11424) <= not (a and b);
    layer5_outputs(11425) <= a xor b;
    layer5_outputs(11426) <= a and b;
    layer5_outputs(11427) <= b;
    layer5_outputs(11428) <= b and not a;
    layer5_outputs(11429) <= a xor b;
    layer5_outputs(11430) <= a or b;
    layer5_outputs(11431) <= a and b;
    layer5_outputs(11432) <= a xor b;
    layer5_outputs(11433) <= not a;
    layer5_outputs(11434) <= not a;
    layer5_outputs(11435) <= a;
    layer5_outputs(11436) <= b;
    layer5_outputs(11437) <= not b or a;
    layer5_outputs(11438) <= '0';
    layer5_outputs(11439) <= b;
    layer5_outputs(11440) <= b;
    layer5_outputs(11441) <= b;
    layer5_outputs(11442) <= a and not b;
    layer5_outputs(11443) <= a;
    layer5_outputs(11444) <= a;
    layer5_outputs(11445) <= not a;
    layer5_outputs(11446) <= a and b;
    layer5_outputs(11447) <= not b;
    layer5_outputs(11448) <= not a or b;
    layer5_outputs(11449) <= a;
    layer5_outputs(11450) <= a or b;
    layer5_outputs(11451) <= a and b;
    layer5_outputs(11452) <= not (a xor b);
    layer5_outputs(11453) <= a;
    layer5_outputs(11454) <= not b;
    layer5_outputs(11455) <= b and not a;
    layer5_outputs(11456) <= not (a or b);
    layer5_outputs(11457) <= not b or a;
    layer5_outputs(11458) <= a or b;
    layer5_outputs(11459) <= a;
    layer5_outputs(11460) <= b;
    layer5_outputs(11461) <= not (a xor b);
    layer5_outputs(11462) <= not (a xor b);
    layer5_outputs(11463) <= not a;
    layer5_outputs(11464) <= a and b;
    layer5_outputs(11465) <= not (a or b);
    layer5_outputs(11466) <= a xor b;
    layer5_outputs(11467) <= not b or a;
    layer5_outputs(11468) <= a or b;
    layer5_outputs(11469) <= not b;
    layer5_outputs(11470) <= not b;
    layer5_outputs(11471) <= a or b;
    layer5_outputs(11472) <= not (a xor b);
    layer5_outputs(11473) <= a;
    layer5_outputs(11474) <= not b or a;
    layer5_outputs(11475) <= a;
    layer5_outputs(11476) <= not (a xor b);
    layer5_outputs(11477) <= not a;
    layer5_outputs(11478) <= not a or b;
    layer5_outputs(11479) <= b;
    layer5_outputs(11480) <= a;
    layer5_outputs(11481) <= a or b;
    layer5_outputs(11482) <= not (a xor b);
    layer5_outputs(11483) <= b and not a;
    layer5_outputs(11484) <= a and not b;
    layer5_outputs(11485) <= '0';
    layer5_outputs(11486) <= a;
    layer5_outputs(11487) <= a xor b;
    layer5_outputs(11488) <= a xor b;
    layer5_outputs(11489) <= a;
    layer5_outputs(11490) <= b and not a;
    layer5_outputs(11491) <= a xor b;
    layer5_outputs(11492) <= a;
    layer5_outputs(11493) <= a and b;
    layer5_outputs(11494) <= a or b;
    layer5_outputs(11495) <= b;
    layer5_outputs(11496) <= not b or a;
    layer5_outputs(11497) <= not b or a;
    layer5_outputs(11498) <= a;
    layer5_outputs(11499) <= not (a xor b);
    layer5_outputs(11500) <= b;
    layer5_outputs(11501) <= not a;
    layer5_outputs(11502) <= a or b;
    layer5_outputs(11503) <= not b or a;
    layer5_outputs(11504) <= not a;
    layer5_outputs(11505) <= not b or a;
    layer5_outputs(11506) <= a and not b;
    layer5_outputs(11507) <= not (a and b);
    layer5_outputs(11508) <= a;
    layer5_outputs(11509) <= not b;
    layer5_outputs(11510) <= a;
    layer5_outputs(11511) <= b and not a;
    layer5_outputs(11512) <= not (a xor b);
    layer5_outputs(11513) <= a xor b;
    layer5_outputs(11514) <= b and not a;
    layer5_outputs(11515) <= not (a or b);
    layer5_outputs(11516) <= not a or b;
    layer5_outputs(11517) <= not (a or b);
    layer5_outputs(11518) <= a and not b;
    layer5_outputs(11519) <= not b;
    layer5_outputs(11520) <= not a;
    layer5_outputs(11521) <= not a or b;
    layer5_outputs(11522) <= '1';
    layer5_outputs(11523) <= not b or a;
    layer5_outputs(11524) <= not b;
    layer5_outputs(11525) <= a and not b;
    layer5_outputs(11526) <= a;
    layer5_outputs(11527) <= a and b;
    layer5_outputs(11528) <= not (a or b);
    layer5_outputs(11529) <= a and not b;
    layer5_outputs(11530) <= a and not b;
    layer5_outputs(11531) <= '1';
    layer5_outputs(11532) <= a xor b;
    layer5_outputs(11533) <= a xor b;
    layer5_outputs(11534) <= not a;
    layer5_outputs(11535) <= not b;
    layer5_outputs(11536) <= not b or a;
    layer5_outputs(11537) <= not a;
    layer5_outputs(11538) <= b;
    layer5_outputs(11539) <= not (a or b);
    layer5_outputs(11540) <= not (a or b);
    layer5_outputs(11541) <= b;
    layer5_outputs(11542) <= b;
    layer5_outputs(11543) <= a or b;
    layer5_outputs(11544) <= a;
    layer5_outputs(11545) <= not a;
    layer5_outputs(11546) <= not (a or b);
    layer5_outputs(11547) <= b;
    layer5_outputs(11548) <= not b;
    layer5_outputs(11549) <= b;
    layer5_outputs(11550) <= not b or a;
    layer5_outputs(11551) <= a xor b;
    layer5_outputs(11552) <= b;
    layer5_outputs(11553) <= b and not a;
    layer5_outputs(11554) <= a and b;
    layer5_outputs(11555) <= a and b;
    layer5_outputs(11556) <= b;
    layer5_outputs(11557) <= a or b;
    layer5_outputs(11558) <= b;
    layer5_outputs(11559) <= b;
    layer5_outputs(11560) <= a and not b;
    layer5_outputs(11561) <= b and not a;
    layer5_outputs(11562) <= a and not b;
    layer5_outputs(11563) <= a and b;
    layer5_outputs(11564) <= not a or b;
    layer5_outputs(11565) <= not (a xor b);
    layer5_outputs(11566) <= a xor b;
    layer5_outputs(11567) <= a;
    layer5_outputs(11568) <= b;
    layer5_outputs(11569) <= not (a xor b);
    layer5_outputs(11570) <= not (a and b);
    layer5_outputs(11571) <= not b;
    layer5_outputs(11572) <= b;
    layer5_outputs(11573) <= not b or a;
    layer5_outputs(11574) <= '0';
    layer5_outputs(11575) <= not a;
    layer5_outputs(11576) <= not b;
    layer5_outputs(11577) <= not (a xor b);
    layer5_outputs(11578) <= a;
    layer5_outputs(11579) <= a;
    layer5_outputs(11580) <= b and not a;
    layer5_outputs(11581) <= not a;
    layer5_outputs(11582) <= not b or a;
    layer5_outputs(11583) <= a;
    layer5_outputs(11584) <= not b;
    layer5_outputs(11585) <= '0';
    layer5_outputs(11586) <= a and b;
    layer5_outputs(11587) <= not b;
    layer5_outputs(11588) <= not b;
    layer5_outputs(11589) <= a;
    layer5_outputs(11590) <= not b;
    layer5_outputs(11591) <= not (a and b);
    layer5_outputs(11592) <= not a or b;
    layer5_outputs(11593) <= not a;
    layer5_outputs(11594) <= a and b;
    layer5_outputs(11595) <= not (a xor b);
    layer5_outputs(11596) <= not (a and b);
    layer5_outputs(11597) <= not (a xor b);
    layer5_outputs(11598) <= not a or b;
    layer5_outputs(11599) <= not (a or b);
    layer5_outputs(11600) <= b and not a;
    layer5_outputs(11601) <= a and not b;
    layer5_outputs(11602) <= not (a xor b);
    layer5_outputs(11603) <= not a;
    layer5_outputs(11604) <= not a or b;
    layer5_outputs(11605) <= a and not b;
    layer5_outputs(11606) <= not a;
    layer5_outputs(11607) <= a or b;
    layer5_outputs(11608) <= not (a xor b);
    layer5_outputs(11609) <= not (a and b);
    layer5_outputs(11610) <= a and not b;
    layer5_outputs(11611) <= not a;
    layer5_outputs(11612) <= a or b;
    layer5_outputs(11613) <= not b;
    layer5_outputs(11614) <= not (a or b);
    layer5_outputs(11615) <= a and b;
    layer5_outputs(11616) <= a xor b;
    layer5_outputs(11617) <= not a or b;
    layer5_outputs(11618) <= a;
    layer5_outputs(11619) <= not (a or b);
    layer5_outputs(11620) <= a and b;
    layer5_outputs(11621) <= not (a and b);
    layer5_outputs(11622) <= a xor b;
    layer5_outputs(11623) <= b;
    layer5_outputs(11624) <= b and not a;
    layer5_outputs(11625) <= not b or a;
    layer5_outputs(11626) <= b;
    layer5_outputs(11627) <= not (a xor b);
    layer5_outputs(11628) <= not (a and b);
    layer5_outputs(11629) <= not a or b;
    layer5_outputs(11630) <= not (a xor b);
    layer5_outputs(11631) <= b and not a;
    layer5_outputs(11632) <= not b or a;
    layer5_outputs(11633) <= a;
    layer5_outputs(11634) <= not b;
    layer5_outputs(11635) <= a;
    layer5_outputs(11636) <= not a;
    layer5_outputs(11637) <= a xor b;
    layer5_outputs(11638) <= b and not a;
    layer5_outputs(11639) <= not (a and b);
    layer5_outputs(11640) <= not b or a;
    layer5_outputs(11641) <= a and not b;
    layer5_outputs(11642) <= a xor b;
    layer5_outputs(11643) <= a or b;
    layer5_outputs(11644) <= not a or b;
    layer5_outputs(11645) <= a;
    layer5_outputs(11646) <= not a;
    layer5_outputs(11647) <= not (a xor b);
    layer5_outputs(11648) <= a and b;
    layer5_outputs(11649) <= not b;
    layer5_outputs(11650) <= not a;
    layer5_outputs(11651) <= not (a and b);
    layer5_outputs(11652) <= b;
    layer5_outputs(11653) <= not b;
    layer5_outputs(11654) <= not b;
    layer5_outputs(11655) <= not (a xor b);
    layer5_outputs(11656) <= not b;
    layer5_outputs(11657) <= not b;
    layer5_outputs(11658) <= not b;
    layer5_outputs(11659) <= a;
    layer5_outputs(11660) <= a;
    layer5_outputs(11661) <= not (a xor b);
    layer5_outputs(11662) <= not a or b;
    layer5_outputs(11663) <= not (a xor b);
    layer5_outputs(11664) <= not b;
    layer5_outputs(11665) <= not a;
    layer5_outputs(11666) <= not b;
    layer5_outputs(11667) <= b;
    layer5_outputs(11668) <= not b;
    layer5_outputs(11669) <= b;
    layer5_outputs(11670) <= not a or b;
    layer5_outputs(11671) <= b;
    layer5_outputs(11672) <= a and b;
    layer5_outputs(11673) <= not b;
    layer5_outputs(11674) <= not (a or b);
    layer5_outputs(11675) <= a xor b;
    layer5_outputs(11676) <= a;
    layer5_outputs(11677) <= not a or b;
    layer5_outputs(11678) <= a and not b;
    layer5_outputs(11679) <= not (a xor b);
    layer5_outputs(11680) <= a or b;
    layer5_outputs(11681) <= not b;
    layer5_outputs(11682) <= not b or a;
    layer5_outputs(11683) <= a or b;
    layer5_outputs(11684) <= a xor b;
    layer5_outputs(11685) <= b;
    layer5_outputs(11686) <= a xor b;
    layer5_outputs(11687) <= not a or b;
    layer5_outputs(11688) <= a or b;
    layer5_outputs(11689) <= a;
    layer5_outputs(11690) <= a xor b;
    layer5_outputs(11691) <= a xor b;
    layer5_outputs(11692) <= a or b;
    layer5_outputs(11693) <= b and not a;
    layer5_outputs(11694) <= b;
    layer5_outputs(11695) <= b and not a;
    layer5_outputs(11696) <= not (a or b);
    layer5_outputs(11697) <= not b;
    layer5_outputs(11698) <= not a;
    layer5_outputs(11699) <= a;
    layer5_outputs(11700) <= a or b;
    layer5_outputs(11701) <= not a;
    layer5_outputs(11702) <= b;
    layer5_outputs(11703) <= b;
    layer5_outputs(11704) <= a xor b;
    layer5_outputs(11705) <= a or b;
    layer5_outputs(11706) <= not (a xor b);
    layer5_outputs(11707) <= a;
    layer5_outputs(11708) <= a;
    layer5_outputs(11709) <= not a;
    layer5_outputs(11710) <= b;
    layer5_outputs(11711) <= a;
    layer5_outputs(11712) <= a and b;
    layer5_outputs(11713) <= not (a xor b);
    layer5_outputs(11714) <= b;
    layer5_outputs(11715) <= a;
    layer5_outputs(11716) <= not b or a;
    layer5_outputs(11717) <= a;
    layer5_outputs(11718) <= a and b;
    layer5_outputs(11719) <= a and not b;
    layer5_outputs(11720) <= a;
    layer5_outputs(11721) <= not b or a;
    layer5_outputs(11722) <= not b;
    layer5_outputs(11723) <= not b;
    layer5_outputs(11724) <= '1';
    layer5_outputs(11725) <= a xor b;
    layer5_outputs(11726) <= not b;
    layer5_outputs(11727) <= a and not b;
    layer5_outputs(11728) <= not a;
    layer5_outputs(11729) <= not (a and b);
    layer5_outputs(11730) <= not a;
    layer5_outputs(11731) <= not b or a;
    layer5_outputs(11732) <= not b;
    layer5_outputs(11733) <= a xor b;
    layer5_outputs(11734) <= a xor b;
    layer5_outputs(11735) <= a;
    layer5_outputs(11736) <= not a;
    layer5_outputs(11737) <= not (a or b);
    layer5_outputs(11738) <= not a;
    layer5_outputs(11739) <= not (a and b);
    layer5_outputs(11740) <= a and b;
    layer5_outputs(11741) <= b;
    layer5_outputs(11742) <= not a;
    layer5_outputs(11743) <= a;
    layer5_outputs(11744) <= not (a or b);
    layer5_outputs(11745) <= not b;
    layer5_outputs(11746) <= b;
    layer5_outputs(11747) <= b;
    layer5_outputs(11748) <= not (a or b);
    layer5_outputs(11749) <= b;
    layer5_outputs(11750) <= a;
    layer5_outputs(11751) <= not a or b;
    layer5_outputs(11752) <= not (a and b);
    layer5_outputs(11753) <= not a;
    layer5_outputs(11754) <= '1';
    layer5_outputs(11755) <= a xor b;
    layer5_outputs(11756) <= not b;
    layer5_outputs(11757) <= not a;
    layer5_outputs(11758) <= not (a or b);
    layer5_outputs(11759) <= not b;
    layer5_outputs(11760) <= a and not b;
    layer5_outputs(11761) <= a xor b;
    layer5_outputs(11762) <= not b or a;
    layer5_outputs(11763) <= not b;
    layer5_outputs(11764) <= not b;
    layer5_outputs(11765) <= not b or a;
    layer5_outputs(11766) <= a or b;
    layer5_outputs(11767) <= b and not a;
    layer5_outputs(11768) <= not b;
    layer5_outputs(11769) <= a or b;
    layer5_outputs(11770) <= a or b;
    layer5_outputs(11771) <= b;
    layer5_outputs(11772) <= a;
    layer5_outputs(11773) <= b;
    layer5_outputs(11774) <= b;
    layer5_outputs(11775) <= not (a xor b);
    layer5_outputs(11776) <= a;
    layer5_outputs(11777) <= b;
    layer5_outputs(11778) <= not (a or b);
    layer5_outputs(11779) <= a xor b;
    layer5_outputs(11780) <= a;
    layer5_outputs(11781) <= b;
    layer5_outputs(11782) <= not (a xor b);
    layer5_outputs(11783) <= not b or a;
    layer5_outputs(11784) <= not b;
    layer5_outputs(11785) <= b;
    layer5_outputs(11786) <= a and not b;
    layer5_outputs(11787) <= b;
    layer5_outputs(11788) <= a;
    layer5_outputs(11789) <= not b;
    layer5_outputs(11790) <= '1';
    layer5_outputs(11791) <= '1';
    layer5_outputs(11792) <= b and not a;
    layer5_outputs(11793) <= not b or a;
    layer5_outputs(11794) <= not b;
    layer5_outputs(11795) <= not (a or b);
    layer5_outputs(11796) <= not a;
    layer5_outputs(11797) <= a;
    layer5_outputs(11798) <= not a;
    layer5_outputs(11799) <= not a or b;
    layer5_outputs(11800) <= b;
    layer5_outputs(11801) <= not b or a;
    layer5_outputs(11802) <= not a;
    layer5_outputs(11803) <= not b;
    layer5_outputs(11804) <= not a;
    layer5_outputs(11805) <= a and not b;
    layer5_outputs(11806) <= b;
    layer5_outputs(11807) <= not (a xor b);
    layer5_outputs(11808) <= b;
    layer5_outputs(11809) <= not a or b;
    layer5_outputs(11810) <= b;
    layer5_outputs(11811) <= not (a xor b);
    layer5_outputs(11812) <= not (a xor b);
    layer5_outputs(11813) <= not (a xor b);
    layer5_outputs(11814) <= a and b;
    layer5_outputs(11815) <= not (a xor b);
    layer5_outputs(11816) <= not b;
    layer5_outputs(11817) <= '1';
    layer5_outputs(11818) <= not a;
    layer5_outputs(11819) <= not (a or b);
    layer5_outputs(11820) <= b;
    layer5_outputs(11821) <= '1';
    layer5_outputs(11822) <= not a or b;
    layer5_outputs(11823) <= not (a xor b);
    layer5_outputs(11824) <= not b or a;
    layer5_outputs(11825) <= not b;
    layer5_outputs(11826) <= b;
    layer5_outputs(11827) <= a;
    layer5_outputs(11828) <= a;
    layer5_outputs(11829) <= not a;
    layer5_outputs(11830) <= b;
    layer5_outputs(11831) <= a and b;
    layer5_outputs(11832) <= b and not a;
    layer5_outputs(11833) <= b;
    layer5_outputs(11834) <= not b;
    layer5_outputs(11835) <= not (a or b);
    layer5_outputs(11836) <= not b or a;
    layer5_outputs(11837) <= not a;
    layer5_outputs(11838) <= not a;
    layer5_outputs(11839) <= not (a or b);
    layer5_outputs(11840) <= not (a or b);
    layer5_outputs(11841) <= not a;
    layer5_outputs(11842) <= b;
    layer5_outputs(11843) <= a or b;
    layer5_outputs(11844) <= not (a and b);
    layer5_outputs(11845) <= a;
    layer5_outputs(11846) <= b;
    layer5_outputs(11847) <= not a;
    layer5_outputs(11848) <= a;
    layer5_outputs(11849) <= not (a xor b);
    layer5_outputs(11850) <= b;
    layer5_outputs(11851) <= not b;
    layer5_outputs(11852) <= a xor b;
    layer5_outputs(11853) <= a and b;
    layer5_outputs(11854) <= not a or b;
    layer5_outputs(11855) <= a and not b;
    layer5_outputs(11856) <= not b;
    layer5_outputs(11857) <= not a;
    layer5_outputs(11858) <= not a;
    layer5_outputs(11859) <= a;
    layer5_outputs(11860) <= a xor b;
    layer5_outputs(11861) <= '0';
    layer5_outputs(11862) <= b;
    layer5_outputs(11863) <= not a;
    layer5_outputs(11864) <= not a;
    layer5_outputs(11865) <= not b;
    layer5_outputs(11866) <= not (a xor b);
    layer5_outputs(11867) <= a;
    layer5_outputs(11868) <= not a or b;
    layer5_outputs(11869) <= not (a and b);
    layer5_outputs(11870) <= not (a or b);
    layer5_outputs(11871) <= not a;
    layer5_outputs(11872) <= a;
    layer5_outputs(11873) <= not (a or b);
    layer5_outputs(11874) <= not a or b;
    layer5_outputs(11875) <= not (a or b);
    layer5_outputs(11876) <= not a or b;
    layer5_outputs(11877) <= a;
    layer5_outputs(11878) <= not a;
    layer5_outputs(11879) <= not (a and b);
    layer5_outputs(11880) <= b;
    layer5_outputs(11881) <= a;
    layer5_outputs(11882) <= b;
    layer5_outputs(11883) <= a and not b;
    layer5_outputs(11884) <= not (a xor b);
    layer5_outputs(11885) <= not b;
    layer5_outputs(11886) <= a;
    layer5_outputs(11887) <= b;
    layer5_outputs(11888) <= a xor b;
    layer5_outputs(11889) <= not (a xor b);
    layer5_outputs(11890) <= not a;
    layer5_outputs(11891) <= a or b;
    layer5_outputs(11892) <= a;
    layer5_outputs(11893) <= not a;
    layer5_outputs(11894) <= a;
    layer5_outputs(11895) <= a and b;
    layer5_outputs(11896) <= a or b;
    layer5_outputs(11897) <= not a or b;
    layer5_outputs(11898) <= not (a xor b);
    layer5_outputs(11899) <= not b;
    layer5_outputs(11900) <= not (a or b);
    layer5_outputs(11901) <= not b;
    layer5_outputs(11902) <= b;
    layer5_outputs(11903) <= a;
    layer5_outputs(11904) <= not a or b;
    layer5_outputs(11905) <= '0';
    layer5_outputs(11906) <= not a;
    layer5_outputs(11907) <= not b;
    layer5_outputs(11908) <= a;
    layer5_outputs(11909) <= a;
    layer5_outputs(11910) <= a and b;
    layer5_outputs(11911) <= not a;
    layer5_outputs(11912) <= a and not b;
    layer5_outputs(11913) <= not (a or b);
    layer5_outputs(11914) <= not (a xor b);
    layer5_outputs(11915) <= not a;
    layer5_outputs(11916) <= not a;
    layer5_outputs(11917) <= b;
    layer5_outputs(11918) <= b;
    layer5_outputs(11919) <= not a;
    layer5_outputs(11920) <= b;
    layer5_outputs(11921) <= a and not b;
    layer5_outputs(11922) <= not a or b;
    layer5_outputs(11923) <= a or b;
    layer5_outputs(11924) <= b;
    layer5_outputs(11925) <= not (a xor b);
    layer5_outputs(11926) <= not a;
    layer5_outputs(11927) <= not (a and b);
    layer5_outputs(11928) <= a;
    layer5_outputs(11929) <= not b or a;
    layer5_outputs(11930) <= b;
    layer5_outputs(11931) <= a;
    layer5_outputs(11932) <= a and b;
    layer5_outputs(11933) <= not (a and b);
    layer5_outputs(11934) <= b;
    layer5_outputs(11935) <= not a;
    layer5_outputs(11936) <= not a or b;
    layer5_outputs(11937) <= b;
    layer5_outputs(11938) <= b and not a;
    layer5_outputs(11939) <= not b;
    layer5_outputs(11940) <= a and not b;
    layer5_outputs(11941) <= a and not b;
    layer5_outputs(11942) <= a xor b;
    layer5_outputs(11943) <= not b or a;
    layer5_outputs(11944) <= not b or a;
    layer5_outputs(11945) <= not b;
    layer5_outputs(11946) <= a or b;
    layer5_outputs(11947) <= a;
    layer5_outputs(11948) <= a or b;
    layer5_outputs(11949) <= b;
    layer5_outputs(11950) <= not (a xor b);
    layer5_outputs(11951) <= b;
    layer5_outputs(11952) <= not (a or b);
    layer5_outputs(11953) <= a or b;
    layer5_outputs(11954) <= a;
    layer5_outputs(11955) <= a xor b;
    layer5_outputs(11956) <= a and not b;
    layer5_outputs(11957) <= not b;
    layer5_outputs(11958) <= not (a xor b);
    layer5_outputs(11959) <= not (a or b);
    layer5_outputs(11960) <= not a;
    layer5_outputs(11961) <= b;
    layer5_outputs(11962) <= a and not b;
    layer5_outputs(11963) <= a;
    layer5_outputs(11964) <= a and not b;
    layer5_outputs(11965) <= not a;
    layer5_outputs(11966) <= a;
    layer5_outputs(11967) <= a;
    layer5_outputs(11968) <= not a or b;
    layer5_outputs(11969) <= not a;
    layer5_outputs(11970) <= b;
    layer5_outputs(11971) <= a and b;
    layer5_outputs(11972) <= not (a and b);
    layer5_outputs(11973) <= a;
    layer5_outputs(11974) <= b;
    layer5_outputs(11975) <= a or b;
    layer5_outputs(11976) <= b;
    layer5_outputs(11977) <= not b;
    layer5_outputs(11978) <= a and b;
    layer5_outputs(11979) <= a and b;
    layer5_outputs(11980) <= a;
    layer5_outputs(11981) <= a or b;
    layer5_outputs(11982) <= a xor b;
    layer5_outputs(11983) <= not (a xor b);
    layer5_outputs(11984) <= not a;
    layer5_outputs(11985) <= not a or b;
    layer5_outputs(11986) <= b;
    layer5_outputs(11987) <= not b;
    layer5_outputs(11988) <= not b or a;
    layer5_outputs(11989) <= b and not a;
    layer5_outputs(11990) <= not (a xor b);
    layer5_outputs(11991) <= not b;
    layer5_outputs(11992) <= not b;
    layer5_outputs(11993) <= not b or a;
    layer5_outputs(11994) <= not (a or b);
    layer5_outputs(11995) <= b;
    layer5_outputs(11996) <= a and b;
    layer5_outputs(11997) <= a xor b;
    layer5_outputs(11998) <= not a;
    layer5_outputs(11999) <= not a;
    layer5_outputs(12000) <= not (a xor b);
    layer5_outputs(12001) <= b;
    layer5_outputs(12002) <= not a or b;
    layer5_outputs(12003) <= not b or a;
    layer5_outputs(12004) <= not a;
    layer5_outputs(12005) <= '1';
    layer5_outputs(12006) <= a;
    layer5_outputs(12007) <= not a or b;
    layer5_outputs(12008) <= not b;
    layer5_outputs(12009) <= not b;
    layer5_outputs(12010) <= a or b;
    layer5_outputs(12011) <= not a or b;
    layer5_outputs(12012) <= not b;
    layer5_outputs(12013) <= a and b;
    layer5_outputs(12014) <= not a;
    layer5_outputs(12015) <= a;
    layer5_outputs(12016) <= not b;
    layer5_outputs(12017) <= not a;
    layer5_outputs(12018) <= not (a xor b);
    layer5_outputs(12019) <= not a;
    layer5_outputs(12020) <= a xor b;
    layer5_outputs(12021) <= not a;
    layer5_outputs(12022) <= a;
    layer5_outputs(12023) <= '0';
    layer5_outputs(12024) <= not b;
    layer5_outputs(12025) <= a xor b;
    layer5_outputs(12026) <= not b;
    layer5_outputs(12027) <= a and not b;
    layer5_outputs(12028) <= a;
    layer5_outputs(12029) <= a or b;
    layer5_outputs(12030) <= a and b;
    layer5_outputs(12031) <= not a;
    layer5_outputs(12032) <= not a or b;
    layer5_outputs(12033) <= a xor b;
    layer5_outputs(12034) <= not (a xor b);
    layer5_outputs(12035) <= a xor b;
    layer5_outputs(12036) <= '0';
    layer5_outputs(12037) <= not a;
    layer5_outputs(12038) <= a xor b;
    layer5_outputs(12039) <= a and not b;
    layer5_outputs(12040) <= not a or b;
    layer5_outputs(12041) <= a and not b;
    layer5_outputs(12042) <= not (a xor b);
    layer5_outputs(12043) <= a;
    layer5_outputs(12044) <= not b;
    layer5_outputs(12045) <= a or b;
    layer5_outputs(12046) <= a or b;
    layer5_outputs(12047) <= a;
    layer5_outputs(12048) <= a and b;
    layer5_outputs(12049) <= not a or b;
    layer5_outputs(12050) <= a xor b;
    layer5_outputs(12051) <= a or b;
    layer5_outputs(12052) <= a;
    layer5_outputs(12053) <= a and b;
    layer5_outputs(12054) <= not a;
    layer5_outputs(12055) <= a xor b;
    layer5_outputs(12056) <= a xor b;
    layer5_outputs(12057) <= b;
    layer5_outputs(12058) <= not a or b;
    layer5_outputs(12059) <= a and not b;
    layer5_outputs(12060) <= not b;
    layer5_outputs(12061) <= b;
    layer5_outputs(12062) <= not b or a;
    layer5_outputs(12063) <= b;
    layer5_outputs(12064) <= not (a and b);
    layer5_outputs(12065) <= not (a and b);
    layer5_outputs(12066) <= b;
    layer5_outputs(12067) <= b;
    layer5_outputs(12068) <= not b;
    layer5_outputs(12069) <= not a;
    layer5_outputs(12070) <= a and not b;
    layer5_outputs(12071) <= a and not b;
    layer5_outputs(12072) <= not (a xor b);
    layer5_outputs(12073) <= b;
    layer5_outputs(12074) <= b;
    layer5_outputs(12075) <= b;
    layer5_outputs(12076) <= b;
    layer5_outputs(12077) <= not (a or b);
    layer5_outputs(12078) <= not a;
    layer5_outputs(12079) <= not a or b;
    layer5_outputs(12080) <= not a;
    layer5_outputs(12081) <= not b;
    layer5_outputs(12082) <= b and not a;
    layer5_outputs(12083) <= a and not b;
    layer5_outputs(12084) <= b;
    layer5_outputs(12085) <= a xor b;
    layer5_outputs(12086) <= a;
    layer5_outputs(12087) <= not (a xor b);
    layer5_outputs(12088) <= not (a or b);
    layer5_outputs(12089) <= not a;
    layer5_outputs(12090) <= not a;
    layer5_outputs(12091) <= a xor b;
    layer5_outputs(12092) <= '1';
    layer5_outputs(12093) <= b;
    layer5_outputs(12094) <= b;
    layer5_outputs(12095) <= not a;
    layer5_outputs(12096) <= not b;
    layer5_outputs(12097) <= not a;
    layer5_outputs(12098) <= not a;
    layer5_outputs(12099) <= not (a or b);
    layer5_outputs(12100) <= not b;
    layer5_outputs(12101) <= not b or a;
    layer5_outputs(12102) <= not (a xor b);
    layer5_outputs(12103) <= not b;
    layer5_outputs(12104) <= b and not a;
    layer5_outputs(12105) <= a;
    layer5_outputs(12106) <= not (a and b);
    layer5_outputs(12107) <= not a;
    layer5_outputs(12108) <= a xor b;
    layer5_outputs(12109) <= not b;
    layer5_outputs(12110) <= a and b;
    layer5_outputs(12111) <= b;
    layer5_outputs(12112) <= b;
    layer5_outputs(12113) <= a and b;
    layer5_outputs(12114) <= a;
    layer5_outputs(12115) <= a;
    layer5_outputs(12116) <= a;
    layer5_outputs(12117) <= not a;
    layer5_outputs(12118) <= not (a xor b);
    layer5_outputs(12119) <= not b;
    layer5_outputs(12120) <= not (a xor b);
    layer5_outputs(12121) <= not b;
    layer5_outputs(12122) <= b and not a;
    layer5_outputs(12123) <= not (a or b);
    layer5_outputs(12124) <= not (a and b);
    layer5_outputs(12125) <= not a or b;
    layer5_outputs(12126) <= not (a xor b);
    layer5_outputs(12127) <= a xor b;
    layer5_outputs(12128) <= b;
    layer5_outputs(12129) <= a or b;
    layer5_outputs(12130) <= a and b;
    layer5_outputs(12131) <= not a or b;
    layer5_outputs(12132) <= a;
    layer5_outputs(12133) <= a;
    layer5_outputs(12134) <= b;
    layer5_outputs(12135) <= not (a xor b);
    layer5_outputs(12136) <= a;
    layer5_outputs(12137) <= '0';
    layer5_outputs(12138) <= not a or b;
    layer5_outputs(12139) <= b;
    layer5_outputs(12140) <= a and b;
    layer5_outputs(12141) <= not b;
    layer5_outputs(12142) <= not b or a;
    layer5_outputs(12143) <= a and b;
    layer5_outputs(12144) <= a xor b;
    layer5_outputs(12145) <= b;
    layer5_outputs(12146) <= a;
    layer5_outputs(12147) <= not b;
    layer5_outputs(12148) <= not (a and b);
    layer5_outputs(12149) <= b;
    layer5_outputs(12150) <= '1';
    layer5_outputs(12151) <= a xor b;
    layer5_outputs(12152) <= b and not a;
    layer5_outputs(12153) <= b and not a;
    layer5_outputs(12154) <= a;
    layer5_outputs(12155) <= not a;
    layer5_outputs(12156) <= a and not b;
    layer5_outputs(12157) <= not (a xor b);
    layer5_outputs(12158) <= a or b;
    layer5_outputs(12159) <= b and not a;
    layer5_outputs(12160) <= a and b;
    layer5_outputs(12161) <= not a or b;
    layer5_outputs(12162) <= b;
    layer5_outputs(12163) <= not (a xor b);
    layer5_outputs(12164) <= a and b;
    layer5_outputs(12165) <= a;
    layer5_outputs(12166) <= not (a and b);
    layer5_outputs(12167) <= not b;
    layer5_outputs(12168) <= not a;
    layer5_outputs(12169) <= b;
    layer5_outputs(12170) <= not a;
    layer5_outputs(12171) <= not (a or b);
    layer5_outputs(12172) <= b;
    layer5_outputs(12173) <= a;
    layer5_outputs(12174) <= a xor b;
    layer5_outputs(12175) <= not a;
    layer5_outputs(12176) <= b;
    layer5_outputs(12177) <= not b;
    layer5_outputs(12178) <= not (a or b);
    layer5_outputs(12179) <= '1';
    layer5_outputs(12180) <= not b;
    layer5_outputs(12181) <= a;
    layer5_outputs(12182) <= a;
    layer5_outputs(12183) <= a;
    layer5_outputs(12184) <= not b;
    layer5_outputs(12185) <= a and not b;
    layer5_outputs(12186) <= a or b;
    layer5_outputs(12187) <= a xor b;
    layer5_outputs(12188) <= b;
    layer5_outputs(12189) <= not b;
    layer5_outputs(12190) <= not a;
    layer5_outputs(12191) <= not a;
    layer5_outputs(12192) <= a or b;
    layer5_outputs(12193) <= a and b;
    layer5_outputs(12194) <= a and not b;
    layer5_outputs(12195) <= b;
    layer5_outputs(12196) <= not (a xor b);
    layer5_outputs(12197) <= '1';
    layer5_outputs(12198) <= a or b;
    layer5_outputs(12199) <= not b;
    layer5_outputs(12200) <= not b;
    layer5_outputs(12201) <= a or b;
    layer5_outputs(12202) <= not b or a;
    layer5_outputs(12203) <= a xor b;
    layer5_outputs(12204) <= not a;
    layer5_outputs(12205) <= not (a xor b);
    layer5_outputs(12206) <= not (a xor b);
    layer5_outputs(12207) <= not a or b;
    layer5_outputs(12208) <= not b;
    layer5_outputs(12209) <= a xor b;
    layer5_outputs(12210) <= b;
    layer5_outputs(12211) <= not a;
    layer5_outputs(12212) <= a and b;
    layer5_outputs(12213) <= not b;
    layer5_outputs(12214) <= a xor b;
    layer5_outputs(12215) <= a;
    layer5_outputs(12216) <= b;
    layer5_outputs(12217) <= b;
    layer5_outputs(12218) <= a;
    layer5_outputs(12219) <= not (a xor b);
    layer5_outputs(12220) <= not (a and b);
    layer5_outputs(12221) <= not (a or b);
    layer5_outputs(12222) <= b;
    layer5_outputs(12223) <= a and b;
    layer5_outputs(12224) <= a;
    layer5_outputs(12225) <= a or b;
    layer5_outputs(12226) <= a xor b;
    layer5_outputs(12227) <= not a;
    layer5_outputs(12228) <= not (a or b);
    layer5_outputs(12229) <= a;
    layer5_outputs(12230) <= not a;
    layer5_outputs(12231) <= not a;
    layer5_outputs(12232) <= not (a or b);
    layer5_outputs(12233) <= not b;
    layer5_outputs(12234) <= not b;
    layer5_outputs(12235) <= not a or b;
    layer5_outputs(12236) <= b;
    layer5_outputs(12237) <= a or b;
    layer5_outputs(12238) <= '1';
    layer5_outputs(12239) <= b;
    layer5_outputs(12240) <= not b;
    layer5_outputs(12241) <= b and not a;
    layer5_outputs(12242) <= a xor b;
    layer5_outputs(12243) <= '0';
    layer5_outputs(12244) <= a and not b;
    layer5_outputs(12245) <= '1';
    layer5_outputs(12246) <= b;
    layer5_outputs(12247) <= not (a xor b);
    layer5_outputs(12248) <= not b;
    layer5_outputs(12249) <= not (a xor b);
    layer5_outputs(12250) <= b;
    layer5_outputs(12251) <= not a;
    layer5_outputs(12252) <= not a;
    layer5_outputs(12253) <= a and not b;
    layer5_outputs(12254) <= a;
    layer5_outputs(12255) <= not (a xor b);
    layer5_outputs(12256) <= not (a or b);
    layer5_outputs(12257) <= not b;
    layer5_outputs(12258) <= '0';
    layer5_outputs(12259) <= not (a and b);
    layer5_outputs(12260) <= not b;
    layer5_outputs(12261) <= not a;
    layer5_outputs(12262) <= a;
    layer5_outputs(12263) <= a;
    layer5_outputs(12264) <= not a or b;
    layer5_outputs(12265) <= b and not a;
    layer5_outputs(12266) <= '0';
    layer5_outputs(12267) <= not b or a;
    layer5_outputs(12268) <= a and not b;
    layer5_outputs(12269) <= a xor b;
    layer5_outputs(12270) <= not (a and b);
    layer5_outputs(12271) <= a or b;
    layer5_outputs(12272) <= a or b;
    layer5_outputs(12273) <= a and not b;
    layer5_outputs(12274) <= a;
    layer5_outputs(12275) <= b;
    layer5_outputs(12276) <= a xor b;
    layer5_outputs(12277) <= a or b;
    layer5_outputs(12278) <= '1';
    layer5_outputs(12279) <= a and not b;
    layer5_outputs(12280) <= not (a xor b);
    layer5_outputs(12281) <= not (a or b);
    layer5_outputs(12282) <= a and b;
    layer5_outputs(12283) <= not (a and b);
    layer5_outputs(12284) <= a;
    layer5_outputs(12285) <= b and not a;
    layer5_outputs(12286) <= not b or a;
    layer5_outputs(12287) <= not b;
    layer5_outputs(12288) <= a and not b;
    layer5_outputs(12289) <= a and not b;
    layer5_outputs(12290) <= '1';
    layer5_outputs(12291) <= not a;
    layer5_outputs(12292) <= b;
    layer5_outputs(12293) <= not (a xor b);
    layer5_outputs(12294) <= not b or a;
    layer5_outputs(12295) <= not a;
    layer5_outputs(12296) <= a and b;
    layer5_outputs(12297) <= a and b;
    layer5_outputs(12298) <= not b;
    layer5_outputs(12299) <= not a or b;
    layer5_outputs(12300) <= not (a and b);
    layer5_outputs(12301) <= a and b;
    layer5_outputs(12302) <= not (a xor b);
    layer5_outputs(12303) <= b and not a;
    layer5_outputs(12304) <= b and not a;
    layer5_outputs(12305) <= not a or b;
    layer5_outputs(12306) <= not b;
    layer5_outputs(12307) <= a;
    layer5_outputs(12308) <= a xor b;
    layer5_outputs(12309) <= b;
    layer5_outputs(12310) <= a and not b;
    layer5_outputs(12311) <= a or b;
    layer5_outputs(12312) <= a;
    layer5_outputs(12313) <= b;
    layer5_outputs(12314) <= a and b;
    layer5_outputs(12315) <= a;
    layer5_outputs(12316) <= not a;
    layer5_outputs(12317) <= b;
    layer5_outputs(12318) <= not b or a;
    layer5_outputs(12319) <= a and not b;
    layer5_outputs(12320) <= not a or b;
    layer5_outputs(12321) <= not (a or b);
    layer5_outputs(12322) <= not (a and b);
    layer5_outputs(12323) <= not b;
    layer5_outputs(12324) <= not a or b;
    layer5_outputs(12325) <= b and not a;
    layer5_outputs(12326) <= a xor b;
    layer5_outputs(12327) <= not (a and b);
    layer5_outputs(12328) <= not b or a;
    layer5_outputs(12329) <= '0';
    layer5_outputs(12330) <= not (a and b);
    layer5_outputs(12331) <= a and not b;
    layer5_outputs(12332) <= not b;
    layer5_outputs(12333) <= not b or a;
    layer5_outputs(12334) <= '0';
    layer5_outputs(12335) <= a xor b;
    layer5_outputs(12336) <= a and b;
    layer5_outputs(12337) <= not a;
    layer5_outputs(12338) <= not a;
    layer5_outputs(12339) <= a or b;
    layer5_outputs(12340) <= a;
    layer5_outputs(12341) <= not a;
    layer5_outputs(12342) <= a or b;
    layer5_outputs(12343) <= not b or a;
    layer5_outputs(12344) <= '1';
    layer5_outputs(12345) <= not b;
    layer5_outputs(12346) <= a or b;
    layer5_outputs(12347) <= a xor b;
    layer5_outputs(12348) <= b;
    layer5_outputs(12349) <= a and b;
    layer5_outputs(12350) <= a and b;
    layer5_outputs(12351) <= b;
    layer5_outputs(12352) <= a;
    layer5_outputs(12353) <= not (a xor b);
    layer5_outputs(12354) <= not (a or b);
    layer5_outputs(12355) <= not a;
    layer5_outputs(12356) <= a and b;
    layer5_outputs(12357) <= a xor b;
    layer5_outputs(12358) <= a;
    layer5_outputs(12359) <= a xor b;
    layer5_outputs(12360) <= a and b;
    layer5_outputs(12361) <= a and b;
    layer5_outputs(12362) <= a;
    layer5_outputs(12363) <= a;
    layer5_outputs(12364) <= a xor b;
    layer5_outputs(12365) <= a xor b;
    layer5_outputs(12366) <= a and b;
    layer5_outputs(12367) <= not a;
    layer5_outputs(12368) <= b and not a;
    layer5_outputs(12369) <= not (a or b);
    layer5_outputs(12370) <= not b or a;
    layer5_outputs(12371) <= not b or a;
    layer5_outputs(12372) <= not (a or b);
    layer5_outputs(12373) <= not a;
    layer5_outputs(12374) <= not a;
    layer5_outputs(12375) <= a and b;
    layer5_outputs(12376) <= '1';
    layer5_outputs(12377) <= not b or a;
    layer5_outputs(12378) <= b;
    layer5_outputs(12379) <= not a;
    layer5_outputs(12380) <= not (a or b);
    layer5_outputs(12381) <= not a;
    layer5_outputs(12382) <= a and b;
    layer5_outputs(12383) <= not a or b;
    layer5_outputs(12384) <= not (a or b);
    layer5_outputs(12385) <= not a or b;
    layer5_outputs(12386) <= a xor b;
    layer5_outputs(12387) <= a;
    layer5_outputs(12388) <= not (a or b);
    layer5_outputs(12389) <= b;
    layer5_outputs(12390) <= a and b;
    layer5_outputs(12391) <= not b;
    layer5_outputs(12392) <= a;
    layer5_outputs(12393) <= not (a or b);
    layer5_outputs(12394) <= not b;
    layer5_outputs(12395) <= a and b;
    layer5_outputs(12396) <= '1';
    layer5_outputs(12397) <= a and not b;
    layer5_outputs(12398) <= b and not a;
    layer5_outputs(12399) <= b and not a;
    layer5_outputs(12400) <= b;
    layer5_outputs(12401) <= not a;
    layer5_outputs(12402) <= b;
    layer5_outputs(12403) <= a and not b;
    layer5_outputs(12404) <= not a;
    layer5_outputs(12405) <= b and not a;
    layer5_outputs(12406) <= not (a xor b);
    layer5_outputs(12407) <= not a;
    layer5_outputs(12408) <= b;
    layer5_outputs(12409) <= not a;
    layer5_outputs(12410) <= not b;
    layer5_outputs(12411) <= b;
    layer5_outputs(12412) <= not a;
    layer5_outputs(12413) <= b;
    layer5_outputs(12414) <= not a or b;
    layer5_outputs(12415) <= not (a xor b);
    layer5_outputs(12416) <= not (a xor b);
    layer5_outputs(12417) <= a;
    layer5_outputs(12418) <= not a;
    layer5_outputs(12419) <= b and not a;
    layer5_outputs(12420) <= not a or b;
    layer5_outputs(12421) <= a;
    layer5_outputs(12422) <= not (a xor b);
    layer5_outputs(12423) <= a and b;
    layer5_outputs(12424) <= not b;
    layer5_outputs(12425) <= a and not b;
    layer5_outputs(12426) <= not a or b;
    layer5_outputs(12427) <= not a;
    layer5_outputs(12428) <= a xor b;
    layer5_outputs(12429) <= not (a xor b);
    layer5_outputs(12430) <= a xor b;
    layer5_outputs(12431) <= not (a or b);
    layer5_outputs(12432) <= b and not a;
    layer5_outputs(12433) <= a;
    layer5_outputs(12434) <= a and b;
    layer5_outputs(12435) <= '0';
    layer5_outputs(12436) <= a and b;
    layer5_outputs(12437) <= b;
    layer5_outputs(12438) <= not b;
    layer5_outputs(12439) <= b;
    layer5_outputs(12440) <= not (a or b);
    layer5_outputs(12441) <= a xor b;
    layer5_outputs(12442) <= not a;
    layer5_outputs(12443) <= not a or b;
    layer5_outputs(12444) <= not b or a;
    layer5_outputs(12445) <= b;
    layer5_outputs(12446) <= not b;
    layer5_outputs(12447) <= b;
    layer5_outputs(12448) <= not (a xor b);
    layer5_outputs(12449) <= not a;
    layer5_outputs(12450) <= not b;
    layer5_outputs(12451) <= a;
    layer5_outputs(12452) <= a and not b;
    layer5_outputs(12453) <= not (a xor b);
    layer5_outputs(12454) <= b and not a;
    layer5_outputs(12455) <= a;
    layer5_outputs(12456) <= not a;
    layer5_outputs(12457) <= a and not b;
    layer5_outputs(12458) <= b;
    layer5_outputs(12459) <= a or b;
    layer5_outputs(12460) <= a or b;
    layer5_outputs(12461) <= a;
    layer5_outputs(12462) <= not a or b;
    layer5_outputs(12463) <= not b;
    layer5_outputs(12464) <= not b;
    layer5_outputs(12465) <= not a or b;
    layer5_outputs(12466) <= not (a xor b);
    layer5_outputs(12467) <= a or b;
    layer5_outputs(12468) <= not a;
    layer5_outputs(12469) <= not b;
    layer5_outputs(12470) <= a;
    layer5_outputs(12471) <= not b;
    layer5_outputs(12472) <= not b;
    layer5_outputs(12473) <= not b;
    layer5_outputs(12474) <= a;
    layer5_outputs(12475) <= not b;
    layer5_outputs(12476) <= not a or b;
    layer5_outputs(12477) <= b;
    layer5_outputs(12478) <= not b;
    layer5_outputs(12479) <= not (a xor b);
    layer5_outputs(12480) <= a;
    layer5_outputs(12481) <= b and not a;
    layer5_outputs(12482) <= a or b;
    layer5_outputs(12483) <= not (a and b);
    layer5_outputs(12484) <= a and b;
    layer5_outputs(12485) <= not b;
    layer5_outputs(12486) <= not b;
    layer5_outputs(12487) <= not b;
    layer5_outputs(12488) <= not b;
    layer5_outputs(12489) <= a xor b;
    layer5_outputs(12490) <= not (a xor b);
    layer5_outputs(12491) <= not a;
    layer5_outputs(12492) <= a xor b;
    layer5_outputs(12493) <= a;
    layer5_outputs(12494) <= not a;
    layer5_outputs(12495) <= a and not b;
    layer5_outputs(12496) <= a and b;
    layer5_outputs(12497) <= a xor b;
    layer5_outputs(12498) <= not b;
    layer5_outputs(12499) <= not a;
    layer5_outputs(12500) <= not b;
    layer5_outputs(12501) <= not a;
    layer5_outputs(12502) <= a;
    layer5_outputs(12503) <= not b;
    layer5_outputs(12504) <= a and not b;
    layer5_outputs(12505) <= not (a xor b);
    layer5_outputs(12506) <= not a or b;
    layer5_outputs(12507) <= not a;
    layer5_outputs(12508) <= a xor b;
    layer5_outputs(12509) <= a xor b;
    layer5_outputs(12510) <= not a;
    layer5_outputs(12511) <= b;
    layer5_outputs(12512) <= not b;
    layer5_outputs(12513) <= not (a xor b);
    layer5_outputs(12514) <= not b or a;
    layer5_outputs(12515) <= not b;
    layer5_outputs(12516) <= a and not b;
    layer5_outputs(12517) <= not b;
    layer5_outputs(12518) <= not a;
    layer5_outputs(12519) <= a;
    layer5_outputs(12520) <= not (a or b);
    layer5_outputs(12521) <= a;
    layer5_outputs(12522) <= not b;
    layer5_outputs(12523) <= not b or a;
    layer5_outputs(12524) <= a;
    layer5_outputs(12525) <= not (a or b);
    layer5_outputs(12526) <= not a;
    layer5_outputs(12527) <= b;
    layer5_outputs(12528) <= not b;
    layer5_outputs(12529) <= not (a and b);
    layer5_outputs(12530) <= b;
    layer5_outputs(12531) <= not b;
    layer5_outputs(12532) <= not b or a;
    layer5_outputs(12533) <= not (a or b);
    layer5_outputs(12534) <= not a;
    layer5_outputs(12535) <= a or b;
    layer5_outputs(12536) <= not b;
    layer5_outputs(12537) <= not b;
    layer5_outputs(12538) <= a xor b;
    layer5_outputs(12539) <= not (a xor b);
    layer5_outputs(12540) <= not (a xor b);
    layer5_outputs(12541) <= not a;
    layer5_outputs(12542) <= not b or a;
    layer5_outputs(12543) <= a and b;
    layer5_outputs(12544) <= '1';
    layer5_outputs(12545) <= not a;
    layer5_outputs(12546) <= not b;
    layer5_outputs(12547) <= b;
    layer5_outputs(12548) <= not (a or b);
    layer5_outputs(12549) <= not (a xor b);
    layer5_outputs(12550) <= a xor b;
    layer5_outputs(12551) <= a;
    layer5_outputs(12552) <= b;
    layer5_outputs(12553) <= not a;
    layer5_outputs(12554) <= a;
    layer5_outputs(12555) <= not (a or b);
    layer5_outputs(12556) <= not b;
    layer5_outputs(12557) <= a;
    layer5_outputs(12558) <= b;
    layer5_outputs(12559) <= not a;
    layer5_outputs(12560) <= b;
    layer5_outputs(12561) <= b;
    layer5_outputs(12562) <= not a;
    layer5_outputs(12563) <= not a;
    layer5_outputs(12564) <= not b;
    layer5_outputs(12565) <= b;
    layer5_outputs(12566) <= not (a or b);
    layer5_outputs(12567) <= a and b;
    layer5_outputs(12568) <= a and not b;
    layer5_outputs(12569) <= not (a or b);
    layer5_outputs(12570) <= not (a or b);
    layer5_outputs(12571) <= not (a or b);
    layer5_outputs(12572) <= not b;
    layer5_outputs(12573) <= not (a and b);
    layer5_outputs(12574) <= b;
    layer5_outputs(12575) <= not b;
    layer5_outputs(12576) <= a xor b;
    layer5_outputs(12577) <= not b or a;
    layer5_outputs(12578) <= '1';
    layer5_outputs(12579) <= not b;
    layer5_outputs(12580) <= b;
    layer5_outputs(12581) <= a;
    layer5_outputs(12582) <= a or b;
    layer5_outputs(12583) <= not b;
    layer5_outputs(12584) <= a or b;
    layer5_outputs(12585) <= a or b;
    layer5_outputs(12586) <= a xor b;
    layer5_outputs(12587) <= not b;
    layer5_outputs(12588) <= a xor b;
    layer5_outputs(12589) <= a;
    layer5_outputs(12590) <= a;
    layer5_outputs(12591) <= a;
    layer5_outputs(12592) <= not (a or b);
    layer5_outputs(12593) <= not b or a;
    layer5_outputs(12594) <= b;
    layer5_outputs(12595) <= a;
    layer5_outputs(12596) <= a;
    layer5_outputs(12597) <= not b;
    layer5_outputs(12598) <= not b;
    layer5_outputs(12599) <= not (a or b);
    layer5_outputs(12600) <= b and not a;
    layer5_outputs(12601) <= not (a and b);
    layer5_outputs(12602) <= not b;
    layer5_outputs(12603) <= not a;
    layer5_outputs(12604) <= b;
    layer5_outputs(12605) <= not a;
    layer5_outputs(12606) <= a xor b;
    layer5_outputs(12607) <= not (a and b);
    layer5_outputs(12608) <= a xor b;
    layer5_outputs(12609) <= not (a and b);
    layer5_outputs(12610) <= not a;
    layer5_outputs(12611) <= b;
    layer5_outputs(12612) <= a;
    layer5_outputs(12613) <= not a;
    layer5_outputs(12614) <= not b;
    layer5_outputs(12615) <= not b or a;
    layer5_outputs(12616) <= not a or b;
    layer5_outputs(12617) <= a and not b;
    layer5_outputs(12618) <= not a;
    layer5_outputs(12619) <= '0';
    layer5_outputs(12620) <= a;
    layer5_outputs(12621) <= not a or b;
    layer5_outputs(12622) <= b;
    layer5_outputs(12623) <= not a;
    layer5_outputs(12624) <= a and not b;
    layer5_outputs(12625) <= a xor b;
    layer5_outputs(12626) <= a and b;
    layer5_outputs(12627) <= not a or b;
    layer5_outputs(12628) <= a and b;
    layer5_outputs(12629) <= a and b;
    layer5_outputs(12630) <= a xor b;
    layer5_outputs(12631) <= not b or a;
    layer5_outputs(12632) <= not a or b;
    layer5_outputs(12633) <= not b;
    layer5_outputs(12634) <= a xor b;
    layer5_outputs(12635) <= a and b;
    layer5_outputs(12636) <= not a;
    layer5_outputs(12637) <= b and not a;
    layer5_outputs(12638) <= '0';
    layer5_outputs(12639) <= b;
    layer5_outputs(12640) <= not (a xor b);
    layer5_outputs(12641) <= a xor b;
    layer5_outputs(12642) <= b;
    layer5_outputs(12643) <= b;
    layer5_outputs(12644) <= not b;
    layer5_outputs(12645) <= a;
    layer5_outputs(12646) <= a;
    layer5_outputs(12647) <= a xor b;
    layer5_outputs(12648) <= not a or b;
    layer5_outputs(12649) <= b;
    layer5_outputs(12650) <= not a;
    layer5_outputs(12651) <= b;
    layer5_outputs(12652) <= not (a or b);
    layer5_outputs(12653) <= not b or a;
    layer5_outputs(12654) <= not b or a;
    layer5_outputs(12655) <= not (a or b);
    layer5_outputs(12656) <= a;
    layer5_outputs(12657) <= not b;
    layer5_outputs(12658) <= not a or b;
    layer5_outputs(12659) <= a;
    layer5_outputs(12660) <= not (a or b);
    layer5_outputs(12661) <= not b;
    layer5_outputs(12662) <= a xor b;
    layer5_outputs(12663) <= not a;
    layer5_outputs(12664) <= not (a and b);
    layer5_outputs(12665) <= not a;
    layer5_outputs(12666) <= b;
    layer5_outputs(12667) <= a and not b;
    layer5_outputs(12668) <= not b or a;
    layer5_outputs(12669) <= not (a xor b);
    layer5_outputs(12670) <= a and not b;
    layer5_outputs(12671) <= a;
    layer5_outputs(12672) <= not b;
    layer5_outputs(12673) <= not b;
    layer5_outputs(12674) <= not b;
    layer5_outputs(12675) <= not a or b;
    layer5_outputs(12676) <= not a;
    layer5_outputs(12677) <= not b;
    layer5_outputs(12678) <= not a;
    layer5_outputs(12679) <= not b;
    layer5_outputs(12680) <= not (a xor b);
    layer5_outputs(12681) <= b;
    layer5_outputs(12682) <= b;
    layer5_outputs(12683) <= not a or b;
    layer5_outputs(12684) <= not a;
    layer5_outputs(12685) <= a;
    layer5_outputs(12686) <= not b;
    layer5_outputs(12687) <= a;
    layer5_outputs(12688) <= not a;
    layer5_outputs(12689) <= '0';
    layer5_outputs(12690) <= not b;
    layer5_outputs(12691) <= b;
    layer5_outputs(12692) <= b;
    layer5_outputs(12693) <= not (a xor b);
    layer5_outputs(12694) <= not (a xor b);
    layer5_outputs(12695) <= b;
    layer5_outputs(12696) <= b;
    layer5_outputs(12697) <= a xor b;
    layer5_outputs(12698) <= not b or a;
    layer5_outputs(12699) <= a;
    layer5_outputs(12700) <= b;
    layer5_outputs(12701) <= a;
    layer5_outputs(12702) <= a and b;
    layer5_outputs(12703) <= not a;
    layer5_outputs(12704) <= a or b;
    layer5_outputs(12705) <= b and not a;
    layer5_outputs(12706) <= b and not a;
    layer5_outputs(12707) <= not a or b;
    layer5_outputs(12708) <= b and not a;
    layer5_outputs(12709) <= b;
    layer5_outputs(12710) <= not b;
    layer5_outputs(12711) <= a;
    layer5_outputs(12712) <= a and not b;
    layer5_outputs(12713) <= a xor b;
    layer5_outputs(12714) <= a;
    layer5_outputs(12715) <= b and not a;
    layer5_outputs(12716) <= a xor b;
    layer5_outputs(12717) <= not (a xor b);
    layer5_outputs(12718) <= not b;
    layer5_outputs(12719) <= b;
    layer5_outputs(12720) <= b and not a;
    layer5_outputs(12721) <= not (a xor b);
    layer5_outputs(12722) <= a and b;
    layer5_outputs(12723) <= not (a and b);
    layer5_outputs(12724) <= not a;
    layer5_outputs(12725) <= a;
    layer5_outputs(12726) <= not (a and b);
    layer5_outputs(12727) <= b;
    layer5_outputs(12728) <= not a;
    layer5_outputs(12729) <= not a;
    layer5_outputs(12730) <= not a;
    layer5_outputs(12731) <= b;
    layer5_outputs(12732) <= not a;
    layer5_outputs(12733) <= a and b;
    layer5_outputs(12734) <= not b or a;
    layer5_outputs(12735) <= not b;
    layer5_outputs(12736) <= b and not a;
    layer5_outputs(12737) <= not a;
    layer5_outputs(12738) <= b and not a;
    layer5_outputs(12739) <= a and not b;
    layer5_outputs(12740) <= not a;
    layer5_outputs(12741) <= b;
    layer5_outputs(12742) <= a xor b;
    layer5_outputs(12743) <= not (a xor b);
    layer5_outputs(12744) <= a;
    layer5_outputs(12745) <= not a or b;
    layer5_outputs(12746) <= not (a xor b);
    layer5_outputs(12747) <= b;
    layer5_outputs(12748) <= a and b;
    layer5_outputs(12749) <= not b;
    layer5_outputs(12750) <= not a;
    layer5_outputs(12751) <= a and not b;
    layer5_outputs(12752) <= a xor b;
    layer5_outputs(12753) <= a xor b;
    layer5_outputs(12754) <= not b;
    layer5_outputs(12755) <= not (a and b);
    layer5_outputs(12756) <= a xor b;
    layer5_outputs(12757) <= not (a xor b);
    layer5_outputs(12758) <= not (a and b);
    layer5_outputs(12759) <= not a or b;
    layer5_outputs(12760) <= b;
    layer5_outputs(12761) <= a or b;
    layer5_outputs(12762) <= not a or b;
    layer5_outputs(12763) <= not a;
    layer5_outputs(12764) <= not b;
    layer5_outputs(12765) <= not b or a;
    layer5_outputs(12766) <= a and not b;
    layer5_outputs(12767) <= a xor b;
    layer5_outputs(12768) <= not (a xor b);
    layer5_outputs(12769) <= a;
    layer5_outputs(12770) <= not a or b;
    layer5_outputs(12771) <= a xor b;
    layer5_outputs(12772) <= not a or b;
    layer5_outputs(12773) <= not (a or b);
    layer5_outputs(12774) <= not b or a;
    layer5_outputs(12775) <= not b;
    layer5_outputs(12776) <= not (a xor b);
    layer5_outputs(12777) <= b;
    layer5_outputs(12778) <= a and not b;
    layer5_outputs(12779) <= not a or b;
    layer5_outputs(12780) <= not a or b;
    layer5_outputs(12781) <= a and b;
    layer5_outputs(12782) <= not (a or b);
    layer5_outputs(12783) <= '1';
    layer5_outputs(12784) <= not a;
    layer5_outputs(12785) <= not a;
    layer5_outputs(12786) <= not b;
    layer5_outputs(12787) <= not b;
    layer5_outputs(12788) <= b;
    layer5_outputs(12789) <= not a;
    layer5_outputs(12790) <= not (a and b);
    layer5_outputs(12791) <= not a or b;
    layer5_outputs(12792) <= a and b;
    layer5_outputs(12793) <= not (a xor b);
    layer5_outputs(12794) <= not b or a;
    layer5_outputs(12795) <= '1';
    layer5_outputs(12796) <= a and b;
    layer5_outputs(12797) <= not b;
    layer5_outputs(12798) <= not b or a;
    layer5_outputs(12799) <= a and not b;
    layer6_outputs(0) <= a and not b;
    layer6_outputs(1) <= not (a xor b);
    layer6_outputs(2) <= not b;
    layer6_outputs(3) <= not (a xor b);
    layer6_outputs(4) <= a and b;
    layer6_outputs(5) <= not (a xor b);
    layer6_outputs(6) <= a and b;
    layer6_outputs(7) <= not a;
    layer6_outputs(8) <= not (a xor b);
    layer6_outputs(9) <= not a;
    layer6_outputs(10) <= b;
    layer6_outputs(11) <= a and b;
    layer6_outputs(12) <= not a;
    layer6_outputs(13) <= not a or b;
    layer6_outputs(14) <= not (a xor b);
    layer6_outputs(15) <= not b;
    layer6_outputs(16) <= not a;
    layer6_outputs(17) <= a or b;
    layer6_outputs(18) <= not a or b;
    layer6_outputs(19) <= a;
    layer6_outputs(20) <= b;
    layer6_outputs(21) <= not a;
    layer6_outputs(22) <= not a;
    layer6_outputs(23) <= not b or a;
    layer6_outputs(24) <= a xor b;
    layer6_outputs(25) <= b and not a;
    layer6_outputs(26) <= b;
    layer6_outputs(27) <= not (a xor b);
    layer6_outputs(28) <= not b;
    layer6_outputs(29) <= a;
    layer6_outputs(30) <= b;
    layer6_outputs(31) <= a xor b;
    layer6_outputs(32) <= a xor b;
    layer6_outputs(33) <= a and b;
    layer6_outputs(34) <= not b;
    layer6_outputs(35) <= not a;
    layer6_outputs(36) <= not a;
    layer6_outputs(37) <= a xor b;
    layer6_outputs(38) <= b and not a;
    layer6_outputs(39) <= not (a xor b);
    layer6_outputs(40) <= a xor b;
    layer6_outputs(41) <= not b;
    layer6_outputs(42) <= a;
    layer6_outputs(43) <= not b or a;
    layer6_outputs(44) <= a and not b;
    layer6_outputs(45) <= a;
    layer6_outputs(46) <= not (a or b);
    layer6_outputs(47) <= a;
    layer6_outputs(48) <= not (a xor b);
    layer6_outputs(49) <= b;
    layer6_outputs(50) <= '0';
    layer6_outputs(51) <= not b;
    layer6_outputs(52) <= a or b;
    layer6_outputs(53) <= b;
    layer6_outputs(54) <= not a;
    layer6_outputs(55) <= not b;
    layer6_outputs(56) <= not (a or b);
    layer6_outputs(57) <= a and b;
    layer6_outputs(58) <= not a or b;
    layer6_outputs(59) <= b and not a;
    layer6_outputs(60) <= b and not a;
    layer6_outputs(61) <= not (a xor b);
    layer6_outputs(62) <= not (a xor b);
    layer6_outputs(63) <= a or b;
    layer6_outputs(64) <= a;
    layer6_outputs(65) <= not b;
    layer6_outputs(66) <= not (a and b);
    layer6_outputs(67) <= a xor b;
    layer6_outputs(68) <= not (a xor b);
    layer6_outputs(69) <= not (a xor b);
    layer6_outputs(70) <= a and not b;
    layer6_outputs(71) <= not b;
    layer6_outputs(72) <= b;
    layer6_outputs(73) <= a xor b;
    layer6_outputs(74) <= not a or b;
    layer6_outputs(75) <= not (a and b);
    layer6_outputs(76) <= not a;
    layer6_outputs(77) <= a or b;
    layer6_outputs(78) <= a;
    layer6_outputs(79) <= b;
    layer6_outputs(80) <= b;
    layer6_outputs(81) <= not a;
    layer6_outputs(82) <= not a;
    layer6_outputs(83) <= not a or b;
    layer6_outputs(84) <= a;
    layer6_outputs(85) <= a xor b;
    layer6_outputs(86) <= not b;
    layer6_outputs(87) <= not (a and b);
    layer6_outputs(88) <= not b;
    layer6_outputs(89) <= a and b;
    layer6_outputs(90) <= not (a and b);
    layer6_outputs(91) <= not a;
    layer6_outputs(92) <= not a or b;
    layer6_outputs(93) <= not b or a;
    layer6_outputs(94) <= not (a xor b);
    layer6_outputs(95) <= not a;
    layer6_outputs(96) <= a or b;
    layer6_outputs(97) <= b;
    layer6_outputs(98) <= a;
    layer6_outputs(99) <= not b;
    layer6_outputs(100) <= not a;
    layer6_outputs(101) <= a xor b;
    layer6_outputs(102) <= b;
    layer6_outputs(103) <= a xor b;
    layer6_outputs(104) <= b;
    layer6_outputs(105) <= b and not a;
    layer6_outputs(106) <= a and b;
    layer6_outputs(107) <= a;
    layer6_outputs(108) <= b and not a;
    layer6_outputs(109) <= '0';
    layer6_outputs(110) <= b and not a;
    layer6_outputs(111) <= not b;
    layer6_outputs(112) <= not (a xor b);
    layer6_outputs(113) <= a and b;
    layer6_outputs(114) <= not a or b;
    layer6_outputs(115) <= a xor b;
    layer6_outputs(116) <= b;
    layer6_outputs(117) <= not b or a;
    layer6_outputs(118) <= '0';
    layer6_outputs(119) <= b and not a;
    layer6_outputs(120) <= not (a xor b);
    layer6_outputs(121) <= a or b;
    layer6_outputs(122) <= b;
    layer6_outputs(123) <= a xor b;
    layer6_outputs(124) <= a xor b;
    layer6_outputs(125) <= not (a xor b);
    layer6_outputs(126) <= b and not a;
    layer6_outputs(127) <= not b;
    layer6_outputs(128) <= not a;
    layer6_outputs(129) <= a or b;
    layer6_outputs(130) <= not (a xor b);
    layer6_outputs(131) <= not b;
    layer6_outputs(132) <= a xor b;
    layer6_outputs(133) <= not a or b;
    layer6_outputs(134) <= a;
    layer6_outputs(135) <= a and not b;
    layer6_outputs(136) <= a or b;
    layer6_outputs(137) <= not b;
    layer6_outputs(138) <= not b;
    layer6_outputs(139) <= a and not b;
    layer6_outputs(140) <= b;
    layer6_outputs(141) <= not b;
    layer6_outputs(142) <= not (a xor b);
    layer6_outputs(143) <= not (a xor b);
    layer6_outputs(144) <= not b;
    layer6_outputs(145) <= not a;
    layer6_outputs(146) <= not b;
    layer6_outputs(147) <= b;
    layer6_outputs(148) <= a xor b;
    layer6_outputs(149) <= not a;
    layer6_outputs(150) <= not b;
    layer6_outputs(151) <= a or b;
    layer6_outputs(152) <= a xor b;
    layer6_outputs(153) <= not a;
    layer6_outputs(154) <= not a;
    layer6_outputs(155) <= b and not a;
    layer6_outputs(156) <= not (a and b);
    layer6_outputs(157) <= not (a xor b);
    layer6_outputs(158) <= b;
    layer6_outputs(159) <= not a or b;
    layer6_outputs(160) <= not a or b;
    layer6_outputs(161) <= not (a xor b);
    layer6_outputs(162) <= b;
    layer6_outputs(163) <= not (a or b);
    layer6_outputs(164) <= b;
    layer6_outputs(165) <= not a;
    layer6_outputs(166) <= not b;
    layer6_outputs(167) <= a xor b;
    layer6_outputs(168) <= not b;
    layer6_outputs(169) <= not (a xor b);
    layer6_outputs(170) <= a and b;
    layer6_outputs(171) <= b;
    layer6_outputs(172) <= not (a xor b);
    layer6_outputs(173) <= a xor b;
    layer6_outputs(174) <= a xor b;
    layer6_outputs(175) <= not b or a;
    layer6_outputs(176) <= not a;
    layer6_outputs(177) <= not (a and b);
    layer6_outputs(178) <= a xor b;
    layer6_outputs(179) <= a;
    layer6_outputs(180) <= a and not b;
    layer6_outputs(181) <= a and b;
    layer6_outputs(182) <= not b;
    layer6_outputs(183) <= not (a xor b);
    layer6_outputs(184) <= a and not b;
    layer6_outputs(185) <= b;
    layer6_outputs(186) <= b and not a;
    layer6_outputs(187) <= a xor b;
    layer6_outputs(188) <= b;
    layer6_outputs(189) <= not (a xor b);
    layer6_outputs(190) <= not (a or b);
    layer6_outputs(191) <= not a or b;
    layer6_outputs(192) <= not (a xor b);
    layer6_outputs(193) <= not (a or b);
    layer6_outputs(194) <= a;
    layer6_outputs(195) <= not (a and b);
    layer6_outputs(196) <= not a;
    layer6_outputs(197) <= a and b;
    layer6_outputs(198) <= a xor b;
    layer6_outputs(199) <= a;
    layer6_outputs(200) <= not a;
    layer6_outputs(201) <= a and not b;
    layer6_outputs(202) <= a or b;
    layer6_outputs(203) <= not a or b;
    layer6_outputs(204) <= not (a and b);
    layer6_outputs(205) <= not (a xor b);
    layer6_outputs(206) <= b;
    layer6_outputs(207) <= b and not a;
    layer6_outputs(208) <= b;
    layer6_outputs(209) <= not a;
    layer6_outputs(210) <= b;
    layer6_outputs(211) <= a;
    layer6_outputs(212) <= not a or b;
    layer6_outputs(213) <= b and not a;
    layer6_outputs(214) <= a and b;
    layer6_outputs(215) <= not a or b;
    layer6_outputs(216) <= a;
    layer6_outputs(217) <= a;
    layer6_outputs(218) <= a;
    layer6_outputs(219) <= a or b;
    layer6_outputs(220) <= a and not b;
    layer6_outputs(221) <= not a;
    layer6_outputs(222) <= b;
    layer6_outputs(223) <= a xor b;
    layer6_outputs(224) <= not (a and b);
    layer6_outputs(225) <= not b or a;
    layer6_outputs(226) <= a;
    layer6_outputs(227) <= not a;
    layer6_outputs(228) <= not a or b;
    layer6_outputs(229) <= a and b;
    layer6_outputs(230) <= not b;
    layer6_outputs(231) <= a;
    layer6_outputs(232) <= b;
    layer6_outputs(233) <= not a;
    layer6_outputs(234) <= '0';
    layer6_outputs(235) <= b and not a;
    layer6_outputs(236) <= a and not b;
    layer6_outputs(237) <= b;
    layer6_outputs(238) <= b and not a;
    layer6_outputs(239) <= b;
    layer6_outputs(240) <= not (a and b);
    layer6_outputs(241) <= not a;
    layer6_outputs(242) <= a or b;
    layer6_outputs(243) <= a and b;
    layer6_outputs(244) <= a;
    layer6_outputs(245) <= not b or a;
    layer6_outputs(246) <= not (a xor b);
    layer6_outputs(247) <= a xor b;
    layer6_outputs(248) <= a xor b;
    layer6_outputs(249) <= not b;
    layer6_outputs(250) <= b;
    layer6_outputs(251) <= b;
    layer6_outputs(252) <= not a;
    layer6_outputs(253) <= not a;
    layer6_outputs(254) <= not b;
    layer6_outputs(255) <= a xor b;
    layer6_outputs(256) <= b;
    layer6_outputs(257) <= not a or b;
    layer6_outputs(258) <= a xor b;
    layer6_outputs(259) <= not a;
    layer6_outputs(260) <= not b or a;
    layer6_outputs(261) <= not (a xor b);
    layer6_outputs(262) <= a and b;
    layer6_outputs(263) <= a and not b;
    layer6_outputs(264) <= not (a and b);
    layer6_outputs(265) <= a xor b;
    layer6_outputs(266) <= a;
    layer6_outputs(267) <= a or b;
    layer6_outputs(268) <= b;
    layer6_outputs(269) <= b;
    layer6_outputs(270) <= a;
    layer6_outputs(271) <= not (a xor b);
    layer6_outputs(272) <= a or b;
    layer6_outputs(273) <= b and not a;
    layer6_outputs(274) <= a;
    layer6_outputs(275) <= a;
    layer6_outputs(276) <= a;
    layer6_outputs(277) <= a xor b;
    layer6_outputs(278) <= a xor b;
    layer6_outputs(279) <= not a;
    layer6_outputs(280) <= a;
    layer6_outputs(281) <= not a;
    layer6_outputs(282) <= '0';
    layer6_outputs(283) <= b and not a;
    layer6_outputs(284) <= not (a xor b);
    layer6_outputs(285) <= a;
    layer6_outputs(286) <= not a;
    layer6_outputs(287) <= not b;
    layer6_outputs(288) <= not (a xor b);
    layer6_outputs(289) <= not a or b;
    layer6_outputs(290) <= b;
    layer6_outputs(291) <= not a;
    layer6_outputs(292) <= not a;
    layer6_outputs(293) <= not (a xor b);
    layer6_outputs(294) <= b and not a;
    layer6_outputs(295) <= a;
    layer6_outputs(296) <= a and b;
    layer6_outputs(297) <= not (a and b);
    layer6_outputs(298) <= a xor b;
    layer6_outputs(299) <= not (a xor b);
    layer6_outputs(300) <= a;
    layer6_outputs(301) <= a xor b;
    layer6_outputs(302) <= a and not b;
    layer6_outputs(303) <= not (a xor b);
    layer6_outputs(304) <= a or b;
    layer6_outputs(305) <= a;
    layer6_outputs(306) <= a and b;
    layer6_outputs(307) <= a;
    layer6_outputs(308) <= not a;
    layer6_outputs(309) <= not (a xor b);
    layer6_outputs(310) <= b;
    layer6_outputs(311) <= b;
    layer6_outputs(312) <= a and not b;
    layer6_outputs(313) <= not b;
    layer6_outputs(314) <= not b;
    layer6_outputs(315) <= not (a or b);
    layer6_outputs(316) <= a and not b;
    layer6_outputs(317) <= a xor b;
    layer6_outputs(318) <= a and not b;
    layer6_outputs(319) <= '0';
    layer6_outputs(320) <= not (a xor b);
    layer6_outputs(321) <= a;
    layer6_outputs(322) <= not a or b;
    layer6_outputs(323) <= not a;
    layer6_outputs(324) <= not b;
    layer6_outputs(325) <= not a;
    layer6_outputs(326) <= not (a xor b);
    layer6_outputs(327) <= not (a or b);
    layer6_outputs(328) <= not (a or b);
    layer6_outputs(329) <= a xor b;
    layer6_outputs(330) <= a xor b;
    layer6_outputs(331) <= a;
    layer6_outputs(332) <= not a or b;
    layer6_outputs(333) <= a;
    layer6_outputs(334) <= not a;
    layer6_outputs(335) <= not b;
    layer6_outputs(336) <= not (a xor b);
    layer6_outputs(337) <= a or b;
    layer6_outputs(338) <= not b;
    layer6_outputs(339) <= a and not b;
    layer6_outputs(340) <= a xor b;
    layer6_outputs(341) <= b;
    layer6_outputs(342) <= not (a and b);
    layer6_outputs(343) <= not a or b;
    layer6_outputs(344) <= b;
    layer6_outputs(345) <= not (a or b);
    layer6_outputs(346) <= a xor b;
    layer6_outputs(347) <= not (a xor b);
    layer6_outputs(348) <= a and not b;
    layer6_outputs(349) <= not b;
    layer6_outputs(350) <= a xor b;
    layer6_outputs(351) <= not b;
    layer6_outputs(352) <= a xor b;
    layer6_outputs(353) <= not a;
    layer6_outputs(354) <= a;
    layer6_outputs(355) <= not (a xor b);
    layer6_outputs(356) <= a xor b;
    layer6_outputs(357) <= b;
    layer6_outputs(358) <= not (a xor b);
    layer6_outputs(359) <= a xor b;
    layer6_outputs(360) <= a;
    layer6_outputs(361) <= a;
    layer6_outputs(362) <= a;
    layer6_outputs(363) <= a;
    layer6_outputs(364) <= not b;
    layer6_outputs(365) <= not b;
    layer6_outputs(366) <= not (a and b);
    layer6_outputs(367) <= b;
    layer6_outputs(368) <= b and not a;
    layer6_outputs(369) <= not b;
    layer6_outputs(370) <= a xor b;
    layer6_outputs(371) <= a;
    layer6_outputs(372) <= b;
    layer6_outputs(373) <= b;
    layer6_outputs(374) <= a xor b;
    layer6_outputs(375) <= not b;
    layer6_outputs(376) <= a xor b;
    layer6_outputs(377) <= a or b;
    layer6_outputs(378) <= not b;
    layer6_outputs(379) <= not (a or b);
    layer6_outputs(380) <= a xor b;
    layer6_outputs(381) <= a or b;
    layer6_outputs(382) <= b;
    layer6_outputs(383) <= not a;
    layer6_outputs(384) <= not a or b;
    layer6_outputs(385) <= b;
    layer6_outputs(386) <= b;
    layer6_outputs(387) <= not b;
    layer6_outputs(388) <= not a;
    layer6_outputs(389) <= not (a xor b);
    layer6_outputs(390) <= not b;
    layer6_outputs(391) <= not b or a;
    layer6_outputs(392) <= not b or a;
    layer6_outputs(393) <= b;
    layer6_outputs(394) <= not (a xor b);
    layer6_outputs(395) <= not a;
    layer6_outputs(396) <= a and not b;
    layer6_outputs(397) <= b;
    layer6_outputs(398) <= not b;
    layer6_outputs(399) <= not a;
    layer6_outputs(400) <= not a;
    layer6_outputs(401) <= not b or a;
    layer6_outputs(402) <= not (a or b);
    layer6_outputs(403) <= a and b;
    layer6_outputs(404) <= b and not a;
    layer6_outputs(405) <= not (a xor b);
    layer6_outputs(406) <= a and b;
    layer6_outputs(407) <= a xor b;
    layer6_outputs(408) <= not (a and b);
    layer6_outputs(409) <= not a or b;
    layer6_outputs(410) <= b;
    layer6_outputs(411) <= not (a xor b);
    layer6_outputs(412) <= not b or a;
    layer6_outputs(413) <= a or b;
    layer6_outputs(414) <= not (a xor b);
    layer6_outputs(415) <= a;
    layer6_outputs(416) <= not a;
    layer6_outputs(417) <= not a;
    layer6_outputs(418) <= not (a or b);
    layer6_outputs(419) <= not a;
    layer6_outputs(420) <= b and not a;
    layer6_outputs(421) <= a or b;
    layer6_outputs(422) <= b and not a;
    layer6_outputs(423) <= a and not b;
    layer6_outputs(424) <= a or b;
    layer6_outputs(425) <= a;
    layer6_outputs(426) <= b;
    layer6_outputs(427) <= a or b;
    layer6_outputs(428) <= a or b;
    layer6_outputs(429) <= not (a xor b);
    layer6_outputs(430) <= not a;
    layer6_outputs(431) <= not (a xor b);
    layer6_outputs(432) <= not a;
    layer6_outputs(433) <= a and b;
    layer6_outputs(434) <= b;
    layer6_outputs(435) <= not (a xor b);
    layer6_outputs(436) <= not (a xor b);
    layer6_outputs(437) <= a or b;
    layer6_outputs(438) <= a xor b;
    layer6_outputs(439) <= a;
    layer6_outputs(440) <= not a;
    layer6_outputs(441) <= not b;
    layer6_outputs(442) <= not b or a;
    layer6_outputs(443) <= not a;
    layer6_outputs(444) <= a;
    layer6_outputs(445) <= b and not a;
    layer6_outputs(446) <= not b;
    layer6_outputs(447) <= b;
    layer6_outputs(448) <= not b;
    layer6_outputs(449) <= b;
    layer6_outputs(450) <= not (a xor b);
    layer6_outputs(451) <= not b or a;
    layer6_outputs(452) <= b;
    layer6_outputs(453) <= b and not a;
    layer6_outputs(454) <= not b;
    layer6_outputs(455) <= a xor b;
    layer6_outputs(456) <= not b;
    layer6_outputs(457) <= a and b;
    layer6_outputs(458) <= a xor b;
    layer6_outputs(459) <= not b;
    layer6_outputs(460) <= not (a or b);
    layer6_outputs(461) <= a and b;
    layer6_outputs(462) <= not (a or b);
    layer6_outputs(463) <= a xor b;
    layer6_outputs(464) <= not a;
    layer6_outputs(465) <= not (a xor b);
    layer6_outputs(466) <= b;
    layer6_outputs(467) <= a;
    layer6_outputs(468) <= a;
    layer6_outputs(469) <= not a;
    layer6_outputs(470) <= a and not b;
    layer6_outputs(471) <= a;
    layer6_outputs(472) <= a xor b;
    layer6_outputs(473) <= not (a or b);
    layer6_outputs(474) <= a;
    layer6_outputs(475) <= a and b;
    layer6_outputs(476) <= b and not a;
    layer6_outputs(477) <= not (a xor b);
    layer6_outputs(478) <= a;
    layer6_outputs(479) <= b;
    layer6_outputs(480) <= a and not b;
    layer6_outputs(481) <= not b or a;
    layer6_outputs(482) <= a;
    layer6_outputs(483) <= a and not b;
    layer6_outputs(484) <= not b or a;
    layer6_outputs(485) <= a or b;
    layer6_outputs(486) <= not b;
    layer6_outputs(487) <= not (a xor b);
    layer6_outputs(488) <= a and b;
    layer6_outputs(489) <= not b;
    layer6_outputs(490) <= not b;
    layer6_outputs(491) <= not a or b;
    layer6_outputs(492) <= b;
    layer6_outputs(493) <= not a;
    layer6_outputs(494) <= not a or b;
    layer6_outputs(495) <= not (a or b);
    layer6_outputs(496) <= a;
    layer6_outputs(497) <= not (a xor b);
    layer6_outputs(498) <= a;
    layer6_outputs(499) <= b;
    layer6_outputs(500) <= not (a xor b);
    layer6_outputs(501) <= b and not a;
    layer6_outputs(502) <= not b;
    layer6_outputs(503) <= b;
    layer6_outputs(504) <= not a;
    layer6_outputs(505) <= not b;
    layer6_outputs(506) <= a;
    layer6_outputs(507) <= not a;
    layer6_outputs(508) <= not a;
    layer6_outputs(509) <= a xor b;
    layer6_outputs(510) <= a;
    layer6_outputs(511) <= b;
    layer6_outputs(512) <= a xor b;
    layer6_outputs(513) <= b;
    layer6_outputs(514) <= not (a xor b);
    layer6_outputs(515) <= a;
    layer6_outputs(516) <= a and b;
    layer6_outputs(517) <= not a;
    layer6_outputs(518) <= b;
    layer6_outputs(519) <= not a;
    layer6_outputs(520) <= a xor b;
    layer6_outputs(521) <= a and b;
    layer6_outputs(522) <= a and not b;
    layer6_outputs(523) <= '0';
    layer6_outputs(524) <= a;
    layer6_outputs(525) <= not a or b;
    layer6_outputs(526) <= a and not b;
    layer6_outputs(527) <= not b;
    layer6_outputs(528) <= a;
    layer6_outputs(529) <= a or b;
    layer6_outputs(530) <= not b or a;
    layer6_outputs(531) <= a;
    layer6_outputs(532) <= a;
    layer6_outputs(533) <= '1';
    layer6_outputs(534) <= not (a and b);
    layer6_outputs(535) <= not a;
    layer6_outputs(536) <= a or b;
    layer6_outputs(537) <= a or b;
    layer6_outputs(538) <= b;
    layer6_outputs(539) <= b;
    layer6_outputs(540) <= a xor b;
    layer6_outputs(541) <= a and b;
    layer6_outputs(542) <= a xor b;
    layer6_outputs(543) <= a xor b;
    layer6_outputs(544) <= a and not b;
    layer6_outputs(545) <= a and not b;
    layer6_outputs(546) <= not a;
    layer6_outputs(547) <= a xor b;
    layer6_outputs(548) <= b;
    layer6_outputs(549) <= b;
    layer6_outputs(550) <= not b;
    layer6_outputs(551) <= a or b;
    layer6_outputs(552) <= not b;
    layer6_outputs(553) <= not (a or b);
    layer6_outputs(554) <= a and b;
    layer6_outputs(555) <= not (a xor b);
    layer6_outputs(556) <= not (a xor b);
    layer6_outputs(557) <= b;
    layer6_outputs(558) <= a xor b;
    layer6_outputs(559) <= a;
    layer6_outputs(560) <= not b;
    layer6_outputs(561) <= b and not a;
    layer6_outputs(562) <= not (a and b);
    layer6_outputs(563) <= a or b;
    layer6_outputs(564) <= not (a or b);
    layer6_outputs(565) <= not b;
    layer6_outputs(566) <= not b or a;
    layer6_outputs(567) <= b;
    layer6_outputs(568) <= b;
    layer6_outputs(569) <= not (a xor b);
    layer6_outputs(570) <= not b or a;
    layer6_outputs(571) <= a;
    layer6_outputs(572) <= not a;
    layer6_outputs(573) <= not (a or b);
    layer6_outputs(574) <= b and not a;
    layer6_outputs(575) <= not b;
    layer6_outputs(576) <= not (a xor b);
    layer6_outputs(577) <= not (a xor b);
    layer6_outputs(578) <= a;
    layer6_outputs(579) <= not b;
    layer6_outputs(580) <= a xor b;
    layer6_outputs(581) <= b and not a;
    layer6_outputs(582) <= b;
    layer6_outputs(583) <= a;
    layer6_outputs(584) <= b and not a;
    layer6_outputs(585) <= not a or b;
    layer6_outputs(586) <= not a or b;
    layer6_outputs(587) <= not a;
    layer6_outputs(588) <= not a or b;
    layer6_outputs(589) <= not a or b;
    layer6_outputs(590) <= not (a and b);
    layer6_outputs(591) <= a xor b;
    layer6_outputs(592) <= b and not a;
    layer6_outputs(593) <= not (a xor b);
    layer6_outputs(594) <= b;
    layer6_outputs(595) <= not a;
    layer6_outputs(596) <= not a;
    layer6_outputs(597) <= a;
    layer6_outputs(598) <= not (a or b);
    layer6_outputs(599) <= a xor b;
    layer6_outputs(600) <= b;
    layer6_outputs(601) <= '1';
    layer6_outputs(602) <= not a;
    layer6_outputs(603) <= not a or b;
    layer6_outputs(604) <= not b or a;
    layer6_outputs(605) <= b;
    layer6_outputs(606) <= a and b;
    layer6_outputs(607) <= not b;
    layer6_outputs(608) <= not b;
    layer6_outputs(609) <= b and not a;
    layer6_outputs(610) <= a xor b;
    layer6_outputs(611) <= not (a or b);
    layer6_outputs(612) <= not (a and b);
    layer6_outputs(613) <= not b;
    layer6_outputs(614) <= not (a xor b);
    layer6_outputs(615) <= a and not b;
    layer6_outputs(616) <= b and not a;
    layer6_outputs(617) <= a xor b;
    layer6_outputs(618) <= a xor b;
    layer6_outputs(619) <= not b;
    layer6_outputs(620) <= not b;
    layer6_outputs(621) <= a xor b;
    layer6_outputs(622) <= not b or a;
    layer6_outputs(623) <= a;
    layer6_outputs(624) <= not a or b;
    layer6_outputs(625) <= b;
    layer6_outputs(626) <= a and b;
    layer6_outputs(627) <= a and not b;
    layer6_outputs(628) <= b and not a;
    layer6_outputs(629) <= '0';
    layer6_outputs(630) <= not (a xor b);
    layer6_outputs(631) <= a and not b;
    layer6_outputs(632) <= not a or b;
    layer6_outputs(633) <= not (a or b);
    layer6_outputs(634) <= b;
    layer6_outputs(635) <= not a;
    layer6_outputs(636) <= not (a and b);
    layer6_outputs(637) <= not a or b;
    layer6_outputs(638) <= not a or b;
    layer6_outputs(639) <= a;
    layer6_outputs(640) <= a;
    layer6_outputs(641) <= a xor b;
    layer6_outputs(642) <= a;
    layer6_outputs(643) <= not (a and b);
    layer6_outputs(644) <= not (a and b);
    layer6_outputs(645) <= a and not b;
    layer6_outputs(646) <= not b;
    layer6_outputs(647) <= not b;
    layer6_outputs(648) <= b and not a;
    layer6_outputs(649) <= a xor b;
    layer6_outputs(650) <= b and not a;
    layer6_outputs(651) <= not (a xor b);
    layer6_outputs(652) <= not b;
    layer6_outputs(653) <= a xor b;
    layer6_outputs(654) <= b;
    layer6_outputs(655) <= not b;
    layer6_outputs(656) <= a;
    layer6_outputs(657) <= b;
    layer6_outputs(658) <= not (a and b);
    layer6_outputs(659) <= a;
    layer6_outputs(660) <= not (a xor b);
    layer6_outputs(661) <= b;
    layer6_outputs(662) <= not a;
    layer6_outputs(663) <= not b or a;
    layer6_outputs(664) <= a or b;
    layer6_outputs(665) <= not (a xor b);
    layer6_outputs(666) <= not b;
    layer6_outputs(667) <= not a;
    layer6_outputs(668) <= not b;
    layer6_outputs(669) <= b;
    layer6_outputs(670) <= not a;
    layer6_outputs(671) <= not b or a;
    layer6_outputs(672) <= not b;
    layer6_outputs(673) <= not (a xor b);
    layer6_outputs(674) <= not (a xor b);
    layer6_outputs(675) <= not (a xor b);
    layer6_outputs(676) <= not (a xor b);
    layer6_outputs(677) <= not a;
    layer6_outputs(678) <= not b;
    layer6_outputs(679) <= not a or b;
    layer6_outputs(680) <= a or b;
    layer6_outputs(681) <= not b;
    layer6_outputs(682) <= b and not a;
    layer6_outputs(683) <= a and b;
    layer6_outputs(684) <= a xor b;
    layer6_outputs(685) <= not (a xor b);
    layer6_outputs(686) <= not a or b;
    layer6_outputs(687) <= not a;
    layer6_outputs(688) <= not a;
    layer6_outputs(689) <= not b;
    layer6_outputs(690) <= b;
    layer6_outputs(691) <= a;
    layer6_outputs(692) <= not (a xor b);
    layer6_outputs(693) <= a;
    layer6_outputs(694) <= not (a or b);
    layer6_outputs(695) <= b and not a;
    layer6_outputs(696) <= not b;
    layer6_outputs(697) <= not (a and b);
    layer6_outputs(698) <= not b or a;
    layer6_outputs(699) <= not b;
    layer6_outputs(700) <= a and b;
    layer6_outputs(701) <= not a;
    layer6_outputs(702) <= not b;
    layer6_outputs(703) <= not (a or b);
    layer6_outputs(704) <= not b;
    layer6_outputs(705) <= a and not b;
    layer6_outputs(706) <= not b;
    layer6_outputs(707) <= not b;
    layer6_outputs(708) <= not b or a;
    layer6_outputs(709) <= not b or a;
    layer6_outputs(710) <= a or b;
    layer6_outputs(711) <= a xor b;
    layer6_outputs(712) <= not (a xor b);
    layer6_outputs(713) <= not b;
    layer6_outputs(714) <= not (a and b);
    layer6_outputs(715) <= not b;
    layer6_outputs(716) <= not a;
    layer6_outputs(717) <= not (a xor b);
    layer6_outputs(718) <= not (a xor b);
    layer6_outputs(719) <= not b;
    layer6_outputs(720) <= not (a xor b);
    layer6_outputs(721) <= '0';
    layer6_outputs(722) <= a xor b;
    layer6_outputs(723) <= b;
    layer6_outputs(724) <= b;
    layer6_outputs(725) <= not b;
    layer6_outputs(726) <= a and not b;
    layer6_outputs(727) <= not b;
    layer6_outputs(728) <= not b;
    layer6_outputs(729) <= not b or a;
    layer6_outputs(730) <= not a;
    layer6_outputs(731) <= a;
    layer6_outputs(732) <= a;
    layer6_outputs(733) <= b;
    layer6_outputs(734) <= a xor b;
    layer6_outputs(735) <= a and not b;
    layer6_outputs(736) <= not b;
    layer6_outputs(737) <= a;
    layer6_outputs(738) <= b;
    layer6_outputs(739) <= a xor b;
    layer6_outputs(740) <= b;
    layer6_outputs(741) <= a;
    layer6_outputs(742) <= a and b;
    layer6_outputs(743) <= b;
    layer6_outputs(744) <= not a or b;
    layer6_outputs(745) <= a xor b;
    layer6_outputs(746) <= not b;
    layer6_outputs(747) <= a xor b;
    layer6_outputs(748) <= b;
    layer6_outputs(749) <= not a;
    layer6_outputs(750) <= not (a xor b);
    layer6_outputs(751) <= not (a xor b);
    layer6_outputs(752) <= not a;
    layer6_outputs(753) <= a;
    layer6_outputs(754) <= not a;
    layer6_outputs(755) <= a or b;
    layer6_outputs(756) <= a and not b;
    layer6_outputs(757) <= b;
    layer6_outputs(758) <= not a;
    layer6_outputs(759) <= a;
    layer6_outputs(760) <= not (a xor b);
    layer6_outputs(761) <= not b;
    layer6_outputs(762) <= not a;
    layer6_outputs(763) <= b and not a;
    layer6_outputs(764) <= b;
    layer6_outputs(765) <= not b;
    layer6_outputs(766) <= a;
    layer6_outputs(767) <= not b;
    layer6_outputs(768) <= b;
    layer6_outputs(769) <= '1';
    layer6_outputs(770) <= a or b;
    layer6_outputs(771) <= not a or b;
    layer6_outputs(772) <= not b or a;
    layer6_outputs(773) <= not b;
    layer6_outputs(774) <= a;
    layer6_outputs(775) <= a;
    layer6_outputs(776) <= a xor b;
    layer6_outputs(777) <= not b;
    layer6_outputs(778) <= not a or b;
    layer6_outputs(779) <= a;
    layer6_outputs(780) <= not (a xor b);
    layer6_outputs(781) <= a and b;
    layer6_outputs(782) <= not (a and b);
    layer6_outputs(783) <= not a;
    layer6_outputs(784) <= not b;
    layer6_outputs(785) <= b;
    layer6_outputs(786) <= b;
    layer6_outputs(787) <= not a or b;
    layer6_outputs(788) <= a;
    layer6_outputs(789) <= b;
    layer6_outputs(790) <= a;
    layer6_outputs(791) <= not b;
    layer6_outputs(792) <= a xor b;
    layer6_outputs(793) <= not (a or b);
    layer6_outputs(794) <= not a;
    layer6_outputs(795) <= b;
    layer6_outputs(796) <= b;
    layer6_outputs(797) <= a;
    layer6_outputs(798) <= a xor b;
    layer6_outputs(799) <= not a or b;
    layer6_outputs(800) <= not (a and b);
    layer6_outputs(801) <= not (a xor b);
    layer6_outputs(802) <= a or b;
    layer6_outputs(803) <= not b;
    layer6_outputs(804) <= a or b;
    layer6_outputs(805) <= a xor b;
    layer6_outputs(806) <= a or b;
    layer6_outputs(807) <= a xor b;
    layer6_outputs(808) <= not a;
    layer6_outputs(809) <= not b;
    layer6_outputs(810) <= not a or b;
    layer6_outputs(811) <= not b;
    layer6_outputs(812) <= b;
    layer6_outputs(813) <= not (a and b);
    layer6_outputs(814) <= not (a or b);
    layer6_outputs(815) <= a or b;
    layer6_outputs(816) <= not b;
    layer6_outputs(817) <= not a;
    layer6_outputs(818) <= a xor b;
    layer6_outputs(819) <= b and not a;
    layer6_outputs(820) <= a xor b;
    layer6_outputs(821) <= a or b;
    layer6_outputs(822) <= '1';
    layer6_outputs(823) <= not a;
    layer6_outputs(824) <= not a;
    layer6_outputs(825) <= not (a and b);
    layer6_outputs(826) <= b and not a;
    layer6_outputs(827) <= a xor b;
    layer6_outputs(828) <= not (a xor b);
    layer6_outputs(829) <= a xor b;
    layer6_outputs(830) <= not (a xor b);
    layer6_outputs(831) <= a;
    layer6_outputs(832) <= not a;
    layer6_outputs(833) <= b;
    layer6_outputs(834) <= '1';
    layer6_outputs(835) <= a and not b;
    layer6_outputs(836) <= not b;
    layer6_outputs(837) <= b;
    layer6_outputs(838) <= b and not a;
    layer6_outputs(839) <= a or b;
    layer6_outputs(840) <= not a;
    layer6_outputs(841) <= a;
    layer6_outputs(842) <= a or b;
    layer6_outputs(843) <= not (a and b);
    layer6_outputs(844) <= not a;
    layer6_outputs(845) <= a;
    layer6_outputs(846) <= a;
    layer6_outputs(847) <= b;
    layer6_outputs(848) <= a;
    layer6_outputs(849) <= a;
    layer6_outputs(850) <= b;
    layer6_outputs(851) <= not a;
    layer6_outputs(852) <= a;
    layer6_outputs(853) <= not (a and b);
    layer6_outputs(854) <= not b;
    layer6_outputs(855) <= not b or a;
    layer6_outputs(856) <= a;
    layer6_outputs(857) <= a xor b;
    layer6_outputs(858) <= not (a or b);
    layer6_outputs(859) <= a and not b;
    layer6_outputs(860) <= not b or a;
    layer6_outputs(861) <= not (a xor b);
    layer6_outputs(862) <= not a or b;
    layer6_outputs(863) <= not (a xor b);
    layer6_outputs(864) <= b;
    layer6_outputs(865) <= not (a or b);
    layer6_outputs(866) <= not (a xor b);
    layer6_outputs(867) <= a and not b;
    layer6_outputs(868) <= not (a and b);
    layer6_outputs(869) <= not b or a;
    layer6_outputs(870) <= b;
    layer6_outputs(871) <= b;
    layer6_outputs(872) <= b;
    layer6_outputs(873) <= a xor b;
    layer6_outputs(874) <= not (a xor b);
    layer6_outputs(875) <= not a;
    layer6_outputs(876) <= a;
    layer6_outputs(877) <= a;
    layer6_outputs(878) <= a;
    layer6_outputs(879) <= not (a or b);
    layer6_outputs(880) <= not b or a;
    layer6_outputs(881) <= a;
    layer6_outputs(882) <= a and b;
    layer6_outputs(883) <= a xor b;
    layer6_outputs(884) <= a or b;
    layer6_outputs(885) <= not b;
    layer6_outputs(886) <= a xor b;
    layer6_outputs(887) <= a xor b;
    layer6_outputs(888) <= b;
    layer6_outputs(889) <= not (a xor b);
    layer6_outputs(890) <= a and b;
    layer6_outputs(891) <= a and not b;
    layer6_outputs(892) <= not a;
    layer6_outputs(893) <= a and not b;
    layer6_outputs(894) <= not (a or b);
    layer6_outputs(895) <= not (a and b);
    layer6_outputs(896) <= a;
    layer6_outputs(897) <= a xor b;
    layer6_outputs(898) <= b;
    layer6_outputs(899) <= a and not b;
    layer6_outputs(900) <= a and not b;
    layer6_outputs(901) <= b;
    layer6_outputs(902) <= not b;
    layer6_outputs(903) <= not (a xor b);
    layer6_outputs(904) <= a;
    layer6_outputs(905) <= not b;
    layer6_outputs(906) <= not a;
    layer6_outputs(907) <= b and not a;
    layer6_outputs(908) <= b and not a;
    layer6_outputs(909) <= a xor b;
    layer6_outputs(910) <= b;
    layer6_outputs(911) <= not (a xor b);
    layer6_outputs(912) <= b;
    layer6_outputs(913) <= not (a and b);
    layer6_outputs(914) <= a;
    layer6_outputs(915) <= not a or b;
    layer6_outputs(916) <= not a;
    layer6_outputs(917) <= not (a xor b);
    layer6_outputs(918) <= b;
    layer6_outputs(919) <= not b or a;
    layer6_outputs(920) <= a;
    layer6_outputs(921) <= a and not b;
    layer6_outputs(922) <= b;
    layer6_outputs(923) <= not b;
    layer6_outputs(924) <= not (a or b);
    layer6_outputs(925) <= a and not b;
    layer6_outputs(926) <= a;
    layer6_outputs(927) <= b;
    layer6_outputs(928) <= a xor b;
    layer6_outputs(929) <= a and not b;
    layer6_outputs(930) <= a;
    layer6_outputs(931) <= not (a or b);
    layer6_outputs(932) <= not b;
    layer6_outputs(933) <= a xor b;
    layer6_outputs(934) <= not (a xor b);
    layer6_outputs(935) <= not a or b;
    layer6_outputs(936) <= b and not a;
    layer6_outputs(937) <= not (a and b);
    layer6_outputs(938) <= not b;
    layer6_outputs(939) <= not a or b;
    layer6_outputs(940) <= b;
    layer6_outputs(941) <= not a;
    layer6_outputs(942) <= a and b;
    layer6_outputs(943) <= not a;
    layer6_outputs(944) <= not b or a;
    layer6_outputs(945) <= not (a xor b);
    layer6_outputs(946) <= a and b;
    layer6_outputs(947) <= a xor b;
    layer6_outputs(948) <= a or b;
    layer6_outputs(949) <= not b or a;
    layer6_outputs(950) <= not a;
    layer6_outputs(951) <= not b;
    layer6_outputs(952) <= a and b;
    layer6_outputs(953) <= not (a or b);
    layer6_outputs(954) <= not a;
    layer6_outputs(955) <= not (a xor b);
    layer6_outputs(956) <= not a;
    layer6_outputs(957) <= not b;
    layer6_outputs(958) <= not a;
    layer6_outputs(959) <= a;
    layer6_outputs(960) <= a;
    layer6_outputs(961) <= b;
    layer6_outputs(962) <= not (a xor b);
    layer6_outputs(963) <= a;
    layer6_outputs(964) <= b;
    layer6_outputs(965) <= a xor b;
    layer6_outputs(966) <= b;
    layer6_outputs(967) <= not b;
    layer6_outputs(968) <= not (a xor b);
    layer6_outputs(969) <= a or b;
    layer6_outputs(970) <= a and b;
    layer6_outputs(971) <= a and not b;
    layer6_outputs(972) <= b and not a;
    layer6_outputs(973) <= b;
    layer6_outputs(974) <= not a;
    layer6_outputs(975) <= b;
    layer6_outputs(976) <= not a;
    layer6_outputs(977) <= a xor b;
    layer6_outputs(978) <= not a;
    layer6_outputs(979) <= not a;
    layer6_outputs(980) <= not (a xor b);
    layer6_outputs(981) <= not a;
    layer6_outputs(982) <= b and not a;
    layer6_outputs(983) <= not b;
    layer6_outputs(984) <= not (a xor b);
    layer6_outputs(985) <= b and not a;
    layer6_outputs(986) <= a;
    layer6_outputs(987) <= not (a or b);
    layer6_outputs(988) <= a and b;
    layer6_outputs(989) <= not a or b;
    layer6_outputs(990) <= not b;
    layer6_outputs(991) <= not (a and b);
    layer6_outputs(992) <= not b;
    layer6_outputs(993) <= not a;
    layer6_outputs(994) <= a or b;
    layer6_outputs(995) <= not (a and b);
    layer6_outputs(996) <= not (a or b);
    layer6_outputs(997) <= a and b;
    layer6_outputs(998) <= a xor b;
    layer6_outputs(999) <= a xor b;
    layer6_outputs(1000) <= not (a and b);
    layer6_outputs(1001) <= a or b;
    layer6_outputs(1002) <= b;
    layer6_outputs(1003) <= b and not a;
    layer6_outputs(1004) <= a or b;
    layer6_outputs(1005) <= not a or b;
    layer6_outputs(1006) <= a or b;
    layer6_outputs(1007) <= a;
    layer6_outputs(1008) <= not a or b;
    layer6_outputs(1009) <= a;
    layer6_outputs(1010) <= a xor b;
    layer6_outputs(1011) <= a and not b;
    layer6_outputs(1012) <= not (a xor b);
    layer6_outputs(1013) <= not (a xor b);
    layer6_outputs(1014) <= not a;
    layer6_outputs(1015) <= not a;
    layer6_outputs(1016) <= not (a xor b);
    layer6_outputs(1017) <= a xor b;
    layer6_outputs(1018) <= b and not a;
    layer6_outputs(1019) <= not (a xor b);
    layer6_outputs(1020) <= not (a and b);
    layer6_outputs(1021) <= b;
    layer6_outputs(1022) <= a and b;
    layer6_outputs(1023) <= not b or a;
    layer6_outputs(1024) <= not a;
    layer6_outputs(1025) <= a or b;
    layer6_outputs(1026) <= b;
    layer6_outputs(1027) <= a;
    layer6_outputs(1028) <= a or b;
    layer6_outputs(1029) <= a and b;
    layer6_outputs(1030) <= a;
    layer6_outputs(1031) <= not (a or b);
    layer6_outputs(1032) <= not (a xor b);
    layer6_outputs(1033) <= b;
    layer6_outputs(1034) <= not (a xor b);
    layer6_outputs(1035) <= not b or a;
    layer6_outputs(1036) <= a and not b;
    layer6_outputs(1037) <= a;
    layer6_outputs(1038) <= a xor b;
    layer6_outputs(1039) <= b;
    layer6_outputs(1040) <= b and not a;
    layer6_outputs(1041) <= not b or a;
    layer6_outputs(1042) <= not a;
    layer6_outputs(1043) <= not (a xor b);
    layer6_outputs(1044) <= not a;
    layer6_outputs(1045) <= not a;
    layer6_outputs(1046) <= not (a xor b);
    layer6_outputs(1047) <= not (a or b);
    layer6_outputs(1048) <= not (a and b);
    layer6_outputs(1049) <= not a;
    layer6_outputs(1050) <= a and not b;
    layer6_outputs(1051) <= b;
    layer6_outputs(1052) <= not b or a;
    layer6_outputs(1053) <= not a or b;
    layer6_outputs(1054) <= a xor b;
    layer6_outputs(1055) <= b;
    layer6_outputs(1056) <= not (a or b);
    layer6_outputs(1057) <= not (a xor b);
    layer6_outputs(1058) <= b;
    layer6_outputs(1059) <= not a;
    layer6_outputs(1060) <= a;
    layer6_outputs(1061) <= not (a xor b);
    layer6_outputs(1062) <= b and not a;
    layer6_outputs(1063) <= a and b;
    layer6_outputs(1064) <= b;
    layer6_outputs(1065) <= not b;
    layer6_outputs(1066) <= not (a and b);
    layer6_outputs(1067) <= not b;
    layer6_outputs(1068) <= a and not b;
    layer6_outputs(1069) <= not (a xor b);
    layer6_outputs(1070) <= a xor b;
    layer6_outputs(1071) <= not a;
    layer6_outputs(1072) <= not b;
    layer6_outputs(1073) <= a xor b;
    layer6_outputs(1074) <= not a;
    layer6_outputs(1075) <= b;
    layer6_outputs(1076) <= a and not b;
    layer6_outputs(1077) <= not a or b;
    layer6_outputs(1078) <= a xor b;
    layer6_outputs(1079) <= a;
    layer6_outputs(1080) <= b;
    layer6_outputs(1081) <= not a;
    layer6_outputs(1082) <= not (a xor b);
    layer6_outputs(1083) <= not (a or b);
    layer6_outputs(1084) <= not a;
    layer6_outputs(1085) <= not b;
    layer6_outputs(1086) <= not b or a;
    layer6_outputs(1087) <= not a or b;
    layer6_outputs(1088) <= a xor b;
    layer6_outputs(1089) <= not b;
    layer6_outputs(1090) <= not (a xor b);
    layer6_outputs(1091) <= a;
    layer6_outputs(1092) <= a xor b;
    layer6_outputs(1093) <= not (a and b);
    layer6_outputs(1094) <= b;
    layer6_outputs(1095) <= b and not a;
    layer6_outputs(1096) <= a and not b;
    layer6_outputs(1097) <= not a or b;
    layer6_outputs(1098) <= a and b;
    layer6_outputs(1099) <= a and b;
    layer6_outputs(1100) <= a and not b;
    layer6_outputs(1101) <= not a;
    layer6_outputs(1102) <= b;
    layer6_outputs(1103) <= b and not a;
    layer6_outputs(1104) <= b;
    layer6_outputs(1105) <= b;
    layer6_outputs(1106) <= not (a xor b);
    layer6_outputs(1107) <= not a or b;
    layer6_outputs(1108) <= not (a or b);
    layer6_outputs(1109) <= not (a xor b);
    layer6_outputs(1110) <= not b;
    layer6_outputs(1111) <= not b;
    layer6_outputs(1112) <= a xor b;
    layer6_outputs(1113) <= not a;
    layer6_outputs(1114) <= a xor b;
    layer6_outputs(1115) <= b;
    layer6_outputs(1116) <= not (a xor b);
    layer6_outputs(1117) <= not b;
    layer6_outputs(1118) <= a xor b;
    layer6_outputs(1119) <= a;
    layer6_outputs(1120) <= not a;
    layer6_outputs(1121) <= a and not b;
    layer6_outputs(1122) <= b;
    layer6_outputs(1123) <= a or b;
    layer6_outputs(1124) <= a xor b;
    layer6_outputs(1125) <= a xor b;
    layer6_outputs(1126) <= a and b;
    layer6_outputs(1127) <= a xor b;
    layer6_outputs(1128) <= a and b;
    layer6_outputs(1129) <= b and not a;
    layer6_outputs(1130) <= a;
    layer6_outputs(1131) <= a or b;
    layer6_outputs(1132) <= not (a or b);
    layer6_outputs(1133) <= b and not a;
    layer6_outputs(1134) <= not (a or b);
    layer6_outputs(1135) <= not (a xor b);
    layer6_outputs(1136) <= a and not b;
    layer6_outputs(1137) <= b;
    layer6_outputs(1138) <= a;
    layer6_outputs(1139) <= a xor b;
    layer6_outputs(1140) <= not (a xor b);
    layer6_outputs(1141) <= not (a and b);
    layer6_outputs(1142) <= a;
    layer6_outputs(1143) <= b;
    layer6_outputs(1144) <= b;
    layer6_outputs(1145) <= b;
    layer6_outputs(1146) <= not (a or b);
    layer6_outputs(1147) <= not (a or b);
    layer6_outputs(1148) <= not b;
    layer6_outputs(1149) <= not b;
    layer6_outputs(1150) <= not (a or b);
    layer6_outputs(1151) <= a and not b;
    layer6_outputs(1152) <= not a or b;
    layer6_outputs(1153) <= a xor b;
    layer6_outputs(1154) <= not b;
    layer6_outputs(1155) <= not b;
    layer6_outputs(1156) <= a and not b;
    layer6_outputs(1157) <= not a;
    layer6_outputs(1158) <= a xor b;
    layer6_outputs(1159) <= a;
    layer6_outputs(1160) <= b and not a;
    layer6_outputs(1161) <= b;
    layer6_outputs(1162) <= a xor b;
    layer6_outputs(1163) <= a xor b;
    layer6_outputs(1164) <= b and not a;
    layer6_outputs(1165) <= a and b;
    layer6_outputs(1166) <= a and b;
    layer6_outputs(1167) <= b;
    layer6_outputs(1168) <= not b or a;
    layer6_outputs(1169) <= not b;
    layer6_outputs(1170) <= not a or b;
    layer6_outputs(1171) <= not b;
    layer6_outputs(1172) <= a and b;
    layer6_outputs(1173) <= not (a or b);
    layer6_outputs(1174) <= b;
    layer6_outputs(1175) <= a;
    layer6_outputs(1176) <= not a;
    layer6_outputs(1177) <= b;
    layer6_outputs(1178) <= a xor b;
    layer6_outputs(1179) <= not b or a;
    layer6_outputs(1180) <= a and b;
    layer6_outputs(1181) <= a xor b;
    layer6_outputs(1182) <= not a;
    layer6_outputs(1183) <= not a;
    layer6_outputs(1184) <= not b;
    layer6_outputs(1185) <= not a or b;
    layer6_outputs(1186) <= not b;
    layer6_outputs(1187) <= a and b;
    layer6_outputs(1188) <= not (a or b);
    layer6_outputs(1189) <= b;
    layer6_outputs(1190) <= a or b;
    layer6_outputs(1191) <= not (a and b);
    layer6_outputs(1192) <= a or b;
    layer6_outputs(1193) <= not (a xor b);
    layer6_outputs(1194) <= a;
    layer6_outputs(1195) <= a xor b;
    layer6_outputs(1196) <= not a or b;
    layer6_outputs(1197) <= not (a xor b);
    layer6_outputs(1198) <= not a or b;
    layer6_outputs(1199) <= not (a or b);
    layer6_outputs(1200) <= not a;
    layer6_outputs(1201) <= a or b;
    layer6_outputs(1202) <= b;
    layer6_outputs(1203) <= not (a and b);
    layer6_outputs(1204) <= a;
    layer6_outputs(1205) <= not b;
    layer6_outputs(1206) <= a xor b;
    layer6_outputs(1207) <= b;
    layer6_outputs(1208) <= not (a xor b);
    layer6_outputs(1209) <= a and not b;
    layer6_outputs(1210) <= not (a xor b);
    layer6_outputs(1211) <= not b;
    layer6_outputs(1212) <= not b;
    layer6_outputs(1213) <= not b;
    layer6_outputs(1214) <= not (a and b);
    layer6_outputs(1215) <= not a or b;
    layer6_outputs(1216) <= not b;
    layer6_outputs(1217) <= not (a and b);
    layer6_outputs(1218) <= not a;
    layer6_outputs(1219) <= a or b;
    layer6_outputs(1220) <= not a or b;
    layer6_outputs(1221) <= b and not a;
    layer6_outputs(1222) <= a;
    layer6_outputs(1223) <= b;
    layer6_outputs(1224) <= b and not a;
    layer6_outputs(1225) <= not b;
    layer6_outputs(1226) <= not b or a;
    layer6_outputs(1227) <= b and not a;
    layer6_outputs(1228) <= not (a xor b);
    layer6_outputs(1229) <= not a or b;
    layer6_outputs(1230) <= b and not a;
    layer6_outputs(1231) <= not (a and b);
    layer6_outputs(1232) <= not b;
    layer6_outputs(1233) <= b;
    layer6_outputs(1234) <= a;
    layer6_outputs(1235) <= a and b;
    layer6_outputs(1236) <= a and not b;
    layer6_outputs(1237) <= a and not b;
    layer6_outputs(1238) <= not b or a;
    layer6_outputs(1239) <= not (a and b);
    layer6_outputs(1240) <= not (a and b);
    layer6_outputs(1241) <= not b or a;
    layer6_outputs(1242) <= not b;
    layer6_outputs(1243) <= a;
    layer6_outputs(1244) <= not a;
    layer6_outputs(1245) <= not (a and b);
    layer6_outputs(1246) <= not b;
    layer6_outputs(1247) <= a and b;
    layer6_outputs(1248) <= a and b;
    layer6_outputs(1249) <= a and not b;
    layer6_outputs(1250) <= not (a and b);
    layer6_outputs(1251) <= a xor b;
    layer6_outputs(1252) <= not a or b;
    layer6_outputs(1253) <= not (a xor b);
    layer6_outputs(1254) <= a xor b;
    layer6_outputs(1255) <= not (a xor b);
    layer6_outputs(1256) <= not a;
    layer6_outputs(1257) <= b;
    layer6_outputs(1258) <= b;
    layer6_outputs(1259) <= not (a or b);
    layer6_outputs(1260) <= not (a or b);
    layer6_outputs(1261) <= a xor b;
    layer6_outputs(1262) <= a xor b;
    layer6_outputs(1263) <= not a or b;
    layer6_outputs(1264) <= not a;
    layer6_outputs(1265) <= a;
    layer6_outputs(1266) <= a xor b;
    layer6_outputs(1267) <= not b or a;
    layer6_outputs(1268) <= not b;
    layer6_outputs(1269) <= '0';
    layer6_outputs(1270) <= not b;
    layer6_outputs(1271) <= not a;
    layer6_outputs(1272) <= not a;
    layer6_outputs(1273) <= not a;
    layer6_outputs(1274) <= not b;
    layer6_outputs(1275) <= not b;
    layer6_outputs(1276) <= a and b;
    layer6_outputs(1277) <= a xor b;
    layer6_outputs(1278) <= not a or b;
    layer6_outputs(1279) <= '0';
    layer6_outputs(1280) <= not a;
    layer6_outputs(1281) <= a xor b;
    layer6_outputs(1282) <= a;
    layer6_outputs(1283) <= not b or a;
    layer6_outputs(1284) <= not (a xor b);
    layer6_outputs(1285) <= not a;
    layer6_outputs(1286) <= not b;
    layer6_outputs(1287) <= a and b;
    layer6_outputs(1288) <= not a or b;
    layer6_outputs(1289) <= not b;
    layer6_outputs(1290) <= b;
    layer6_outputs(1291) <= a;
    layer6_outputs(1292) <= not a;
    layer6_outputs(1293) <= a xor b;
    layer6_outputs(1294) <= a and not b;
    layer6_outputs(1295) <= b;
    layer6_outputs(1296) <= a and b;
    layer6_outputs(1297) <= a and b;
    layer6_outputs(1298) <= not b;
    layer6_outputs(1299) <= not b;
    layer6_outputs(1300) <= a;
    layer6_outputs(1301) <= not a or b;
    layer6_outputs(1302) <= not b;
    layer6_outputs(1303) <= not a;
    layer6_outputs(1304) <= not (a xor b);
    layer6_outputs(1305) <= a and not b;
    layer6_outputs(1306) <= b and not a;
    layer6_outputs(1307) <= a;
    layer6_outputs(1308) <= not b;
    layer6_outputs(1309) <= not a or b;
    layer6_outputs(1310) <= not b;
    layer6_outputs(1311) <= a xor b;
    layer6_outputs(1312) <= a and not b;
    layer6_outputs(1313) <= not (a or b);
    layer6_outputs(1314) <= b;
    layer6_outputs(1315) <= a;
    layer6_outputs(1316) <= not (a and b);
    layer6_outputs(1317) <= not b;
    layer6_outputs(1318) <= not a or b;
    layer6_outputs(1319) <= a and not b;
    layer6_outputs(1320) <= a;
    layer6_outputs(1321) <= not (a or b);
    layer6_outputs(1322) <= not b;
    layer6_outputs(1323) <= not b;
    layer6_outputs(1324) <= not (a xor b);
    layer6_outputs(1325) <= a xor b;
    layer6_outputs(1326) <= not (a and b);
    layer6_outputs(1327) <= a xor b;
    layer6_outputs(1328) <= not (a and b);
    layer6_outputs(1329) <= not (a or b);
    layer6_outputs(1330) <= a and not b;
    layer6_outputs(1331) <= a;
    layer6_outputs(1332) <= not (a xor b);
    layer6_outputs(1333) <= a xor b;
    layer6_outputs(1334) <= b;
    layer6_outputs(1335) <= not (a xor b);
    layer6_outputs(1336) <= b and not a;
    layer6_outputs(1337) <= a and not b;
    layer6_outputs(1338) <= a xor b;
    layer6_outputs(1339) <= not a;
    layer6_outputs(1340) <= not a;
    layer6_outputs(1341) <= a xor b;
    layer6_outputs(1342) <= a and not b;
    layer6_outputs(1343) <= a xor b;
    layer6_outputs(1344) <= not a;
    layer6_outputs(1345) <= b;
    layer6_outputs(1346) <= not b;
    layer6_outputs(1347) <= a xor b;
    layer6_outputs(1348) <= a;
    layer6_outputs(1349) <= not (a xor b);
    layer6_outputs(1350) <= not b or a;
    layer6_outputs(1351) <= not a;
    layer6_outputs(1352) <= not (a xor b);
    layer6_outputs(1353) <= not (a xor b);
    layer6_outputs(1354) <= not b;
    layer6_outputs(1355) <= not a;
    layer6_outputs(1356) <= a xor b;
    layer6_outputs(1357) <= b and not a;
    layer6_outputs(1358) <= a xor b;
    layer6_outputs(1359) <= b;
    layer6_outputs(1360) <= b;
    layer6_outputs(1361) <= a xor b;
    layer6_outputs(1362) <= not (a or b);
    layer6_outputs(1363) <= a and b;
    layer6_outputs(1364) <= not (a xor b);
    layer6_outputs(1365) <= not b or a;
    layer6_outputs(1366) <= a and b;
    layer6_outputs(1367) <= a and not b;
    layer6_outputs(1368) <= not b;
    layer6_outputs(1369) <= not b;
    layer6_outputs(1370) <= not a;
    layer6_outputs(1371) <= a;
    layer6_outputs(1372) <= a and not b;
    layer6_outputs(1373) <= a or b;
    layer6_outputs(1374) <= not a or b;
    layer6_outputs(1375) <= not (a xor b);
    layer6_outputs(1376) <= not b or a;
    layer6_outputs(1377) <= b;
    layer6_outputs(1378) <= not b;
    layer6_outputs(1379) <= a and not b;
    layer6_outputs(1380) <= a and not b;
    layer6_outputs(1381) <= not (a xor b);
    layer6_outputs(1382) <= a or b;
    layer6_outputs(1383) <= b;
    layer6_outputs(1384) <= b and not a;
    layer6_outputs(1385) <= a xor b;
    layer6_outputs(1386) <= not (a xor b);
    layer6_outputs(1387) <= b;
    layer6_outputs(1388) <= b;
    layer6_outputs(1389) <= a;
    layer6_outputs(1390) <= not a;
    layer6_outputs(1391) <= not b;
    layer6_outputs(1392) <= a and b;
    layer6_outputs(1393) <= b;
    layer6_outputs(1394) <= a;
    layer6_outputs(1395) <= b;
    layer6_outputs(1396) <= a or b;
    layer6_outputs(1397) <= not b;
    layer6_outputs(1398) <= not b;
    layer6_outputs(1399) <= not (a xor b);
    layer6_outputs(1400) <= a;
    layer6_outputs(1401) <= b and not a;
    layer6_outputs(1402) <= a;
    layer6_outputs(1403) <= not b;
    layer6_outputs(1404) <= not b;
    layer6_outputs(1405) <= b;
    layer6_outputs(1406) <= not b;
    layer6_outputs(1407) <= a or b;
    layer6_outputs(1408) <= not (a xor b);
    layer6_outputs(1409) <= not b;
    layer6_outputs(1410) <= not (a and b);
    layer6_outputs(1411) <= not a or b;
    layer6_outputs(1412) <= not (a xor b);
    layer6_outputs(1413) <= a xor b;
    layer6_outputs(1414) <= b;
    layer6_outputs(1415) <= a or b;
    layer6_outputs(1416) <= b;
    layer6_outputs(1417) <= not (a xor b);
    layer6_outputs(1418) <= a;
    layer6_outputs(1419) <= not b;
    layer6_outputs(1420) <= not (a xor b);
    layer6_outputs(1421) <= not (a and b);
    layer6_outputs(1422) <= not (a xor b);
    layer6_outputs(1423) <= not (a xor b);
    layer6_outputs(1424) <= not b or a;
    layer6_outputs(1425) <= b and not a;
    layer6_outputs(1426) <= not b;
    layer6_outputs(1427) <= not (a xor b);
    layer6_outputs(1428) <= a and not b;
    layer6_outputs(1429) <= not (a or b);
    layer6_outputs(1430) <= a or b;
    layer6_outputs(1431) <= a or b;
    layer6_outputs(1432) <= not a or b;
    layer6_outputs(1433) <= not (a xor b);
    layer6_outputs(1434) <= not a;
    layer6_outputs(1435) <= not a;
    layer6_outputs(1436) <= not b;
    layer6_outputs(1437) <= a or b;
    layer6_outputs(1438) <= not a;
    layer6_outputs(1439) <= a or b;
    layer6_outputs(1440) <= a and not b;
    layer6_outputs(1441) <= a xor b;
    layer6_outputs(1442) <= not (a or b);
    layer6_outputs(1443) <= b;
    layer6_outputs(1444) <= not a;
    layer6_outputs(1445) <= a or b;
    layer6_outputs(1446) <= '1';
    layer6_outputs(1447) <= a;
    layer6_outputs(1448) <= not b;
    layer6_outputs(1449) <= b;
    layer6_outputs(1450) <= b and not a;
    layer6_outputs(1451) <= not b;
    layer6_outputs(1452) <= a xor b;
    layer6_outputs(1453) <= not (a xor b);
    layer6_outputs(1454) <= b and not a;
    layer6_outputs(1455) <= not a;
    layer6_outputs(1456) <= a;
    layer6_outputs(1457) <= not b;
    layer6_outputs(1458) <= not b;
    layer6_outputs(1459) <= b and not a;
    layer6_outputs(1460) <= not a or b;
    layer6_outputs(1461) <= not (a xor b);
    layer6_outputs(1462) <= not (a xor b);
    layer6_outputs(1463) <= a xor b;
    layer6_outputs(1464) <= b;
    layer6_outputs(1465) <= b and not a;
    layer6_outputs(1466) <= not a;
    layer6_outputs(1467) <= a or b;
    layer6_outputs(1468) <= a and not b;
    layer6_outputs(1469) <= not (a xor b);
    layer6_outputs(1470) <= a;
    layer6_outputs(1471) <= a xor b;
    layer6_outputs(1472) <= not (a or b);
    layer6_outputs(1473) <= not b;
    layer6_outputs(1474) <= not b;
    layer6_outputs(1475) <= not (a xor b);
    layer6_outputs(1476) <= a xor b;
    layer6_outputs(1477) <= not (a xor b);
    layer6_outputs(1478) <= not b;
    layer6_outputs(1479) <= b;
    layer6_outputs(1480) <= not b or a;
    layer6_outputs(1481) <= a and b;
    layer6_outputs(1482) <= a xor b;
    layer6_outputs(1483) <= not (a xor b);
    layer6_outputs(1484) <= not (a xor b);
    layer6_outputs(1485) <= b;
    layer6_outputs(1486) <= not b or a;
    layer6_outputs(1487) <= not b;
    layer6_outputs(1488) <= not b;
    layer6_outputs(1489) <= a;
    layer6_outputs(1490) <= not b;
    layer6_outputs(1491) <= b;
    layer6_outputs(1492) <= a xor b;
    layer6_outputs(1493) <= not (a xor b);
    layer6_outputs(1494) <= b;
    layer6_outputs(1495) <= b;
    layer6_outputs(1496) <= not b;
    layer6_outputs(1497) <= not (a xor b);
    layer6_outputs(1498) <= not b;
    layer6_outputs(1499) <= a and not b;
    layer6_outputs(1500) <= a;
    layer6_outputs(1501) <= '1';
    layer6_outputs(1502) <= a;
    layer6_outputs(1503) <= not (a or b);
    layer6_outputs(1504) <= a and not b;
    layer6_outputs(1505) <= b and not a;
    layer6_outputs(1506) <= not b;
    layer6_outputs(1507) <= b;
    layer6_outputs(1508) <= not a;
    layer6_outputs(1509) <= not a or b;
    layer6_outputs(1510) <= not a;
    layer6_outputs(1511) <= b;
    layer6_outputs(1512) <= '0';
    layer6_outputs(1513) <= not b;
    layer6_outputs(1514) <= not b;
    layer6_outputs(1515) <= not (a xor b);
    layer6_outputs(1516) <= a xor b;
    layer6_outputs(1517) <= b and not a;
    layer6_outputs(1518) <= not b or a;
    layer6_outputs(1519) <= b;
    layer6_outputs(1520) <= a and b;
    layer6_outputs(1521) <= a or b;
    layer6_outputs(1522) <= not a;
    layer6_outputs(1523) <= a and not b;
    layer6_outputs(1524) <= not b;
    layer6_outputs(1525) <= not (a xor b);
    layer6_outputs(1526) <= not a or b;
    layer6_outputs(1527) <= not a;
    layer6_outputs(1528) <= b and not a;
    layer6_outputs(1529) <= not (a xor b);
    layer6_outputs(1530) <= not (a or b);
    layer6_outputs(1531) <= a xor b;
    layer6_outputs(1532) <= not a;
    layer6_outputs(1533) <= not a;
    layer6_outputs(1534) <= not a;
    layer6_outputs(1535) <= a;
    layer6_outputs(1536) <= a;
    layer6_outputs(1537) <= not (a or b);
    layer6_outputs(1538) <= a xor b;
    layer6_outputs(1539) <= a xor b;
    layer6_outputs(1540) <= a;
    layer6_outputs(1541) <= a and not b;
    layer6_outputs(1542) <= a;
    layer6_outputs(1543) <= not b;
    layer6_outputs(1544) <= a xor b;
    layer6_outputs(1545) <= not a;
    layer6_outputs(1546) <= a and not b;
    layer6_outputs(1547) <= a xor b;
    layer6_outputs(1548) <= a;
    layer6_outputs(1549) <= not b;
    layer6_outputs(1550) <= not b or a;
    layer6_outputs(1551) <= a xor b;
    layer6_outputs(1552) <= a or b;
    layer6_outputs(1553) <= a xor b;
    layer6_outputs(1554) <= b;
    layer6_outputs(1555) <= not (a and b);
    layer6_outputs(1556) <= not a;
    layer6_outputs(1557) <= a;
    layer6_outputs(1558) <= a;
    layer6_outputs(1559) <= a xor b;
    layer6_outputs(1560) <= not (a xor b);
    layer6_outputs(1561) <= b;
    layer6_outputs(1562) <= not (a xor b);
    layer6_outputs(1563) <= not a;
    layer6_outputs(1564) <= not b;
    layer6_outputs(1565) <= a xor b;
    layer6_outputs(1566) <= not a;
    layer6_outputs(1567) <= b and not a;
    layer6_outputs(1568) <= b and not a;
    layer6_outputs(1569) <= a;
    layer6_outputs(1570) <= b;
    layer6_outputs(1571) <= not b;
    layer6_outputs(1572) <= not a or b;
    layer6_outputs(1573) <= not b;
    layer6_outputs(1574) <= a;
    layer6_outputs(1575) <= b and not a;
    layer6_outputs(1576) <= a and b;
    layer6_outputs(1577) <= a and b;
    layer6_outputs(1578) <= b;
    layer6_outputs(1579) <= b;
    layer6_outputs(1580) <= not (a xor b);
    layer6_outputs(1581) <= a and not b;
    layer6_outputs(1582) <= a;
    layer6_outputs(1583) <= a and b;
    layer6_outputs(1584) <= not a;
    layer6_outputs(1585) <= a;
    layer6_outputs(1586) <= a;
    layer6_outputs(1587) <= a and b;
    layer6_outputs(1588) <= a;
    layer6_outputs(1589) <= not b;
    layer6_outputs(1590) <= b;
    layer6_outputs(1591) <= not b;
    layer6_outputs(1592) <= not b;
    layer6_outputs(1593) <= b;
    layer6_outputs(1594) <= a;
    layer6_outputs(1595) <= a or b;
    layer6_outputs(1596) <= a or b;
    layer6_outputs(1597) <= a and b;
    layer6_outputs(1598) <= a or b;
    layer6_outputs(1599) <= a and not b;
    layer6_outputs(1600) <= a xor b;
    layer6_outputs(1601) <= not (a or b);
    layer6_outputs(1602) <= a;
    layer6_outputs(1603) <= b;
    layer6_outputs(1604) <= a xor b;
    layer6_outputs(1605) <= not (a xor b);
    layer6_outputs(1606) <= not b;
    layer6_outputs(1607) <= not a;
    layer6_outputs(1608) <= b;
    layer6_outputs(1609) <= not (a and b);
    layer6_outputs(1610) <= b and not a;
    layer6_outputs(1611) <= a xor b;
    layer6_outputs(1612) <= b;
    layer6_outputs(1613) <= a or b;
    layer6_outputs(1614) <= b;
    layer6_outputs(1615) <= not b;
    layer6_outputs(1616) <= not a;
    layer6_outputs(1617) <= not a or b;
    layer6_outputs(1618) <= a xor b;
    layer6_outputs(1619) <= b;
    layer6_outputs(1620) <= b and not a;
    layer6_outputs(1621) <= b;
    layer6_outputs(1622) <= not b or a;
    layer6_outputs(1623) <= b;
    layer6_outputs(1624) <= a or b;
    layer6_outputs(1625) <= not b or a;
    layer6_outputs(1626) <= a xor b;
    layer6_outputs(1627) <= not a;
    layer6_outputs(1628) <= not b or a;
    layer6_outputs(1629) <= not (a and b);
    layer6_outputs(1630) <= not b;
    layer6_outputs(1631) <= not a;
    layer6_outputs(1632) <= b;
    layer6_outputs(1633) <= a xor b;
    layer6_outputs(1634) <= a and not b;
    layer6_outputs(1635) <= not (a xor b);
    layer6_outputs(1636) <= not a;
    layer6_outputs(1637) <= b and not a;
    layer6_outputs(1638) <= not a or b;
    layer6_outputs(1639) <= a or b;
    layer6_outputs(1640) <= a;
    layer6_outputs(1641) <= not b or a;
    layer6_outputs(1642) <= a and not b;
    layer6_outputs(1643) <= a;
    layer6_outputs(1644) <= a xor b;
    layer6_outputs(1645) <= b and not a;
    layer6_outputs(1646) <= a xor b;
    layer6_outputs(1647) <= a xor b;
    layer6_outputs(1648) <= not (a xor b);
    layer6_outputs(1649) <= not b;
    layer6_outputs(1650) <= a or b;
    layer6_outputs(1651) <= not a;
    layer6_outputs(1652) <= b and not a;
    layer6_outputs(1653) <= a xor b;
    layer6_outputs(1654) <= not b;
    layer6_outputs(1655) <= not (a xor b);
    layer6_outputs(1656) <= not b or a;
    layer6_outputs(1657) <= not (a and b);
    layer6_outputs(1658) <= not b;
    layer6_outputs(1659) <= not a or b;
    layer6_outputs(1660) <= not a;
    layer6_outputs(1661) <= a;
    layer6_outputs(1662) <= not b;
    layer6_outputs(1663) <= not (a xor b);
    layer6_outputs(1664) <= not (a or b);
    layer6_outputs(1665) <= a and b;
    layer6_outputs(1666) <= not b or a;
    layer6_outputs(1667) <= b;
    layer6_outputs(1668) <= a and b;
    layer6_outputs(1669) <= not b;
    layer6_outputs(1670) <= a;
    layer6_outputs(1671) <= b;
    layer6_outputs(1672) <= not (a xor b);
    layer6_outputs(1673) <= a xor b;
    layer6_outputs(1674) <= a;
    layer6_outputs(1675) <= a xor b;
    layer6_outputs(1676) <= a;
    layer6_outputs(1677) <= not b or a;
    layer6_outputs(1678) <= not a;
    layer6_outputs(1679) <= not a;
    layer6_outputs(1680) <= not (a xor b);
    layer6_outputs(1681) <= a or b;
    layer6_outputs(1682) <= not a;
    layer6_outputs(1683) <= not (a xor b);
    layer6_outputs(1684) <= a xor b;
    layer6_outputs(1685) <= not b;
    layer6_outputs(1686) <= a;
    layer6_outputs(1687) <= not b;
    layer6_outputs(1688) <= not (a or b);
    layer6_outputs(1689) <= a;
    layer6_outputs(1690) <= not (a xor b);
    layer6_outputs(1691) <= not a or b;
    layer6_outputs(1692) <= not b;
    layer6_outputs(1693) <= a;
    layer6_outputs(1694) <= not a;
    layer6_outputs(1695) <= not b;
    layer6_outputs(1696) <= not (a and b);
    layer6_outputs(1697) <= not (a and b);
    layer6_outputs(1698) <= a and b;
    layer6_outputs(1699) <= a xor b;
    layer6_outputs(1700) <= not a;
    layer6_outputs(1701) <= a xor b;
    layer6_outputs(1702) <= a xor b;
    layer6_outputs(1703) <= not (a and b);
    layer6_outputs(1704) <= a xor b;
    layer6_outputs(1705) <= not (a xor b);
    layer6_outputs(1706) <= not b or a;
    layer6_outputs(1707) <= not (a and b);
    layer6_outputs(1708) <= a xor b;
    layer6_outputs(1709) <= not (a xor b);
    layer6_outputs(1710) <= not a;
    layer6_outputs(1711) <= a or b;
    layer6_outputs(1712) <= a;
    layer6_outputs(1713) <= a;
    layer6_outputs(1714) <= b and not a;
    layer6_outputs(1715) <= a xor b;
    layer6_outputs(1716) <= not a;
    layer6_outputs(1717) <= not b or a;
    layer6_outputs(1718) <= a xor b;
    layer6_outputs(1719) <= not a;
    layer6_outputs(1720) <= '1';
    layer6_outputs(1721) <= a;
    layer6_outputs(1722) <= a xor b;
    layer6_outputs(1723) <= b;
    layer6_outputs(1724) <= not b or a;
    layer6_outputs(1725) <= not b;
    layer6_outputs(1726) <= not b or a;
    layer6_outputs(1727) <= not b;
    layer6_outputs(1728) <= not a or b;
    layer6_outputs(1729) <= b;
    layer6_outputs(1730) <= a or b;
    layer6_outputs(1731) <= not (a xor b);
    layer6_outputs(1732) <= not a;
    layer6_outputs(1733) <= a;
    layer6_outputs(1734) <= not a;
    layer6_outputs(1735) <= a or b;
    layer6_outputs(1736) <= not (a or b);
    layer6_outputs(1737) <= not a;
    layer6_outputs(1738) <= a;
    layer6_outputs(1739) <= not b;
    layer6_outputs(1740) <= a xor b;
    layer6_outputs(1741) <= a;
    layer6_outputs(1742) <= not b;
    layer6_outputs(1743) <= a and not b;
    layer6_outputs(1744) <= a;
    layer6_outputs(1745) <= b and not a;
    layer6_outputs(1746) <= not (a or b);
    layer6_outputs(1747) <= a xor b;
    layer6_outputs(1748) <= b and not a;
    layer6_outputs(1749) <= a xor b;
    layer6_outputs(1750) <= b;
    layer6_outputs(1751) <= b;
    layer6_outputs(1752) <= not a;
    layer6_outputs(1753) <= b and not a;
    layer6_outputs(1754) <= a xor b;
    layer6_outputs(1755) <= not b;
    layer6_outputs(1756) <= b;
    layer6_outputs(1757) <= a;
    layer6_outputs(1758) <= a and not b;
    layer6_outputs(1759) <= not a;
    layer6_outputs(1760) <= a;
    layer6_outputs(1761) <= not a;
    layer6_outputs(1762) <= a xor b;
    layer6_outputs(1763) <= a or b;
    layer6_outputs(1764) <= not a or b;
    layer6_outputs(1765) <= not b;
    layer6_outputs(1766) <= b;
    layer6_outputs(1767) <= a;
    layer6_outputs(1768) <= not b;
    layer6_outputs(1769) <= not (a and b);
    layer6_outputs(1770) <= not (a xor b);
    layer6_outputs(1771) <= not b;
    layer6_outputs(1772) <= a and b;
    layer6_outputs(1773) <= a;
    layer6_outputs(1774) <= not a;
    layer6_outputs(1775) <= not (a or b);
    layer6_outputs(1776) <= b;
    layer6_outputs(1777) <= a xor b;
    layer6_outputs(1778) <= b;
    layer6_outputs(1779) <= b;
    layer6_outputs(1780) <= not a;
    layer6_outputs(1781) <= not a;
    layer6_outputs(1782) <= b;
    layer6_outputs(1783) <= not a or b;
    layer6_outputs(1784) <= not b;
    layer6_outputs(1785) <= a;
    layer6_outputs(1786) <= b;
    layer6_outputs(1787) <= not (a xor b);
    layer6_outputs(1788) <= b;
    layer6_outputs(1789) <= a and not b;
    layer6_outputs(1790) <= not b or a;
    layer6_outputs(1791) <= a xor b;
    layer6_outputs(1792) <= a and b;
    layer6_outputs(1793) <= a;
    layer6_outputs(1794) <= a;
    layer6_outputs(1795) <= not a or b;
    layer6_outputs(1796) <= a and b;
    layer6_outputs(1797) <= a and not b;
    layer6_outputs(1798) <= a or b;
    layer6_outputs(1799) <= not b;
    layer6_outputs(1800) <= a;
    layer6_outputs(1801) <= not (a xor b);
    layer6_outputs(1802) <= not b;
    layer6_outputs(1803) <= not (a and b);
    layer6_outputs(1804) <= not a;
    layer6_outputs(1805) <= a xor b;
    layer6_outputs(1806) <= not b;
    layer6_outputs(1807) <= not a;
    layer6_outputs(1808) <= not (a or b);
    layer6_outputs(1809) <= b and not a;
    layer6_outputs(1810) <= not b;
    layer6_outputs(1811) <= not b;
    layer6_outputs(1812) <= not b;
    layer6_outputs(1813) <= not (a or b);
    layer6_outputs(1814) <= b;
    layer6_outputs(1815) <= not a;
    layer6_outputs(1816) <= b;
    layer6_outputs(1817) <= not a;
    layer6_outputs(1818) <= a;
    layer6_outputs(1819) <= a and b;
    layer6_outputs(1820) <= not a or b;
    layer6_outputs(1821) <= not b or a;
    layer6_outputs(1822) <= a or b;
    layer6_outputs(1823) <= not (a or b);
    layer6_outputs(1824) <= not b;
    layer6_outputs(1825) <= not a;
    layer6_outputs(1826) <= not (a and b);
    layer6_outputs(1827) <= not b;
    layer6_outputs(1828) <= b;
    layer6_outputs(1829) <= a and not b;
    layer6_outputs(1830) <= not b;
    layer6_outputs(1831) <= a;
    layer6_outputs(1832) <= not b;
    layer6_outputs(1833) <= b and not a;
    layer6_outputs(1834) <= a and b;
    layer6_outputs(1835) <= not (a and b);
    layer6_outputs(1836) <= a;
    layer6_outputs(1837) <= not a or b;
    layer6_outputs(1838) <= a xor b;
    layer6_outputs(1839) <= b;
    layer6_outputs(1840) <= not b or a;
    layer6_outputs(1841) <= not a;
    layer6_outputs(1842) <= a and b;
    layer6_outputs(1843) <= b;
    layer6_outputs(1844) <= b;
    layer6_outputs(1845) <= a xor b;
    layer6_outputs(1846) <= b;
    layer6_outputs(1847) <= not a or b;
    layer6_outputs(1848) <= a xor b;
    layer6_outputs(1849) <= not b or a;
    layer6_outputs(1850) <= a xor b;
    layer6_outputs(1851) <= not b or a;
    layer6_outputs(1852) <= a;
    layer6_outputs(1853) <= a;
    layer6_outputs(1854) <= not b or a;
    layer6_outputs(1855) <= not (a or b);
    layer6_outputs(1856) <= a;
    layer6_outputs(1857) <= not a;
    layer6_outputs(1858) <= not a;
    layer6_outputs(1859) <= a and b;
    layer6_outputs(1860) <= not b or a;
    layer6_outputs(1861) <= b and not a;
    layer6_outputs(1862) <= b and not a;
    layer6_outputs(1863) <= a and b;
    layer6_outputs(1864) <= a or b;
    layer6_outputs(1865) <= b;
    layer6_outputs(1866) <= not (a and b);
    layer6_outputs(1867) <= not b;
    layer6_outputs(1868) <= not (a and b);
    layer6_outputs(1869) <= b;
    layer6_outputs(1870) <= not (a and b);
    layer6_outputs(1871) <= not b;
    layer6_outputs(1872) <= a;
    layer6_outputs(1873) <= not b or a;
    layer6_outputs(1874) <= not b or a;
    layer6_outputs(1875) <= a;
    layer6_outputs(1876) <= not (a xor b);
    layer6_outputs(1877) <= '0';
    layer6_outputs(1878) <= a and not b;
    layer6_outputs(1879) <= b and not a;
    layer6_outputs(1880) <= a or b;
    layer6_outputs(1881) <= b and not a;
    layer6_outputs(1882) <= a or b;
    layer6_outputs(1883) <= not (a xor b);
    layer6_outputs(1884) <= not b;
    layer6_outputs(1885) <= not (a and b);
    layer6_outputs(1886) <= not b;
    layer6_outputs(1887) <= not a;
    layer6_outputs(1888) <= not a or b;
    layer6_outputs(1889) <= b;
    layer6_outputs(1890) <= a and not b;
    layer6_outputs(1891) <= a and b;
    layer6_outputs(1892) <= not a;
    layer6_outputs(1893) <= not a;
    layer6_outputs(1894) <= a;
    layer6_outputs(1895) <= not a;
    layer6_outputs(1896) <= a;
    layer6_outputs(1897) <= a;
    layer6_outputs(1898) <= not (a xor b);
    layer6_outputs(1899) <= b;
    layer6_outputs(1900) <= not a;
    layer6_outputs(1901) <= not a;
    layer6_outputs(1902) <= not a;
    layer6_outputs(1903) <= a and not b;
    layer6_outputs(1904) <= not a;
    layer6_outputs(1905) <= not b;
    layer6_outputs(1906) <= not b;
    layer6_outputs(1907) <= a;
    layer6_outputs(1908) <= a;
    layer6_outputs(1909) <= a;
    layer6_outputs(1910) <= not (a xor b);
    layer6_outputs(1911) <= not a;
    layer6_outputs(1912) <= not b;
    layer6_outputs(1913) <= not (a xor b);
    layer6_outputs(1914) <= a xor b;
    layer6_outputs(1915) <= a;
    layer6_outputs(1916) <= not a;
    layer6_outputs(1917) <= '1';
    layer6_outputs(1918) <= not b;
    layer6_outputs(1919) <= not a;
    layer6_outputs(1920) <= not b;
    layer6_outputs(1921) <= not b;
    layer6_outputs(1922) <= not (a and b);
    layer6_outputs(1923) <= not a;
    layer6_outputs(1924) <= not a or b;
    layer6_outputs(1925) <= a;
    layer6_outputs(1926) <= b;
    layer6_outputs(1927) <= not (a or b);
    layer6_outputs(1928) <= b;
    layer6_outputs(1929) <= b and not a;
    layer6_outputs(1930) <= a and b;
    layer6_outputs(1931) <= a;
    layer6_outputs(1932) <= not (a xor b);
    layer6_outputs(1933) <= not b or a;
    layer6_outputs(1934) <= not (a or b);
    layer6_outputs(1935) <= not (a and b);
    layer6_outputs(1936) <= not b;
    layer6_outputs(1937) <= '0';
    layer6_outputs(1938) <= not (a and b);
    layer6_outputs(1939) <= a and b;
    layer6_outputs(1940) <= not a;
    layer6_outputs(1941) <= not b;
    layer6_outputs(1942) <= not b or a;
    layer6_outputs(1943) <= a;
    layer6_outputs(1944) <= a and not b;
    layer6_outputs(1945) <= a;
    layer6_outputs(1946) <= a xor b;
    layer6_outputs(1947) <= not (a or b);
    layer6_outputs(1948) <= not (a xor b);
    layer6_outputs(1949) <= not b;
    layer6_outputs(1950) <= not b or a;
    layer6_outputs(1951) <= not (a xor b);
    layer6_outputs(1952) <= a;
    layer6_outputs(1953) <= b;
    layer6_outputs(1954) <= not (a xor b);
    layer6_outputs(1955) <= a xor b;
    layer6_outputs(1956) <= not (a xor b);
    layer6_outputs(1957) <= not (a xor b);
    layer6_outputs(1958) <= a xor b;
    layer6_outputs(1959) <= a;
    layer6_outputs(1960) <= not b or a;
    layer6_outputs(1961) <= a and b;
    layer6_outputs(1962) <= not a;
    layer6_outputs(1963) <= not b;
    layer6_outputs(1964) <= a or b;
    layer6_outputs(1965) <= not b;
    layer6_outputs(1966) <= not b;
    layer6_outputs(1967) <= b;
    layer6_outputs(1968) <= b;
    layer6_outputs(1969) <= a xor b;
    layer6_outputs(1970) <= a;
    layer6_outputs(1971) <= not a;
    layer6_outputs(1972) <= a and b;
    layer6_outputs(1973) <= a xor b;
    layer6_outputs(1974) <= not a;
    layer6_outputs(1975) <= a xor b;
    layer6_outputs(1976) <= not a;
    layer6_outputs(1977) <= not b or a;
    layer6_outputs(1978) <= not a;
    layer6_outputs(1979) <= b;
    layer6_outputs(1980) <= b;
    layer6_outputs(1981) <= not a or b;
    layer6_outputs(1982) <= a and b;
    layer6_outputs(1983) <= not a;
    layer6_outputs(1984) <= not (a xor b);
    layer6_outputs(1985) <= not b;
    layer6_outputs(1986) <= a and b;
    layer6_outputs(1987) <= not a or b;
    layer6_outputs(1988) <= a or b;
    layer6_outputs(1989) <= a xor b;
    layer6_outputs(1990) <= a xor b;
    layer6_outputs(1991) <= b;
    layer6_outputs(1992) <= b;
    layer6_outputs(1993) <= not (a or b);
    layer6_outputs(1994) <= b and not a;
    layer6_outputs(1995) <= not a;
    layer6_outputs(1996) <= a xor b;
    layer6_outputs(1997) <= not (a or b);
    layer6_outputs(1998) <= not (a and b);
    layer6_outputs(1999) <= not a;
    layer6_outputs(2000) <= b;
    layer6_outputs(2001) <= not b;
    layer6_outputs(2002) <= b;
    layer6_outputs(2003) <= not b;
    layer6_outputs(2004) <= not (a and b);
    layer6_outputs(2005) <= not (a or b);
    layer6_outputs(2006) <= not (a or b);
    layer6_outputs(2007) <= not a;
    layer6_outputs(2008) <= a;
    layer6_outputs(2009) <= not a or b;
    layer6_outputs(2010) <= not a;
    layer6_outputs(2011) <= a;
    layer6_outputs(2012) <= not b;
    layer6_outputs(2013) <= not (a and b);
    layer6_outputs(2014) <= b;
    layer6_outputs(2015) <= not (a xor b);
    layer6_outputs(2016) <= b;
    layer6_outputs(2017) <= not b;
    layer6_outputs(2018) <= not b;
    layer6_outputs(2019) <= a;
    layer6_outputs(2020) <= not a;
    layer6_outputs(2021) <= a xor b;
    layer6_outputs(2022) <= not b;
    layer6_outputs(2023) <= not a or b;
    layer6_outputs(2024) <= not (a xor b);
    layer6_outputs(2025) <= not a;
    layer6_outputs(2026) <= not b or a;
    layer6_outputs(2027) <= b;
    layer6_outputs(2028) <= not a or b;
    layer6_outputs(2029) <= not a or b;
    layer6_outputs(2030) <= a xor b;
    layer6_outputs(2031) <= not b;
    layer6_outputs(2032) <= not a;
    layer6_outputs(2033) <= not a;
    layer6_outputs(2034) <= not b or a;
    layer6_outputs(2035) <= not (a xor b);
    layer6_outputs(2036) <= b and not a;
    layer6_outputs(2037) <= a xor b;
    layer6_outputs(2038) <= not (a xor b);
    layer6_outputs(2039) <= not b;
    layer6_outputs(2040) <= a xor b;
    layer6_outputs(2041) <= not (a xor b);
    layer6_outputs(2042) <= not (a xor b);
    layer6_outputs(2043) <= not b;
    layer6_outputs(2044) <= not a or b;
    layer6_outputs(2045) <= a xor b;
    layer6_outputs(2046) <= a;
    layer6_outputs(2047) <= not (a xor b);
    layer6_outputs(2048) <= not (a xor b);
    layer6_outputs(2049) <= not a;
    layer6_outputs(2050) <= a xor b;
    layer6_outputs(2051) <= b;
    layer6_outputs(2052) <= '1';
    layer6_outputs(2053) <= not a or b;
    layer6_outputs(2054) <= a;
    layer6_outputs(2055) <= not b or a;
    layer6_outputs(2056) <= a or b;
    layer6_outputs(2057) <= b;
    layer6_outputs(2058) <= b;
    layer6_outputs(2059) <= b;
    layer6_outputs(2060) <= a;
    layer6_outputs(2061) <= not b;
    layer6_outputs(2062) <= b;
    layer6_outputs(2063) <= a or b;
    layer6_outputs(2064) <= a xor b;
    layer6_outputs(2065) <= not b;
    layer6_outputs(2066) <= not a;
    layer6_outputs(2067) <= not b;
    layer6_outputs(2068) <= b and not a;
    layer6_outputs(2069) <= a;
    layer6_outputs(2070) <= not a;
    layer6_outputs(2071) <= not a or b;
    layer6_outputs(2072) <= b;
    layer6_outputs(2073) <= a and b;
    layer6_outputs(2074) <= not a;
    layer6_outputs(2075) <= not (a or b);
    layer6_outputs(2076) <= not b;
    layer6_outputs(2077) <= a xor b;
    layer6_outputs(2078) <= not a;
    layer6_outputs(2079) <= not a;
    layer6_outputs(2080) <= not (a xor b);
    layer6_outputs(2081) <= not (a xor b);
    layer6_outputs(2082) <= not (a xor b);
    layer6_outputs(2083) <= not b;
    layer6_outputs(2084) <= not b or a;
    layer6_outputs(2085) <= not (a xor b);
    layer6_outputs(2086) <= not b;
    layer6_outputs(2087) <= not a;
    layer6_outputs(2088) <= not a;
    layer6_outputs(2089) <= not (a xor b);
    layer6_outputs(2090) <= not b;
    layer6_outputs(2091) <= not b;
    layer6_outputs(2092) <= a or b;
    layer6_outputs(2093) <= a and b;
    layer6_outputs(2094) <= a and b;
    layer6_outputs(2095) <= not b or a;
    layer6_outputs(2096) <= not (a xor b);
    layer6_outputs(2097) <= not b;
    layer6_outputs(2098) <= not a;
    layer6_outputs(2099) <= a;
    layer6_outputs(2100) <= a xor b;
    layer6_outputs(2101) <= b;
    layer6_outputs(2102) <= a and not b;
    layer6_outputs(2103) <= a;
    layer6_outputs(2104) <= b and not a;
    layer6_outputs(2105) <= not a;
    layer6_outputs(2106) <= b and not a;
    layer6_outputs(2107) <= not a or b;
    layer6_outputs(2108) <= a;
    layer6_outputs(2109) <= b;
    layer6_outputs(2110) <= a or b;
    layer6_outputs(2111) <= a xor b;
    layer6_outputs(2112) <= not (a and b);
    layer6_outputs(2113) <= a xor b;
    layer6_outputs(2114) <= not b;
    layer6_outputs(2115) <= not a or b;
    layer6_outputs(2116) <= not a;
    layer6_outputs(2117) <= not (a xor b);
    layer6_outputs(2118) <= not (a and b);
    layer6_outputs(2119) <= a xor b;
    layer6_outputs(2120) <= not a;
    layer6_outputs(2121) <= b;
    layer6_outputs(2122) <= not (a or b);
    layer6_outputs(2123) <= not a;
    layer6_outputs(2124) <= not a;
    layer6_outputs(2125) <= a or b;
    layer6_outputs(2126) <= not (a xor b);
    layer6_outputs(2127) <= not a;
    layer6_outputs(2128) <= b and not a;
    layer6_outputs(2129) <= not a;
    layer6_outputs(2130) <= not (a or b);
    layer6_outputs(2131) <= a;
    layer6_outputs(2132) <= a xor b;
    layer6_outputs(2133) <= not a;
    layer6_outputs(2134) <= not (a xor b);
    layer6_outputs(2135) <= not b;
    layer6_outputs(2136) <= not b;
    layer6_outputs(2137) <= not (a and b);
    layer6_outputs(2138) <= b;
    layer6_outputs(2139) <= not b;
    layer6_outputs(2140) <= a;
    layer6_outputs(2141) <= a;
    layer6_outputs(2142) <= a xor b;
    layer6_outputs(2143) <= a;
    layer6_outputs(2144) <= b;
    layer6_outputs(2145) <= b;
    layer6_outputs(2146) <= not b;
    layer6_outputs(2147) <= not (a xor b);
    layer6_outputs(2148) <= not a;
    layer6_outputs(2149) <= a xor b;
    layer6_outputs(2150) <= not b;
    layer6_outputs(2151) <= not b;
    layer6_outputs(2152) <= not (a xor b);
    layer6_outputs(2153) <= not a;
    layer6_outputs(2154) <= not b;
    layer6_outputs(2155) <= a xor b;
    layer6_outputs(2156) <= not b;
    layer6_outputs(2157) <= b and not a;
    layer6_outputs(2158) <= not (a xor b);
    layer6_outputs(2159) <= a or b;
    layer6_outputs(2160) <= not (a xor b);
    layer6_outputs(2161) <= not b;
    layer6_outputs(2162) <= not (a xor b);
    layer6_outputs(2163) <= b and not a;
    layer6_outputs(2164) <= not b or a;
    layer6_outputs(2165) <= a and b;
    layer6_outputs(2166) <= a or b;
    layer6_outputs(2167) <= not a;
    layer6_outputs(2168) <= a xor b;
    layer6_outputs(2169) <= a xor b;
    layer6_outputs(2170) <= not a;
    layer6_outputs(2171) <= not a;
    layer6_outputs(2172) <= a xor b;
    layer6_outputs(2173) <= b and not a;
    layer6_outputs(2174) <= a;
    layer6_outputs(2175) <= b and not a;
    layer6_outputs(2176) <= not a or b;
    layer6_outputs(2177) <= a and not b;
    layer6_outputs(2178) <= not b or a;
    layer6_outputs(2179) <= a and b;
    layer6_outputs(2180) <= a or b;
    layer6_outputs(2181) <= not b;
    layer6_outputs(2182) <= a;
    layer6_outputs(2183) <= not a or b;
    layer6_outputs(2184) <= a xor b;
    layer6_outputs(2185) <= not b;
    layer6_outputs(2186) <= not (a xor b);
    layer6_outputs(2187) <= not b;
    layer6_outputs(2188) <= not a or b;
    layer6_outputs(2189) <= not (a xor b);
    layer6_outputs(2190) <= not (a xor b);
    layer6_outputs(2191) <= a and not b;
    layer6_outputs(2192) <= a;
    layer6_outputs(2193) <= not a or b;
    layer6_outputs(2194) <= a or b;
    layer6_outputs(2195) <= a;
    layer6_outputs(2196) <= b;
    layer6_outputs(2197) <= a xor b;
    layer6_outputs(2198) <= not (a or b);
    layer6_outputs(2199) <= not a;
    layer6_outputs(2200) <= not b;
    layer6_outputs(2201) <= a or b;
    layer6_outputs(2202) <= a and b;
    layer6_outputs(2203) <= a;
    layer6_outputs(2204) <= not a or b;
    layer6_outputs(2205) <= a and b;
    layer6_outputs(2206) <= b and not a;
    layer6_outputs(2207) <= a;
    layer6_outputs(2208) <= a and b;
    layer6_outputs(2209) <= not (a xor b);
    layer6_outputs(2210) <= not (a or b);
    layer6_outputs(2211) <= not (a xor b);
    layer6_outputs(2212) <= not a or b;
    layer6_outputs(2213) <= a;
    layer6_outputs(2214) <= '1';
    layer6_outputs(2215) <= not a;
    layer6_outputs(2216) <= a xor b;
    layer6_outputs(2217) <= not b;
    layer6_outputs(2218) <= a;
    layer6_outputs(2219) <= not (a xor b);
    layer6_outputs(2220) <= not b or a;
    layer6_outputs(2221) <= a and not b;
    layer6_outputs(2222) <= a and not b;
    layer6_outputs(2223) <= a xor b;
    layer6_outputs(2224) <= a and b;
    layer6_outputs(2225) <= not (a xor b);
    layer6_outputs(2226) <= not b;
    layer6_outputs(2227) <= not a;
    layer6_outputs(2228) <= a;
    layer6_outputs(2229) <= a or b;
    layer6_outputs(2230) <= b;
    layer6_outputs(2231) <= not a;
    layer6_outputs(2232) <= not b;
    layer6_outputs(2233) <= a xor b;
    layer6_outputs(2234) <= a xor b;
    layer6_outputs(2235) <= a or b;
    layer6_outputs(2236) <= a and not b;
    layer6_outputs(2237) <= not b;
    layer6_outputs(2238) <= not a;
    layer6_outputs(2239) <= a and not b;
    layer6_outputs(2240) <= not b;
    layer6_outputs(2241) <= a and not b;
    layer6_outputs(2242) <= not a;
    layer6_outputs(2243) <= a and b;
    layer6_outputs(2244) <= not (a and b);
    layer6_outputs(2245) <= not (a and b);
    layer6_outputs(2246) <= not (a xor b);
    layer6_outputs(2247) <= b;
    layer6_outputs(2248) <= a and not b;
    layer6_outputs(2249) <= not (a xor b);
    layer6_outputs(2250) <= b and not a;
    layer6_outputs(2251) <= '1';
    layer6_outputs(2252) <= not a or b;
    layer6_outputs(2253) <= a xor b;
    layer6_outputs(2254) <= not b;
    layer6_outputs(2255) <= not (a and b);
    layer6_outputs(2256) <= not (a and b);
    layer6_outputs(2257) <= a or b;
    layer6_outputs(2258) <= a and b;
    layer6_outputs(2259) <= not b or a;
    layer6_outputs(2260) <= a and not b;
    layer6_outputs(2261) <= not a or b;
    layer6_outputs(2262) <= a;
    layer6_outputs(2263) <= not b;
    layer6_outputs(2264) <= not (a and b);
    layer6_outputs(2265) <= not b or a;
    layer6_outputs(2266) <= not (a xor b);
    layer6_outputs(2267) <= '0';
    layer6_outputs(2268) <= not (a xor b);
    layer6_outputs(2269) <= a;
    layer6_outputs(2270) <= not a;
    layer6_outputs(2271) <= a or b;
    layer6_outputs(2272) <= a;
    layer6_outputs(2273) <= b;
    layer6_outputs(2274) <= not (a or b);
    layer6_outputs(2275) <= not b or a;
    layer6_outputs(2276) <= a xor b;
    layer6_outputs(2277) <= a;
    layer6_outputs(2278) <= a;
    layer6_outputs(2279) <= a or b;
    layer6_outputs(2280) <= a and b;
    layer6_outputs(2281) <= b;
    layer6_outputs(2282) <= a or b;
    layer6_outputs(2283) <= a and not b;
    layer6_outputs(2284) <= b and not a;
    layer6_outputs(2285) <= not b;
    layer6_outputs(2286) <= not a;
    layer6_outputs(2287) <= b;
    layer6_outputs(2288) <= not (a xor b);
    layer6_outputs(2289) <= not (a and b);
    layer6_outputs(2290) <= not (a xor b);
    layer6_outputs(2291) <= not (a or b);
    layer6_outputs(2292) <= not (a xor b);
    layer6_outputs(2293) <= b;
    layer6_outputs(2294) <= not a or b;
    layer6_outputs(2295) <= a and b;
    layer6_outputs(2296) <= a;
    layer6_outputs(2297) <= a and not b;
    layer6_outputs(2298) <= a xor b;
    layer6_outputs(2299) <= not b;
    layer6_outputs(2300) <= not (a xor b);
    layer6_outputs(2301) <= a and b;
    layer6_outputs(2302) <= not b or a;
    layer6_outputs(2303) <= not b;
    layer6_outputs(2304) <= not b;
    layer6_outputs(2305) <= a xor b;
    layer6_outputs(2306) <= not (a and b);
    layer6_outputs(2307) <= not (a or b);
    layer6_outputs(2308) <= not b;
    layer6_outputs(2309) <= b;
    layer6_outputs(2310) <= not b;
    layer6_outputs(2311) <= not a;
    layer6_outputs(2312) <= not (a xor b);
    layer6_outputs(2313) <= b;
    layer6_outputs(2314) <= a or b;
    layer6_outputs(2315) <= not a;
    layer6_outputs(2316) <= a or b;
    layer6_outputs(2317) <= a;
    layer6_outputs(2318) <= not a;
    layer6_outputs(2319) <= b;
    layer6_outputs(2320) <= not a or b;
    layer6_outputs(2321) <= b;
    layer6_outputs(2322) <= a;
    layer6_outputs(2323) <= a;
    layer6_outputs(2324) <= not b;
    layer6_outputs(2325) <= a xor b;
    layer6_outputs(2326) <= not b;
    layer6_outputs(2327) <= a and not b;
    layer6_outputs(2328) <= not (a or b);
    layer6_outputs(2329) <= not a or b;
    layer6_outputs(2330) <= a and b;
    layer6_outputs(2331) <= not b;
    layer6_outputs(2332) <= not a or b;
    layer6_outputs(2333) <= a or b;
    layer6_outputs(2334) <= not b;
    layer6_outputs(2335) <= a xor b;
    layer6_outputs(2336) <= a xor b;
    layer6_outputs(2337) <= b;
    layer6_outputs(2338) <= b;
    layer6_outputs(2339) <= a xor b;
    layer6_outputs(2340) <= a;
    layer6_outputs(2341) <= not b;
    layer6_outputs(2342) <= a and b;
    layer6_outputs(2343) <= a xor b;
    layer6_outputs(2344) <= not b or a;
    layer6_outputs(2345) <= not (a xor b);
    layer6_outputs(2346) <= b;
    layer6_outputs(2347) <= not (a and b);
    layer6_outputs(2348) <= '1';
    layer6_outputs(2349) <= a;
    layer6_outputs(2350) <= not (a and b);
    layer6_outputs(2351) <= not a;
    layer6_outputs(2352) <= not a;
    layer6_outputs(2353) <= a;
    layer6_outputs(2354) <= not b or a;
    layer6_outputs(2355) <= not a;
    layer6_outputs(2356) <= not (a xor b);
    layer6_outputs(2357) <= not (a or b);
    layer6_outputs(2358) <= not a;
    layer6_outputs(2359) <= a;
    layer6_outputs(2360) <= a and b;
    layer6_outputs(2361) <= b;
    layer6_outputs(2362) <= b;
    layer6_outputs(2363) <= a or b;
    layer6_outputs(2364) <= not (a xor b);
    layer6_outputs(2365) <= a xor b;
    layer6_outputs(2366) <= not a;
    layer6_outputs(2367) <= not a;
    layer6_outputs(2368) <= a xor b;
    layer6_outputs(2369) <= b;
    layer6_outputs(2370) <= b;
    layer6_outputs(2371) <= a xor b;
    layer6_outputs(2372) <= b;
    layer6_outputs(2373) <= b;
    layer6_outputs(2374) <= not (a xor b);
    layer6_outputs(2375) <= not a;
    layer6_outputs(2376) <= not (a xor b);
    layer6_outputs(2377) <= a and not b;
    layer6_outputs(2378) <= a xor b;
    layer6_outputs(2379) <= not (a xor b);
    layer6_outputs(2380) <= a;
    layer6_outputs(2381) <= not (a and b);
    layer6_outputs(2382) <= not b;
    layer6_outputs(2383) <= a and b;
    layer6_outputs(2384) <= a and not b;
    layer6_outputs(2385) <= a and not b;
    layer6_outputs(2386) <= b;
    layer6_outputs(2387) <= not a or b;
    layer6_outputs(2388) <= a;
    layer6_outputs(2389) <= a and b;
    layer6_outputs(2390) <= a;
    layer6_outputs(2391) <= b;
    layer6_outputs(2392) <= not a;
    layer6_outputs(2393) <= not a;
    layer6_outputs(2394) <= a or b;
    layer6_outputs(2395) <= not (a and b);
    layer6_outputs(2396) <= not (a xor b);
    layer6_outputs(2397) <= not b;
    layer6_outputs(2398) <= not b;
    layer6_outputs(2399) <= a or b;
    layer6_outputs(2400) <= a;
    layer6_outputs(2401) <= b;
    layer6_outputs(2402) <= a;
    layer6_outputs(2403) <= b and not a;
    layer6_outputs(2404) <= not (a xor b);
    layer6_outputs(2405) <= a or b;
    layer6_outputs(2406) <= not a;
    layer6_outputs(2407) <= a xor b;
    layer6_outputs(2408) <= not b;
    layer6_outputs(2409) <= not a;
    layer6_outputs(2410) <= a xor b;
    layer6_outputs(2411) <= a xor b;
    layer6_outputs(2412) <= a;
    layer6_outputs(2413) <= not a or b;
    layer6_outputs(2414) <= b;
    layer6_outputs(2415) <= a xor b;
    layer6_outputs(2416) <= a and b;
    layer6_outputs(2417) <= not (a xor b);
    layer6_outputs(2418) <= not b;
    layer6_outputs(2419) <= not (a or b);
    layer6_outputs(2420) <= a and b;
    layer6_outputs(2421) <= a;
    layer6_outputs(2422) <= b;
    layer6_outputs(2423) <= not a or b;
    layer6_outputs(2424) <= not b;
    layer6_outputs(2425) <= a xor b;
    layer6_outputs(2426) <= not a;
    layer6_outputs(2427) <= not a;
    layer6_outputs(2428) <= b;
    layer6_outputs(2429) <= not (a xor b);
    layer6_outputs(2430) <= b;
    layer6_outputs(2431) <= not a;
    layer6_outputs(2432) <= not a;
    layer6_outputs(2433) <= a xor b;
    layer6_outputs(2434) <= a and b;
    layer6_outputs(2435) <= b;
    layer6_outputs(2436) <= a;
    layer6_outputs(2437) <= a xor b;
    layer6_outputs(2438) <= not a;
    layer6_outputs(2439) <= not (a xor b);
    layer6_outputs(2440) <= a;
    layer6_outputs(2441) <= b;
    layer6_outputs(2442) <= a or b;
    layer6_outputs(2443) <= a;
    layer6_outputs(2444) <= not a;
    layer6_outputs(2445) <= a xor b;
    layer6_outputs(2446) <= not (a and b);
    layer6_outputs(2447) <= b and not a;
    layer6_outputs(2448) <= a and not b;
    layer6_outputs(2449) <= not (a xor b);
    layer6_outputs(2450) <= not (a xor b);
    layer6_outputs(2451) <= not (a or b);
    layer6_outputs(2452) <= b;
    layer6_outputs(2453) <= not (a xor b);
    layer6_outputs(2454) <= b;
    layer6_outputs(2455) <= b;
    layer6_outputs(2456) <= a or b;
    layer6_outputs(2457) <= not a or b;
    layer6_outputs(2458) <= a xor b;
    layer6_outputs(2459) <= not (a xor b);
    layer6_outputs(2460) <= not a;
    layer6_outputs(2461) <= not b;
    layer6_outputs(2462) <= b and not a;
    layer6_outputs(2463) <= not b;
    layer6_outputs(2464) <= a and b;
    layer6_outputs(2465) <= a and not b;
    layer6_outputs(2466) <= not a;
    layer6_outputs(2467) <= b;
    layer6_outputs(2468) <= b;
    layer6_outputs(2469) <= a xor b;
    layer6_outputs(2470) <= a;
    layer6_outputs(2471) <= a;
    layer6_outputs(2472) <= a xor b;
    layer6_outputs(2473) <= not (a xor b);
    layer6_outputs(2474) <= not (a or b);
    layer6_outputs(2475) <= a xor b;
    layer6_outputs(2476) <= a or b;
    layer6_outputs(2477) <= not b;
    layer6_outputs(2478) <= a;
    layer6_outputs(2479) <= a or b;
    layer6_outputs(2480) <= b;
    layer6_outputs(2481) <= not (a xor b);
    layer6_outputs(2482) <= not a;
    layer6_outputs(2483) <= a;
    layer6_outputs(2484) <= not b;
    layer6_outputs(2485) <= b;
    layer6_outputs(2486) <= a xor b;
    layer6_outputs(2487) <= not (a xor b);
    layer6_outputs(2488) <= a and not b;
    layer6_outputs(2489) <= a xor b;
    layer6_outputs(2490) <= a and b;
    layer6_outputs(2491) <= not (a xor b);
    layer6_outputs(2492) <= not (a xor b);
    layer6_outputs(2493) <= not (a xor b);
    layer6_outputs(2494) <= a and b;
    layer6_outputs(2495) <= not a;
    layer6_outputs(2496) <= b and not a;
    layer6_outputs(2497) <= a and b;
    layer6_outputs(2498) <= a xor b;
    layer6_outputs(2499) <= not a or b;
    layer6_outputs(2500) <= not a;
    layer6_outputs(2501) <= not a;
    layer6_outputs(2502) <= a;
    layer6_outputs(2503) <= not a;
    layer6_outputs(2504) <= not (a xor b);
    layer6_outputs(2505) <= a xor b;
    layer6_outputs(2506) <= not (a xor b);
    layer6_outputs(2507) <= not (a and b);
    layer6_outputs(2508) <= not a or b;
    layer6_outputs(2509) <= not b or a;
    layer6_outputs(2510) <= a;
    layer6_outputs(2511) <= not (a and b);
    layer6_outputs(2512) <= a or b;
    layer6_outputs(2513) <= a and not b;
    layer6_outputs(2514) <= a xor b;
    layer6_outputs(2515) <= not (a xor b);
    layer6_outputs(2516) <= b and not a;
    layer6_outputs(2517) <= not (a xor b);
    layer6_outputs(2518) <= a xor b;
    layer6_outputs(2519) <= not a;
    layer6_outputs(2520) <= a xor b;
    layer6_outputs(2521) <= a xor b;
    layer6_outputs(2522) <= not (a xor b);
    layer6_outputs(2523) <= a or b;
    layer6_outputs(2524) <= a xor b;
    layer6_outputs(2525) <= a and not b;
    layer6_outputs(2526) <= b;
    layer6_outputs(2527) <= not (a and b);
    layer6_outputs(2528) <= not (a xor b);
    layer6_outputs(2529) <= a;
    layer6_outputs(2530) <= a;
    layer6_outputs(2531) <= not b or a;
    layer6_outputs(2532) <= not (a xor b);
    layer6_outputs(2533) <= a xor b;
    layer6_outputs(2534) <= not (a xor b);
    layer6_outputs(2535) <= a xor b;
    layer6_outputs(2536) <= not b or a;
    layer6_outputs(2537) <= not (a or b);
    layer6_outputs(2538) <= a;
    layer6_outputs(2539) <= not a or b;
    layer6_outputs(2540) <= not b or a;
    layer6_outputs(2541) <= a;
    layer6_outputs(2542) <= a;
    layer6_outputs(2543) <= a or b;
    layer6_outputs(2544) <= a;
    layer6_outputs(2545) <= a;
    layer6_outputs(2546) <= b;
    layer6_outputs(2547) <= b;
    layer6_outputs(2548) <= not (a and b);
    layer6_outputs(2549) <= a or b;
    layer6_outputs(2550) <= not (a and b);
    layer6_outputs(2551) <= a and not b;
    layer6_outputs(2552) <= a;
    layer6_outputs(2553) <= a xor b;
    layer6_outputs(2554) <= '0';
    layer6_outputs(2555) <= not b;
    layer6_outputs(2556) <= not a;
    layer6_outputs(2557) <= not (a xor b);
    layer6_outputs(2558) <= not (a and b);
    layer6_outputs(2559) <= a xor b;
    layer6_outputs(2560) <= a or b;
    layer6_outputs(2561) <= not a or b;
    layer6_outputs(2562) <= not (a xor b);
    layer6_outputs(2563) <= b;
    layer6_outputs(2564) <= not a;
    layer6_outputs(2565) <= a;
    layer6_outputs(2566) <= not (a and b);
    layer6_outputs(2567) <= not (a xor b);
    layer6_outputs(2568) <= not a;
    layer6_outputs(2569) <= not a or b;
    layer6_outputs(2570) <= b and not a;
    layer6_outputs(2571) <= a or b;
    layer6_outputs(2572) <= not a;
    layer6_outputs(2573) <= a;
    layer6_outputs(2574) <= a;
    layer6_outputs(2575) <= a and b;
    layer6_outputs(2576) <= not b or a;
    layer6_outputs(2577) <= a xor b;
    layer6_outputs(2578) <= a xor b;
    layer6_outputs(2579) <= not (a and b);
    layer6_outputs(2580) <= a xor b;
    layer6_outputs(2581) <= not (a or b);
    layer6_outputs(2582) <= not (a and b);
    layer6_outputs(2583) <= not (a and b);
    layer6_outputs(2584) <= a;
    layer6_outputs(2585) <= not b;
    layer6_outputs(2586) <= a xor b;
    layer6_outputs(2587) <= not (a xor b);
    layer6_outputs(2588) <= not a;
    layer6_outputs(2589) <= not a;
    layer6_outputs(2590) <= not b;
    layer6_outputs(2591) <= not a;
    layer6_outputs(2592) <= not a;
    layer6_outputs(2593) <= a;
    layer6_outputs(2594) <= not a;
    layer6_outputs(2595) <= a and b;
    layer6_outputs(2596) <= not b or a;
    layer6_outputs(2597) <= not b;
    layer6_outputs(2598) <= a xor b;
    layer6_outputs(2599) <= a xor b;
    layer6_outputs(2600) <= not b;
    layer6_outputs(2601) <= not b or a;
    layer6_outputs(2602) <= a xor b;
    layer6_outputs(2603) <= not b;
    layer6_outputs(2604) <= not b;
    layer6_outputs(2605) <= a xor b;
    layer6_outputs(2606) <= not (a and b);
    layer6_outputs(2607) <= not a;
    layer6_outputs(2608) <= not (a xor b);
    layer6_outputs(2609) <= a and b;
    layer6_outputs(2610) <= b;
    layer6_outputs(2611) <= a or b;
    layer6_outputs(2612) <= not a;
    layer6_outputs(2613) <= not b;
    layer6_outputs(2614) <= not b;
    layer6_outputs(2615) <= not b;
    layer6_outputs(2616) <= a;
    layer6_outputs(2617) <= not b;
    layer6_outputs(2618) <= not (a xor b);
    layer6_outputs(2619) <= a xor b;
    layer6_outputs(2620) <= not b;
    layer6_outputs(2621) <= a xor b;
    layer6_outputs(2622) <= a xor b;
    layer6_outputs(2623) <= not b;
    layer6_outputs(2624) <= not b;
    layer6_outputs(2625) <= a xor b;
    layer6_outputs(2626) <= b;
    layer6_outputs(2627) <= a and b;
    layer6_outputs(2628) <= a xor b;
    layer6_outputs(2629) <= not a;
    layer6_outputs(2630) <= not a;
    layer6_outputs(2631) <= not b;
    layer6_outputs(2632) <= not (a or b);
    layer6_outputs(2633) <= not (a xor b);
    layer6_outputs(2634) <= a;
    layer6_outputs(2635) <= '1';
    layer6_outputs(2636) <= b;
    layer6_outputs(2637) <= a;
    layer6_outputs(2638) <= not (a xor b);
    layer6_outputs(2639) <= a or b;
    layer6_outputs(2640) <= not a;
    layer6_outputs(2641) <= a;
    layer6_outputs(2642) <= a;
    layer6_outputs(2643) <= a or b;
    layer6_outputs(2644) <= a or b;
    layer6_outputs(2645) <= not (a or b);
    layer6_outputs(2646) <= not (a xor b);
    layer6_outputs(2647) <= not (a and b);
    layer6_outputs(2648) <= not (a or b);
    layer6_outputs(2649) <= a xor b;
    layer6_outputs(2650) <= a xor b;
    layer6_outputs(2651) <= b;
    layer6_outputs(2652) <= not (a or b);
    layer6_outputs(2653) <= a;
    layer6_outputs(2654) <= a xor b;
    layer6_outputs(2655) <= not (a xor b);
    layer6_outputs(2656) <= a;
    layer6_outputs(2657) <= '1';
    layer6_outputs(2658) <= b;
    layer6_outputs(2659) <= a;
    layer6_outputs(2660) <= not a;
    layer6_outputs(2661) <= not b or a;
    layer6_outputs(2662) <= a;
    layer6_outputs(2663) <= not a or b;
    layer6_outputs(2664) <= not a;
    layer6_outputs(2665) <= b;
    layer6_outputs(2666) <= not (a or b);
    layer6_outputs(2667) <= not a or b;
    layer6_outputs(2668) <= not a;
    layer6_outputs(2669) <= a xor b;
    layer6_outputs(2670) <= a;
    layer6_outputs(2671) <= not (a xor b);
    layer6_outputs(2672) <= a;
    layer6_outputs(2673) <= b;
    layer6_outputs(2674) <= a xor b;
    layer6_outputs(2675) <= not b or a;
    layer6_outputs(2676) <= a;
    layer6_outputs(2677) <= not (a or b);
    layer6_outputs(2678) <= not a or b;
    layer6_outputs(2679) <= a;
    layer6_outputs(2680) <= not (a and b);
    layer6_outputs(2681) <= not b;
    layer6_outputs(2682) <= a and not b;
    layer6_outputs(2683) <= not (a xor b);
    layer6_outputs(2684) <= b;
    layer6_outputs(2685) <= not a;
    layer6_outputs(2686) <= not b;
    layer6_outputs(2687) <= not a;
    layer6_outputs(2688) <= not (a xor b);
    layer6_outputs(2689) <= not (a and b);
    layer6_outputs(2690) <= b and not a;
    layer6_outputs(2691) <= not (a and b);
    layer6_outputs(2692) <= not (a xor b);
    layer6_outputs(2693) <= a and b;
    layer6_outputs(2694) <= not a;
    layer6_outputs(2695) <= not b;
    layer6_outputs(2696) <= b and not a;
    layer6_outputs(2697) <= not (a and b);
    layer6_outputs(2698) <= b and not a;
    layer6_outputs(2699) <= not a;
    layer6_outputs(2700) <= a and b;
    layer6_outputs(2701) <= a and b;
    layer6_outputs(2702) <= a;
    layer6_outputs(2703) <= not (a or b);
    layer6_outputs(2704) <= not a;
    layer6_outputs(2705) <= b;
    layer6_outputs(2706) <= not (a xor b);
    layer6_outputs(2707) <= not b;
    layer6_outputs(2708) <= b;
    layer6_outputs(2709) <= not (a xor b);
    layer6_outputs(2710) <= a;
    layer6_outputs(2711) <= a;
    layer6_outputs(2712) <= a or b;
    layer6_outputs(2713) <= not (a xor b);
    layer6_outputs(2714) <= not (a xor b);
    layer6_outputs(2715) <= not a or b;
    layer6_outputs(2716) <= b;
    layer6_outputs(2717) <= a xor b;
    layer6_outputs(2718) <= not b or a;
    layer6_outputs(2719) <= a and not b;
    layer6_outputs(2720) <= not (a and b);
    layer6_outputs(2721) <= a and not b;
    layer6_outputs(2722) <= not b or a;
    layer6_outputs(2723) <= b;
    layer6_outputs(2724) <= not (a xor b);
    layer6_outputs(2725) <= a;
    layer6_outputs(2726) <= a and not b;
    layer6_outputs(2727) <= not (a xor b);
    layer6_outputs(2728) <= not b or a;
    layer6_outputs(2729) <= not b;
    layer6_outputs(2730) <= not b;
    layer6_outputs(2731) <= b;
    layer6_outputs(2732) <= not a;
    layer6_outputs(2733) <= a xor b;
    layer6_outputs(2734) <= b;
    layer6_outputs(2735) <= not (a and b);
    layer6_outputs(2736) <= b and not a;
    layer6_outputs(2737) <= not a;
    layer6_outputs(2738) <= a and b;
    layer6_outputs(2739) <= not b;
    layer6_outputs(2740) <= not a;
    layer6_outputs(2741) <= not (a xor b);
    layer6_outputs(2742) <= b;
    layer6_outputs(2743) <= not a or b;
    layer6_outputs(2744) <= a xor b;
    layer6_outputs(2745) <= not (a and b);
    layer6_outputs(2746) <= a and b;
    layer6_outputs(2747) <= not a;
    layer6_outputs(2748) <= b and not a;
    layer6_outputs(2749) <= b;
    layer6_outputs(2750) <= a xor b;
    layer6_outputs(2751) <= a and not b;
    layer6_outputs(2752) <= not a;
    layer6_outputs(2753) <= not a;
    layer6_outputs(2754) <= b;
    layer6_outputs(2755) <= b;
    layer6_outputs(2756) <= not a;
    layer6_outputs(2757) <= a xor b;
    layer6_outputs(2758) <= not (a and b);
    layer6_outputs(2759) <= b;
    layer6_outputs(2760) <= not a;
    layer6_outputs(2761) <= b;
    layer6_outputs(2762) <= a and not b;
    layer6_outputs(2763) <= a;
    layer6_outputs(2764) <= not a;
    layer6_outputs(2765) <= b;
    layer6_outputs(2766) <= not (a or b);
    layer6_outputs(2767) <= not (a or b);
    layer6_outputs(2768) <= not (a xor b);
    layer6_outputs(2769) <= not (a and b);
    layer6_outputs(2770) <= not a;
    layer6_outputs(2771) <= a;
    layer6_outputs(2772) <= not (a xor b);
    layer6_outputs(2773) <= not (a and b);
    layer6_outputs(2774) <= not a or b;
    layer6_outputs(2775) <= b;
    layer6_outputs(2776) <= a or b;
    layer6_outputs(2777) <= not a;
    layer6_outputs(2778) <= a;
    layer6_outputs(2779) <= b;
    layer6_outputs(2780) <= a and not b;
    layer6_outputs(2781) <= not (a xor b);
    layer6_outputs(2782) <= a and b;
    layer6_outputs(2783) <= a;
    layer6_outputs(2784) <= a or b;
    layer6_outputs(2785) <= a and b;
    layer6_outputs(2786) <= a and not b;
    layer6_outputs(2787) <= a xor b;
    layer6_outputs(2788) <= a;
    layer6_outputs(2789) <= a or b;
    layer6_outputs(2790) <= b;
    layer6_outputs(2791) <= not b;
    layer6_outputs(2792) <= a and not b;
    layer6_outputs(2793) <= not (a xor b);
    layer6_outputs(2794) <= not (a xor b);
    layer6_outputs(2795) <= not (a or b);
    layer6_outputs(2796) <= a and not b;
    layer6_outputs(2797) <= a;
    layer6_outputs(2798) <= not (a xor b);
    layer6_outputs(2799) <= not a;
    layer6_outputs(2800) <= a or b;
    layer6_outputs(2801) <= not a;
    layer6_outputs(2802) <= not a;
    layer6_outputs(2803) <= b;
    layer6_outputs(2804) <= a and b;
    layer6_outputs(2805) <= a;
    layer6_outputs(2806) <= not (a xor b);
    layer6_outputs(2807) <= not a;
    layer6_outputs(2808) <= not (a xor b);
    layer6_outputs(2809) <= a and b;
    layer6_outputs(2810) <= a;
    layer6_outputs(2811) <= '0';
    layer6_outputs(2812) <= not b;
    layer6_outputs(2813) <= a;
    layer6_outputs(2814) <= not b;
    layer6_outputs(2815) <= a xor b;
    layer6_outputs(2816) <= a xor b;
    layer6_outputs(2817) <= not (a xor b);
    layer6_outputs(2818) <= not (a or b);
    layer6_outputs(2819) <= a;
    layer6_outputs(2820) <= not (a or b);
    layer6_outputs(2821) <= a and b;
    layer6_outputs(2822) <= b and not a;
    layer6_outputs(2823) <= b;
    layer6_outputs(2824) <= not (a and b);
    layer6_outputs(2825) <= not (a or b);
    layer6_outputs(2826) <= not (a or b);
    layer6_outputs(2827) <= a;
    layer6_outputs(2828) <= not b;
    layer6_outputs(2829) <= not a;
    layer6_outputs(2830) <= not (a or b);
    layer6_outputs(2831) <= not (a xor b);
    layer6_outputs(2832) <= a or b;
    layer6_outputs(2833) <= not a;
    layer6_outputs(2834) <= not (a xor b);
    layer6_outputs(2835) <= b;
    layer6_outputs(2836) <= not a;
    layer6_outputs(2837) <= b and not a;
    layer6_outputs(2838) <= not (a xor b);
    layer6_outputs(2839) <= not (a xor b);
    layer6_outputs(2840) <= not a;
    layer6_outputs(2841) <= not b;
    layer6_outputs(2842) <= not a;
    layer6_outputs(2843) <= not a;
    layer6_outputs(2844) <= a;
    layer6_outputs(2845) <= b;
    layer6_outputs(2846) <= not a;
    layer6_outputs(2847) <= a;
    layer6_outputs(2848) <= b;
    layer6_outputs(2849) <= not b;
    layer6_outputs(2850) <= not a or b;
    layer6_outputs(2851) <= not (a xor b);
    layer6_outputs(2852) <= b;
    layer6_outputs(2853) <= a xor b;
    layer6_outputs(2854) <= not a;
    layer6_outputs(2855) <= not b or a;
    layer6_outputs(2856) <= not b;
    layer6_outputs(2857) <= not a or b;
    layer6_outputs(2858) <= a;
    layer6_outputs(2859) <= b and not a;
    layer6_outputs(2860) <= a and b;
    layer6_outputs(2861) <= not a;
    layer6_outputs(2862) <= not (a xor b);
    layer6_outputs(2863) <= not a;
    layer6_outputs(2864) <= b;
    layer6_outputs(2865) <= not (a xor b);
    layer6_outputs(2866) <= not b;
    layer6_outputs(2867) <= a or b;
    layer6_outputs(2868) <= '0';
    layer6_outputs(2869) <= not b;
    layer6_outputs(2870) <= not (a or b);
    layer6_outputs(2871) <= a;
    layer6_outputs(2872) <= not (a xor b);
    layer6_outputs(2873) <= not (a and b);
    layer6_outputs(2874) <= b;
    layer6_outputs(2875) <= a;
    layer6_outputs(2876) <= b;
    layer6_outputs(2877) <= a;
    layer6_outputs(2878) <= b;
    layer6_outputs(2879) <= '1';
    layer6_outputs(2880) <= a and not b;
    layer6_outputs(2881) <= a or b;
    layer6_outputs(2882) <= '0';
    layer6_outputs(2883) <= not a or b;
    layer6_outputs(2884) <= a;
    layer6_outputs(2885) <= not b or a;
    layer6_outputs(2886) <= not a or b;
    layer6_outputs(2887) <= not b;
    layer6_outputs(2888) <= a;
    layer6_outputs(2889) <= '1';
    layer6_outputs(2890) <= not b;
    layer6_outputs(2891) <= not (a xor b);
    layer6_outputs(2892) <= not a;
    layer6_outputs(2893) <= not b;
    layer6_outputs(2894) <= a;
    layer6_outputs(2895) <= b;
    layer6_outputs(2896) <= not b;
    layer6_outputs(2897) <= a xor b;
    layer6_outputs(2898) <= not (a xor b);
    layer6_outputs(2899) <= b;
    layer6_outputs(2900) <= b;
    layer6_outputs(2901) <= not b;
    layer6_outputs(2902) <= not (a xor b);
    layer6_outputs(2903) <= a and not b;
    layer6_outputs(2904) <= a;
    layer6_outputs(2905) <= b and not a;
    layer6_outputs(2906) <= not b;
    layer6_outputs(2907) <= b;
    layer6_outputs(2908) <= a and b;
    layer6_outputs(2909) <= b;
    layer6_outputs(2910) <= a or b;
    layer6_outputs(2911) <= not b or a;
    layer6_outputs(2912) <= not (a xor b);
    layer6_outputs(2913) <= a xor b;
    layer6_outputs(2914) <= a or b;
    layer6_outputs(2915) <= not (a xor b);
    layer6_outputs(2916) <= b;
    layer6_outputs(2917) <= a;
    layer6_outputs(2918) <= not a;
    layer6_outputs(2919) <= not (a xor b);
    layer6_outputs(2920) <= not a;
    layer6_outputs(2921) <= not (a or b);
    layer6_outputs(2922) <= b;
    layer6_outputs(2923) <= a xor b;
    layer6_outputs(2924) <= not b;
    layer6_outputs(2925) <= not (a xor b);
    layer6_outputs(2926) <= not a or b;
    layer6_outputs(2927) <= not (a or b);
    layer6_outputs(2928) <= a;
    layer6_outputs(2929) <= not b;
    layer6_outputs(2930) <= not a;
    layer6_outputs(2931) <= a;
    layer6_outputs(2932) <= not a or b;
    layer6_outputs(2933) <= b;
    layer6_outputs(2934) <= a xor b;
    layer6_outputs(2935) <= not a;
    layer6_outputs(2936) <= not a;
    layer6_outputs(2937) <= a;
    layer6_outputs(2938) <= b;
    layer6_outputs(2939) <= a or b;
    layer6_outputs(2940) <= not a;
    layer6_outputs(2941) <= not (a xor b);
    layer6_outputs(2942) <= not (a and b);
    layer6_outputs(2943) <= a xor b;
    layer6_outputs(2944) <= b and not a;
    layer6_outputs(2945) <= not b or a;
    layer6_outputs(2946) <= a and b;
    layer6_outputs(2947) <= not a;
    layer6_outputs(2948) <= a and b;
    layer6_outputs(2949) <= not (a xor b);
    layer6_outputs(2950) <= not (a or b);
    layer6_outputs(2951) <= not (a xor b);
    layer6_outputs(2952) <= not b;
    layer6_outputs(2953) <= not b;
    layer6_outputs(2954) <= not a;
    layer6_outputs(2955) <= not b;
    layer6_outputs(2956) <= not a;
    layer6_outputs(2957) <= a and not b;
    layer6_outputs(2958) <= not a;
    layer6_outputs(2959) <= not b or a;
    layer6_outputs(2960) <= a xor b;
    layer6_outputs(2961) <= a and not b;
    layer6_outputs(2962) <= a and b;
    layer6_outputs(2963) <= b;
    layer6_outputs(2964) <= not (a xor b);
    layer6_outputs(2965) <= a xor b;
    layer6_outputs(2966) <= not a;
    layer6_outputs(2967) <= a;
    layer6_outputs(2968) <= not (a or b);
    layer6_outputs(2969) <= a xor b;
    layer6_outputs(2970) <= not b;
    layer6_outputs(2971) <= b;
    layer6_outputs(2972) <= not (a xor b);
    layer6_outputs(2973) <= not a;
    layer6_outputs(2974) <= a;
    layer6_outputs(2975) <= b;
    layer6_outputs(2976) <= not (a xor b);
    layer6_outputs(2977) <= not (a and b);
    layer6_outputs(2978) <= a and b;
    layer6_outputs(2979) <= a;
    layer6_outputs(2980) <= b;
    layer6_outputs(2981) <= a xor b;
    layer6_outputs(2982) <= not a;
    layer6_outputs(2983) <= not b;
    layer6_outputs(2984) <= a;
    layer6_outputs(2985) <= a;
    layer6_outputs(2986) <= not (a and b);
    layer6_outputs(2987) <= not (a xor b);
    layer6_outputs(2988) <= '1';
    layer6_outputs(2989) <= a;
    layer6_outputs(2990) <= b;
    layer6_outputs(2991) <= not b;
    layer6_outputs(2992) <= b;
    layer6_outputs(2993) <= not (a or b);
    layer6_outputs(2994) <= not (a xor b);
    layer6_outputs(2995) <= not b;
    layer6_outputs(2996) <= a;
    layer6_outputs(2997) <= a;
    layer6_outputs(2998) <= not b;
    layer6_outputs(2999) <= a;
    layer6_outputs(3000) <= b;
    layer6_outputs(3001) <= a xor b;
    layer6_outputs(3002) <= a;
    layer6_outputs(3003) <= not (a xor b);
    layer6_outputs(3004) <= a or b;
    layer6_outputs(3005) <= not b;
    layer6_outputs(3006) <= a xor b;
    layer6_outputs(3007) <= a and not b;
    layer6_outputs(3008) <= a xor b;
    layer6_outputs(3009) <= not b;
    layer6_outputs(3010) <= a;
    layer6_outputs(3011) <= not a or b;
    layer6_outputs(3012) <= b;
    layer6_outputs(3013) <= not b;
    layer6_outputs(3014) <= a and not b;
    layer6_outputs(3015) <= not (a xor b);
    layer6_outputs(3016) <= a xor b;
    layer6_outputs(3017) <= not a;
    layer6_outputs(3018) <= not (a and b);
    layer6_outputs(3019) <= not b or a;
    layer6_outputs(3020) <= a;
    layer6_outputs(3021) <= not b;
    layer6_outputs(3022) <= a and not b;
    layer6_outputs(3023) <= not b;
    layer6_outputs(3024) <= b and not a;
    layer6_outputs(3025) <= not b;
    layer6_outputs(3026) <= b and not a;
    layer6_outputs(3027) <= a xor b;
    layer6_outputs(3028) <= a;
    layer6_outputs(3029) <= b and not a;
    layer6_outputs(3030) <= not (a xor b);
    layer6_outputs(3031) <= a and not b;
    layer6_outputs(3032) <= b and not a;
    layer6_outputs(3033) <= b and not a;
    layer6_outputs(3034) <= not a;
    layer6_outputs(3035) <= not (a or b);
    layer6_outputs(3036) <= a and not b;
    layer6_outputs(3037) <= a and b;
    layer6_outputs(3038) <= not (a xor b);
    layer6_outputs(3039) <= not (a or b);
    layer6_outputs(3040) <= a or b;
    layer6_outputs(3041) <= not b or a;
    layer6_outputs(3042) <= b;
    layer6_outputs(3043) <= a and not b;
    layer6_outputs(3044) <= not b;
    layer6_outputs(3045) <= a xor b;
    layer6_outputs(3046) <= a or b;
    layer6_outputs(3047) <= not a;
    layer6_outputs(3048) <= not b;
    layer6_outputs(3049) <= b;
    layer6_outputs(3050) <= not a or b;
    layer6_outputs(3051) <= a xor b;
    layer6_outputs(3052) <= a and b;
    layer6_outputs(3053) <= a;
    layer6_outputs(3054) <= not (a and b);
    layer6_outputs(3055) <= a and b;
    layer6_outputs(3056) <= b;
    layer6_outputs(3057) <= a xor b;
    layer6_outputs(3058) <= a xor b;
    layer6_outputs(3059) <= a;
    layer6_outputs(3060) <= b;
    layer6_outputs(3061) <= not a;
    layer6_outputs(3062) <= not b;
    layer6_outputs(3063) <= b;
    layer6_outputs(3064) <= b and not a;
    layer6_outputs(3065) <= not a or b;
    layer6_outputs(3066) <= not (a or b);
    layer6_outputs(3067) <= not a;
    layer6_outputs(3068) <= not a;
    layer6_outputs(3069) <= a xor b;
    layer6_outputs(3070) <= not b or a;
    layer6_outputs(3071) <= a xor b;
    layer6_outputs(3072) <= not a;
    layer6_outputs(3073) <= a or b;
    layer6_outputs(3074) <= a or b;
    layer6_outputs(3075) <= a xor b;
    layer6_outputs(3076) <= not (a xor b);
    layer6_outputs(3077) <= not a or b;
    layer6_outputs(3078) <= b;
    layer6_outputs(3079) <= '1';
    layer6_outputs(3080) <= a and b;
    layer6_outputs(3081) <= not a;
    layer6_outputs(3082) <= a xor b;
    layer6_outputs(3083) <= b;
    layer6_outputs(3084) <= not (a xor b);
    layer6_outputs(3085) <= a xor b;
    layer6_outputs(3086) <= a and not b;
    layer6_outputs(3087) <= not a;
    layer6_outputs(3088) <= not a or b;
    layer6_outputs(3089) <= not a or b;
    layer6_outputs(3090) <= not b or a;
    layer6_outputs(3091) <= not a;
    layer6_outputs(3092) <= b;
    layer6_outputs(3093) <= not b;
    layer6_outputs(3094) <= a;
    layer6_outputs(3095) <= not (a or b);
    layer6_outputs(3096) <= a;
    layer6_outputs(3097) <= not a;
    layer6_outputs(3098) <= not a;
    layer6_outputs(3099) <= a and b;
    layer6_outputs(3100) <= not a or b;
    layer6_outputs(3101) <= not b;
    layer6_outputs(3102) <= a;
    layer6_outputs(3103) <= b;
    layer6_outputs(3104) <= not a or b;
    layer6_outputs(3105) <= a;
    layer6_outputs(3106) <= a and b;
    layer6_outputs(3107) <= not a;
    layer6_outputs(3108) <= not b;
    layer6_outputs(3109) <= b;
    layer6_outputs(3110) <= not a;
    layer6_outputs(3111) <= not b;
    layer6_outputs(3112) <= not a or b;
    layer6_outputs(3113) <= b;
    layer6_outputs(3114) <= a xor b;
    layer6_outputs(3115) <= not a or b;
    layer6_outputs(3116) <= not a;
    layer6_outputs(3117) <= not b;
    layer6_outputs(3118) <= not b;
    layer6_outputs(3119) <= not (a or b);
    layer6_outputs(3120) <= not a;
    layer6_outputs(3121) <= b;
    layer6_outputs(3122) <= not a or b;
    layer6_outputs(3123) <= a and b;
    layer6_outputs(3124) <= b;
    layer6_outputs(3125) <= not b;
    layer6_outputs(3126) <= not b;
    layer6_outputs(3127) <= not b;
    layer6_outputs(3128) <= a;
    layer6_outputs(3129) <= a or b;
    layer6_outputs(3130) <= a or b;
    layer6_outputs(3131) <= a;
    layer6_outputs(3132) <= a and not b;
    layer6_outputs(3133) <= a or b;
    layer6_outputs(3134) <= not (a xor b);
    layer6_outputs(3135) <= not (a xor b);
    layer6_outputs(3136) <= a xor b;
    layer6_outputs(3137) <= b;
    layer6_outputs(3138) <= b;
    layer6_outputs(3139) <= a and not b;
    layer6_outputs(3140) <= a or b;
    layer6_outputs(3141) <= not b;
    layer6_outputs(3142) <= not a or b;
    layer6_outputs(3143) <= b;
    layer6_outputs(3144) <= a and not b;
    layer6_outputs(3145) <= not b;
    layer6_outputs(3146) <= a xor b;
    layer6_outputs(3147) <= not a;
    layer6_outputs(3148) <= a;
    layer6_outputs(3149) <= not a;
    layer6_outputs(3150) <= not b or a;
    layer6_outputs(3151) <= not (a xor b);
    layer6_outputs(3152) <= '1';
    layer6_outputs(3153) <= not (a and b);
    layer6_outputs(3154) <= b;
    layer6_outputs(3155) <= not a;
    layer6_outputs(3156) <= not a;
    layer6_outputs(3157) <= not b;
    layer6_outputs(3158) <= a xor b;
    layer6_outputs(3159) <= not (a and b);
    layer6_outputs(3160) <= a or b;
    layer6_outputs(3161) <= not b;
    layer6_outputs(3162) <= not (a xor b);
    layer6_outputs(3163) <= not (a and b);
    layer6_outputs(3164) <= not a or b;
    layer6_outputs(3165) <= b;
    layer6_outputs(3166) <= not (a or b);
    layer6_outputs(3167) <= a;
    layer6_outputs(3168) <= not b;
    layer6_outputs(3169) <= a xor b;
    layer6_outputs(3170) <= a;
    layer6_outputs(3171) <= not (a and b);
    layer6_outputs(3172) <= a;
    layer6_outputs(3173) <= not a;
    layer6_outputs(3174) <= not b;
    layer6_outputs(3175) <= not (a or b);
    layer6_outputs(3176) <= not a or b;
    layer6_outputs(3177) <= not (a xor b);
    layer6_outputs(3178) <= a or b;
    layer6_outputs(3179) <= not b;
    layer6_outputs(3180) <= a xor b;
    layer6_outputs(3181) <= b;
    layer6_outputs(3182) <= not (a or b);
    layer6_outputs(3183) <= not b;
    layer6_outputs(3184) <= not b;
    layer6_outputs(3185) <= a xor b;
    layer6_outputs(3186) <= not b;
    layer6_outputs(3187) <= a xor b;
    layer6_outputs(3188) <= not a;
    layer6_outputs(3189) <= a and b;
    layer6_outputs(3190) <= not b;
    layer6_outputs(3191) <= not (a xor b);
    layer6_outputs(3192) <= '0';
    layer6_outputs(3193) <= not a;
    layer6_outputs(3194) <= not a;
    layer6_outputs(3195) <= b;
    layer6_outputs(3196) <= a or b;
    layer6_outputs(3197) <= not (a or b);
    layer6_outputs(3198) <= not (a or b);
    layer6_outputs(3199) <= not b;
    layer6_outputs(3200) <= not a;
    layer6_outputs(3201) <= not (a or b);
    layer6_outputs(3202) <= b and not a;
    layer6_outputs(3203) <= b;
    layer6_outputs(3204) <= a;
    layer6_outputs(3205) <= b;
    layer6_outputs(3206) <= a or b;
    layer6_outputs(3207) <= not b;
    layer6_outputs(3208) <= a xor b;
    layer6_outputs(3209) <= a;
    layer6_outputs(3210) <= a or b;
    layer6_outputs(3211) <= a and b;
    layer6_outputs(3212) <= a and not b;
    layer6_outputs(3213) <= a and not b;
    layer6_outputs(3214) <= a xor b;
    layer6_outputs(3215) <= a and not b;
    layer6_outputs(3216) <= not a;
    layer6_outputs(3217) <= b;
    layer6_outputs(3218) <= not b or a;
    layer6_outputs(3219) <= a and not b;
    layer6_outputs(3220) <= not b or a;
    layer6_outputs(3221) <= b;
    layer6_outputs(3222) <= not b;
    layer6_outputs(3223) <= not a;
    layer6_outputs(3224) <= not (a and b);
    layer6_outputs(3225) <= not a;
    layer6_outputs(3226) <= b;
    layer6_outputs(3227) <= not a;
    layer6_outputs(3228) <= not b or a;
    layer6_outputs(3229) <= b;
    layer6_outputs(3230) <= not (a xor b);
    layer6_outputs(3231) <= not a or b;
    layer6_outputs(3232) <= a;
    layer6_outputs(3233) <= not (a xor b);
    layer6_outputs(3234) <= b;
    layer6_outputs(3235) <= b and not a;
    layer6_outputs(3236) <= not (a and b);
    layer6_outputs(3237) <= a or b;
    layer6_outputs(3238) <= not a;
    layer6_outputs(3239) <= not a or b;
    layer6_outputs(3240) <= b;
    layer6_outputs(3241) <= not b;
    layer6_outputs(3242) <= not a;
    layer6_outputs(3243) <= not (a xor b);
    layer6_outputs(3244) <= not (a xor b);
    layer6_outputs(3245) <= not a;
    layer6_outputs(3246) <= not a or b;
    layer6_outputs(3247) <= not a;
    layer6_outputs(3248) <= b;
    layer6_outputs(3249) <= a and b;
    layer6_outputs(3250) <= a;
    layer6_outputs(3251) <= a;
    layer6_outputs(3252) <= b;
    layer6_outputs(3253) <= not a;
    layer6_outputs(3254) <= '0';
    layer6_outputs(3255) <= not a;
    layer6_outputs(3256) <= not b;
    layer6_outputs(3257) <= not a;
    layer6_outputs(3258) <= b;
    layer6_outputs(3259) <= not b or a;
    layer6_outputs(3260) <= not a;
    layer6_outputs(3261) <= a xor b;
    layer6_outputs(3262) <= not (a xor b);
    layer6_outputs(3263) <= not a;
    layer6_outputs(3264) <= a xor b;
    layer6_outputs(3265) <= b;
    layer6_outputs(3266) <= a;
    layer6_outputs(3267) <= a;
    layer6_outputs(3268) <= not b;
    layer6_outputs(3269) <= a and b;
    layer6_outputs(3270) <= not b;
    layer6_outputs(3271) <= b;
    layer6_outputs(3272) <= not (a and b);
    layer6_outputs(3273) <= not (a or b);
    layer6_outputs(3274) <= a;
    layer6_outputs(3275) <= a xor b;
    layer6_outputs(3276) <= a xor b;
    layer6_outputs(3277) <= not b;
    layer6_outputs(3278) <= not a;
    layer6_outputs(3279) <= a xor b;
    layer6_outputs(3280) <= not a;
    layer6_outputs(3281) <= not b;
    layer6_outputs(3282) <= not a;
    layer6_outputs(3283) <= not (a xor b);
    layer6_outputs(3284) <= not a;
    layer6_outputs(3285) <= b and not a;
    layer6_outputs(3286) <= a and not b;
    layer6_outputs(3287) <= b;
    layer6_outputs(3288) <= not (a xor b);
    layer6_outputs(3289) <= not b;
    layer6_outputs(3290) <= not (a or b);
    layer6_outputs(3291) <= not (a xor b);
    layer6_outputs(3292) <= not b;
    layer6_outputs(3293) <= a xor b;
    layer6_outputs(3294) <= not (a and b);
    layer6_outputs(3295) <= not a or b;
    layer6_outputs(3296) <= a xor b;
    layer6_outputs(3297) <= not a;
    layer6_outputs(3298) <= not (a and b);
    layer6_outputs(3299) <= a xor b;
    layer6_outputs(3300) <= not b;
    layer6_outputs(3301) <= not b;
    layer6_outputs(3302) <= a;
    layer6_outputs(3303) <= not b;
    layer6_outputs(3304) <= not (a or b);
    layer6_outputs(3305) <= not b;
    layer6_outputs(3306) <= not b;
    layer6_outputs(3307) <= a and b;
    layer6_outputs(3308) <= a;
    layer6_outputs(3309) <= b;
    layer6_outputs(3310) <= not a;
    layer6_outputs(3311) <= a and not b;
    layer6_outputs(3312) <= not (a xor b);
    layer6_outputs(3313) <= not b or a;
    layer6_outputs(3314) <= not (a xor b);
    layer6_outputs(3315) <= a and not b;
    layer6_outputs(3316) <= a xor b;
    layer6_outputs(3317) <= not (a xor b);
    layer6_outputs(3318) <= a;
    layer6_outputs(3319) <= not (a xor b);
    layer6_outputs(3320) <= not (a xor b);
    layer6_outputs(3321) <= a and not b;
    layer6_outputs(3322) <= not b;
    layer6_outputs(3323) <= not b;
    layer6_outputs(3324) <= not (a and b);
    layer6_outputs(3325) <= b;
    layer6_outputs(3326) <= a and b;
    layer6_outputs(3327) <= a xor b;
    layer6_outputs(3328) <= a xor b;
    layer6_outputs(3329) <= b;
    layer6_outputs(3330) <= a;
    layer6_outputs(3331) <= a;
    layer6_outputs(3332) <= not (a xor b);
    layer6_outputs(3333) <= not a or b;
    layer6_outputs(3334) <= not a;
    layer6_outputs(3335) <= a xor b;
    layer6_outputs(3336) <= b;
    layer6_outputs(3337) <= not b;
    layer6_outputs(3338) <= not b;
    layer6_outputs(3339) <= not a;
    layer6_outputs(3340) <= a;
    layer6_outputs(3341) <= b;
    layer6_outputs(3342) <= not a;
    layer6_outputs(3343) <= not b or a;
    layer6_outputs(3344) <= not a;
    layer6_outputs(3345) <= not (a or b);
    layer6_outputs(3346) <= not a;
    layer6_outputs(3347) <= a and not b;
    layer6_outputs(3348) <= not (a or b);
    layer6_outputs(3349) <= a and not b;
    layer6_outputs(3350) <= not a;
    layer6_outputs(3351) <= a and b;
    layer6_outputs(3352) <= a;
    layer6_outputs(3353) <= a and b;
    layer6_outputs(3354) <= not b or a;
    layer6_outputs(3355) <= not (a xor b);
    layer6_outputs(3356) <= a;
    layer6_outputs(3357) <= not (a and b);
    layer6_outputs(3358) <= not a;
    layer6_outputs(3359) <= not a;
    layer6_outputs(3360) <= not (a xor b);
    layer6_outputs(3361) <= not (a xor b);
    layer6_outputs(3362) <= a or b;
    layer6_outputs(3363) <= b;
    layer6_outputs(3364) <= not a;
    layer6_outputs(3365) <= not (a and b);
    layer6_outputs(3366) <= not a;
    layer6_outputs(3367) <= not (a xor b);
    layer6_outputs(3368) <= a;
    layer6_outputs(3369) <= not b;
    layer6_outputs(3370) <= a;
    layer6_outputs(3371) <= a or b;
    layer6_outputs(3372) <= not (a xor b);
    layer6_outputs(3373) <= not a or b;
    layer6_outputs(3374) <= b and not a;
    layer6_outputs(3375) <= b;
    layer6_outputs(3376) <= not b;
    layer6_outputs(3377) <= not a;
    layer6_outputs(3378) <= a xor b;
    layer6_outputs(3379) <= not (a and b);
    layer6_outputs(3380) <= b;
    layer6_outputs(3381) <= a;
    layer6_outputs(3382) <= a xor b;
    layer6_outputs(3383) <= a and not b;
    layer6_outputs(3384) <= '1';
    layer6_outputs(3385) <= not b;
    layer6_outputs(3386) <= a or b;
    layer6_outputs(3387) <= a xor b;
    layer6_outputs(3388) <= a;
    layer6_outputs(3389) <= a or b;
    layer6_outputs(3390) <= not b;
    layer6_outputs(3391) <= not b;
    layer6_outputs(3392) <= not (a or b);
    layer6_outputs(3393) <= b;
    layer6_outputs(3394) <= b;
    layer6_outputs(3395) <= not (a xor b);
    layer6_outputs(3396) <= a;
    layer6_outputs(3397) <= a and not b;
    layer6_outputs(3398) <= not a;
    layer6_outputs(3399) <= not (a or b);
    layer6_outputs(3400) <= not a;
    layer6_outputs(3401) <= a xor b;
    layer6_outputs(3402) <= a;
    layer6_outputs(3403) <= not b;
    layer6_outputs(3404) <= not (a and b);
    layer6_outputs(3405) <= not a;
    layer6_outputs(3406) <= a;
    layer6_outputs(3407) <= a and b;
    layer6_outputs(3408) <= not a;
    layer6_outputs(3409) <= b and not a;
    layer6_outputs(3410) <= b;
    layer6_outputs(3411) <= not a;
    layer6_outputs(3412) <= a and b;
    layer6_outputs(3413) <= a xor b;
    layer6_outputs(3414) <= not (a and b);
    layer6_outputs(3415) <= a and not b;
    layer6_outputs(3416) <= not (a and b);
    layer6_outputs(3417) <= a;
    layer6_outputs(3418) <= a xor b;
    layer6_outputs(3419) <= a;
    layer6_outputs(3420) <= not b;
    layer6_outputs(3421) <= a and b;
    layer6_outputs(3422) <= not a;
    layer6_outputs(3423) <= not a;
    layer6_outputs(3424) <= a;
    layer6_outputs(3425) <= b;
    layer6_outputs(3426) <= a xor b;
    layer6_outputs(3427) <= a xor b;
    layer6_outputs(3428) <= a and not b;
    layer6_outputs(3429) <= not a;
    layer6_outputs(3430) <= not b;
    layer6_outputs(3431) <= not (a or b);
    layer6_outputs(3432) <= not a or b;
    layer6_outputs(3433) <= a xor b;
    layer6_outputs(3434) <= not b;
    layer6_outputs(3435) <= a;
    layer6_outputs(3436) <= b;
    layer6_outputs(3437) <= not a;
    layer6_outputs(3438) <= not (a xor b);
    layer6_outputs(3439) <= a xor b;
    layer6_outputs(3440) <= not a;
    layer6_outputs(3441) <= b and not a;
    layer6_outputs(3442) <= not a;
    layer6_outputs(3443) <= a xor b;
    layer6_outputs(3444) <= b and not a;
    layer6_outputs(3445) <= a;
    layer6_outputs(3446) <= not (a and b);
    layer6_outputs(3447) <= a;
    layer6_outputs(3448) <= not b;
    layer6_outputs(3449) <= not a;
    layer6_outputs(3450) <= a and not b;
    layer6_outputs(3451) <= not a;
    layer6_outputs(3452) <= not (a xor b);
    layer6_outputs(3453) <= a and b;
    layer6_outputs(3454) <= a and b;
    layer6_outputs(3455) <= a and not b;
    layer6_outputs(3456) <= a xor b;
    layer6_outputs(3457) <= a and not b;
    layer6_outputs(3458) <= not a or b;
    layer6_outputs(3459) <= a;
    layer6_outputs(3460) <= not (a xor b);
    layer6_outputs(3461) <= not b;
    layer6_outputs(3462) <= a xor b;
    layer6_outputs(3463) <= not a;
    layer6_outputs(3464) <= a or b;
    layer6_outputs(3465) <= a and not b;
    layer6_outputs(3466) <= not b;
    layer6_outputs(3467) <= not (a and b);
    layer6_outputs(3468) <= not a;
    layer6_outputs(3469) <= not b;
    layer6_outputs(3470) <= b;
    layer6_outputs(3471) <= a xor b;
    layer6_outputs(3472) <= not b or a;
    layer6_outputs(3473) <= not a;
    layer6_outputs(3474) <= not a or b;
    layer6_outputs(3475) <= not (a xor b);
    layer6_outputs(3476) <= not b;
    layer6_outputs(3477) <= a xor b;
    layer6_outputs(3478) <= a;
    layer6_outputs(3479) <= b;
    layer6_outputs(3480) <= not a or b;
    layer6_outputs(3481) <= a and not b;
    layer6_outputs(3482) <= not b;
    layer6_outputs(3483) <= b;
    layer6_outputs(3484) <= a and b;
    layer6_outputs(3485) <= not a;
    layer6_outputs(3486) <= not b;
    layer6_outputs(3487) <= not b or a;
    layer6_outputs(3488) <= b and not a;
    layer6_outputs(3489) <= a xor b;
    layer6_outputs(3490) <= a and b;
    layer6_outputs(3491) <= not b or a;
    layer6_outputs(3492) <= a xor b;
    layer6_outputs(3493) <= b;
    layer6_outputs(3494) <= not b;
    layer6_outputs(3495) <= a xor b;
    layer6_outputs(3496) <= a xor b;
    layer6_outputs(3497) <= not b;
    layer6_outputs(3498) <= not b;
    layer6_outputs(3499) <= a or b;
    layer6_outputs(3500) <= b;
    layer6_outputs(3501) <= not a;
    layer6_outputs(3502) <= a;
    layer6_outputs(3503) <= not (a or b);
    layer6_outputs(3504) <= not (a xor b);
    layer6_outputs(3505) <= not b;
    layer6_outputs(3506) <= b;
    layer6_outputs(3507) <= not b;
    layer6_outputs(3508) <= a and b;
    layer6_outputs(3509) <= a;
    layer6_outputs(3510) <= not a;
    layer6_outputs(3511) <= not a;
    layer6_outputs(3512) <= not (a or b);
    layer6_outputs(3513) <= a;
    layer6_outputs(3514) <= not (a and b);
    layer6_outputs(3515) <= not (a xor b);
    layer6_outputs(3516) <= not (a xor b);
    layer6_outputs(3517) <= not a;
    layer6_outputs(3518) <= a;
    layer6_outputs(3519) <= a xor b;
    layer6_outputs(3520) <= a;
    layer6_outputs(3521) <= a;
    layer6_outputs(3522) <= a and not b;
    layer6_outputs(3523) <= not b;
    layer6_outputs(3524) <= a and not b;
    layer6_outputs(3525) <= not b;
    layer6_outputs(3526) <= not a or b;
    layer6_outputs(3527) <= b;
    layer6_outputs(3528) <= a;
    layer6_outputs(3529) <= a and not b;
    layer6_outputs(3530) <= a;
    layer6_outputs(3531) <= b;
    layer6_outputs(3532) <= a xor b;
    layer6_outputs(3533) <= b;
    layer6_outputs(3534) <= not (a xor b);
    layer6_outputs(3535) <= a;
    layer6_outputs(3536) <= not b;
    layer6_outputs(3537) <= not a;
    layer6_outputs(3538) <= not (a xor b);
    layer6_outputs(3539) <= not b;
    layer6_outputs(3540) <= b;
    layer6_outputs(3541) <= b and not a;
    layer6_outputs(3542) <= a xor b;
    layer6_outputs(3543) <= b and not a;
    layer6_outputs(3544) <= not a;
    layer6_outputs(3545) <= a xor b;
    layer6_outputs(3546) <= not (a or b);
    layer6_outputs(3547) <= a xor b;
    layer6_outputs(3548) <= not a;
    layer6_outputs(3549) <= not (a or b);
    layer6_outputs(3550) <= b;
    layer6_outputs(3551) <= not a;
    layer6_outputs(3552) <= a;
    layer6_outputs(3553) <= a;
    layer6_outputs(3554) <= not a or b;
    layer6_outputs(3555) <= a;
    layer6_outputs(3556) <= a or b;
    layer6_outputs(3557) <= not (a and b);
    layer6_outputs(3558) <= not b;
    layer6_outputs(3559) <= not b or a;
    layer6_outputs(3560) <= not b;
    layer6_outputs(3561) <= a xor b;
    layer6_outputs(3562) <= a and not b;
    layer6_outputs(3563) <= not (a xor b);
    layer6_outputs(3564) <= b;
    layer6_outputs(3565) <= not a or b;
    layer6_outputs(3566) <= not (a or b);
    layer6_outputs(3567) <= a;
    layer6_outputs(3568) <= a;
    layer6_outputs(3569) <= a;
    layer6_outputs(3570) <= a or b;
    layer6_outputs(3571) <= not a;
    layer6_outputs(3572) <= not a;
    layer6_outputs(3573) <= a and not b;
    layer6_outputs(3574) <= b;
    layer6_outputs(3575) <= not a;
    layer6_outputs(3576) <= a;
    layer6_outputs(3577) <= not (a xor b);
    layer6_outputs(3578) <= not (a or b);
    layer6_outputs(3579) <= not (a or b);
    layer6_outputs(3580) <= not a;
    layer6_outputs(3581) <= b;
    layer6_outputs(3582) <= not a;
    layer6_outputs(3583) <= not a;
    layer6_outputs(3584) <= a;
    layer6_outputs(3585) <= a or b;
    layer6_outputs(3586) <= a;
    layer6_outputs(3587) <= not (a xor b);
    layer6_outputs(3588) <= a xor b;
    layer6_outputs(3589) <= a;
    layer6_outputs(3590) <= not a;
    layer6_outputs(3591) <= b;
    layer6_outputs(3592) <= not a or b;
    layer6_outputs(3593) <= not (a xor b);
    layer6_outputs(3594) <= not a;
    layer6_outputs(3595) <= not a;
    layer6_outputs(3596) <= b;
    layer6_outputs(3597) <= not (a xor b);
    layer6_outputs(3598) <= a xor b;
    layer6_outputs(3599) <= not (a xor b);
    layer6_outputs(3600) <= b;
    layer6_outputs(3601) <= a or b;
    layer6_outputs(3602) <= not (a and b);
    layer6_outputs(3603) <= not (a xor b);
    layer6_outputs(3604) <= not (a and b);
    layer6_outputs(3605) <= a;
    layer6_outputs(3606) <= a and not b;
    layer6_outputs(3607) <= a;
    layer6_outputs(3608) <= a;
    layer6_outputs(3609) <= not a;
    layer6_outputs(3610) <= a xor b;
    layer6_outputs(3611) <= b and not a;
    layer6_outputs(3612) <= a xor b;
    layer6_outputs(3613) <= not b;
    layer6_outputs(3614) <= a;
    layer6_outputs(3615) <= a and not b;
    layer6_outputs(3616) <= a;
    layer6_outputs(3617) <= not a or b;
    layer6_outputs(3618) <= a;
    layer6_outputs(3619) <= not b;
    layer6_outputs(3620) <= not a or b;
    layer6_outputs(3621) <= not b;
    layer6_outputs(3622) <= not a;
    layer6_outputs(3623) <= b and not a;
    layer6_outputs(3624) <= not (a or b);
    layer6_outputs(3625) <= not a;
    layer6_outputs(3626) <= not a;
    layer6_outputs(3627) <= b and not a;
    layer6_outputs(3628) <= b and not a;
    layer6_outputs(3629) <= b;
    layer6_outputs(3630) <= not a;
    layer6_outputs(3631) <= b;
    layer6_outputs(3632) <= a or b;
    layer6_outputs(3633) <= not a;
    layer6_outputs(3634) <= a or b;
    layer6_outputs(3635) <= not a or b;
    layer6_outputs(3636) <= b and not a;
    layer6_outputs(3637) <= b;
    layer6_outputs(3638) <= a xor b;
    layer6_outputs(3639) <= b;
    layer6_outputs(3640) <= not (a xor b);
    layer6_outputs(3641) <= a;
    layer6_outputs(3642) <= not b;
    layer6_outputs(3643) <= not a;
    layer6_outputs(3644) <= not (a xor b);
    layer6_outputs(3645) <= not b or a;
    layer6_outputs(3646) <= '1';
    layer6_outputs(3647) <= not b;
    layer6_outputs(3648) <= not a;
    layer6_outputs(3649) <= a and not b;
    layer6_outputs(3650) <= a xor b;
    layer6_outputs(3651) <= b and not a;
    layer6_outputs(3652) <= not b;
    layer6_outputs(3653) <= a and not b;
    layer6_outputs(3654) <= not a;
    layer6_outputs(3655) <= not (a xor b);
    layer6_outputs(3656) <= a xor b;
    layer6_outputs(3657) <= not (a or b);
    layer6_outputs(3658) <= not (a xor b);
    layer6_outputs(3659) <= a;
    layer6_outputs(3660) <= b;
    layer6_outputs(3661) <= not a;
    layer6_outputs(3662) <= a and b;
    layer6_outputs(3663) <= not a;
    layer6_outputs(3664) <= not a;
    layer6_outputs(3665) <= not b or a;
    layer6_outputs(3666) <= not a or b;
    layer6_outputs(3667) <= not a;
    layer6_outputs(3668) <= not (a and b);
    layer6_outputs(3669) <= not (a xor b);
    layer6_outputs(3670) <= a xor b;
    layer6_outputs(3671) <= not (a and b);
    layer6_outputs(3672) <= '0';
    layer6_outputs(3673) <= not (a and b);
    layer6_outputs(3674) <= not b or a;
    layer6_outputs(3675) <= not a;
    layer6_outputs(3676) <= not a;
    layer6_outputs(3677) <= not a;
    layer6_outputs(3678) <= a xor b;
    layer6_outputs(3679) <= b and not a;
    layer6_outputs(3680) <= a;
    layer6_outputs(3681) <= not b;
    layer6_outputs(3682) <= a and not b;
    layer6_outputs(3683) <= not b;
    layer6_outputs(3684) <= a and not b;
    layer6_outputs(3685) <= not a;
    layer6_outputs(3686) <= not (a xor b);
    layer6_outputs(3687) <= not (a or b);
    layer6_outputs(3688) <= not b;
    layer6_outputs(3689) <= b;
    layer6_outputs(3690) <= a xor b;
    layer6_outputs(3691) <= a or b;
    layer6_outputs(3692) <= b;
    layer6_outputs(3693) <= a and not b;
    layer6_outputs(3694) <= a or b;
    layer6_outputs(3695) <= b;
    layer6_outputs(3696) <= a xor b;
    layer6_outputs(3697) <= not (a or b);
    layer6_outputs(3698) <= not (a xor b);
    layer6_outputs(3699) <= a;
    layer6_outputs(3700) <= not (a and b);
    layer6_outputs(3701) <= not (a or b);
    layer6_outputs(3702) <= b;
    layer6_outputs(3703) <= not (a or b);
    layer6_outputs(3704) <= a;
    layer6_outputs(3705) <= not a;
    layer6_outputs(3706) <= not (a or b);
    layer6_outputs(3707) <= a and b;
    layer6_outputs(3708) <= not (a xor b);
    layer6_outputs(3709) <= a and not b;
    layer6_outputs(3710) <= not a;
    layer6_outputs(3711) <= not a or b;
    layer6_outputs(3712) <= b;
    layer6_outputs(3713) <= a and not b;
    layer6_outputs(3714) <= a;
    layer6_outputs(3715) <= a;
    layer6_outputs(3716) <= a and b;
    layer6_outputs(3717) <= not b;
    layer6_outputs(3718) <= a;
    layer6_outputs(3719) <= a;
    layer6_outputs(3720) <= b;
    layer6_outputs(3721) <= a xor b;
    layer6_outputs(3722) <= a or b;
    layer6_outputs(3723) <= a xor b;
    layer6_outputs(3724) <= a xor b;
    layer6_outputs(3725) <= a;
    layer6_outputs(3726) <= a and b;
    layer6_outputs(3727) <= not (a xor b);
    layer6_outputs(3728) <= a and b;
    layer6_outputs(3729) <= a or b;
    layer6_outputs(3730) <= not (a xor b);
    layer6_outputs(3731) <= not (a xor b);
    layer6_outputs(3732) <= a and b;
    layer6_outputs(3733) <= a;
    layer6_outputs(3734) <= b;
    layer6_outputs(3735) <= not b;
    layer6_outputs(3736) <= a xor b;
    layer6_outputs(3737) <= a and not b;
    layer6_outputs(3738) <= a;
    layer6_outputs(3739) <= not b or a;
    layer6_outputs(3740) <= not (a or b);
    layer6_outputs(3741) <= not (a xor b);
    layer6_outputs(3742) <= not a;
    layer6_outputs(3743) <= a or b;
    layer6_outputs(3744) <= not a;
    layer6_outputs(3745) <= a or b;
    layer6_outputs(3746) <= a and b;
    layer6_outputs(3747) <= a and not b;
    layer6_outputs(3748) <= not b;
    layer6_outputs(3749) <= not b or a;
    layer6_outputs(3750) <= a;
    layer6_outputs(3751) <= not a or b;
    layer6_outputs(3752) <= a xor b;
    layer6_outputs(3753) <= not a;
    layer6_outputs(3754) <= a;
    layer6_outputs(3755) <= a xor b;
    layer6_outputs(3756) <= not a;
    layer6_outputs(3757) <= b and not a;
    layer6_outputs(3758) <= a xor b;
    layer6_outputs(3759) <= not a;
    layer6_outputs(3760) <= not a;
    layer6_outputs(3761) <= a xor b;
    layer6_outputs(3762) <= b and not a;
    layer6_outputs(3763) <= not b;
    layer6_outputs(3764) <= not (a or b);
    layer6_outputs(3765) <= b and not a;
    layer6_outputs(3766) <= '1';
    layer6_outputs(3767) <= a xor b;
    layer6_outputs(3768) <= not (a xor b);
    layer6_outputs(3769) <= a and not b;
    layer6_outputs(3770) <= not (a and b);
    layer6_outputs(3771) <= not a or b;
    layer6_outputs(3772) <= b;
    layer6_outputs(3773) <= b and not a;
    layer6_outputs(3774) <= b;
    layer6_outputs(3775) <= not a;
    layer6_outputs(3776) <= not (a xor b);
    layer6_outputs(3777) <= a xor b;
    layer6_outputs(3778) <= not (a xor b);
    layer6_outputs(3779) <= not b;
    layer6_outputs(3780) <= a xor b;
    layer6_outputs(3781) <= a and b;
    layer6_outputs(3782) <= not a or b;
    layer6_outputs(3783) <= not a;
    layer6_outputs(3784) <= a;
    layer6_outputs(3785) <= a and not b;
    layer6_outputs(3786) <= not a;
    layer6_outputs(3787) <= not (a and b);
    layer6_outputs(3788) <= b;
    layer6_outputs(3789) <= not (a xor b);
    layer6_outputs(3790) <= not b;
    layer6_outputs(3791) <= not b or a;
    layer6_outputs(3792) <= a and b;
    layer6_outputs(3793) <= not (a and b);
    layer6_outputs(3794) <= not a;
    layer6_outputs(3795) <= b and not a;
    layer6_outputs(3796) <= a and not b;
    layer6_outputs(3797) <= a and b;
    layer6_outputs(3798) <= a;
    layer6_outputs(3799) <= b;
    layer6_outputs(3800) <= '1';
    layer6_outputs(3801) <= not a;
    layer6_outputs(3802) <= not b;
    layer6_outputs(3803) <= b;
    layer6_outputs(3804) <= a or b;
    layer6_outputs(3805) <= a xor b;
    layer6_outputs(3806) <= a xor b;
    layer6_outputs(3807) <= a and not b;
    layer6_outputs(3808) <= b;
    layer6_outputs(3809) <= a;
    layer6_outputs(3810) <= a;
    layer6_outputs(3811) <= not a;
    layer6_outputs(3812) <= not (a and b);
    layer6_outputs(3813) <= a and b;
    layer6_outputs(3814) <= a and b;
    layer6_outputs(3815) <= not a;
    layer6_outputs(3816) <= not b;
    layer6_outputs(3817) <= not (a xor b);
    layer6_outputs(3818) <= b and not a;
    layer6_outputs(3819) <= not a;
    layer6_outputs(3820) <= not a;
    layer6_outputs(3821) <= not a;
    layer6_outputs(3822) <= not (a and b);
    layer6_outputs(3823) <= not a;
    layer6_outputs(3824) <= not a;
    layer6_outputs(3825) <= a;
    layer6_outputs(3826) <= not b;
    layer6_outputs(3827) <= not a or b;
    layer6_outputs(3828) <= not a;
    layer6_outputs(3829) <= b and not a;
    layer6_outputs(3830) <= b and not a;
    layer6_outputs(3831) <= a and b;
    layer6_outputs(3832) <= not a;
    layer6_outputs(3833) <= b;
    layer6_outputs(3834) <= a and not b;
    layer6_outputs(3835) <= a xor b;
    layer6_outputs(3836) <= a xor b;
    layer6_outputs(3837) <= a;
    layer6_outputs(3838) <= not (a or b);
    layer6_outputs(3839) <= not (a or b);
    layer6_outputs(3840) <= a;
    layer6_outputs(3841) <= a xor b;
    layer6_outputs(3842) <= b;
    layer6_outputs(3843) <= not a;
    layer6_outputs(3844) <= not a;
    layer6_outputs(3845) <= b and not a;
    layer6_outputs(3846) <= not a;
    layer6_outputs(3847) <= a xor b;
    layer6_outputs(3848) <= not b;
    layer6_outputs(3849) <= not b;
    layer6_outputs(3850) <= b and not a;
    layer6_outputs(3851) <= a and b;
    layer6_outputs(3852) <= not (a xor b);
    layer6_outputs(3853) <= not (a xor b);
    layer6_outputs(3854) <= b and not a;
    layer6_outputs(3855) <= a;
    layer6_outputs(3856) <= a;
    layer6_outputs(3857) <= not (a and b);
    layer6_outputs(3858) <= a xor b;
    layer6_outputs(3859) <= not (a xor b);
    layer6_outputs(3860) <= not b;
    layer6_outputs(3861) <= not b;
    layer6_outputs(3862) <= a and not b;
    layer6_outputs(3863) <= not (a xor b);
    layer6_outputs(3864) <= a and b;
    layer6_outputs(3865) <= not (a or b);
    layer6_outputs(3866) <= not b or a;
    layer6_outputs(3867) <= b;
    layer6_outputs(3868) <= not (a xor b);
    layer6_outputs(3869) <= not b;
    layer6_outputs(3870) <= b;
    layer6_outputs(3871) <= a xor b;
    layer6_outputs(3872) <= not (a xor b);
    layer6_outputs(3873) <= not b or a;
    layer6_outputs(3874) <= a or b;
    layer6_outputs(3875) <= not a or b;
    layer6_outputs(3876) <= b;
    layer6_outputs(3877) <= a;
    layer6_outputs(3878) <= b;
    layer6_outputs(3879) <= not a;
    layer6_outputs(3880) <= a xor b;
    layer6_outputs(3881) <= b;
    layer6_outputs(3882) <= a xor b;
    layer6_outputs(3883) <= not a;
    layer6_outputs(3884) <= not (a xor b);
    layer6_outputs(3885) <= not (a xor b);
    layer6_outputs(3886) <= not b;
    layer6_outputs(3887) <= a;
    layer6_outputs(3888) <= a;
    layer6_outputs(3889) <= b;
    layer6_outputs(3890) <= a;
    layer6_outputs(3891) <= a;
    layer6_outputs(3892) <= not (a or b);
    layer6_outputs(3893) <= a xor b;
    layer6_outputs(3894) <= a;
    layer6_outputs(3895) <= a and b;
    layer6_outputs(3896) <= not b;
    layer6_outputs(3897) <= a or b;
    layer6_outputs(3898) <= not a;
    layer6_outputs(3899) <= a;
    layer6_outputs(3900) <= not a;
    layer6_outputs(3901) <= not b or a;
    layer6_outputs(3902) <= a or b;
    layer6_outputs(3903) <= not (a xor b);
    layer6_outputs(3904) <= not b or a;
    layer6_outputs(3905) <= not b;
    layer6_outputs(3906) <= a;
    layer6_outputs(3907) <= not a;
    layer6_outputs(3908) <= not (a xor b);
    layer6_outputs(3909) <= b;
    layer6_outputs(3910) <= not b;
    layer6_outputs(3911) <= not a;
    layer6_outputs(3912) <= not b or a;
    layer6_outputs(3913) <= a xor b;
    layer6_outputs(3914) <= not a or b;
    layer6_outputs(3915) <= not a;
    layer6_outputs(3916) <= not b;
    layer6_outputs(3917) <= not a or b;
    layer6_outputs(3918) <= not (a and b);
    layer6_outputs(3919) <= not a;
    layer6_outputs(3920) <= not a;
    layer6_outputs(3921) <= a;
    layer6_outputs(3922) <= not b;
    layer6_outputs(3923) <= not b;
    layer6_outputs(3924) <= a and b;
    layer6_outputs(3925) <= not (a or b);
    layer6_outputs(3926) <= b and not a;
    layer6_outputs(3927) <= not a;
    layer6_outputs(3928) <= a;
    layer6_outputs(3929) <= a xor b;
    layer6_outputs(3930) <= not b;
    layer6_outputs(3931) <= b and not a;
    layer6_outputs(3932) <= a;
    layer6_outputs(3933) <= a;
    layer6_outputs(3934) <= a xor b;
    layer6_outputs(3935) <= not b or a;
    layer6_outputs(3936) <= not a;
    layer6_outputs(3937) <= not a or b;
    layer6_outputs(3938) <= a xor b;
    layer6_outputs(3939) <= not a;
    layer6_outputs(3940) <= b;
    layer6_outputs(3941) <= not b;
    layer6_outputs(3942) <= not a;
    layer6_outputs(3943) <= not (a and b);
    layer6_outputs(3944) <= a;
    layer6_outputs(3945) <= not (a xor b);
    layer6_outputs(3946) <= a or b;
    layer6_outputs(3947) <= not a;
    layer6_outputs(3948) <= b;
    layer6_outputs(3949) <= a xor b;
    layer6_outputs(3950) <= not (a xor b);
    layer6_outputs(3951) <= b;
    layer6_outputs(3952) <= not a;
    layer6_outputs(3953) <= not (a xor b);
    layer6_outputs(3954) <= b;
    layer6_outputs(3955) <= not a;
    layer6_outputs(3956) <= b;
    layer6_outputs(3957) <= a xor b;
    layer6_outputs(3958) <= not a;
    layer6_outputs(3959) <= a and b;
    layer6_outputs(3960) <= not (a xor b);
    layer6_outputs(3961) <= a and not b;
    layer6_outputs(3962) <= a;
    layer6_outputs(3963) <= a xor b;
    layer6_outputs(3964) <= a xor b;
    layer6_outputs(3965) <= b;
    layer6_outputs(3966) <= not a or b;
    layer6_outputs(3967) <= b and not a;
    layer6_outputs(3968) <= not (a xor b);
    layer6_outputs(3969) <= not a;
    layer6_outputs(3970) <= a;
    layer6_outputs(3971) <= a and b;
    layer6_outputs(3972) <= b and not a;
    layer6_outputs(3973) <= not a;
    layer6_outputs(3974) <= not a;
    layer6_outputs(3975) <= a and not b;
    layer6_outputs(3976) <= a and b;
    layer6_outputs(3977) <= not b;
    layer6_outputs(3978) <= not a or b;
    layer6_outputs(3979) <= a or b;
    layer6_outputs(3980) <= a or b;
    layer6_outputs(3981) <= a;
    layer6_outputs(3982) <= not a or b;
    layer6_outputs(3983) <= not b;
    layer6_outputs(3984) <= not b;
    layer6_outputs(3985) <= not a or b;
    layer6_outputs(3986) <= b;
    layer6_outputs(3987) <= not b;
    layer6_outputs(3988) <= not a;
    layer6_outputs(3989) <= b and not a;
    layer6_outputs(3990) <= not b;
    layer6_outputs(3991) <= a;
    layer6_outputs(3992) <= not b or a;
    layer6_outputs(3993) <= not b;
    layer6_outputs(3994) <= not (a or b);
    layer6_outputs(3995) <= not b;
    layer6_outputs(3996) <= not b;
    layer6_outputs(3997) <= not b or a;
    layer6_outputs(3998) <= b;
    layer6_outputs(3999) <= not b or a;
    layer6_outputs(4000) <= not (a xor b);
    layer6_outputs(4001) <= a and b;
    layer6_outputs(4002) <= not a or b;
    layer6_outputs(4003) <= not a;
    layer6_outputs(4004) <= a;
    layer6_outputs(4005) <= not (a and b);
    layer6_outputs(4006) <= not b;
    layer6_outputs(4007) <= not a;
    layer6_outputs(4008) <= not a or b;
    layer6_outputs(4009) <= a and not b;
    layer6_outputs(4010) <= a and b;
    layer6_outputs(4011) <= a and not b;
    layer6_outputs(4012) <= not (a xor b);
    layer6_outputs(4013) <= not (a xor b);
    layer6_outputs(4014) <= not b;
    layer6_outputs(4015) <= a xor b;
    layer6_outputs(4016) <= b;
    layer6_outputs(4017) <= not (a and b);
    layer6_outputs(4018) <= a;
    layer6_outputs(4019) <= not (a xor b);
    layer6_outputs(4020) <= not a;
    layer6_outputs(4021) <= not b;
    layer6_outputs(4022) <= not b or a;
    layer6_outputs(4023) <= a;
    layer6_outputs(4024) <= a xor b;
    layer6_outputs(4025) <= b;
    layer6_outputs(4026) <= a;
    layer6_outputs(4027) <= a xor b;
    layer6_outputs(4028) <= not b or a;
    layer6_outputs(4029) <= a;
    layer6_outputs(4030) <= not b or a;
    layer6_outputs(4031) <= not a;
    layer6_outputs(4032) <= a xor b;
    layer6_outputs(4033) <= a xor b;
    layer6_outputs(4034) <= a and b;
    layer6_outputs(4035) <= not a;
    layer6_outputs(4036) <= a;
    layer6_outputs(4037) <= a or b;
    layer6_outputs(4038) <= '0';
    layer6_outputs(4039) <= not (a or b);
    layer6_outputs(4040) <= not (a xor b);
    layer6_outputs(4041) <= not (a xor b);
    layer6_outputs(4042) <= a;
    layer6_outputs(4043) <= a or b;
    layer6_outputs(4044) <= a xor b;
    layer6_outputs(4045) <= a xor b;
    layer6_outputs(4046) <= a xor b;
    layer6_outputs(4047) <= not (a or b);
    layer6_outputs(4048) <= a or b;
    layer6_outputs(4049) <= a and not b;
    layer6_outputs(4050) <= not b or a;
    layer6_outputs(4051) <= not a;
    layer6_outputs(4052) <= not (a or b);
    layer6_outputs(4053) <= a;
    layer6_outputs(4054) <= not b;
    layer6_outputs(4055) <= a and not b;
    layer6_outputs(4056) <= not a or b;
    layer6_outputs(4057) <= not b;
    layer6_outputs(4058) <= not b;
    layer6_outputs(4059) <= not (a and b);
    layer6_outputs(4060) <= a;
    layer6_outputs(4061) <= a xor b;
    layer6_outputs(4062) <= a xor b;
    layer6_outputs(4063) <= not (a and b);
    layer6_outputs(4064) <= not (a xor b);
    layer6_outputs(4065) <= a;
    layer6_outputs(4066) <= not (a or b);
    layer6_outputs(4067) <= not b;
    layer6_outputs(4068) <= a xor b;
    layer6_outputs(4069) <= a xor b;
    layer6_outputs(4070) <= not a or b;
    layer6_outputs(4071) <= a;
    layer6_outputs(4072) <= a xor b;
    layer6_outputs(4073) <= b;
    layer6_outputs(4074) <= not (a and b);
    layer6_outputs(4075) <= b;
    layer6_outputs(4076) <= not b;
    layer6_outputs(4077) <= b and not a;
    layer6_outputs(4078) <= not b;
    layer6_outputs(4079) <= b;
    layer6_outputs(4080) <= a xor b;
    layer6_outputs(4081) <= b;
    layer6_outputs(4082) <= not a;
    layer6_outputs(4083) <= b;
    layer6_outputs(4084) <= a;
    layer6_outputs(4085) <= a and not b;
    layer6_outputs(4086) <= not b;
    layer6_outputs(4087) <= not (a xor b);
    layer6_outputs(4088) <= not b;
    layer6_outputs(4089) <= not a or b;
    layer6_outputs(4090) <= not a;
    layer6_outputs(4091) <= a;
    layer6_outputs(4092) <= not (a or b);
    layer6_outputs(4093) <= a;
    layer6_outputs(4094) <= not (a or b);
    layer6_outputs(4095) <= not a or b;
    layer6_outputs(4096) <= not (a xor b);
    layer6_outputs(4097) <= not a or b;
    layer6_outputs(4098) <= not b or a;
    layer6_outputs(4099) <= not (a xor b);
    layer6_outputs(4100) <= a xor b;
    layer6_outputs(4101) <= not b;
    layer6_outputs(4102) <= not b;
    layer6_outputs(4103) <= not (a or b);
    layer6_outputs(4104) <= a;
    layer6_outputs(4105) <= not a;
    layer6_outputs(4106) <= a;
    layer6_outputs(4107) <= not a or b;
    layer6_outputs(4108) <= not b or a;
    layer6_outputs(4109) <= a xor b;
    layer6_outputs(4110) <= not b;
    layer6_outputs(4111) <= not (a xor b);
    layer6_outputs(4112) <= not b;
    layer6_outputs(4113) <= not b;
    layer6_outputs(4114) <= not b;
    layer6_outputs(4115) <= not a;
    layer6_outputs(4116) <= not b or a;
    layer6_outputs(4117) <= not (a xor b);
    layer6_outputs(4118) <= not b;
    layer6_outputs(4119) <= not b;
    layer6_outputs(4120) <= not b;
    layer6_outputs(4121) <= not a;
    layer6_outputs(4122) <= not (a xor b);
    layer6_outputs(4123) <= not b;
    layer6_outputs(4124) <= a;
    layer6_outputs(4125) <= b;
    layer6_outputs(4126) <= a xor b;
    layer6_outputs(4127) <= a;
    layer6_outputs(4128) <= not (a xor b);
    layer6_outputs(4129) <= not a;
    layer6_outputs(4130) <= b and not a;
    layer6_outputs(4131) <= b;
    layer6_outputs(4132) <= a;
    layer6_outputs(4133) <= not (a or b);
    layer6_outputs(4134) <= a xor b;
    layer6_outputs(4135) <= not b or a;
    layer6_outputs(4136) <= not b or a;
    layer6_outputs(4137) <= not a;
    layer6_outputs(4138) <= not (a xor b);
    layer6_outputs(4139) <= a xor b;
    layer6_outputs(4140) <= a;
    layer6_outputs(4141) <= not a;
    layer6_outputs(4142) <= not b or a;
    layer6_outputs(4143) <= not b;
    layer6_outputs(4144) <= b and not a;
    layer6_outputs(4145) <= not a;
    layer6_outputs(4146) <= a;
    layer6_outputs(4147) <= not (a and b);
    layer6_outputs(4148) <= not (a xor b);
    layer6_outputs(4149) <= a and not b;
    layer6_outputs(4150) <= not b;
    layer6_outputs(4151) <= not (a xor b);
    layer6_outputs(4152) <= a and not b;
    layer6_outputs(4153) <= not a;
    layer6_outputs(4154) <= b;
    layer6_outputs(4155) <= a xor b;
    layer6_outputs(4156) <= a and b;
    layer6_outputs(4157) <= not a or b;
    layer6_outputs(4158) <= not b;
    layer6_outputs(4159) <= not (a xor b);
    layer6_outputs(4160) <= a;
    layer6_outputs(4161) <= not (a xor b);
    layer6_outputs(4162) <= a xor b;
    layer6_outputs(4163) <= a and not b;
    layer6_outputs(4164) <= a xor b;
    layer6_outputs(4165) <= a or b;
    layer6_outputs(4166) <= not a or b;
    layer6_outputs(4167) <= a;
    layer6_outputs(4168) <= a or b;
    layer6_outputs(4169) <= a and b;
    layer6_outputs(4170) <= not (a xor b);
    layer6_outputs(4171) <= not (a and b);
    layer6_outputs(4172) <= a;
    layer6_outputs(4173) <= a and b;
    layer6_outputs(4174) <= not (a xor b);
    layer6_outputs(4175) <= not (a and b);
    layer6_outputs(4176) <= b and not a;
    layer6_outputs(4177) <= a;
    layer6_outputs(4178) <= not (a xor b);
    layer6_outputs(4179) <= not a or b;
    layer6_outputs(4180) <= a and b;
    layer6_outputs(4181) <= not (a or b);
    layer6_outputs(4182) <= not (a xor b);
    layer6_outputs(4183) <= b;
    layer6_outputs(4184) <= not (a xor b);
    layer6_outputs(4185) <= not (a xor b);
    layer6_outputs(4186) <= not (a and b);
    layer6_outputs(4187) <= not (a xor b);
    layer6_outputs(4188) <= not (a xor b);
    layer6_outputs(4189) <= not b;
    layer6_outputs(4190) <= a and b;
    layer6_outputs(4191) <= not (a xor b);
    layer6_outputs(4192) <= not (a xor b);
    layer6_outputs(4193) <= not (a xor b);
    layer6_outputs(4194) <= a;
    layer6_outputs(4195) <= not b;
    layer6_outputs(4196) <= not (a xor b);
    layer6_outputs(4197) <= b;
    layer6_outputs(4198) <= not b or a;
    layer6_outputs(4199) <= not (a xor b);
    layer6_outputs(4200) <= a xor b;
    layer6_outputs(4201) <= not a or b;
    layer6_outputs(4202) <= a xor b;
    layer6_outputs(4203) <= not b;
    layer6_outputs(4204) <= not b or a;
    layer6_outputs(4205) <= not (a or b);
    layer6_outputs(4206) <= not (a and b);
    layer6_outputs(4207) <= b and not a;
    layer6_outputs(4208) <= b and not a;
    layer6_outputs(4209) <= not (a xor b);
    layer6_outputs(4210) <= not (a and b);
    layer6_outputs(4211) <= not (a and b);
    layer6_outputs(4212) <= a xor b;
    layer6_outputs(4213) <= not b or a;
    layer6_outputs(4214) <= a;
    layer6_outputs(4215) <= b;
    layer6_outputs(4216) <= a;
    layer6_outputs(4217) <= not (a xor b);
    layer6_outputs(4218) <= a;
    layer6_outputs(4219) <= not (a or b);
    layer6_outputs(4220) <= not (a xor b);
    layer6_outputs(4221) <= not (a xor b);
    layer6_outputs(4222) <= not b;
    layer6_outputs(4223) <= a;
    layer6_outputs(4224) <= b and not a;
    layer6_outputs(4225) <= not b;
    layer6_outputs(4226) <= b;
    layer6_outputs(4227) <= b;
    layer6_outputs(4228) <= a or b;
    layer6_outputs(4229) <= not b;
    layer6_outputs(4230) <= not (a and b);
    layer6_outputs(4231) <= a xor b;
    layer6_outputs(4232) <= a;
    layer6_outputs(4233) <= not (a xor b);
    layer6_outputs(4234) <= a xor b;
    layer6_outputs(4235) <= b;
    layer6_outputs(4236) <= a xor b;
    layer6_outputs(4237) <= not (a xor b);
    layer6_outputs(4238) <= a;
    layer6_outputs(4239) <= not (a xor b);
    layer6_outputs(4240) <= not (a xor b);
    layer6_outputs(4241) <= a xor b;
    layer6_outputs(4242) <= not a;
    layer6_outputs(4243) <= a and b;
    layer6_outputs(4244) <= b;
    layer6_outputs(4245) <= a;
    layer6_outputs(4246) <= not a or b;
    layer6_outputs(4247) <= not a or b;
    layer6_outputs(4248) <= a xor b;
    layer6_outputs(4249) <= not (a xor b);
    layer6_outputs(4250) <= not b;
    layer6_outputs(4251) <= not b or a;
    layer6_outputs(4252) <= not a or b;
    layer6_outputs(4253) <= b;
    layer6_outputs(4254) <= not a or b;
    layer6_outputs(4255) <= not (a xor b);
    layer6_outputs(4256) <= a;
    layer6_outputs(4257) <= a or b;
    layer6_outputs(4258) <= a;
    layer6_outputs(4259) <= b;
    layer6_outputs(4260) <= not a;
    layer6_outputs(4261) <= not (a xor b);
    layer6_outputs(4262) <= b and not a;
    layer6_outputs(4263) <= a;
    layer6_outputs(4264) <= b;
    layer6_outputs(4265) <= not b;
    layer6_outputs(4266) <= a and not b;
    layer6_outputs(4267) <= not (a xor b);
    layer6_outputs(4268) <= not a;
    layer6_outputs(4269) <= not (a xor b);
    layer6_outputs(4270) <= a;
    layer6_outputs(4271) <= not (a or b);
    layer6_outputs(4272) <= not a;
    layer6_outputs(4273) <= not b;
    layer6_outputs(4274) <= not (a xor b);
    layer6_outputs(4275) <= a;
    layer6_outputs(4276) <= not (a xor b);
    layer6_outputs(4277) <= not b;
    layer6_outputs(4278) <= b and not a;
    layer6_outputs(4279) <= not (a xor b);
    layer6_outputs(4280) <= a and b;
    layer6_outputs(4281) <= not (a or b);
    layer6_outputs(4282) <= not (a xor b);
    layer6_outputs(4283) <= a xor b;
    layer6_outputs(4284) <= not a or b;
    layer6_outputs(4285) <= not (a xor b);
    layer6_outputs(4286) <= b;
    layer6_outputs(4287) <= a and not b;
    layer6_outputs(4288) <= a and not b;
    layer6_outputs(4289) <= b and not a;
    layer6_outputs(4290) <= a;
    layer6_outputs(4291) <= not (a and b);
    layer6_outputs(4292) <= a;
    layer6_outputs(4293) <= not (a or b);
    layer6_outputs(4294) <= not b or a;
    layer6_outputs(4295) <= a;
    layer6_outputs(4296) <= a;
    layer6_outputs(4297) <= a xor b;
    layer6_outputs(4298) <= a;
    layer6_outputs(4299) <= a and b;
    layer6_outputs(4300) <= not a;
    layer6_outputs(4301) <= not a;
    layer6_outputs(4302) <= not a;
    layer6_outputs(4303) <= '1';
    layer6_outputs(4304) <= not a;
    layer6_outputs(4305) <= not b;
    layer6_outputs(4306) <= a xor b;
    layer6_outputs(4307) <= a xor b;
    layer6_outputs(4308) <= not b;
    layer6_outputs(4309) <= a;
    layer6_outputs(4310) <= not (a xor b);
    layer6_outputs(4311) <= not a;
    layer6_outputs(4312) <= not a;
    layer6_outputs(4313) <= not a;
    layer6_outputs(4314) <= not a;
    layer6_outputs(4315) <= b;
    layer6_outputs(4316) <= a;
    layer6_outputs(4317) <= a and not b;
    layer6_outputs(4318) <= not (a xor b);
    layer6_outputs(4319) <= not (a xor b);
    layer6_outputs(4320) <= not (a and b);
    layer6_outputs(4321) <= a;
    layer6_outputs(4322) <= not (a and b);
    layer6_outputs(4323) <= b;
    layer6_outputs(4324) <= not b;
    layer6_outputs(4325) <= a;
    layer6_outputs(4326) <= a;
    layer6_outputs(4327) <= a;
    layer6_outputs(4328) <= a xor b;
    layer6_outputs(4329) <= a;
    layer6_outputs(4330) <= b;
    layer6_outputs(4331) <= not a;
    layer6_outputs(4332) <= not b;
    layer6_outputs(4333) <= not b or a;
    layer6_outputs(4334) <= not (a or b);
    layer6_outputs(4335) <= a;
    layer6_outputs(4336) <= not (a xor b);
    layer6_outputs(4337) <= not (a and b);
    layer6_outputs(4338) <= a or b;
    layer6_outputs(4339) <= not (a and b);
    layer6_outputs(4340) <= a;
    layer6_outputs(4341) <= not (a xor b);
    layer6_outputs(4342) <= not a;
    layer6_outputs(4343) <= a;
    layer6_outputs(4344) <= b;
    layer6_outputs(4345) <= not b;
    layer6_outputs(4346) <= not (a xor b);
    layer6_outputs(4347) <= a xor b;
    layer6_outputs(4348) <= a or b;
    layer6_outputs(4349) <= not a;
    layer6_outputs(4350) <= not (a or b);
    layer6_outputs(4351) <= a;
    layer6_outputs(4352) <= not (a xor b);
    layer6_outputs(4353) <= not b;
    layer6_outputs(4354) <= not b;
    layer6_outputs(4355) <= not b;
    layer6_outputs(4356) <= a and b;
    layer6_outputs(4357) <= not (a xor b);
    layer6_outputs(4358) <= a or b;
    layer6_outputs(4359) <= not a;
    layer6_outputs(4360) <= not (a and b);
    layer6_outputs(4361) <= not b;
    layer6_outputs(4362) <= not (a xor b);
    layer6_outputs(4363) <= b;
    layer6_outputs(4364) <= a;
    layer6_outputs(4365) <= not (a and b);
    layer6_outputs(4366) <= not (a or b);
    layer6_outputs(4367) <= b and not a;
    layer6_outputs(4368) <= not b;
    layer6_outputs(4369) <= b;
    layer6_outputs(4370) <= not (a or b);
    layer6_outputs(4371) <= b and not a;
    layer6_outputs(4372) <= not (a xor b);
    layer6_outputs(4373) <= not b;
    layer6_outputs(4374) <= a xor b;
    layer6_outputs(4375) <= a xor b;
    layer6_outputs(4376) <= a;
    layer6_outputs(4377) <= not (a or b);
    layer6_outputs(4378) <= a;
    layer6_outputs(4379) <= not (a xor b);
    layer6_outputs(4380) <= b and not a;
    layer6_outputs(4381) <= a;
    layer6_outputs(4382) <= a and b;
    layer6_outputs(4383) <= not b;
    layer6_outputs(4384) <= not b;
    layer6_outputs(4385) <= not a;
    layer6_outputs(4386) <= not (a and b);
    layer6_outputs(4387) <= not (a and b);
    layer6_outputs(4388) <= a or b;
    layer6_outputs(4389) <= not (a or b);
    layer6_outputs(4390) <= a and b;
    layer6_outputs(4391) <= b and not a;
    layer6_outputs(4392) <= not a;
    layer6_outputs(4393) <= a or b;
    layer6_outputs(4394) <= b;
    layer6_outputs(4395) <= not a;
    layer6_outputs(4396) <= a or b;
    layer6_outputs(4397) <= a xor b;
    layer6_outputs(4398) <= not (a xor b);
    layer6_outputs(4399) <= a;
    layer6_outputs(4400) <= a xor b;
    layer6_outputs(4401) <= a;
    layer6_outputs(4402) <= a xor b;
    layer6_outputs(4403) <= not (a and b);
    layer6_outputs(4404) <= not (a and b);
    layer6_outputs(4405) <= a;
    layer6_outputs(4406) <= not a;
    layer6_outputs(4407) <= not b;
    layer6_outputs(4408) <= not (a or b);
    layer6_outputs(4409) <= not (a and b);
    layer6_outputs(4410) <= b;
    layer6_outputs(4411) <= b and not a;
    layer6_outputs(4412) <= not a;
    layer6_outputs(4413) <= not (a and b);
    layer6_outputs(4414) <= a;
    layer6_outputs(4415) <= not (a and b);
    layer6_outputs(4416) <= b;
    layer6_outputs(4417) <= not b;
    layer6_outputs(4418) <= not a;
    layer6_outputs(4419) <= not b or a;
    layer6_outputs(4420) <= a and b;
    layer6_outputs(4421) <= not a;
    layer6_outputs(4422) <= not a;
    layer6_outputs(4423) <= a;
    layer6_outputs(4424) <= not b;
    layer6_outputs(4425) <= b and not a;
    layer6_outputs(4426) <= not (a xor b);
    layer6_outputs(4427) <= b;
    layer6_outputs(4428) <= b and not a;
    layer6_outputs(4429) <= not b;
    layer6_outputs(4430) <= not b;
    layer6_outputs(4431) <= b;
    layer6_outputs(4432) <= a xor b;
    layer6_outputs(4433) <= a and b;
    layer6_outputs(4434) <= not (a xor b);
    layer6_outputs(4435) <= a and not b;
    layer6_outputs(4436) <= a;
    layer6_outputs(4437) <= not (a xor b);
    layer6_outputs(4438) <= not b or a;
    layer6_outputs(4439) <= a;
    layer6_outputs(4440) <= a;
    layer6_outputs(4441) <= not b;
    layer6_outputs(4442) <= not a;
    layer6_outputs(4443) <= a;
    layer6_outputs(4444) <= a or b;
    layer6_outputs(4445) <= b;
    layer6_outputs(4446) <= not b;
    layer6_outputs(4447) <= a and b;
    layer6_outputs(4448) <= not b;
    layer6_outputs(4449) <= not (a xor b);
    layer6_outputs(4450) <= not (a xor b);
    layer6_outputs(4451) <= a and b;
    layer6_outputs(4452) <= a or b;
    layer6_outputs(4453) <= a or b;
    layer6_outputs(4454) <= not (a xor b);
    layer6_outputs(4455) <= not a or b;
    layer6_outputs(4456) <= not a or b;
    layer6_outputs(4457) <= not b;
    layer6_outputs(4458) <= a xor b;
    layer6_outputs(4459) <= b;
    layer6_outputs(4460) <= not a;
    layer6_outputs(4461) <= a xor b;
    layer6_outputs(4462) <= a xor b;
    layer6_outputs(4463) <= not b;
    layer6_outputs(4464) <= not b or a;
    layer6_outputs(4465) <= b and not a;
    layer6_outputs(4466) <= not a or b;
    layer6_outputs(4467) <= not a;
    layer6_outputs(4468) <= a;
    layer6_outputs(4469) <= not a;
    layer6_outputs(4470) <= b;
    layer6_outputs(4471) <= a xor b;
    layer6_outputs(4472) <= b;
    layer6_outputs(4473) <= a xor b;
    layer6_outputs(4474) <= a xor b;
    layer6_outputs(4475) <= a xor b;
    layer6_outputs(4476) <= not a;
    layer6_outputs(4477) <= not (a xor b);
    layer6_outputs(4478) <= b;
    layer6_outputs(4479) <= not (a xor b);
    layer6_outputs(4480) <= a xor b;
    layer6_outputs(4481) <= not (a xor b);
    layer6_outputs(4482) <= not a or b;
    layer6_outputs(4483) <= not a;
    layer6_outputs(4484) <= not (a and b);
    layer6_outputs(4485) <= not b or a;
    layer6_outputs(4486) <= not (a or b);
    layer6_outputs(4487) <= a;
    layer6_outputs(4488) <= not (a or b);
    layer6_outputs(4489) <= b;
    layer6_outputs(4490) <= not (a or b);
    layer6_outputs(4491) <= not b;
    layer6_outputs(4492) <= b;
    layer6_outputs(4493) <= a;
    layer6_outputs(4494) <= a;
    layer6_outputs(4495) <= not b;
    layer6_outputs(4496) <= not b;
    layer6_outputs(4497) <= a;
    layer6_outputs(4498) <= a and b;
    layer6_outputs(4499) <= a or b;
    layer6_outputs(4500) <= not b or a;
    layer6_outputs(4501) <= not (a xor b);
    layer6_outputs(4502) <= b;
    layer6_outputs(4503) <= a and b;
    layer6_outputs(4504) <= a xor b;
    layer6_outputs(4505) <= not a;
    layer6_outputs(4506) <= not a or b;
    layer6_outputs(4507) <= a;
    layer6_outputs(4508) <= not b or a;
    layer6_outputs(4509) <= a;
    layer6_outputs(4510) <= not (a and b);
    layer6_outputs(4511) <= not a;
    layer6_outputs(4512) <= a;
    layer6_outputs(4513) <= not (a xor b);
    layer6_outputs(4514) <= a or b;
    layer6_outputs(4515) <= a;
    layer6_outputs(4516) <= a;
    layer6_outputs(4517) <= not b;
    layer6_outputs(4518) <= not (a and b);
    layer6_outputs(4519) <= not a or b;
    layer6_outputs(4520) <= a xor b;
    layer6_outputs(4521) <= a and not b;
    layer6_outputs(4522) <= not b;
    layer6_outputs(4523) <= not a;
    layer6_outputs(4524) <= b;
    layer6_outputs(4525) <= a;
    layer6_outputs(4526) <= not (a and b);
    layer6_outputs(4527) <= a;
    layer6_outputs(4528) <= not a or b;
    layer6_outputs(4529) <= not b;
    layer6_outputs(4530) <= b;
    layer6_outputs(4531) <= a or b;
    layer6_outputs(4532) <= not (a xor b);
    layer6_outputs(4533) <= not (a or b);
    layer6_outputs(4534) <= not (a xor b);
    layer6_outputs(4535) <= a and b;
    layer6_outputs(4536) <= b;
    layer6_outputs(4537) <= a;
    layer6_outputs(4538) <= b;
    layer6_outputs(4539) <= not b;
    layer6_outputs(4540) <= a or b;
    layer6_outputs(4541) <= a or b;
    layer6_outputs(4542) <= not (a xor b);
    layer6_outputs(4543) <= a and b;
    layer6_outputs(4544) <= b;
    layer6_outputs(4545) <= b;
    layer6_outputs(4546) <= a;
    layer6_outputs(4547) <= not (a xor b);
    layer6_outputs(4548) <= a;
    layer6_outputs(4549) <= b and not a;
    layer6_outputs(4550) <= not a or b;
    layer6_outputs(4551) <= not (a and b);
    layer6_outputs(4552) <= a xor b;
    layer6_outputs(4553) <= not a;
    layer6_outputs(4554) <= b and not a;
    layer6_outputs(4555) <= a xor b;
    layer6_outputs(4556) <= not a;
    layer6_outputs(4557) <= a or b;
    layer6_outputs(4558) <= not b;
    layer6_outputs(4559) <= a;
    layer6_outputs(4560) <= b;
    layer6_outputs(4561) <= a;
    layer6_outputs(4562) <= not b;
    layer6_outputs(4563) <= a and not b;
    layer6_outputs(4564) <= not b;
    layer6_outputs(4565) <= not a;
    layer6_outputs(4566) <= not (a xor b);
    layer6_outputs(4567) <= not a or b;
    layer6_outputs(4568) <= not b;
    layer6_outputs(4569) <= not b;
    layer6_outputs(4570) <= not a;
    layer6_outputs(4571) <= a xor b;
    layer6_outputs(4572) <= not a;
    layer6_outputs(4573) <= b and not a;
    layer6_outputs(4574) <= a xor b;
    layer6_outputs(4575) <= not a;
    layer6_outputs(4576) <= not a;
    layer6_outputs(4577) <= a or b;
    layer6_outputs(4578) <= not (a or b);
    layer6_outputs(4579) <= a and not b;
    layer6_outputs(4580) <= a and b;
    layer6_outputs(4581) <= not (a xor b);
    layer6_outputs(4582) <= not b;
    layer6_outputs(4583) <= a or b;
    layer6_outputs(4584) <= not a;
    layer6_outputs(4585) <= not (a xor b);
    layer6_outputs(4586) <= not a;
    layer6_outputs(4587) <= not a or b;
    layer6_outputs(4588) <= a xor b;
    layer6_outputs(4589) <= not b;
    layer6_outputs(4590) <= a or b;
    layer6_outputs(4591) <= a and b;
    layer6_outputs(4592) <= a;
    layer6_outputs(4593) <= a xor b;
    layer6_outputs(4594) <= not b;
    layer6_outputs(4595) <= a xor b;
    layer6_outputs(4596) <= a;
    layer6_outputs(4597) <= a;
    layer6_outputs(4598) <= b;
    layer6_outputs(4599) <= not a;
    layer6_outputs(4600) <= b and not a;
    layer6_outputs(4601) <= not a;
    layer6_outputs(4602) <= not b or a;
    layer6_outputs(4603) <= a or b;
    layer6_outputs(4604) <= a xor b;
    layer6_outputs(4605) <= not (a xor b);
    layer6_outputs(4606) <= a and not b;
    layer6_outputs(4607) <= not (a xor b);
    layer6_outputs(4608) <= a and not b;
    layer6_outputs(4609) <= a xor b;
    layer6_outputs(4610) <= a xor b;
    layer6_outputs(4611) <= a and b;
    layer6_outputs(4612) <= b;
    layer6_outputs(4613) <= b;
    layer6_outputs(4614) <= b;
    layer6_outputs(4615) <= not a;
    layer6_outputs(4616) <= a;
    layer6_outputs(4617) <= not (a or b);
    layer6_outputs(4618) <= a;
    layer6_outputs(4619) <= a or b;
    layer6_outputs(4620) <= a;
    layer6_outputs(4621) <= not a or b;
    layer6_outputs(4622) <= a and b;
    layer6_outputs(4623) <= not b;
    layer6_outputs(4624) <= a xor b;
    layer6_outputs(4625) <= a and b;
    layer6_outputs(4626) <= not (a xor b);
    layer6_outputs(4627) <= not b or a;
    layer6_outputs(4628) <= not a;
    layer6_outputs(4629) <= a;
    layer6_outputs(4630) <= not (a or b);
    layer6_outputs(4631) <= not b;
    layer6_outputs(4632) <= not b;
    layer6_outputs(4633) <= b;
    layer6_outputs(4634) <= not (a xor b);
    layer6_outputs(4635) <= a xor b;
    layer6_outputs(4636) <= a and not b;
    layer6_outputs(4637) <= not b or a;
    layer6_outputs(4638) <= not a;
    layer6_outputs(4639) <= not (a xor b);
    layer6_outputs(4640) <= not a or b;
    layer6_outputs(4641) <= not (a xor b);
    layer6_outputs(4642) <= a xor b;
    layer6_outputs(4643) <= not b or a;
    layer6_outputs(4644) <= not a;
    layer6_outputs(4645) <= not (a and b);
    layer6_outputs(4646) <= a xor b;
    layer6_outputs(4647) <= not a or b;
    layer6_outputs(4648) <= a xor b;
    layer6_outputs(4649) <= a xor b;
    layer6_outputs(4650) <= a xor b;
    layer6_outputs(4651) <= a xor b;
    layer6_outputs(4652) <= a and b;
    layer6_outputs(4653) <= a;
    layer6_outputs(4654) <= a xor b;
    layer6_outputs(4655) <= not b;
    layer6_outputs(4656) <= a;
    layer6_outputs(4657) <= not (a xor b);
    layer6_outputs(4658) <= not (a xor b);
    layer6_outputs(4659) <= a;
    layer6_outputs(4660) <= b;
    layer6_outputs(4661) <= b;
    layer6_outputs(4662) <= a and not b;
    layer6_outputs(4663) <= not b;
    layer6_outputs(4664) <= b;
    layer6_outputs(4665) <= a xor b;
    layer6_outputs(4666) <= b;
    layer6_outputs(4667) <= not (a or b);
    layer6_outputs(4668) <= a xor b;
    layer6_outputs(4669) <= b;
    layer6_outputs(4670) <= a or b;
    layer6_outputs(4671) <= not a;
    layer6_outputs(4672) <= b;
    layer6_outputs(4673) <= not a;
    layer6_outputs(4674) <= a xor b;
    layer6_outputs(4675) <= not b or a;
    layer6_outputs(4676) <= not b;
    layer6_outputs(4677) <= not a or b;
    layer6_outputs(4678) <= a or b;
    layer6_outputs(4679) <= not a or b;
    layer6_outputs(4680) <= a or b;
    layer6_outputs(4681) <= not (a xor b);
    layer6_outputs(4682) <= a;
    layer6_outputs(4683) <= b;
    layer6_outputs(4684) <= a;
    layer6_outputs(4685) <= b;
    layer6_outputs(4686) <= b and not a;
    layer6_outputs(4687) <= a;
    layer6_outputs(4688) <= not a;
    layer6_outputs(4689) <= b and not a;
    layer6_outputs(4690) <= b;
    layer6_outputs(4691) <= b;
    layer6_outputs(4692) <= b and not a;
    layer6_outputs(4693) <= not b;
    layer6_outputs(4694) <= a;
    layer6_outputs(4695) <= not b;
    layer6_outputs(4696) <= not a;
    layer6_outputs(4697) <= not (a xor b);
    layer6_outputs(4698) <= not a;
    layer6_outputs(4699) <= a or b;
    layer6_outputs(4700) <= not a;
    layer6_outputs(4701) <= not a;
    layer6_outputs(4702) <= a or b;
    layer6_outputs(4703) <= not b;
    layer6_outputs(4704) <= b and not a;
    layer6_outputs(4705) <= not a;
    layer6_outputs(4706) <= b;
    layer6_outputs(4707) <= not b;
    layer6_outputs(4708) <= a xor b;
    layer6_outputs(4709) <= not a;
    layer6_outputs(4710) <= not b;
    layer6_outputs(4711) <= a;
    layer6_outputs(4712) <= a;
    layer6_outputs(4713) <= not (a xor b);
    layer6_outputs(4714) <= a xor b;
    layer6_outputs(4715) <= not b or a;
    layer6_outputs(4716) <= not (a or b);
    layer6_outputs(4717) <= not a;
    layer6_outputs(4718) <= not a or b;
    layer6_outputs(4719) <= a xor b;
    layer6_outputs(4720) <= not (a and b);
    layer6_outputs(4721) <= not b or a;
    layer6_outputs(4722) <= a;
    layer6_outputs(4723) <= b;
    layer6_outputs(4724) <= not b or a;
    layer6_outputs(4725) <= not (a or b);
    layer6_outputs(4726) <= not (a xor b);
    layer6_outputs(4727) <= not b;
    layer6_outputs(4728) <= not (a and b);
    layer6_outputs(4729) <= not (a xor b);
    layer6_outputs(4730) <= not a or b;
    layer6_outputs(4731) <= not b;
    layer6_outputs(4732) <= b;
    layer6_outputs(4733) <= not (a or b);
    layer6_outputs(4734) <= not b;
    layer6_outputs(4735) <= not (a and b);
    layer6_outputs(4736) <= not a;
    layer6_outputs(4737) <= not a or b;
    layer6_outputs(4738) <= b and not a;
    layer6_outputs(4739) <= not (a xor b);
    layer6_outputs(4740) <= not b or a;
    layer6_outputs(4741) <= a;
    layer6_outputs(4742) <= a and not b;
    layer6_outputs(4743) <= not a or b;
    layer6_outputs(4744) <= not b;
    layer6_outputs(4745) <= not a;
    layer6_outputs(4746) <= not (a xor b);
    layer6_outputs(4747) <= a;
    layer6_outputs(4748) <= a or b;
    layer6_outputs(4749) <= not (a and b);
    layer6_outputs(4750) <= not (a or b);
    layer6_outputs(4751) <= not a;
    layer6_outputs(4752) <= a or b;
    layer6_outputs(4753) <= a xor b;
    layer6_outputs(4754) <= not a;
    layer6_outputs(4755) <= not b;
    layer6_outputs(4756) <= a;
    layer6_outputs(4757) <= not b;
    layer6_outputs(4758) <= not a;
    layer6_outputs(4759) <= not (a xor b);
    layer6_outputs(4760) <= a xor b;
    layer6_outputs(4761) <= not a or b;
    layer6_outputs(4762) <= a xor b;
    layer6_outputs(4763) <= a xor b;
    layer6_outputs(4764) <= a xor b;
    layer6_outputs(4765) <= a xor b;
    layer6_outputs(4766) <= a xor b;
    layer6_outputs(4767) <= b;
    layer6_outputs(4768) <= a;
    layer6_outputs(4769) <= a and b;
    layer6_outputs(4770) <= b;
    layer6_outputs(4771) <= not b;
    layer6_outputs(4772) <= not (a xor b);
    layer6_outputs(4773) <= not b;
    layer6_outputs(4774) <= a and b;
    layer6_outputs(4775) <= not a or b;
    layer6_outputs(4776) <= not b or a;
    layer6_outputs(4777) <= not (a xor b);
    layer6_outputs(4778) <= a;
    layer6_outputs(4779) <= not b;
    layer6_outputs(4780) <= not a or b;
    layer6_outputs(4781) <= a or b;
    layer6_outputs(4782) <= a;
    layer6_outputs(4783) <= not a;
    layer6_outputs(4784) <= a;
    layer6_outputs(4785) <= a xor b;
    layer6_outputs(4786) <= not (a xor b);
    layer6_outputs(4787) <= not a;
    layer6_outputs(4788) <= a;
    layer6_outputs(4789) <= not (a or b);
    layer6_outputs(4790) <= not b;
    layer6_outputs(4791) <= a or b;
    layer6_outputs(4792) <= a;
    layer6_outputs(4793) <= a and not b;
    layer6_outputs(4794) <= not b;
    layer6_outputs(4795) <= b;
    layer6_outputs(4796) <= a and not b;
    layer6_outputs(4797) <= a xor b;
    layer6_outputs(4798) <= not (a or b);
    layer6_outputs(4799) <= a or b;
    layer6_outputs(4800) <= a and not b;
    layer6_outputs(4801) <= a or b;
    layer6_outputs(4802) <= not (a or b);
    layer6_outputs(4803) <= b;
    layer6_outputs(4804) <= not a;
    layer6_outputs(4805) <= not (a or b);
    layer6_outputs(4806) <= not b;
    layer6_outputs(4807) <= not (a or b);
    layer6_outputs(4808) <= a or b;
    layer6_outputs(4809) <= not a;
    layer6_outputs(4810) <= a;
    layer6_outputs(4811) <= not b;
    layer6_outputs(4812) <= not b or a;
    layer6_outputs(4813) <= b;
    layer6_outputs(4814) <= not a;
    layer6_outputs(4815) <= not (a xor b);
    layer6_outputs(4816) <= not (a xor b);
    layer6_outputs(4817) <= not b;
    layer6_outputs(4818) <= not b;
    layer6_outputs(4819) <= a;
    layer6_outputs(4820) <= a or b;
    layer6_outputs(4821) <= not a;
    layer6_outputs(4822) <= not (a xor b);
    layer6_outputs(4823) <= a and not b;
    layer6_outputs(4824) <= not a;
    layer6_outputs(4825) <= b;
    layer6_outputs(4826) <= not b;
    layer6_outputs(4827) <= not (a or b);
    layer6_outputs(4828) <= b and not a;
    layer6_outputs(4829) <= a and b;
    layer6_outputs(4830) <= a xor b;
    layer6_outputs(4831) <= not a or b;
    layer6_outputs(4832) <= not (a xor b);
    layer6_outputs(4833) <= not (a xor b);
    layer6_outputs(4834) <= not a;
    layer6_outputs(4835) <= not b;
    layer6_outputs(4836) <= b and not a;
    layer6_outputs(4837) <= not b;
    layer6_outputs(4838) <= a;
    layer6_outputs(4839) <= a and b;
    layer6_outputs(4840) <= a and not b;
    layer6_outputs(4841) <= not b or a;
    layer6_outputs(4842) <= a xor b;
    layer6_outputs(4843) <= not (a and b);
    layer6_outputs(4844) <= a;
    layer6_outputs(4845) <= a or b;
    layer6_outputs(4846) <= a and not b;
    layer6_outputs(4847) <= not b;
    layer6_outputs(4848) <= not b;
    layer6_outputs(4849) <= a or b;
    layer6_outputs(4850) <= a xor b;
    layer6_outputs(4851) <= not b;
    layer6_outputs(4852) <= not (a xor b);
    layer6_outputs(4853) <= a and not b;
    layer6_outputs(4854) <= not (a xor b);
    layer6_outputs(4855) <= a and not b;
    layer6_outputs(4856) <= not (a or b);
    layer6_outputs(4857) <= a or b;
    layer6_outputs(4858) <= not b;
    layer6_outputs(4859) <= b;
    layer6_outputs(4860) <= a xor b;
    layer6_outputs(4861) <= not a;
    layer6_outputs(4862) <= a xor b;
    layer6_outputs(4863) <= not b or a;
    layer6_outputs(4864) <= a xor b;
    layer6_outputs(4865) <= a or b;
    layer6_outputs(4866) <= not (a xor b);
    layer6_outputs(4867) <= not (a xor b);
    layer6_outputs(4868) <= not b;
    layer6_outputs(4869) <= b and not a;
    layer6_outputs(4870) <= not a or b;
    layer6_outputs(4871) <= b;
    layer6_outputs(4872) <= a;
    layer6_outputs(4873) <= not a;
    layer6_outputs(4874) <= a;
    layer6_outputs(4875) <= not (a xor b);
    layer6_outputs(4876) <= b and not a;
    layer6_outputs(4877) <= a;
    layer6_outputs(4878) <= a xor b;
    layer6_outputs(4879) <= a xor b;
    layer6_outputs(4880) <= a or b;
    layer6_outputs(4881) <= not (a xor b);
    layer6_outputs(4882) <= not b or a;
    layer6_outputs(4883) <= not (a or b);
    layer6_outputs(4884) <= b;
    layer6_outputs(4885) <= not a;
    layer6_outputs(4886) <= not b;
    layer6_outputs(4887) <= b;
    layer6_outputs(4888) <= b;
    layer6_outputs(4889) <= b and not a;
    layer6_outputs(4890) <= not (a and b);
    layer6_outputs(4891) <= not a or b;
    layer6_outputs(4892) <= not (a and b);
    layer6_outputs(4893) <= a xor b;
    layer6_outputs(4894) <= a;
    layer6_outputs(4895) <= not b;
    layer6_outputs(4896) <= not a;
    layer6_outputs(4897) <= a;
    layer6_outputs(4898) <= b;
    layer6_outputs(4899) <= a and not b;
    layer6_outputs(4900) <= a;
    layer6_outputs(4901) <= a xor b;
    layer6_outputs(4902) <= not a;
    layer6_outputs(4903) <= a;
    layer6_outputs(4904) <= not a;
    layer6_outputs(4905) <= a xor b;
    layer6_outputs(4906) <= a;
    layer6_outputs(4907) <= not b or a;
    layer6_outputs(4908) <= not b or a;
    layer6_outputs(4909) <= not (a and b);
    layer6_outputs(4910) <= not a;
    layer6_outputs(4911) <= a;
    layer6_outputs(4912) <= not (a or b);
    layer6_outputs(4913) <= not a;
    layer6_outputs(4914) <= a or b;
    layer6_outputs(4915) <= not a or b;
    layer6_outputs(4916) <= not b;
    layer6_outputs(4917) <= not (a and b);
    layer6_outputs(4918) <= a and not b;
    layer6_outputs(4919) <= a or b;
    layer6_outputs(4920) <= b;
    layer6_outputs(4921) <= not b or a;
    layer6_outputs(4922) <= a;
    layer6_outputs(4923) <= a xor b;
    layer6_outputs(4924) <= a or b;
    layer6_outputs(4925) <= not a;
    layer6_outputs(4926) <= not (a xor b);
    layer6_outputs(4927) <= b and not a;
    layer6_outputs(4928) <= not (a xor b);
    layer6_outputs(4929) <= a;
    layer6_outputs(4930) <= not b;
    layer6_outputs(4931) <= a xor b;
    layer6_outputs(4932) <= not a or b;
    layer6_outputs(4933) <= not b;
    layer6_outputs(4934) <= not (a xor b);
    layer6_outputs(4935) <= not (a or b);
    layer6_outputs(4936) <= not b;
    layer6_outputs(4937) <= b;
    layer6_outputs(4938) <= a xor b;
    layer6_outputs(4939) <= not b or a;
    layer6_outputs(4940) <= a;
    layer6_outputs(4941) <= a and b;
    layer6_outputs(4942) <= not (a xor b);
    layer6_outputs(4943) <= b;
    layer6_outputs(4944) <= not b or a;
    layer6_outputs(4945) <= not b;
    layer6_outputs(4946) <= b;
    layer6_outputs(4947) <= b;
    layer6_outputs(4948) <= b;
    layer6_outputs(4949) <= not a;
    layer6_outputs(4950) <= not b;
    layer6_outputs(4951) <= b;
    layer6_outputs(4952) <= not (a and b);
    layer6_outputs(4953) <= not a;
    layer6_outputs(4954) <= a;
    layer6_outputs(4955) <= not (a xor b);
    layer6_outputs(4956) <= not (a xor b);
    layer6_outputs(4957) <= not b;
    layer6_outputs(4958) <= a xor b;
    layer6_outputs(4959) <= not (a xor b);
    layer6_outputs(4960) <= not (a xor b);
    layer6_outputs(4961) <= a or b;
    layer6_outputs(4962) <= a and not b;
    layer6_outputs(4963) <= b;
    layer6_outputs(4964) <= a and not b;
    layer6_outputs(4965) <= a;
    layer6_outputs(4966) <= a xor b;
    layer6_outputs(4967) <= not b or a;
    layer6_outputs(4968) <= a and b;
    layer6_outputs(4969) <= b;
    layer6_outputs(4970) <= a xor b;
    layer6_outputs(4971) <= a;
    layer6_outputs(4972) <= not (a or b);
    layer6_outputs(4973) <= a xor b;
    layer6_outputs(4974) <= a xor b;
    layer6_outputs(4975) <= not a;
    layer6_outputs(4976) <= not a;
    layer6_outputs(4977) <= a xor b;
    layer6_outputs(4978) <= b;
    layer6_outputs(4979) <= a xor b;
    layer6_outputs(4980) <= a and not b;
    layer6_outputs(4981) <= b;
    layer6_outputs(4982) <= not (a or b);
    layer6_outputs(4983) <= a and not b;
    layer6_outputs(4984) <= b;
    layer6_outputs(4985) <= a xor b;
    layer6_outputs(4986) <= a and b;
    layer6_outputs(4987) <= not b;
    layer6_outputs(4988) <= a and not b;
    layer6_outputs(4989) <= not (a or b);
    layer6_outputs(4990) <= b and not a;
    layer6_outputs(4991) <= b;
    layer6_outputs(4992) <= a and not b;
    layer6_outputs(4993) <= not (a xor b);
    layer6_outputs(4994) <= not b or a;
    layer6_outputs(4995) <= not b or a;
    layer6_outputs(4996) <= not b;
    layer6_outputs(4997) <= b;
    layer6_outputs(4998) <= a;
    layer6_outputs(4999) <= not a or b;
    layer6_outputs(5000) <= b;
    layer6_outputs(5001) <= not b;
    layer6_outputs(5002) <= not a;
    layer6_outputs(5003) <= not (a or b);
    layer6_outputs(5004) <= a xor b;
    layer6_outputs(5005) <= not (a xor b);
    layer6_outputs(5006) <= not b;
    layer6_outputs(5007) <= not (a xor b);
    layer6_outputs(5008) <= not a;
    layer6_outputs(5009) <= not a;
    layer6_outputs(5010) <= a;
    layer6_outputs(5011) <= not (a and b);
    layer6_outputs(5012) <= b;
    layer6_outputs(5013) <= not (a or b);
    layer6_outputs(5014) <= not a;
    layer6_outputs(5015) <= a;
    layer6_outputs(5016) <= not (a and b);
    layer6_outputs(5017) <= not a;
    layer6_outputs(5018) <= a;
    layer6_outputs(5019) <= a;
    layer6_outputs(5020) <= b;
    layer6_outputs(5021) <= not a;
    layer6_outputs(5022) <= not a;
    layer6_outputs(5023) <= not (a xor b);
    layer6_outputs(5024) <= a xor b;
    layer6_outputs(5025) <= a or b;
    layer6_outputs(5026) <= b and not a;
    layer6_outputs(5027) <= not (a xor b);
    layer6_outputs(5028) <= not a or b;
    layer6_outputs(5029) <= a;
    layer6_outputs(5030) <= not a;
    layer6_outputs(5031) <= b;
    layer6_outputs(5032) <= not a;
    layer6_outputs(5033) <= not (a and b);
    layer6_outputs(5034) <= not (a or b);
    layer6_outputs(5035) <= not (a xor b);
    layer6_outputs(5036) <= b;
    layer6_outputs(5037) <= not (a xor b);
    layer6_outputs(5038) <= not (a or b);
    layer6_outputs(5039) <= b;
    layer6_outputs(5040) <= not b;
    layer6_outputs(5041) <= not b;
    layer6_outputs(5042) <= not a or b;
    layer6_outputs(5043) <= b;
    layer6_outputs(5044) <= a xor b;
    layer6_outputs(5045) <= b;
    layer6_outputs(5046) <= not a;
    layer6_outputs(5047) <= a;
    layer6_outputs(5048) <= not (a and b);
    layer6_outputs(5049) <= not b or a;
    layer6_outputs(5050) <= not (a and b);
    layer6_outputs(5051) <= a and not b;
    layer6_outputs(5052) <= a;
    layer6_outputs(5053) <= not b;
    layer6_outputs(5054) <= not b;
    layer6_outputs(5055) <= not (a xor b);
    layer6_outputs(5056) <= '0';
    layer6_outputs(5057) <= not (a and b);
    layer6_outputs(5058) <= not (a xor b);
    layer6_outputs(5059) <= not (a xor b);
    layer6_outputs(5060) <= a xor b;
    layer6_outputs(5061) <= b;
    layer6_outputs(5062) <= not b;
    layer6_outputs(5063) <= not b or a;
    layer6_outputs(5064) <= a;
    layer6_outputs(5065) <= not a;
    layer6_outputs(5066) <= a;
    layer6_outputs(5067) <= not a;
    layer6_outputs(5068) <= not (a or b);
    layer6_outputs(5069) <= not (a or b);
    layer6_outputs(5070) <= not a or b;
    layer6_outputs(5071) <= b;
    layer6_outputs(5072) <= not (a or b);
    layer6_outputs(5073) <= not (a xor b);
    layer6_outputs(5074) <= b;
    layer6_outputs(5075) <= not a;
    layer6_outputs(5076) <= not (a xor b);
    layer6_outputs(5077) <= a or b;
    layer6_outputs(5078) <= not a or b;
    layer6_outputs(5079) <= not a;
    layer6_outputs(5080) <= not (a and b);
    layer6_outputs(5081) <= b;
    layer6_outputs(5082) <= '0';
    layer6_outputs(5083) <= not (a or b);
    layer6_outputs(5084) <= not b;
    layer6_outputs(5085) <= b;
    layer6_outputs(5086) <= not (a and b);
    layer6_outputs(5087) <= a xor b;
    layer6_outputs(5088) <= not a;
    layer6_outputs(5089) <= not (a xor b);
    layer6_outputs(5090) <= a xor b;
    layer6_outputs(5091) <= a or b;
    layer6_outputs(5092) <= not a;
    layer6_outputs(5093) <= not a;
    layer6_outputs(5094) <= not b;
    layer6_outputs(5095) <= a;
    layer6_outputs(5096) <= not a;
    layer6_outputs(5097) <= not (a xor b);
    layer6_outputs(5098) <= a;
    layer6_outputs(5099) <= not b or a;
    layer6_outputs(5100) <= not (a xor b);
    layer6_outputs(5101) <= b and not a;
    layer6_outputs(5102) <= a xor b;
    layer6_outputs(5103) <= a xor b;
    layer6_outputs(5104) <= not a;
    layer6_outputs(5105) <= a xor b;
    layer6_outputs(5106) <= not (a xor b);
    layer6_outputs(5107) <= a;
    layer6_outputs(5108) <= a;
    layer6_outputs(5109) <= a xor b;
    layer6_outputs(5110) <= a or b;
    layer6_outputs(5111) <= not b;
    layer6_outputs(5112) <= not (a xor b);
    layer6_outputs(5113) <= a;
    layer6_outputs(5114) <= not b or a;
    layer6_outputs(5115) <= a xor b;
    layer6_outputs(5116) <= a;
    layer6_outputs(5117) <= not a or b;
    layer6_outputs(5118) <= not (a or b);
    layer6_outputs(5119) <= not b;
    layer6_outputs(5120) <= a;
    layer6_outputs(5121) <= a and not b;
    layer6_outputs(5122) <= not a;
    layer6_outputs(5123) <= b;
    layer6_outputs(5124) <= not b;
    layer6_outputs(5125) <= a;
    layer6_outputs(5126) <= b;
    layer6_outputs(5127) <= a;
    layer6_outputs(5128) <= not (a xor b);
    layer6_outputs(5129) <= a xor b;
    layer6_outputs(5130) <= b;
    layer6_outputs(5131) <= not (a and b);
    layer6_outputs(5132) <= not a;
    layer6_outputs(5133) <= not a;
    layer6_outputs(5134) <= not a;
    layer6_outputs(5135) <= not a or b;
    layer6_outputs(5136) <= a xor b;
    layer6_outputs(5137) <= not (a xor b);
    layer6_outputs(5138) <= not b;
    layer6_outputs(5139) <= a;
    layer6_outputs(5140) <= not b;
    layer6_outputs(5141) <= not b;
    layer6_outputs(5142) <= not b;
    layer6_outputs(5143) <= a or b;
    layer6_outputs(5144) <= not (a xor b);
    layer6_outputs(5145) <= not a;
    layer6_outputs(5146) <= not a or b;
    layer6_outputs(5147) <= b;
    layer6_outputs(5148) <= not b;
    layer6_outputs(5149) <= a xor b;
    layer6_outputs(5150) <= not (a xor b);
    layer6_outputs(5151) <= b;
    layer6_outputs(5152) <= not (a xor b);
    layer6_outputs(5153) <= b and not a;
    layer6_outputs(5154) <= a xor b;
    layer6_outputs(5155) <= a and b;
    layer6_outputs(5156) <= not (a xor b);
    layer6_outputs(5157) <= not a;
    layer6_outputs(5158) <= not b;
    layer6_outputs(5159) <= a;
    layer6_outputs(5160) <= b and not a;
    layer6_outputs(5161) <= a xor b;
    layer6_outputs(5162) <= not a;
    layer6_outputs(5163) <= not a or b;
    layer6_outputs(5164) <= not (a and b);
    layer6_outputs(5165) <= a and b;
    layer6_outputs(5166) <= a or b;
    layer6_outputs(5167) <= not (a or b);
    layer6_outputs(5168) <= b;
    layer6_outputs(5169) <= not (a and b);
    layer6_outputs(5170) <= not (a or b);
    layer6_outputs(5171) <= not b;
    layer6_outputs(5172) <= not (a xor b);
    layer6_outputs(5173) <= b;
    layer6_outputs(5174) <= b;
    layer6_outputs(5175) <= not (a or b);
    layer6_outputs(5176) <= not a;
    layer6_outputs(5177) <= b;
    layer6_outputs(5178) <= not a;
    layer6_outputs(5179) <= a;
    layer6_outputs(5180) <= a;
    layer6_outputs(5181) <= a xor b;
    layer6_outputs(5182) <= not (a and b);
    layer6_outputs(5183) <= a and not b;
    layer6_outputs(5184) <= '0';
    layer6_outputs(5185) <= b and not a;
    layer6_outputs(5186) <= not b;
    layer6_outputs(5187) <= a;
    layer6_outputs(5188) <= not b or a;
    layer6_outputs(5189) <= not b or a;
    layer6_outputs(5190) <= not a or b;
    layer6_outputs(5191) <= not (a xor b);
    layer6_outputs(5192) <= b;
    layer6_outputs(5193) <= not b;
    layer6_outputs(5194) <= a xor b;
    layer6_outputs(5195) <= not (a and b);
    layer6_outputs(5196) <= not (a or b);
    layer6_outputs(5197) <= b;
    layer6_outputs(5198) <= a and b;
    layer6_outputs(5199) <= not a or b;
    layer6_outputs(5200) <= a xor b;
    layer6_outputs(5201) <= not a;
    layer6_outputs(5202) <= b;
    layer6_outputs(5203) <= b and not a;
    layer6_outputs(5204) <= a;
    layer6_outputs(5205) <= not (a xor b);
    layer6_outputs(5206) <= b;
    layer6_outputs(5207) <= a and not b;
    layer6_outputs(5208) <= not (a or b);
    layer6_outputs(5209) <= not b;
    layer6_outputs(5210) <= not (a xor b);
    layer6_outputs(5211) <= b and not a;
    layer6_outputs(5212) <= b;
    layer6_outputs(5213) <= not a;
    layer6_outputs(5214) <= not b;
    layer6_outputs(5215) <= b and not a;
    layer6_outputs(5216) <= not (a xor b);
    layer6_outputs(5217) <= not b;
    layer6_outputs(5218) <= not a;
    layer6_outputs(5219) <= b;
    layer6_outputs(5220) <= not (a and b);
    layer6_outputs(5221) <= not a;
    layer6_outputs(5222) <= not a;
    layer6_outputs(5223) <= a;
    layer6_outputs(5224) <= a and b;
    layer6_outputs(5225) <= not a or b;
    layer6_outputs(5226) <= not b;
    layer6_outputs(5227) <= not (a or b);
    layer6_outputs(5228) <= b;
    layer6_outputs(5229) <= b;
    layer6_outputs(5230) <= a;
    layer6_outputs(5231) <= not b or a;
    layer6_outputs(5232) <= not (a and b);
    layer6_outputs(5233) <= b;
    layer6_outputs(5234) <= a xor b;
    layer6_outputs(5235) <= not (a xor b);
    layer6_outputs(5236) <= a;
    layer6_outputs(5237) <= not (a xor b);
    layer6_outputs(5238) <= not (a or b);
    layer6_outputs(5239) <= not b;
    layer6_outputs(5240) <= a or b;
    layer6_outputs(5241) <= a xor b;
    layer6_outputs(5242) <= b;
    layer6_outputs(5243) <= b;
    layer6_outputs(5244) <= a xor b;
    layer6_outputs(5245) <= b;
    layer6_outputs(5246) <= not a or b;
    layer6_outputs(5247) <= not (a and b);
    layer6_outputs(5248) <= not a;
    layer6_outputs(5249) <= a or b;
    layer6_outputs(5250) <= a;
    layer6_outputs(5251) <= not (a xor b);
    layer6_outputs(5252) <= not b;
    layer6_outputs(5253) <= not (a xor b);
    layer6_outputs(5254) <= a and not b;
    layer6_outputs(5255) <= not a;
    layer6_outputs(5256) <= b;
    layer6_outputs(5257) <= not (a or b);
    layer6_outputs(5258) <= a and not b;
    layer6_outputs(5259) <= a or b;
    layer6_outputs(5260) <= b and not a;
    layer6_outputs(5261) <= not (a and b);
    layer6_outputs(5262) <= not (a or b);
    layer6_outputs(5263) <= not a;
    layer6_outputs(5264) <= not a or b;
    layer6_outputs(5265) <= a;
    layer6_outputs(5266) <= not (a xor b);
    layer6_outputs(5267) <= not b;
    layer6_outputs(5268) <= a;
    layer6_outputs(5269) <= b and not a;
    layer6_outputs(5270) <= b;
    layer6_outputs(5271) <= not (a xor b);
    layer6_outputs(5272) <= a and not b;
    layer6_outputs(5273) <= not b;
    layer6_outputs(5274) <= b;
    layer6_outputs(5275) <= not b;
    layer6_outputs(5276) <= a and b;
    layer6_outputs(5277) <= a and b;
    layer6_outputs(5278) <= b and not a;
    layer6_outputs(5279) <= a;
    layer6_outputs(5280) <= not b;
    layer6_outputs(5281) <= not a;
    layer6_outputs(5282) <= a xor b;
    layer6_outputs(5283) <= a xor b;
    layer6_outputs(5284) <= not (a and b);
    layer6_outputs(5285) <= not b or a;
    layer6_outputs(5286) <= a;
    layer6_outputs(5287) <= b;
    layer6_outputs(5288) <= a xor b;
    layer6_outputs(5289) <= a or b;
    layer6_outputs(5290) <= a and b;
    layer6_outputs(5291) <= a and b;
    layer6_outputs(5292) <= not b;
    layer6_outputs(5293) <= not a;
    layer6_outputs(5294) <= not b or a;
    layer6_outputs(5295) <= not b;
    layer6_outputs(5296) <= a and b;
    layer6_outputs(5297) <= not (a or b);
    layer6_outputs(5298) <= not (a or b);
    layer6_outputs(5299) <= not a;
    layer6_outputs(5300) <= a;
    layer6_outputs(5301) <= not a;
    layer6_outputs(5302) <= a;
    layer6_outputs(5303) <= not a or b;
    layer6_outputs(5304) <= not b;
    layer6_outputs(5305) <= not a or b;
    layer6_outputs(5306) <= not (a xor b);
    layer6_outputs(5307) <= not b;
    layer6_outputs(5308) <= a xor b;
    layer6_outputs(5309) <= not b;
    layer6_outputs(5310) <= not a or b;
    layer6_outputs(5311) <= not a;
    layer6_outputs(5312) <= a;
    layer6_outputs(5313) <= not a or b;
    layer6_outputs(5314) <= b;
    layer6_outputs(5315) <= b;
    layer6_outputs(5316) <= not b;
    layer6_outputs(5317) <= not b;
    layer6_outputs(5318) <= not (a and b);
    layer6_outputs(5319) <= not b;
    layer6_outputs(5320) <= b;
    layer6_outputs(5321) <= not b or a;
    layer6_outputs(5322) <= not (a or b);
    layer6_outputs(5323) <= not (a and b);
    layer6_outputs(5324) <= b;
    layer6_outputs(5325) <= not a or b;
    layer6_outputs(5326) <= not (a xor b);
    layer6_outputs(5327) <= a and b;
    layer6_outputs(5328) <= not (a and b);
    layer6_outputs(5329) <= not a;
    layer6_outputs(5330) <= not b;
    layer6_outputs(5331) <= '0';
    layer6_outputs(5332) <= not b;
    layer6_outputs(5333) <= not (a or b);
    layer6_outputs(5334) <= a;
    layer6_outputs(5335) <= not (a xor b);
    layer6_outputs(5336) <= a and b;
    layer6_outputs(5337) <= a or b;
    layer6_outputs(5338) <= not a;
    layer6_outputs(5339) <= a xor b;
    layer6_outputs(5340) <= a or b;
    layer6_outputs(5341) <= not (a xor b);
    layer6_outputs(5342) <= not a or b;
    layer6_outputs(5343) <= b;
    layer6_outputs(5344) <= a and b;
    layer6_outputs(5345) <= a or b;
    layer6_outputs(5346) <= not (a or b);
    layer6_outputs(5347) <= not a;
    layer6_outputs(5348) <= not (a xor b);
    layer6_outputs(5349) <= not a;
    layer6_outputs(5350) <= b and not a;
    layer6_outputs(5351) <= not a or b;
    layer6_outputs(5352) <= b and not a;
    layer6_outputs(5353) <= a or b;
    layer6_outputs(5354) <= not (a xor b);
    layer6_outputs(5355) <= a xor b;
    layer6_outputs(5356) <= not b or a;
    layer6_outputs(5357) <= not (a xor b);
    layer6_outputs(5358) <= b;
    layer6_outputs(5359) <= '1';
    layer6_outputs(5360) <= a;
    layer6_outputs(5361) <= b;
    layer6_outputs(5362) <= b;
    layer6_outputs(5363) <= not a;
    layer6_outputs(5364) <= a xor b;
    layer6_outputs(5365) <= not (a xor b);
    layer6_outputs(5366) <= b and not a;
    layer6_outputs(5367) <= not (a xor b);
    layer6_outputs(5368) <= not a;
    layer6_outputs(5369) <= a and b;
    layer6_outputs(5370) <= not b;
    layer6_outputs(5371) <= b and not a;
    layer6_outputs(5372) <= not b;
    layer6_outputs(5373) <= a or b;
    layer6_outputs(5374) <= a xor b;
    layer6_outputs(5375) <= not a;
    layer6_outputs(5376) <= b;
    layer6_outputs(5377) <= not a;
    layer6_outputs(5378) <= a or b;
    layer6_outputs(5379) <= a and b;
    layer6_outputs(5380) <= a xor b;
    layer6_outputs(5381) <= a and b;
    layer6_outputs(5382) <= a or b;
    layer6_outputs(5383) <= not (a or b);
    layer6_outputs(5384) <= not a or b;
    layer6_outputs(5385) <= not (a and b);
    layer6_outputs(5386) <= not a;
    layer6_outputs(5387) <= a and b;
    layer6_outputs(5388) <= a or b;
    layer6_outputs(5389) <= a and b;
    layer6_outputs(5390) <= not a or b;
    layer6_outputs(5391) <= b;
    layer6_outputs(5392) <= a xor b;
    layer6_outputs(5393) <= not a;
    layer6_outputs(5394) <= not (a or b);
    layer6_outputs(5395) <= not (a xor b);
    layer6_outputs(5396) <= not a or b;
    layer6_outputs(5397) <= not (a xor b);
    layer6_outputs(5398) <= a and not b;
    layer6_outputs(5399) <= not (a xor b);
    layer6_outputs(5400) <= a xor b;
    layer6_outputs(5401) <= a or b;
    layer6_outputs(5402) <= a xor b;
    layer6_outputs(5403) <= a xor b;
    layer6_outputs(5404) <= not a;
    layer6_outputs(5405) <= a;
    layer6_outputs(5406) <= b and not a;
    layer6_outputs(5407) <= b and not a;
    layer6_outputs(5408) <= not (a and b);
    layer6_outputs(5409) <= a;
    layer6_outputs(5410) <= not b;
    layer6_outputs(5411) <= a xor b;
    layer6_outputs(5412) <= not (a or b);
    layer6_outputs(5413) <= not (a or b);
    layer6_outputs(5414) <= b;
    layer6_outputs(5415) <= a;
    layer6_outputs(5416) <= a xor b;
    layer6_outputs(5417) <= a xor b;
    layer6_outputs(5418) <= a;
    layer6_outputs(5419) <= not b or a;
    layer6_outputs(5420) <= not (a and b);
    layer6_outputs(5421) <= not b;
    layer6_outputs(5422) <= a xor b;
    layer6_outputs(5423) <= b;
    layer6_outputs(5424) <= not a;
    layer6_outputs(5425) <= a xor b;
    layer6_outputs(5426) <= a xor b;
    layer6_outputs(5427) <= b;
    layer6_outputs(5428) <= a xor b;
    layer6_outputs(5429) <= '0';
    layer6_outputs(5430) <= not a or b;
    layer6_outputs(5431) <= not a;
    layer6_outputs(5432) <= b;
    layer6_outputs(5433) <= not a or b;
    layer6_outputs(5434) <= a;
    layer6_outputs(5435) <= not (a or b);
    layer6_outputs(5436) <= a and b;
    layer6_outputs(5437) <= not (a xor b);
    layer6_outputs(5438) <= a and b;
    layer6_outputs(5439) <= b and not a;
    layer6_outputs(5440) <= a;
    layer6_outputs(5441) <= a xor b;
    layer6_outputs(5442) <= not (a xor b);
    layer6_outputs(5443) <= a and b;
    layer6_outputs(5444) <= not (a and b);
    layer6_outputs(5445) <= not b;
    layer6_outputs(5446) <= a xor b;
    layer6_outputs(5447) <= a xor b;
    layer6_outputs(5448) <= b;
    layer6_outputs(5449) <= not (a and b);
    layer6_outputs(5450) <= a xor b;
    layer6_outputs(5451) <= a xor b;
    layer6_outputs(5452) <= not (a xor b);
    layer6_outputs(5453) <= b;
    layer6_outputs(5454) <= not b or a;
    layer6_outputs(5455) <= a;
    layer6_outputs(5456) <= a;
    layer6_outputs(5457) <= b;
    layer6_outputs(5458) <= b;
    layer6_outputs(5459) <= a xor b;
    layer6_outputs(5460) <= b and not a;
    layer6_outputs(5461) <= not b;
    layer6_outputs(5462) <= a and b;
    layer6_outputs(5463) <= not b or a;
    layer6_outputs(5464) <= a;
    layer6_outputs(5465) <= a xor b;
    layer6_outputs(5466) <= a xor b;
    layer6_outputs(5467) <= not a;
    layer6_outputs(5468) <= not a;
    layer6_outputs(5469) <= a and not b;
    layer6_outputs(5470) <= b and not a;
    layer6_outputs(5471) <= b and not a;
    layer6_outputs(5472) <= a;
    layer6_outputs(5473) <= not b;
    layer6_outputs(5474) <= not a;
    layer6_outputs(5475) <= not a;
    layer6_outputs(5476) <= not (a xor b);
    layer6_outputs(5477) <= not a;
    layer6_outputs(5478) <= not (a xor b);
    layer6_outputs(5479) <= not b;
    layer6_outputs(5480) <= '1';
    layer6_outputs(5481) <= not (a and b);
    layer6_outputs(5482) <= '1';
    layer6_outputs(5483) <= not (a and b);
    layer6_outputs(5484) <= b and not a;
    layer6_outputs(5485) <= not b or a;
    layer6_outputs(5486) <= b;
    layer6_outputs(5487) <= a;
    layer6_outputs(5488) <= not b;
    layer6_outputs(5489) <= a and b;
    layer6_outputs(5490) <= not (a and b);
    layer6_outputs(5491) <= a or b;
    layer6_outputs(5492) <= b and not a;
    layer6_outputs(5493) <= b and not a;
    layer6_outputs(5494) <= a;
    layer6_outputs(5495) <= a;
    layer6_outputs(5496) <= b;
    layer6_outputs(5497) <= not (a or b);
    layer6_outputs(5498) <= a and b;
    layer6_outputs(5499) <= a or b;
    layer6_outputs(5500) <= b and not a;
    layer6_outputs(5501) <= a and b;
    layer6_outputs(5502) <= not (a and b);
    layer6_outputs(5503) <= a or b;
    layer6_outputs(5504) <= not a;
    layer6_outputs(5505) <= b;
    layer6_outputs(5506) <= b;
    layer6_outputs(5507) <= not a or b;
    layer6_outputs(5508) <= a;
    layer6_outputs(5509) <= a xor b;
    layer6_outputs(5510) <= a and b;
    layer6_outputs(5511) <= not a or b;
    layer6_outputs(5512) <= b;
    layer6_outputs(5513) <= not (a xor b);
    layer6_outputs(5514) <= not (a xor b);
    layer6_outputs(5515) <= b;
    layer6_outputs(5516) <= not (a xor b);
    layer6_outputs(5517) <= a or b;
    layer6_outputs(5518) <= b;
    layer6_outputs(5519) <= a and not b;
    layer6_outputs(5520) <= not a;
    layer6_outputs(5521) <= not b;
    layer6_outputs(5522) <= a;
    layer6_outputs(5523) <= not a;
    layer6_outputs(5524) <= a or b;
    layer6_outputs(5525) <= a xor b;
    layer6_outputs(5526) <= b;
    layer6_outputs(5527) <= a xor b;
    layer6_outputs(5528) <= b;
    layer6_outputs(5529) <= not a;
    layer6_outputs(5530) <= a xor b;
    layer6_outputs(5531) <= not (a xor b);
    layer6_outputs(5532) <= a and b;
    layer6_outputs(5533) <= a;
    layer6_outputs(5534) <= a;
    layer6_outputs(5535) <= not b or a;
    layer6_outputs(5536) <= b and not a;
    layer6_outputs(5537) <= a or b;
    layer6_outputs(5538) <= a xor b;
    layer6_outputs(5539) <= not (a xor b);
    layer6_outputs(5540) <= not (a xor b);
    layer6_outputs(5541) <= b;
    layer6_outputs(5542) <= b;
    layer6_outputs(5543) <= b;
    layer6_outputs(5544) <= a xor b;
    layer6_outputs(5545) <= a or b;
    layer6_outputs(5546) <= not a;
    layer6_outputs(5547) <= not (a and b);
    layer6_outputs(5548) <= a xor b;
    layer6_outputs(5549) <= not a;
    layer6_outputs(5550) <= not (a xor b);
    layer6_outputs(5551) <= b;
    layer6_outputs(5552) <= b and not a;
    layer6_outputs(5553) <= not a;
    layer6_outputs(5554) <= not (a and b);
    layer6_outputs(5555) <= not (a or b);
    layer6_outputs(5556) <= b and not a;
    layer6_outputs(5557) <= b and not a;
    layer6_outputs(5558) <= a xor b;
    layer6_outputs(5559) <= a and b;
    layer6_outputs(5560) <= not b;
    layer6_outputs(5561) <= b and not a;
    layer6_outputs(5562) <= a and b;
    layer6_outputs(5563) <= not a;
    layer6_outputs(5564) <= not a or b;
    layer6_outputs(5565) <= b and not a;
    layer6_outputs(5566) <= a xor b;
    layer6_outputs(5567) <= not b or a;
    layer6_outputs(5568) <= not b;
    layer6_outputs(5569) <= not b;
    layer6_outputs(5570) <= not a;
    layer6_outputs(5571) <= a;
    layer6_outputs(5572) <= not (a and b);
    layer6_outputs(5573) <= not (a xor b);
    layer6_outputs(5574) <= not a or b;
    layer6_outputs(5575) <= a;
    layer6_outputs(5576) <= a;
    layer6_outputs(5577) <= not a;
    layer6_outputs(5578) <= not b;
    layer6_outputs(5579) <= a;
    layer6_outputs(5580) <= not a;
    layer6_outputs(5581) <= b;
    layer6_outputs(5582) <= a xor b;
    layer6_outputs(5583) <= a;
    layer6_outputs(5584) <= a or b;
    layer6_outputs(5585) <= a;
    layer6_outputs(5586) <= b and not a;
    layer6_outputs(5587) <= a;
    layer6_outputs(5588) <= a or b;
    layer6_outputs(5589) <= not b;
    layer6_outputs(5590) <= not (a or b);
    layer6_outputs(5591) <= b and not a;
    layer6_outputs(5592) <= b;
    layer6_outputs(5593) <= b;
    layer6_outputs(5594) <= b;
    layer6_outputs(5595) <= a;
    layer6_outputs(5596) <= not a;
    layer6_outputs(5597) <= b;
    layer6_outputs(5598) <= not (a xor b);
    layer6_outputs(5599) <= a and not b;
    layer6_outputs(5600) <= not b;
    layer6_outputs(5601) <= not a or b;
    layer6_outputs(5602) <= a and b;
    layer6_outputs(5603) <= b;
    layer6_outputs(5604) <= a xor b;
    layer6_outputs(5605) <= b and not a;
    layer6_outputs(5606) <= a xor b;
    layer6_outputs(5607) <= b;
    layer6_outputs(5608) <= not b;
    layer6_outputs(5609) <= a and b;
    layer6_outputs(5610) <= a xor b;
    layer6_outputs(5611) <= a or b;
    layer6_outputs(5612) <= a;
    layer6_outputs(5613) <= '1';
    layer6_outputs(5614) <= not (a xor b);
    layer6_outputs(5615) <= a xor b;
    layer6_outputs(5616) <= not a;
    layer6_outputs(5617) <= a and not b;
    layer6_outputs(5618) <= not a;
    layer6_outputs(5619) <= not a;
    layer6_outputs(5620) <= a or b;
    layer6_outputs(5621) <= not a;
    layer6_outputs(5622) <= not (a or b);
    layer6_outputs(5623) <= a xor b;
    layer6_outputs(5624) <= b and not a;
    layer6_outputs(5625) <= '0';
    layer6_outputs(5626) <= not a;
    layer6_outputs(5627) <= a and b;
    layer6_outputs(5628) <= not a;
    layer6_outputs(5629) <= '0';
    layer6_outputs(5630) <= not b or a;
    layer6_outputs(5631) <= not a or b;
    layer6_outputs(5632) <= not a;
    layer6_outputs(5633) <= not b;
    layer6_outputs(5634) <= not (a xor b);
    layer6_outputs(5635) <= not a;
    layer6_outputs(5636) <= not b;
    layer6_outputs(5637) <= a xor b;
    layer6_outputs(5638) <= not b;
    layer6_outputs(5639) <= a and b;
    layer6_outputs(5640) <= not b;
    layer6_outputs(5641) <= not b or a;
    layer6_outputs(5642) <= a;
    layer6_outputs(5643) <= not (a xor b);
    layer6_outputs(5644) <= a or b;
    layer6_outputs(5645) <= not b;
    layer6_outputs(5646) <= not (a and b);
    layer6_outputs(5647) <= not (a xor b);
    layer6_outputs(5648) <= b;
    layer6_outputs(5649) <= not a or b;
    layer6_outputs(5650) <= not b;
    layer6_outputs(5651) <= not (a xor b);
    layer6_outputs(5652) <= a or b;
    layer6_outputs(5653) <= not a or b;
    layer6_outputs(5654) <= not b or a;
    layer6_outputs(5655) <= not (a and b);
    layer6_outputs(5656) <= not (a and b);
    layer6_outputs(5657) <= not (a xor b);
    layer6_outputs(5658) <= not (a xor b);
    layer6_outputs(5659) <= a;
    layer6_outputs(5660) <= not b;
    layer6_outputs(5661) <= a and not b;
    layer6_outputs(5662) <= a xor b;
    layer6_outputs(5663) <= a and b;
    layer6_outputs(5664) <= b;
    layer6_outputs(5665) <= not b;
    layer6_outputs(5666) <= not (a xor b);
    layer6_outputs(5667) <= not b or a;
    layer6_outputs(5668) <= not (a xor b);
    layer6_outputs(5669) <= b;
    layer6_outputs(5670) <= a;
    layer6_outputs(5671) <= a or b;
    layer6_outputs(5672) <= a and b;
    layer6_outputs(5673) <= b;
    layer6_outputs(5674) <= b;
    layer6_outputs(5675) <= a;
    layer6_outputs(5676) <= a xor b;
    layer6_outputs(5677) <= b;
    layer6_outputs(5678) <= not (a and b);
    layer6_outputs(5679) <= a;
    layer6_outputs(5680) <= a and b;
    layer6_outputs(5681) <= a xor b;
    layer6_outputs(5682) <= not b;
    layer6_outputs(5683) <= a;
    layer6_outputs(5684) <= a xor b;
    layer6_outputs(5685) <= a and b;
    layer6_outputs(5686) <= not (a xor b);
    layer6_outputs(5687) <= a;
    layer6_outputs(5688) <= not a;
    layer6_outputs(5689) <= not (a and b);
    layer6_outputs(5690) <= not a;
    layer6_outputs(5691) <= not (a or b);
    layer6_outputs(5692) <= a or b;
    layer6_outputs(5693) <= not b;
    layer6_outputs(5694) <= a or b;
    layer6_outputs(5695) <= a;
    layer6_outputs(5696) <= b and not a;
    layer6_outputs(5697) <= not a;
    layer6_outputs(5698) <= a or b;
    layer6_outputs(5699) <= not b or a;
    layer6_outputs(5700) <= not b;
    layer6_outputs(5701) <= b;
    layer6_outputs(5702) <= a;
    layer6_outputs(5703) <= not (a xor b);
    layer6_outputs(5704) <= not b;
    layer6_outputs(5705) <= not b or a;
    layer6_outputs(5706) <= not a;
    layer6_outputs(5707) <= not b or a;
    layer6_outputs(5708) <= not (a or b);
    layer6_outputs(5709) <= not a;
    layer6_outputs(5710) <= a or b;
    layer6_outputs(5711) <= a and b;
    layer6_outputs(5712) <= not b;
    layer6_outputs(5713) <= a and b;
    layer6_outputs(5714) <= not (a or b);
    layer6_outputs(5715) <= not a;
    layer6_outputs(5716) <= b and not a;
    layer6_outputs(5717) <= not b;
    layer6_outputs(5718) <= b;
    layer6_outputs(5719) <= a and b;
    layer6_outputs(5720) <= not b;
    layer6_outputs(5721) <= a;
    layer6_outputs(5722) <= not b;
    layer6_outputs(5723) <= not a;
    layer6_outputs(5724) <= a xor b;
    layer6_outputs(5725) <= not (a xor b);
    layer6_outputs(5726) <= a;
    layer6_outputs(5727) <= not b;
    layer6_outputs(5728) <= a xor b;
    layer6_outputs(5729) <= b;
    layer6_outputs(5730) <= not b;
    layer6_outputs(5731) <= a xor b;
    layer6_outputs(5732) <= not b;
    layer6_outputs(5733) <= not a;
    layer6_outputs(5734) <= not b or a;
    layer6_outputs(5735) <= a;
    layer6_outputs(5736) <= a;
    layer6_outputs(5737) <= a xor b;
    layer6_outputs(5738) <= b;
    layer6_outputs(5739) <= b and not a;
    layer6_outputs(5740) <= not (a or b);
    layer6_outputs(5741) <= not a;
    layer6_outputs(5742) <= not a or b;
    layer6_outputs(5743) <= a or b;
    layer6_outputs(5744) <= a and not b;
    layer6_outputs(5745) <= not a;
    layer6_outputs(5746) <= a;
    layer6_outputs(5747) <= b;
    layer6_outputs(5748) <= b and not a;
    layer6_outputs(5749) <= a;
    layer6_outputs(5750) <= not a;
    layer6_outputs(5751) <= b and not a;
    layer6_outputs(5752) <= not b or a;
    layer6_outputs(5753) <= a or b;
    layer6_outputs(5754) <= a;
    layer6_outputs(5755) <= a and b;
    layer6_outputs(5756) <= a;
    layer6_outputs(5757) <= not b or a;
    layer6_outputs(5758) <= not a or b;
    layer6_outputs(5759) <= a and not b;
    layer6_outputs(5760) <= b;
    layer6_outputs(5761) <= not b;
    layer6_outputs(5762) <= a or b;
    layer6_outputs(5763) <= not (a or b);
    layer6_outputs(5764) <= b;
    layer6_outputs(5765) <= a xor b;
    layer6_outputs(5766) <= a;
    layer6_outputs(5767) <= a and b;
    layer6_outputs(5768) <= a and b;
    layer6_outputs(5769) <= b and not a;
    layer6_outputs(5770) <= not b or a;
    layer6_outputs(5771) <= not a;
    layer6_outputs(5772) <= not (a xor b);
    layer6_outputs(5773) <= a;
    layer6_outputs(5774) <= a;
    layer6_outputs(5775) <= not (a and b);
    layer6_outputs(5776) <= not (a or b);
    layer6_outputs(5777) <= not b or a;
    layer6_outputs(5778) <= a;
    layer6_outputs(5779) <= '1';
    layer6_outputs(5780) <= not a or b;
    layer6_outputs(5781) <= b;
    layer6_outputs(5782) <= not (a and b);
    layer6_outputs(5783) <= a;
    layer6_outputs(5784) <= b;
    layer6_outputs(5785) <= a or b;
    layer6_outputs(5786) <= b;
    layer6_outputs(5787) <= not a;
    layer6_outputs(5788) <= not (a xor b);
    layer6_outputs(5789) <= '1';
    layer6_outputs(5790) <= not a or b;
    layer6_outputs(5791) <= a xor b;
    layer6_outputs(5792) <= not b;
    layer6_outputs(5793) <= b;
    layer6_outputs(5794) <= a xor b;
    layer6_outputs(5795) <= not (a and b);
    layer6_outputs(5796) <= not a;
    layer6_outputs(5797) <= a and b;
    layer6_outputs(5798) <= a and b;
    layer6_outputs(5799) <= not (a or b);
    layer6_outputs(5800) <= a and b;
    layer6_outputs(5801) <= b;
    layer6_outputs(5802) <= not a;
    layer6_outputs(5803) <= b;
    layer6_outputs(5804) <= not a;
    layer6_outputs(5805) <= a;
    layer6_outputs(5806) <= not b;
    layer6_outputs(5807) <= a and not b;
    layer6_outputs(5808) <= not (a xor b);
    layer6_outputs(5809) <= not b;
    layer6_outputs(5810) <= b;
    layer6_outputs(5811) <= b;
    layer6_outputs(5812) <= a and not b;
    layer6_outputs(5813) <= a xor b;
    layer6_outputs(5814) <= not (a xor b);
    layer6_outputs(5815) <= a and b;
    layer6_outputs(5816) <= b;
    layer6_outputs(5817) <= a;
    layer6_outputs(5818) <= a and b;
    layer6_outputs(5819) <= b;
    layer6_outputs(5820) <= not b;
    layer6_outputs(5821) <= not b;
    layer6_outputs(5822) <= b;
    layer6_outputs(5823) <= b;
    layer6_outputs(5824) <= not b;
    layer6_outputs(5825) <= not b;
    layer6_outputs(5826) <= b;
    layer6_outputs(5827) <= not (a xor b);
    layer6_outputs(5828) <= a xor b;
    layer6_outputs(5829) <= b and not a;
    layer6_outputs(5830) <= not b or a;
    layer6_outputs(5831) <= a;
    layer6_outputs(5832) <= a and b;
    layer6_outputs(5833) <= a xor b;
    layer6_outputs(5834) <= not a;
    layer6_outputs(5835) <= not b;
    layer6_outputs(5836) <= a xor b;
    layer6_outputs(5837) <= a and not b;
    layer6_outputs(5838) <= not a or b;
    layer6_outputs(5839) <= a and b;
    layer6_outputs(5840) <= not a;
    layer6_outputs(5841) <= a;
    layer6_outputs(5842) <= not a;
    layer6_outputs(5843) <= b;
    layer6_outputs(5844) <= b;
    layer6_outputs(5845) <= b;
    layer6_outputs(5846) <= b;
    layer6_outputs(5847) <= b and not a;
    layer6_outputs(5848) <= not a;
    layer6_outputs(5849) <= a and not b;
    layer6_outputs(5850) <= b;
    layer6_outputs(5851) <= not b or a;
    layer6_outputs(5852) <= not (a or b);
    layer6_outputs(5853) <= b and not a;
    layer6_outputs(5854) <= a and b;
    layer6_outputs(5855) <= not b;
    layer6_outputs(5856) <= a and not b;
    layer6_outputs(5857) <= not (a xor b);
    layer6_outputs(5858) <= not a;
    layer6_outputs(5859) <= a or b;
    layer6_outputs(5860) <= a;
    layer6_outputs(5861) <= not b or a;
    layer6_outputs(5862) <= a;
    layer6_outputs(5863) <= not b;
    layer6_outputs(5864) <= not b;
    layer6_outputs(5865) <= b and not a;
    layer6_outputs(5866) <= b;
    layer6_outputs(5867) <= b;
    layer6_outputs(5868) <= not (a xor b);
    layer6_outputs(5869) <= not (a or b);
    layer6_outputs(5870) <= not b;
    layer6_outputs(5871) <= b and not a;
    layer6_outputs(5872) <= not b;
    layer6_outputs(5873) <= a or b;
    layer6_outputs(5874) <= a;
    layer6_outputs(5875) <= a;
    layer6_outputs(5876) <= b;
    layer6_outputs(5877) <= not (a and b);
    layer6_outputs(5878) <= not b or a;
    layer6_outputs(5879) <= a or b;
    layer6_outputs(5880) <= a and b;
    layer6_outputs(5881) <= not a;
    layer6_outputs(5882) <= not b;
    layer6_outputs(5883) <= not b or a;
    layer6_outputs(5884) <= a and b;
    layer6_outputs(5885) <= b;
    layer6_outputs(5886) <= not (a and b);
    layer6_outputs(5887) <= b;
    layer6_outputs(5888) <= a or b;
    layer6_outputs(5889) <= a xor b;
    layer6_outputs(5890) <= b;
    layer6_outputs(5891) <= not a;
    layer6_outputs(5892) <= not b;
    layer6_outputs(5893) <= a xor b;
    layer6_outputs(5894) <= not b;
    layer6_outputs(5895) <= not b;
    layer6_outputs(5896) <= b;
    layer6_outputs(5897) <= b;
    layer6_outputs(5898) <= not a;
    layer6_outputs(5899) <= b;
    layer6_outputs(5900) <= not a;
    layer6_outputs(5901) <= not a;
    layer6_outputs(5902) <= not a;
    layer6_outputs(5903) <= not b;
    layer6_outputs(5904) <= b;
    layer6_outputs(5905) <= not b or a;
    layer6_outputs(5906) <= b and not a;
    layer6_outputs(5907) <= a;
    layer6_outputs(5908) <= not (a xor b);
    layer6_outputs(5909) <= a xor b;
    layer6_outputs(5910) <= a xor b;
    layer6_outputs(5911) <= b and not a;
    layer6_outputs(5912) <= not (a and b);
    layer6_outputs(5913) <= not a;
    layer6_outputs(5914) <= a;
    layer6_outputs(5915) <= a;
    layer6_outputs(5916) <= not a;
    layer6_outputs(5917) <= not a;
    layer6_outputs(5918) <= a xor b;
    layer6_outputs(5919) <= not b;
    layer6_outputs(5920) <= a;
    layer6_outputs(5921) <= a or b;
    layer6_outputs(5922) <= not (a xor b);
    layer6_outputs(5923) <= not a or b;
    layer6_outputs(5924) <= b and not a;
    layer6_outputs(5925) <= a xor b;
    layer6_outputs(5926) <= not (a xor b);
    layer6_outputs(5927) <= a;
    layer6_outputs(5928) <= not a or b;
    layer6_outputs(5929) <= a xor b;
    layer6_outputs(5930) <= not a;
    layer6_outputs(5931) <= not b;
    layer6_outputs(5932) <= a or b;
    layer6_outputs(5933) <= a;
    layer6_outputs(5934) <= not b;
    layer6_outputs(5935) <= not b;
    layer6_outputs(5936) <= a;
    layer6_outputs(5937) <= b;
    layer6_outputs(5938) <= a;
    layer6_outputs(5939) <= not a or b;
    layer6_outputs(5940) <= not b;
    layer6_outputs(5941) <= not (a and b);
    layer6_outputs(5942) <= a xor b;
    layer6_outputs(5943) <= a and b;
    layer6_outputs(5944) <= a and not b;
    layer6_outputs(5945) <= a and b;
    layer6_outputs(5946) <= a xor b;
    layer6_outputs(5947) <= not b;
    layer6_outputs(5948) <= b;
    layer6_outputs(5949) <= b;
    layer6_outputs(5950) <= a xor b;
    layer6_outputs(5951) <= not a;
    layer6_outputs(5952) <= b;
    layer6_outputs(5953) <= b;
    layer6_outputs(5954) <= a xor b;
    layer6_outputs(5955) <= b;
    layer6_outputs(5956) <= a xor b;
    layer6_outputs(5957) <= a;
    layer6_outputs(5958) <= not a;
    layer6_outputs(5959) <= not (a and b);
    layer6_outputs(5960) <= not (a or b);
    layer6_outputs(5961) <= not a;
    layer6_outputs(5962) <= b;
    layer6_outputs(5963) <= b;
    layer6_outputs(5964) <= b;
    layer6_outputs(5965) <= b;
    layer6_outputs(5966) <= not b;
    layer6_outputs(5967) <= a and b;
    layer6_outputs(5968) <= not a or b;
    layer6_outputs(5969) <= b;
    layer6_outputs(5970) <= not (a xor b);
    layer6_outputs(5971) <= a and not b;
    layer6_outputs(5972) <= not a;
    layer6_outputs(5973) <= b;
    layer6_outputs(5974) <= not a or b;
    layer6_outputs(5975) <= a xor b;
    layer6_outputs(5976) <= not b;
    layer6_outputs(5977) <= a and b;
    layer6_outputs(5978) <= not b;
    layer6_outputs(5979) <= a xor b;
    layer6_outputs(5980) <= not a;
    layer6_outputs(5981) <= a xor b;
    layer6_outputs(5982) <= not b or a;
    layer6_outputs(5983) <= a or b;
    layer6_outputs(5984) <= not (a xor b);
    layer6_outputs(5985) <= not a;
    layer6_outputs(5986) <= b and not a;
    layer6_outputs(5987) <= not a;
    layer6_outputs(5988) <= not (a or b);
    layer6_outputs(5989) <= not a;
    layer6_outputs(5990) <= not (a xor b);
    layer6_outputs(5991) <= not a;
    layer6_outputs(5992) <= not a or b;
    layer6_outputs(5993) <= a;
    layer6_outputs(5994) <= a;
    layer6_outputs(5995) <= not a or b;
    layer6_outputs(5996) <= a and not b;
    layer6_outputs(5997) <= b;
    layer6_outputs(5998) <= not (a and b);
    layer6_outputs(5999) <= a and not b;
    layer6_outputs(6000) <= not (a or b);
    layer6_outputs(6001) <= not b;
    layer6_outputs(6002) <= b;
    layer6_outputs(6003) <= a xor b;
    layer6_outputs(6004) <= not (a xor b);
    layer6_outputs(6005) <= b;
    layer6_outputs(6006) <= not a or b;
    layer6_outputs(6007) <= not (a xor b);
    layer6_outputs(6008) <= not b;
    layer6_outputs(6009) <= a xor b;
    layer6_outputs(6010) <= a and b;
    layer6_outputs(6011) <= not (a xor b);
    layer6_outputs(6012) <= a;
    layer6_outputs(6013) <= a xor b;
    layer6_outputs(6014) <= not (a xor b);
    layer6_outputs(6015) <= not (a and b);
    layer6_outputs(6016) <= not (a xor b);
    layer6_outputs(6017) <= a xor b;
    layer6_outputs(6018) <= not b or a;
    layer6_outputs(6019) <= b;
    layer6_outputs(6020) <= a xor b;
    layer6_outputs(6021) <= not (a xor b);
    layer6_outputs(6022) <= not a;
    layer6_outputs(6023) <= not (a and b);
    layer6_outputs(6024) <= not (a or b);
    layer6_outputs(6025) <= not a;
    layer6_outputs(6026) <= a and b;
    layer6_outputs(6027) <= a xor b;
    layer6_outputs(6028) <= a;
    layer6_outputs(6029) <= not a;
    layer6_outputs(6030) <= a and b;
    layer6_outputs(6031) <= not (a or b);
    layer6_outputs(6032) <= not b or a;
    layer6_outputs(6033) <= not b or a;
    layer6_outputs(6034) <= a;
    layer6_outputs(6035) <= not a or b;
    layer6_outputs(6036) <= not b;
    layer6_outputs(6037) <= not b;
    layer6_outputs(6038) <= not b;
    layer6_outputs(6039) <= a or b;
    layer6_outputs(6040) <= not a or b;
    layer6_outputs(6041) <= not (a and b);
    layer6_outputs(6042) <= b and not a;
    layer6_outputs(6043) <= not (a or b);
    layer6_outputs(6044) <= not b;
    layer6_outputs(6045) <= not b;
    layer6_outputs(6046) <= not (a or b);
    layer6_outputs(6047) <= a xor b;
    layer6_outputs(6048) <= a;
    layer6_outputs(6049) <= a;
    layer6_outputs(6050) <= b;
    layer6_outputs(6051) <= a;
    layer6_outputs(6052) <= a and b;
    layer6_outputs(6053) <= not b;
    layer6_outputs(6054) <= a and b;
    layer6_outputs(6055) <= b and not a;
    layer6_outputs(6056) <= a;
    layer6_outputs(6057) <= a and b;
    layer6_outputs(6058) <= a and not b;
    layer6_outputs(6059) <= not (a xor b);
    layer6_outputs(6060) <= not b or a;
    layer6_outputs(6061) <= b;
    layer6_outputs(6062) <= not a;
    layer6_outputs(6063) <= b;
    layer6_outputs(6064) <= a;
    layer6_outputs(6065) <= not a;
    layer6_outputs(6066) <= a xor b;
    layer6_outputs(6067) <= not (a xor b);
    layer6_outputs(6068) <= a xor b;
    layer6_outputs(6069) <= not b or a;
    layer6_outputs(6070) <= not b;
    layer6_outputs(6071) <= a and not b;
    layer6_outputs(6072) <= not a or b;
    layer6_outputs(6073) <= not (a or b);
    layer6_outputs(6074) <= not a;
    layer6_outputs(6075) <= a and not b;
    layer6_outputs(6076) <= not b;
    layer6_outputs(6077) <= a xor b;
    layer6_outputs(6078) <= b;
    layer6_outputs(6079) <= a;
    layer6_outputs(6080) <= not (a xor b);
    layer6_outputs(6081) <= not (a and b);
    layer6_outputs(6082) <= b;
    layer6_outputs(6083) <= a and not b;
    layer6_outputs(6084) <= not (a xor b);
    layer6_outputs(6085) <= a;
    layer6_outputs(6086) <= a and not b;
    layer6_outputs(6087) <= b;
    layer6_outputs(6088) <= a and b;
    layer6_outputs(6089) <= not a;
    layer6_outputs(6090) <= a and not b;
    layer6_outputs(6091) <= b and not a;
    layer6_outputs(6092) <= b;
    layer6_outputs(6093) <= not b;
    layer6_outputs(6094) <= not b;
    layer6_outputs(6095) <= not a;
    layer6_outputs(6096) <= b and not a;
    layer6_outputs(6097) <= not a or b;
    layer6_outputs(6098) <= b;
    layer6_outputs(6099) <= b;
    layer6_outputs(6100) <= not (a xor b);
    layer6_outputs(6101) <= not (a xor b);
    layer6_outputs(6102) <= not (a or b);
    layer6_outputs(6103) <= b;
    layer6_outputs(6104) <= not a;
    layer6_outputs(6105) <= b;
    layer6_outputs(6106) <= a or b;
    layer6_outputs(6107) <= a xor b;
    layer6_outputs(6108) <= a xor b;
    layer6_outputs(6109) <= a xor b;
    layer6_outputs(6110) <= not a;
    layer6_outputs(6111) <= not b;
    layer6_outputs(6112) <= not a;
    layer6_outputs(6113) <= not a;
    layer6_outputs(6114) <= not b;
    layer6_outputs(6115) <= not b;
    layer6_outputs(6116) <= '1';
    layer6_outputs(6117) <= a xor b;
    layer6_outputs(6118) <= not (a and b);
    layer6_outputs(6119) <= not b;
    layer6_outputs(6120) <= a;
    layer6_outputs(6121) <= b;
    layer6_outputs(6122) <= a;
    layer6_outputs(6123) <= not (a and b);
    layer6_outputs(6124) <= not b;
    layer6_outputs(6125) <= a and not b;
    layer6_outputs(6126) <= a;
    layer6_outputs(6127) <= not b;
    layer6_outputs(6128) <= a and b;
    layer6_outputs(6129) <= a xor b;
    layer6_outputs(6130) <= not a or b;
    layer6_outputs(6131) <= a and b;
    layer6_outputs(6132) <= not b;
    layer6_outputs(6133) <= not a;
    layer6_outputs(6134) <= a and not b;
    layer6_outputs(6135) <= a and b;
    layer6_outputs(6136) <= not b;
    layer6_outputs(6137) <= a;
    layer6_outputs(6138) <= not a;
    layer6_outputs(6139) <= not b;
    layer6_outputs(6140) <= not b;
    layer6_outputs(6141) <= a;
    layer6_outputs(6142) <= b;
    layer6_outputs(6143) <= not b;
    layer6_outputs(6144) <= a;
    layer6_outputs(6145) <= b;
    layer6_outputs(6146) <= not (a or b);
    layer6_outputs(6147) <= not a;
    layer6_outputs(6148) <= not a;
    layer6_outputs(6149) <= a;
    layer6_outputs(6150) <= not b or a;
    layer6_outputs(6151) <= b and not a;
    layer6_outputs(6152) <= not (a xor b);
    layer6_outputs(6153) <= not (a xor b);
    layer6_outputs(6154) <= not (a xor b);
    layer6_outputs(6155) <= a xor b;
    layer6_outputs(6156) <= not a or b;
    layer6_outputs(6157) <= not (a or b);
    layer6_outputs(6158) <= not b;
    layer6_outputs(6159) <= a and not b;
    layer6_outputs(6160) <= a;
    layer6_outputs(6161) <= not a;
    layer6_outputs(6162) <= not a;
    layer6_outputs(6163) <= not (a and b);
    layer6_outputs(6164) <= b and not a;
    layer6_outputs(6165) <= not a;
    layer6_outputs(6166) <= a;
    layer6_outputs(6167) <= not a;
    layer6_outputs(6168) <= not (a xor b);
    layer6_outputs(6169) <= '1';
    layer6_outputs(6170) <= not a or b;
    layer6_outputs(6171) <= b and not a;
    layer6_outputs(6172) <= b;
    layer6_outputs(6173) <= not b;
    layer6_outputs(6174) <= not a;
    layer6_outputs(6175) <= a;
    layer6_outputs(6176) <= not (a xor b);
    layer6_outputs(6177) <= a and b;
    layer6_outputs(6178) <= not (a or b);
    layer6_outputs(6179) <= b;
    layer6_outputs(6180) <= not (a or b);
    layer6_outputs(6181) <= not b;
    layer6_outputs(6182) <= not (a and b);
    layer6_outputs(6183) <= a xor b;
    layer6_outputs(6184) <= not (a or b);
    layer6_outputs(6185) <= not a or b;
    layer6_outputs(6186) <= a;
    layer6_outputs(6187) <= a xor b;
    layer6_outputs(6188) <= not a or b;
    layer6_outputs(6189) <= not (a or b);
    layer6_outputs(6190) <= a or b;
    layer6_outputs(6191) <= a;
    layer6_outputs(6192) <= a;
    layer6_outputs(6193) <= not a;
    layer6_outputs(6194) <= a or b;
    layer6_outputs(6195) <= b and not a;
    layer6_outputs(6196) <= a and b;
    layer6_outputs(6197) <= not b;
    layer6_outputs(6198) <= not (a xor b);
    layer6_outputs(6199) <= b;
    layer6_outputs(6200) <= a xor b;
    layer6_outputs(6201) <= b and not a;
    layer6_outputs(6202) <= not a;
    layer6_outputs(6203) <= not (a xor b);
    layer6_outputs(6204) <= a and not b;
    layer6_outputs(6205) <= a;
    layer6_outputs(6206) <= b and not a;
    layer6_outputs(6207) <= not a or b;
    layer6_outputs(6208) <= not (a or b);
    layer6_outputs(6209) <= not (a xor b);
    layer6_outputs(6210) <= not a;
    layer6_outputs(6211) <= not a;
    layer6_outputs(6212) <= a;
    layer6_outputs(6213) <= a and b;
    layer6_outputs(6214) <= not a;
    layer6_outputs(6215) <= not b or a;
    layer6_outputs(6216) <= not a or b;
    layer6_outputs(6217) <= a;
    layer6_outputs(6218) <= not (a xor b);
    layer6_outputs(6219) <= not a;
    layer6_outputs(6220) <= not (a or b);
    layer6_outputs(6221) <= not a or b;
    layer6_outputs(6222) <= not (a xor b);
    layer6_outputs(6223) <= a xor b;
    layer6_outputs(6224) <= not b;
    layer6_outputs(6225) <= b and not a;
    layer6_outputs(6226) <= b;
    layer6_outputs(6227) <= b;
    layer6_outputs(6228) <= b;
    layer6_outputs(6229) <= not (a or b);
    layer6_outputs(6230) <= not a;
    layer6_outputs(6231) <= not a or b;
    layer6_outputs(6232) <= not a;
    layer6_outputs(6233) <= a;
    layer6_outputs(6234) <= not (a xor b);
    layer6_outputs(6235) <= not b;
    layer6_outputs(6236) <= not a or b;
    layer6_outputs(6237) <= not a or b;
    layer6_outputs(6238) <= not b;
    layer6_outputs(6239) <= not a;
    layer6_outputs(6240) <= b and not a;
    layer6_outputs(6241) <= not (a xor b);
    layer6_outputs(6242) <= not b;
    layer6_outputs(6243) <= not (a or b);
    layer6_outputs(6244) <= b;
    layer6_outputs(6245) <= a xor b;
    layer6_outputs(6246) <= a and not b;
    layer6_outputs(6247) <= not (a xor b);
    layer6_outputs(6248) <= a xor b;
    layer6_outputs(6249) <= not b;
    layer6_outputs(6250) <= not (a or b);
    layer6_outputs(6251) <= not b or a;
    layer6_outputs(6252) <= not (a xor b);
    layer6_outputs(6253) <= not (a xor b);
    layer6_outputs(6254) <= a;
    layer6_outputs(6255) <= not (a xor b);
    layer6_outputs(6256) <= not (a xor b);
    layer6_outputs(6257) <= a;
    layer6_outputs(6258) <= not b;
    layer6_outputs(6259) <= a xor b;
    layer6_outputs(6260) <= b;
    layer6_outputs(6261) <= not (a or b);
    layer6_outputs(6262) <= a xor b;
    layer6_outputs(6263) <= not (a xor b);
    layer6_outputs(6264) <= not b;
    layer6_outputs(6265) <= a and not b;
    layer6_outputs(6266) <= b;
    layer6_outputs(6267) <= a;
    layer6_outputs(6268) <= not b;
    layer6_outputs(6269) <= not b;
    layer6_outputs(6270) <= not b;
    layer6_outputs(6271) <= b and not a;
    layer6_outputs(6272) <= not b;
    layer6_outputs(6273) <= not b;
    layer6_outputs(6274) <= not a;
    layer6_outputs(6275) <= b;
    layer6_outputs(6276) <= '1';
    layer6_outputs(6277) <= not (a or b);
    layer6_outputs(6278) <= a and b;
    layer6_outputs(6279) <= b and not a;
    layer6_outputs(6280) <= not a or b;
    layer6_outputs(6281) <= not a;
    layer6_outputs(6282) <= not b;
    layer6_outputs(6283) <= b;
    layer6_outputs(6284) <= a or b;
    layer6_outputs(6285) <= not (a or b);
    layer6_outputs(6286) <= not (a xor b);
    layer6_outputs(6287) <= not b;
    layer6_outputs(6288) <= not (a xor b);
    layer6_outputs(6289) <= not (a or b);
    layer6_outputs(6290) <= not a;
    layer6_outputs(6291) <= not (a xor b);
    layer6_outputs(6292) <= not a or b;
    layer6_outputs(6293) <= a and not b;
    layer6_outputs(6294) <= b;
    layer6_outputs(6295) <= not a;
    layer6_outputs(6296) <= a xor b;
    layer6_outputs(6297) <= b;
    layer6_outputs(6298) <= a;
    layer6_outputs(6299) <= a xor b;
    layer6_outputs(6300) <= a or b;
    layer6_outputs(6301) <= a;
    layer6_outputs(6302) <= not b;
    layer6_outputs(6303) <= not (a xor b);
    layer6_outputs(6304) <= b;
    layer6_outputs(6305) <= not a;
    layer6_outputs(6306) <= a;
    layer6_outputs(6307) <= a or b;
    layer6_outputs(6308) <= not (a and b);
    layer6_outputs(6309) <= b;
    layer6_outputs(6310) <= a and not b;
    layer6_outputs(6311) <= not b or a;
    layer6_outputs(6312) <= not (a xor b);
    layer6_outputs(6313) <= b and not a;
    layer6_outputs(6314) <= not b;
    layer6_outputs(6315) <= b;
    layer6_outputs(6316) <= not a;
    layer6_outputs(6317) <= a;
    layer6_outputs(6318) <= not a;
    layer6_outputs(6319) <= b;
    layer6_outputs(6320) <= a;
    layer6_outputs(6321) <= a and b;
    layer6_outputs(6322) <= b and not a;
    layer6_outputs(6323) <= not b or a;
    layer6_outputs(6324) <= b;
    layer6_outputs(6325) <= not (a xor b);
    layer6_outputs(6326) <= a and not b;
    layer6_outputs(6327) <= b and not a;
    layer6_outputs(6328) <= a and b;
    layer6_outputs(6329) <= not (a or b);
    layer6_outputs(6330) <= b and not a;
    layer6_outputs(6331) <= not (a or b);
    layer6_outputs(6332) <= not (a xor b);
    layer6_outputs(6333) <= a;
    layer6_outputs(6334) <= not b;
    layer6_outputs(6335) <= not (a or b);
    layer6_outputs(6336) <= not b or a;
    layer6_outputs(6337) <= a;
    layer6_outputs(6338) <= not b;
    layer6_outputs(6339) <= a and b;
    layer6_outputs(6340) <= a and not b;
    layer6_outputs(6341) <= a xor b;
    layer6_outputs(6342) <= a or b;
    layer6_outputs(6343) <= not a;
    layer6_outputs(6344) <= not b;
    layer6_outputs(6345) <= not b;
    layer6_outputs(6346) <= b;
    layer6_outputs(6347) <= a xor b;
    layer6_outputs(6348) <= a or b;
    layer6_outputs(6349) <= a xor b;
    layer6_outputs(6350) <= not b;
    layer6_outputs(6351) <= not a;
    layer6_outputs(6352) <= not a or b;
    layer6_outputs(6353) <= a xor b;
    layer6_outputs(6354) <= '0';
    layer6_outputs(6355) <= a xor b;
    layer6_outputs(6356) <= not a;
    layer6_outputs(6357) <= not a;
    layer6_outputs(6358) <= a or b;
    layer6_outputs(6359) <= not a;
    layer6_outputs(6360) <= not b or a;
    layer6_outputs(6361) <= not a or b;
    layer6_outputs(6362) <= not (a xor b);
    layer6_outputs(6363) <= a;
    layer6_outputs(6364) <= not b or a;
    layer6_outputs(6365) <= not b;
    layer6_outputs(6366) <= not (a xor b);
    layer6_outputs(6367) <= a or b;
    layer6_outputs(6368) <= a and not b;
    layer6_outputs(6369) <= not a;
    layer6_outputs(6370) <= a or b;
    layer6_outputs(6371) <= a xor b;
    layer6_outputs(6372) <= b;
    layer6_outputs(6373) <= a xor b;
    layer6_outputs(6374) <= not b;
    layer6_outputs(6375) <= not b;
    layer6_outputs(6376) <= not a or b;
    layer6_outputs(6377) <= '0';
    layer6_outputs(6378) <= not (a xor b);
    layer6_outputs(6379) <= a and b;
    layer6_outputs(6380) <= b;
    layer6_outputs(6381) <= not (a xor b);
    layer6_outputs(6382) <= not (a and b);
    layer6_outputs(6383) <= not a;
    layer6_outputs(6384) <= a;
    layer6_outputs(6385) <= not b;
    layer6_outputs(6386) <= a xor b;
    layer6_outputs(6387) <= a and not b;
    layer6_outputs(6388) <= not (a xor b);
    layer6_outputs(6389) <= a xor b;
    layer6_outputs(6390) <= not (a and b);
    layer6_outputs(6391) <= a and not b;
    layer6_outputs(6392) <= not a;
    layer6_outputs(6393) <= b;
    layer6_outputs(6394) <= a or b;
    layer6_outputs(6395) <= not (a xor b);
    layer6_outputs(6396) <= not a;
    layer6_outputs(6397) <= not b;
    layer6_outputs(6398) <= a xor b;
    layer6_outputs(6399) <= b;
    layer6_outputs(6400) <= a or b;
    layer6_outputs(6401) <= a and not b;
    layer6_outputs(6402) <= a xor b;
    layer6_outputs(6403) <= b;
    layer6_outputs(6404) <= a xor b;
    layer6_outputs(6405) <= not b or a;
    layer6_outputs(6406) <= a and not b;
    layer6_outputs(6407) <= not a;
    layer6_outputs(6408) <= not (a xor b);
    layer6_outputs(6409) <= a and b;
    layer6_outputs(6410) <= b;
    layer6_outputs(6411) <= not (a and b);
    layer6_outputs(6412) <= not a;
    layer6_outputs(6413) <= a;
    layer6_outputs(6414) <= a and not b;
    layer6_outputs(6415) <= a xor b;
    layer6_outputs(6416) <= b;
    layer6_outputs(6417) <= a;
    layer6_outputs(6418) <= b;
    layer6_outputs(6419) <= a or b;
    layer6_outputs(6420) <= not a;
    layer6_outputs(6421) <= b and not a;
    layer6_outputs(6422) <= not b;
    layer6_outputs(6423) <= not b;
    layer6_outputs(6424) <= not (a or b);
    layer6_outputs(6425) <= not (a or b);
    layer6_outputs(6426) <= not (a xor b);
    layer6_outputs(6427) <= not (a xor b);
    layer6_outputs(6428) <= not (a or b);
    layer6_outputs(6429) <= a;
    layer6_outputs(6430) <= a;
    layer6_outputs(6431) <= not a or b;
    layer6_outputs(6432) <= a;
    layer6_outputs(6433) <= not b;
    layer6_outputs(6434) <= not b or a;
    layer6_outputs(6435) <= not a;
    layer6_outputs(6436) <= not (a and b);
    layer6_outputs(6437) <= not a or b;
    layer6_outputs(6438) <= not a;
    layer6_outputs(6439) <= not a or b;
    layer6_outputs(6440) <= b;
    layer6_outputs(6441) <= not b;
    layer6_outputs(6442) <= not b;
    layer6_outputs(6443) <= not (a xor b);
    layer6_outputs(6444) <= not b;
    layer6_outputs(6445) <= b;
    layer6_outputs(6446) <= b and not a;
    layer6_outputs(6447) <= b;
    layer6_outputs(6448) <= a and not b;
    layer6_outputs(6449) <= not a;
    layer6_outputs(6450) <= b;
    layer6_outputs(6451) <= not b or a;
    layer6_outputs(6452) <= a or b;
    layer6_outputs(6453) <= a xor b;
    layer6_outputs(6454) <= not (a and b);
    layer6_outputs(6455) <= a xor b;
    layer6_outputs(6456) <= a and b;
    layer6_outputs(6457) <= a xor b;
    layer6_outputs(6458) <= not (a xor b);
    layer6_outputs(6459) <= not a or b;
    layer6_outputs(6460) <= b and not a;
    layer6_outputs(6461) <= a xor b;
    layer6_outputs(6462) <= not (a xor b);
    layer6_outputs(6463) <= not (a xor b);
    layer6_outputs(6464) <= not (a xor b);
    layer6_outputs(6465) <= b;
    layer6_outputs(6466) <= not a;
    layer6_outputs(6467) <= not (a and b);
    layer6_outputs(6468) <= a;
    layer6_outputs(6469) <= not b;
    layer6_outputs(6470) <= a and b;
    layer6_outputs(6471) <= not b;
    layer6_outputs(6472) <= not a;
    layer6_outputs(6473) <= a and not b;
    layer6_outputs(6474) <= a xor b;
    layer6_outputs(6475) <= b;
    layer6_outputs(6476) <= b and not a;
    layer6_outputs(6477) <= not a;
    layer6_outputs(6478) <= not b or a;
    layer6_outputs(6479) <= not (a xor b);
    layer6_outputs(6480) <= b;
    layer6_outputs(6481) <= a and b;
    layer6_outputs(6482) <= a or b;
    layer6_outputs(6483) <= a;
    layer6_outputs(6484) <= b;
    layer6_outputs(6485) <= not b;
    layer6_outputs(6486) <= a;
    layer6_outputs(6487) <= not b;
    layer6_outputs(6488) <= a xor b;
    layer6_outputs(6489) <= a and not b;
    layer6_outputs(6490) <= not (a or b);
    layer6_outputs(6491) <= not (a and b);
    layer6_outputs(6492) <= a and b;
    layer6_outputs(6493) <= a xor b;
    layer6_outputs(6494) <= not (a xor b);
    layer6_outputs(6495) <= not (a xor b);
    layer6_outputs(6496) <= not a;
    layer6_outputs(6497) <= not b or a;
    layer6_outputs(6498) <= not a;
    layer6_outputs(6499) <= not a;
    layer6_outputs(6500) <= not (a xor b);
    layer6_outputs(6501) <= a xor b;
    layer6_outputs(6502) <= not (a xor b);
    layer6_outputs(6503) <= b;
    layer6_outputs(6504) <= b;
    layer6_outputs(6505) <= not (a and b);
    layer6_outputs(6506) <= not (a xor b);
    layer6_outputs(6507) <= b;
    layer6_outputs(6508) <= a xor b;
    layer6_outputs(6509) <= b;
    layer6_outputs(6510) <= a xor b;
    layer6_outputs(6511) <= not a;
    layer6_outputs(6512) <= not b;
    layer6_outputs(6513) <= a and not b;
    layer6_outputs(6514) <= a and b;
    layer6_outputs(6515) <= '1';
    layer6_outputs(6516) <= a;
    layer6_outputs(6517) <= b and not a;
    layer6_outputs(6518) <= a and not b;
    layer6_outputs(6519) <= b;
    layer6_outputs(6520) <= not a;
    layer6_outputs(6521) <= a and b;
    layer6_outputs(6522) <= b;
    layer6_outputs(6523) <= a;
    layer6_outputs(6524) <= not (a xor b);
    layer6_outputs(6525) <= not (a or b);
    layer6_outputs(6526) <= not a;
    layer6_outputs(6527) <= not b;
    layer6_outputs(6528) <= a xor b;
    layer6_outputs(6529) <= not a;
    layer6_outputs(6530) <= a xor b;
    layer6_outputs(6531) <= b and not a;
    layer6_outputs(6532) <= not b or a;
    layer6_outputs(6533) <= b and not a;
    layer6_outputs(6534) <= b;
    layer6_outputs(6535) <= a xor b;
    layer6_outputs(6536) <= not b;
    layer6_outputs(6537) <= not (a and b);
    layer6_outputs(6538) <= a or b;
    layer6_outputs(6539) <= not (a or b);
    layer6_outputs(6540) <= b;
    layer6_outputs(6541) <= a;
    layer6_outputs(6542) <= a xor b;
    layer6_outputs(6543) <= a and not b;
    layer6_outputs(6544) <= a;
    layer6_outputs(6545) <= not (a xor b);
    layer6_outputs(6546) <= not a;
    layer6_outputs(6547) <= a xor b;
    layer6_outputs(6548) <= a and not b;
    layer6_outputs(6549) <= b and not a;
    layer6_outputs(6550) <= a;
    layer6_outputs(6551) <= b;
    layer6_outputs(6552) <= not (a or b);
    layer6_outputs(6553) <= not b;
    layer6_outputs(6554) <= a or b;
    layer6_outputs(6555) <= not a;
    layer6_outputs(6556) <= not a or b;
    layer6_outputs(6557) <= not a or b;
    layer6_outputs(6558) <= not a;
    layer6_outputs(6559) <= b;
    layer6_outputs(6560) <= a or b;
    layer6_outputs(6561) <= not b;
    layer6_outputs(6562) <= not a or b;
    layer6_outputs(6563) <= not a or b;
    layer6_outputs(6564) <= a and b;
    layer6_outputs(6565) <= b and not a;
    layer6_outputs(6566) <= not a;
    layer6_outputs(6567) <= not b;
    layer6_outputs(6568) <= b;
    layer6_outputs(6569) <= b;
    layer6_outputs(6570) <= not b or a;
    layer6_outputs(6571) <= not (a and b);
    layer6_outputs(6572) <= not b;
    layer6_outputs(6573) <= a xor b;
    layer6_outputs(6574) <= not (a xor b);
    layer6_outputs(6575) <= not a;
    layer6_outputs(6576) <= not a;
    layer6_outputs(6577) <= not (a xor b);
    layer6_outputs(6578) <= a or b;
    layer6_outputs(6579) <= not (a xor b);
    layer6_outputs(6580) <= '1';
    layer6_outputs(6581) <= a and not b;
    layer6_outputs(6582) <= not a;
    layer6_outputs(6583) <= not b;
    layer6_outputs(6584) <= not (a xor b);
    layer6_outputs(6585) <= not a;
    layer6_outputs(6586) <= not a;
    layer6_outputs(6587) <= a;
    layer6_outputs(6588) <= a;
    layer6_outputs(6589) <= not b;
    layer6_outputs(6590) <= b;
    layer6_outputs(6591) <= not (a xor b);
    layer6_outputs(6592) <= not a;
    layer6_outputs(6593) <= not (a or b);
    layer6_outputs(6594) <= not (a xor b);
    layer6_outputs(6595) <= a and b;
    layer6_outputs(6596) <= a;
    layer6_outputs(6597) <= not (a xor b);
    layer6_outputs(6598) <= not a;
    layer6_outputs(6599) <= not (a xor b);
    layer6_outputs(6600) <= not b;
    layer6_outputs(6601) <= not b;
    layer6_outputs(6602) <= a and b;
    layer6_outputs(6603) <= not (a and b);
    layer6_outputs(6604) <= a;
    layer6_outputs(6605) <= a or b;
    layer6_outputs(6606) <= not (a and b);
    layer6_outputs(6607) <= not a;
    layer6_outputs(6608) <= a or b;
    layer6_outputs(6609) <= a and b;
    layer6_outputs(6610) <= not (a xor b);
    layer6_outputs(6611) <= a;
    layer6_outputs(6612) <= not a;
    layer6_outputs(6613) <= not b;
    layer6_outputs(6614) <= b;
    layer6_outputs(6615) <= a xor b;
    layer6_outputs(6616) <= not a;
    layer6_outputs(6617) <= a or b;
    layer6_outputs(6618) <= a and not b;
    layer6_outputs(6619) <= a;
    layer6_outputs(6620) <= not (a xor b);
    layer6_outputs(6621) <= not a;
    layer6_outputs(6622) <= not b;
    layer6_outputs(6623) <= a xor b;
    layer6_outputs(6624) <= not b;
    layer6_outputs(6625) <= a or b;
    layer6_outputs(6626) <= not (a xor b);
    layer6_outputs(6627) <= not a;
    layer6_outputs(6628) <= a and b;
    layer6_outputs(6629) <= not b or a;
    layer6_outputs(6630) <= not a;
    layer6_outputs(6631) <= a and not b;
    layer6_outputs(6632) <= a and b;
    layer6_outputs(6633) <= a and b;
    layer6_outputs(6634) <= a and not b;
    layer6_outputs(6635) <= a;
    layer6_outputs(6636) <= b and not a;
    layer6_outputs(6637) <= a;
    layer6_outputs(6638) <= a;
    layer6_outputs(6639) <= a;
    layer6_outputs(6640) <= b;
    layer6_outputs(6641) <= a xor b;
    layer6_outputs(6642) <= a or b;
    layer6_outputs(6643) <= not (a xor b);
    layer6_outputs(6644) <= a or b;
    layer6_outputs(6645) <= a xor b;
    layer6_outputs(6646) <= not b;
    layer6_outputs(6647) <= not a;
    layer6_outputs(6648) <= not a;
    layer6_outputs(6649) <= a and b;
    layer6_outputs(6650) <= not b or a;
    layer6_outputs(6651) <= not a;
    layer6_outputs(6652) <= not a;
    layer6_outputs(6653) <= not a;
    layer6_outputs(6654) <= not (a or b);
    layer6_outputs(6655) <= b;
    layer6_outputs(6656) <= not b or a;
    layer6_outputs(6657) <= not (a xor b);
    layer6_outputs(6658) <= not a;
    layer6_outputs(6659) <= b and not a;
    layer6_outputs(6660) <= b and not a;
    layer6_outputs(6661) <= not (a xor b);
    layer6_outputs(6662) <= not b;
    layer6_outputs(6663) <= a and b;
    layer6_outputs(6664) <= a xor b;
    layer6_outputs(6665) <= not b;
    layer6_outputs(6666) <= not b;
    layer6_outputs(6667) <= a xor b;
    layer6_outputs(6668) <= not b;
    layer6_outputs(6669) <= not (a xor b);
    layer6_outputs(6670) <= not a or b;
    layer6_outputs(6671) <= a and not b;
    layer6_outputs(6672) <= a or b;
    layer6_outputs(6673) <= b;
    layer6_outputs(6674) <= a and b;
    layer6_outputs(6675) <= not (a xor b);
    layer6_outputs(6676) <= not b or a;
    layer6_outputs(6677) <= a xor b;
    layer6_outputs(6678) <= not (a xor b);
    layer6_outputs(6679) <= a;
    layer6_outputs(6680) <= a;
    layer6_outputs(6681) <= not b or a;
    layer6_outputs(6682) <= a;
    layer6_outputs(6683) <= a xor b;
    layer6_outputs(6684) <= b;
    layer6_outputs(6685) <= not a;
    layer6_outputs(6686) <= a or b;
    layer6_outputs(6687) <= a and not b;
    layer6_outputs(6688) <= not a or b;
    layer6_outputs(6689) <= a;
    layer6_outputs(6690) <= not b;
    layer6_outputs(6691) <= a or b;
    layer6_outputs(6692) <= not (a and b);
    layer6_outputs(6693) <= b and not a;
    layer6_outputs(6694) <= not a;
    layer6_outputs(6695) <= b;
    layer6_outputs(6696) <= not (a xor b);
    layer6_outputs(6697) <= not (a and b);
    layer6_outputs(6698) <= not b;
    layer6_outputs(6699) <= not (a xor b);
    layer6_outputs(6700) <= a xor b;
    layer6_outputs(6701) <= not b;
    layer6_outputs(6702) <= a;
    layer6_outputs(6703) <= b;
    layer6_outputs(6704) <= b;
    layer6_outputs(6705) <= a and not b;
    layer6_outputs(6706) <= b;
    layer6_outputs(6707) <= not a;
    layer6_outputs(6708) <= a and b;
    layer6_outputs(6709) <= b and not a;
    layer6_outputs(6710) <= a xor b;
    layer6_outputs(6711) <= not (a xor b);
    layer6_outputs(6712) <= b;
    layer6_outputs(6713) <= not b;
    layer6_outputs(6714) <= a xor b;
    layer6_outputs(6715) <= b and not a;
    layer6_outputs(6716) <= not b or a;
    layer6_outputs(6717) <= not a;
    layer6_outputs(6718) <= a and not b;
    layer6_outputs(6719) <= b;
    layer6_outputs(6720) <= '0';
    layer6_outputs(6721) <= b;
    layer6_outputs(6722) <= not a;
    layer6_outputs(6723) <= b and not a;
    layer6_outputs(6724) <= not a;
    layer6_outputs(6725) <= b;
    layer6_outputs(6726) <= not a;
    layer6_outputs(6727) <= not a or b;
    layer6_outputs(6728) <= not b;
    layer6_outputs(6729) <= not (a xor b);
    layer6_outputs(6730) <= not b;
    layer6_outputs(6731) <= not a or b;
    layer6_outputs(6732) <= not (a xor b);
    layer6_outputs(6733) <= a and b;
    layer6_outputs(6734) <= b;
    layer6_outputs(6735) <= not b;
    layer6_outputs(6736) <= not a;
    layer6_outputs(6737) <= a xor b;
    layer6_outputs(6738) <= not a;
    layer6_outputs(6739) <= not a;
    layer6_outputs(6740) <= not (a xor b);
    layer6_outputs(6741) <= b and not a;
    layer6_outputs(6742) <= a xor b;
    layer6_outputs(6743) <= not (a and b);
    layer6_outputs(6744) <= a;
    layer6_outputs(6745) <= a;
    layer6_outputs(6746) <= not a or b;
    layer6_outputs(6747) <= not b;
    layer6_outputs(6748) <= a xor b;
    layer6_outputs(6749) <= not a or b;
    layer6_outputs(6750) <= not a;
    layer6_outputs(6751) <= not (a xor b);
    layer6_outputs(6752) <= not (a and b);
    layer6_outputs(6753) <= a or b;
    layer6_outputs(6754) <= a xor b;
    layer6_outputs(6755) <= a xor b;
    layer6_outputs(6756) <= not b;
    layer6_outputs(6757) <= not (a xor b);
    layer6_outputs(6758) <= not a;
    layer6_outputs(6759) <= a and not b;
    layer6_outputs(6760) <= not b;
    layer6_outputs(6761) <= not a or b;
    layer6_outputs(6762) <= not (a and b);
    layer6_outputs(6763) <= a and not b;
    layer6_outputs(6764) <= not a;
    layer6_outputs(6765) <= not b;
    layer6_outputs(6766) <= not b or a;
    layer6_outputs(6767) <= not b;
    layer6_outputs(6768) <= a and b;
    layer6_outputs(6769) <= a or b;
    layer6_outputs(6770) <= not a or b;
    layer6_outputs(6771) <= not b;
    layer6_outputs(6772) <= a and b;
    layer6_outputs(6773) <= b;
    layer6_outputs(6774) <= b;
    layer6_outputs(6775) <= a and b;
    layer6_outputs(6776) <= b;
    layer6_outputs(6777) <= not (a xor b);
    layer6_outputs(6778) <= not (a or b);
    layer6_outputs(6779) <= not b;
    layer6_outputs(6780) <= a and b;
    layer6_outputs(6781) <= a;
    layer6_outputs(6782) <= b;
    layer6_outputs(6783) <= a or b;
    layer6_outputs(6784) <= b;
    layer6_outputs(6785) <= not b or a;
    layer6_outputs(6786) <= not (a and b);
    layer6_outputs(6787) <= not a or b;
    layer6_outputs(6788) <= not a;
    layer6_outputs(6789) <= not b;
    layer6_outputs(6790) <= a xor b;
    layer6_outputs(6791) <= '0';
    layer6_outputs(6792) <= a xor b;
    layer6_outputs(6793) <= b;
    layer6_outputs(6794) <= b;
    layer6_outputs(6795) <= '1';
    layer6_outputs(6796) <= a or b;
    layer6_outputs(6797) <= a or b;
    layer6_outputs(6798) <= a;
    layer6_outputs(6799) <= not a or b;
    layer6_outputs(6800) <= a and b;
    layer6_outputs(6801) <= not b;
    layer6_outputs(6802) <= not a;
    layer6_outputs(6803) <= not b or a;
    layer6_outputs(6804) <= a;
    layer6_outputs(6805) <= a or b;
    layer6_outputs(6806) <= b and not a;
    layer6_outputs(6807) <= b;
    layer6_outputs(6808) <= b;
    layer6_outputs(6809) <= not a;
    layer6_outputs(6810) <= b and not a;
    layer6_outputs(6811) <= not (a and b);
    layer6_outputs(6812) <= a and not b;
    layer6_outputs(6813) <= not b;
    layer6_outputs(6814) <= a and b;
    layer6_outputs(6815) <= a and not b;
    layer6_outputs(6816) <= not (a xor b);
    layer6_outputs(6817) <= not a;
    layer6_outputs(6818) <= a;
    layer6_outputs(6819) <= not b;
    layer6_outputs(6820) <= a and not b;
    layer6_outputs(6821) <= not (a xor b);
    layer6_outputs(6822) <= not (a xor b);
    layer6_outputs(6823) <= not b;
    layer6_outputs(6824) <= not b or a;
    layer6_outputs(6825) <= not b;
    layer6_outputs(6826) <= a;
    layer6_outputs(6827) <= not (a or b);
    layer6_outputs(6828) <= not (a or b);
    layer6_outputs(6829) <= b;
    layer6_outputs(6830) <= not (a xor b);
    layer6_outputs(6831) <= a and b;
    layer6_outputs(6832) <= b;
    layer6_outputs(6833) <= a or b;
    layer6_outputs(6834) <= a xor b;
    layer6_outputs(6835) <= a and not b;
    layer6_outputs(6836) <= not (a xor b);
    layer6_outputs(6837) <= not (a xor b);
    layer6_outputs(6838) <= a or b;
    layer6_outputs(6839) <= not a or b;
    layer6_outputs(6840) <= a xor b;
    layer6_outputs(6841) <= a and b;
    layer6_outputs(6842) <= not (a or b);
    layer6_outputs(6843) <= b;
    layer6_outputs(6844) <= b;
    layer6_outputs(6845) <= b;
    layer6_outputs(6846) <= a xor b;
    layer6_outputs(6847) <= not (a xor b);
    layer6_outputs(6848) <= b and not a;
    layer6_outputs(6849) <= a;
    layer6_outputs(6850) <= not (a and b);
    layer6_outputs(6851) <= a xor b;
    layer6_outputs(6852) <= b;
    layer6_outputs(6853) <= not a;
    layer6_outputs(6854) <= b;
    layer6_outputs(6855) <= a xor b;
    layer6_outputs(6856) <= not b;
    layer6_outputs(6857) <= a xor b;
    layer6_outputs(6858) <= not b or a;
    layer6_outputs(6859) <= b;
    layer6_outputs(6860) <= '1';
    layer6_outputs(6861) <= not b or a;
    layer6_outputs(6862) <= b;
    layer6_outputs(6863) <= not b;
    layer6_outputs(6864) <= a or b;
    layer6_outputs(6865) <= a;
    layer6_outputs(6866) <= not (a or b);
    layer6_outputs(6867) <= a and b;
    layer6_outputs(6868) <= not (a or b);
    layer6_outputs(6869) <= not (a or b);
    layer6_outputs(6870) <= b;
    layer6_outputs(6871) <= not a;
    layer6_outputs(6872) <= not a;
    layer6_outputs(6873) <= not (a xor b);
    layer6_outputs(6874) <= not (a xor b);
    layer6_outputs(6875) <= a or b;
    layer6_outputs(6876) <= not (a and b);
    layer6_outputs(6877) <= a and b;
    layer6_outputs(6878) <= not b;
    layer6_outputs(6879) <= a or b;
    layer6_outputs(6880) <= not (a xor b);
    layer6_outputs(6881) <= not b or a;
    layer6_outputs(6882) <= not a;
    layer6_outputs(6883) <= a or b;
    layer6_outputs(6884) <= not (a xor b);
    layer6_outputs(6885) <= a xor b;
    layer6_outputs(6886) <= a xor b;
    layer6_outputs(6887) <= not a;
    layer6_outputs(6888) <= a xor b;
    layer6_outputs(6889) <= not a;
    layer6_outputs(6890) <= a xor b;
    layer6_outputs(6891) <= not (a xor b);
    layer6_outputs(6892) <= a or b;
    layer6_outputs(6893) <= not a or b;
    layer6_outputs(6894) <= a and not b;
    layer6_outputs(6895) <= not b;
    layer6_outputs(6896) <= a xor b;
    layer6_outputs(6897) <= not a;
    layer6_outputs(6898) <= not b or a;
    layer6_outputs(6899) <= not b;
    layer6_outputs(6900) <= not (a xor b);
    layer6_outputs(6901) <= a;
    layer6_outputs(6902) <= not (a xor b);
    layer6_outputs(6903) <= not (a xor b);
    layer6_outputs(6904) <= not (a xor b);
    layer6_outputs(6905) <= a and not b;
    layer6_outputs(6906) <= not (a or b);
    layer6_outputs(6907) <= not a;
    layer6_outputs(6908) <= not b;
    layer6_outputs(6909) <= a or b;
    layer6_outputs(6910) <= not (a xor b);
    layer6_outputs(6911) <= a and b;
    layer6_outputs(6912) <= a and b;
    layer6_outputs(6913) <= not b;
    layer6_outputs(6914) <= not b;
    layer6_outputs(6915) <= not b;
    layer6_outputs(6916) <= b;
    layer6_outputs(6917) <= a and not b;
    layer6_outputs(6918) <= not (a xor b);
    layer6_outputs(6919) <= b;
    layer6_outputs(6920) <= not a;
    layer6_outputs(6921) <= a xor b;
    layer6_outputs(6922) <= not (a xor b);
    layer6_outputs(6923) <= a and b;
    layer6_outputs(6924) <= not a;
    layer6_outputs(6925) <= not (a xor b);
    layer6_outputs(6926) <= b;
    layer6_outputs(6927) <= not b;
    layer6_outputs(6928) <= not a;
    layer6_outputs(6929) <= not b or a;
    layer6_outputs(6930) <= not (a xor b);
    layer6_outputs(6931) <= a and b;
    layer6_outputs(6932) <= not a or b;
    layer6_outputs(6933) <= not a or b;
    layer6_outputs(6934) <= b and not a;
    layer6_outputs(6935) <= not b;
    layer6_outputs(6936) <= a or b;
    layer6_outputs(6937) <= not a;
    layer6_outputs(6938) <= b;
    layer6_outputs(6939) <= a or b;
    layer6_outputs(6940) <= a;
    layer6_outputs(6941) <= not b or a;
    layer6_outputs(6942) <= not b;
    layer6_outputs(6943) <= not (a or b);
    layer6_outputs(6944) <= not (a or b);
    layer6_outputs(6945) <= not a;
    layer6_outputs(6946) <= not (a xor b);
    layer6_outputs(6947) <= not a;
    layer6_outputs(6948) <= not b;
    layer6_outputs(6949) <= a xor b;
    layer6_outputs(6950) <= not (a xor b);
    layer6_outputs(6951) <= not (a xor b);
    layer6_outputs(6952) <= not a or b;
    layer6_outputs(6953) <= a;
    layer6_outputs(6954) <= a xor b;
    layer6_outputs(6955) <= not (a or b);
    layer6_outputs(6956) <= a;
    layer6_outputs(6957) <= a;
    layer6_outputs(6958) <= a xor b;
    layer6_outputs(6959) <= a and not b;
    layer6_outputs(6960) <= a xor b;
    layer6_outputs(6961) <= a xor b;
    layer6_outputs(6962) <= b and not a;
    layer6_outputs(6963) <= '0';
    layer6_outputs(6964) <= not (a xor b);
    layer6_outputs(6965) <= not a or b;
    layer6_outputs(6966) <= a and not b;
    layer6_outputs(6967) <= not a or b;
    layer6_outputs(6968) <= b and not a;
    layer6_outputs(6969) <= not (a xor b);
    layer6_outputs(6970) <= a and b;
    layer6_outputs(6971) <= a;
    layer6_outputs(6972) <= not b or a;
    layer6_outputs(6973) <= not (a xor b);
    layer6_outputs(6974) <= not (a xor b);
    layer6_outputs(6975) <= b;
    layer6_outputs(6976) <= not (a or b);
    layer6_outputs(6977) <= b and not a;
    layer6_outputs(6978) <= not b or a;
    layer6_outputs(6979) <= b;
    layer6_outputs(6980) <= not a or b;
    layer6_outputs(6981) <= a;
    layer6_outputs(6982) <= not (a xor b);
    layer6_outputs(6983) <= not a;
    layer6_outputs(6984) <= b and not a;
    layer6_outputs(6985) <= a and not b;
    layer6_outputs(6986) <= not (a xor b);
    layer6_outputs(6987) <= a xor b;
    layer6_outputs(6988) <= not (a xor b);
    layer6_outputs(6989) <= not a;
    layer6_outputs(6990) <= a;
    layer6_outputs(6991) <= b;
    layer6_outputs(6992) <= a xor b;
    layer6_outputs(6993) <= a xor b;
    layer6_outputs(6994) <= a xor b;
    layer6_outputs(6995) <= b;
    layer6_outputs(6996) <= not (a xor b);
    layer6_outputs(6997) <= not b;
    layer6_outputs(6998) <= not (a or b);
    layer6_outputs(6999) <= not a or b;
    layer6_outputs(7000) <= a xor b;
    layer6_outputs(7001) <= not (a and b);
    layer6_outputs(7002) <= not a or b;
    layer6_outputs(7003) <= b;
    layer6_outputs(7004) <= not a;
    layer6_outputs(7005) <= not b or a;
    layer6_outputs(7006) <= b and not a;
    layer6_outputs(7007) <= not a or b;
    layer6_outputs(7008) <= not b or a;
    layer6_outputs(7009) <= a xor b;
    layer6_outputs(7010) <= not b or a;
    layer6_outputs(7011) <= not a or b;
    layer6_outputs(7012) <= not b;
    layer6_outputs(7013) <= a;
    layer6_outputs(7014) <= not b;
    layer6_outputs(7015) <= not (a xor b);
    layer6_outputs(7016) <= a xor b;
    layer6_outputs(7017) <= a;
    layer6_outputs(7018) <= not (a xor b);
    layer6_outputs(7019) <= a and not b;
    layer6_outputs(7020) <= not (a and b);
    layer6_outputs(7021) <= not (a or b);
    layer6_outputs(7022) <= not (a xor b);
    layer6_outputs(7023) <= a or b;
    layer6_outputs(7024) <= not b or a;
    layer6_outputs(7025) <= b;
    layer6_outputs(7026) <= a or b;
    layer6_outputs(7027) <= not a or b;
    layer6_outputs(7028) <= b;
    layer6_outputs(7029) <= not a;
    layer6_outputs(7030) <= not b;
    layer6_outputs(7031) <= a and not b;
    layer6_outputs(7032) <= not (a xor b);
    layer6_outputs(7033) <= a;
    layer6_outputs(7034) <= not b;
    layer6_outputs(7035) <= not b;
    layer6_outputs(7036) <= a xor b;
    layer6_outputs(7037) <= a;
    layer6_outputs(7038) <= not (a or b);
    layer6_outputs(7039) <= not (a xor b);
    layer6_outputs(7040) <= not a or b;
    layer6_outputs(7041) <= a xor b;
    layer6_outputs(7042) <= not (a xor b);
    layer6_outputs(7043) <= not (a or b);
    layer6_outputs(7044) <= b and not a;
    layer6_outputs(7045) <= not b or a;
    layer6_outputs(7046) <= b and not a;
    layer6_outputs(7047) <= not b;
    layer6_outputs(7048) <= not a or b;
    layer6_outputs(7049) <= not a;
    layer6_outputs(7050) <= '0';
    layer6_outputs(7051) <= a xor b;
    layer6_outputs(7052) <= not a;
    layer6_outputs(7053) <= a xor b;
    layer6_outputs(7054) <= b;
    layer6_outputs(7055) <= not a;
    layer6_outputs(7056) <= a xor b;
    layer6_outputs(7057) <= a;
    layer6_outputs(7058) <= not a;
    layer6_outputs(7059) <= not a;
    layer6_outputs(7060) <= not a;
    layer6_outputs(7061) <= not a;
    layer6_outputs(7062) <= a;
    layer6_outputs(7063) <= not b;
    layer6_outputs(7064) <= a and b;
    layer6_outputs(7065) <= a and b;
    layer6_outputs(7066) <= not (a xor b);
    layer6_outputs(7067) <= b;
    layer6_outputs(7068) <= not a;
    layer6_outputs(7069) <= a and not b;
    layer6_outputs(7070) <= a and b;
    layer6_outputs(7071) <= not a;
    layer6_outputs(7072) <= b;
    layer6_outputs(7073) <= not a;
    layer6_outputs(7074) <= not b;
    layer6_outputs(7075) <= not (a xor b);
    layer6_outputs(7076) <= not (a xor b);
    layer6_outputs(7077) <= b;
    layer6_outputs(7078) <= b;
    layer6_outputs(7079) <= not b;
    layer6_outputs(7080) <= a xor b;
    layer6_outputs(7081) <= a or b;
    layer6_outputs(7082) <= b and not a;
    layer6_outputs(7083) <= not b or a;
    layer6_outputs(7084) <= not b or a;
    layer6_outputs(7085) <= a;
    layer6_outputs(7086) <= not (a or b);
    layer6_outputs(7087) <= not b or a;
    layer6_outputs(7088) <= a;
    layer6_outputs(7089) <= not a;
    layer6_outputs(7090) <= b and not a;
    layer6_outputs(7091) <= not b;
    layer6_outputs(7092) <= a and b;
    layer6_outputs(7093) <= a;
    layer6_outputs(7094) <= not a or b;
    layer6_outputs(7095) <= not a;
    layer6_outputs(7096) <= a;
    layer6_outputs(7097) <= not b;
    layer6_outputs(7098) <= b and not a;
    layer6_outputs(7099) <= a xor b;
    layer6_outputs(7100) <= b and not a;
    layer6_outputs(7101) <= not (a and b);
    layer6_outputs(7102) <= a;
    layer6_outputs(7103) <= not b;
    layer6_outputs(7104) <= b;
    layer6_outputs(7105) <= a xor b;
    layer6_outputs(7106) <= a and b;
    layer6_outputs(7107) <= not a;
    layer6_outputs(7108) <= not a;
    layer6_outputs(7109) <= a xor b;
    layer6_outputs(7110) <= not a;
    layer6_outputs(7111) <= not (a and b);
    layer6_outputs(7112) <= a;
    layer6_outputs(7113) <= not a or b;
    layer6_outputs(7114) <= not b;
    layer6_outputs(7115) <= a xor b;
    layer6_outputs(7116) <= a xor b;
    layer6_outputs(7117) <= not b;
    layer6_outputs(7118) <= a xor b;
    layer6_outputs(7119) <= a and b;
    layer6_outputs(7120) <= a;
    layer6_outputs(7121) <= a and not b;
    layer6_outputs(7122) <= not (a and b);
    layer6_outputs(7123) <= a;
    layer6_outputs(7124) <= a;
    layer6_outputs(7125) <= a;
    layer6_outputs(7126) <= not (a xor b);
    layer6_outputs(7127) <= b;
    layer6_outputs(7128) <= b;
    layer6_outputs(7129) <= a xor b;
    layer6_outputs(7130) <= a and b;
    layer6_outputs(7131) <= b;
    layer6_outputs(7132) <= not (a and b);
    layer6_outputs(7133) <= not (a and b);
    layer6_outputs(7134) <= a;
    layer6_outputs(7135) <= not (a xor b);
    layer6_outputs(7136) <= a or b;
    layer6_outputs(7137) <= not (a or b);
    layer6_outputs(7138) <= not b;
    layer6_outputs(7139) <= a xor b;
    layer6_outputs(7140) <= not b;
    layer6_outputs(7141) <= not a or b;
    layer6_outputs(7142) <= a;
    layer6_outputs(7143) <= not b;
    layer6_outputs(7144) <= not (a and b);
    layer6_outputs(7145) <= b and not a;
    layer6_outputs(7146) <= not a;
    layer6_outputs(7147) <= not a;
    layer6_outputs(7148) <= a;
    layer6_outputs(7149) <= not (a xor b);
    layer6_outputs(7150) <= not a;
    layer6_outputs(7151) <= a xor b;
    layer6_outputs(7152) <= b;
    layer6_outputs(7153) <= not b or a;
    layer6_outputs(7154) <= a;
    layer6_outputs(7155) <= b;
    layer6_outputs(7156) <= a xor b;
    layer6_outputs(7157) <= a xor b;
    layer6_outputs(7158) <= not a;
    layer6_outputs(7159) <= a;
    layer6_outputs(7160) <= a and not b;
    layer6_outputs(7161) <= a xor b;
    layer6_outputs(7162) <= a;
    layer6_outputs(7163) <= a;
    layer6_outputs(7164) <= not a or b;
    layer6_outputs(7165) <= not b;
    layer6_outputs(7166) <= not a;
    layer6_outputs(7167) <= not a or b;
    layer6_outputs(7168) <= not b;
    layer6_outputs(7169) <= not b;
    layer6_outputs(7170) <= a xor b;
    layer6_outputs(7171) <= b;
    layer6_outputs(7172) <= a xor b;
    layer6_outputs(7173) <= not b;
    layer6_outputs(7174) <= a xor b;
    layer6_outputs(7175) <= not b;
    layer6_outputs(7176) <= b;
    layer6_outputs(7177) <= not (a xor b);
    layer6_outputs(7178) <= a xor b;
    layer6_outputs(7179) <= a or b;
    layer6_outputs(7180) <= not (a xor b);
    layer6_outputs(7181) <= not (a xor b);
    layer6_outputs(7182) <= not b;
    layer6_outputs(7183) <= a;
    layer6_outputs(7184) <= not (a xor b);
    layer6_outputs(7185) <= not a;
    layer6_outputs(7186) <= not b;
    layer6_outputs(7187) <= b;
    layer6_outputs(7188) <= a xor b;
    layer6_outputs(7189) <= b;
    layer6_outputs(7190) <= not a;
    layer6_outputs(7191) <= a and not b;
    layer6_outputs(7192) <= a xor b;
    layer6_outputs(7193) <= not a or b;
    layer6_outputs(7194) <= not a;
    layer6_outputs(7195) <= not b;
    layer6_outputs(7196) <= a and b;
    layer6_outputs(7197) <= not a;
    layer6_outputs(7198) <= not b;
    layer6_outputs(7199) <= not b;
    layer6_outputs(7200) <= b;
    layer6_outputs(7201) <= a or b;
    layer6_outputs(7202) <= a;
    layer6_outputs(7203) <= a xor b;
    layer6_outputs(7204) <= not a or b;
    layer6_outputs(7205) <= not (a xor b);
    layer6_outputs(7206) <= b and not a;
    layer6_outputs(7207) <= a xor b;
    layer6_outputs(7208) <= a;
    layer6_outputs(7209) <= not b;
    layer6_outputs(7210) <= not a or b;
    layer6_outputs(7211) <= not (a or b);
    layer6_outputs(7212) <= not (a and b);
    layer6_outputs(7213) <= a or b;
    layer6_outputs(7214) <= not b;
    layer6_outputs(7215) <= not a;
    layer6_outputs(7216) <= b and not a;
    layer6_outputs(7217) <= b;
    layer6_outputs(7218) <= not (a xor b);
    layer6_outputs(7219) <= not (a or b);
    layer6_outputs(7220) <= not (a and b);
    layer6_outputs(7221) <= b;
    layer6_outputs(7222) <= a or b;
    layer6_outputs(7223) <= not a or b;
    layer6_outputs(7224) <= a;
    layer6_outputs(7225) <= a or b;
    layer6_outputs(7226) <= not b;
    layer6_outputs(7227) <= not (a or b);
    layer6_outputs(7228) <= a xor b;
    layer6_outputs(7229) <= not (a or b);
    layer6_outputs(7230) <= b;
    layer6_outputs(7231) <= a xor b;
    layer6_outputs(7232) <= a and not b;
    layer6_outputs(7233) <= a xor b;
    layer6_outputs(7234) <= b;
    layer6_outputs(7235) <= a or b;
    layer6_outputs(7236) <= not b or a;
    layer6_outputs(7237) <= not a or b;
    layer6_outputs(7238) <= a xor b;
    layer6_outputs(7239) <= not a or b;
    layer6_outputs(7240) <= not (a xor b);
    layer6_outputs(7241) <= not (a and b);
    layer6_outputs(7242) <= not a;
    layer6_outputs(7243) <= not (a xor b);
    layer6_outputs(7244) <= b and not a;
    layer6_outputs(7245) <= '1';
    layer6_outputs(7246) <= not a;
    layer6_outputs(7247) <= a and b;
    layer6_outputs(7248) <= not (a xor b);
    layer6_outputs(7249) <= b;
    layer6_outputs(7250) <= a and not b;
    layer6_outputs(7251) <= b;
    layer6_outputs(7252) <= b;
    layer6_outputs(7253) <= b;
    layer6_outputs(7254) <= not a;
    layer6_outputs(7255) <= not (a xor b);
    layer6_outputs(7256) <= not (a xor b);
    layer6_outputs(7257) <= not a;
    layer6_outputs(7258) <= a xor b;
    layer6_outputs(7259) <= a;
    layer6_outputs(7260) <= not a;
    layer6_outputs(7261) <= a;
    layer6_outputs(7262) <= a or b;
    layer6_outputs(7263) <= b and not a;
    layer6_outputs(7264) <= not a;
    layer6_outputs(7265) <= not a;
    layer6_outputs(7266) <= not (a xor b);
    layer6_outputs(7267) <= b;
    layer6_outputs(7268) <= not a or b;
    layer6_outputs(7269) <= a xor b;
    layer6_outputs(7270) <= a and not b;
    layer6_outputs(7271) <= not a;
    layer6_outputs(7272) <= not b or a;
    layer6_outputs(7273) <= a or b;
    layer6_outputs(7274) <= a and not b;
    layer6_outputs(7275) <= a xor b;
    layer6_outputs(7276) <= not a or b;
    layer6_outputs(7277) <= a;
    layer6_outputs(7278) <= b;
    layer6_outputs(7279) <= not b;
    layer6_outputs(7280) <= not a;
    layer6_outputs(7281) <= b;
    layer6_outputs(7282) <= a or b;
    layer6_outputs(7283) <= b;
    layer6_outputs(7284) <= b;
    layer6_outputs(7285) <= a and b;
    layer6_outputs(7286) <= a xor b;
    layer6_outputs(7287) <= not b;
    layer6_outputs(7288) <= b;
    layer6_outputs(7289) <= not a;
    layer6_outputs(7290) <= a xor b;
    layer6_outputs(7291) <= a;
    layer6_outputs(7292) <= not b;
    layer6_outputs(7293) <= a xor b;
    layer6_outputs(7294) <= a xor b;
    layer6_outputs(7295) <= not b;
    layer6_outputs(7296) <= not b;
    layer6_outputs(7297) <= a;
    layer6_outputs(7298) <= a and b;
    layer6_outputs(7299) <= not a;
    layer6_outputs(7300) <= a or b;
    layer6_outputs(7301) <= not (a or b);
    layer6_outputs(7302) <= a and b;
    layer6_outputs(7303) <= not a;
    layer6_outputs(7304) <= a xor b;
    layer6_outputs(7305) <= not a;
    layer6_outputs(7306) <= not (a xor b);
    layer6_outputs(7307) <= a;
    layer6_outputs(7308) <= not b;
    layer6_outputs(7309) <= a;
    layer6_outputs(7310) <= a and not b;
    layer6_outputs(7311) <= a;
    layer6_outputs(7312) <= not a;
    layer6_outputs(7313) <= a xor b;
    layer6_outputs(7314) <= not (a and b);
    layer6_outputs(7315) <= a and b;
    layer6_outputs(7316) <= '1';
    layer6_outputs(7317) <= not (a and b);
    layer6_outputs(7318) <= not a;
    layer6_outputs(7319) <= b;
    layer6_outputs(7320) <= a;
    layer6_outputs(7321) <= b;
    layer6_outputs(7322) <= not (a or b);
    layer6_outputs(7323) <= a;
    layer6_outputs(7324) <= a;
    layer6_outputs(7325) <= not a;
    layer6_outputs(7326) <= a;
    layer6_outputs(7327) <= b;
    layer6_outputs(7328) <= not a;
    layer6_outputs(7329) <= not b or a;
    layer6_outputs(7330) <= not a;
    layer6_outputs(7331) <= a xor b;
    layer6_outputs(7332) <= b;
    layer6_outputs(7333) <= not b;
    layer6_outputs(7334) <= a;
    layer6_outputs(7335) <= not (a xor b);
    layer6_outputs(7336) <= not a or b;
    layer6_outputs(7337) <= not a;
    layer6_outputs(7338) <= b and not a;
    layer6_outputs(7339) <= b;
    layer6_outputs(7340) <= a;
    layer6_outputs(7341) <= not b;
    layer6_outputs(7342) <= a;
    layer6_outputs(7343) <= a xor b;
    layer6_outputs(7344) <= a xor b;
    layer6_outputs(7345) <= not b;
    layer6_outputs(7346) <= a;
    layer6_outputs(7347) <= not (a and b);
    layer6_outputs(7348) <= b and not a;
    layer6_outputs(7349) <= a and b;
    layer6_outputs(7350) <= a xor b;
    layer6_outputs(7351) <= b and not a;
    layer6_outputs(7352) <= not b;
    layer6_outputs(7353) <= b;
    layer6_outputs(7354) <= b;
    layer6_outputs(7355) <= a and not b;
    layer6_outputs(7356) <= not (a xor b);
    layer6_outputs(7357) <= not a;
    layer6_outputs(7358) <= a;
    layer6_outputs(7359) <= a or b;
    layer6_outputs(7360) <= not a;
    layer6_outputs(7361) <= not b;
    layer6_outputs(7362) <= not a or b;
    layer6_outputs(7363) <= a and not b;
    layer6_outputs(7364) <= not a;
    layer6_outputs(7365) <= not (a and b);
    layer6_outputs(7366) <= a;
    layer6_outputs(7367) <= not b;
    layer6_outputs(7368) <= a;
    layer6_outputs(7369) <= not b;
    layer6_outputs(7370) <= a;
    layer6_outputs(7371) <= not (a and b);
    layer6_outputs(7372) <= a xor b;
    layer6_outputs(7373) <= not b;
    layer6_outputs(7374) <= not a or b;
    layer6_outputs(7375) <= a and not b;
    layer6_outputs(7376) <= not b;
    layer6_outputs(7377) <= not b or a;
    layer6_outputs(7378) <= not b;
    layer6_outputs(7379) <= a xor b;
    layer6_outputs(7380) <= not a or b;
    layer6_outputs(7381) <= a xor b;
    layer6_outputs(7382) <= a and not b;
    layer6_outputs(7383) <= not b;
    layer6_outputs(7384) <= not (a or b);
    layer6_outputs(7385) <= b and not a;
    layer6_outputs(7386) <= b;
    layer6_outputs(7387) <= not a;
    layer6_outputs(7388) <= not a;
    layer6_outputs(7389) <= a and b;
    layer6_outputs(7390) <= a or b;
    layer6_outputs(7391) <= not (a and b);
    layer6_outputs(7392) <= a;
    layer6_outputs(7393) <= not b;
    layer6_outputs(7394) <= not b or a;
    layer6_outputs(7395) <= a;
    layer6_outputs(7396) <= b;
    layer6_outputs(7397) <= a xor b;
    layer6_outputs(7398) <= a and not b;
    layer6_outputs(7399) <= a or b;
    layer6_outputs(7400) <= not b;
    layer6_outputs(7401) <= a and b;
    layer6_outputs(7402) <= a and b;
    layer6_outputs(7403) <= a or b;
    layer6_outputs(7404) <= a;
    layer6_outputs(7405) <= not (a or b);
    layer6_outputs(7406) <= not (a xor b);
    layer6_outputs(7407) <= not a or b;
    layer6_outputs(7408) <= a or b;
    layer6_outputs(7409) <= not a or b;
    layer6_outputs(7410) <= b;
    layer6_outputs(7411) <= b and not a;
    layer6_outputs(7412) <= not (a xor b);
    layer6_outputs(7413) <= b;
    layer6_outputs(7414) <= not b;
    layer6_outputs(7415) <= b and not a;
    layer6_outputs(7416) <= not (a xor b);
    layer6_outputs(7417) <= b and not a;
    layer6_outputs(7418) <= not (a xor b);
    layer6_outputs(7419) <= a or b;
    layer6_outputs(7420) <= a and b;
    layer6_outputs(7421) <= b;
    layer6_outputs(7422) <= a;
    layer6_outputs(7423) <= b and not a;
    layer6_outputs(7424) <= not a or b;
    layer6_outputs(7425) <= b;
    layer6_outputs(7426) <= not b or a;
    layer6_outputs(7427) <= not (a and b);
    layer6_outputs(7428) <= not (a and b);
    layer6_outputs(7429) <= a xor b;
    layer6_outputs(7430) <= b and not a;
    layer6_outputs(7431) <= a or b;
    layer6_outputs(7432) <= '1';
    layer6_outputs(7433) <= not (a or b);
    layer6_outputs(7434) <= a;
    layer6_outputs(7435) <= not a;
    layer6_outputs(7436) <= not b or a;
    layer6_outputs(7437) <= b;
    layer6_outputs(7438) <= not (a and b);
    layer6_outputs(7439) <= not (a xor b);
    layer6_outputs(7440) <= not (a xor b);
    layer6_outputs(7441) <= not (a and b);
    layer6_outputs(7442) <= not b;
    layer6_outputs(7443) <= a;
    layer6_outputs(7444) <= a and b;
    layer6_outputs(7445) <= a;
    layer6_outputs(7446) <= not b;
    layer6_outputs(7447) <= a xor b;
    layer6_outputs(7448) <= not a;
    layer6_outputs(7449) <= a or b;
    layer6_outputs(7450) <= not a;
    layer6_outputs(7451) <= not b;
    layer6_outputs(7452) <= not b;
    layer6_outputs(7453) <= a and not b;
    layer6_outputs(7454) <= '0';
    layer6_outputs(7455) <= not b;
    layer6_outputs(7456) <= not a;
    layer6_outputs(7457) <= not b or a;
    layer6_outputs(7458) <= '1';
    layer6_outputs(7459) <= a;
    layer6_outputs(7460) <= a xor b;
    layer6_outputs(7461) <= not b or a;
    layer6_outputs(7462) <= not b or a;
    layer6_outputs(7463) <= not (a or b);
    layer6_outputs(7464) <= not b or a;
    layer6_outputs(7465) <= a;
    layer6_outputs(7466) <= not a;
    layer6_outputs(7467) <= a;
    layer6_outputs(7468) <= not b;
    layer6_outputs(7469) <= not a or b;
    layer6_outputs(7470) <= b;
    layer6_outputs(7471) <= not (a xor b);
    layer6_outputs(7472) <= not a or b;
    layer6_outputs(7473) <= not b;
    layer6_outputs(7474) <= b;
    layer6_outputs(7475) <= a xor b;
    layer6_outputs(7476) <= not a;
    layer6_outputs(7477) <= b;
    layer6_outputs(7478) <= a and not b;
    layer6_outputs(7479) <= a;
    layer6_outputs(7480) <= not (a xor b);
    layer6_outputs(7481) <= not (a or b);
    layer6_outputs(7482) <= b;
    layer6_outputs(7483) <= not (a xor b);
    layer6_outputs(7484) <= not a;
    layer6_outputs(7485) <= not (a xor b);
    layer6_outputs(7486) <= a and b;
    layer6_outputs(7487) <= not a or b;
    layer6_outputs(7488) <= b;
    layer6_outputs(7489) <= not (a xor b);
    layer6_outputs(7490) <= a;
    layer6_outputs(7491) <= b and not a;
    layer6_outputs(7492) <= a xor b;
    layer6_outputs(7493) <= a xor b;
    layer6_outputs(7494) <= not (a xor b);
    layer6_outputs(7495) <= a xor b;
    layer6_outputs(7496) <= not a;
    layer6_outputs(7497) <= not b;
    layer6_outputs(7498) <= b;
    layer6_outputs(7499) <= not a;
    layer6_outputs(7500) <= not (a and b);
    layer6_outputs(7501) <= a xor b;
    layer6_outputs(7502) <= not b;
    layer6_outputs(7503) <= not b;
    layer6_outputs(7504) <= b;
    layer6_outputs(7505) <= not a;
    layer6_outputs(7506) <= '1';
    layer6_outputs(7507) <= b;
    layer6_outputs(7508) <= not (a and b);
    layer6_outputs(7509) <= not (a and b);
    layer6_outputs(7510) <= a or b;
    layer6_outputs(7511) <= b;
    layer6_outputs(7512) <= b;
    layer6_outputs(7513) <= not a;
    layer6_outputs(7514) <= a xor b;
    layer6_outputs(7515) <= not (a xor b);
    layer6_outputs(7516) <= not (a and b);
    layer6_outputs(7517) <= not (a xor b);
    layer6_outputs(7518) <= not b;
    layer6_outputs(7519) <= a or b;
    layer6_outputs(7520) <= not b;
    layer6_outputs(7521) <= a;
    layer6_outputs(7522) <= a or b;
    layer6_outputs(7523) <= not (a xor b);
    layer6_outputs(7524) <= not b;
    layer6_outputs(7525) <= not b;
    layer6_outputs(7526) <= a;
    layer6_outputs(7527) <= a and b;
    layer6_outputs(7528) <= not a or b;
    layer6_outputs(7529) <= not b or a;
    layer6_outputs(7530) <= not b or a;
    layer6_outputs(7531) <= not a;
    layer6_outputs(7532) <= not (a xor b);
    layer6_outputs(7533) <= not (a or b);
    layer6_outputs(7534) <= not (a xor b);
    layer6_outputs(7535) <= not (a xor b);
    layer6_outputs(7536) <= a;
    layer6_outputs(7537) <= b;
    layer6_outputs(7538) <= not b;
    layer6_outputs(7539) <= a;
    layer6_outputs(7540) <= not (a xor b);
    layer6_outputs(7541) <= not a;
    layer6_outputs(7542) <= not b;
    layer6_outputs(7543) <= a xor b;
    layer6_outputs(7544) <= not b;
    layer6_outputs(7545) <= not (a xor b);
    layer6_outputs(7546) <= not a;
    layer6_outputs(7547) <= not b or a;
    layer6_outputs(7548) <= b and not a;
    layer6_outputs(7549) <= a and b;
    layer6_outputs(7550) <= a or b;
    layer6_outputs(7551) <= a xor b;
    layer6_outputs(7552) <= not (a xor b);
    layer6_outputs(7553) <= a;
    layer6_outputs(7554) <= not (a and b);
    layer6_outputs(7555) <= not (a or b);
    layer6_outputs(7556) <= not (a xor b);
    layer6_outputs(7557) <= not b;
    layer6_outputs(7558) <= a xor b;
    layer6_outputs(7559) <= a xor b;
    layer6_outputs(7560) <= a and not b;
    layer6_outputs(7561) <= a;
    layer6_outputs(7562) <= not a;
    layer6_outputs(7563) <= '0';
    layer6_outputs(7564) <= a and not b;
    layer6_outputs(7565) <= a xor b;
    layer6_outputs(7566) <= a;
    layer6_outputs(7567) <= not b or a;
    layer6_outputs(7568) <= a xor b;
    layer6_outputs(7569) <= not (a xor b);
    layer6_outputs(7570) <= not (a and b);
    layer6_outputs(7571) <= not (a xor b);
    layer6_outputs(7572) <= a and b;
    layer6_outputs(7573) <= a or b;
    layer6_outputs(7574) <= not a;
    layer6_outputs(7575) <= not b;
    layer6_outputs(7576) <= not (a and b);
    layer6_outputs(7577) <= b;
    layer6_outputs(7578) <= b;
    layer6_outputs(7579) <= a xor b;
    layer6_outputs(7580) <= not a or b;
    layer6_outputs(7581) <= a xor b;
    layer6_outputs(7582) <= a or b;
    layer6_outputs(7583) <= b;
    layer6_outputs(7584) <= not b;
    layer6_outputs(7585) <= not (a xor b);
    layer6_outputs(7586) <= a xor b;
    layer6_outputs(7587) <= not (a xor b);
    layer6_outputs(7588) <= b;
    layer6_outputs(7589) <= not (a xor b);
    layer6_outputs(7590) <= not (a xor b);
    layer6_outputs(7591) <= not (a xor b);
    layer6_outputs(7592) <= not (a xor b);
    layer6_outputs(7593) <= b and not a;
    layer6_outputs(7594) <= not a;
    layer6_outputs(7595) <= b and not a;
    layer6_outputs(7596) <= not (a xor b);
    layer6_outputs(7597) <= a or b;
    layer6_outputs(7598) <= a;
    layer6_outputs(7599) <= not a;
    layer6_outputs(7600) <= not a;
    layer6_outputs(7601) <= b;
    layer6_outputs(7602) <= not b;
    layer6_outputs(7603) <= a;
    layer6_outputs(7604) <= not b;
    layer6_outputs(7605) <= a;
    layer6_outputs(7606) <= not b;
    layer6_outputs(7607) <= not (a xor b);
    layer6_outputs(7608) <= not (a or b);
    layer6_outputs(7609) <= not a;
    layer6_outputs(7610) <= a or b;
    layer6_outputs(7611) <= b;
    layer6_outputs(7612) <= not b;
    layer6_outputs(7613) <= not b;
    layer6_outputs(7614) <= not (a xor b);
    layer6_outputs(7615) <= a;
    layer6_outputs(7616) <= not b;
    layer6_outputs(7617) <= not a;
    layer6_outputs(7618) <= not b;
    layer6_outputs(7619) <= not a;
    layer6_outputs(7620) <= a;
    layer6_outputs(7621) <= not (a and b);
    layer6_outputs(7622) <= b;
    layer6_outputs(7623) <= not (a xor b);
    layer6_outputs(7624) <= not a;
    layer6_outputs(7625) <= not (a xor b);
    layer6_outputs(7626) <= b;
    layer6_outputs(7627) <= a and not b;
    layer6_outputs(7628) <= a and b;
    layer6_outputs(7629) <= not b or a;
    layer6_outputs(7630) <= a and b;
    layer6_outputs(7631) <= a and b;
    layer6_outputs(7632) <= a;
    layer6_outputs(7633) <= a and b;
    layer6_outputs(7634) <= not a;
    layer6_outputs(7635) <= not b or a;
    layer6_outputs(7636) <= b and not a;
    layer6_outputs(7637) <= not (a xor b);
    layer6_outputs(7638) <= not (a and b);
    layer6_outputs(7639) <= b;
    layer6_outputs(7640) <= a and not b;
    layer6_outputs(7641) <= a xor b;
    layer6_outputs(7642) <= not (a xor b);
    layer6_outputs(7643) <= not (a xor b);
    layer6_outputs(7644) <= b and not a;
    layer6_outputs(7645) <= not a;
    layer6_outputs(7646) <= a and b;
    layer6_outputs(7647) <= a;
    layer6_outputs(7648) <= not (a and b);
    layer6_outputs(7649) <= not a or b;
    layer6_outputs(7650) <= not b;
    layer6_outputs(7651) <= not (a xor b);
    layer6_outputs(7652) <= b;
    layer6_outputs(7653) <= not (a xor b);
    layer6_outputs(7654) <= b and not a;
    layer6_outputs(7655) <= not b;
    layer6_outputs(7656) <= not a or b;
    layer6_outputs(7657) <= not b;
    layer6_outputs(7658) <= b;
    layer6_outputs(7659) <= not (a and b);
    layer6_outputs(7660) <= '1';
    layer6_outputs(7661) <= not (a xor b);
    layer6_outputs(7662) <= a xor b;
    layer6_outputs(7663) <= b;
    layer6_outputs(7664) <= a or b;
    layer6_outputs(7665) <= a;
    layer6_outputs(7666) <= not (a xor b);
    layer6_outputs(7667) <= a and not b;
    layer6_outputs(7668) <= b;
    layer6_outputs(7669) <= not (a and b);
    layer6_outputs(7670) <= not a;
    layer6_outputs(7671) <= not (a and b);
    layer6_outputs(7672) <= a xor b;
    layer6_outputs(7673) <= b;
    layer6_outputs(7674) <= not a or b;
    layer6_outputs(7675) <= b and not a;
    layer6_outputs(7676) <= not a;
    layer6_outputs(7677) <= a xor b;
    layer6_outputs(7678) <= not (a xor b);
    layer6_outputs(7679) <= b;
    layer6_outputs(7680) <= not b;
    layer6_outputs(7681) <= b and not a;
    layer6_outputs(7682) <= a xor b;
    layer6_outputs(7683) <= not a;
    layer6_outputs(7684) <= a or b;
    layer6_outputs(7685) <= b and not a;
    layer6_outputs(7686) <= a xor b;
    layer6_outputs(7687) <= not a;
    layer6_outputs(7688) <= '1';
    layer6_outputs(7689) <= a;
    layer6_outputs(7690) <= not (a or b);
    layer6_outputs(7691) <= not (a xor b);
    layer6_outputs(7692) <= a xor b;
    layer6_outputs(7693) <= not b or a;
    layer6_outputs(7694) <= not a;
    layer6_outputs(7695) <= not b;
    layer6_outputs(7696) <= not (a xor b);
    layer6_outputs(7697) <= a and not b;
    layer6_outputs(7698) <= b and not a;
    layer6_outputs(7699) <= a xor b;
    layer6_outputs(7700) <= b and not a;
    layer6_outputs(7701) <= b;
    layer6_outputs(7702) <= a xor b;
    layer6_outputs(7703) <= not (a or b);
    layer6_outputs(7704) <= a;
    layer6_outputs(7705) <= b;
    layer6_outputs(7706) <= b and not a;
    layer6_outputs(7707) <= not b or a;
    layer6_outputs(7708) <= a xor b;
    layer6_outputs(7709) <= a;
    layer6_outputs(7710) <= not (a or b);
    layer6_outputs(7711) <= not b;
    layer6_outputs(7712) <= not (a and b);
    layer6_outputs(7713) <= a and not b;
    layer6_outputs(7714) <= a xor b;
    layer6_outputs(7715) <= not b or a;
    layer6_outputs(7716) <= a xor b;
    layer6_outputs(7717) <= not b or a;
    layer6_outputs(7718) <= not a;
    layer6_outputs(7719) <= not a;
    layer6_outputs(7720) <= not a;
    layer6_outputs(7721) <= b;
    layer6_outputs(7722) <= a;
    layer6_outputs(7723) <= not a;
    layer6_outputs(7724) <= a and b;
    layer6_outputs(7725) <= not a;
    layer6_outputs(7726) <= a and b;
    layer6_outputs(7727) <= a;
    layer6_outputs(7728) <= not a;
    layer6_outputs(7729) <= a xor b;
    layer6_outputs(7730) <= a or b;
    layer6_outputs(7731) <= not (a and b);
    layer6_outputs(7732) <= a xor b;
    layer6_outputs(7733) <= b and not a;
    layer6_outputs(7734) <= b;
    layer6_outputs(7735) <= b and not a;
    layer6_outputs(7736) <= not a;
    layer6_outputs(7737) <= a xor b;
    layer6_outputs(7738) <= b;
    layer6_outputs(7739) <= not (a xor b);
    layer6_outputs(7740) <= not (a xor b);
    layer6_outputs(7741) <= a;
    layer6_outputs(7742) <= a;
    layer6_outputs(7743) <= not b or a;
    layer6_outputs(7744) <= not b;
    layer6_outputs(7745) <= a;
    layer6_outputs(7746) <= a xor b;
    layer6_outputs(7747) <= not b;
    layer6_outputs(7748) <= a xor b;
    layer6_outputs(7749) <= not b;
    layer6_outputs(7750) <= a xor b;
    layer6_outputs(7751) <= b;
    layer6_outputs(7752) <= not (a or b);
    layer6_outputs(7753) <= not b;
    layer6_outputs(7754) <= not (a or b);
    layer6_outputs(7755) <= not a or b;
    layer6_outputs(7756) <= b and not a;
    layer6_outputs(7757) <= not a or b;
    layer6_outputs(7758) <= b;
    layer6_outputs(7759) <= a;
    layer6_outputs(7760) <= not b;
    layer6_outputs(7761) <= not (a and b);
    layer6_outputs(7762) <= not b;
    layer6_outputs(7763) <= a or b;
    layer6_outputs(7764) <= not (a or b);
    layer6_outputs(7765) <= b;
    layer6_outputs(7766) <= not (a xor b);
    layer6_outputs(7767) <= b;
    layer6_outputs(7768) <= a;
    layer6_outputs(7769) <= not a;
    layer6_outputs(7770) <= not a;
    layer6_outputs(7771) <= not b;
    layer6_outputs(7772) <= b;
    layer6_outputs(7773) <= not b;
    layer6_outputs(7774) <= a and not b;
    layer6_outputs(7775) <= not a;
    layer6_outputs(7776) <= not a;
    layer6_outputs(7777) <= b;
    layer6_outputs(7778) <= a;
    layer6_outputs(7779) <= not a;
    layer6_outputs(7780) <= b and not a;
    layer6_outputs(7781) <= not a;
    layer6_outputs(7782) <= b and not a;
    layer6_outputs(7783) <= a;
    layer6_outputs(7784) <= b;
    layer6_outputs(7785) <= not (a and b);
    layer6_outputs(7786) <= not (a xor b);
    layer6_outputs(7787) <= b;
    layer6_outputs(7788) <= not (a xor b);
    layer6_outputs(7789) <= not a;
    layer6_outputs(7790) <= not (a xor b);
    layer6_outputs(7791) <= a xor b;
    layer6_outputs(7792) <= b;
    layer6_outputs(7793) <= not a;
    layer6_outputs(7794) <= a xor b;
    layer6_outputs(7795) <= not b or a;
    layer6_outputs(7796) <= not b;
    layer6_outputs(7797) <= a and b;
    layer6_outputs(7798) <= not a;
    layer6_outputs(7799) <= not a;
    layer6_outputs(7800) <= a;
    layer6_outputs(7801) <= not b;
    layer6_outputs(7802) <= not a;
    layer6_outputs(7803) <= a xor b;
    layer6_outputs(7804) <= not b or a;
    layer6_outputs(7805) <= not (a xor b);
    layer6_outputs(7806) <= not (a or b);
    layer6_outputs(7807) <= not b or a;
    layer6_outputs(7808) <= a and b;
    layer6_outputs(7809) <= not a;
    layer6_outputs(7810) <= a and not b;
    layer6_outputs(7811) <= b;
    layer6_outputs(7812) <= not (a xor b);
    layer6_outputs(7813) <= not (a or b);
    layer6_outputs(7814) <= b and not a;
    layer6_outputs(7815) <= b;
    layer6_outputs(7816) <= not b;
    layer6_outputs(7817) <= not b;
    layer6_outputs(7818) <= not b;
    layer6_outputs(7819) <= not b;
    layer6_outputs(7820) <= not (a xor b);
    layer6_outputs(7821) <= b;
    layer6_outputs(7822) <= b;
    layer6_outputs(7823) <= a;
    layer6_outputs(7824) <= a;
    layer6_outputs(7825) <= not a;
    layer6_outputs(7826) <= not b or a;
    layer6_outputs(7827) <= a xor b;
    layer6_outputs(7828) <= b;
    layer6_outputs(7829) <= not a;
    layer6_outputs(7830) <= not (a xor b);
    layer6_outputs(7831) <= a xor b;
    layer6_outputs(7832) <= a;
    layer6_outputs(7833) <= a xor b;
    layer6_outputs(7834) <= b;
    layer6_outputs(7835) <= not a;
    layer6_outputs(7836) <= not b;
    layer6_outputs(7837) <= not (a xor b);
    layer6_outputs(7838) <= not b;
    layer6_outputs(7839) <= a;
    layer6_outputs(7840) <= not a;
    layer6_outputs(7841) <= b;
    layer6_outputs(7842) <= not (a or b);
    layer6_outputs(7843) <= not b;
    layer6_outputs(7844) <= not b;
    layer6_outputs(7845) <= not b;
    layer6_outputs(7846) <= a or b;
    layer6_outputs(7847) <= not a;
    layer6_outputs(7848) <= not b;
    layer6_outputs(7849) <= a xor b;
    layer6_outputs(7850) <= not (a xor b);
    layer6_outputs(7851) <= b;
    layer6_outputs(7852) <= a;
    layer6_outputs(7853) <= a;
    layer6_outputs(7854) <= not (a xor b);
    layer6_outputs(7855) <= not (a xor b);
    layer6_outputs(7856) <= not (a xor b);
    layer6_outputs(7857) <= a;
    layer6_outputs(7858) <= not a or b;
    layer6_outputs(7859) <= not b;
    layer6_outputs(7860) <= not (a and b);
    layer6_outputs(7861) <= a and not b;
    layer6_outputs(7862) <= not a;
    layer6_outputs(7863) <= not a;
    layer6_outputs(7864) <= not (a xor b);
    layer6_outputs(7865) <= not b;
    layer6_outputs(7866) <= not b;
    layer6_outputs(7867) <= not (a xor b);
    layer6_outputs(7868) <= a xor b;
    layer6_outputs(7869) <= b;
    layer6_outputs(7870) <= not b or a;
    layer6_outputs(7871) <= a xor b;
    layer6_outputs(7872) <= not a;
    layer6_outputs(7873) <= a and b;
    layer6_outputs(7874) <= not a or b;
    layer6_outputs(7875) <= not a;
    layer6_outputs(7876) <= not b;
    layer6_outputs(7877) <= not (a xor b);
    layer6_outputs(7878) <= not a;
    layer6_outputs(7879) <= a and not b;
    layer6_outputs(7880) <= not (a xor b);
    layer6_outputs(7881) <= not a;
    layer6_outputs(7882) <= a xor b;
    layer6_outputs(7883) <= a or b;
    layer6_outputs(7884) <= a and not b;
    layer6_outputs(7885) <= b;
    layer6_outputs(7886) <= not b;
    layer6_outputs(7887) <= not a or b;
    layer6_outputs(7888) <= a xor b;
    layer6_outputs(7889) <= not (a and b);
    layer6_outputs(7890) <= a or b;
    layer6_outputs(7891) <= b and not a;
    layer6_outputs(7892) <= not (a and b);
    layer6_outputs(7893) <= a;
    layer6_outputs(7894) <= not (a xor b);
    layer6_outputs(7895) <= a xor b;
    layer6_outputs(7896) <= not (a or b);
    layer6_outputs(7897) <= not (a or b);
    layer6_outputs(7898) <= a;
    layer6_outputs(7899) <= not b;
    layer6_outputs(7900) <= a;
    layer6_outputs(7901) <= a xor b;
    layer6_outputs(7902) <= not b or a;
    layer6_outputs(7903) <= not (a xor b);
    layer6_outputs(7904) <= b;
    layer6_outputs(7905) <= not a;
    layer6_outputs(7906) <= a xor b;
    layer6_outputs(7907) <= a;
    layer6_outputs(7908) <= not b;
    layer6_outputs(7909) <= b;
    layer6_outputs(7910) <= not a;
    layer6_outputs(7911) <= not b or a;
    layer6_outputs(7912) <= not b;
    layer6_outputs(7913) <= a;
    layer6_outputs(7914) <= a xor b;
    layer6_outputs(7915) <= a xor b;
    layer6_outputs(7916) <= b;
    layer6_outputs(7917) <= a xor b;
    layer6_outputs(7918) <= b;
    layer6_outputs(7919) <= a xor b;
    layer6_outputs(7920) <= not a or b;
    layer6_outputs(7921) <= not b;
    layer6_outputs(7922) <= not a or b;
    layer6_outputs(7923) <= not a;
    layer6_outputs(7924) <= b;
    layer6_outputs(7925) <= a or b;
    layer6_outputs(7926) <= a;
    layer6_outputs(7927) <= a xor b;
    layer6_outputs(7928) <= a xor b;
    layer6_outputs(7929) <= b;
    layer6_outputs(7930) <= b;
    layer6_outputs(7931) <= not b or a;
    layer6_outputs(7932) <= not b;
    layer6_outputs(7933) <= not (a xor b);
    layer6_outputs(7934) <= not a;
    layer6_outputs(7935) <= a xor b;
    layer6_outputs(7936) <= not (a xor b);
    layer6_outputs(7937) <= not (a and b);
    layer6_outputs(7938) <= b and not a;
    layer6_outputs(7939) <= b;
    layer6_outputs(7940) <= not (a and b);
    layer6_outputs(7941) <= b;
    layer6_outputs(7942) <= not a or b;
    layer6_outputs(7943) <= not b;
    layer6_outputs(7944) <= a or b;
    layer6_outputs(7945) <= not (a xor b);
    layer6_outputs(7946) <= not b or a;
    layer6_outputs(7947) <= not (a xor b);
    layer6_outputs(7948) <= not a;
    layer6_outputs(7949) <= b and not a;
    layer6_outputs(7950) <= a and not b;
    layer6_outputs(7951) <= b;
    layer6_outputs(7952) <= not b;
    layer6_outputs(7953) <= a;
    layer6_outputs(7954) <= not a or b;
    layer6_outputs(7955) <= a;
    layer6_outputs(7956) <= a or b;
    layer6_outputs(7957) <= b and not a;
    layer6_outputs(7958) <= '1';
    layer6_outputs(7959) <= not (a and b);
    layer6_outputs(7960) <= not a or b;
    layer6_outputs(7961) <= not b;
    layer6_outputs(7962) <= a or b;
    layer6_outputs(7963) <= b;
    layer6_outputs(7964) <= a and b;
    layer6_outputs(7965) <= not b or a;
    layer6_outputs(7966) <= a;
    layer6_outputs(7967) <= a or b;
    layer6_outputs(7968) <= a;
    layer6_outputs(7969) <= a;
    layer6_outputs(7970) <= b;
    layer6_outputs(7971) <= a xor b;
    layer6_outputs(7972) <= a;
    layer6_outputs(7973) <= not b;
    layer6_outputs(7974) <= not a;
    layer6_outputs(7975) <= a xor b;
    layer6_outputs(7976) <= not a or b;
    layer6_outputs(7977) <= a;
    layer6_outputs(7978) <= not (a xor b);
    layer6_outputs(7979) <= not b;
    layer6_outputs(7980) <= a or b;
    layer6_outputs(7981) <= not (a xor b);
    layer6_outputs(7982) <= not (a xor b);
    layer6_outputs(7983) <= not a;
    layer6_outputs(7984) <= b;
    layer6_outputs(7985) <= not a;
    layer6_outputs(7986) <= not a or b;
    layer6_outputs(7987) <= a xor b;
    layer6_outputs(7988) <= a and b;
    layer6_outputs(7989) <= not b or a;
    layer6_outputs(7990) <= a;
    layer6_outputs(7991) <= not (a or b);
    layer6_outputs(7992) <= not a;
    layer6_outputs(7993) <= not a or b;
    layer6_outputs(7994) <= b;
    layer6_outputs(7995) <= not (a xor b);
    layer6_outputs(7996) <= not b;
    layer6_outputs(7997) <= a;
    layer6_outputs(7998) <= a xor b;
    layer6_outputs(7999) <= not b or a;
    layer6_outputs(8000) <= not (a and b);
    layer6_outputs(8001) <= a xor b;
    layer6_outputs(8002) <= not a;
    layer6_outputs(8003) <= not (a xor b);
    layer6_outputs(8004) <= not a;
    layer6_outputs(8005) <= b;
    layer6_outputs(8006) <= not a;
    layer6_outputs(8007) <= not (a or b);
    layer6_outputs(8008) <= not b or a;
    layer6_outputs(8009) <= not (a xor b);
    layer6_outputs(8010) <= a xor b;
    layer6_outputs(8011) <= a xor b;
    layer6_outputs(8012) <= not (a xor b);
    layer6_outputs(8013) <= not b;
    layer6_outputs(8014) <= not (a xor b);
    layer6_outputs(8015) <= not (a xor b);
    layer6_outputs(8016) <= not (a xor b);
    layer6_outputs(8017) <= b;
    layer6_outputs(8018) <= a xor b;
    layer6_outputs(8019) <= not b or a;
    layer6_outputs(8020) <= a;
    layer6_outputs(8021) <= not (a xor b);
    layer6_outputs(8022) <= a or b;
    layer6_outputs(8023) <= not a or b;
    layer6_outputs(8024) <= b and not a;
    layer6_outputs(8025) <= a;
    layer6_outputs(8026) <= not (a xor b);
    layer6_outputs(8027) <= a or b;
    layer6_outputs(8028) <= not a;
    layer6_outputs(8029) <= not b;
    layer6_outputs(8030) <= not b;
    layer6_outputs(8031) <= a xor b;
    layer6_outputs(8032) <= a and b;
    layer6_outputs(8033) <= a and b;
    layer6_outputs(8034) <= not (a xor b);
    layer6_outputs(8035) <= a and b;
    layer6_outputs(8036) <= b;
    layer6_outputs(8037) <= not b or a;
    layer6_outputs(8038) <= a or b;
    layer6_outputs(8039) <= b;
    layer6_outputs(8040) <= b;
    layer6_outputs(8041) <= b;
    layer6_outputs(8042) <= a xor b;
    layer6_outputs(8043) <= not (a and b);
    layer6_outputs(8044) <= not (a xor b);
    layer6_outputs(8045) <= not b or a;
    layer6_outputs(8046) <= a and b;
    layer6_outputs(8047) <= not b;
    layer6_outputs(8048) <= not (a xor b);
    layer6_outputs(8049) <= not a or b;
    layer6_outputs(8050) <= a;
    layer6_outputs(8051) <= a and not b;
    layer6_outputs(8052) <= b and not a;
    layer6_outputs(8053) <= a;
    layer6_outputs(8054) <= not b;
    layer6_outputs(8055) <= b;
    layer6_outputs(8056) <= b and not a;
    layer6_outputs(8057) <= a and b;
    layer6_outputs(8058) <= a xor b;
    layer6_outputs(8059) <= not a;
    layer6_outputs(8060) <= a or b;
    layer6_outputs(8061) <= not b;
    layer6_outputs(8062) <= a xor b;
    layer6_outputs(8063) <= not b;
    layer6_outputs(8064) <= a and b;
    layer6_outputs(8065) <= b;
    layer6_outputs(8066) <= not (a xor b);
    layer6_outputs(8067) <= a;
    layer6_outputs(8068) <= a xor b;
    layer6_outputs(8069) <= not b or a;
    layer6_outputs(8070) <= not a;
    layer6_outputs(8071) <= not b;
    layer6_outputs(8072) <= a and not b;
    layer6_outputs(8073) <= not (a and b);
    layer6_outputs(8074) <= a or b;
    layer6_outputs(8075) <= a xor b;
    layer6_outputs(8076) <= b;
    layer6_outputs(8077) <= not b;
    layer6_outputs(8078) <= a;
    layer6_outputs(8079) <= a;
    layer6_outputs(8080) <= b;
    layer6_outputs(8081) <= not (a xor b);
    layer6_outputs(8082) <= a;
    layer6_outputs(8083) <= not (a xor b);
    layer6_outputs(8084) <= a;
    layer6_outputs(8085) <= a xor b;
    layer6_outputs(8086) <= not (a or b);
    layer6_outputs(8087) <= b;
    layer6_outputs(8088) <= b and not a;
    layer6_outputs(8089) <= a and not b;
    layer6_outputs(8090) <= not b;
    layer6_outputs(8091) <= not b or a;
    layer6_outputs(8092) <= not a;
    layer6_outputs(8093) <= not (a xor b);
    layer6_outputs(8094) <= not (a xor b);
    layer6_outputs(8095) <= not a;
    layer6_outputs(8096) <= b;
    layer6_outputs(8097) <= not (a or b);
    layer6_outputs(8098) <= a or b;
    layer6_outputs(8099) <= b;
    layer6_outputs(8100) <= b and not a;
    layer6_outputs(8101) <= not (a xor b);
    layer6_outputs(8102) <= not (a xor b);
    layer6_outputs(8103) <= a or b;
    layer6_outputs(8104) <= a;
    layer6_outputs(8105) <= not a;
    layer6_outputs(8106) <= a;
    layer6_outputs(8107) <= a xor b;
    layer6_outputs(8108) <= a and not b;
    layer6_outputs(8109) <= not b;
    layer6_outputs(8110) <= a xor b;
    layer6_outputs(8111) <= not a or b;
    layer6_outputs(8112) <= a xor b;
    layer6_outputs(8113) <= not (a and b);
    layer6_outputs(8114) <= a xor b;
    layer6_outputs(8115) <= not b or a;
    layer6_outputs(8116) <= a;
    layer6_outputs(8117) <= not b;
    layer6_outputs(8118) <= not a;
    layer6_outputs(8119) <= not (a xor b);
    layer6_outputs(8120) <= not b;
    layer6_outputs(8121) <= b;
    layer6_outputs(8122) <= a and not b;
    layer6_outputs(8123) <= a xor b;
    layer6_outputs(8124) <= a;
    layer6_outputs(8125) <= not a or b;
    layer6_outputs(8126) <= a and not b;
    layer6_outputs(8127) <= not (a xor b);
    layer6_outputs(8128) <= not (a xor b);
    layer6_outputs(8129) <= not (a xor b);
    layer6_outputs(8130) <= not (a and b);
    layer6_outputs(8131) <= a;
    layer6_outputs(8132) <= not b;
    layer6_outputs(8133) <= not b;
    layer6_outputs(8134) <= a xor b;
    layer6_outputs(8135) <= not a;
    layer6_outputs(8136) <= b;
    layer6_outputs(8137) <= not a;
    layer6_outputs(8138) <= a;
    layer6_outputs(8139) <= a xor b;
    layer6_outputs(8140) <= not a or b;
    layer6_outputs(8141) <= not (a xor b);
    layer6_outputs(8142) <= a xor b;
    layer6_outputs(8143) <= not b;
    layer6_outputs(8144) <= not (a xor b);
    layer6_outputs(8145) <= not a;
    layer6_outputs(8146) <= not b;
    layer6_outputs(8147) <= not a;
    layer6_outputs(8148) <= a or b;
    layer6_outputs(8149) <= a xor b;
    layer6_outputs(8150) <= not b;
    layer6_outputs(8151) <= a and not b;
    layer6_outputs(8152) <= a xor b;
    layer6_outputs(8153) <= not b;
    layer6_outputs(8154) <= not b;
    layer6_outputs(8155) <= a and not b;
    layer6_outputs(8156) <= not a;
    layer6_outputs(8157) <= not a;
    layer6_outputs(8158) <= b;
    layer6_outputs(8159) <= a;
    layer6_outputs(8160) <= not (a or b);
    layer6_outputs(8161) <= a xor b;
    layer6_outputs(8162) <= not (a xor b);
    layer6_outputs(8163) <= not a;
    layer6_outputs(8164) <= a and b;
    layer6_outputs(8165) <= a and not b;
    layer6_outputs(8166) <= a and not b;
    layer6_outputs(8167) <= a and b;
    layer6_outputs(8168) <= a xor b;
    layer6_outputs(8169) <= not a;
    layer6_outputs(8170) <= not a or b;
    layer6_outputs(8171) <= not b or a;
    layer6_outputs(8172) <= not (a xor b);
    layer6_outputs(8173) <= b;
    layer6_outputs(8174) <= not a;
    layer6_outputs(8175) <= a xor b;
    layer6_outputs(8176) <= not (a and b);
    layer6_outputs(8177) <= not a or b;
    layer6_outputs(8178) <= not a or b;
    layer6_outputs(8179) <= b;
    layer6_outputs(8180) <= a and b;
    layer6_outputs(8181) <= b and not a;
    layer6_outputs(8182) <= a;
    layer6_outputs(8183) <= b;
    layer6_outputs(8184) <= not b or a;
    layer6_outputs(8185) <= not (a and b);
    layer6_outputs(8186) <= a xor b;
    layer6_outputs(8187) <= a xor b;
    layer6_outputs(8188) <= a and b;
    layer6_outputs(8189) <= not (a and b);
    layer6_outputs(8190) <= a;
    layer6_outputs(8191) <= not b;
    layer6_outputs(8192) <= b;
    layer6_outputs(8193) <= a xor b;
    layer6_outputs(8194) <= not a;
    layer6_outputs(8195) <= not b;
    layer6_outputs(8196) <= b and not a;
    layer6_outputs(8197) <= not (a xor b);
    layer6_outputs(8198) <= not (a xor b);
    layer6_outputs(8199) <= a xor b;
    layer6_outputs(8200) <= a and not b;
    layer6_outputs(8201) <= a;
    layer6_outputs(8202) <= a and b;
    layer6_outputs(8203) <= b;
    layer6_outputs(8204) <= '1';
    layer6_outputs(8205) <= a and b;
    layer6_outputs(8206) <= not (a xor b);
    layer6_outputs(8207) <= b;
    layer6_outputs(8208) <= a xor b;
    layer6_outputs(8209) <= a;
    layer6_outputs(8210) <= b and not a;
    layer6_outputs(8211) <= b;
    layer6_outputs(8212) <= not b;
    layer6_outputs(8213) <= not (a or b);
    layer6_outputs(8214) <= not (a or b);
    layer6_outputs(8215) <= not b;
    layer6_outputs(8216) <= not (a and b);
    layer6_outputs(8217) <= a;
    layer6_outputs(8218) <= not a;
    layer6_outputs(8219) <= not b;
    layer6_outputs(8220) <= not a;
    layer6_outputs(8221) <= not a or b;
    layer6_outputs(8222) <= not a;
    layer6_outputs(8223) <= b;
    layer6_outputs(8224) <= a and b;
    layer6_outputs(8225) <= b and not a;
    layer6_outputs(8226) <= a xor b;
    layer6_outputs(8227) <= a;
    layer6_outputs(8228) <= not a;
    layer6_outputs(8229) <= not a;
    layer6_outputs(8230) <= a;
    layer6_outputs(8231) <= a xor b;
    layer6_outputs(8232) <= not (a or b);
    layer6_outputs(8233) <= a xor b;
    layer6_outputs(8234) <= not a;
    layer6_outputs(8235) <= not (a or b);
    layer6_outputs(8236) <= not b;
    layer6_outputs(8237) <= b;
    layer6_outputs(8238) <= a;
    layer6_outputs(8239) <= b;
    layer6_outputs(8240) <= b;
    layer6_outputs(8241) <= not b;
    layer6_outputs(8242) <= a or b;
    layer6_outputs(8243) <= a xor b;
    layer6_outputs(8244) <= not a;
    layer6_outputs(8245) <= a xor b;
    layer6_outputs(8246) <= b;
    layer6_outputs(8247) <= a and b;
    layer6_outputs(8248) <= a xor b;
    layer6_outputs(8249) <= not a;
    layer6_outputs(8250) <= a or b;
    layer6_outputs(8251) <= b;
    layer6_outputs(8252) <= a and not b;
    layer6_outputs(8253) <= not b or a;
    layer6_outputs(8254) <= b;
    layer6_outputs(8255) <= b and not a;
    layer6_outputs(8256) <= b and not a;
    layer6_outputs(8257) <= not (a or b);
    layer6_outputs(8258) <= not b or a;
    layer6_outputs(8259) <= not (a and b);
    layer6_outputs(8260) <= not b;
    layer6_outputs(8261) <= a;
    layer6_outputs(8262) <= a xor b;
    layer6_outputs(8263) <= '1';
    layer6_outputs(8264) <= not a;
    layer6_outputs(8265) <= b and not a;
    layer6_outputs(8266) <= not b;
    layer6_outputs(8267) <= a xor b;
    layer6_outputs(8268) <= a or b;
    layer6_outputs(8269) <= not b;
    layer6_outputs(8270) <= not (a xor b);
    layer6_outputs(8271) <= b;
    layer6_outputs(8272) <= a;
    layer6_outputs(8273) <= not a;
    layer6_outputs(8274) <= b;
    layer6_outputs(8275) <= not (a or b);
    layer6_outputs(8276) <= not (a xor b);
    layer6_outputs(8277) <= not (a and b);
    layer6_outputs(8278) <= not b;
    layer6_outputs(8279) <= not b;
    layer6_outputs(8280) <= b and not a;
    layer6_outputs(8281) <= not a;
    layer6_outputs(8282) <= b;
    layer6_outputs(8283) <= not a;
    layer6_outputs(8284) <= b;
    layer6_outputs(8285) <= a or b;
    layer6_outputs(8286) <= not (a xor b);
    layer6_outputs(8287) <= a and not b;
    layer6_outputs(8288) <= a xor b;
    layer6_outputs(8289) <= b;
    layer6_outputs(8290) <= not a;
    layer6_outputs(8291) <= not (a xor b);
    layer6_outputs(8292) <= a and not b;
    layer6_outputs(8293) <= b;
    layer6_outputs(8294) <= not b or a;
    layer6_outputs(8295) <= b;
    layer6_outputs(8296) <= '1';
    layer6_outputs(8297) <= not (a xor b);
    layer6_outputs(8298) <= not (a xor b);
    layer6_outputs(8299) <= b;
    layer6_outputs(8300) <= not b;
    layer6_outputs(8301) <= not (a or b);
    layer6_outputs(8302) <= not b or a;
    layer6_outputs(8303) <= not b or a;
    layer6_outputs(8304) <= a;
    layer6_outputs(8305) <= not b or a;
    layer6_outputs(8306) <= b;
    layer6_outputs(8307) <= not b;
    layer6_outputs(8308) <= not b;
    layer6_outputs(8309) <= not (a and b);
    layer6_outputs(8310) <= b and not a;
    layer6_outputs(8311) <= b and not a;
    layer6_outputs(8312) <= b and not a;
    layer6_outputs(8313) <= not (a xor b);
    layer6_outputs(8314) <= not a;
    layer6_outputs(8315) <= b;
    layer6_outputs(8316) <= a;
    layer6_outputs(8317) <= not a;
    layer6_outputs(8318) <= a;
    layer6_outputs(8319) <= b;
    layer6_outputs(8320) <= a and not b;
    layer6_outputs(8321) <= b and not a;
    layer6_outputs(8322) <= not (a and b);
    layer6_outputs(8323) <= not a;
    layer6_outputs(8324) <= not a;
    layer6_outputs(8325) <= not (a xor b);
    layer6_outputs(8326) <= b;
    layer6_outputs(8327) <= not a or b;
    layer6_outputs(8328) <= not a;
    layer6_outputs(8329) <= a or b;
    layer6_outputs(8330) <= a;
    layer6_outputs(8331) <= not (a xor b);
    layer6_outputs(8332) <= a;
    layer6_outputs(8333) <= not b;
    layer6_outputs(8334) <= not (a xor b);
    layer6_outputs(8335) <= not a or b;
    layer6_outputs(8336) <= a xor b;
    layer6_outputs(8337) <= not b;
    layer6_outputs(8338) <= a and b;
    layer6_outputs(8339) <= not b;
    layer6_outputs(8340) <= '1';
    layer6_outputs(8341) <= not b or a;
    layer6_outputs(8342) <= not b or a;
    layer6_outputs(8343) <= not (a and b);
    layer6_outputs(8344) <= not (a xor b);
    layer6_outputs(8345) <= a;
    layer6_outputs(8346) <= a and b;
    layer6_outputs(8347) <= not b or a;
    layer6_outputs(8348) <= a;
    layer6_outputs(8349) <= not a;
    layer6_outputs(8350) <= a and b;
    layer6_outputs(8351) <= a and b;
    layer6_outputs(8352) <= a;
    layer6_outputs(8353) <= not a or b;
    layer6_outputs(8354) <= not b or a;
    layer6_outputs(8355) <= not b;
    layer6_outputs(8356) <= a and not b;
    layer6_outputs(8357) <= not b or a;
    layer6_outputs(8358) <= not b;
    layer6_outputs(8359) <= '0';
    layer6_outputs(8360) <= a;
    layer6_outputs(8361) <= not (a xor b);
    layer6_outputs(8362) <= a or b;
    layer6_outputs(8363) <= not (a xor b);
    layer6_outputs(8364) <= a;
    layer6_outputs(8365) <= not a;
    layer6_outputs(8366) <= not a or b;
    layer6_outputs(8367) <= a;
    layer6_outputs(8368) <= not a;
    layer6_outputs(8369) <= '0';
    layer6_outputs(8370) <= b;
    layer6_outputs(8371) <= b;
    layer6_outputs(8372) <= not b or a;
    layer6_outputs(8373) <= not (a and b);
    layer6_outputs(8374) <= not (a xor b);
    layer6_outputs(8375) <= not (a and b);
    layer6_outputs(8376) <= b and not a;
    layer6_outputs(8377) <= a xor b;
    layer6_outputs(8378) <= b;
    layer6_outputs(8379) <= not (a xor b);
    layer6_outputs(8380) <= a and b;
    layer6_outputs(8381) <= not a or b;
    layer6_outputs(8382) <= a or b;
    layer6_outputs(8383) <= b;
    layer6_outputs(8384) <= b and not a;
    layer6_outputs(8385) <= b;
    layer6_outputs(8386) <= a;
    layer6_outputs(8387) <= not b or a;
    layer6_outputs(8388) <= not (a xor b);
    layer6_outputs(8389) <= '1';
    layer6_outputs(8390) <= not (a xor b);
    layer6_outputs(8391) <= not (a xor b);
    layer6_outputs(8392) <= not (a xor b);
    layer6_outputs(8393) <= not (a xor b);
    layer6_outputs(8394) <= a xor b;
    layer6_outputs(8395) <= a or b;
    layer6_outputs(8396) <= not b or a;
    layer6_outputs(8397) <= a and b;
    layer6_outputs(8398) <= b;
    layer6_outputs(8399) <= not b;
    layer6_outputs(8400) <= b;
    layer6_outputs(8401) <= b;
    layer6_outputs(8402) <= not (a xor b);
    layer6_outputs(8403) <= not b;
    layer6_outputs(8404) <= a xor b;
    layer6_outputs(8405) <= not (a xor b);
    layer6_outputs(8406) <= not (a xor b);
    layer6_outputs(8407) <= a xor b;
    layer6_outputs(8408) <= a and not b;
    layer6_outputs(8409) <= not b;
    layer6_outputs(8410) <= '0';
    layer6_outputs(8411) <= b;
    layer6_outputs(8412) <= not b or a;
    layer6_outputs(8413) <= b and not a;
    layer6_outputs(8414) <= b and not a;
    layer6_outputs(8415) <= not (a and b);
    layer6_outputs(8416) <= b;
    layer6_outputs(8417) <= b and not a;
    layer6_outputs(8418) <= not a;
    layer6_outputs(8419) <= not (a xor b);
    layer6_outputs(8420) <= not (a or b);
    layer6_outputs(8421) <= not (a or b);
    layer6_outputs(8422) <= a and b;
    layer6_outputs(8423) <= not b;
    layer6_outputs(8424) <= a;
    layer6_outputs(8425) <= a;
    layer6_outputs(8426) <= b;
    layer6_outputs(8427) <= b and not a;
    layer6_outputs(8428) <= a;
    layer6_outputs(8429) <= not a;
    layer6_outputs(8430) <= a xor b;
    layer6_outputs(8431) <= not b or a;
    layer6_outputs(8432) <= not (a xor b);
    layer6_outputs(8433) <= a and b;
    layer6_outputs(8434) <= not a;
    layer6_outputs(8435) <= '1';
    layer6_outputs(8436) <= a;
    layer6_outputs(8437) <= not (a xor b);
    layer6_outputs(8438) <= a and not b;
    layer6_outputs(8439) <= not b;
    layer6_outputs(8440) <= not (a or b);
    layer6_outputs(8441) <= not a;
    layer6_outputs(8442) <= not b;
    layer6_outputs(8443) <= not b;
    layer6_outputs(8444) <= not b or a;
    layer6_outputs(8445) <= not b;
    layer6_outputs(8446) <= not a;
    layer6_outputs(8447) <= not a;
    layer6_outputs(8448) <= a xor b;
    layer6_outputs(8449) <= not b;
    layer6_outputs(8450) <= not (a xor b);
    layer6_outputs(8451) <= a xor b;
    layer6_outputs(8452) <= not (a or b);
    layer6_outputs(8453) <= not (a or b);
    layer6_outputs(8454) <= b;
    layer6_outputs(8455) <= b;
    layer6_outputs(8456) <= not a;
    layer6_outputs(8457) <= b;
    layer6_outputs(8458) <= not b;
    layer6_outputs(8459) <= b and not a;
    layer6_outputs(8460) <= not (a xor b);
    layer6_outputs(8461) <= not a or b;
    layer6_outputs(8462) <= a;
    layer6_outputs(8463) <= a;
    layer6_outputs(8464) <= a;
    layer6_outputs(8465) <= not (a xor b);
    layer6_outputs(8466) <= b and not a;
    layer6_outputs(8467) <= a and b;
    layer6_outputs(8468) <= not b or a;
    layer6_outputs(8469) <= not a;
    layer6_outputs(8470) <= a xor b;
    layer6_outputs(8471) <= b;
    layer6_outputs(8472) <= not (a and b);
    layer6_outputs(8473) <= a;
    layer6_outputs(8474) <= not (a xor b);
    layer6_outputs(8475) <= not b;
    layer6_outputs(8476) <= not a;
    layer6_outputs(8477) <= b;
    layer6_outputs(8478) <= not a or b;
    layer6_outputs(8479) <= a;
    layer6_outputs(8480) <= a;
    layer6_outputs(8481) <= not a;
    layer6_outputs(8482) <= not a or b;
    layer6_outputs(8483) <= not b or a;
    layer6_outputs(8484) <= a;
    layer6_outputs(8485) <= not b;
    layer6_outputs(8486) <= not (a xor b);
    layer6_outputs(8487) <= a and b;
    layer6_outputs(8488) <= b;
    layer6_outputs(8489) <= a and b;
    layer6_outputs(8490) <= not b;
    layer6_outputs(8491) <= a;
    layer6_outputs(8492) <= a;
    layer6_outputs(8493) <= a;
    layer6_outputs(8494) <= not (a or b);
    layer6_outputs(8495) <= a;
    layer6_outputs(8496) <= a;
    layer6_outputs(8497) <= a and b;
    layer6_outputs(8498) <= a or b;
    layer6_outputs(8499) <= not (a xor b);
    layer6_outputs(8500) <= not b or a;
    layer6_outputs(8501) <= a;
    layer6_outputs(8502) <= not a;
    layer6_outputs(8503) <= a;
    layer6_outputs(8504) <= not b;
    layer6_outputs(8505) <= not a or b;
    layer6_outputs(8506) <= not b;
    layer6_outputs(8507) <= not a;
    layer6_outputs(8508) <= a xor b;
    layer6_outputs(8509) <= not (a xor b);
    layer6_outputs(8510) <= b;
    layer6_outputs(8511) <= b;
    layer6_outputs(8512) <= a;
    layer6_outputs(8513) <= not (a and b);
    layer6_outputs(8514) <= b and not a;
    layer6_outputs(8515) <= a;
    layer6_outputs(8516) <= a xor b;
    layer6_outputs(8517) <= not a;
    layer6_outputs(8518) <= not (a and b);
    layer6_outputs(8519) <= b;
    layer6_outputs(8520) <= not b;
    layer6_outputs(8521) <= a;
    layer6_outputs(8522) <= b and not a;
    layer6_outputs(8523) <= not a;
    layer6_outputs(8524) <= a and not b;
    layer6_outputs(8525) <= not b;
    layer6_outputs(8526) <= not (a xor b);
    layer6_outputs(8527) <= not a or b;
    layer6_outputs(8528) <= not b;
    layer6_outputs(8529) <= '1';
    layer6_outputs(8530) <= a;
    layer6_outputs(8531) <= b and not a;
    layer6_outputs(8532) <= a and b;
    layer6_outputs(8533) <= not a or b;
    layer6_outputs(8534) <= b;
    layer6_outputs(8535) <= not b;
    layer6_outputs(8536) <= a and not b;
    layer6_outputs(8537) <= not b or a;
    layer6_outputs(8538) <= not (a xor b);
    layer6_outputs(8539) <= not a;
    layer6_outputs(8540) <= a;
    layer6_outputs(8541) <= not (a and b);
    layer6_outputs(8542) <= a and not b;
    layer6_outputs(8543) <= not (a or b);
    layer6_outputs(8544) <= a or b;
    layer6_outputs(8545) <= b;
    layer6_outputs(8546) <= b;
    layer6_outputs(8547) <= a xor b;
    layer6_outputs(8548) <= not a;
    layer6_outputs(8549) <= b;
    layer6_outputs(8550) <= b;
    layer6_outputs(8551) <= b and not a;
    layer6_outputs(8552) <= a and not b;
    layer6_outputs(8553) <= not b;
    layer6_outputs(8554) <= b;
    layer6_outputs(8555) <= not (a and b);
    layer6_outputs(8556) <= not (a or b);
    layer6_outputs(8557) <= not b;
    layer6_outputs(8558) <= b;
    layer6_outputs(8559) <= b;
    layer6_outputs(8560) <= a xor b;
    layer6_outputs(8561) <= b;
    layer6_outputs(8562) <= b;
    layer6_outputs(8563) <= a;
    layer6_outputs(8564) <= a;
    layer6_outputs(8565) <= a;
    layer6_outputs(8566) <= not (a xor b);
    layer6_outputs(8567) <= b;
    layer6_outputs(8568) <= not a or b;
    layer6_outputs(8569) <= a and b;
    layer6_outputs(8570) <= not (a xor b);
    layer6_outputs(8571) <= not (a and b);
    layer6_outputs(8572) <= a and b;
    layer6_outputs(8573) <= not (a and b);
    layer6_outputs(8574) <= not a or b;
    layer6_outputs(8575) <= not a;
    layer6_outputs(8576) <= not a;
    layer6_outputs(8577) <= a or b;
    layer6_outputs(8578) <= b;
    layer6_outputs(8579) <= b;
    layer6_outputs(8580) <= a xor b;
    layer6_outputs(8581) <= not b;
    layer6_outputs(8582) <= not b;
    layer6_outputs(8583) <= not (a xor b);
    layer6_outputs(8584) <= b;
    layer6_outputs(8585) <= a xor b;
    layer6_outputs(8586) <= b;
    layer6_outputs(8587) <= b and not a;
    layer6_outputs(8588) <= not (a and b);
    layer6_outputs(8589) <= a xor b;
    layer6_outputs(8590) <= not a;
    layer6_outputs(8591) <= a xor b;
    layer6_outputs(8592) <= not a;
    layer6_outputs(8593) <= not (a xor b);
    layer6_outputs(8594) <= not a;
    layer6_outputs(8595) <= a and not b;
    layer6_outputs(8596) <= not (a xor b);
    layer6_outputs(8597) <= a xor b;
    layer6_outputs(8598) <= not b;
    layer6_outputs(8599) <= a and b;
    layer6_outputs(8600) <= a;
    layer6_outputs(8601) <= a and not b;
    layer6_outputs(8602) <= a;
    layer6_outputs(8603) <= a;
    layer6_outputs(8604) <= not a or b;
    layer6_outputs(8605) <= not a;
    layer6_outputs(8606) <= a and not b;
    layer6_outputs(8607) <= not (a or b);
    layer6_outputs(8608) <= b and not a;
    layer6_outputs(8609) <= a;
    layer6_outputs(8610) <= a;
    layer6_outputs(8611) <= b and not a;
    layer6_outputs(8612) <= a;
    layer6_outputs(8613) <= not a;
    layer6_outputs(8614) <= not a or b;
    layer6_outputs(8615) <= a;
    layer6_outputs(8616) <= not a;
    layer6_outputs(8617) <= b;
    layer6_outputs(8618) <= not b;
    layer6_outputs(8619) <= not a or b;
    layer6_outputs(8620) <= a xor b;
    layer6_outputs(8621) <= a and not b;
    layer6_outputs(8622) <= a xor b;
    layer6_outputs(8623) <= a xor b;
    layer6_outputs(8624) <= a;
    layer6_outputs(8625) <= not b;
    layer6_outputs(8626) <= not b;
    layer6_outputs(8627) <= not a or b;
    layer6_outputs(8628) <= not (a xor b);
    layer6_outputs(8629) <= a and b;
    layer6_outputs(8630) <= a;
    layer6_outputs(8631) <= b and not a;
    layer6_outputs(8632) <= not a or b;
    layer6_outputs(8633) <= '0';
    layer6_outputs(8634) <= not b or a;
    layer6_outputs(8635) <= b and not a;
    layer6_outputs(8636) <= not b or a;
    layer6_outputs(8637) <= a xor b;
    layer6_outputs(8638) <= a and b;
    layer6_outputs(8639) <= a xor b;
    layer6_outputs(8640) <= a and not b;
    layer6_outputs(8641) <= not (a xor b);
    layer6_outputs(8642) <= a xor b;
    layer6_outputs(8643) <= not b or a;
    layer6_outputs(8644) <= not (a or b);
    layer6_outputs(8645) <= b;
    layer6_outputs(8646) <= not a;
    layer6_outputs(8647) <= b;
    layer6_outputs(8648) <= a;
    layer6_outputs(8649) <= not b;
    layer6_outputs(8650) <= a xor b;
    layer6_outputs(8651) <= a;
    layer6_outputs(8652) <= not a;
    layer6_outputs(8653) <= not a or b;
    layer6_outputs(8654) <= a and b;
    layer6_outputs(8655) <= not a or b;
    layer6_outputs(8656) <= a and not b;
    layer6_outputs(8657) <= b;
    layer6_outputs(8658) <= b;
    layer6_outputs(8659) <= a;
    layer6_outputs(8660) <= not (a xor b);
    layer6_outputs(8661) <= a xor b;
    layer6_outputs(8662) <= a xor b;
    layer6_outputs(8663) <= not a;
    layer6_outputs(8664) <= not (a and b);
    layer6_outputs(8665) <= a xor b;
    layer6_outputs(8666) <= b;
    layer6_outputs(8667) <= not (a xor b);
    layer6_outputs(8668) <= b;
    layer6_outputs(8669) <= a xor b;
    layer6_outputs(8670) <= not a or b;
    layer6_outputs(8671) <= not b or a;
    layer6_outputs(8672) <= a xor b;
    layer6_outputs(8673) <= not a or b;
    layer6_outputs(8674) <= a;
    layer6_outputs(8675) <= not a;
    layer6_outputs(8676) <= a;
    layer6_outputs(8677) <= a or b;
    layer6_outputs(8678) <= not a or b;
    layer6_outputs(8679) <= not b;
    layer6_outputs(8680) <= a;
    layer6_outputs(8681) <= a;
    layer6_outputs(8682) <= not (a xor b);
    layer6_outputs(8683) <= not b;
    layer6_outputs(8684) <= not a or b;
    layer6_outputs(8685) <= b and not a;
    layer6_outputs(8686) <= not (a xor b);
    layer6_outputs(8687) <= not (a or b);
    layer6_outputs(8688) <= a;
    layer6_outputs(8689) <= not a;
    layer6_outputs(8690) <= a and not b;
    layer6_outputs(8691) <= not (a and b);
    layer6_outputs(8692) <= a;
    layer6_outputs(8693) <= not (a xor b);
    layer6_outputs(8694) <= b;
    layer6_outputs(8695) <= a;
    layer6_outputs(8696) <= a;
    layer6_outputs(8697) <= not (a or b);
    layer6_outputs(8698) <= b;
    layer6_outputs(8699) <= a;
    layer6_outputs(8700) <= b;
    layer6_outputs(8701) <= a;
    layer6_outputs(8702) <= not a;
    layer6_outputs(8703) <= a and not b;
    layer6_outputs(8704) <= a and b;
    layer6_outputs(8705) <= a and not b;
    layer6_outputs(8706) <= not a;
    layer6_outputs(8707) <= not (a xor b);
    layer6_outputs(8708) <= not b;
    layer6_outputs(8709) <= not a or b;
    layer6_outputs(8710) <= not a;
    layer6_outputs(8711) <= b;
    layer6_outputs(8712) <= a and b;
    layer6_outputs(8713) <= not a;
    layer6_outputs(8714) <= a;
    layer6_outputs(8715) <= not a;
    layer6_outputs(8716) <= not (a and b);
    layer6_outputs(8717) <= not (a or b);
    layer6_outputs(8718) <= a and not b;
    layer6_outputs(8719) <= a and b;
    layer6_outputs(8720) <= not b;
    layer6_outputs(8721) <= a or b;
    layer6_outputs(8722) <= a and b;
    layer6_outputs(8723) <= not (a or b);
    layer6_outputs(8724) <= a and b;
    layer6_outputs(8725) <= a xor b;
    layer6_outputs(8726) <= not b;
    layer6_outputs(8727) <= a and b;
    layer6_outputs(8728) <= a or b;
    layer6_outputs(8729) <= a;
    layer6_outputs(8730) <= a;
    layer6_outputs(8731) <= not (a or b);
    layer6_outputs(8732) <= not (a xor b);
    layer6_outputs(8733) <= not (a xor b);
    layer6_outputs(8734) <= not a;
    layer6_outputs(8735) <= not (a xor b);
    layer6_outputs(8736) <= a or b;
    layer6_outputs(8737) <= not b;
    layer6_outputs(8738) <= a;
    layer6_outputs(8739) <= not b;
    layer6_outputs(8740) <= not b;
    layer6_outputs(8741) <= a and b;
    layer6_outputs(8742) <= a;
    layer6_outputs(8743) <= b;
    layer6_outputs(8744) <= not b;
    layer6_outputs(8745) <= not a or b;
    layer6_outputs(8746) <= not b;
    layer6_outputs(8747) <= b and not a;
    layer6_outputs(8748) <= a xor b;
    layer6_outputs(8749) <= not b or a;
    layer6_outputs(8750) <= a;
    layer6_outputs(8751) <= not a or b;
    layer6_outputs(8752) <= not b;
    layer6_outputs(8753) <= b;
    layer6_outputs(8754) <= not a;
    layer6_outputs(8755) <= b;
    layer6_outputs(8756) <= not (a or b);
    layer6_outputs(8757) <= not (a xor b);
    layer6_outputs(8758) <= a and b;
    layer6_outputs(8759) <= a or b;
    layer6_outputs(8760) <= b;
    layer6_outputs(8761) <= a xor b;
    layer6_outputs(8762) <= a xor b;
    layer6_outputs(8763) <= a and not b;
    layer6_outputs(8764) <= not (a and b);
    layer6_outputs(8765) <= not (a xor b);
    layer6_outputs(8766) <= not b;
    layer6_outputs(8767) <= b;
    layer6_outputs(8768) <= a xor b;
    layer6_outputs(8769) <= a and not b;
    layer6_outputs(8770) <= not (a or b);
    layer6_outputs(8771) <= '0';
    layer6_outputs(8772) <= not b or a;
    layer6_outputs(8773) <= a or b;
    layer6_outputs(8774) <= not (a or b);
    layer6_outputs(8775) <= b;
    layer6_outputs(8776) <= not a;
    layer6_outputs(8777) <= not a;
    layer6_outputs(8778) <= not (a xor b);
    layer6_outputs(8779) <= not b;
    layer6_outputs(8780) <= a;
    layer6_outputs(8781) <= not a;
    layer6_outputs(8782) <= b;
    layer6_outputs(8783) <= a;
    layer6_outputs(8784) <= a and not b;
    layer6_outputs(8785) <= not b;
    layer6_outputs(8786) <= a and b;
    layer6_outputs(8787) <= not (a and b);
    layer6_outputs(8788) <= b and not a;
    layer6_outputs(8789) <= not a;
    layer6_outputs(8790) <= not b;
    layer6_outputs(8791) <= not (a xor b);
    layer6_outputs(8792) <= a xor b;
    layer6_outputs(8793) <= not b or a;
    layer6_outputs(8794) <= not (a and b);
    layer6_outputs(8795) <= not a;
    layer6_outputs(8796) <= not a;
    layer6_outputs(8797) <= a or b;
    layer6_outputs(8798) <= a;
    layer6_outputs(8799) <= not a;
    layer6_outputs(8800) <= not (a xor b);
    layer6_outputs(8801) <= not b or a;
    layer6_outputs(8802) <= not (a or b);
    layer6_outputs(8803) <= a and not b;
    layer6_outputs(8804) <= not (a xor b);
    layer6_outputs(8805) <= a and not b;
    layer6_outputs(8806) <= not a or b;
    layer6_outputs(8807) <= a or b;
    layer6_outputs(8808) <= not b;
    layer6_outputs(8809) <= a xor b;
    layer6_outputs(8810) <= not b;
    layer6_outputs(8811) <= not a or b;
    layer6_outputs(8812) <= a;
    layer6_outputs(8813) <= not a;
    layer6_outputs(8814) <= a or b;
    layer6_outputs(8815) <= not (a xor b);
    layer6_outputs(8816) <= not (a xor b);
    layer6_outputs(8817) <= a;
    layer6_outputs(8818) <= a xor b;
    layer6_outputs(8819) <= a xor b;
    layer6_outputs(8820) <= a xor b;
    layer6_outputs(8821) <= not (a or b);
    layer6_outputs(8822) <= not a;
    layer6_outputs(8823) <= b;
    layer6_outputs(8824) <= b;
    layer6_outputs(8825) <= a;
    layer6_outputs(8826) <= not a;
    layer6_outputs(8827) <= a;
    layer6_outputs(8828) <= a or b;
    layer6_outputs(8829) <= b and not a;
    layer6_outputs(8830) <= a xor b;
    layer6_outputs(8831) <= a;
    layer6_outputs(8832) <= not b or a;
    layer6_outputs(8833) <= not (a and b);
    layer6_outputs(8834) <= a;
    layer6_outputs(8835) <= not (a and b);
    layer6_outputs(8836) <= not a;
    layer6_outputs(8837) <= not b;
    layer6_outputs(8838) <= b;
    layer6_outputs(8839) <= not a;
    layer6_outputs(8840) <= b;
    layer6_outputs(8841) <= a;
    layer6_outputs(8842) <= a xor b;
    layer6_outputs(8843) <= b;
    layer6_outputs(8844) <= a;
    layer6_outputs(8845) <= a xor b;
    layer6_outputs(8846) <= not a;
    layer6_outputs(8847) <= not (a xor b);
    layer6_outputs(8848) <= b;
    layer6_outputs(8849) <= b;
    layer6_outputs(8850) <= a;
    layer6_outputs(8851) <= b;
    layer6_outputs(8852) <= a and b;
    layer6_outputs(8853) <= not b;
    layer6_outputs(8854) <= not a;
    layer6_outputs(8855) <= a and not b;
    layer6_outputs(8856) <= a;
    layer6_outputs(8857) <= a xor b;
    layer6_outputs(8858) <= a or b;
    layer6_outputs(8859) <= not b or a;
    layer6_outputs(8860) <= a;
    layer6_outputs(8861) <= b;
    layer6_outputs(8862) <= a;
    layer6_outputs(8863) <= a or b;
    layer6_outputs(8864) <= b;
    layer6_outputs(8865) <= not b or a;
    layer6_outputs(8866) <= b and not a;
    layer6_outputs(8867) <= b;
    layer6_outputs(8868) <= not b;
    layer6_outputs(8869) <= a or b;
    layer6_outputs(8870) <= a;
    layer6_outputs(8871) <= b;
    layer6_outputs(8872) <= not (a xor b);
    layer6_outputs(8873) <= a xor b;
    layer6_outputs(8874) <= not (a xor b);
    layer6_outputs(8875) <= b;
    layer6_outputs(8876) <= not (a xor b);
    layer6_outputs(8877) <= not (a xor b);
    layer6_outputs(8878) <= not a;
    layer6_outputs(8879) <= b and not a;
    layer6_outputs(8880) <= not b;
    layer6_outputs(8881) <= not (a and b);
    layer6_outputs(8882) <= b;
    layer6_outputs(8883) <= not b;
    layer6_outputs(8884) <= not a or b;
    layer6_outputs(8885) <= a and not b;
    layer6_outputs(8886) <= not (a xor b);
    layer6_outputs(8887) <= b;
    layer6_outputs(8888) <= a or b;
    layer6_outputs(8889) <= not (a and b);
    layer6_outputs(8890) <= not b or a;
    layer6_outputs(8891) <= a;
    layer6_outputs(8892) <= a xor b;
    layer6_outputs(8893) <= a and not b;
    layer6_outputs(8894) <= b;
    layer6_outputs(8895) <= a xor b;
    layer6_outputs(8896) <= a xor b;
    layer6_outputs(8897) <= not a;
    layer6_outputs(8898) <= not (a or b);
    layer6_outputs(8899) <= not a or b;
    layer6_outputs(8900) <= not (a xor b);
    layer6_outputs(8901) <= not b or a;
    layer6_outputs(8902) <= not (a xor b);
    layer6_outputs(8903) <= b;
    layer6_outputs(8904) <= a;
    layer6_outputs(8905) <= a;
    layer6_outputs(8906) <= a and not b;
    layer6_outputs(8907) <= not (a and b);
    layer6_outputs(8908) <= not b;
    layer6_outputs(8909) <= a;
    layer6_outputs(8910) <= not b;
    layer6_outputs(8911) <= not (a xor b);
    layer6_outputs(8912) <= a xor b;
    layer6_outputs(8913) <= b and not a;
    layer6_outputs(8914) <= not a;
    layer6_outputs(8915) <= not b;
    layer6_outputs(8916) <= a or b;
    layer6_outputs(8917) <= b and not a;
    layer6_outputs(8918) <= not b;
    layer6_outputs(8919) <= a;
    layer6_outputs(8920) <= not a;
    layer6_outputs(8921) <= a;
    layer6_outputs(8922) <= not (a xor b);
    layer6_outputs(8923) <= a and b;
    layer6_outputs(8924) <= not (a and b);
    layer6_outputs(8925) <= a;
    layer6_outputs(8926) <= a and b;
    layer6_outputs(8927) <= not b;
    layer6_outputs(8928) <= a or b;
    layer6_outputs(8929) <= not (a xor b);
    layer6_outputs(8930) <= a xor b;
    layer6_outputs(8931) <= a xor b;
    layer6_outputs(8932) <= b;
    layer6_outputs(8933) <= a and b;
    layer6_outputs(8934) <= a xor b;
    layer6_outputs(8935) <= not a;
    layer6_outputs(8936) <= not a;
    layer6_outputs(8937) <= not (a xor b);
    layer6_outputs(8938) <= not (a xor b);
    layer6_outputs(8939) <= b;
    layer6_outputs(8940) <= a or b;
    layer6_outputs(8941) <= b and not a;
    layer6_outputs(8942) <= not a or b;
    layer6_outputs(8943) <= not a;
    layer6_outputs(8944) <= b;
    layer6_outputs(8945) <= not (a and b);
    layer6_outputs(8946) <= not a;
    layer6_outputs(8947) <= b;
    layer6_outputs(8948) <= not b;
    layer6_outputs(8949) <= a xor b;
    layer6_outputs(8950) <= a;
    layer6_outputs(8951) <= a;
    layer6_outputs(8952) <= b;
    layer6_outputs(8953) <= not b or a;
    layer6_outputs(8954) <= a and b;
    layer6_outputs(8955) <= not (a or b);
    layer6_outputs(8956) <= not (a or b);
    layer6_outputs(8957) <= not b;
    layer6_outputs(8958) <= not (a xor b);
    layer6_outputs(8959) <= not (a xor b);
    layer6_outputs(8960) <= not b;
    layer6_outputs(8961) <= a and not b;
    layer6_outputs(8962) <= not (a xor b);
    layer6_outputs(8963) <= not (a xor b);
    layer6_outputs(8964) <= not (a xor b);
    layer6_outputs(8965) <= b;
    layer6_outputs(8966) <= not (a xor b);
    layer6_outputs(8967) <= a and b;
    layer6_outputs(8968) <= not (a xor b);
    layer6_outputs(8969) <= not (a xor b);
    layer6_outputs(8970) <= a and b;
    layer6_outputs(8971) <= not b;
    layer6_outputs(8972) <= a and not b;
    layer6_outputs(8973) <= not b or a;
    layer6_outputs(8974) <= not b;
    layer6_outputs(8975) <= a xor b;
    layer6_outputs(8976) <= not a;
    layer6_outputs(8977) <= a xor b;
    layer6_outputs(8978) <= not b;
    layer6_outputs(8979) <= a and b;
    layer6_outputs(8980) <= not (a xor b);
    layer6_outputs(8981) <= a and b;
    layer6_outputs(8982) <= a;
    layer6_outputs(8983) <= b;
    layer6_outputs(8984) <= not (a and b);
    layer6_outputs(8985) <= a or b;
    layer6_outputs(8986) <= b;
    layer6_outputs(8987) <= b and not a;
    layer6_outputs(8988) <= b and not a;
    layer6_outputs(8989) <= a;
    layer6_outputs(8990) <= not (a xor b);
    layer6_outputs(8991) <= a and b;
    layer6_outputs(8992) <= b;
    layer6_outputs(8993) <= not a;
    layer6_outputs(8994) <= a;
    layer6_outputs(8995) <= not b;
    layer6_outputs(8996) <= b;
    layer6_outputs(8997) <= a;
    layer6_outputs(8998) <= b;
    layer6_outputs(8999) <= not (a xor b);
    layer6_outputs(9000) <= not (a xor b);
    layer6_outputs(9001) <= not a;
    layer6_outputs(9002) <= b and not a;
    layer6_outputs(9003) <= a xor b;
    layer6_outputs(9004) <= b;
    layer6_outputs(9005) <= not a;
    layer6_outputs(9006) <= not (a xor b);
    layer6_outputs(9007) <= not (a and b);
    layer6_outputs(9008) <= a xor b;
    layer6_outputs(9009) <= a xor b;
    layer6_outputs(9010) <= a and not b;
    layer6_outputs(9011) <= a or b;
    layer6_outputs(9012) <= a xor b;
    layer6_outputs(9013) <= a xor b;
    layer6_outputs(9014) <= not (a xor b);
    layer6_outputs(9015) <= not (a or b);
    layer6_outputs(9016) <= not a;
    layer6_outputs(9017) <= a;
    layer6_outputs(9018) <= not (a and b);
    layer6_outputs(9019) <= not (a or b);
    layer6_outputs(9020) <= a;
    layer6_outputs(9021) <= not a;
    layer6_outputs(9022) <= not a;
    layer6_outputs(9023) <= not b;
    layer6_outputs(9024) <= a;
    layer6_outputs(9025) <= a or b;
    layer6_outputs(9026) <= a;
    layer6_outputs(9027) <= b and not a;
    layer6_outputs(9028) <= not (a xor b);
    layer6_outputs(9029) <= not b;
    layer6_outputs(9030) <= not a;
    layer6_outputs(9031) <= not (a or b);
    layer6_outputs(9032) <= not a;
    layer6_outputs(9033) <= not a;
    layer6_outputs(9034) <= not a;
    layer6_outputs(9035) <= b;
    layer6_outputs(9036) <= a and not b;
    layer6_outputs(9037) <= a and not b;
    layer6_outputs(9038) <= not a;
    layer6_outputs(9039) <= not a or b;
    layer6_outputs(9040) <= '1';
    layer6_outputs(9041) <= b;
    layer6_outputs(9042) <= not b or a;
    layer6_outputs(9043) <= not b or a;
    layer6_outputs(9044) <= not b;
    layer6_outputs(9045) <= a or b;
    layer6_outputs(9046) <= not (a xor b);
    layer6_outputs(9047) <= not (a and b);
    layer6_outputs(9048) <= not b;
    layer6_outputs(9049) <= a xor b;
    layer6_outputs(9050) <= b;
    layer6_outputs(9051) <= not (a and b);
    layer6_outputs(9052) <= b;
    layer6_outputs(9053) <= a xor b;
    layer6_outputs(9054) <= a or b;
    layer6_outputs(9055) <= not b;
    layer6_outputs(9056) <= not (a and b);
    layer6_outputs(9057) <= not (a or b);
    layer6_outputs(9058) <= not (a xor b);
    layer6_outputs(9059) <= a and b;
    layer6_outputs(9060) <= not a or b;
    layer6_outputs(9061) <= not (a xor b);
    layer6_outputs(9062) <= a;
    layer6_outputs(9063) <= not (a xor b);
    layer6_outputs(9064) <= not (a xor b);
    layer6_outputs(9065) <= not (a or b);
    layer6_outputs(9066) <= b and not a;
    layer6_outputs(9067) <= a;
    layer6_outputs(9068) <= b;
    layer6_outputs(9069) <= a;
    layer6_outputs(9070) <= not (a xor b);
    layer6_outputs(9071) <= a and not b;
    layer6_outputs(9072) <= not a;
    layer6_outputs(9073) <= a and not b;
    layer6_outputs(9074) <= a and not b;
    layer6_outputs(9075) <= a;
    layer6_outputs(9076) <= not a or b;
    layer6_outputs(9077) <= a or b;
    layer6_outputs(9078) <= not (a or b);
    layer6_outputs(9079) <= b;
    layer6_outputs(9080) <= a and b;
    layer6_outputs(9081) <= a;
    layer6_outputs(9082) <= a xor b;
    layer6_outputs(9083) <= not b;
    layer6_outputs(9084) <= not (a xor b);
    layer6_outputs(9085) <= a;
    layer6_outputs(9086) <= not (a xor b);
    layer6_outputs(9087) <= a xor b;
    layer6_outputs(9088) <= b;
    layer6_outputs(9089) <= b;
    layer6_outputs(9090) <= b;
    layer6_outputs(9091) <= a xor b;
    layer6_outputs(9092) <= a;
    layer6_outputs(9093) <= a or b;
    layer6_outputs(9094) <= not (a or b);
    layer6_outputs(9095) <= not (a xor b);
    layer6_outputs(9096) <= b and not a;
    layer6_outputs(9097) <= a xor b;
    layer6_outputs(9098) <= not b or a;
    layer6_outputs(9099) <= not b;
    layer6_outputs(9100) <= not (a xor b);
    layer6_outputs(9101) <= not (a xor b);
    layer6_outputs(9102) <= not a;
    layer6_outputs(9103) <= a or b;
    layer6_outputs(9104) <= '0';
    layer6_outputs(9105) <= a xor b;
    layer6_outputs(9106) <= not a;
    layer6_outputs(9107) <= a xor b;
    layer6_outputs(9108) <= not b or a;
    layer6_outputs(9109) <= not b or a;
    layer6_outputs(9110) <= not (a or b);
    layer6_outputs(9111) <= a and b;
    layer6_outputs(9112) <= a and b;
    layer6_outputs(9113) <= b;
    layer6_outputs(9114) <= a;
    layer6_outputs(9115) <= b;
    layer6_outputs(9116) <= a;
    layer6_outputs(9117) <= a or b;
    layer6_outputs(9118) <= not b;
    layer6_outputs(9119) <= a;
    layer6_outputs(9120) <= not a;
    layer6_outputs(9121) <= not (a xor b);
    layer6_outputs(9122) <= not b;
    layer6_outputs(9123) <= not (a and b);
    layer6_outputs(9124) <= a;
    layer6_outputs(9125) <= not a;
    layer6_outputs(9126) <= not a;
    layer6_outputs(9127) <= not b;
    layer6_outputs(9128) <= not b;
    layer6_outputs(9129) <= a xor b;
    layer6_outputs(9130) <= b and not a;
    layer6_outputs(9131) <= not (a xor b);
    layer6_outputs(9132) <= not (a and b);
    layer6_outputs(9133) <= not (a and b);
    layer6_outputs(9134) <= not (a xor b);
    layer6_outputs(9135) <= a xor b;
    layer6_outputs(9136) <= a;
    layer6_outputs(9137) <= b;
    layer6_outputs(9138) <= not (a xor b);
    layer6_outputs(9139) <= not (a or b);
    layer6_outputs(9140) <= b;
    layer6_outputs(9141) <= a and not b;
    layer6_outputs(9142) <= b and not a;
    layer6_outputs(9143) <= a xor b;
    layer6_outputs(9144) <= a xor b;
    layer6_outputs(9145) <= a xor b;
    layer6_outputs(9146) <= not a;
    layer6_outputs(9147) <= a and not b;
    layer6_outputs(9148) <= a;
    layer6_outputs(9149) <= not a;
    layer6_outputs(9150) <= a;
    layer6_outputs(9151) <= a xor b;
    layer6_outputs(9152) <= a and not b;
    layer6_outputs(9153) <= b;
    layer6_outputs(9154) <= a;
    layer6_outputs(9155) <= a;
    layer6_outputs(9156) <= not (a or b);
    layer6_outputs(9157) <= not (a xor b);
    layer6_outputs(9158) <= not a;
    layer6_outputs(9159) <= not (a or b);
    layer6_outputs(9160) <= not (a and b);
    layer6_outputs(9161) <= not (a xor b);
    layer6_outputs(9162) <= a or b;
    layer6_outputs(9163) <= a xor b;
    layer6_outputs(9164) <= not b;
    layer6_outputs(9165) <= not a;
    layer6_outputs(9166) <= not b;
    layer6_outputs(9167) <= not a;
    layer6_outputs(9168) <= a xor b;
    layer6_outputs(9169) <= not a;
    layer6_outputs(9170) <= a;
    layer6_outputs(9171) <= not a or b;
    layer6_outputs(9172) <= not (a xor b);
    layer6_outputs(9173) <= b;
    layer6_outputs(9174) <= not b;
    layer6_outputs(9175) <= '0';
    layer6_outputs(9176) <= not (a xor b);
    layer6_outputs(9177) <= a;
    layer6_outputs(9178) <= not a;
    layer6_outputs(9179) <= a xor b;
    layer6_outputs(9180) <= not a;
    layer6_outputs(9181) <= not b;
    layer6_outputs(9182) <= b;
    layer6_outputs(9183) <= a xor b;
    layer6_outputs(9184) <= not a;
    layer6_outputs(9185) <= not b;
    layer6_outputs(9186) <= b;
    layer6_outputs(9187) <= not b;
    layer6_outputs(9188) <= a;
    layer6_outputs(9189) <= a or b;
    layer6_outputs(9190) <= not a;
    layer6_outputs(9191) <= a;
    layer6_outputs(9192) <= b;
    layer6_outputs(9193) <= b and not a;
    layer6_outputs(9194) <= not a;
    layer6_outputs(9195) <= a xor b;
    layer6_outputs(9196) <= a xor b;
    layer6_outputs(9197) <= b and not a;
    layer6_outputs(9198) <= not b;
    layer6_outputs(9199) <= not a;
    layer6_outputs(9200) <= b;
    layer6_outputs(9201) <= b;
    layer6_outputs(9202) <= a xor b;
    layer6_outputs(9203) <= not a;
    layer6_outputs(9204) <= not (a xor b);
    layer6_outputs(9205) <= a;
    layer6_outputs(9206) <= a;
    layer6_outputs(9207) <= a;
    layer6_outputs(9208) <= a xor b;
    layer6_outputs(9209) <= b;
    layer6_outputs(9210) <= a and not b;
    layer6_outputs(9211) <= a and b;
    layer6_outputs(9212) <= not (a and b);
    layer6_outputs(9213) <= b and not a;
    layer6_outputs(9214) <= not (a and b);
    layer6_outputs(9215) <= a or b;
    layer6_outputs(9216) <= a xor b;
    layer6_outputs(9217) <= not a or b;
    layer6_outputs(9218) <= b;
    layer6_outputs(9219) <= not (a xor b);
    layer6_outputs(9220) <= not a;
    layer6_outputs(9221) <= a;
    layer6_outputs(9222) <= a or b;
    layer6_outputs(9223) <= a xor b;
    layer6_outputs(9224) <= a or b;
    layer6_outputs(9225) <= b;
    layer6_outputs(9226) <= b;
    layer6_outputs(9227) <= a;
    layer6_outputs(9228) <= not b or a;
    layer6_outputs(9229) <= not b or a;
    layer6_outputs(9230) <= not (a xor b);
    layer6_outputs(9231) <= not b or a;
    layer6_outputs(9232) <= a xor b;
    layer6_outputs(9233) <= not a or b;
    layer6_outputs(9234) <= not b;
    layer6_outputs(9235) <= a;
    layer6_outputs(9236) <= not a;
    layer6_outputs(9237) <= a xor b;
    layer6_outputs(9238) <= not a;
    layer6_outputs(9239) <= not b or a;
    layer6_outputs(9240) <= a xor b;
    layer6_outputs(9241) <= not (a and b);
    layer6_outputs(9242) <= '0';
    layer6_outputs(9243) <= not (a xor b);
    layer6_outputs(9244) <= not a;
    layer6_outputs(9245) <= a;
    layer6_outputs(9246) <= a xor b;
    layer6_outputs(9247) <= not (a xor b);
    layer6_outputs(9248) <= a;
    layer6_outputs(9249) <= not b;
    layer6_outputs(9250) <= not (a and b);
    layer6_outputs(9251) <= not a;
    layer6_outputs(9252) <= not (a xor b);
    layer6_outputs(9253) <= a xor b;
    layer6_outputs(9254) <= not a;
    layer6_outputs(9255) <= a and not b;
    layer6_outputs(9256) <= a;
    layer6_outputs(9257) <= a;
    layer6_outputs(9258) <= a and not b;
    layer6_outputs(9259) <= b;
    layer6_outputs(9260) <= not a;
    layer6_outputs(9261) <= b;
    layer6_outputs(9262) <= not (a xor b);
    layer6_outputs(9263) <= not (a and b);
    layer6_outputs(9264) <= a;
    layer6_outputs(9265) <= b;
    layer6_outputs(9266) <= b;
    layer6_outputs(9267) <= not b;
    layer6_outputs(9268) <= b and not a;
    layer6_outputs(9269) <= not b or a;
    layer6_outputs(9270) <= not (a or b);
    layer6_outputs(9271) <= a xor b;
    layer6_outputs(9272) <= b and not a;
    layer6_outputs(9273) <= a;
    layer6_outputs(9274) <= not a;
    layer6_outputs(9275) <= a;
    layer6_outputs(9276) <= a and not b;
    layer6_outputs(9277) <= a xor b;
    layer6_outputs(9278) <= not b;
    layer6_outputs(9279) <= not (a or b);
    layer6_outputs(9280) <= a or b;
    layer6_outputs(9281) <= not b;
    layer6_outputs(9282) <= b;
    layer6_outputs(9283) <= not a;
    layer6_outputs(9284) <= not a;
    layer6_outputs(9285) <= not b;
    layer6_outputs(9286) <= not a;
    layer6_outputs(9287) <= b;
    layer6_outputs(9288) <= not b or a;
    layer6_outputs(9289) <= not (a xor b);
    layer6_outputs(9290) <= not b;
    layer6_outputs(9291) <= '0';
    layer6_outputs(9292) <= a and b;
    layer6_outputs(9293) <= not a or b;
    layer6_outputs(9294) <= a xor b;
    layer6_outputs(9295) <= a xor b;
    layer6_outputs(9296) <= not (a or b);
    layer6_outputs(9297) <= b;
    layer6_outputs(9298) <= not a;
    layer6_outputs(9299) <= not (a xor b);
    layer6_outputs(9300) <= not b;
    layer6_outputs(9301) <= a xor b;
    layer6_outputs(9302) <= b;
    layer6_outputs(9303) <= a and not b;
    layer6_outputs(9304) <= not a or b;
    layer6_outputs(9305) <= b and not a;
    layer6_outputs(9306) <= a xor b;
    layer6_outputs(9307) <= a;
    layer6_outputs(9308) <= a;
    layer6_outputs(9309) <= not a;
    layer6_outputs(9310) <= a xor b;
    layer6_outputs(9311) <= not a or b;
    layer6_outputs(9312) <= not b or a;
    layer6_outputs(9313) <= not (a and b);
    layer6_outputs(9314) <= not b;
    layer6_outputs(9315) <= not b;
    layer6_outputs(9316) <= a xor b;
    layer6_outputs(9317) <= not a;
    layer6_outputs(9318) <= a and not b;
    layer6_outputs(9319) <= not (a or b);
    layer6_outputs(9320) <= not (a and b);
    layer6_outputs(9321) <= not b;
    layer6_outputs(9322) <= not (a or b);
    layer6_outputs(9323) <= a or b;
    layer6_outputs(9324) <= not a;
    layer6_outputs(9325) <= not b;
    layer6_outputs(9326) <= a xor b;
    layer6_outputs(9327) <= a xor b;
    layer6_outputs(9328) <= not b;
    layer6_outputs(9329) <= not b or a;
    layer6_outputs(9330) <= b and not a;
    layer6_outputs(9331) <= not (a xor b);
    layer6_outputs(9332) <= b and not a;
    layer6_outputs(9333) <= a;
    layer6_outputs(9334) <= not a;
    layer6_outputs(9335) <= b;
    layer6_outputs(9336) <= not (a xor b);
    layer6_outputs(9337) <= not (a and b);
    layer6_outputs(9338) <= not (a xor b);
    layer6_outputs(9339) <= a;
    layer6_outputs(9340) <= b and not a;
    layer6_outputs(9341) <= not (a xor b);
    layer6_outputs(9342) <= not (a and b);
    layer6_outputs(9343) <= not a or b;
    layer6_outputs(9344) <= not b or a;
    layer6_outputs(9345) <= not (a and b);
    layer6_outputs(9346) <= b;
    layer6_outputs(9347) <= not a;
    layer6_outputs(9348) <= not b;
    layer6_outputs(9349) <= not b;
    layer6_outputs(9350) <= b;
    layer6_outputs(9351) <= b and not a;
    layer6_outputs(9352) <= not (a xor b);
    layer6_outputs(9353) <= not a or b;
    layer6_outputs(9354) <= a or b;
    layer6_outputs(9355) <= a;
    layer6_outputs(9356) <= not b;
    layer6_outputs(9357) <= a xor b;
    layer6_outputs(9358) <= b;
    layer6_outputs(9359) <= a or b;
    layer6_outputs(9360) <= not (a or b);
    layer6_outputs(9361) <= a;
    layer6_outputs(9362) <= not a;
    layer6_outputs(9363) <= b;
    layer6_outputs(9364) <= a;
    layer6_outputs(9365) <= not (a and b);
    layer6_outputs(9366) <= not b or a;
    layer6_outputs(9367) <= not (a xor b);
    layer6_outputs(9368) <= not (a xor b);
    layer6_outputs(9369) <= a and b;
    layer6_outputs(9370) <= not (a and b);
    layer6_outputs(9371) <= not a;
    layer6_outputs(9372) <= a xor b;
    layer6_outputs(9373) <= a;
    layer6_outputs(9374) <= not (a xor b);
    layer6_outputs(9375) <= not (a xor b);
    layer6_outputs(9376) <= a or b;
    layer6_outputs(9377) <= not b;
    layer6_outputs(9378) <= b and not a;
    layer6_outputs(9379) <= not b;
    layer6_outputs(9380) <= not a;
    layer6_outputs(9381) <= not b;
    layer6_outputs(9382) <= a xor b;
    layer6_outputs(9383) <= not a;
    layer6_outputs(9384) <= b and not a;
    layer6_outputs(9385) <= a and b;
    layer6_outputs(9386) <= b;
    layer6_outputs(9387) <= not b;
    layer6_outputs(9388) <= b and not a;
    layer6_outputs(9389) <= not a;
    layer6_outputs(9390) <= not a or b;
    layer6_outputs(9391) <= not b or a;
    layer6_outputs(9392) <= not b;
    layer6_outputs(9393) <= not (a and b);
    layer6_outputs(9394) <= not b;
    layer6_outputs(9395) <= a;
    layer6_outputs(9396) <= b and not a;
    layer6_outputs(9397) <= a;
    layer6_outputs(9398) <= not b;
    layer6_outputs(9399) <= not a;
    layer6_outputs(9400) <= '0';
    layer6_outputs(9401) <= not (a xor b);
    layer6_outputs(9402) <= not a;
    layer6_outputs(9403) <= b and not a;
    layer6_outputs(9404) <= not b or a;
    layer6_outputs(9405) <= not b or a;
    layer6_outputs(9406) <= a xor b;
    layer6_outputs(9407) <= a;
    layer6_outputs(9408) <= not a or b;
    layer6_outputs(9409) <= b;
    layer6_outputs(9410) <= b and not a;
    layer6_outputs(9411) <= not a;
    layer6_outputs(9412) <= not b;
    layer6_outputs(9413) <= not b;
    layer6_outputs(9414) <= a;
    layer6_outputs(9415) <= not a;
    layer6_outputs(9416) <= a and not b;
    layer6_outputs(9417) <= not (a or b);
    layer6_outputs(9418) <= not b;
    layer6_outputs(9419) <= a;
    layer6_outputs(9420) <= a xor b;
    layer6_outputs(9421) <= a xor b;
    layer6_outputs(9422) <= b;
    layer6_outputs(9423) <= b and not a;
    layer6_outputs(9424) <= a and not b;
    layer6_outputs(9425) <= b;
    layer6_outputs(9426) <= not b;
    layer6_outputs(9427) <= not b;
    layer6_outputs(9428) <= not a;
    layer6_outputs(9429) <= not (a xor b);
    layer6_outputs(9430) <= not b;
    layer6_outputs(9431) <= not (a xor b);
    layer6_outputs(9432) <= a xor b;
    layer6_outputs(9433) <= not (a xor b);
    layer6_outputs(9434) <= b;
    layer6_outputs(9435) <= not (a xor b);
    layer6_outputs(9436) <= not (a xor b);
    layer6_outputs(9437) <= b;
    layer6_outputs(9438) <= not (a or b);
    layer6_outputs(9439) <= not (a or b);
    layer6_outputs(9440) <= not a;
    layer6_outputs(9441) <= a xor b;
    layer6_outputs(9442) <= a xor b;
    layer6_outputs(9443) <= b and not a;
    layer6_outputs(9444) <= not b;
    layer6_outputs(9445) <= not (a or b);
    layer6_outputs(9446) <= not b;
    layer6_outputs(9447) <= a xor b;
    layer6_outputs(9448) <= not b;
    layer6_outputs(9449) <= not a;
    layer6_outputs(9450) <= a xor b;
    layer6_outputs(9451) <= not b;
    layer6_outputs(9452) <= b;
    layer6_outputs(9453) <= a;
    layer6_outputs(9454) <= not b;
    layer6_outputs(9455) <= not a or b;
    layer6_outputs(9456) <= a;
    layer6_outputs(9457) <= not (a or b);
    layer6_outputs(9458) <= a and not b;
    layer6_outputs(9459) <= a xor b;
    layer6_outputs(9460) <= not b or a;
    layer6_outputs(9461) <= not b;
    layer6_outputs(9462) <= a or b;
    layer6_outputs(9463) <= not (a xor b);
    layer6_outputs(9464) <= a or b;
    layer6_outputs(9465) <= a and not b;
    layer6_outputs(9466) <= not (a xor b);
    layer6_outputs(9467) <= b;
    layer6_outputs(9468) <= not b or a;
    layer6_outputs(9469) <= a or b;
    layer6_outputs(9470) <= a or b;
    layer6_outputs(9471) <= a;
    layer6_outputs(9472) <= b;
    layer6_outputs(9473) <= a and b;
    layer6_outputs(9474) <= not a;
    layer6_outputs(9475) <= not (a or b);
    layer6_outputs(9476) <= a;
    layer6_outputs(9477) <= a xor b;
    layer6_outputs(9478) <= not b;
    layer6_outputs(9479) <= not b or a;
    layer6_outputs(9480) <= not a;
    layer6_outputs(9481) <= a and not b;
    layer6_outputs(9482) <= not (a xor b);
    layer6_outputs(9483) <= not b;
    layer6_outputs(9484) <= not a;
    layer6_outputs(9485) <= a;
    layer6_outputs(9486) <= not a or b;
    layer6_outputs(9487) <= not b;
    layer6_outputs(9488) <= not (a xor b);
    layer6_outputs(9489) <= b;
    layer6_outputs(9490) <= not (a or b);
    layer6_outputs(9491) <= a xor b;
    layer6_outputs(9492) <= a or b;
    layer6_outputs(9493) <= a xor b;
    layer6_outputs(9494) <= a;
    layer6_outputs(9495) <= a;
    layer6_outputs(9496) <= a and b;
    layer6_outputs(9497) <= a xor b;
    layer6_outputs(9498) <= b;
    layer6_outputs(9499) <= not b;
    layer6_outputs(9500) <= a;
    layer6_outputs(9501) <= not b or a;
    layer6_outputs(9502) <= a xor b;
    layer6_outputs(9503) <= a and not b;
    layer6_outputs(9504) <= not (a xor b);
    layer6_outputs(9505) <= a;
    layer6_outputs(9506) <= a;
    layer6_outputs(9507) <= a or b;
    layer6_outputs(9508) <= not a;
    layer6_outputs(9509) <= not a;
    layer6_outputs(9510) <= not a;
    layer6_outputs(9511) <= not a or b;
    layer6_outputs(9512) <= a;
    layer6_outputs(9513) <= a xor b;
    layer6_outputs(9514) <= a and b;
    layer6_outputs(9515) <= not (a and b);
    layer6_outputs(9516) <= not b;
    layer6_outputs(9517) <= a;
    layer6_outputs(9518) <= a xor b;
    layer6_outputs(9519) <= b;
    layer6_outputs(9520) <= not a or b;
    layer6_outputs(9521) <= b and not a;
    layer6_outputs(9522) <= not a;
    layer6_outputs(9523) <= b;
    layer6_outputs(9524) <= not a;
    layer6_outputs(9525) <= not a;
    layer6_outputs(9526) <= not (a and b);
    layer6_outputs(9527) <= not b;
    layer6_outputs(9528) <= a xor b;
    layer6_outputs(9529) <= a;
    layer6_outputs(9530) <= a xor b;
    layer6_outputs(9531) <= not a;
    layer6_outputs(9532) <= not a;
    layer6_outputs(9533) <= a xor b;
    layer6_outputs(9534) <= a;
    layer6_outputs(9535) <= b;
    layer6_outputs(9536) <= a xor b;
    layer6_outputs(9537) <= not a or b;
    layer6_outputs(9538) <= not b or a;
    layer6_outputs(9539) <= not b;
    layer6_outputs(9540) <= a;
    layer6_outputs(9541) <= not (a xor b);
    layer6_outputs(9542) <= a;
    layer6_outputs(9543) <= not (a and b);
    layer6_outputs(9544) <= a and b;
    layer6_outputs(9545) <= a and not b;
    layer6_outputs(9546) <= not a;
    layer6_outputs(9547) <= not b or a;
    layer6_outputs(9548) <= b and not a;
    layer6_outputs(9549) <= a;
    layer6_outputs(9550) <= not b;
    layer6_outputs(9551) <= a;
    layer6_outputs(9552) <= a;
    layer6_outputs(9553) <= a or b;
    layer6_outputs(9554) <= a xor b;
    layer6_outputs(9555) <= b and not a;
    layer6_outputs(9556) <= not b;
    layer6_outputs(9557) <= a or b;
    layer6_outputs(9558) <= a;
    layer6_outputs(9559) <= a;
    layer6_outputs(9560) <= b;
    layer6_outputs(9561) <= not (a xor b);
    layer6_outputs(9562) <= a xor b;
    layer6_outputs(9563) <= b;
    layer6_outputs(9564) <= not (a xor b);
    layer6_outputs(9565) <= a or b;
    layer6_outputs(9566) <= a or b;
    layer6_outputs(9567) <= a xor b;
    layer6_outputs(9568) <= b;
    layer6_outputs(9569) <= not a;
    layer6_outputs(9570) <= not b;
    layer6_outputs(9571) <= a and not b;
    layer6_outputs(9572) <= not a;
    layer6_outputs(9573) <= not a;
    layer6_outputs(9574) <= a or b;
    layer6_outputs(9575) <= b;
    layer6_outputs(9576) <= b;
    layer6_outputs(9577) <= b;
    layer6_outputs(9578) <= b and not a;
    layer6_outputs(9579) <= a xor b;
    layer6_outputs(9580) <= not a;
    layer6_outputs(9581) <= a and b;
    layer6_outputs(9582) <= b and not a;
    layer6_outputs(9583) <= not b;
    layer6_outputs(9584) <= b;
    layer6_outputs(9585) <= a or b;
    layer6_outputs(9586) <= a or b;
    layer6_outputs(9587) <= not a;
    layer6_outputs(9588) <= not a;
    layer6_outputs(9589) <= a and not b;
    layer6_outputs(9590) <= '0';
    layer6_outputs(9591) <= a or b;
    layer6_outputs(9592) <= not (a xor b);
    layer6_outputs(9593) <= a or b;
    layer6_outputs(9594) <= a xor b;
    layer6_outputs(9595) <= not (a xor b);
    layer6_outputs(9596) <= not a;
    layer6_outputs(9597) <= b;
    layer6_outputs(9598) <= a;
    layer6_outputs(9599) <= not (a xor b);
    layer6_outputs(9600) <= b;
    layer6_outputs(9601) <= a or b;
    layer6_outputs(9602) <= not a;
    layer6_outputs(9603) <= b and not a;
    layer6_outputs(9604) <= not b;
    layer6_outputs(9605) <= a;
    layer6_outputs(9606) <= not b;
    layer6_outputs(9607) <= a;
    layer6_outputs(9608) <= a;
    layer6_outputs(9609) <= b and not a;
    layer6_outputs(9610) <= not (a and b);
    layer6_outputs(9611) <= a;
    layer6_outputs(9612) <= a;
    layer6_outputs(9613) <= not (a xor b);
    layer6_outputs(9614) <= a or b;
    layer6_outputs(9615) <= a xor b;
    layer6_outputs(9616) <= not a;
    layer6_outputs(9617) <= a xor b;
    layer6_outputs(9618) <= a;
    layer6_outputs(9619) <= not a or b;
    layer6_outputs(9620) <= not (a and b);
    layer6_outputs(9621) <= not b;
    layer6_outputs(9622) <= not (a xor b);
    layer6_outputs(9623) <= not b or a;
    layer6_outputs(9624) <= a xor b;
    layer6_outputs(9625) <= a;
    layer6_outputs(9626) <= a;
    layer6_outputs(9627) <= b and not a;
    layer6_outputs(9628) <= not b or a;
    layer6_outputs(9629) <= a xor b;
    layer6_outputs(9630) <= not b;
    layer6_outputs(9631) <= b;
    layer6_outputs(9632) <= a;
    layer6_outputs(9633) <= not a;
    layer6_outputs(9634) <= a and b;
    layer6_outputs(9635) <= not b;
    layer6_outputs(9636) <= a;
    layer6_outputs(9637) <= a;
    layer6_outputs(9638) <= not (a xor b);
    layer6_outputs(9639) <= not b;
    layer6_outputs(9640) <= a or b;
    layer6_outputs(9641) <= not b or a;
    layer6_outputs(9642) <= not (a and b);
    layer6_outputs(9643) <= not a;
    layer6_outputs(9644) <= a or b;
    layer6_outputs(9645) <= not (a xor b);
    layer6_outputs(9646) <= a xor b;
    layer6_outputs(9647) <= not b or a;
    layer6_outputs(9648) <= a and not b;
    layer6_outputs(9649) <= not a;
    layer6_outputs(9650) <= a xor b;
    layer6_outputs(9651) <= b and not a;
    layer6_outputs(9652) <= a;
    layer6_outputs(9653) <= b;
    layer6_outputs(9654) <= b and not a;
    layer6_outputs(9655) <= b;
    layer6_outputs(9656) <= not (a xor b);
    layer6_outputs(9657) <= not (a xor b);
    layer6_outputs(9658) <= b;
    layer6_outputs(9659) <= not a;
    layer6_outputs(9660) <= not (a xor b);
    layer6_outputs(9661) <= a or b;
    layer6_outputs(9662) <= a;
    layer6_outputs(9663) <= b and not a;
    layer6_outputs(9664) <= not b;
    layer6_outputs(9665) <= a and not b;
    layer6_outputs(9666) <= not (a and b);
    layer6_outputs(9667) <= not a;
    layer6_outputs(9668) <= not (a xor b);
    layer6_outputs(9669) <= b;
    layer6_outputs(9670) <= a;
    layer6_outputs(9671) <= not b or a;
    layer6_outputs(9672) <= a;
    layer6_outputs(9673) <= not a;
    layer6_outputs(9674) <= not b;
    layer6_outputs(9675) <= not (a xor b);
    layer6_outputs(9676) <= not b;
    layer6_outputs(9677) <= a xor b;
    layer6_outputs(9678) <= a;
    layer6_outputs(9679) <= not (a xor b);
    layer6_outputs(9680) <= b;
    layer6_outputs(9681) <= a;
    layer6_outputs(9682) <= not (a xor b);
    layer6_outputs(9683) <= not a or b;
    layer6_outputs(9684) <= not a;
    layer6_outputs(9685) <= b;
    layer6_outputs(9686) <= not a;
    layer6_outputs(9687) <= b and not a;
    layer6_outputs(9688) <= b;
    layer6_outputs(9689) <= a and b;
    layer6_outputs(9690) <= a xor b;
    layer6_outputs(9691) <= a xor b;
    layer6_outputs(9692) <= not a or b;
    layer6_outputs(9693) <= b;
    layer6_outputs(9694) <= a;
    layer6_outputs(9695) <= a and not b;
    layer6_outputs(9696) <= not a;
    layer6_outputs(9697) <= not (a and b);
    layer6_outputs(9698) <= a and not b;
    layer6_outputs(9699) <= a;
    layer6_outputs(9700) <= a and b;
    layer6_outputs(9701) <= a or b;
    layer6_outputs(9702) <= not a;
    layer6_outputs(9703) <= a and not b;
    layer6_outputs(9704) <= b;
    layer6_outputs(9705) <= not a;
    layer6_outputs(9706) <= not a;
    layer6_outputs(9707) <= a and b;
    layer6_outputs(9708) <= b;
    layer6_outputs(9709) <= b;
    layer6_outputs(9710) <= a or b;
    layer6_outputs(9711) <= not a;
    layer6_outputs(9712) <= a and not b;
    layer6_outputs(9713) <= a;
    layer6_outputs(9714) <= not (a xor b);
    layer6_outputs(9715) <= not (a xor b);
    layer6_outputs(9716) <= not (a and b);
    layer6_outputs(9717) <= a xor b;
    layer6_outputs(9718) <= not a;
    layer6_outputs(9719) <= a xor b;
    layer6_outputs(9720) <= not (a xor b);
    layer6_outputs(9721) <= a;
    layer6_outputs(9722) <= a;
    layer6_outputs(9723) <= not (a xor b);
    layer6_outputs(9724) <= a and not b;
    layer6_outputs(9725) <= a;
    layer6_outputs(9726) <= b and not a;
    layer6_outputs(9727) <= not a;
    layer6_outputs(9728) <= a and not b;
    layer6_outputs(9729) <= not (a and b);
    layer6_outputs(9730) <= b and not a;
    layer6_outputs(9731) <= not (a xor b);
    layer6_outputs(9732) <= not a;
    layer6_outputs(9733) <= not b;
    layer6_outputs(9734) <= not (a xor b);
    layer6_outputs(9735) <= not b;
    layer6_outputs(9736) <= a or b;
    layer6_outputs(9737) <= a xor b;
    layer6_outputs(9738) <= not (a and b);
    layer6_outputs(9739) <= not b;
    layer6_outputs(9740) <= not b;
    layer6_outputs(9741) <= not b or a;
    layer6_outputs(9742) <= not (a xor b);
    layer6_outputs(9743) <= not (a xor b);
    layer6_outputs(9744) <= a;
    layer6_outputs(9745) <= not b;
    layer6_outputs(9746) <= b;
    layer6_outputs(9747) <= not b;
    layer6_outputs(9748) <= not (a or b);
    layer6_outputs(9749) <= a;
    layer6_outputs(9750) <= not (a xor b);
    layer6_outputs(9751) <= a;
    layer6_outputs(9752) <= a and not b;
    layer6_outputs(9753) <= a and b;
    layer6_outputs(9754) <= not (a xor b);
    layer6_outputs(9755) <= not b;
    layer6_outputs(9756) <= not (a xor b);
    layer6_outputs(9757) <= a;
    layer6_outputs(9758) <= a xor b;
    layer6_outputs(9759) <= a and not b;
    layer6_outputs(9760) <= a;
    layer6_outputs(9761) <= not b or a;
    layer6_outputs(9762) <= b and not a;
    layer6_outputs(9763) <= not (a xor b);
    layer6_outputs(9764) <= not a or b;
    layer6_outputs(9765) <= not a;
    layer6_outputs(9766) <= not b;
    layer6_outputs(9767) <= not b;
    layer6_outputs(9768) <= a and b;
    layer6_outputs(9769) <= a or b;
    layer6_outputs(9770) <= not a;
    layer6_outputs(9771) <= not (a or b);
    layer6_outputs(9772) <= b;
    layer6_outputs(9773) <= not a or b;
    layer6_outputs(9774) <= not b;
    layer6_outputs(9775) <= a xor b;
    layer6_outputs(9776) <= a xor b;
    layer6_outputs(9777) <= not b or a;
    layer6_outputs(9778) <= not (a xor b);
    layer6_outputs(9779) <= a xor b;
    layer6_outputs(9780) <= not b;
    layer6_outputs(9781) <= b;
    layer6_outputs(9782) <= not (a and b);
    layer6_outputs(9783) <= a and b;
    layer6_outputs(9784) <= not b or a;
    layer6_outputs(9785) <= a;
    layer6_outputs(9786) <= b and not a;
    layer6_outputs(9787) <= b;
    layer6_outputs(9788) <= not a;
    layer6_outputs(9789) <= a;
    layer6_outputs(9790) <= a and b;
    layer6_outputs(9791) <= not (a xor b);
    layer6_outputs(9792) <= not b;
    layer6_outputs(9793) <= b;
    layer6_outputs(9794) <= not a;
    layer6_outputs(9795) <= a;
    layer6_outputs(9796) <= not b or a;
    layer6_outputs(9797) <= not b;
    layer6_outputs(9798) <= not (a or b);
    layer6_outputs(9799) <= not b;
    layer6_outputs(9800) <= '0';
    layer6_outputs(9801) <= b;
    layer6_outputs(9802) <= a;
    layer6_outputs(9803) <= a xor b;
    layer6_outputs(9804) <= not b;
    layer6_outputs(9805) <= b;
    layer6_outputs(9806) <= a and b;
    layer6_outputs(9807) <= a xor b;
    layer6_outputs(9808) <= not (a xor b);
    layer6_outputs(9809) <= a;
    layer6_outputs(9810) <= not b or a;
    layer6_outputs(9811) <= not a;
    layer6_outputs(9812) <= a;
    layer6_outputs(9813) <= not (a xor b);
    layer6_outputs(9814) <= not b;
    layer6_outputs(9815) <= not b or a;
    layer6_outputs(9816) <= not (a xor b);
    layer6_outputs(9817) <= not (a and b);
    layer6_outputs(9818) <= b;
    layer6_outputs(9819) <= b;
    layer6_outputs(9820) <= '0';
    layer6_outputs(9821) <= b;
    layer6_outputs(9822) <= a and not b;
    layer6_outputs(9823) <= b;
    layer6_outputs(9824) <= not a or b;
    layer6_outputs(9825) <= a;
    layer6_outputs(9826) <= a and not b;
    layer6_outputs(9827) <= not (a xor b);
    layer6_outputs(9828) <= a xor b;
    layer6_outputs(9829) <= not a;
    layer6_outputs(9830) <= not (a and b);
    layer6_outputs(9831) <= not (a xor b);
    layer6_outputs(9832) <= not b;
    layer6_outputs(9833) <= b and not a;
    layer6_outputs(9834) <= not a;
    layer6_outputs(9835) <= not (a or b);
    layer6_outputs(9836) <= b and not a;
    layer6_outputs(9837) <= not (a xor b);
    layer6_outputs(9838) <= a or b;
    layer6_outputs(9839) <= a or b;
    layer6_outputs(9840) <= a or b;
    layer6_outputs(9841) <= not b;
    layer6_outputs(9842) <= not a or b;
    layer6_outputs(9843) <= not (a xor b);
    layer6_outputs(9844) <= a;
    layer6_outputs(9845) <= b;
    layer6_outputs(9846) <= not (a xor b);
    layer6_outputs(9847) <= b and not a;
    layer6_outputs(9848) <= a and b;
    layer6_outputs(9849) <= not a or b;
    layer6_outputs(9850) <= not (a xor b);
    layer6_outputs(9851) <= not b or a;
    layer6_outputs(9852) <= a and not b;
    layer6_outputs(9853) <= a;
    layer6_outputs(9854) <= not b;
    layer6_outputs(9855) <= a;
    layer6_outputs(9856) <= a and not b;
    layer6_outputs(9857) <= a or b;
    layer6_outputs(9858) <= not (a xor b);
    layer6_outputs(9859) <= not b or a;
    layer6_outputs(9860) <= not (a xor b);
    layer6_outputs(9861) <= not a or b;
    layer6_outputs(9862) <= a xor b;
    layer6_outputs(9863) <= not b;
    layer6_outputs(9864) <= b;
    layer6_outputs(9865) <= a xor b;
    layer6_outputs(9866) <= a;
    layer6_outputs(9867) <= a and b;
    layer6_outputs(9868) <= not a or b;
    layer6_outputs(9869) <= not a or b;
    layer6_outputs(9870) <= not (a and b);
    layer6_outputs(9871) <= not a or b;
    layer6_outputs(9872) <= a and b;
    layer6_outputs(9873) <= a xor b;
    layer6_outputs(9874) <= b;
    layer6_outputs(9875) <= not (a or b);
    layer6_outputs(9876) <= not (a and b);
    layer6_outputs(9877) <= not b;
    layer6_outputs(9878) <= a;
    layer6_outputs(9879) <= not (a and b);
    layer6_outputs(9880) <= not (a xor b);
    layer6_outputs(9881) <= a xor b;
    layer6_outputs(9882) <= a and not b;
    layer6_outputs(9883) <= not a or b;
    layer6_outputs(9884) <= not a;
    layer6_outputs(9885) <= a xor b;
    layer6_outputs(9886) <= a and not b;
    layer6_outputs(9887) <= a xor b;
    layer6_outputs(9888) <= not (a and b);
    layer6_outputs(9889) <= not a;
    layer6_outputs(9890) <= not b;
    layer6_outputs(9891) <= not b;
    layer6_outputs(9892) <= b;
    layer6_outputs(9893) <= not (a or b);
    layer6_outputs(9894) <= a or b;
    layer6_outputs(9895) <= not b;
    layer6_outputs(9896) <= a and not b;
    layer6_outputs(9897) <= a and not b;
    layer6_outputs(9898) <= b;
    layer6_outputs(9899) <= b;
    layer6_outputs(9900) <= a and b;
    layer6_outputs(9901) <= b;
    layer6_outputs(9902) <= not a;
    layer6_outputs(9903) <= b;
    layer6_outputs(9904) <= a and not b;
    layer6_outputs(9905) <= not b or a;
    layer6_outputs(9906) <= a and b;
    layer6_outputs(9907) <= a or b;
    layer6_outputs(9908) <= a and not b;
    layer6_outputs(9909) <= b;
    layer6_outputs(9910) <= not (a xor b);
    layer6_outputs(9911) <= not a;
    layer6_outputs(9912) <= not a or b;
    layer6_outputs(9913) <= not a;
    layer6_outputs(9914) <= not a;
    layer6_outputs(9915) <= not (a or b);
    layer6_outputs(9916) <= a xor b;
    layer6_outputs(9917) <= a xor b;
    layer6_outputs(9918) <= a xor b;
    layer6_outputs(9919) <= a;
    layer6_outputs(9920) <= not b;
    layer6_outputs(9921) <= a xor b;
    layer6_outputs(9922) <= b and not a;
    layer6_outputs(9923) <= not (a or b);
    layer6_outputs(9924) <= a xor b;
    layer6_outputs(9925) <= a;
    layer6_outputs(9926) <= a xor b;
    layer6_outputs(9927) <= not a;
    layer6_outputs(9928) <= a and b;
    layer6_outputs(9929) <= not (a xor b);
    layer6_outputs(9930) <= a;
    layer6_outputs(9931) <= not b;
    layer6_outputs(9932) <= b;
    layer6_outputs(9933) <= a and b;
    layer6_outputs(9934) <= a xor b;
    layer6_outputs(9935) <= not b or a;
    layer6_outputs(9936) <= b;
    layer6_outputs(9937) <= not b;
    layer6_outputs(9938) <= a;
    layer6_outputs(9939) <= a xor b;
    layer6_outputs(9940) <= b;
    layer6_outputs(9941) <= not b;
    layer6_outputs(9942) <= a;
    layer6_outputs(9943) <= not b or a;
    layer6_outputs(9944) <= not a or b;
    layer6_outputs(9945) <= b;
    layer6_outputs(9946) <= a or b;
    layer6_outputs(9947) <= b;
    layer6_outputs(9948) <= b and not a;
    layer6_outputs(9949) <= a xor b;
    layer6_outputs(9950) <= not (a and b);
    layer6_outputs(9951) <= b and not a;
    layer6_outputs(9952) <= not (a and b);
    layer6_outputs(9953) <= a or b;
    layer6_outputs(9954) <= a and not b;
    layer6_outputs(9955) <= not (a xor b);
    layer6_outputs(9956) <= not a;
    layer6_outputs(9957) <= a xor b;
    layer6_outputs(9958) <= b and not a;
    layer6_outputs(9959) <= not b;
    layer6_outputs(9960) <= not (a xor b);
    layer6_outputs(9961) <= a;
    layer6_outputs(9962) <= a xor b;
    layer6_outputs(9963) <= not a;
    layer6_outputs(9964) <= not b;
    layer6_outputs(9965) <= a or b;
    layer6_outputs(9966) <= not b;
    layer6_outputs(9967) <= b and not a;
    layer6_outputs(9968) <= not a;
    layer6_outputs(9969) <= b;
    layer6_outputs(9970) <= not (a or b);
    layer6_outputs(9971) <= b and not a;
    layer6_outputs(9972) <= not (a xor b);
    layer6_outputs(9973) <= not (a or b);
    layer6_outputs(9974) <= not (a xor b);
    layer6_outputs(9975) <= a xor b;
    layer6_outputs(9976) <= a and not b;
    layer6_outputs(9977) <= a xor b;
    layer6_outputs(9978) <= b and not a;
    layer6_outputs(9979) <= b;
    layer6_outputs(9980) <= not (a xor b);
    layer6_outputs(9981) <= a;
    layer6_outputs(9982) <= a xor b;
    layer6_outputs(9983) <= b and not a;
    layer6_outputs(9984) <= b and not a;
    layer6_outputs(9985) <= b;
    layer6_outputs(9986) <= a xor b;
    layer6_outputs(9987) <= not (a or b);
    layer6_outputs(9988) <= not b or a;
    layer6_outputs(9989) <= b;
    layer6_outputs(9990) <= b;
    layer6_outputs(9991) <= b;
    layer6_outputs(9992) <= not b;
    layer6_outputs(9993) <= not (a or b);
    layer6_outputs(9994) <= a xor b;
    layer6_outputs(9995) <= not (a xor b);
    layer6_outputs(9996) <= not (a xor b);
    layer6_outputs(9997) <= not a;
    layer6_outputs(9998) <= b and not a;
    layer6_outputs(9999) <= not a;
    layer6_outputs(10000) <= not a or b;
    layer6_outputs(10001) <= a xor b;
    layer6_outputs(10002) <= not (a and b);
    layer6_outputs(10003) <= not (a and b);
    layer6_outputs(10004) <= not (a and b);
    layer6_outputs(10005) <= not (a xor b);
    layer6_outputs(10006) <= a xor b;
    layer6_outputs(10007) <= a xor b;
    layer6_outputs(10008) <= not a;
    layer6_outputs(10009) <= not (a or b);
    layer6_outputs(10010) <= not (a and b);
    layer6_outputs(10011) <= b;
    layer6_outputs(10012) <= a xor b;
    layer6_outputs(10013) <= a and not b;
    layer6_outputs(10014) <= not a;
    layer6_outputs(10015) <= '0';
    layer6_outputs(10016) <= a and not b;
    layer6_outputs(10017) <= a xor b;
    layer6_outputs(10018) <= a xor b;
    layer6_outputs(10019) <= a xor b;
    layer6_outputs(10020) <= not (a or b);
    layer6_outputs(10021) <= b;
    layer6_outputs(10022) <= a;
    layer6_outputs(10023) <= a;
    layer6_outputs(10024) <= not a;
    layer6_outputs(10025) <= not b;
    layer6_outputs(10026) <= not (a xor b);
    layer6_outputs(10027) <= not a;
    layer6_outputs(10028) <= not a;
    layer6_outputs(10029) <= a and b;
    layer6_outputs(10030) <= not a or b;
    layer6_outputs(10031) <= not a;
    layer6_outputs(10032) <= a and not b;
    layer6_outputs(10033) <= not a;
    layer6_outputs(10034) <= not b;
    layer6_outputs(10035) <= not b;
    layer6_outputs(10036) <= a xor b;
    layer6_outputs(10037) <= not b or a;
    layer6_outputs(10038) <= not a or b;
    layer6_outputs(10039) <= not (a xor b);
    layer6_outputs(10040) <= not (a or b);
    layer6_outputs(10041) <= a xor b;
    layer6_outputs(10042) <= b;
    layer6_outputs(10043) <= a xor b;
    layer6_outputs(10044) <= a;
    layer6_outputs(10045) <= not (a and b);
    layer6_outputs(10046) <= not b or a;
    layer6_outputs(10047) <= not b or a;
    layer6_outputs(10048) <= b;
    layer6_outputs(10049) <= not (a xor b);
    layer6_outputs(10050) <= not a or b;
    layer6_outputs(10051) <= b;
    layer6_outputs(10052) <= not b or a;
    layer6_outputs(10053) <= not a;
    layer6_outputs(10054) <= not b or a;
    layer6_outputs(10055) <= a and b;
    layer6_outputs(10056) <= a;
    layer6_outputs(10057) <= b;
    layer6_outputs(10058) <= not a;
    layer6_outputs(10059) <= not (a and b);
    layer6_outputs(10060) <= '1';
    layer6_outputs(10061) <= not (a or b);
    layer6_outputs(10062) <= not (a and b);
    layer6_outputs(10063) <= a and b;
    layer6_outputs(10064) <= a xor b;
    layer6_outputs(10065) <= not (a xor b);
    layer6_outputs(10066) <= not (a xor b);
    layer6_outputs(10067) <= a;
    layer6_outputs(10068) <= b and not a;
    layer6_outputs(10069) <= a xor b;
    layer6_outputs(10070) <= not b;
    layer6_outputs(10071) <= a and not b;
    layer6_outputs(10072) <= not b;
    layer6_outputs(10073) <= a xor b;
    layer6_outputs(10074) <= not (a and b);
    layer6_outputs(10075) <= not a;
    layer6_outputs(10076) <= not (a xor b);
    layer6_outputs(10077) <= not (a and b);
    layer6_outputs(10078) <= not a or b;
    layer6_outputs(10079) <= b;
    layer6_outputs(10080) <= not (a or b);
    layer6_outputs(10081) <= not (a and b);
    layer6_outputs(10082) <= not a or b;
    layer6_outputs(10083) <= a;
    layer6_outputs(10084) <= a and not b;
    layer6_outputs(10085) <= a or b;
    layer6_outputs(10086) <= not (a and b);
    layer6_outputs(10087) <= a and b;
    layer6_outputs(10088) <= not (a xor b);
    layer6_outputs(10089) <= a xor b;
    layer6_outputs(10090) <= b;
    layer6_outputs(10091) <= not a;
    layer6_outputs(10092) <= not (a xor b);
    layer6_outputs(10093) <= not b or a;
    layer6_outputs(10094) <= b;
    layer6_outputs(10095) <= a and not b;
    layer6_outputs(10096) <= b;
    layer6_outputs(10097) <= a xor b;
    layer6_outputs(10098) <= a and b;
    layer6_outputs(10099) <= not b;
    layer6_outputs(10100) <= a and b;
    layer6_outputs(10101) <= b;
    layer6_outputs(10102) <= a xor b;
    layer6_outputs(10103) <= not a or b;
    layer6_outputs(10104) <= a;
    layer6_outputs(10105) <= a and b;
    layer6_outputs(10106) <= a;
    layer6_outputs(10107) <= not a;
    layer6_outputs(10108) <= not b;
    layer6_outputs(10109) <= not a;
    layer6_outputs(10110) <= not b;
    layer6_outputs(10111) <= not a or b;
    layer6_outputs(10112) <= b and not a;
    layer6_outputs(10113) <= not b or a;
    layer6_outputs(10114) <= not b;
    layer6_outputs(10115) <= not a or b;
    layer6_outputs(10116) <= a and b;
    layer6_outputs(10117) <= not (a xor b);
    layer6_outputs(10118) <= not (a or b);
    layer6_outputs(10119) <= not b;
    layer6_outputs(10120) <= '0';
    layer6_outputs(10121) <= not b or a;
    layer6_outputs(10122) <= not a or b;
    layer6_outputs(10123) <= a and not b;
    layer6_outputs(10124) <= a and not b;
    layer6_outputs(10125) <= a xor b;
    layer6_outputs(10126) <= a and b;
    layer6_outputs(10127) <= not (a xor b);
    layer6_outputs(10128) <= not a or b;
    layer6_outputs(10129) <= a;
    layer6_outputs(10130) <= not a;
    layer6_outputs(10131) <= not b;
    layer6_outputs(10132) <= not (a xor b);
    layer6_outputs(10133) <= a;
    layer6_outputs(10134) <= b and not a;
    layer6_outputs(10135) <= not (a xor b);
    layer6_outputs(10136) <= not (a xor b);
    layer6_outputs(10137) <= a xor b;
    layer6_outputs(10138) <= not a;
    layer6_outputs(10139) <= a;
    layer6_outputs(10140) <= not b;
    layer6_outputs(10141) <= not b;
    layer6_outputs(10142) <= a;
    layer6_outputs(10143) <= not a or b;
    layer6_outputs(10144) <= a xor b;
    layer6_outputs(10145) <= b and not a;
    layer6_outputs(10146) <= not a or b;
    layer6_outputs(10147) <= not b;
    layer6_outputs(10148) <= a xor b;
    layer6_outputs(10149) <= not b or a;
    layer6_outputs(10150) <= not (a xor b);
    layer6_outputs(10151) <= a xor b;
    layer6_outputs(10152) <= a xor b;
    layer6_outputs(10153) <= not a;
    layer6_outputs(10154) <= not a;
    layer6_outputs(10155) <= not a;
    layer6_outputs(10156) <= not b;
    layer6_outputs(10157) <= a or b;
    layer6_outputs(10158) <= not a;
    layer6_outputs(10159) <= not a;
    layer6_outputs(10160) <= a;
    layer6_outputs(10161) <= not (a xor b);
    layer6_outputs(10162) <= not a;
    layer6_outputs(10163) <= b;
    layer6_outputs(10164) <= not (a xor b);
    layer6_outputs(10165) <= not b;
    layer6_outputs(10166) <= not (a or b);
    layer6_outputs(10167) <= a;
    layer6_outputs(10168) <= not a;
    layer6_outputs(10169) <= a;
    layer6_outputs(10170) <= not (a xor b);
    layer6_outputs(10171) <= a or b;
    layer6_outputs(10172) <= b;
    layer6_outputs(10173) <= not b;
    layer6_outputs(10174) <= a xor b;
    layer6_outputs(10175) <= a and not b;
    layer6_outputs(10176) <= not a;
    layer6_outputs(10177) <= a;
    layer6_outputs(10178) <= a;
    layer6_outputs(10179) <= not (a xor b);
    layer6_outputs(10180) <= a xor b;
    layer6_outputs(10181) <= b and not a;
    layer6_outputs(10182) <= a xor b;
    layer6_outputs(10183) <= not b;
    layer6_outputs(10184) <= not b;
    layer6_outputs(10185) <= not a;
    layer6_outputs(10186) <= b and not a;
    layer6_outputs(10187) <= b and not a;
    layer6_outputs(10188) <= a;
    layer6_outputs(10189) <= a;
    layer6_outputs(10190) <= b and not a;
    layer6_outputs(10191) <= b;
    layer6_outputs(10192) <= not a or b;
    layer6_outputs(10193) <= not b;
    layer6_outputs(10194) <= not a or b;
    layer6_outputs(10195) <= a;
    layer6_outputs(10196) <= b;
    layer6_outputs(10197) <= b;
    layer6_outputs(10198) <= a;
    layer6_outputs(10199) <= not (a and b);
    layer6_outputs(10200) <= a xor b;
    layer6_outputs(10201) <= b;
    layer6_outputs(10202) <= b and not a;
    layer6_outputs(10203) <= not a;
    layer6_outputs(10204) <= a;
    layer6_outputs(10205) <= not a;
    layer6_outputs(10206) <= not b or a;
    layer6_outputs(10207) <= b;
    layer6_outputs(10208) <= not b;
    layer6_outputs(10209) <= b;
    layer6_outputs(10210) <= b;
    layer6_outputs(10211) <= not a;
    layer6_outputs(10212) <= not a or b;
    layer6_outputs(10213) <= '1';
    layer6_outputs(10214) <= not (a xor b);
    layer6_outputs(10215) <= not (a xor b);
    layer6_outputs(10216) <= b;
    layer6_outputs(10217) <= not a;
    layer6_outputs(10218) <= not (a xor b);
    layer6_outputs(10219) <= not a or b;
    layer6_outputs(10220) <= b;
    layer6_outputs(10221) <= a or b;
    layer6_outputs(10222) <= not a or b;
    layer6_outputs(10223) <= a;
    layer6_outputs(10224) <= not b;
    layer6_outputs(10225) <= not a;
    layer6_outputs(10226) <= a or b;
    layer6_outputs(10227) <= not a;
    layer6_outputs(10228) <= b;
    layer6_outputs(10229) <= not a;
    layer6_outputs(10230) <= a xor b;
    layer6_outputs(10231) <= a xor b;
    layer6_outputs(10232) <= not (a or b);
    layer6_outputs(10233) <= not (a and b);
    layer6_outputs(10234) <= b;
    layer6_outputs(10235) <= a;
    layer6_outputs(10236) <= a and not b;
    layer6_outputs(10237) <= not b;
    layer6_outputs(10238) <= not (a xor b);
    layer6_outputs(10239) <= a xor b;
    layer6_outputs(10240) <= a;
    layer6_outputs(10241) <= a;
    layer6_outputs(10242) <= not (a or b);
    layer6_outputs(10243) <= a and b;
    layer6_outputs(10244) <= not a;
    layer6_outputs(10245) <= not (a and b);
    layer6_outputs(10246) <= not b;
    layer6_outputs(10247) <= not b;
    layer6_outputs(10248) <= a;
    layer6_outputs(10249) <= b and not a;
    layer6_outputs(10250) <= a and b;
    layer6_outputs(10251) <= a;
    layer6_outputs(10252) <= a and not b;
    layer6_outputs(10253) <= b and not a;
    layer6_outputs(10254) <= a xor b;
    layer6_outputs(10255) <= '1';
    layer6_outputs(10256) <= a;
    layer6_outputs(10257) <= a;
    layer6_outputs(10258) <= a;
    layer6_outputs(10259) <= a and not b;
    layer6_outputs(10260) <= not (a xor b);
    layer6_outputs(10261) <= '1';
    layer6_outputs(10262) <= a xor b;
    layer6_outputs(10263) <= not b;
    layer6_outputs(10264) <= a;
    layer6_outputs(10265) <= a or b;
    layer6_outputs(10266) <= b and not a;
    layer6_outputs(10267) <= b;
    layer6_outputs(10268) <= b and not a;
    layer6_outputs(10269) <= a xor b;
    layer6_outputs(10270) <= not a or b;
    layer6_outputs(10271) <= not b;
    layer6_outputs(10272) <= b;
    layer6_outputs(10273) <= not (a xor b);
    layer6_outputs(10274) <= b;
    layer6_outputs(10275) <= not b or a;
    layer6_outputs(10276) <= not b;
    layer6_outputs(10277) <= not b;
    layer6_outputs(10278) <= a xor b;
    layer6_outputs(10279) <= a;
    layer6_outputs(10280) <= a or b;
    layer6_outputs(10281) <= not (a xor b);
    layer6_outputs(10282) <= a;
    layer6_outputs(10283) <= b;
    layer6_outputs(10284) <= not (a xor b);
    layer6_outputs(10285) <= a xor b;
    layer6_outputs(10286) <= not a;
    layer6_outputs(10287) <= a;
    layer6_outputs(10288) <= not a;
    layer6_outputs(10289) <= not a;
    layer6_outputs(10290) <= not (a xor b);
    layer6_outputs(10291) <= not (a xor b);
    layer6_outputs(10292) <= a and not b;
    layer6_outputs(10293) <= not b or a;
    layer6_outputs(10294) <= not a;
    layer6_outputs(10295) <= a;
    layer6_outputs(10296) <= a xor b;
    layer6_outputs(10297) <= a;
    layer6_outputs(10298) <= b;
    layer6_outputs(10299) <= b and not a;
    layer6_outputs(10300) <= a and b;
    layer6_outputs(10301) <= a;
    layer6_outputs(10302) <= a;
    layer6_outputs(10303) <= not (a xor b);
    layer6_outputs(10304) <= not a or b;
    layer6_outputs(10305) <= a and not b;
    layer6_outputs(10306) <= a xor b;
    layer6_outputs(10307) <= not (a and b);
    layer6_outputs(10308) <= a;
    layer6_outputs(10309) <= not (a xor b);
    layer6_outputs(10310) <= a and not b;
    layer6_outputs(10311) <= a xor b;
    layer6_outputs(10312) <= a xor b;
    layer6_outputs(10313) <= a and b;
    layer6_outputs(10314) <= a and not b;
    layer6_outputs(10315) <= not (a xor b);
    layer6_outputs(10316) <= not (a or b);
    layer6_outputs(10317) <= a xor b;
    layer6_outputs(10318) <= not a;
    layer6_outputs(10319) <= a;
    layer6_outputs(10320) <= b;
    layer6_outputs(10321) <= not (a xor b);
    layer6_outputs(10322) <= a and not b;
    layer6_outputs(10323) <= not b or a;
    layer6_outputs(10324) <= a and not b;
    layer6_outputs(10325) <= b;
    layer6_outputs(10326) <= not b;
    layer6_outputs(10327) <= a xor b;
    layer6_outputs(10328) <= not (a xor b);
    layer6_outputs(10329) <= a or b;
    layer6_outputs(10330) <= a and not b;
    layer6_outputs(10331) <= not b;
    layer6_outputs(10332) <= b;
    layer6_outputs(10333) <= not a;
    layer6_outputs(10334) <= b;
    layer6_outputs(10335) <= a or b;
    layer6_outputs(10336) <= not (a xor b);
    layer6_outputs(10337) <= b;
    layer6_outputs(10338) <= not (a xor b);
    layer6_outputs(10339) <= not (a xor b);
    layer6_outputs(10340) <= not b or a;
    layer6_outputs(10341) <= not (a and b);
    layer6_outputs(10342) <= a;
    layer6_outputs(10343) <= not a or b;
    layer6_outputs(10344) <= a or b;
    layer6_outputs(10345) <= b;
    layer6_outputs(10346) <= a xor b;
    layer6_outputs(10347) <= b;
    layer6_outputs(10348) <= not b;
    layer6_outputs(10349) <= a xor b;
    layer6_outputs(10350) <= not b;
    layer6_outputs(10351) <= not b or a;
    layer6_outputs(10352) <= a;
    layer6_outputs(10353) <= not (a xor b);
    layer6_outputs(10354) <= b;
    layer6_outputs(10355) <= not (a or b);
    layer6_outputs(10356) <= b;
    layer6_outputs(10357) <= not (a or b);
    layer6_outputs(10358) <= not a;
    layer6_outputs(10359) <= not a;
    layer6_outputs(10360) <= not (a xor b);
    layer6_outputs(10361) <= a;
    layer6_outputs(10362) <= a or b;
    layer6_outputs(10363) <= a or b;
    layer6_outputs(10364) <= not a;
    layer6_outputs(10365) <= b;
    layer6_outputs(10366) <= b and not a;
    layer6_outputs(10367) <= not b;
    layer6_outputs(10368) <= not b;
    layer6_outputs(10369) <= a xor b;
    layer6_outputs(10370) <= a;
    layer6_outputs(10371) <= not (a or b);
    layer6_outputs(10372) <= not (a xor b);
    layer6_outputs(10373) <= a and not b;
    layer6_outputs(10374) <= a and not b;
    layer6_outputs(10375) <= b;
    layer6_outputs(10376) <= a;
    layer6_outputs(10377) <= not (a xor b);
    layer6_outputs(10378) <= a;
    layer6_outputs(10379) <= a;
    layer6_outputs(10380) <= not (a xor b);
    layer6_outputs(10381) <= not a or b;
    layer6_outputs(10382) <= not a;
    layer6_outputs(10383) <= not a or b;
    layer6_outputs(10384) <= not b;
    layer6_outputs(10385) <= a;
    layer6_outputs(10386) <= not (a xor b);
    layer6_outputs(10387) <= not a;
    layer6_outputs(10388) <= a xor b;
    layer6_outputs(10389) <= a xor b;
    layer6_outputs(10390) <= a;
    layer6_outputs(10391) <= a xor b;
    layer6_outputs(10392) <= a;
    layer6_outputs(10393) <= a xor b;
    layer6_outputs(10394) <= a;
    layer6_outputs(10395) <= not (a xor b);
    layer6_outputs(10396) <= b;
    layer6_outputs(10397) <= not (a xor b);
    layer6_outputs(10398) <= not b or a;
    layer6_outputs(10399) <= a;
    layer6_outputs(10400) <= not (a and b);
    layer6_outputs(10401) <= not (a xor b);
    layer6_outputs(10402) <= a;
    layer6_outputs(10403) <= a and b;
    layer6_outputs(10404) <= not (a xor b);
    layer6_outputs(10405) <= b and not a;
    layer6_outputs(10406) <= not b;
    layer6_outputs(10407) <= not (a and b);
    layer6_outputs(10408) <= a;
    layer6_outputs(10409) <= b;
    layer6_outputs(10410) <= a;
    layer6_outputs(10411) <= a xor b;
    layer6_outputs(10412) <= a or b;
    layer6_outputs(10413) <= not b;
    layer6_outputs(10414) <= b;
    layer6_outputs(10415) <= not (a xor b);
    layer6_outputs(10416) <= a;
    layer6_outputs(10417) <= not a;
    layer6_outputs(10418) <= not (a xor b);
    layer6_outputs(10419) <= not b or a;
    layer6_outputs(10420) <= not a;
    layer6_outputs(10421) <= not a;
    layer6_outputs(10422) <= not a or b;
    layer6_outputs(10423) <= a or b;
    layer6_outputs(10424) <= a xor b;
    layer6_outputs(10425) <= not a;
    layer6_outputs(10426) <= a and b;
    layer6_outputs(10427) <= not (a xor b);
    layer6_outputs(10428) <= not b;
    layer6_outputs(10429) <= not a;
    layer6_outputs(10430) <= b;
    layer6_outputs(10431) <= not b;
    layer6_outputs(10432) <= b and not a;
    layer6_outputs(10433) <= a;
    layer6_outputs(10434) <= not b;
    layer6_outputs(10435) <= '1';
    layer6_outputs(10436) <= not (a xor b);
    layer6_outputs(10437) <= not a or b;
    layer6_outputs(10438) <= not (a and b);
    layer6_outputs(10439) <= a and b;
    layer6_outputs(10440) <= not (a xor b);
    layer6_outputs(10441) <= a and not b;
    layer6_outputs(10442) <= a or b;
    layer6_outputs(10443) <= not b or a;
    layer6_outputs(10444) <= not b or a;
    layer6_outputs(10445) <= not b or a;
    layer6_outputs(10446) <= a;
    layer6_outputs(10447) <= a;
    layer6_outputs(10448) <= not (a xor b);
    layer6_outputs(10449) <= a and not b;
    layer6_outputs(10450) <= not a;
    layer6_outputs(10451) <= b;
    layer6_outputs(10452) <= not b or a;
    layer6_outputs(10453) <= b;
    layer6_outputs(10454) <= not b;
    layer6_outputs(10455) <= not (a or b);
    layer6_outputs(10456) <= a;
    layer6_outputs(10457) <= b;
    layer6_outputs(10458) <= a xor b;
    layer6_outputs(10459) <= not b;
    layer6_outputs(10460) <= not a;
    layer6_outputs(10461) <= not a;
    layer6_outputs(10462) <= b;
    layer6_outputs(10463) <= a xor b;
    layer6_outputs(10464) <= a;
    layer6_outputs(10465) <= a xor b;
    layer6_outputs(10466) <= not b;
    layer6_outputs(10467) <= a and not b;
    layer6_outputs(10468) <= a xor b;
    layer6_outputs(10469) <= not (a xor b);
    layer6_outputs(10470) <= not a;
    layer6_outputs(10471) <= not a;
    layer6_outputs(10472) <= not a;
    layer6_outputs(10473) <= not b;
    layer6_outputs(10474) <= not (a and b);
    layer6_outputs(10475) <= not a or b;
    layer6_outputs(10476) <= b;
    layer6_outputs(10477) <= not (a xor b);
    layer6_outputs(10478) <= a and not b;
    layer6_outputs(10479) <= a xor b;
    layer6_outputs(10480) <= a;
    layer6_outputs(10481) <= b;
    layer6_outputs(10482) <= b;
    layer6_outputs(10483) <= a or b;
    layer6_outputs(10484) <= not a;
    layer6_outputs(10485) <= not b;
    layer6_outputs(10486) <= not a;
    layer6_outputs(10487) <= not a or b;
    layer6_outputs(10488) <= not a;
    layer6_outputs(10489) <= a and b;
    layer6_outputs(10490) <= not b;
    layer6_outputs(10491) <= not a or b;
    layer6_outputs(10492) <= not (a xor b);
    layer6_outputs(10493) <= not b;
    layer6_outputs(10494) <= '1';
    layer6_outputs(10495) <= not (a or b);
    layer6_outputs(10496) <= not (a or b);
    layer6_outputs(10497) <= not (a or b);
    layer6_outputs(10498) <= not (a xor b);
    layer6_outputs(10499) <= not b;
    layer6_outputs(10500) <= not b or a;
    layer6_outputs(10501) <= not b;
    layer6_outputs(10502) <= not b;
    layer6_outputs(10503) <= a and not b;
    layer6_outputs(10504) <= a;
    layer6_outputs(10505) <= not b;
    layer6_outputs(10506) <= not a or b;
    layer6_outputs(10507) <= not a;
    layer6_outputs(10508) <= not b or a;
    layer6_outputs(10509) <= not b;
    layer6_outputs(10510) <= not b;
    layer6_outputs(10511) <= not (a xor b);
    layer6_outputs(10512) <= b;
    layer6_outputs(10513) <= a or b;
    layer6_outputs(10514) <= b and not a;
    layer6_outputs(10515) <= b;
    layer6_outputs(10516) <= a xor b;
    layer6_outputs(10517) <= a;
    layer6_outputs(10518) <= not b;
    layer6_outputs(10519) <= not (a or b);
    layer6_outputs(10520) <= a xor b;
    layer6_outputs(10521) <= not (a or b);
    layer6_outputs(10522) <= not (a xor b);
    layer6_outputs(10523) <= b;
    layer6_outputs(10524) <= not b;
    layer6_outputs(10525) <= not a;
    layer6_outputs(10526) <= a and not b;
    layer6_outputs(10527) <= b;
    layer6_outputs(10528) <= not a;
    layer6_outputs(10529) <= b;
    layer6_outputs(10530) <= a;
    layer6_outputs(10531) <= not a or b;
    layer6_outputs(10532) <= not (a xor b);
    layer6_outputs(10533) <= a and not b;
    layer6_outputs(10534) <= a or b;
    layer6_outputs(10535) <= a xor b;
    layer6_outputs(10536) <= not (a xor b);
    layer6_outputs(10537) <= b and not a;
    layer6_outputs(10538) <= not (a or b);
    layer6_outputs(10539) <= b;
    layer6_outputs(10540) <= a;
    layer6_outputs(10541) <= b;
    layer6_outputs(10542) <= not (a and b);
    layer6_outputs(10543) <= a xor b;
    layer6_outputs(10544) <= not a;
    layer6_outputs(10545) <= not a or b;
    layer6_outputs(10546) <= not b;
    layer6_outputs(10547) <= a xor b;
    layer6_outputs(10548) <= b;
    layer6_outputs(10549) <= a and b;
    layer6_outputs(10550) <= b;
    layer6_outputs(10551) <= a or b;
    layer6_outputs(10552) <= '0';
    layer6_outputs(10553) <= a xor b;
    layer6_outputs(10554) <= b and not a;
    layer6_outputs(10555) <= b;
    layer6_outputs(10556) <= not a or b;
    layer6_outputs(10557) <= not a;
    layer6_outputs(10558) <= not b or a;
    layer6_outputs(10559) <= not (a and b);
    layer6_outputs(10560) <= not a;
    layer6_outputs(10561) <= b and not a;
    layer6_outputs(10562) <= b and not a;
    layer6_outputs(10563) <= a and b;
    layer6_outputs(10564) <= a and not b;
    layer6_outputs(10565) <= a and b;
    layer6_outputs(10566) <= not (a and b);
    layer6_outputs(10567) <= not b;
    layer6_outputs(10568) <= not a;
    layer6_outputs(10569) <= b;
    layer6_outputs(10570) <= a and not b;
    layer6_outputs(10571) <= not a;
    layer6_outputs(10572) <= not a;
    layer6_outputs(10573) <= not a;
    layer6_outputs(10574) <= not b;
    layer6_outputs(10575) <= a or b;
    layer6_outputs(10576) <= not (a and b);
    layer6_outputs(10577) <= b;
    layer6_outputs(10578) <= not b;
    layer6_outputs(10579) <= not (a xor b);
    layer6_outputs(10580) <= a xor b;
    layer6_outputs(10581) <= not a;
    layer6_outputs(10582) <= not (a or b);
    layer6_outputs(10583) <= not (a or b);
    layer6_outputs(10584) <= a and b;
    layer6_outputs(10585) <= b;
    layer6_outputs(10586) <= a and b;
    layer6_outputs(10587) <= not a;
    layer6_outputs(10588) <= not b or a;
    layer6_outputs(10589) <= a;
    layer6_outputs(10590) <= b;
    layer6_outputs(10591) <= b and not a;
    layer6_outputs(10592) <= not (a xor b);
    layer6_outputs(10593) <= not a or b;
    layer6_outputs(10594) <= b;
    layer6_outputs(10595) <= a or b;
    layer6_outputs(10596) <= a xor b;
    layer6_outputs(10597) <= not b;
    layer6_outputs(10598) <= not a or b;
    layer6_outputs(10599) <= not (a xor b);
    layer6_outputs(10600) <= not a;
    layer6_outputs(10601) <= a and b;
    layer6_outputs(10602) <= not b or a;
    layer6_outputs(10603) <= not a or b;
    layer6_outputs(10604) <= not a;
    layer6_outputs(10605) <= a xor b;
    layer6_outputs(10606) <= not a or b;
    layer6_outputs(10607) <= a;
    layer6_outputs(10608) <= not (a and b);
    layer6_outputs(10609) <= b;
    layer6_outputs(10610) <= not a or b;
    layer6_outputs(10611) <= not b or a;
    layer6_outputs(10612) <= not b;
    layer6_outputs(10613) <= not b;
    layer6_outputs(10614) <= a;
    layer6_outputs(10615) <= a and b;
    layer6_outputs(10616) <= not b;
    layer6_outputs(10617) <= not b or a;
    layer6_outputs(10618) <= not a;
    layer6_outputs(10619) <= a;
    layer6_outputs(10620) <= not a;
    layer6_outputs(10621) <= b and not a;
    layer6_outputs(10622) <= a;
    layer6_outputs(10623) <= not a;
    layer6_outputs(10624) <= not b;
    layer6_outputs(10625) <= not (a or b);
    layer6_outputs(10626) <= not a;
    layer6_outputs(10627) <= a;
    layer6_outputs(10628) <= not a;
    layer6_outputs(10629) <= not b;
    layer6_outputs(10630) <= a xor b;
    layer6_outputs(10631) <= not b;
    layer6_outputs(10632) <= not (a xor b);
    layer6_outputs(10633) <= b;
    layer6_outputs(10634) <= not (a xor b);
    layer6_outputs(10635) <= b;
    layer6_outputs(10636) <= not (a xor b);
    layer6_outputs(10637) <= not a;
    layer6_outputs(10638) <= a;
    layer6_outputs(10639) <= a or b;
    layer6_outputs(10640) <= a;
    layer6_outputs(10641) <= not (a xor b);
    layer6_outputs(10642) <= not (a xor b);
    layer6_outputs(10643) <= not b or a;
    layer6_outputs(10644) <= a;
    layer6_outputs(10645) <= b;
    layer6_outputs(10646) <= not (a xor b);
    layer6_outputs(10647) <= a;
    layer6_outputs(10648) <= a;
    layer6_outputs(10649) <= a and not b;
    layer6_outputs(10650) <= b and not a;
    layer6_outputs(10651) <= not (a xor b);
    layer6_outputs(10652) <= not b;
    layer6_outputs(10653) <= a xor b;
    layer6_outputs(10654) <= b and not a;
    layer6_outputs(10655) <= not a;
    layer6_outputs(10656) <= b and not a;
    layer6_outputs(10657) <= b;
    layer6_outputs(10658) <= a xor b;
    layer6_outputs(10659) <= not b;
    layer6_outputs(10660) <= not a;
    layer6_outputs(10661) <= not a;
    layer6_outputs(10662) <= not b;
    layer6_outputs(10663) <= a and b;
    layer6_outputs(10664) <= not a;
    layer6_outputs(10665) <= a xor b;
    layer6_outputs(10666) <= b;
    layer6_outputs(10667) <= b and not a;
    layer6_outputs(10668) <= a xor b;
    layer6_outputs(10669) <= not a;
    layer6_outputs(10670) <= not a;
    layer6_outputs(10671) <= not b or a;
    layer6_outputs(10672) <= b;
    layer6_outputs(10673) <= not b;
    layer6_outputs(10674) <= not (a xor b);
    layer6_outputs(10675) <= not (a and b);
    layer6_outputs(10676) <= b;
    layer6_outputs(10677) <= '0';
    layer6_outputs(10678) <= b;
    layer6_outputs(10679) <= not b;
    layer6_outputs(10680) <= not a;
    layer6_outputs(10681) <= a xor b;
    layer6_outputs(10682) <= b;
    layer6_outputs(10683) <= not a;
    layer6_outputs(10684) <= a xor b;
    layer6_outputs(10685) <= b;
    layer6_outputs(10686) <= b;
    layer6_outputs(10687) <= a and not b;
    layer6_outputs(10688) <= a and not b;
    layer6_outputs(10689) <= not a;
    layer6_outputs(10690) <= not a;
    layer6_outputs(10691) <= not a;
    layer6_outputs(10692) <= not (a xor b);
    layer6_outputs(10693) <= not (a or b);
    layer6_outputs(10694) <= not b;
    layer6_outputs(10695) <= a xor b;
    layer6_outputs(10696) <= not (a xor b);
    layer6_outputs(10697) <= not a or b;
    layer6_outputs(10698) <= b;
    layer6_outputs(10699) <= a xor b;
    layer6_outputs(10700) <= a xor b;
    layer6_outputs(10701) <= a xor b;
    layer6_outputs(10702) <= a or b;
    layer6_outputs(10703) <= not a or b;
    layer6_outputs(10704) <= not a or b;
    layer6_outputs(10705) <= not a;
    layer6_outputs(10706) <= not (a xor b);
    layer6_outputs(10707) <= not b;
    layer6_outputs(10708) <= not b or a;
    layer6_outputs(10709) <= a and b;
    layer6_outputs(10710) <= not a;
    layer6_outputs(10711) <= a and b;
    layer6_outputs(10712) <= a and not b;
    layer6_outputs(10713) <= a xor b;
    layer6_outputs(10714) <= a xor b;
    layer6_outputs(10715) <= not (a or b);
    layer6_outputs(10716) <= not a;
    layer6_outputs(10717) <= a;
    layer6_outputs(10718) <= b;
    layer6_outputs(10719) <= not (a xor b);
    layer6_outputs(10720) <= a and b;
    layer6_outputs(10721) <= a;
    layer6_outputs(10722) <= not a;
    layer6_outputs(10723) <= a;
    layer6_outputs(10724) <= b;
    layer6_outputs(10725) <= b and not a;
    layer6_outputs(10726) <= not b or a;
    layer6_outputs(10727) <= not b or a;
    layer6_outputs(10728) <= b and not a;
    layer6_outputs(10729) <= a;
    layer6_outputs(10730) <= not b;
    layer6_outputs(10731) <= not (a xor b);
    layer6_outputs(10732) <= a xor b;
    layer6_outputs(10733) <= not a;
    layer6_outputs(10734) <= a xor b;
    layer6_outputs(10735) <= a;
    layer6_outputs(10736) <= not a;
    layer6_outputs(10737) <= b and not a;
    layer6_outputs(10738) <= a xor b;
    layer6_outputs(10739) <= not b or a;
    layer6_outputs(10740) <= b;
    layer6_outputs(10741) <= not b;
    layer6_outputs(10742) <= not b;
    layer6_outputs(10743) <= a xor b;
    layer6_outputs(10744) <= b;
    layer6_outputs(10745) <= not (a and b);
    layer6_outputs(10746) <= b;
    layer6_outputs(10747) <= not a;
    layer6_outputs(10748) <= not a;
    layer6_outputs(10749) <= b;
    layer6_outputs(10750) <= not a or b;
    layer6_outputs(10751) <= b;
    layer6_outputs(10752) <= not (a xor b);
    layer6_outputs(10753) <= a or b;
    layer6_outputs(10754) <= a xor b;
    layer6_outputs(10755) <= not a or b;
    layer6_outputs(10756) <= not (a xor b);
    layer6_outputs(10757) <= not b or a;
    layer6_outputs(10758) <= a;
    layer6_outputs(10759) <= not a;
    layer6_outputs(10760) <= not (a and b);
    layer6_outputs(10761) <= a xor b;
    layer6_outputs(10762) <= not b or a;
    layer6_outputs(10763) <= a xor b;
    layer6_outputs(10764) <= a;
    layer6_outputs(10765) <= not (a and b);
    layer6_outputs(10766) <= a or b;
    layer6_outputs(10767) <= b;
    layer6_outputs(10768) <= a;
    layer6_outputs(10769) <= not (a xor b);
    layer6_outputs(10770) <= not a;
    layer6_outputs(10771) <= not a or b;
    layer6_outputs(10772) <= not a;
    layer6_outputs(10773) <= not b;
    layer6_outputs(10774) <= not b or a;
    layer6_outputs(10775) <= a and b;
    layer6_outputs(10776) <= a and not b;
    layer6_outputs(10777) <= a xor b;
    layer6_outputs(10778) <= a and b;
    layer6_outputs(10779) <= not a or b;
    layer6_outputs(10780) <= not a;
    layer6_outputs(10781) <= b;
    layer6_outputs(10782) <= not b or a;
    layer6_outputs(10783) <= a and not b;
    layer6_outputs(10784) <= a;
    layer6_outputs(10785) <= not (a and b);
    layer6_outputs(10786) <= not b;
    layer6_outputs(10787) <= not a;
    layer6_outputs(10788) <= not (a xor b);
    layer6_outputs(10789) <= not b;
    layer6_outputs(10790) <= a and b;
    layer6_outputs(10791) <= not a;
    layer6_outputs(10792) <= b;
    layer6_outputs(10793) <= not (a or b);
    layer6_outputs(10794) <= not (a xor b);
    layer6_outputs(10795) <= a;
    layer6_outputs(10796) <= a or b;
    layer6_outputs(10797) <= not (a or b);
    layer6_outputs(10798) <= a;
    layer6_outputs(10799) <= not (a or b);
    layer6_outputs(10800) <= not (a or b);
    layer6_outputs(10801) <= not a;
    layer6_outputs(10802) <= not (a xor b);
    layer6_outputs(10803) <= not a;
    layer6_outputs(10804) <= not a;
    layer6_outputs(10805) <= a and not b;
    layer6_outputs(10806) <= a and not b;
    layer6_outputs(10807) <= a and b;
    layer6_outputs(10808) <= b;
    layer6_outputs(10809) <= b;
    layer6_outputs(10810) <= b;
    layer6_outputs(10811) <= b;
    layer6_outputs(10812) <= b;
    layer6_outputs(10813) <= not a or b;
    layer6_outputs(10814) <= a and not b;
    layer6_outputs(10815) <= a xor b;
    layer6_outputs(10816) <= not b;
    layer6_outputs(10817) <= not b;
    layer6_outputs(10818) <= not b or a;
    layer6_outputs(10819) <= a;
    layer6_outputs(10820) <= b;
    layer6_outputs(10821) <= not b or a;
    layer6_outputs(10822) <= a or b;
    layer6_outputs(10823) <= a and not b;
    layer6_outputs(10824) <= b and not a;
    layer6_outputs(10825) <= a xor b;
    layer6_outputs(10826) <= not a or b;
    layer6_outputs(10827) <= not b;
    layer6_outputs(10828) <= not (a xor b);
    layer6_outputs(10829) <= not a;
    layer6_outputs(10830) <= not a;
    layer6_outputs(10831) <= a xor b;
    layer6_outputs(10832) <= b;
    layer6_outputs(10833) <= not a or b;
    layer6_outputs(10834) <= a;
    layer6_outputs(10835) <= not b or a;
    layer6_outputs(10836) <= not b or a;
    layer6_outputs(10837) <= not (a or b);
    layer6_outputs(10838) <= not b;
    layer6_outputs(10839) <= b and not a;
    layer6_outputs(10840) <= b;
    layer6_outputs(10841) <= not b;
    layer6_outputs(10842) <= a;
    layer6_outputs(10843) <= a xor b;
    layer6_outputs(10844) <= a and b;
    layer6_outputs(10845) <= a or b;
    layer6_outputs(10846) <= a;
    layer6_outputs(10847) <= a and b;
    layer6_outputs(10848) <= a and not b;
    layer6_outputs(10849) <= a or b;
    layer6_outputs(10850) <= not a;
    layer6_outputs(10851) <= not a;
    layer6_outputs(10852) <= a and b;
    layer6_outputs(10853) <= not a or b;
    layer6_outputs(10854) <= not b or a;
    layer6_outputs(10855) <= a xor b;
    layer6_outputs(10856) <= not (a xor b);
    layer6_outputs(10857) <= a and not b;
    layer6_outputs(10858) <= not a;
    layer6_outputs(10859) <= not b;
    layer6_outputs(10860) <= b;
    layer6_outputs(10861) <= not a or b;
    layer6_outputs(10862) <= b;
    layer6_outputs(10863) <= b and not a;
    layer6_outputs(10864) <= b;
    layer6_outputs(10865) <= a and not b;
    layer6_outputs(10866) <= not a;
    layer6_outputs(10867) <= not (a xor b);
    layer6_outputs(10868) <= not a;
    layer6_outputs(10869) <= b and not a;
    layer6_outputs(10870) <= a;
    layer6_outputs(10871) <= a;
    layer6_outputs(10872) <= b;
    layer6_outputs(10873) <= not b;
    layer6_outputs(10874) <= not a;
    layer6_outputs(10875) <= not b;
    layer6_outputs(10876) <= a or b;
    layer6_outputs(10877) <= a or b;
    layer6_outputs(10878) <= not (a xor b);
    layer6_outputs(10879) <= a;
    layer6_outputs(10880) <= a xor b;
    layer6_outputs(10881) <= a xor b;
    layer6_outputs(10882) <= not a;
    layer6_outputs(10883) <= not b;
    layer6_outputs(10884) <= a or b;
    layer6_outputs(10885) <= not (a and b);
    layer6_outputs(10886) <= not a;
    layer6_outputs(10887) <= a;
    layer6_outputs(10888) <= a or b;
    layer6_outputs(10889) <= a;
    layer6_outputs(10890) <= b;
    layer6_outputs(10891) <= not (a or b);
    layer6_outputs(10892) <= '0';
    layer6_outputs(10893) <= b;
    layer6_outputs(10894) <= not b;
    layer6_outputs(10895) <= b;
    layer6_outputs(10896) <= not (a or b);
    layer6_outputs(10897) <= a and b;
    layer6_outputs(10898) <= not (a xor b);
    layer6_outputs(10899) <= a xor b;
    layer6_outputs(10900) <= not a;
    layer6_outputs(10901) <= not (a xor b);
    layer6_outputs(10902) <= not (a and b);
    layer6_outputs(10903) <= a and b;
    layer6_outputs(10904) <= not b;
    layer6_outputs(10905) <= not (a and b);
    layer6_outputs(10906) <= not a;
    layer6_outputs(10907) <= not a;
    layer6_outputs(10908) <= a;
    layer6_outputs(10909) <= b;
    layer6_outputs(10910) <= a and not b;
    layer6_outputs(10911) <= not b;
    layer6_outputs(10912) <= not b or a;
    layer6_outputs(10913) <= not b;
    layer6_outputs(10914) <= not b;
    layer6_outputs(10915) <= not (a xor b);
    layer6_outputs(10916) <= a xor b;
    layer6_outputs(10917) <= a and b;
    layer6_outputs(10918) <= a xor b;
    layer6_outputs(10919) <= not b;
    layer6_outputs(10920) <= a;
    layer6_outputs(10921) <= not (a xor b);
    layer6_outputs(10922) <= not a or b;
    layer6_outputs(10923) <= b;
    layer6_outputs(10924) <= b;
    layer6_outputs(10925) <= a;
    layer6_outputs(10926) <= not (a and b);
    layer6_outputs(10927) <= a;
    layer6_outputs(10928) <= b and not a;
    layer6_outputs(10929) <= not (a and b);
    layer6_outputs(10930) <= not (a or b);
    layer6_outputs(10931) <= not (a xor b);
    layer6_outputs(10932) <= a;
    layer6_outputs(10933) <= a;
    layer6_outputs(10934) <= not (a or b);
    layer6_outputs(10935) <= not b or a;
    layer6_outputs(10936) <= a and not b;
    layer6_outputs(10937) <= a and not b;
    layer6_outputs(10938) <= b;
    layer6_outputs(10939) <= a;
    layer6_outputs(10940) <= a xor b;
    layer6_outputs(10941) <= not a or b;
    layer6_outputs(10942) <= a or b;
    layer6_outputs(10943) <= a;
    layer6_outputs(10944) <= a and not b;
    layer6_outputs(10945) <= b;
    layer6_outputs(10946) <= not b;
    layer6_outputs(10947) <= not (a xor b);
    layer6_outputs(10948) <= b and not a;
    layer6_outputs(10949) <= a and b;
    layer6_outputs(10950) <= not b;
    layer6_outputs(10951) <= not (a xor b);
    layer6_outputs(10952) <= b and not a;
    layer6_outputs(10953) <= a or b;
    layer6_outputs(10954) <= b;
    layer6_outputs(10955) <= a;
    layer6_outputs(10956) <= not (a xor b);
    layer6_outputs(10957) <= not b or a;
    layer6_outputs(10958) <= a xor b;
    layer6_outputs(10959) <= not a or b;
    layer6_outputs(10960) <= b;
    layer6_outputs(10961) <= a xor b;
    layer6_outputs(10962) <= not a;
    layer6_outputs(10963) <= not b;
    layer6_outputs(10964) <= not (a xor b);
    layer6_outputs(10965) <= a and not b;
    layer6_outputs(10966) <= not (a or b);
    layer6_outputs(10967) <= not (a xor b);
    layer6_outputs(10968) <= not (a and b);
    layer6_outputs(10969) <= a xor b;
    layer6_outputs(10970) <= a xor b;
    layer6_outputs(10971) <= not (a xor b);
    layer6_outputs(10972) <= not b;
    layer6_outputs(10973) <= a;
    layer6_outputs(10974) <= not (a or b);
    layer6_outputs(10975) <= not b;
    layer6_outputs(10976) <= not a;
    layer6_outputs(10977) <= not b;
    layer6_outputs(10978) <= not a;
    layer6_outputs(10979) <= b;
    layer6_outputs(10980) <= a;
    layer6_outputs(10981) <= b and not a;
    layer6_outputs(10982) <= not (a and b);
    layer6_outputs(10983) <= not (a or b);
    layer6_outputs(10984) <= a;
    layer6_outputs(10985) <= a;
    layer6_outputs(10986) <= b;
    layer6_outputs(10987) <= not b;
    layer6_outputs(10988) <= b;
    layer6_outputs(10989) <= a xor b;
    layer6_outputs(10990) <= b;
    layer6_outputs(10991) <= not (a xor b);
    layer6_outputs(10992) <= a or b;
    layer6_outputs(10993) <= b;
    layer6_outputs(10994) <= a xor b;
    layer6_outputs(10995) <= a;
    layer6_outputs(10996) <= b;
    layer6_outputs(10997) <= not (a xor b);
    layer6_outputs(10998) <= not a;
    layer6_outputs(10999) <= b;
    layer6_outputs(11000) <= a xor b;
    layer6_outputs(11001) <= not a;
    layer6_outputs(11002) <= not (a and b);
    layer6_outputs(11003) <= not (a and b);
    layer6_outputs(11004) <= b;
    layer6_outputs(11005) <= not b;
    layer6_outputs(11006) <= a;
    layer6_outputs(11007) <= a;
    layer6_outputs(11008) <= not a;
    layer6_outputs(11009) <= b;
    layer6_outputs(11010) <= not b;
    layer6_outputs(11011) <= not (a xor b);
    layer6_outputs(11012) <= not b;
    layer6_outputs(11013) <= a and b;
    layer6_outputs(11014) <= not a or b;
    layer6_outputs(11015) <= a and not b;
    layer6_outputs(11016) <= b and not a;
    layer6_outputs(11017) <= b;
    layer6_outputs(11018) <= not (a xor b);
    layer6_outputs(11019) <= not a;
    layer6_outputs(11020) <= not (a and b);
    layer6_outputs(11021) <= '0';
    layer6_outputs(11022) <= a xor b;
    layer6_outputs(11023) <= not (a and b);
    layer6_outputs(11024) <= a and b;
    layer6_outputs(11025) <= not (a or b);
    layer6_outputs(11026) <= a;
    layer6_outputs(11027) <= b;
    layer6_outputs(11028) <= a;
    layer6_outputs(11029) <= not (a xor b);
    layer6_outputs(11030) <= not b;
    layer6_outputs(11031) <= a or b;
    layer6_outputs(11032) <= not a;
    layer6_outputs(11033) <= a;
    layer6_outputs(11034) <= not b;
    layer6_outputs(11035) <= b;
    layer6_outputs(11036) <= b;
    layer6_outputs(11037) <= b and not a;
    layer6_outputs(11038) <= not a;
    layer6_outputs(11039) <= b and not a;
    layer6_outputs(11040) <= a or b;
    layer6_outputs(11041) <= not (a or b);
    layer6_outputs(11042) <= not (a or b);
    layer6_outputs(11043) <= b;
    layer6_outputs(11044) <= a and b;
    layer6_outputs(11045) <= not b;
    layer6_outputs(11046) <= not (a xor b);
    layer6_outputs(11047) <= not b or a;
    layer6_outputs(11048) <= b;
    layer6_outputs(11049) <= not b;
    layer6_outputs(11050) <= a xor b;
    layer6_outputs(11051) <= a xor b;
    layer6_outputs(11052) <= a xor b;
    layer6_outputs(11053) <= not a;
    layer6_outputs(11054) <= not (a or b);
    layer6_outputs(11055) <= not (a and b);
    layer6_outputs(11056) <= a xor b;
    layer6_outputs(11057) <= a;
    layer6_outputs(11058) <= a;
    layer6_outputs(11059) <= not (a xor b);
    layer6_outputs(11060) <= a;
    layer6_outputs(11061) <= a;
    layer6_outputs(11062) <= not (a and b);
    layer6_outputs(11063) <= not b or a;
    layer6_outputs(11064) <= a and not b;
    layer6_outputs(11065) <= not a;
    layer6_outputs(11066) <= a xor b;
    layer6_outputs(11067) <= b and not a;
    layer6_outputs(11068) <= a xor b;
    layer6_outputs(11069) <= not b;
    layer6_outputs(11070) <= not (a xor b);
    layer6_outputs(11071) <= not b or a;
    layer6_outputs(11072) <= not (a xor b);
    layer6_outputs(11073) <= not (a xor b);
    layer6_outputs(11074) <= a xor b;
    layer6_outputs(11075) <= not a;
    layer6_outputs(11076) <= a and not b;
    layer6_outputs(11077) <= not (a and b);
    layer6_outputs(11078) <= b and not a;
    layer6_outputs(11079) <= a;
    layer6_outputs(11080) <= not b;
    layer6_outputs(11081) <= not (a and b);
    layer6_outputs(11082) <= not (a xor b);
    layer6_outputs(11083) <= not (a and b);
    layer6_outputs(11084) <= a;
    layer6_outputs(11085) <= b;
    layer6_outputs(11086) <= not a or b;
    layer6_outputs(11087) <= not a;
    layer6_outputs(11088) <= a xor b;
    layer6_outputs(11089) <= not a;
    layer6_outputs(11090) <= not (a xor b);
    layer6_outputs(11091) <= a xor b;
    layer6_outputs(11092) <= not (a xor b);
    layer6_outputs(11093) <= a xor b;
    layer6_outputs(11094) <= a xor b;
    layer6_outputs(11095) <= not (a xor b);
    layer6_outputs(11096) <= a;
    layer6_outputs(11097) <= a xor b;
    layer6_outputs(11098) <= b;
    layer6_outputs(11099) <= a;
    layer6_outputs(11100) <= not b or a;
    layer6_outputs(11101) <= not (a xor b);
    layer6_outputs(11102) <= a;
    layer6_outputs(11103) <= a;
    layer6_outputs(11104) <= not b;
    layer6_outputs(11105) <= not b or a;
    layer6_outputs(11106) <= not (a or b);
    layer6_outputs(11107) <= not b or a;
    layer6_outputs(11108) <= a;
    layer6_outputs(11109) <= not (a and b);
    layer6_outputs(11110) <= not a or b;
    layer6_outputs(11111) <= not (a and b);
    layer6_outputs(11112) <= not b;
    layer6_outputs(11113) <= not b or a;
    layer6_outputs(11114) <= a or b;
    layer6_outputs(11115) <= not (a and b);
    layer6_outputs(11116) <= not b or a;
    layer6_outputs(11117) <= a and b;
    layer6_outputs(11118) <= not (a xor b);
    layer6_outputs(11119) <= not b;
    layer6_outputs(11120) <= not a;
    layer6_outputs(11121) <= not (a and b);
    layer6_outputs(11122) <= not a or b;
    layer6_outputs(11123) <= a;
    layer6_outputs(11124) <= not b or a;
    layer6_outputs(11125) <= not b;
    layer6_outputs(11126) <= not b;
    layer6_outputs(11127) <= not a;
    layer6_outputs(11128) <= b;
    layer6_outputs(11129) <= not (a xor b);
    layer6_outputs(11130) <= not a;
    layer6_outputs(11131) <= a xor b;
    layer6_outputs(11132) <= a xor b;
    layer6_outputs(11133) <= a or b;
    layer6_outputs(11134) <= not b;
    layer6_outputs(11135) <= not b;
    layer6_outputs(11136) <= a or b;
    layer6_outputs(11137) <= b and not a;
    layer6_outputs(11138) <= not b or a;
    layer6_outputs(11139) <= not (a xor b);
    layer6_outputs(11140) <= a and not b;
    layer6_outputs(11141) <= a xor b;
    layer6_outputs(11142) <= not b;
    layer6_outputs(11143) <= b;
    layer6_outputs(11144) <= not (a xor b);
    layer6_outputs(11145) <= not (a xor b);
    layer6_outputs(11146) <= not a;
    layer6_outputs(11147) <= not (a xor b);
    layer6_outputs(11148) <= b;
    layer6_outputs(11149) <= a and b;
    layer6_outputs(11150) <= a and b;
    layer6_outputs(11151) <= b and not a;
    layer6_outputs(11152) <= a;
    layer6_outputs(11153) <= b;
    layer6_outputs(11154) <= a;
    layer6_outputs(11155) <= not a or b;
    layer6_outputs(11156) <= b and not a;
    layer6_outputs(11157) <= not (a or b);
    layer6_outputs(11158) <= not (a or b);
    layer6_outputs(11159) <= a xor b;
    layer6_outputs(11160) <= a xor b;
    layer6_outputs(11161) <= not a;
    layer6_outputs(11162) <= not a or b;
    layer6_outputs(11163) <= a;
    layer6_outputs(11164) <= not (a xor b);
    layer6_outputs(11165) <= not (a xor b);
    layer6_outputs(11166) <= b;
    layer6_outputs(11167) <= not b or a;
    layer6_outputs(11168) <= a;
    layer6_outputs(11169) <= not (a or b);
    layer6_outputs(11170) <= b and not a;
    layer6_outputs(11171) <= not b;
    layer6_outputs(11172) <= not b;
    layer6_outputs(11173) <= a and not b;
    layer6_outputs(11174) <= b;
    layer6_outputs(11175) <= a xor b;
    layer6_outputs(11176) <= a;
    layer6_outputs(11177) <= not a or b;
    layer6_outputs(11178) <= a;
    layer6_outputs(11179) <= not (a and b);
    layer6_outputs(11180) <= not a;
    layer6_outputs(11181) <= not a;
    layer6_outputs(11182) <= not (a xor b);
    layer6_outputs(11183) <= not a or b;
    layer6_outputs(11184) <= not b or a;
    layer6_outputs(11185) <= not (a xor b);
    layer6_outputs(11186) <= not b;
    layer6_outputs(11187) <= not (a or b);
    layer6_outputs(11188) <= not a;
    layer6_outputs(11189) <= b;
    layer6_outputs(11190) <= not a or b;
    layer6_outputs(11191) <= not (a or b);
    layer6_outputs(11192) <= a;
    layer6_outputs(11193) <= a xor b;
    layer6_outputs(11194) <= b and not a;
    layer6_outputs(11195) <= b and not a;
    layer6_outputs(11196) <= a xor b;
    layer6_outputs(11197) <= not (a xor b);
    layer6_outputs(11198) <= a and not b;
    layer6_outputs(11199) <= not b or a;
    layer6_outputs(11200) <= a and not b;
    layer6_outputs(11201) <= a xor b;
    layer6_outputs(11202) <= a xor b;
    layer6_outputs(11203) <= a xor b;
    layer6_outputs(11204) <= not a;
    layer6_outputs(11205) <= not (a xor b);
    layer6_outputs(11206) <= not (a xor b);
    layer6_outputs(11207) <= a and not b;
    layer6_outputs(11208) <= a xor b;
    layer6_outputs(11209) <= not (a and b);
    layer6_outputs(11210) <= a xor b;
    layer6_outputs(11211) <= a;
    layer6_outputs(11212) <= not (a or b);
    layer6_outputs(11213) <= b;
    layer6_outputs(11214) <= a;
    layer6_outputs(11215) <= not a;
    layer6_outputs(11216) <= a;
    layer6_outputs(11217) <= b;
    layer6_outputs(11218) <= not a;
    layer6_outputs(11219) <= not (a xor b);
    layer6_outputs(11220) <= b;
    layer6_outputs(11221) <= not (a xor b);
    layer6_outputs(11222) <= not b;
    layer6_outputs(11223) <= not a;
    layer6_outputs(11224) <= a and b;
    layer6_outputs(11225) <= not a or b;
    layer6_outputs(11226) <= not a or b;
    layer6_outputs(11227) <= not a or b;
    layer6_outputs(11228) <= not (a xor b);
    layer6_outputs(11229) <= not (a xor b);
    layer6_outputs(11230) <= not (a or b);
    layer6_outputs(11231) <= not b;
    layer6_outputs(11232) <= a;
    layer6_outputs(11233) <= b;
    layer6_outputs(11234) <= not a;
    layer6_outputs(11235) <= a;
    layer6_outputs(11236) <= b and not a;
    layer6_outputs(11237) <= a xor b;
    layer6_outputs(11238) <= a and not b;
    layer6_outputs(11239) <= a or b;
    layer6_outputs(11240) <= not a or b;
    layer6_outputs(11241) <= a;
    layer6_outputs(11242) <= not a;
    layer6_outputs(11243) <= not a;
    layer6_outputs(11244) <= not b;
    layer6_outputs(11245) <= b;
    layer6_outputs(11246) <= a and b;
    layer6_outputs(11247) <= not (a xor b);
    layer6_outputs(11248) <= not b;
    layer6_outputs(11249) <= not a;
    layer6_outputs(11250) <= a and not b;
    layer6_outputs(11251) <= a;
    layer6_outputs(11252) <= not (a xor b);
    layer6_outputs(11253) <= a or b;
    layer6_outputs(11254) <= a;
    layer6_outputs(11255) <= not (a xor b);
    layer6_outputs(11256) <= not b;
    layer6_outputs(11257) <= a;
    layer6_outputs(11258) <= b and not a;
    layer6_outputs(11259) <= a xor b;
    layer6_outputs(11260) <= a;
    layer6_outputs(11261) <= a xor b;
    layer6_outputs(11262) <= a and not b;
    layer6_outputs(11263) <= not (a or b);
    layer6_outputs(11264) <= not (a xor b);
    layer6_outputs(11265) <= a and not b;
    layer6_outputs(11266) <= not (a xor b);
    layer6_outputs(11267) <= b;
    layer6_outputs(11268) <= not (a and b);
    layer6_outputs(11269) <= a or b;
    layer6_outputs(11270) <= a xor b;
    layer6_outputs(11271) <= not (a and b);
    layer6_outputs(11272) <= a or b;
    layer6_outputs(11273) <= not a;
    layer6_outputs(11274) <= a;
    layer6_outputs(11275) <= a;
    layer6_outputs(11276) <= b;
    layer6_outputs(11277) <= b and not a;
    layer6_outputs(11278) <= a;
    layer6_outputs(11279) <= b;
    layer6_outputs(11280) <= a;
    layer6_outputs(11281) <= a;
    layer6_outputs(11282) <= not a or b;
    layer6_outputs(11283) <= not a;
    layer6_outputs(11284) <= a;
    layer6_outputs(11285) <= not a or b;
    layer6_outputs(11286) <= not (a xor b);
    layer6_outputs(11287) <= a xor b;
    layer6_outputs(11288) <= not a;
    layer6_outputs(11289) <= a and not b;
    layer6_outputs(11290) <= not a;
    layer6_outputs(11291) <= b and not a;
    layer6_outputs(11292) <= b and not a;
    layer6_outputs(11293) <= a xor b;
    layer6_outputs(11294) <= a and b;
    layer6_outputs(11295) <= a xor b;
    layer6_outputs(11296) <= not a or b;
    layer6_outputs(11297) <= b;
    layer6_outputs(11298) <= not b;
    layer6_outputs(11299) <= a or b;
    layer6_outputs(11300) <= not b or a;
    layer6_outputs(11301) <= not (a xor b);
    layer6_outputs(11302) <= a;
    layer6_outputs(11303) <= not a or b;
    layer6_outputs(11304) <= not b;
    layer6_outputs(11305) <= not (a xor b);
    layer6_outputs(11306) <= not a;
    layer6_outputs(11307) <= b and not a;
    layer6_outputs(11308) <= a xor b;
    layer6_outputs(11309) <= a;
    layer6_outputs(11310) <= a xor b;
    layer6_outputs(11311) <= not b;
    layer6_outputs(11312) <= a xor b;
    layer6_outputs(11313) <= not (a or b);
    layer6_outputs(11314) <= b;
    layer6_outputs(11315) <= a xor b;
    layer6_outputs(11316) <= not a;
    layer6_outputs(11317) <= b;
    layer6_outputs(11318) <= not a;
    layer6_outputs(11319) <= a;
    layer6_outputs(11320) <= b;
    layer6_outputs(11321) <= a and b;
    layer6_outputs(11322) <= not (a xor b);
    layer6_outputs(11323) <= a xor b;
    layer6_outputs(11324) <= a;
    layer6_outputs(11325) <= not b;
    layer6_outputs(11326) <= b;
    layer6_outputs(11327) <= not b or a;
    layer6_outputs(11328) <= not a;
    layer6_outputs(11329) <= not a;
    layer6_outputs(11330) <= a xor b;
    layer6_outputs(11331) <= a xor b;
    layer6_outputs(11332) <= not a or b;
    layer6_outputs(11333) <= not b;
    layer6_outputs(11334) <= not (a and b);
    layer6_outputs(11335) <= not (a xor b);
    layer6_outputs(11336) <= not (a xor b);
    layer6_outputs(11337) <= not b;
    layer6_outputs(11338) <= b;
    layer6_outputs(11339) <= not a;
    layer6_outputs(11340) <= a;
    layer6_outputs(11341) <= b;
    layer6_outputs(11342) <= b and not a;
    layer6_outputs(11343) <= b;
    layer6_outputs(11344) <= not b or a;
    layer6_outputs(11345) <= not b or a;
    layer6_outputs(11346) <= b;
    layer6_outputs(11347) <= a and b;
    layer6_outputs(11348) <= not (a and b);
    layer6_outputs(11349) <= a;
    layer6_outputs(11350) <= not b;
    layer6_outputs(11351) <= a and b;
    layer6_outputs(11352) <= not (a or b);
    layer6_outputs(11353) <= not b or a;
    layer6_outputs(11354) <= a and b;
    layer6_outputs(11355) <= not a;
    layer6_outputs(11356) <= not b or a;
    layer6_outputs(11357) <= not (a or b);
    layer6_outputs(11358) <= not a;
    layer6_outputs(11359) <= a;
    layer6_outputs(11360) <= not b;
    layer6_outputs(11361) <= a;
    layer6_outputs(11362) <= not (a and b);
    layer6_outputs(11363) <= not a;
    layer6_outputs(11364) <= b;
    layer6_outputs(11365) <= not (a xor b);
    layer6_outputs(11366) <= not a or b;
    layer6_outputs(11367) <= not b or a;
    layer6_outputs(11368) <= a xor b;
    layer6_outputs(11369) <= a xor b;
    layer6_outputs(11370) <= a and b;
    layer6_outputs(11371) <= a and b;
    layer6_outputs(11372) <= not b;
    layer6_outputs(11373) <= b and not a;
    layer6_outputs(11374) <= not (a or b);
    layer6_outputs(11375) <= not b;
    layer6_outputs(11376) <= b;
    layer6_outputs(11377) <= b;
    layer6_outputs(11378) <= not (a or b);
    layer6_outputs(11379) <= a and not b;
    layer6_outputs(11380) <= a and not b;
    layer6_outputs(11381) <= not a;
    layer6_outputs(11382) <= not (a xor b);
    layer6_outputs(11383) <= a;
    layer6_outputs(11384) <= not (a xor b);
    layer6_outputs(11385) <= a xor b;
    layer6_outputs(11386) <= not (a or b);
    layer6_outputs(11387) <= a and not b;
    layer6_outputs(11388) <= b and not a;
    layer6_outputs(11389) <= not (a xor b);
    layer6_outputs(11390) <= not b or a;
    layer6_outputs(11391) <= not a;
    layer6_outputs(11392) <= a xor b;
    layer6_outputs(11393) <= a;
    layer6_outputs(11394) <= not b;
    layer6_outputs(11395) <= a xor b;
    layer6_outputs(11396) <= a xor b;
    layer6_outputs(11397) <= not a;
    layer6_outputs(11398) <= a xor b;
    layer6_outputs(11399) <= not a or b;
    layer6_outputs(11400) <= b;
    layer6_outputs(11401) <= a or b;
    layer6_outputs(11402) <= not b;
    layer6_outputs(11403) <= a;
    layer6_outputs(11404) <= a xor b;
    layer6_outputs(11405) <= a;
    layer6_outputs(11406) <= not (a or b);
    layer6_outputs(11407) <= b;
    layer6_outputs(11408) <= a xor b;
    layer6_outputs(11409) <= a xor b;
    layer6_outputs(11410) <= a xor b;
    layer6_outputs(11411) <= not a;
    layer6_outputs(11412) <= a and not b;
    layer6_outputs(11413) <= a;
    layer6_outputs(11414) <= a xor b;
    layer6_outputs(11415) <= not (a and b);
    layer6_outputs(11416) <= a xor b;
    layer6_outputs(11417) <= not a or b;
    layer6_outputs(11418) <= a or b;
    layer6_outputs(11419) <= a or b;
    layer6_outputs(11420) <= not a or b;
    layer6_outputs(11421) <= not b;
    layer6_outputs(11422) <= b;
    layer6_outputs(11423) <= not (a xor b);
    layer6_outputs(11424) <= not (a xor b);
    layer6_outputs(11425) <= not a;
    layer6_outputs(11426) <= not (a xor b);
    layer6_outputs(11427) <= not a or b;
    layer6_outputs(11428) <= not (a xor b);
    layer6_outputs(11429) <= not b;
    layer6_outputs(11430) <= not b;
    layer6_outputs(11431) <= not b or a;
    layer6_outputs(11432) <= not (a xor b);
    layer6_outputs(11433) <= not b;
    layer6_outputs(11434) <= a;
    layer6_outputs(11435) <= not (a and b);
    layer6_outputs(11436) <= not a;
    layer6_outputs(11437) <= a;
    layer6_outputs(11438) <= not (a or b);
    layer6_outputs(11439) <= not a;
    layer6_outputs(11440) <= a or b;
    layer6_outputs(11441) <= '0';
    layer6_outputs(11442) <= b;
    layer6_outputs(11443) <= a xor b;
    layer6_outputs(11444) <= not b;
    layer6_outputs(11445) <= not a or b;
    layer6_outputs(11446) <= not a;
    layer6_outputs(11447) <= not (a and b);
    layer6_outputs(11448) <= not (a xor b);
    layer6_outputs(11449) <= b;
    layer6_outputs(11450) <= not b;
    layer6_outputs(11451) <= a xor b;
    layer6_outputs(11452) <= a and b;
    layer6_outputs(11453) <= b and not a;
    layer6_outputs(11454) <= a;
    layer6_outputs(11455) <= not b or a;
    layer6_outputs(11456) <= a;
    layer6_outputs(11457) <= a xor b;
    layer6_outputs(11458) <= a;
    layer6_outputs(11459) <= not a;
    layer6_outputs(11460) <= not (a or b);
    layer6_outputs(11461) <= not b;
    layer6_outputs(11462) <= a or b;
    layer6_outputs(11463) <= a xor b;
    layer6_outputs(11464) <= not b;
    layer6_outputs(11465) <= a;
    layer6_outputs(11466) <= b;
    layer6_outputs(11467) <= not a;
    layer6_outputs(11468) <= a xor b;
    layer6_outputs(11469) <= b;
    layer6_outputs(11470) <= a and not b;
    layer6_outputs(11471) <= not a;
    layer6_outputs(11472) <= a and b;
    layer6_outputs(11473) <= b;
    layer6_outputs(11474) <= not (a or b);
    layer6_outputs(11475) <= not (a or b);
    layer6_outputs(11476) <= not (a xor b);
    layer6_outputs(11477) <= a xor b;
    layer6_outputs(11478) <= not a;
    layer6_outputs(11479) <= b;
    layer6_outputs(11480) <= not (a xor b);
    layer6_outputs(11481) <= a xor b;
    layer6_outputs(11482) <= not a;
    layer6_outputs(11483) <= '1';
    layer6_outputs(11484) <= not a;
    layer6_outputs(11485) <= a;
    layer6_outputs(11486) <= not a;
    layer6_outputs(11487) <= not b;
    layer6_outputs(11488) <= a or b;
    layer6_outputs(11489) <= not b;
    layer6_outputs(11490) <= a;
    layer6_outputs(11491) <= not (a or b);
    layer6_outputs(11492) <= a or b;
    layer6_outputs(11493) <= not (a or b);
    layer6_outputs(11494) <= not a;
    layer6_outputs(11495) <= not a or b;
    layer6_outputs(11496) <= not a or b;
    layer6_outputs(11497) <= b and not a;
    layer6_outputs(11498) <= not a;
    layer6_outputs(11499) <= b and not a;
    layer6_outputs(11500) <= not b;
    layer6_outputs(11501) <= b;
    layer6_outputs(11502) <= not (a xor b);
    layer6_outputs(11503) <= a xor b;
    layer6_outputs(11504) <= not a;
    layer6_outputs(11505) <= a and not b;
    layer6_outputs(11506) <= not (a or b);
    layer6_outputs(11507) <= not (a and b);
    layer6_outputs(11508) <= a;
    layer6_outputs(11509) <= not (a xor b);
    layer6_outputs(11510) <= not (a xor b);
    layer6_outputs(11511) <= not b or a;
    layer6_outputs(11512) <= a or b;
    layer6_outputs(11513) <= not (a xor b);
    layer6_outputs(11514) <= not b;
    layer6_outputs(11515) <= b;
    layer6_outputs(11516) <= not a or b;
    layer6_outputs(11517) <= not a or b;
    layer6_outputs(11518) <= a xor b;
    layer6_outputs(11519) <= b;
    layer6_outputs(11520) <= not (a or b);
    layer6_outputs(11521) <= not (a xor b);
    layer6_outputs(11522) <= not a or b;
    layer6_outputs(11523) <= a xor b;
    layer6_outputs(11524) <= a and b;
    layer6_outputs(11525) <= a xor b;
    layer6_outputs(11526) <= a and not b;
    layer6_outputs(11527) <= not a;
    layer6_outputs(11528) <= b;
    layer6_outputs(11529) <= not b;
    layer6_outputs(11530) <= a xor b;
    layer6_outputs(11531) <= b;
    layer6_outputs(11532) <= a and not b;
    layer6_outputs(11533) <= not (a xor b);
    layer6_outputs(11534) <= a and b;
    layer6_outputs(11535) <= not b;
    layer6_outputs(11536) <= b;
    layer6_outputs(11537) <= b;
    layer6_outputs(11538) <= b;
    layer6_outputs(11539) <= not (a xor b);
    layer6_outputs(11540) <= not (a xor b);
    layer6_outputs(11541) <= not b;
    layer6_outputs(11542) <= b and not a;
    layer6_outputs(11543) <= b;
    layer6_outputs(11544) <= a;
    layer6_outputs(11545) <= not (a xor b);
    layer6_outputs(11546) <= not (a or b);
    layer6_outputs(11547) <= not b or a;
    layer6_outputs(11548) <= not a;
    layer6_outputs(11549) <= not (a and b);
    layer6_outputs(11550) <= a;
    layer6_outputs(11551) <= not (a xor b);
    layer6_outputs(11552) <= '0';
    layer6_outputs(11553) <= not a;
    layer6_outputs(11554) <= a or b;
    layer6_outputs(11555) <= not b;
    layer6_outputs(11556) <= a;
    layer6_outputs(11557) <= not (a and b);
    layer6_outputs(11558) <= not a;
    layer6_outputs(11559) <= not (a xor b);
    layer6_outputs(11560) <= not b or a;
    layer6_outputs(11561) <= not (a xor b);
    layer6_outputs(11562) <= not a;
    layer6_outputs(11563) <= a and not b;
    layer6_outputs(11564) <= not (a or b);
    layer6_outputs(11565) <= a xor b;
    layer6_outputs(11566) <= a xor b;
    layer6_outputs(11567) <= not a;
    layer6_outputs(11568) <= a;
    layer6_outputs(11569) <= a xor b;
    layer6_outputs(11570) <= not (a or b);
    layer6_outputs(11571) <= a and b;
    layer6_outputs(11572) <= b;
    layer6_outputs(11573) <= a xor b;
    layer6_outputs(11574) <= not b;
    layer6_outputs(11575) <= not (a or b);
    layer6_outputs(11576) <= not (a and b);
    layer6_outputs(11577) <= a and not b;
    layer6_outputs(11578) <= b;
    layer6_outputs(11579) <= not a;
    layer6_outputs(11580) <= not b;
    layer6_outputs(11581) <= a and b;
    layer6_outputs(11582) <= b;
    layer6_outputs(11583) <= a and b;
    layer6_outputs(11584) <= not a;
    layer6_outputs(11585) <= a;
    layer6_outputs(11586) <= not (a xor b);
    layer6_outputs(11587) <= b;
    layer6_outputs(11588) <= a or b;
    layer6_outputs(11589) <= b;
    layer6_outputs(11590) <= not a;
    layer6_outputs(11591) <= b;
    layer6_outputs(11592) <= a xor b;
    layer6_outputs(11593) <= a xor b;
    layer6_outputs(11594) <= a or b;
    layer6_outputs(11595) <= b;
    layer6_outputs(11596) <= a;
    layer6_outputs(11597) <= not a;
    layer6_outputs(11598) <= a or b;
    layer6_outputs(11599) <= b;
    layer6_outputs(11600) <= b and not a;
    layer6_outputs(11601) <= a;
    layer6_outputs(11602) <= not (a and b);
    layer6_outputs(11603) <= not b;
    layer6_outputs(11604) <= a;
    layer6_outputs(11605) <= a;
    layer6_outputs(11606) <= not a;
    layer6_outputs(11607) <= not b;
    layer6_outputs(11608) <= not b;
    layer6_outputs(11609) <= not a;
    layer6_outputs(11610) <= a;
    layer6_outputs(11611) <= not b;
    layer6_outputs(11612) <= b;
    layer6_outputs(11613) <= not a or b;
    layer6_outputs(11614) <= not a or b;
    layer6_outputs(11615) <= b;
    layer6_outputs(11616) <= not (a or b);
    layer6_outputs(11617) <= not (a xor b);
    layer6_outputs(11618) <= b;
    layer6_outputs(11619) <= a;
    layer6_outputs(11620) <= a;
    layer6_outputs(11621) <= not (a and b);
    layer6_outputs(11622) <= b;
    layer6_outputs(11623) <= a xor b;
    layer6_outputs(11624) <= b and not a;
    layer6_outputs(11625) <= b;
    layer6_outputs(11626) <= b;
    layer6_outputs(11627) <= b;
    layer6_outputs(11628) <= a or b;
    layer6_outputs(11629) <= not (a and b);
    layer6_outputs(11630) <= a;
    layer6_outputs(11631) <= b;
    layer6_outputs(11632) <= not a;
    layer6_outputs(11633) <= a xor b;
    layer6_outputs(11634) <= a and not b;
    layer6_outputs(11635) <= not (a xor b);
    layer6_outputs(11636) <= not (a and b);
    layer6_outputs(11637) <= not (a xor b);
    layer6_outputs(11638) <= a;
    layer6_outputs(11639) <= not a or b;
    layer6_outputs(11640) <= not a;
    layer6_outputs(11641) <= not (a xor b);
    layer6_outputs(11642) <= not a or b;
    layer6_outputs(11643) <= not (a or b);
    layer6_outputs(11644) <= b;
    layer6_outputs(11645) <= not b;
    layer6_outputs(11646) <= a;
    layer6_outputs(11647) <= a;
    layer6_outputs(11648) <= a;
    layer6_outputs(11649) <= b;
    layer6_outputs(11650) <= not (a and b);
    layer6_outputs(11651) <= b;
    layer6_outputs(11652) <= not (a or b);
    layer6_outputs(11653) <= a or b;
    layer6_outputs(11654) <= not a;
    layer6_outputs(11655) <= not a;
    layer6_outputs(11656) <= not (a or b);
    layer6_outputs(11657) <= a xor b;
    layer6_outputs(11658) <= not (a or b);
    layer6_outputs(11659) <= not (a xor b);
    layer6_outputs(11660) <= a xor b;
    layer6_outputs(11661) <= not a;
    layer6_outputs(11662) <= not (a or b);
    layer6_outputs(11663) <= not (a or b);
    layer6_outputs(11664) <= a or b;
    layer6_outputs(11665) <= b;
    layer6_outputs(11666) <= not b or a;
    layer6_outputs(11667) <= not a or b;
    layer6_outputs(11668) <= a;
    layer6_outputs(11669) <= not b;
    layer6_outputs(11670) <= a and b;
    layer6_outputs(11671) <= a and not b;
    layer6_outputs(11672) <= a;
    layer6_outputs(11673) <= b;
    layer6_outputs(11674) <= not a;
    layer6_outputs(11675) <= b;
    layer6_outputs(11676) <= a or b;
    layer6_outputs(11677) <= a xor b;
    layer6_outputs(11678) <= b;
    layer6_outputs(11679) <= not b;
    layer6_outputs(11680) <= not b;
    layer6_outputs(11681) <= a xor b;
    layer6_outputs(11682) <= not b or a;
    layer6_outputs(11683) <= not b or a;
    layer6_outputs(11684) <= not b;
    layer6_outputs(11685) <= not (a or b);
    layer6_outputs(11686) <= not (a xor b);
    layer6_outputs(11687) <= not (a or b);
    layer6_outputs(11688) <= a or b;
    layer6_outputs(11689) <= b;
    layer6_outputs(11690) <= not a;
    layer6_outputs(11691) <= a xor b;
    layer6_outputs(11692) <= b;
    layer6_outputs(11693) <= not (a xor b);
    layer6_outputs(11694) <= not b;
    layer6_outputs(11695) <= not a;
    layer6_outputs(11696) <= not (a and b);
    layer6_outputs(11697) <= not a;
    layer6_outputs(11698) <= a or b;
    layer6_outputs(11699) <= not (a or b);
    layer6_outputs(11700) <= not b;
    layer6_outputs(11701) <= not (a or b);
    layer6_outputs(11702) <= a xor b;
    layer6_outputs(11703) <= not (a xor b);
    layer6_outputs(11704) <= not b;
    layer6_outputs(11705) <= a xor b;
    layer6_outputs(11706) <= a and not b;
    layer6_outputs(11707) <= not a;
    layer6_outputs(11708) <= a xor b;
    layer6_outputs(11709) <= a or b;
    layer6_outputs(11710) <= a xor b;
    layer6_outputs(11711) <= a;
    layer6_outputs(11712) <= not a;
    layer6_outputs(11713) <= a xor b;
    layer6_outputs(11714) <= not a;
    layer6_outputs(11715) <= not (a and b);
    layer6_outputs(11716) <= not a or b;
    layer6_outputs(11717) <= not (a xor b);
    layer6_outputs(11718) <= a xor b;
    layer6_outputs(11719) <= not a;
    layer6_outputs(11720) <= not b or a;
    layer6_outputs(11721) <= not a;
    layer6_outputs(11722) <= a xor b;
    layer6_outputs(11723) <= a or b;
    layer6_outputs(11724) <= a;
    layer6_outputs(11725) <= not a;
    layer6_outputs(11726) <= b;
    layer6_outputs(11727) <= not b;
    layer6_outputs(11728) <= not a;
    layer6_outputs(11729) <= a;
    layer6_outputs(11730) <= not b or a;
    layer6_outputs(11731) <= not b;
    layer6_outputs(11732) <= not b;
    layer6_outputs(11733) <= a;
    layer6_outputs(11734) <= not (a or b);
    layer6_outputs(11735) <= a and b;
    layer6_outputs(11736) <= b and not a;
    layer6_outputs(11737) <= not b;
    layer6_outputs(11738) <= not b;
    layer6_outputs(11739) <= not (a or b);
    layer6_outputs(11740) <= not b;
    layer6_outputs(11741) <= b;
    layer6_outputs(11742) <= not b;
    layer6_outputs(11743) <= not (a or b);
    layer6_outputs(11744) <= b;
    layer6_outputs(11745) <= b;
    layer6_outputs(11746) <= a and not b;
    layer6_outputs(11747) <= a xor b;
    layer6_outputs(11748) <= b;
    layer6_outputs(11749) <= not b;
    layer6_outputs(11750) <= not b;
    layer6_outputs(11751) <= a xor b;
    layer6_outputs(11752) <= a xor b;
    layer6_outputs(11753) <= a;
    layer6_outputs(11754) <= not (a xor b);
    layer6_outputs(11755) <= not (a xor b);
    layer6_outputs(11756) <= not (a or b);
    layer6_outputs(11757) <= b;
    layer6_outputs(11758) <= not b;
    layer6_outputs(11759) <= a and b;
    layer6_outputs(11760) <= not a;
    layer6_outputs(11761) <= not a;
    layer6_outputs(11762) <= a;
    layer6_outputs(11763) <= a or b;
    layer6_outputs(11764) <= not a;
    layer6_outputs(11765) <= b;
    layer6_outputs(11766) <= b;
    layer6_outputs(11767) <= not b;
    layer6_outputs(11768) <= not (a xor b);
    layer6_outputs(11769) <= b;
    layer6_outputs(11770) <= a xor b;
    layer6_outputs(11771) <= b;
    layer6_outputs(11772) <= not a;
    layer6_outputs(11773) <= a;
    layer6_outputs(11774) <= not (a xor b);
    layer6_outputs(11775) <= a xor b;
    layer6_outputs(11776) <= not a;
    layer6_outputs(11777) <= b;
    layer6_outputs(11778) <= not a;
    layer6_outputs(11779) <= not b or a;
    layer6_outputs(11780) <= a and b;
    layer6_outputs(11781) <= a and not b;
    layer6_outputs(11782) <= not (a or b);
    layer6_outputs(11783) <= not b;
    layer6_outputs(11784) <= '0';
    layer6_outputs(11785) <= not b or a;
    layer6_outputs(11786) <= not (a xor b);
    layer6_outputs(11787) <= not (a and b);
    layer6_outputs(11788) <= b and not a;
    layer6_outputs(11789) <= not (a or b);
    layer6_outputs(11790) <= not (a xor b);
    layer6_outputs(11791) <= not (a xor b);
    layer6_outputs(11792) <= not b;
    layer6_outputs(11793) <= not b;
    layer6_outputs(11794) <= not b;
    layer6_outputs(11795) <= a and not b;
    layer6_outputs(11796) <= not b;
    layer6_outputs(11797) <= a or b;
    layer6_outputs(11798) <= a xor b;
    layer6_outputs(11799) <= not (a xor b);
    layer6_outputs(11800) <= a xor b;
    layer6_outputs(11801) <= not b;
    layer6_outputs(11802) <= not (a xor b);
    layer6_outputs(11803) <= not (a xor b);
    layer6_outputs(11804) <= b;
    layer6_outputs(11805) <= not (a xor b);
    layer6_outputs(11806) <= a and b;
    layer6_outputs(11807) <= a xor b;
    layer6_outputs(11808) <= not b;
    layer6_outputs(11809) <= a;
    layer6_outputs(11810) <= a xor b;
    layer6_outputs(11811) <= not b;
    layer6_outputs(11812) <= a and b;
    layer6_outputs(11813) <= a or b;
    layer6_outputs(11814) <= not b;
    layer6_outputs(11815) <= not a;
    layer6_outputs(11816) <= b;
    layer6_outputs(11817) <= not a or b;
    layer6_outputs(11818) <= not (a xor b);
    layer6_outputs(11819) <= b and not a;
    layer6_outputs(11820) <= a xor b;
    layer6_outputs(11821) <= b;
    layer6_outputs(11822) <= not (a or b);
    layer6_outputs(11823) <= not a;
    layer6_outputs(11824) <= '1';
    layer6_outputs(11825) <= a;
    layer6_outputs(11826) <= not (a or b);
    layer6_outputs(11827) <= not (a and b);
    layer6_outputs(11828) <= not b;
    layer6_outputs(11829) <= a;
    layer6_outputs(11830) <= b;
    layer6_outputs(11831) <= not (a xor b);
    layer6_outputs(11832) <= a and b;
    layer6_outputs(11833) <= not a;
    layer6_outputs(11834) <= not (a xor b);
    layer6_outputs(11835) <= a xor b;
    layer6_outputs(11836) <= not a or b;
    layer6_outputs(11837) <= a and b;
    layer6_outputs(11838) <= a and not b;
    layer6_outputs(11839) <= not (a and b);
    layer6_outputs(11840) <= not (a or b);
    layer6_outputs(11841) <= not (a and b);
    layer6_outputs(11842) <= not (a and b);
    layer6_outputs(11843) <= not a or b;
    layer6_outputs(11844) <= a and not b;
    layer6_outputs(11845) <= not a;
    layer6_outputs(11846) <= b and not a;
    layer6_outputs(11847) <= b and not a;
    layer6_outputs(11848) <= b;
    layer6_outputs(11849) <= not b;
    layer6_outputs(11850) <= not b;
    layer6_outputs(11851) <= b and not a;
    layer6_outputs(11852) <= '0';
    layer6_outputs(11853) <= not (a xor b);
    layer6_outputs(11854) <= not b;
    layer6_outputs(11855) <= a and not b;
    layer6_outputs(11856) <= not a;
    layer6_outputs(11857) <= b and not a;
    layer6_outputs(11858) <= not a or b;
    layer6_outputs(11859) <= a or b;
    layer6_outputs(11860) <= not a;
    layer6_outputs(11861) <= not (a xor b);
    layer6_outputs(11862) <= not b or a;
    layer6_outputs(11863) <= not b or a;
    layer6_outputs(11864) <= not b or a;
    layer6_outputs(11865) <= not a;
    layer6_outputs(11866) <= a xor b;
    layer6_outputs(11867) <= not b;
    layer6_outputs(11868) <= not b;
    layer6_outputs(11869) <= not a;
    layer6_outputs(11870) <= not a;
    layer6_outputs(11871) <= a;
    layer6_outputs(11872) <= not b;
    layer6_outputs(11873) <= a xor b;
    layer6_outputs(11874) <= not b;
    layer6_outputs(11875) <= b and not a;
    layer6_outputs(11876) <= a;
    layer6_outputs(11877) <= not b or a;
    layer6_outputs(11878) <= a;
    layer6_outputs(11879) <= not b;
    layer6_outputs(11880) <= not (a or b);
    layer6_outputs(11881) <= a;
    layer6_outputs(11882) <= not b or a;
    layer6_outputs(11883) <= not b;
    layer6_outputs(11884) <= a;
    layer6_outputs(11885) <= not a;
    layer6_outputs(11886) <= a or b;
    layer6_outputs(11887) <= a;
    layer6_outputs(11888) <= not (a xor b);
    layer6_outputs(11889) <= '1';
    layer6_outputs(11890) <= a xor b;
    layer6_outputs(11891) <= not b or a;
    layer6_outputs(11892) <= a and not b;
    layer6_outputs(11893) <= not (a xor b);
    layer6_outputs(11894) <= not b or a;
    layer6_outputs(11895) <= a and not b;
    layer6_outputs(11896) <= not a;
    layer6_outputs(11897) <= b;
    layer6_outputs(11898) <= a and not b;
    layer6_outputs(11899) <= a;
    layer6_outputs(11900) <= a;
    layer6_outputs(11901) <= b;
    layer6_outputs(11902) <= a xor b;
    layer6_outputs(11903) <= not b;
    layer6_outputs(11904) <= b;
    layer6_outputs(11905) <= b and not a;
    layer6_outputs(11906) <= not a or b;
    layer6_outputs(11907) <= not a;
    layer6_outputs(11908) <= a;
    layer6_outputs(11909) <= not b;
    layer6_outputs(11910) <= a xor b;
    layer6_outputs(11911) <= b;
    layer6_outputs(11912) <= not b;
    layer6_outputs(11913) <= not b;
    layer6_outputs(11914) <= a;
    layer6_outputs(11915) <= not (a or b);
    layer6_outputs(11916) <= not (a xor b);
    layer6_outputs(11917) <= a and not b;
    layer6_outputs(11918) <= not (a and b);
    layer6_outputs(11919) <= not a;
    layer6_outputs(11920) <= not a or b;
    layer6_outputs(11921) <= b;
    layer6_outputs(11922) <= not (a and b);
    layer6_outputs(11923) <= not a;
    layer6_outputs(11924) <= a and b;
    layer6_outputs(11925) <= not a or b;
    layer6_outputs(11926) <= not a;
    layer6_outputs(11927) <= b;
    layer6_outputs(11928) <= a xor b;
    layer6_outputs(11929) <= not a;
    layer6_outputs(11930) <= not (a xor b);
    layer6_outputs(11931) <= a xor b;
    layer6_outputs(11932) <= not b;
    layer6_outputs(11933) <= b;
    layer6_outputs(11934) <= not b;
    layer6_outputs(11935) <= not a;
    layer6_outputs(11936) <= not (a and b);
    layer6_outputs(11937) <= not b;
    layer6_outputs(11938) <= a;
    layer6_outputs(11939) <= a;
    layer6_outputs(11940) <= not a;
    layer6_outputs(11941) <= b;
    layer6_outputs(11942) <= not b;
    layer6_outputs(11943) <= not (a xor b);
    layer6_outputs(11944) <= a xor b;
    layer6_outputs(11945) <= a;
    layer6_outputs(11946) <= a xor b;
    layer6_outputs(11947) <= a and not b;
    layer6_outputs(11948) <= not b or a;
    layer6_outputs(11949) <= a;
    layer6_outputs(11950) <= '0';
    layer6_outputs(11951) <= b and not a;
    layer6_outputs(11952) <= not (a xor b);
    layer6_outputs(11953) <= b;
    layer6_outputs(11954) <= a xor b;
    layer6_outputs(11955) <= not a;
    layer6_outputs(11956) <= a xor b;
    layer6_outputs(11957) <= b;
    layer6_outputs(11958) <= b;
    layer6_outputs(11959) <= b and not a;
    layer6_outputs(11960) <= b;
    layer6_outputs(11961) <= not b or a;
    layer6_outputs(11962) <= not b;
    layer6_outputs(11963) <= a xor b;
    layer6_outputs(11964) <= b;
    layer6_outputs(11965) <= not (a xor b);
    layer6_outputs(11966) <= not a;
    layer6_outputs(11967) <= a xor b;
    layer6_outputs(11968) <= not (a xor b);
    layer6_outputs(11969) <= a;
    layer6_outputs(11970) <= not (a or b);
    layer6_outputs(11971) <= a xor b;
    layer6_outputs(11972) <= a and not b;
    layer6_outputs(11973) <= not (a or b);
    layer6_outputs(11974) <= not a;
    layer6_outputs(11975) <= b and not a;
    layer6_outputs(11976) <= b;
    layer6_outputs(11977) <= b;
    layer6_outputs(11978) <= a and b;
    layer6_outputs(11979) <= a xor b;
    layer6_outputs(11980) <= not (a xor b);
    layer6_outputs(11981) <= not b or a;
    layer6_outputs(11982) <= not b;
    layer6_outputs(11983) <= not a;
    layer6_outputs(11984) <= not (a or b);
    layer6_outputs(11985) <= not a;
    layer6_outputs(11986) <= a;
    layer6_outputs(11987) <= a xor b;
    layer6_outputs(11988) <= not (a or b);
    layer6_outputs(11989) <= not a;
    layer6_outputs(11990) <= not b;
    layer6_outputs(11991) <= not (a xor b);
    layer6_outputs(11992) <= b;
    layer6_outputs(11993) <= '0';
    layer6_outputs(11994) <= not a;
    layer6_outputs(11995) <= a;
    layer6_outputs(11996) <= not b or a;
    layer6_outputs(11997) <= not b;
    layer6_outputs(11998) <= a xor b;
    layer6_outputs(11999) <= not (a and b);
    layer6_outputs(12000) <= a;
    layer6_outputs(12001) <= a;
    layer6_outputs(12002) <= not (a and b);
    layer6_outputs(12003) <= a;
    layer6_outputs(12004) <= not (a and b);
    layer6_outputs(12005) <= a xor b;
    layer6_outputs(12006) <= a xor b;
    layer6_outputs(12007) <= not b or a;
    layer6_outputs(12008) <= not a;
    layer6_outputs(12009) <= not b;
    layer6_outputs(12010) <= b and not a;
    layer6_outputs(12011) <= not a;
    layer6_outputs(12012) <= not (a or b);
    layer6_outputs(12013) <= a and not b;
    layer6_outputs(12014) <= not b;
    layer6_outputs(12015) <= not b or a;
    layer6_outputs(12016) <= not (a xor b);
    layer6_outputs(12017) <= not a or b;
    layer6_outputs(12018) <= a;
    layer6_outputs(12019) <= not a;
    layer6_outputs(12020) <= '1';
    layer6_outputs(12021) <= not b;
    layer6_outputs(12022) <= not a;
    layer6_outputs(12023) <= a;
    layer6_outputs(12024) <= not b;
    layer6_outputs(12025) <= not (a xor b);
    layer6_outputs(12026) <= not b or a;
    layer6_outputs(12027) <= a;
    layer6_outputs(12028) <= not b;
    layer6_outputs(12029) <= b;
    layer6_outputs(12030) <= not a;
    layer6_outputs(12031) <= a;
    layer6_outputs(12032) <= a and b;
    layer6_outputs(12033) <= not a;
    layer6_outputs(12034) <= a;
    layer6_outputs(12035) <= a or b;
    layer6_outputs(12036) <= not (a xor b);
    layer6_outputs(12037) <= a xor b;
    layer6_outputs(12038) <= not b;
    layer6_outputs(12039) <= not (a xor b);
    layer6_outputs(12040) <= a and not b;
    layer6_outputs(12041) <= b;
    layer6_outputs(12042) <= not a;
    layer6_outputs(12043) <= a;
    layer6_outputs(12044) <= not b or a;
    layer6_outputs(12045) <= b;
    layer6_outputs(12046) <= a;
    layer6_outputs(12047) <= not (a and b);
    layer6_outputs(12048) <= a;
    layer6_outputs(12049) <= a xor b;
    layer6_outputs(12050) <= not (a xor b);
    layer6_outputs(12051) <= a and not b;
    layer6_outputs(12052) <= a;
    layer6_outputs(12053) <= not (a or b);
    layer6_outputs(12054) <= not (a xor b);
    layer6_outputs(12055) <= a;
    layer6_outputs(12056) <= not b;
    layer6_outputs(12057) <= b;
    layer6_outputs(12058) <= b;
    layer6_outputs(12059) <= not a or b;
    layer6_outputs(12060) <= a;
    layer6_outputs(12061) <= not a;
    layer6_outputs(12062) <= b;
    layer6_outputs(12063) <= a or b;
    layer6_outputs(12064) <= not b or a;
    layer6_outputs(12065) <= not a;
    layer6_outputs(12066) <= not a or b;
    layer6_outputs(12067) <= b;
    layer6_outputs(12068) <= a xor b;
    layer6_outputs(12069) <= not b;
    layer6_outputs(12070) <= not b or a;
    layer6_outputs(12071) <= b;
    layer6_outputs(12072) <= b;
    layer6_outputs(12073) <= a and not b;
    layer6_outputs(12074) <= a and b;
    layer6_outputs(12075) <= b and not a;
    layer6_outputs(12076) <= b;
    layer6_outputs(12077) <= b and not a;
    layer6_outputs(12078) <= b;
    layer6_outputs(12079) <= a and not b;
    layer6_outputs(12080) <= not a or b;
    layer6_outputs(12081) <= a;
    layer6_outputs(12082) <= a;
    layer6_outputs(12083) <= not (a xor b);
    layer6_outputs(12084) <= a xor b;
    layer6_outputs(12085) <= a and b;
    layer6_outputs(12086) <= b;
    layer6_outputs(12087) <= a xor b;
    layer6_outputs(12088) <= a xor b;
    layer6_outputs(12089) <= a or b;
    layer6_outputs(12090) <= not b or a;
    layer6_outputs(12091) <= not a;
    layer6_outputs(12092) <= a;
    layer6_outputs(12093) <= not a;
    layer6_outputs(12094) <= a or b;
    layer6_outputs(12095) <= a xor b;
    layer6_outputs(12096) <= a xor b;
    layer6_outputs(12097) <= not b or a;
    layer6_outputs(12098) <= not b or a;
    layer6_outputs(12099) <= not b;
    layer6_outputs(12100) <= a and not b;
    layer6_outputs(12101) <= b and not a;
    layer6_outputs(12102) <= a and b;
    layer6_outputs(12103) <= a and not b;
    layer6_outputs(12104) <= b;
    layer6_outputs(12105) <= not a;
    layer6_outputs(12106) <= b;
    layer6_outputs(12107) <= b and not a;
    layer6_outputs(12108) <= a or b;
    layer6_outputs(12109) <= a and not b;
    layer6_outputs(12110) <= not a;
    layer6_outputs(12111) <= not a or b;
    layer6_outputs(12112) <= b;
    layer6_outputs(12113) <= not (a or b);
    layer6_outputs(12114) <= a xor b;
    layer6_outputs(12115) <= not b;
    layer6_outputs(12116) <= a or b;
    layer6_outputs(12117) <= a xor b;
    layer6_outputs(12118) <= b;
    layer6_outputs(12119) <= a;
    layer6_outputs(12120) <= not (a and b);
    layer6_outputs(12121) <= '0';
    layer6_outputs(12122) <= not a;
    layer6_outputs(12123) <= not a;
    layer6_outputs(12124) <= a xor b;
    layer6_outputs(12125) <= not (a or b);
    layer6_outputs(12126) <= not a or b;
    layer6_outputs(12127) <= b and not a;
    layer6_outputs(12128) <= '1';
    layer6_outputs(12129) <= b and not a;
    layer6_outputs(12130) <= not b or a;
    layer6_outputs(12131) <= b;
    layer6_outputs(12132) <= b;
    layer6_outputs(12133) <= a xor b;
    layer6_outputs(12134) <= not b;
    layer6_outputs(12135) <= b;
    layer6_outputs(12136) <= a or b;
    layer6_outputs(12137) <= a and b;
    layer6_outputs(12138) <= not a;
    layer6_outputs(12139) <= not b;
    layer6_outputs(12140) <= not a;
    layer6_outputs(12141) <= not (a xor b);
    layer6_outputs(12142) <= a xor b;
    layer6_outputs(12143) <= a and b;
    layer6_outputs(12144) <= b and not a;
    layer6_outputs(12145) <= a or b;
    layer6_outputs(12146) <= a and not b;
    layer6_outputs(12147) <= b and not a;
    layer6_outputs(12148) <= a;
    layer6_outputs(12149) <= b;
    layer6_outputs(12150) <= a and not b;
    layer6_outputs(12151) <= not (a xor b);
    layer6_outputs(12152) <= not b;
    layer6_outputs(12153) <= b;
    layer6_outputs(12154) <= not b;
    layer6_outputs(12155) <= not a;
    layer6_outputs(12156) <= b and not a;
    layer6_outputs(12157) <= not a or b;
    layer6_outputs(12158) <= a;
    layer6_outputs(12159) <= b;
    layer6_outputs(12160) <= not (a or b);
    layer6_outputs(12161) <= b;
    layer6_outputs(12162) <= not (a and b);
    layer6_outputs(12163) <= not (a xor b);
    layer6_outputs(12164) <= a;
    layer6_outputs(12165) <= not (a xor b);
    layer6_outputs(12166) <= not (a and b);
    layer6_outputs(12167) <= not (a and b);
    layer6_outputs(12168) <= not (a and b);
    layer6_outputs(12169) <= not a or b;
    layer6_outputs(12170) <= not (a xor b);
    layer6_outputs(12171) <= not a;
    layer6_outputs(12172) <= a xor b;
    layer6_outputs(12173) <= not (a xor b);
    layer6_outputs(12174) <= not b;
    layer6_outputs(12175) <= a or b;
    layer6_outputs(12176) <= not a;
    layer6_outputs(12177) <= a xor b;
    layer6_outputs(12178) <= a and not b;
    layer6_outputs(12179) <= a;
    layer6_outputs(12180) <= b;
    layer6_outputs(12181) <= not a or b;
    layer6_outputs(12182) <= not a or b;
    layer6_outputs(12183) <= not (a and b);
    layer6_outputs(12184) <= b and not a;
    layer6_outputs(12185) <= a;
    layer6_outputs(12186) <= not (a and b);
    layer6_outputs(12187) <= a xor b;
    layer6_outputs(12188) <= a;
    layer6_outputs(12189) <= not a;
    layer6_outputs(12190) <= not b;
    layer6_outputs(12191) <= not a;
    layer6_outputs(12192) <= not (a or b);
    layer6_outputs(12193) <= b;
    layer6_outputs(12194) <= a xor b;
    layer6_outputs(12195) <= b and not a;
    layer6_outputs(12196) <= a xor b;
    layer6_outputs(12197) <= a;
    layer6_outputs(12198) <= not b;
    layer6_outputs(12199) <= b and not a;
    layer6_outputs(12200) <= '0';
    layer6_outputs(12201) <= not (a xor b);
    layer6_outputs(12202) <= not (a or b);
    layer6_outputs(12203) <= not (a xor b);
    layer6_outputs(12204) <= not (a or b);
    layer6_outputs(12205) <= b;
    layer6_outputs(12206) <= not (a xor b);
    layer6_outputs(12207) <= not b;
    layer6_outputs(12208) <= not a or b;
    layer6_outputs(12209) <= a;
    layer6_outputs(12210) <= not a;
    layer6_outputs(12211) <= not (a or b);
    layer6_outputs(12212) <= not a;
    layer6_outputs(12213) <= not a;
    layer6_outputs(12214) <= b;
    layer6_outputs(12215) <= not (a xor b);
    layer6_outputs(12216) <= b;
    layer6_outputs(12217) <= a;
    layer6_outputs(12218) <= not b;
    layer6_outputs(12219) <= not a;
    layer6_outputs(12220) <= a xor b;
    layer6_outputs(12221) <= not a or b;
    layer6_outputs(12222) <= not (a xor b);
    layer6_outputs(12223) <= not b or a;
    layer6_outputs(12224) <= b and not a;
    layer6_outputs(12225) <= a;
    layer6_outputs(12226) <= a or b;
    layer6_outputs(12227) <= not b;
    layer6_outputs(12228) <= not b or a;
    layer6_outputs(12229) <= a;
    layer6_outputs(12230) <= not b;
    layer6_outputs(12231) <= not b;
    layer6_outputs(12232) <= not b;
    layer6_outputs(12233) <= not a;
    layer6_outputs(12234) <= not b;
    layer6_outputs(12235) <= not a;
    layer6_outputs(12236) <= not b;
    layer6_outputs(12237) <= a;
    layer6_outputs(12238) <= not b;
    layer6_outputs(12239) <= not (a or b);
    layer6_outputs(12240) <= a or b;
    layer6_outputs(12241) <= not (a or b);
    layer6_outputs(12242) <= not (a xor b);
    layer6_outputs(12243) <= not b;
    layer6_outputs(12244) <= a;
    layer6_outputs(12245) <= not b or a;
    layer6_outputs(12246) <= not (a xor b);
    layer6_outputs(12247) <= a;
    layer6_outputs(12248) <= not (a and b);
    layer6_outputs(12249) <= not (a xor b);
    layer6_outputs(12250) <= a or b;
    layer6_outputs(12251) <= a xor b;
    layer6_outputs(12252) <= a;
    layer6_outputs(12253) <= not (a and b);
    layer6_outputs(12254) <= not b;
    layer6_outputs(12255) <= not a;
    layer6_outputs(12256) <= a xor b;
    layer6_outputs(12257) <= a xor b;
    layer6_outputs(12258) <= b;
    layer6_outputs(12259) <= not a;
    layer6_outputs(12260) <= a;
    layer6_outputs(12261) <= not a;
    layer6_outputs(12262) <= not (a xor b);
    layer6_outputs(12263) <= a xor b;
    layer6_outputs(12264) <= not a;
    layer6_outputs(12265) <= b;
    layer6_outputs(12266) <= not b;
    layer6_outputs(12267) <= b;
    layer6_outputs(12268) <= a;
    layer6_outputs(12269) <= a;
    layer6_outputs(12270) <= b;
    layer6_outputs(12271) <= b;
    layer6_outputs(12272) <= a xor b;
    layer6_outputs(12273) <= a xor b;
    layer6_outputs(12274) <= a xor b;
    layer6_outputs(12275) <= not a;
    layer6_outputs(12276) <= b;
    layer6_outputs(12277) <= not a or b;
    layer6_outputs(12278) <= not a;
    layer6_outputs(12279) <= not b or a;
    layer6_outputs(12280) <= a and not b;
    layer6_outputs(12281) <= not (a xor b);
    layer6_outputs(12282) <= not (a xor b);
    layer6_outputs(12283) <= not b;
    layer6_outputs(12284) <= b;
    layer6_outputs(12285) <= not b;
    layer6_outputs(12286) <= a xor b;
    layer6_outputs(12287) <= b;
    layer6_outputs(12288) <= b and not a;
    layer6_outputs(12289) <= a or b;
    layer6_outputs(12290) <= not (a and b);
    layer6_outputs(12291) <= not (a or b);
    layer6_outputs(12292) <= a;
    layer6_outputs(12293) <= a and b;
    layer6_outputs(12294) <= a xor b;
    layer6_outputs(12295) <= b;
    layer6_outputs(12296) <= not (a xor b);
    layer6_outputs(12297) <= a;
    layer6_outputs(12298) <= not b;
    layer6_outputs(12299) <= not b or a;
    layer6_outputs(12300) <= a;
    layer6_outputs(12301) <= b;
    layer6_outputs(12302) <= not (a xor b);
    layer6_outputs(12303) <= b;
    layer6_outputs(12304) <= not b;
    layer6_outputs(12305) <= a;
    layer6_outputs(12306) <= not a;
    layer6_outputs(12307) <= a and b;
    layer6_outputs(12308) <= a or b;
    layer6_outputs(12309) <= b;
    layer6_outputs(12310) <= not (a xor b);
    layer6_outputs(12311) <= a;
    layer6_outputs(12312) <= not b;
    layer6_outputs(12313) <= not (a xor b);
    layer6_outputs(12314) <= a and not b;
    layer6_outputs(12315) <= a;
    layer6_outputs(12316) <= not b or a;
    layer6_outputs(12317) <= a;
    layer6_outputs(12318) <= a and not b;
    layer6_outputs(12319) <= not (a xor b);
    layer6_outputs(12320) <= not (a or b);
    layer6_outputs(12321) <= a;
    layer6_outputs(12322) <= a or b;
    layer6_outputs(12323) <= not a;
    layer6_outputs(12324) <= not a;
    layer6_outputs(12325) <= a xor b;
    layer6_outputs(12326) <= not b;
    layer6_outputs(12327) <= not b or a;
    layer6_outputs(12328) <= b;
    layer6_outputs(12329) <= b;
    layer6_outputs(12330) <= not (a xor b);
    layer6_outputs(12331) <= a xor b;
    layer6_outputs(12332) <= b;
    layer6_outputs(12333) <= not a or b;
    layer6_outputs(12334) <= not (a and b);
    layer6_outputs(12335) <= not (a and b);
    layer6_outputs(12336) <= not (a xor b);
    layer6_outputs(12337) <= not b;
    layer6_outputs(12338) <= not b;
    layer6_outputs(12339) <= b;
    layer6_outputs(12340) <= b and not a;
    layer6_outputs(12341) <= b;
    layer6_outputs(12342) <= not b;
    layer6_outputs(12343) <= b and not a;
    layer6_outputs(12344) <= b;
    layer6_outputs(12345) <= b;
    layer6_outputs(12346) <= b;
    layer6_outputs(12347) <= a and b;
    layer6_outputs(12348) <= not b;
    layer6_outputs(12349) <= not a;
    layer6_outputs(12350) <= not (a and b);
    layer6_outputs(12351) <= a;
    layer6_outputs(12352) <= not a;
    layer6_outputs(12353) <= a xor b;
    layer6_outputs(12354) <= not a or b;
    layer6_outputs(12355) <= not a;
    layer6_outputs(12356) <= a;
    layer6_outputs(12357) <= not b or a;
    layer6_outputs(12358) <= not (a xor b);
    layer6_outputs(12359) <= not b or a;
    layer6_outputs(12360) <= not b;
    layer6_outputs(12361) <= b;
    layer6_outputs(12362) <= not (a and b);
    layer6_outputs(12363) <= a and not b;
    layer6_outputs(12364) <= a xor b;
    layer6_outputs(12365) <= a;
    layer6_outputs(12366) <= b;
    layer6_outputs(12367) <= not a;
    layer6_outputs(12368) <= not a or b;
    layer6_outputs(12369) <= not a;
    layer6_outputs(12370) <= a and b;
    layer6_outputs(12371) <= not b;
    layer6_outputs(12372) <= a xor b;
    layer6_outputs(12373) <= b;
    layer6_outputs(12374) <= a and not b;
    layer6_outputs(12375) <= a;
    layer6_outputs(12376) <= not (a xor b);
    layer6_outputs(12377) <= b and not a;
    layer6_outputs(12378) <= a;
    layer6_outputs(12379) <= a;
    layer6_outputs(12380) <= not a;
    layer6_outputs(12381) <= not a;
    layer6_outputs(12382) <= b and not a;
    layer6_outputs(12383) <= a;
    layer6_outputs(12384) <= a;
    layer6_outputs(12385) <= a;
    layer6_outputs(12386) <= not (a xor b);
    layer6_outputs(12387) <= not (a xor b);
    layer6_outputs(12388) <= a xor b;
    layer6_outputs(12389) <= not (a or b);
    layer6_outputs(12390) <= not a or b;
    layer6_outputs(12391) <= b;
    layer6_outputs(12392) <= b;
    layer6_outputs(12393) <= b and not a;
    layer6_outputs(12394) <= not a;
    layer6_outputs(12395) <= not b;
    layer6_outputs(12396) <= not (a or b);
    layer6_outputs(12397) <= b;
    layer6_outputs(12398) <= not b or a;
    layer6_outputs(12399) <= not (a xor b);
    layer6_outputs(12400) <= not b;
    layer6_outputs(12401) <= a xor b;
    layer6_outputs(12402) <= not (a and b);
    layer6_outputs(12403) <= a xor b;
    layer6_outputs(12404) <= b;
    layer6_outputs(12405) <= not b;
    layer6_outputs(12406) <= not b or a;
    layer6_outputs(12407) <= not a;
    layer6_outputs(12408) <= not b;
    layer6_outputs(12409) <= not a;
    layer6_outputs(12410) <= a xor b;
    layer6_outputs(12411) <= not (a xor b);
    layer6_outputs(12412) <= b;
    layer6_outputs(12413) <= not b;
    layer6_outputs(12414) <= not (a or b);
    layer6_outputs(12415) <= b and not a;
    layer6_outputs(12416) <= a xor b;
    layer6_outputs(12417) <= not a;
    layer6_outputs(12418) <= not (a xor b);
    layer6_outputs(12419) <= not a;
    layer6_outputs(12420) <= not (a xor b);
    layer6_outputs(12421) <= not (a xor b);
    layer6_outputs(12422) <= not (a or b);
    layer6_outputs(12423) <= a;
    layer6_outputs(12424) <= a and not b;
    layer6_outputs(12425) <= not a or b;
    layer6_outputs(12426) <= not (a or b);
    layer6_outputs(12427) <= a or b;
    layer6_outputs(12428) <= not b;
    layer6_outputs(12429) <= not a or b;
    layer6_outputs(12430) <= not (a xor b);
    layer6_outputs(12431) <= not a;
    layer6_outputs(12432) <= not (a xor b);
    layer6_outputs(12433) <= not (a or b);
    layer6_outputs(12434) <= not (a or b);
    layer6_outputs(12435) <= not (a xor b);
    layer6_outputs(12436) <= not b or a;
    layer6_outputs(12437) <= not a or b;
    layer6_outputs(12438) <= not a;
    layer6_outputs(12439) <= a xor b;
    layer6_outputs(12440) <= b;
    layer6_outputs(12441) <= '0';
    layer6_outputs(12442) <= not (a xor b);
    layer6_outputs(12443) <= not (a xor b);
    layer6_outputs(12444) <= not (a xor b);
    layer6_outputs(12445) <= a xor b;
    layer6_outputs(12446) <= not (a or b);
    layer6_outputs(12447) <= not b or a;
    layer6_outputs(12448) <= not (a xor b);
    layer6_outputs(12449) <= a and b;
    layer6_outputs(12450) <= not a;
    layer6_outputs(12451) <= not (a xor b);
    layer6_outputs(12452) <= not (a xor b);
    layer6_outputs(12453) <= not b;
    layer6_outputs(12454) <= not (a xor b);
    layer6_outputs(12455) <= a and not b;
    layer6_outputs(12456) <= a and not b;
    layer6_outputs(12457) <= a and not b;
    layer6_outputs(12458) <= not (a and b);
    layer6_outputs(12459) <= a and not b;
    layer6_outputs(12460) <= b;
    layer6_outputs(12461) <= not a or b;
    layer6_outputs(12462) <= not a or b;
    layer6_outputs(12463) <= a;
    layer6_outputs(12464) <= not a;
    layer6_outputs(12465) <= not b;
    layer6_outputs(12466) <= a;
    layer6_outputs(12467) <= a xor b;
    layer6_outputs(12468) <= not (a and b);
    layer6_outputs(12469) <= a;
    layer6_outputs(12470) <= a and b;
    layer6_outputs(12471) <= not b or a;
    layer6_outputs(12472) <= not a;
    layer6_outputs(12473) <= not a or b;
    layer6_outputs(12474) <= not b or a;
    layer6_outputs(12475) <= not (a xor b);
    layer6_outputs(12476) <= not (a or b);
    layer6_outputs(12477) <= a;
    layer6_outputs(12478) <= a and b;
    layer6_outputs(12479) <= b;
    layer6_outputs(12480) <= not a;
    layer6_outputs(12481) <= b and not a;
    layer6_outputs(12482) <= b and not a;
    layer6_outputs(12483) <= a and not b;
    layer6_outputs(12484) <= not a;
    layer6_outputs(12485) <= a and b;
    layer6_outputs(12486) <= not (a or b);
    layer6_outputs(12487) <= a xor b;
    layer6_outputs(12488) <= a;
    layer6_outputs(12489) <= a and b;
    layer6_outputs(12490) <= a and b;
    layer6_outputs(12491) <= b and not a;
    layer6_outputs(12492) <= a or b;
    layer6_outputs(12493) <= not b or a;
    layer6_outputs(12494) <= a;
    layer6_outputs(12495) <= not a;
    layer6_outputs(12496) <= a xor b;
    layer6_outputs(12497) <= not (a and b);
    layer6_outputs(12498) <= a;
    layer6_outputs(12499) <= a and b;
    layer6_outputs(12500) <= not (a and b);
    layer6_outputs(12501) <= '0';
    layer6_outputs(12502) <= a xor b;
    layer6_outputs(12503) <= a or b;
    layer6_outputs(12504) <= not b;
    layer6_outputs(12505) <= a or b;
    layer6_outputs(12506) <= b;
    layer6_outputs(12507) <= not (a or b);
    layer6_outputs(12508) <= not b or a;
    layer6_outputs(12509) <= not (a xor b);
    layer6_outputs(12510) <= not a;
    layer6_outputs(12511) <= not a;
    layer6_outputs(12512) <= a;
    layer6_outputs(12513) <= not (a xor b);
    layer6_outputs(12514) <= a;
    layer6_outputs(12515) <= b;
    layer6_outputs(12516) <= a or b;
    layer6_outputs(12517) <= not b;
    layer6_outputs(12518) <= not a;
    layer6_outputs(12519) <= not a;
    layer6_outputs(12520) <= b;
    layer6_outputs(12521) <= not (a xor b);
    layer6_outputs(12522) <= b;
    layer6_outputs(12523) <= a;
    layer6_outputs(12524) <= a;
    layer6_outputs(12525) <= b and not a;
    layer6_outputs(12526) <= not a;
    layer6_outputs(12527) <= not (a and b);
    layer6_outputs(12528) <= a xor b;
    layer6_outputs(12529) <= not (a xor b);
    layer6_outputs(12530) <= b and not a;
    layer6_outputs(12531) <= a;
    layer6_outputs(12532) <= b and not a;
    layer6_outputs(12533) <= b and not a;
    layer6_outputs(12534) <= not b;
    layer6_outputs(12535) <= not (a xor b);
    layer6_outputs(12536) <= a xor b;
    layer6_outputs(12537) <= not (a or b);
    layer6_outputs(12538) <= not a;
    layer6_outputs(12539) <= not a or b;
    layer6_outputs(12540) <= not (a xor b);
    layer6_outputs(12541) <= not a;
    layer6_outputs(12542) <= a;
    layer6_outputs(12543) <= b;
    layer6_outputs(12544) <= not a or b;
    layer6_outputs(12545) <= a and b;
    layer6_outputs(12546) <= a and not b;
    layer6_outputs(12547) <= a and b;
    layer6_outputs(12548) <= not (a and b);
    layer6_outputs(12549) <= not a;
    layer6_outputs(12550) <= not b or a;
    layer6_outputs(12551) <= a and not b;
    layer6_outputs(12552) <= a or b;
    layer6_outputs(12553) <= a and not b;
    layer6_outputs(12554) <= b and not a;
    layer6_outputs(12555) <= not a;
    layer6_outputs(12556) <= b;
    layer6_outputs(12557) <= a and not b;
    layer6_outputs(12558) <= b;
    layer6_outputs(12559) <= not a;
    layer6_outputs(12560) <= b and not a;
    layer6_outputs(12561) <= b;
    layer6_outputs(12562) <= not (a and b);
    layer6_outputs(12563) <= not (a xor b);
    layer6_outputs(12564) <= not b;
    layer6_outputs(12565) <= not (a xor b);
    layer6_outputs(12566) <= a;
    layer6_outputs(12567) <= b and not a;
    layer6_outputs(12568) <= a xor b;
    layer6_outputs(12569) <= a and b;
    layer6_outputs(12570) <= b and not a;
    layer6_outputs(12571) <= not b;
    layer6_outputs(12572) <= a xor b;
    layer6_outputs(12573) <= not (a xor b);
    layer6_outputs(12574) <= not a;
    layer6_outputs(12575) <= b;
    layer6_outputs(12576) <= a and not b;
    layer6_outputs(12577) <= not (a xor b);
    layer6_outputs(12578) <= not b or a;
    layer6_outputs(12579) <= a;
    layer6_outputs(12580) <= not b or a;
    layer6_outputs(12581) <= not (a xor b);
    layer6_outputs(12582) <= not a;
    layer6_outputs(12583) <= not a or b;
    layer6_outputs(12584) <= b and not a;
    layer6_outputs(12585) <= not a or b;
    layer6_outputs(12586) <= not a;
    layer6_outputs(12587) <= a and b;
    layer6_outputs(12588) <= not a;
    layer6_outputs(12589) <= not (a xor b);
    layer6_outputs(12590) <= not a;
    layer6_outputs(12591) <= not a or b;
    layer6_outputs(12592) <= '1';
    layer6_outputs(12593) <= b;
    layer6_outputs(12594) <= b;
    layer6_outputs(12595) <= not b;
    layer6_outputs(12596) <= not (a or b);
    layer6_outputs(12597) <= b;
    layer6_outputs(12598) <= not a or b;
    layer6_outputs(12599) <= b;
    layer6_outputs(12600) <= b;
    layer6_outputs(12601) <= a and b;
    layer6_outputs(12602) <= b;
    layer6_outputs(12603) <= a xor b;
    layer6_outputs(12604) <= a or b;
    layer6_outputs(12605) <= a;
    layer6_outputs(12606) <= not (a or b);
    layer6_outputs(12607) <= a;
    layer6_outputs(12608) <= '0';
    layer6_outputs(12609) <= not b or a;
    layer6_outputs(12610) <= a and b;
    layer6_outputs(12611) <= not (a xor b);
    layer6_outputs(12612) <= not (a xor b);
    layer6_outputs(12613) <= b;
    layer6_outputs(12614) <= not (a xor b);
    layer6_outputs(12615) <= not a;
    layer6_outputs(12616) <= not a;
    layer6_outputs(12617) <= not b or a;
    layer6_outputs(12618) <= a;
    layer6_outputs(12619) <= b;
    layer6_outputs(12620) <= not b;
    layer6_outputs(12621) <= a and not b;
    layer6_outputs(12622) <= a;
    layer6_outputs(12623) <= not b;
    layer6_outputs(12624) <= b;
    layer6_outputs(12625) <= b;
    layer6_outputs(12626) <= not a;
    layer6_outputs(12627) <= not (a xor b);
    layer6_outputs(12628) <= not a;
    layer6_outputs(12629) <= not a or b;
    layer6_outputs(12630) <= not b or a;
    layer6_outputs(12631) <= a and not b;
    layer6_outputs(12632) <= not b or a;
    layer6_outputs(12633) <= not b;
    layer6_outputs(12634) <= not b or a;
    layer6_outputs(12635) <= a;
    layer6_outputs(12636) <= a and b;
    layer6_outputs(12637) <= b;
    layer6_outputs(12638) <= b;
    layer6_outputs(12639) <= b;
    layer6_outputs(12640) <= a;
    layer6_outputs(12641) <= not (a or b);
    layer6_outputs(12642) <= not (a or b);
    layer6_outputs(12643) <= a xor b;
    layer6_outputs(12644) <= a;
    layer6_outputs(12645) <= not b or a;
    layer6_outputs(12646) <= not b;
    layer6_outputs(12647) <= a;
    layer6_outputs(12648) <= not b;
    layer6_outputs(12649) <= a;
    layer6_outputs(12650) <= a;
    layer6_outputs(12651) <= not a;
    layer6_outputs(12652) <= not (a xor b);
    layer6_outputs(12653) <= a xor b;
    layer6_outputs(12654) <= not (a xor b);
    layer6_outputs(12655) <= not b;
    layer6_outputs(12656) <= not (a xor b);
    layer6_outputs(12657) <= not a;
    layer6_outputs(12658) <= not b;
    layer6_outputs(12659) <= not (a xor b);
    layer6_outputs(12660) <= a xor b;
    layer6_outputs(12661) <= a xor b;
    layer6_outputs(12662) <= a xor b;
    layer6_outputs(12663) <= a;
    layer6_outputs(12664) <= not a;
    layer6_outputs(12665) <= b and not a;
    layer6_outputs(12666) <= not b;
    layer6_outputs(12667) <= a;
    layer6_outputs(12668) <= b and not a;
    layer6_outputs(12669) <= a xor b;
    layer6_outputs(12670) <= not b or a;
    layer6_outputs(12671) <= not (a or b);
    layer6_outputs(12672) <= not a;
    layer6_outputs(12673) <= b and not a;
    layer6_outputs(12674) <= a;
    layer6_outputs(12675) <= a xor b;
    layer6_outputs(12676) <= not (a and b);
    layer6_outputs(12677) <= b;
    layer6_outputs(12678) <= a xor b;
    layer6_outputs(12679) <= a;
    layer6_outputs(12680) <= not a or b;
    layer6_outputs(12681) <= not b;
    layer6_outputs(12682) <= not b;
    layer6_outputs(12683) <= b;
    layer6_outputs(12684) <= not a;
    layer6_outputs(12685) <= a and b;
    layer6_outputs(12686) <= not (a or b);
    layer6_outputs(12687) <= not a;
    layer6_outputs(12688) <= not a or b;
    layer6_outputs(12689) <= not b;
    layer6_outputs(12690) <= not (a xor b);
    layer6_outputs(12691) <= not a;
    layer6_outputs(12692) <= not (a and b);
    layer6_outputs(12693) <= not (a and b);
    layer6_outputs(12694) <= a or b;
    layer6_outputs(12695) <= a xor b;
    layer6_outputs(12696) <= not a or b;
    layer6_outputs(12697) <= a;
    layer6_outputs(12698) <= b;
    layer6_outputs(12699) <= not (a xor b);
    layer6_outputs(12700) <= a;
    layer6_outputs(12701) <= b;
    layer6_outputs(12702) <= a or b;
    layer6_outputs(12703) <= not (a and b);
    layer6_outputs(12704) <= not b or a;
    layer6_outputs(12705) <= not a or b;
    layer6_outputs(12706) <= a and not b;
    layer6_outputs(12707) <= not b or a;
    layer6_outputs(12708) <= a and b;
    layer6_outputs(12709) <= a xor b;
    layer6_outputs(12710) <= not (a xor b);
    layer6_outputs(12711) <= not a;
    layer6_outputs(12712) <= not (a or b);
    layer6_outputs(12713) <= not (a xor b);
    layer6_outputs(12714) <= not b;
    layer6_outputs(12715) <= a;
    layer6_outputs(12716) <= a xor b;
    layer6_outputs(12717) <= a xor b;
    layer6_outputs(12718) <= b;
    layer6_outputs(12719) <= a xor b;
    layer6_outputs(12720) <= not (a or b);
    layer6_outputs(12721) <= a;
    layer6_outputs(12722) <= b;
    layer6_outputs(12723) <= not a;
    layer6_outputs(12724) <= a xor b;
    layer6_outputs(12725) <= a or b;
    layer6_outputs(12726) <= not b;
    layer6_outputs(12727) <= not b;
    layer6_outputs(12728) <= a and not b;
    layer6_outputs(12729) <= a or b;
    layer6_outputs(12730) <= a;
    layer6_outputs(12731) <= not (a or b);
    layer6_outputs(12732) <= a and not b;
    layer6_outputs(12733) <= not b;
    layer6_outputs(12734) <= not b or a;
    layer6_outputs(12735) <= not a;
    layer6_outputs(12736) <= a and not b;
    layer6_outputs(12737) <= not b;
    layer6_outputs(12738) <= b;
    layer6_outputs(12739) <= not b;
    layer6_outputs(12740) <= b and not a;
    layer6_outputs(12741) <= not a;
    layer6_outputs(12742) <= a or b;
    layer6_outputs(12743) <= not a;
    layer6_outputs(12744) <= not a or b;
    layer6_outputs(12745) <= not b;
    layer6_outputs(12746) <= not b;
    layer6_outputs(12747) <= not (a xor b);
    layer6_outputs(12748) <= a xor b;
    layer6_outputs(12749) <= not a;
    layer6_outputs(12750) <= not (a and b);
    layer6_outputs(12751) <= a and b;
    layer6_outputs(12752) <= b;
    layer6_outputs(12753) <= a xor b;
    layer6_outputs(12754) <= not (a and b);
    layer6_outputs(12755) <= not (a xor b);
    layer6_outputs(12756) <= not b or a;
    layer6_outputs(12757) <= a and not b;
    layer6_outputs(12758) <= a xor b;
    layer6_outputs(12759) <= not b;
    layer6_outputs(12760) <= not (a xor b);
    layer6_outputs(12761) <= not a;
    layer6_outputs(12762) <= not (a and b);
    layer6_outputs(12763) <= not b or a;
    layer6_outputs(12764) <= b;
    layer6_outputs(12765) <= a or b;
    layer6_outputs(12766) <= not b;
    layer6_outputs(12767) <= b;
    layer6_outputs(12768) <= b;
    layer6_outputs(12769) <= b;
    layer6_outputs(12770) <= not b or a;
    layer6_outputs(12771) <= not a;
    layer6_outputs(12772) <= not (a and b);
    layer6_outputs(12773) <= b and not a;
    layer6_outputs(12774) <= not (a xor b);
    layer6_outputs(12775) <= a xor b;
    layer6_outputs(12776) <= b;
    layer6_outputs(12777) <= not a;
    layer6_outputs(12778) <= b;
    layer6_outputs(12779) <= not (a xor b);
    layer6_outputs(12780) <= b;
    layer6_outputs(12781) <= b;
    layer6_outputs(12782) <= b;
    layer6_outputs(12783) <= a and not b;
    layer6_outputs(12784) <= not (a or b);
    layer6_outputs(12785) <= b and not a;
    layer6_outputs(12786) <= b;
    layer6_outputs(12787) <= not b;
    layer6_outputs(12788) <= not b;
    layer6_outputs(12789) <= a and not b;
    layer6_outputs(12790) <= not b or a;
    layer6_outputs(12791) <= not a;
    layer6_outputs(12792) <= not a;
    layer6_outputs(12793) <= b;
    layer6_outputs(12794) <= not (a xor b);
    layer6_outputs(12795) <= not a or b;
    layer6_outputs(12796) <= not (a xor b);
    layer6_outputs(12797) <= not a;
    layer6_outputs(12798) <= not (a xor b);
    layer6_outputs(12799) <= not a;
    outputs(0) <= b;
    outputs(1) <= a xor b;
    outputs(2) <= a or b;
    outputs(3) <= a xor b;
    outputs(4) <= not (a or b);
    outputs(5) <= a and not b;
    outputs(6) <= a and b;
    outputs(7) <= a;
    outputs(8) <= not a;
    outputs(9) <= a xor b;
    outputs(10) <= not b;
    outputs(11) <= b and not a;
    outputs(12) <= a and b;
    outputs(13) <= b;
    outputs(14) <= a or b;
    outputs(15) <= a xor b;
    outputs(16) <= not (a xor b);
    outputs(17) <= not (a xor b);
    outputs(18) <= b;
    outputs(19) <= b;
    outputs(20) <= not a;
    outputs(21) <= not (a xor b);
    outputs(22) <= a;
    outputs(23) <= not b;
    outputs(24) <= not (a or b);
    outputs(25) <= not (a xor b);
    outputs(26) <= a and b;
    outputs(27) <= a xor b;
    outputs(28) <= b;
    outputs(29) <= b and not a;
    outputs(30) <= b and not a;
    outputs(31) <= a xor b;
    outputs(32) <= a or b;
    outputs(33) <= a;
    outputs(34) <= not a;
    outputs(35) <= a;
    outputs(36) <= a or b;
    outputs(37) <= not (a or b);
    outputs(38) <= not b;
    outputs(39) <= a xor b;
    outputs(40) <= not b;
    outputs(41) <= a and not b;
    outputs(42) <= not (a xor b);
    outputs(43) <= a and b;
    outputs(44) <= not (a xor b);
    outputs(45) <= b;
    outputs(46) <= not b;
    outputs(47) <= a xor b;
    outputs(48) <= b and not a;
    outputs(49) <= a;
    outputs(50) <= not (a xor b);
    outputs(51) <= b;
    outputs(52) <= not (a or b);
    outputs(53) <= a xor b;
    outputs(54) <= not (a or b);
    outputs(55) <= a xor b;
    outputs(56) <= a and b;
    outputs(57) <= b;
    outputs(58) <= a and b;
    outputs(59) <= not a;
    outputs(60) <= not (a or b);
    outputs(61) <= a and not b;
    outputs(62) <= a and b;
    outputs(63) <= a xor b;
    outputs(64) <= a;
    outputs(65) <= not (a xor b);
    outputs(66) <= not a;
    outputs(67) <= b;
    outputs(68) <= not a;
    outputs(69) <= a;
    outputs(70) <= not (a or b);
    outputs(71) <= not a;
    outputs(72) <= not a;
    outputs(73) <= not b;
    outputs(74) <= not b;
    outputs(75) <= not b;
    outputs(76) <= not (a xor b);
    outputs(77) <= not (a xor b);
    outputs(78) <= not (a or b);
    outputs(79) <= not b;
    outputs(80) <= not a;
    outputs(81) <= b;
    outputs(82) <= a xor b;
    outputs(83) <= not (a or b);
    outputs(84) <= a;
    outputs(85) <= b;
    outputs(86) <= b and not a;
    outputs(87) <= a and not b;
    outputs(88) <= a;
    outputs(89) <= not a;
    outputs(90) <= not a;
    outputs(91) <= not (a xor b);
    outputs(92) <= a and b;
    outputs(93) <= not (a or b);
    outputs(94) <= a xor b;
    outputs(95) <= not (a or b);
    outputs(96) <= not a or b;
    outputs(97) <= not b;
    outputs(98) <= not (a xor b);
    outputs(99) <= not a;
    outputs(100) <= a or b;
    outputs(101) <= not b;
    outputs(102) <= a xor b;
    outputs(103) <= a;
    outputs(104) <= a xor b;
    outputs(105) <= a;
    outputs(106) <= not a;
    outputs(107) <= not (a or b);
    outputs(108) <= a xor b;
    outputs(109) <= not a;
    outputs(110) <= a xor b;
    outputs(111) <= not a;
    outputs(112) <= not b;
    outputs(113) <= b;
    outputs(114) <= a xor b;
    outputs(115) <= not (a xor b);
    outputs(116) <= not b;
    outputs(117) <= not b;
    outputs(118) <= a;
    outputs(119) <= a xor b;
    outputs(120) <= a;
    outputs(121) <= not (a xor b);
    outputs(122) <= not b;
    outputs(123) <= not a;
    outputs(124) <= a;
    outputs(125) <= not (a and b);
    outputs(126) <= not (a xor b);
    outputs(127) <= b;
    outputs(128) <= not (a xor b);
    outputs(129) <= a and not b;
    outputs(130) <= a xor b;
    outputs(131) <= b;
    outputs(132) <= b;
    outputs(133) <= not a;
    outputs(134) <= not b;
    outputs(135) <= not (a xor b);
    outputs(136) <= a xor b;
    outputs(137) <= b;
    outputs(138) <= a and b;
    outputs(139) <= not a;
    outputs(140) <= not (a xor b);
    outputs(141) <= not b;
    outputs(142) <= not b;
    outputs(143) <= not a or b;
    outputs(144) <= b;
    outputs(145) <= not (a xor b);
    outputs(146) <= a;
    outputs(147) <= a xor b;
    outputs(148) <= b;
    outputs(149) <= a;
    outputs(150) <= not a or b;
    outputs(151) <= not b;
    outputs(152) <= a;
    outputs(153) <= a;
    outputs(154) <= not a;
    outputs(155) <= not (a xor b);
    outputs(156) <= not (a xor b);
    outputs(157) <= a xor b;
    outputs(158) <= not a or b;
    outputs(159) <= b;
    outputs(160) <= not a or b;
    outputs(161) <= not a;
    outputs(162) <= b and not a;
    outputs(163) <= not (a xor b);
    outputs(164) <= not (a or b);
    outputs(165) <= not (a or b);
    outputs(166) <= not (a xor b);
    outputs(167) <= b;
    outputs(168) <= not (a or b);
    outputs(169) <= not a;
    outputs(170) <= a or b;
    outputs(171) <= a and b;
    outputs(172) <= not (a and b);
    outputs(173) <= b;
    outputs(174) <= not (a xor b);
    outputs(175) <= a or b;
    outputs(176) <= b;
    outputs(177) <= not a;
    outputs(178) <= not (a and b);
    outputs(179) <= a;
    outputs(180) <= not a;
    outputs(181) <= a;
    outputs(182) <= not (a xor b);
    outputs(183) <= b and not a;
    outputs(184) <= a;
    outputs(185) <= not a;
    outputs(186) <= a and not b;
    outputs(187) <= a xor b;
    outputs(188) <= a or b;
    outputs(189) <= a;
    outputs(190) <= b;
    outputs(191) <= not a;
    outputs(192) <= not (a xor b);
    outputs(193) <= b;
    outputs(194) <= b and not a;
    outputs(195) <= not (a or b);
    outputs(196) <= not a;
    outputs(197) <= a and not b;
    outputs(198) <= a xor b;
    outputs(199) <= b;
    outputs(200) <= not a or b;
    outputs(201) <= not (a xor b);
    outputs(202) <= a xor b;
    outputs(203) <= a and b;
    outputs(204) <= a;
    outputs(205) <= not (a or b);
    outputs(206) <= not b;
    outputs(207) <= not (a xor b);
    outputs(208) <= not a;
    outputs(209) <= a;
    outputs(210) <= not (a xor b);
    outputs(211) <= a xor b;
    outputs(212) <= '1';
    outputs(213) <= not b;
    outputs(214) <= not b or a;
    outputs(215) <= a or b;
    outputs(216) <= not (a xor b);
    outputs(217) <= not (a xor b);
    outputs(218) <= not (a xor b);
    outputs(219) <= not (a xor b);
    outputs(220) <= not (a xor b);
    outputs(221) <= a and not b;
    outputs(222) <= a xor b;
    outputs(223) <= not a;
    outputs(224) <= not (a xor b);
    outputs(225) <= a and b;
    outputs(226) <= a;
    outputs(227) <= a;
    outputs(228) <= b;
    outputs(229) <= a;
    outputs(230) <= a;
    outputs(231) <= not a;
    outputs(232) <= a xor b;
    outputs(233) <= not (a xor b);
    outputs(234) <= not (a xor b);
    outputs(235) <= not b;
    outputs(236) <= not b;
    outputs(237) <= a and not b;
    outputs(238) <= not a;
    outputs(239) <= a xor b;
    outputs(240) <= a;
    outputs(241) <= a xor b;
    outputs(242) <= not b;
    outputs(243) <= a;
    outputs(244) <= b;
    outputs(245) <= not a;
    outputs(246) <= not (a xor b);
    outputs(247) <= not b or a;
    outputs(248) <= a;
    outputs(249) <= not a;
    outputs(250) <= not b;
    outputs(251) <= not (a xor b);
    outputs(252) <= a;
    outputs(253) <= not b;
    outputs(254) <= a xor b;
    outputs(255) <= b;
    outputs(256) <= not a;
    outputs(257) <= b;
    outputs(258) <= a and not b;
    outputs(259) <= not (a xor b);
    outputs(260) <= a;
    outputs(261) <= a xor b;
    outputs(262) <= not a;
    outputs(263) <= b and not a;
    outputs(264) <= a;
    outputs(265) <= not b;
    outputs(266) <= a and not b;
    outputs(267) <= not (a xor b);
    outputs(268) <= not a;
    outputs(269) <= not a;
    outputs(270) <= a or b;
    outputs(271) <= not (a or b);
    outputs(272) <= a;
    outputs(273) <= b;
    outputs(274) <= not b;
    outputs(275) <= not a;
    outputs(276) <= not (a xor b);
    outputs(277) <= not a or b;
    outputs(278) <= a xor b;
    outputs(279) <= not a;
    outputs(280) <= not (a or b);
    outputs(281) <= a and b;
    outputs(282) <= a xor b;
    outputs(283) <= not (a xor b);
    outputs(284) <= b;
    outputs(285) <= b;
    outputs(286) <= not (a xor b);
    outputs(287) <= not b;
    outputs(288) <= not b;
    outputs(289) <= a xor b;
    outputs(290) <= b;
    outputs(291) <= a xor b;
    outputs(292) <= a xor b;
    outputs(293) <= a xor b;
    outputs(294) <= a xor b;
    outputs(295) <= not b or a;
    outputs(296) <= a or b;
    outputs(297) <= not b;
    outputs(298) <= a xor b;
    outputs(299) <= not b;
    outputs(300) <= a xor b;
    outputs(301) <= not a;
    outputs(302) <= not (a xor b);
    outputs(303) <= a;
    outputs(304) <= a xor b;
    outputs(305) <= a;
    outputs(306) <= not b;
    outputs(307) <= a and b;
    outputs(308) <= a xor b;
    outputs(309) <= not (a and b);
    outputs(310) <= a or b;
    outputs(311) <= a xor b;
    outputs(312) <= b and not a;
    outputs(313) <= a xor b;
    outputs(314) <= b;
    outputs(315) <= not (a xor b);
    outputs(316) <= not a;
    outputs(317) <= a;
    outputs(318) <= not (a xor b);
    outputs(319) <= not b or a;
    outputs(320) <= not b;
    outputs(321) <= b;
    outputs(322) <= a;
    outputs(323) <= not (a xor b);
    outputs(324) <= a xor b;
    outputs(325) <= not (a or b);
    outputs(326) <= not (a and b);
    outputs(327) <= not (a xor b);
    outputs(328) <= not b;
    outputs(329) <= a;
    outputs(330) <= a xor b;
    outputs(331) <= not (a xor b);
    outputs(332) <= a xor b;
    outputs(333) <= a;
    outputs(334) <= b;
    outputs(335) <= b;
    outputs(336) <= a xor b;
    outputs(337) <= a;
    outputs(338) <= a and not b;
    outputs(339) <= not (a xor b);
    outputs(340) <= a or b;
    outputs(341) <= a xor b;
    outputs(342) <= a and b;
    outputs(343) <= b and not a;
    outputs(344) <= b;
    outputs(345) <= not b;
    outputs(346) <= a;
    outputs(347) <= a and b;
    outputs(348) <= b;
    outputs(349) <= not (a and b);
    outputs(350) <= not a;
    outputs(351) <= not b or a;
    outputs(352) <= a;
    outputs(353) <= not a;
    outputs(354) <= a;
    outputs(355) <= not b;
    outputs(356) <= not (a xor b);
    outputs(357) <= b;
    outputs(358) <= b;
    outputs(359) <= b;
    outputs(360) <= not (a xor b);
    outputs(361) <= not b;
    outputs(362) <= not (a xor b);
    outputs(363) <= not b;
    outputs(364) <= not b or a;
    outputs(365) <= b;
    outputs(366) <= a or b;
    outputs(367) <= not b;
    outputs(368) <= not b;
    outputs(369) <= not (a xor b);
    outputs(370) <= b;
    outputs(371) <= not b;
    outputs(372) <= a and not b;
    outputs(373) <= not (a xor b);
    outputs(374) <= b;
    outputs(375) <= b and not a;
    outputs(376) <= not a;
    outputs(377) <= not (a xor b);
    outputs(378) <= not (a and b);
    outputs(379) <= b;
    outputs(380) <= b;
    outputs(381) <= a and b;
    outputs(382) <= not (a xor b);
    outputs(383) <= not b;
    outputs(384) <= not a;
    outputs(385) <= not (a xor b);
    outputs(386) <= not (a xor b);
    outputs(387) <= b;
    outputs(388) <= a xor b;
    outputs(389) <= a;
    outputs(390) <= not a;
    outputs(391) <= not b;
    outputs(392) <= a;
    outputs(393) <= not (a xor b);
    outputs(394) <= a;
    outputs(395) <= a and not b;
    outputs(396) <= a xor b;
    outputs(397) <= a and not b;
    outputs(398) <= not b;
    outputs(399) <= not b;
    outputs(400) <= not a;
    outputs(401) <= a;
    outputs(402) <= not a;
    outputs(403) <= b;
    outputs(404) <= a;
    outputs(405) <= not (a xor b);
    outputs(406) <= not (a xor b);
    outputs(407) <= not (a and b);
    outputs(408) <= not (a xor b);
    outputs(409) <= b;
    outputs(410) <= a xor b;
    outputs(411) <= not b or a;
    outputs(412) <= not (a xor b);
    outputs(413) <= a xor b;
    outputs(414) <= a;
    outputs(415) <= b;
    outputs(416) <= a xor b;
    outputs(417) <= b;
    outputs(418) <= a and b;
    outputs(419) <= not b;
    outputs(420) <= not (a or b);
    outputs(421) <= not (a or b);
    outputs(422) <= a xor b;
    outputs(423) <= b;
    outputs(424) <= a xor b;
    outputs(425) <= b;
    outputs(426) <= b;
    outputs(427) <= not a or b;
    outputs(428) <= a xor b;
    outputs(429) <= a xor b;
    outputs(430) <= not (a xor b);
    outputs(431) <= b;
    outputs(432) <= a;
    outputs(433) <= not a;
    outputs(434) <= not a;
    outputs(435) <= not (a xor b);
    outputs(436) <= b;
    outputs(437) <= not a;
    outputs(438) <= b;
    outputs(439) <= a;
    outputs(440) <= b;
    outputs(441) <= not (a and b);
    outputs(442) <= b;
    outputs(443) <= not a;
    outputs(444) <= b;
    outputs(445) <= not (a xor b);
    outputs(446) <= not a;
    outputs(447) <= a;
    outputs(448) <= a;
    outputs(449) <= not b;
    outputs(450) <= b and not a;
    outputs(451) <= not b or a;
    outputs(452) <= a;
    outputs(453) <= b;
    outputs(454) <= not a;
    outputs(455) <= not (a or b);
    outputs(456) <= not a;
    outputs(457) <= not b;
    outputs(458) <= a xor b;
    outputs(459) <= a;
    outputs(460) <= not a;
    outputs(461) <= not (a and b);
    outputs(462) <= b;
    outputs(463) <= not b;
    outputs(464) <= a or b;
    outputs(465) <= not (a xor b);
    outputs(466) <= a xor b;
    outputs(467) <= not b;
    outputs(468) <= not (a xor b);
    outputs(469) <= not b;
    outputs(470) <= not a;
    outputs(471) <= not b;
    outputs(472) <= a;
    outputs(473) <= not a;
    outputs(474) <= not a;
    outputs(475) <= a and not b;
    outputs(476) <= not b;
    outputs(477) <= b;
    outputs(478) <= not a;
    outputs(479) <= a xor b;
    outputs(480) <= b;
    outputs(481) <= a;
    outputs(482) <= a and b;
    outputs(483) <= a xor b;
    outputs(484) <= a;
    outputs(485) <= a;
    outputs(486) <= not (a xor b);
    outputs(487) <= b;
    outputs(488) <= a or b;
    outputs(489) <= a xor b;
    outputs(490) <= not b;
    outputs(491) <= not (a xor b);
    outputs(492) <= a xor b;
    outputs(493) <= a;
    outputs(494) <= not (a xor b);
    outputs(495) <= not (a xor b);
    outputs(496) <= a and not b;
    outputs(497) <= b;
    outputs(498) <= not b;
    outputs(499) <= a and not b;
    outputs(500) <= not (a xor b);
    outputs(501) <= not a;
    outputs(502) <= not (a or b);
    outputs(503) <= not (a xor b);
    outputs(504) <= not (a xor b);
    outputs(505) <= a;
    outputs(506) <= a xor b;
    outputs(507) <= b;
    outputs(508) <= not (a or b);
    outputs(509) <= not b or a;
    outputs(510) <= not a;
    outputs(511) <= not b;
    outputs(512) <= a and b;
    outputs(513) <= a and b;
    outputs(514) <= a or b;
    outputs(515) <= not (a xor b);
    outputs(516) <= b;
    outputs(517) <= not b;
    outputs(518) <= a xor b;
    outputs(519) <= not (a xor b);
    outputs(520) <= a;
    outputs(521) <= a xor b;
    outputs(522) <= not a;
    outputs(523) <= not (a or b);
    outputs(524) <= not (a xor b);
    outputs(525) <= not b;
    outputs(526) <= a and b;
    outputs(527) <= a and not b;
    outputs(528) <= a and b;
    outputs(529) <= b and not a;
    outputs(530) <= not (a xor b);
    outputs(531) <= a;
    outputs(532) <= a;
    outputs(533) <= a xor b;
    outputs(534) <= not a;
    outputs(535) <= b;
    outputs(536) <= b;
    outputs(537) <= a xor b;
    outputs(538) <= a and not b;
    outputs(539) <= not a;
    outputs(540) <= a;
    outputs(541) <= a xor b;
    outputs(542) <= not b;
    outputs(543) <= b;
    outputs(544) <= b and not a;
    outputs(545) <= not (a xor b);
    outputs(546) <= a and not b;
    outputs(547) <= b and not a;
    outputs(548) <= b;
    outputs(549) <= a xor b;
    outputs(550) <= a;
    outputs(551) <= b;
    outputs(552) <= b;
    outputs(553) <= not b;
    outputs(554) <= not b;
    outputs(555) <= not a;
    outputs(556) <= a;
    outputs(557) <= not b;
    outputs(558) <= not (a xor b);
    outputs(559) <= not a or b;
    outputs(560) <= not b;
    outputs(561) <= not b or a;
    outputs(562) <= a and not b;
    outputs(563) <= a;
    outputs(564) <= a;
    outputs(565) <= a xor b;
    outputs(566) <= not (a xor b);
    outputs(567) <= not b;
    outputs(568) <= a and b;
    outputs(569) <= not a;
    outputs(570) <= a;
    outputs(571) <= not a;
    outputs(572) <= a xor b;
    outputs(573) <= not b;
    outputs(574) <= not a;
    outputs(575) <= not a;
    outputs(576) <= b;
    outputs(577) <= a xor b;
    outputs(578) <= not (a or b);
    outputs(579) <= not (a xor b);
    outputs(580) <= b and not a;
    outputs(581) <= not (a and b);
    outputs(582) <= not a or b;
    outputs(583) <= not (a or b);
    outputs(584) <= not (a xor b);
    outputs(585) <= b;
    outputs(586) <= b;
    outputs(587) <= a xor b;
    outputs(588) <= not (a xor b);
    outputs(589) <= not a;
    outputs(590) <= b;
    outputs(591) <= b;
    outputs(592) <= not a;
    outputs(593) <= not b or a;
    outputs(594) <= not a;
    outputs(595) <= b and not a;
    outputs(596) <= a xor b;
    outputs(597) <= not (a or b);
    outputs(598) <= a xor b;
    outputs(599) <= a and b;
    outputs(600) <= not a;
    outputs(601) <= not (a xor b);
    outputs(602) <= not a;
    outputs(603) <= a xor b;
    outputs(604) <= not (a xor b);
    outputs(605) <= not (a xor b);
    outputs(606) <= a xor b;
    outputs(607) <= b;
    outputs(608) <= not (a and b);
    outputs(609) <= a xor b;
    outputs(610) <= b;
    outputs(611) <= b and not a;
    outputs(612) <= a and b;
    outputs(613) <= b;
    outputs(614) <= not (a and b);
    outputs(615) <= a and not b;
    outputs(616) <= a;
    outputs(617) <= not b;
    outputs(618) <= not (a xor b);
    outputs(619) <= not b;
    outputs(620) <= not a;
    outputs(621) <= a or b;
    outputs(622) <= a;
    outputs(623) <= not (a or b);
    outputs(624) <= a;
    outputs(625) <= not a;
    outputs(626) <= a;
    outputs(627) <= b and not a;
    outputs(628) <= not a;
    outputs(629) <= b;
    outputs(630) <= not b;
    outputs(631) <= a xor b;
    outputs(632) <= b;
    outputs(633) <= a xor b;
    outputs(634) <= b;
    outputs(635) <= b;
    outputs(636) <= not (a or b);
    outputs(637) <= not (a xor b);
    outputs(638) <= b and not a;
    outputs(639) <= a xor b;
    outputs(640) <= not b or a;
    outputs(641) <= a xor b;
    outputs(642) <= a xor b;
    outputs(643) <= not a;
    outputs(644) <= a xor b;
    outputs(645) <= a xor b;
    outputs(646) <= not b;
    outputs(647) <= not b;
    outputs(648) <= a xor b;
    outputs(649) <= not a;
    outputs(650) <= a;
    outputs(651) <= a and b;
    outputs(652) <= not a or b;
    outputs(653) <= a and not b;
    outputs(654) <= b;
    outputs(655) <= b;
    outputs(656) <= not (a xor b);
    outputs(657) <= not (a xor b);
    outputs(658) <= b and not a;
    outputs(659) <= a or b;
    outputs(660) <= not (a or b);
    outputs(661) <= not a;
    outputs(662) <= not b;
    outputs(663) <= not b;
    outputs(664) <= not (a xor b);
    outputs(665) <= a xor b;
    outputs(666) <= a xor b;
    outputs(667) <= a;
    outputs(668) <= a and b;
    outputs(669) <= a;
    outputs(670) <= b;
    outputs(671) <= a xor b;
    outputs(672) <= a xor b;
    outputs(673) <= a xor b;
    outputs(674) <= not a;
    outputs(675) <= b and not a;
    outputs(676) <= a or b;
    outputs(677) <= not b;
    outputs(678) <= a and not b;
    outputs(679) <= a xor b;
    outputs(680) <= b and not a;
    outputs(681) <= a and not b;
    outputs(682) <= b;
    outputs(683) <= not (a xor b);
    outputs(684) <= not b;
    outputs(685) <= not a;
    outputs(686) <= a xor b;
    outputs(687) <= not (a xor b);
    outputs(688) <= not (a and b);
    outputs(689) <= not b;
    outputs(690) <= a and not b;
    outputs(691) <= not b;
    outputs(692) <= not (a and b);
    outputs(693) <= not a;
    outputs(694) <= not b;
    outputs(695) <= not a;
    outputs(696) <= b and not a;
    outputs(697) <= not (a xor b);
    outputs(698) <= a xor b;
    outputs(699) <= a xor b;
    outputs(700) <= not a;
    outputs(701) <= not b;
    outputs(702) <= not b;
    outputs(703) <= not (a xor b);
    outputs(704) <= not b;
    outputs(705) <= not (a or b);
    outputs(706) <= a and b;
    outputs(707) <= not (a or b);
    outputs(708) <= not a;
    outputs(709) <= not (a xor b);
    outputs(710) <= not (a xor b);
    outputs(711) <= not a;
    outputs(712) <= not b;
    outputs(713) <= a;
    outputs(714) <= a and b;
    outputs(715) <= not (a xor b);
    outputs(716) <= b;
    outputs(717) <= not (a xor b);
    outputs(718) <= a;
    outputs(719) <= not b or a;
    outputs(720) <= a xor b;
    outputs(721) <= b and not a;
    outputs(722) <= not a;
    outputs(723) <= b;
    outputs(724) <= a xor b;
    outputs(725) <= a and b;
    outputs(726) <= a;
    outputs(727) <= a and b;
    outputs(728) <= not (a xor b);
    outputs(729) <= not a;
    outputs(730) <= a xor b;
    outputs(731) <= not a;
    outputs(732) <= not b;
    outputs(733) <= a xor b;
    outputs(734) <= not b or a;
    outputs(735) <= b;
    outputs(736) <= not a or b;
    outputs(737) <= a and b;
    outputs(738) <= a xor b;
    outputs(739) <= a xor b;
    outputs(740) <= not b;
    outputs(741) <= a;
    outputs(742) <= not (a xor b);
    outputs(743) <= a xor b;
    outputs(744) <= a and b;
    outputs(745) <= not a;
    outputs(746) <= b;
    outputs(747) <= a and b;
    outputs(748) <= a xor b;
    outputs(749) <= not b;
    outputs(750) <= b and not a;
    outputs(751) <= not (a or b);
    outputs(752) <= not (a xor b);
    outputs(753) <= b and not a;
    outputs(754) <= not a;
    outputs(755) <= not b;
    outputs(756) <= not b;
    outputs(757) <= a xor b;
    outputs(758) <= a xor b;
    outputs(759) <= a xor b;
    outputs(760) <= a and not b;
    outputs(761) <= not (a xor b);
    outputs(762) <= a xor b;
    outputs(763) <= not (a xor b);
    outputs(764) <= a;
    outputs(765) <= b;
    outputs(766) <= not (a xor b);
    outputs(767) <= b;
    outputs(768) <= b;
    outputs(769) <= not a;
    outputs(770) <= b;
    outputs(771) <= not b or a;
    outputs(772) <= b;
    outputs(773) <= not (a or b);
    outputs(774) <= a or b;
    outputs(775) <= not a or b;
    outputs(776) <= a xor b;
    outputs(777) <= b;
    outputs(778) <= not b;
    outputs(779) <= not b;
    outputs(780) <= a;
    outputs(781) <= b;
    outputs(782) <= a xor b;
    outputs(783) <= a xor b;
    outputs(784) <= b;
    outputs(785) <= a xor b;
    outputs(786) <= not a;
    outputs(787) <= b and not a;
    outputs(788) <= a xor b;
    outputs(789) <= a;
    outputs(790) <= b;
    outputs(791) <= not (a xor b);
    outputs(792) <= not a;
    outputs(793) <= a;
    outputs(794) <= b;
    outputs(795) <= a xor b;
    outputs(796) <= a xor b;
    outputs(797) <= b;
    outputs(798) <= not a;
    outputs(799) <= a;
    outputs(800) <= a;
    outputs(801) <= not b or a;
    outputs(802) <= b;
    outputs(803) <= not (a xor b);
    outputs(804) <= a;
    outputs(805) <= not a;
    outputs(806) <= a;
    outputs(807) <= a xor b;
    outputs(808) <= b and not a;
    outputs(809) <= not a;
    outputs(810) <= a;
    outputs(811) <= not b;
    outputs(812) <= a;
    outputs(813) <= a;
    outputs(814) <= not b;
    outputs(815) <= not (a xor b);
    outputs(816) <= a and not b;
    outputs(817) <= not b;
    outputs(818) <= not (a xor b);
    outputs(819) <= not a;
    outputs(820) <= b;
    outputs(821) <= a;
    outputs(822) <= not a;
    outputs(823) <= not b;
    outputs(824) <= not a;
    outputs(825) <= not a;
    outputs(826) <= a and not b;
    outputs(827) <= not b;
    outputs(828) <= not a;
    outputs(829) <= not b;
    outputs(830) <= not b;
    outputs(831) <= not (a xor b);
    outputs(832) <= a or b;
    outputs(833) <= not a;
    outputs(834) <= b;
    outputs(835) <= not a or b;
    outputs(836) <= a and not b;
    outputs(837) <= not a;
    outputs(838) <= a xor b;
    outputs(839) <= b;
    outputs(840) <= a and not b;
    outputs(841) <= not a;
    outputs(842) <= a;
    outputs(843) <= not (a xor b);
    outputs(844) <= not (a xor b);
    outputs(845) <= a;
    outputs(846) <= not a or b;
    outputs(847) <= a;
    outputs(848) <= a xor b;
    outputs(849) <= a;
    outputs(850) <= not (a or b);
    outputs(851) <= not b or a;
    outputs(852) <= not b or a;
    outputs(853) <= b and not a;
    outputs(854) <= b;
    outputs(855) <= not (a or b);
    outputs(856) <= not (a xor b);
    outputs(857) <= b and not a;
    outputs(858) <= a xor b;
    outputs(859) <= not (a xor b);
    outputs(860) <= not a;
    outputs(861) <= a xor b;
    outputs(862) <= not (a xor b);
    outputs(863) <= b and not a;
    outputs(864) <= a or b;
    outputs(865) <= not (a xor b);
    outputs(866) <= not b;
    outputs(867) <= not (a xor b);
    outputs(868) <= not b;
    outputs(869) <= not b;
    outputs(870) <= a and b;
    outputs(871) <= a;
    outputs(872) <= not a;
    outputs(873) <= b;
    outputs(874) <= b;
    outputs(875) <= a and b;
    outputs(876) <= not b or a;
    outputs(877) <= not (a xor b);
    outputs(878) <= a;
    outputs(879) <= not b;
    outputs(880) <= not a or b;
    outputs(881) <= a xor b;
    outputs(882) <= a;
    outputs(883) <= a xor b;
    outputs(884) <= not (a xor b);
    outputs(885) <= not a;
    outputs(886) <= b;
    outputs(887) <= a;
    outputs(888) <= not a;
    outputs(889) <= not b;
    outputs(890) <= a;
    outputs(891) <= a;
    outputs(892) <= not (a xor b);
    outputs(893) <= a;
    outputs(894) <= not b or a;
    outputs(895) <= not a;
    outputs(896) <= not (a xor b);
    outputs(897) <= a;
    outputs(898) <= not a;
    outputs(899) <= a xor b;
    outputs(900) <= b;
    outputs(901) <= a and not b;
    outputs(902) <= b;
    outputs(903) <= b;
    outputs(904) <= a xor b;
    outputs(905) <= a and b;
    outputs(906) <= a xor b;
    outputs(907) <= b;
    outputs(908) <= not (a and b);
    outputs(909) <= a;
    outputs(910) <= a xor b;
    outputs(911) <= b;
    outputs(912) <= not b;
    outputs(913) <= not a;
    outputs(914) <= not b;
    outputs(915) <= not b;
    outputs(916) <= a and b;
    outputs(917) <= a xor b;
    outputs(918) <= not a;
    outputs(919) <= not a;
    outputs(920) <= not b;
    outputs(921) <= a xor b;
    outputs(922) <= b;
    outputs(923) <= a and b;
    outputs(924) <= b;
    outputs(925) <= not b;
    outputs(926) <= not a;
    outputs(927) <= a xor b;
    outputs(928) <= a and b;
    outputs(929) <= not a;
    outputs(930) <= a;
    outputs(931) <= not b;
    outputs(932) <= a and b;
    outputs(933) <= a or b;
    outputs(934) <= not a;
    outputs(935) <= a xor b;
    outputs(936) <= not a;
    outputs(937) <= not b;
    outputs(938) <= not (a xor b);
    outputs(939) <= not (a or b);
    outputs(940) <= a xor b;
    outputs(941) <= a;
    outputs(942) <= a and b;
    outputs(943) <= not a;
    outputs(944) <= a xor b;
    outputs(945) <= a;
    outputs(946) <= a xor b;
    outputs(947) <= a;
    outputs(948) <= not (a xor b);
    outputs(949) <= not (a xor b);
    outputs(950) <= a and b;
    outputs(951) <= not (a and b);
    outputs(952) <= not (a or b);
    outputs(953) <= b and not a;
    outputs(954) <= b and not a;
    outputs(955) <= not b;
    outputs(956) <= not b;
    outputs(957) <= a;
    outputs(958) <= not b;
    outputs(959) <= not (a xor b);
    outputs(960) <= a and b;
    outputs(961) <= a;
    outputs(962) <= not b;
    outputs(963) <= a and not b;
    outputs(964) <= not b;
    outputs(965) <= not b;
    outputs(966) <= b and not a;
    outputs(967) <= a;
    outputs(968) <= not (a xor b);
    outputs(969) <= not (a xor b);
    outputs(970) <= b;
    outputs(971) <= a and b;
    outputs(972) <= b;
    outputs(973) <= not a;
    outputs(974) <= not a;
    outputs(975) <= a xor b;
    outputs(976) <= not b;
    outputs(977) <= not (a xor b);
    outputs(978) <= not (a xor b);
    outputs(979) <= not a;
    outputs(980) <= a and not b;
    outputs(981) <= not a;
    outputs(982) <= b and not a;
    outputs(983) <= not a;
    outputs(984) <= a;
    outputs(985) <= not (a and b);
    outputs(986) <= not a;
    outputs(987) <= not b;
    outputs(988) <= not b;
    outputs(989) <= a or b;
    outputs(990) <= a;
    outputs(991) <= b;
    outputs(992) <= a xor b;
    outputs(993) <= not (a xor b);
    outputs(994) <= not a;
    outputs(995) <= a;
    outputs(996) <= not a;
    outputs(997) <= a and b;
    outputs(998) <= b;
    outputs(999) <= a xor b;
    outputs(1000) <= a xor b;
    outputs(1001) <= b;
    outputs(1002) <= a xor b;
    outputs(1003) <= b;
    outputs(1004) <= not (a xor b);
    outputs(1005) <= not (a xor b);
    outputs(1006) <= not a;
    outputs(1007) <= not a;
    outputs(1008) <= not (a xor b);
    outputs(1009) <= a and not b;
    outputs(1010) <= not b;
    outputs(1011) <= a;
    outputs(1012) <= a xor b;
    outputs(1013) <= b;
    outputs(1014) <= not b;
    outputs(1015) <= not b;
    outputs(1016) <= a;
    outputs(1017) <= not b or a;
    outputs(1018) <= not (a xor b);
    outputs(1019) <= not a or b;
    outputs(1020) <= b;
    outputs(1021) <= not (a xor b);
    outputs(1022) <= not a;
    outputs(1023) <= not b;
    outputs(1024) <= b and not a;
    outputs(1025) <= not (a xor b);
    outputs(1026) <= b;
    outputs(1027) <= a xor b;
    outputs(1028) <= not a or b;
    outputs(1029) <= a xor b;
    outputs(1030) <= not (a xor b);
    outputs(1031) <= not b;
    outputs(1032) <= not (a or b);
    outputs(1033) <= a xor b;
    outputs(1034) <= a xor b;
    outputs(1035) <= not a;
    outputs(1036) <= a;
    outputs(1037) <= b and not a;
    outputs(1038) <= a xor b;
    outputs(1039) <= not (a or b);
    outputs(1040) <= not a;
    outputs(1041) <= a;
    outputs(1042) <= not a;
    outputs(1043) <= not b;
    outputs(1044) <= a xor b;
    outputs(1045) <= not (a xor b);
    outputs(1046) <= b and not a;
    outputs(1047) <= not (a xor b);
    outputs(1048) <= not (a xor b);
    outputs(1049) <= not (a xor b);
    outputs(1050) <= a xor b;
    outputs(1051) <= a and not b;
    outputs(1052) <= not b;
    outputs(1053) <= a xor b;
    outputs(1054) <= not a;
    outputs(1055) <= a;
    outputs(1056) <= b;
    outputs(1057) <= a and not b;
    outputs(1058) <= not a or b;
    outputs(1059) <= a xor b;
    outputs(1060) <= not b;
    outputs(1061) <= a xor b;
    outputs(1062) <= not (a or b);
    outputs(1063) <= a and not b;
    outputs(1064) <= not (a xor b);
    outputs(1065) <= a and not b;
    outputs(1066) <= not b;
    outputs(1067) <= not a;
    outputs(1068) <= not b;
    outputs(1069) <= not (a xor b);
    outputs(1070) <= not b or a;
    outputs(1071) <= a and not b;
    outputs(1072) <= not (a and b);
    outputs(1073) <= b;
    outputs(1074) <= not a;
    outputs(1075) <= not a;
    outputs(1076) <= not (a xor b);
    outputs(1077) <= not (a xor b);
    outputs(1078) <= a and b;
    outputs(1079) <= a;
    outputs(1080) <= not a;
    outputs(1081) <= not a;
    outputs(1082) <= not a;
    outputs(1083) <= a xor b;
    outputs(1084) <= not (a or b);
    outputs(1085) <= b and not a;
    outputs(1086) <= a;
    outputs(1087) <= not b;
    outputs(1088) <= not a;
    outputs(1089) <= a xor b;
    outputs(1090) <= a xor b;
    outputs(1091) <= not (a xor b);
    outputs(1092) <= not (a xor b);
    outputs(1093) <= not (a xor b);
    outputs(1094) <= b and not a;
    outputs(1095) <= not (a or b);
    outputs(1096) <= a xor b;
    outputs(1097) <= a;
    outputs(1098) <= a xor b;
    outputs(1099) <= not b;
    outputs(1100) <= b;
    outputs(1101) <= a and b;
    outputs(1102) <= a;
    outputs(1103) <= not (a xor b);
    outputs(1104) <= b;
    outputs(1105) <= not b;
    outputs(1106) <= a xor b;
    outputs(1107) <= a;
    outputs(1108) <= not b;
    outputs(1109) <= not a;
    outputs(1110) <= not (a xor b);
    outputs(1111) <= not (a or b);
    outputs(1112) <= not b;
    outputs(1113) <= a and b;
    outputs(1114) <= not b;
    outputs(1115) <= a xor b;
    outputs(1116) <= b and not a;
    outputs(1117) <= a;
    outputs(1118) <= a xor b;
    outputs(1119) <= not (a and b);
    outputs(1120) <= not (a xor b);
    outputs(1121) <= not b;
    outputs(1122) <= not (a or b);
    outputs(1123) <= a;
    outputs(1124) <= not (a xor b);
    outputs(1125) <= b;
    outputs(1126) <= b;
    outputs(1127) <= not (a or b);
    outputs(1128) <= not (a or b);
    outputs(1129) <= a xor b;
    outputs(1130) <= a;
    outputs(1131) <= a;
    outputs(1132) <= b and not a;
    outputs(1133) <= a;
    outputs(1134) <= not a;
    outputs(1135) <= a and not b;
    outputs(1136) <= a xor b;
    outputs(1137) <= not (a xor b);
    outputs(1138) <= not (a xor b);
    outputs(1139) <= a and b;
    outputs(1140) <= a and b;
    outputs(1141) <= not (a and b);
    outputs(1142) <= a xor b;
    outputs(1143) <= not (a xor b);
    outputs(1144) <= not b;
    outputs(1145) <= not a or b;
    outputs(1146) <= b;
    outputs(1147) <= not a;
    outputs(1148) <= not b;
    outputs(1149) <= not a;
    outputs(1150) <= a and not b;
    outputs(1151) <= not b;
    outputs(1152) <= b and not a;
    outputs(1153) <= not (a xor b);
    outputs(1154) <= not a;
    outputs(1155) <= a xor b;
    outputs(1156) <= not (a or b);
    outputs(1157) <= not a;
    outputs(1158) <= not (a xor b);
    outputs(1159) <= a;
    outputs(1160) <= not (a xor b);
    outputs(1161) <= not (a xor b);
    outputs(1162) <= a and b;
    outputs(1163) <= not a;
    outputs(1164) <= a xor b;
    outputs(1165) <= not b;
    outputs(1166) <= not a;
    outputs(1167) <= not (a xor b);
    outputs(1168) <= a;
    outputs(1169) <= not a;
    outputs(1170) <= b;
    outputs(1171) <= b and not a;
    outputs(1172) <= not a;
    outputs(1173) <= a xor b;
    outputs(1174) <= not a;
    outputs(1175) <= b and not a;
    outputs(1176) <= not (a xor b);
    outputs(1177) <= a xor b;
    outputs(1178) <= a xor b;
    outputs(1179) <= b;
    outputs(1180) <= a and b;
    outputs(1181) <= not b;
    outputs(1182) <= not a;
    outputs(1183) <= not a;
    outputs(1184) <= not a;
    outputs(1185) <= not (a xor b);
    outputs(1186) <= a xor b;
    outputs(1187) <= a;
    outputs(1188) <= not a;
    outputs(1189) <= a xor b;
    outputs(1190) <= b and not a;
    outputs(1191) <= not (a xor b);
    outputs(1192) <= a and b;
    outputs(1193) <= a;
    outputs(1194) <= not a;
    outputs(1195) <= not b;
    outputs(1196) <= not (a xor b);
    outputs(1197) <= not b or a;
    outputs(1198) <= b;
    outputs(1199) <= a;
    outputs(1200) <= a;
    outputs(1201) <= not a;
    outputs(1202) <= not a;
    outputs(1203) <= a;
    outputs(1204) <= a xor b;
    outputs(1205) <= not (a xor b);
    outputs(1206) <= a xor b;
    outputs(1207) <= not (a xor b);
    outputs(1208) <= b;
    outputs(1209) <= not a;
    outputs(1210) <= a;
    outputs(1211) <= not (a xor b);
    outputs(1212) <= b;
    outputs(1213) <= not b;
    outputs(1214) <= not a;
    outputs(1215) <= not b;
    outputs(1216) <= a xor b;
    outputs(1217) <= a and b;
    outputs(1218) <= not (a and b);
    outputs(1219) <= not b;
    outputs(1220) <= a xor b;
    outputs(1221) <= not (a xor b);
    outputs(1222) <= a and not b;
    outputs(1223) <= a;
    outputs(1224) <= not a or b;
    outputs(1225) <= not a;
    outputs(1226) <= not (a xor b);
    outputs(1227) <= not a;
    outputs(1228) <= not b;
    outputs(1229) <= b;
    outputs(1230) <= a;
    outputs(1231) <= not (a xor b);
    outputs(1232) <= not a;
    outputs(1233) <= not a;
    outputs(1234) <= a xor b;
    outputs(1235) <= not (a xor b);
    outputs(1236) <= b;
    outputs(1237) <= b;
    outputs(1238) <= b;
    outputs(1239) <= a;
    outputs(1240) <= not b;
    outputs(1241) <= a xor b;
    outputs(1242) <= b;
    outputs(1243) <= not (a xor b);
    outputs(1244) <= a xor b;
    outputs(1245) <= a xor b;
    outputs(1246) <= b;
    outputs(1247) <= b;
    outputs(1248) <= a and not b;
    outputs(1249) <= not (a xor b);
    outputs(1250) <= not (a xor b);
    outputs(1251) <= a xor b;
    outputs(1252) <= a;
    outputs(1253) <= not a or b;
    outputs(1254) <= b and not a;
    outputs(1255) <= a;
    outputs(1256) <= a or b;
    outputs(1257) <= not b;
    outputs(1258) <= not (a xor b);
    outputs(1259) <= a xor b;
    outputs(1260) <= not (a or b);
    outputs(1261) <= a;
    outputs(1262) <= a xor b;
    outputs(1263) <= a xor b;
    outputs(1264) <= not a;
    outputs(1265) <= not (a xor b);
    outputs(1266) <= not a;
    outputs(1267) <= not b or a;
    outputs(1268) <= not a;
    outputs(1269) <= a xor b;
    outputs(1270) <= b and not a;
    outputs(1271) <= not a;
    outputs(1272) <= not a;
    outputs(1273) <= not b;
    outputs(1274) <= a xor b;
    outputs(1275) <= not b;
    outputs(1276) <= not a or b;
    outputs(1277) <= not (a xor b);
    outputs(1278) <= not a;
    outputs(1279) <= not a;
    outputs(1280) <= not (a xor b);
    outputs(1281) <= a xor b;
    outputs(1282) <= not (a xor b);
    outputs(1283) <= b and not a;
    outputs(1284) <= b and not a;
    outputs(1285) <= not (a xor b);
    outputs(1286) <= a and b;
    outputs(1287) <= not (a xor b);
    outputs(1288) <= not a;
    outputs(1289) <= not b;
    outputs(1290) <= not (a xor b);
    outputs(1291) <= a xor b;
    outputs(1292) <= a xor b;
    outputs(1293) <= not a;
    outputs(1294) <= a xor b;
    outputs(1295) <= a xor b;
    outputs(1296) <= b;
    outputs(1297) <= b;
    outputs(1298) <= b;
    outputs(1299) <= a and b;
    outputs(1300) <= a;
    outputs(1301) <= not a;
    outputs(1302) <= a and not b;
    outputs(1303) <= '0';
    outputs(1304) <= not a or b;
    outputs(1305) <= not a;
    outputs(1306) <= b and not a;
    outputs(1307) <= a xor b;
    outputs(1308) <= b and not a;
    outputs(1309) <= a xor b;
    outputs(1310) <= a;
    outputs(1311) <= '0';
    outputs(1312) <= not b;
    outputs(1313) <= a xor b;
    outputs(1314) <= not (a xor b);
    outputs(1315) <= not (a xor b);
    outputs(1316) <= a;
    outputs(1317) <= not (a xor b);
    outputs(1318) <= not a;
    outputs(1319) <= not b or a;
    outputs(1320) <= not (a xor b);
    outputs(1321) <= a and b;
    outputs(1322) <= not (a xor b);
    outputs(1323) <= a;
    outputs(1324) <= b and not a;
    outputs(1325) <= a;
    outputs(1326) <= b;
    outputs(1327) <= not (a xor b);
    outputs(1328) <= a xor b;
    outputs(1329) <= b and not a;
    outputs(1330) <= b and not a;
    outputs(1331) <= a and not b;
    outputs(1332) <= a xor b;
    outputs(1333) <= b;
    outputs(1334) <= not (a xor b);
    outputs(1335) <= not b;
    outputs(1336) <= a xor b;
    outputs(1337) <= b;
    outputs(1338) <= not (a xor b);
    outputs(1339) <= not (a xor b);
    outputs(1340) <= a;
    outputs(1341) <= not (a xor b);
    outputs(1342) <= b;
    outputs(1343) <= b and not a;
    outputs(1344) <= a and b;
    outputs(1345) <= a xor b;
    outputs(1346) <= a and not b;
    outputs(1347) <= a;
    outputs(1348) <= a xor b;
    outputs(1349) <= a xor b;
    outputs(1350) <= a and b;
    outputs(1351) <= not (a xor b);
    outputs(1352) <= not b;
    outputs(1353) <= a xor b;
    outputs(1354) <= not b;
    outputs(1355) <= a and b;
    outputs(1356) <= not a;
    outputs(1357) <= not (a xor b);
    outputs(1358) <= not b;
    outputs(1359) <= a xor b;
    outputs(1360) <= b and not a;
    outputs(1361) <= a xor b;
    outputs(1362) <= a;
    outputs(1363) <= not b;
    outputs(1364) <= not a;
    outputs(1365) <= b;
    outputs(1366) <= not a;
    outputs(1367) <= not a;
    outputs(1368) <= a;
    outputs(1369) <= a or b;
    outputs(1370) <= a and not b;
    outputs(1371) <= not (a xor b);
    outputs(1372) <= a;
    outputs(1373) <= not (a or b);
    outputs(1374) <= not (a xor b);
    outputs(1375) <= not (a or b);
    outputs(1376) <= not b;
    outputs(1377) <= a;
    outputs(1378) <= b;
    outputs(1379) <= a xor b;
    outputs(1380) <= a xor b;
    outputs(1381) <= b;
    outputs(1382) <= a or b;
    outputs(1383) <= a;
    outputs(1384) <= a;
    outputs(1385) <= not (a xor b);
    outputs(1386) <= b;
    outputs(1387) <= not a or b;
    outputs(1388) <= not a;
    outputs(1389) <= not a;
    outputs(1390) <= a xor b;
    outputs(1391) <= not (a xor b);
    outputs(1392) <= not b;
    outputs(1393) <= a;
    outputs(1394) <= b;
    outputs(1395) <= not a or b;
    outputs(1396) <= not a;
    outputs(1397) <= a xor b;
    outputs(1398) <= a and b;
    outputs(1399) <= not (a xor b);
    outputs(1400) <= not a;
    outputs(1401) <= a;
    outputs(1402) <= not b;
    outputs(1403) <= b and not a;
    outputs(1404) <= a xor b;
    outputs(1405) <= not (a xor b);
    outputs(1406) <= a;
    outputs(1407) <= not b;
    outputs(1408) <= not a;
    outputs(1409) <= not (a xor b);
    outputs(1410) <= b;
    outputs(1411) <= a;
    outputs(1412) <= a and not b;
    outputs(1413) <= b;
    outputs(1414) <= b;
    outputs(1415) <= b;
    outputs(1416) <= not (a xor b);
    outputs(1417) <= a and not b;
    outputs(1418) <= not (a xor b);
    outputs(1419) <= b;
    outputs(1420) <= a xor b;
    outputs(1421) <= a;
    outputs(1422) <= a;
    outputs(1423) <= a and b;
    outputs(1424) <= a xor b;
    outputs(1425) <= not b;
    outputs(1426) <= not (a or b);
    outputs(1427) <= a;
    outputs(1428) <= not (a or b);
    outputs(1429) <= not a;
    outputs(1430) <= a and b;
    outputs(1431) <= a xor b;
    outputs(1432) <= a xor b;
    outputs(1433) <= a or b;
    outputs(1434) <= not (a or b);
    outputs(1435) <= b;
    outputs(1436) <= b and not a;
    outputs(1437) <= not a;
    outputs(1438) <= not (a xor b);
    outputs(1439) <= not (a xor b);
    outputs(1440) <= b;
    outputs(1441) <= b and not a;
    outputs(1442) <= a xor b;
    outputs(1443) <= a;
    outputs(1444) <= a and not b;
    outputs(1445) <= a xor b;
    outputs(1446) <= not (a xor b);
    outputs(1447) <= not b;
    outputs(1448) <= not (a xor b);
    outputs(1449) <= not a or b;
    outputs(1450) <= not b;
    outputs(1451) <= not (a xor b);
    outputs(1452) <= a xor b;
    outputs(1453) <= not (a xor b);
    outputs(1454) <= not b;
    outputs(1455) <= not (a xor b);
    outputs(1456) <= not (a xor b);
    outputs(1457) <= a or b;
    outputs(1458) <= b and not a;
    outputs(1459) <= a;
    outputs(1460) <= not (a xor b);
    outputs(1461) <= not b;
    outputs(1462) <= a xor b;
    outputs(1463) <= a;
    outputs(1464) <= not (a xor b);
    outputs(1465) <= a and not b;
    outputs(1466) <= not a;
    outputs(1467) <= a xor b;
    outputs(1468) <= not a;
    outputs(1469) <= a;
    outputs(1470) <= not (a or b);
    outputs(1471) <= a xor b;
    outputs(1472) <= a;
    outputs(1473) <= not (a xor b);
    outputs(1474) <= a xor b;
    outputs(1475) <= a xor b;
    outputs(1476) <= not (a xor b);
    outputs(1477) <= b;
    outputs(1478) <= a and b;
    outputs(1479) <= not b;
    outputs(1480) <= not a;
    outputs(1481) <= a xor b;
    outputs(1482) <= not (a and b);
    outputs(1483) <= not a;
    outputs(1484) <= b;
    outputs(1485) <= '0';
    outputs(1486) <= not (a xor b);
    outputs(1487) <= b;
    outputs(1488) <= b;
    outputs(1489) <= not (a or b);
    outputs(1490) <= a xor b;
    outputs(1491) <= a and b;
    outputs(1492) <= not a;
    outputs(1493) <= not (a xor b);
    outputs(1494) <= not b;
    outputs(1495) <= a xor b;
    outputs(1496) <= a xor b;
    outputs(1497) <= a;
    outputs(1498) <= not b;
    outputs(1499) <= not b;
    outputs(1500) <= not a;
    outputs(1501) <= a and not b;
    outputs(1502) <= not b;
    outputs(1503) <= not (a or b);
    outputs(1504) <= a xor b;
    outputs(1505) <= not a;
    outputs(1506) <= not a;
    outputs(1507) <= not b;
    outputs(1508) <= a xor b;
    outputs(1509) <= not (a xor b);
    outputs(1510) <= a and not b;
    outputs(1511) <= a and b;
    outputs(1512) <= b;
    outputs(1513) <= a xor b;
    outputs(1514) <= not b;
    outputs(1515) <= not b;
    outputs(1516) <= b and not a;
    outputs(1517) <= a xor b;
    outputs(1518) <= a and b;
    outputs(1519) <= b and not a;
    outputs(1520) <= b and not a;
    outputs(1521) <= a;
    outputs(1522) <= a xor b;
    outputs(1523) <= a;
    outputs(1524) <= not (a or b);
    outputs(1525) <= b;
    outputs(1526) <= not (a xor b);
    outputs(1527) <= not b or a;
    outputs(1528) <= not b;
    outputs(1529) <= a xor b;
    outputs(1530) <= not (a or b);
    outputs(1531) <= b;
    outputs(1532) <= b and not a;
    outputs(1533) <= a and b;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= not (a xor b);
    outputs(1536) <= a;
    outputs(1537) <= not b;
    outputs(1538) <= not (a or b);
    outputs(1539) <= not b;
    outputs(1540) <= not (a or b);
    outputs(1541) <= a xor b;
    outputs(1542) <= a and b;
    outputs(1543) <= b;
    outputs(1544) <= b;
    outputs(1545) <= not (a or b);
    outputs(1546) <= not (a and b);
    outputs(1547) <= not a;
    outputs(1548) <= a;
    outputs(1549) <= not b;
    outputs(1550) <= a xor b;
    outputs(1551) <= not (a xor b);
    outputs(1552) <= not (a xor b);
    outputs(1553) <= not (a or b);
    outputs(1554) <= not a;
    outputs(1555) <= not (a xor b);
    outputs(1556) <= not a;
    outputs(1557) <= b;
    outputs(1558) <= b;
    outputs(1559) <= a xor b;
    outputs(1560) <= a;
    outputs(1561) <= not (a xor b);
    outputs(1562) <= a and b;
    outputs(1563) <= a and not b;
    outputs(1564) <= not a;
    outputs(1565) <= not a;
    outputs(1566) <= not b;
    outputs(1567) <= not (a xor b);
    outputs(1568) <= not (a or b);
    outputs(1569) <= not a;
    outputs(1570) <= not a;
    outputs(1571) <= a and b;
    outputs(1572) <= b;
    outputs(1573) <= a xor b;
    outputs(1574) <= a xor b;
    outputs(1575) <= not a;
    outputs(1576) <= a xor b;
    outputs(1577) <= a xor b;
    outputs(1578) <= not b;
    outputs(1579) <= a and b;
    outputs(1580) <= not (a and b);
    outputs(1581) <= a xor b;
    outputs(1582) <= not (a xor b);
    outputs(1583) <= not (a xor b);
    outputs(1584) <= not (a and b);
    outputs(1585) <= a or b;
    outputs(1586) <= b and not a;
    outputs(1587) <= not a;
    outputs(1588) <= a;
    outputs(1589) <= not a;
    outputs(1590) <= a;
    outputs(1591) <= b;
    outputs(1592) <= not b;
    outputs(1593) <= not a;
    outputs(1594) <= not b;
    outputs(1595) <= not b;
    outputs(1596) <= a xor b;
    outputs(1597) <= a and b;
    outputs(1598) <= a and not b;
    outputs(1599) <= a and b;
    outputs(1600) <= a;
    outputs(1601) <= a and not b;
    outputs(1602) <= not (a xor b);
    outputs(1603) <= a xor b;
    outputs(1604) <= a xor b;
    outputs(1605) <= not (a xor b);
    outputs(1606) <= a and b;
    outputs(1607) <= not b;
    outputs(1608) <= a xor b;
    outputs(1609) <= a xor b;
    outputs(1610) <= a xor b;
    outputs(1611) <= a and b;
    outputs(1612) <= not b;
    outputs(1613) <= b;
    outputs(1614) <= b;
    outputs(1615) <= a xor b;
    outputs(1616) <= a xor b;
    outputs(1617) <= b;
    outputs(1618) <= a xor b;
    outputs(1619) <= a;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= a xor b;
    outputs(1622) <= b;
    outputs(1623) <= b;
    outputs(1624) <= a and b;
    outputs(1625) <= a xor b;
    outputs(1626) <= b;
    outputs(1627) <= not b;
    outputs(1628) <= not (a xor b);
    outputs(1629) <= a xor b;
    outputs(1630) <= b;
    outputs(1631) <= a and b;
    outputs(1632) <= b and not a;
    outputs(1633) <= b;
    outputs(1634) <= not b;
    outputs(1635) <= not (a and b);
    outputs(1636) <= not a;
    outputs(1637) <= a xor b;
    outputs(1638) <= b;
    outputs(1639) <= not a;
    outputs(1640) <= a and b;
    outputs(1641) <= not a;
    outputs(1642) <= a xor b;
    outputs(1643) <= not (a xor b);
    outputs(1644) <= not b;
    outputs(1645) <= a and b;
    outputs(1646) <= a and not b;
    outputs(1647) <= not (a xor b);
    outputs(1648) <= not (a xor b);
    outputs(1649) <= a and b;
    outputs(1650) <= not a;
    outputs(1651) <= not (a xor b);
    outputs(1652) <= not (a xor b);
    outputs(1653) <= b;
    outputs(1654) <= b;
    outputs(1655) <= a and not b;
    outputs(1656) <= not (a xor b);
    outputs(1657) <= not (a or b);
    outputs(1658) <= b;
    outputs(1659) <= a xor b;
    outputs(1660) <= not a;
    outputs(1661) <= not (a and b);
    outputs(1662) <= not (a xor b);
    outputs(1663) <= a xor b;
    outputs(1664) <= not b;
    outputs(1665) <= not (a xor b);
    outputs(1666) <= a;
    outputs(1667) <= a xor b;
    outputs(1668) <= not b;
    outputs(1669) <= not (a or b);
    outputs(1670) <= a;
    outputs(1671) <= not b or a;
    outputs(1672) <= not (a xor b);
    outputs(1673) <= b;
    outputs(1674) <= a and b;
    outputs(1675) <= a and b;
    outputs(1676) <= not a;
    outputs(1677) <= a;
    outputs(1678) <= not (a or b);
    outputs(1679) <= not (a xor b);
    outputs(1680) <= a;
    outputs(1681) <= a;
    outputs(1682) <= a and not b;
    outputs(1683) <= not (a xor b);
    outputs(1684) <= not (a xor b);
    outputs(1685) <= a;
    outputs(1686) <= a;
    outputs(1687) <= a;
    outputs(1688) <= not a;
    outputs(1689) <= not a;
    outputs(1690) <= b;
    outputs(1691) <= a;
    outputs(1692) <= not b;
    outputs(1693) <= not (a xor b);
    outputs(1694) <= not (a and b);
    outputs(1695) <= not a;
    outputs(1696) <= a xor b;
    outputs(1697) <= not b;
    outputs(1698) <= a xor b;
    outputs(1699) <= not (a xor b);
    outputs(1700) <= not b;
    outputs(1701) <= not a;
    outputs(1702) <= not a;
    outputs(1703) <= not (a xor b);
    outputs(1704) <= not b;
    outputs(1705) <= a;
    outputs(1706) <= a and b;
    outputs(1707) <= not a;
    outputs(1708) <= b;
    outputs(1709) <= not b;
    outputs(1710) <= a xor b;
    outputs(1711) <= a xor b;
    outputs(1712) <= a xor b;
    outputs(1713) <= a xor b;
    outputs(1714) <= a;
    outputs(1715) <= not (a xor b);
    outputs(1716) <= not (a or b);
    outputs(1717) <= b;
    outputs(1718) <= b and not a;
    outputs(1719) <= not (a xor b);
    outputs(1720) <= not a;
    outputs(1721) <= a and not b;
    outputs(1722) <= b and not a;
    outputs(1723) <= b;
    outputs(1724) <= not (a xor b);
    outputs(1725) <= not (a xor b);
    outputs(1726) <= a and not b;
    outputs(1727) <= not (a xor b);
    outputs(1728) <= not a;
    outputs(1729) <= a xor b;
    outputs(1730) <= not (a xor b);
    outputs(1731) <= not (a xor b);
    outputs(1732) <= b;
    outputs(1733) <= not (a xor b);
    outputs(1734) <= a xor b;
    outputs(1735) <= not (a xor b);
    outputs(1736) <= not (a or b);
    outputs(1737) <= b;
    outputs(1738) <= not b;
    outputs(1739) <= not (a xor b);
    outputs(1740) <= b;
    outputs(1741) <= a xor b;
    outputs(1742) <= not (a xor b);
    outputs(1743) <= not a;
    outputs(1744) <= a;
    outputs(1745) <= a xor b;
    outputs(1746) <= not b;
    outputs(1747) <= a xor b;
    outputs(1748) <= b;
    outputs(1749) <= a and b;
    outputs(1750) <= b;
    outputs(1751) <= not a;
    outputs(1752) <= a;
    outputs(1753) <= a;
    outputs(1754) <= not a;
    outputs(1755) <= a;
    outputs(1756) <= a;
    outputs(1757) <= a xor b;
    outputs(1758) <= a xor b;
    outputs(1759) <= not b or a;
    outputs(1760) <= not b;
    outputs(1761) <= a and not b;
    outputs(1762) <= a;
    outputs(1763) <= a and not b;
    outputs(1764) <= a;
    outputs(1765) <= b;
    outputs(1766) <= b and not a;
    outputs(1767) <= not (a xor b);
    outputs(1768) <= a xor b;
    outputs(1769) <= not (a xor b);
    outputs(1770) <= a xor b;
    outputs(1771) <= not (a xor b);
    outputs(1772) <= a;
    outputs(1773) <= b and not a;
    outputs(1774) <= b;
    outputs(1775) <= not (a xor b);
    outputs(1776) <= not (a xor b);
    outputs(1777) <= not (a or b);
    outputs(1778) <= b;
    outputs(1779) <= not (a xor b);
    outputs(1780) <= a;
    outputs(1781) <= b;
    outputs(1782) <= b and not a;
    outputs(1783) <= a;
    outputs(1784) <= not (a or b);
    outputs(1785) <= not b;
    outputs(1786) <= not a;
    outputs(1787) <= not (a xor b);
    outputs(1788) <= not (a xor b);
    outputs(1789) <= b and not a;
    outputs(1790) <= a xor b;
    outputs(1791) <= b;
    outputs(1792) <= b and not a;
    outputs(1793) <= not b;
    outputs(1794) <= a;
    outputs(1795) <= not a;
    outputs(1796) <= a;
    outputs(1797) <= a;
    outputs(1798) <= '0';
    outputs(1799) <= a;
    outputs(1800) <= not a;
    outputs(1801) <= b;
    outputs(1802) <= a xor b;
    outputs(1803) <= b and not a;
    outputs(1804) <= not b;
    outputs(1805) <= not a;
    outputs(1806) <= not (a xor b);
    outputs(1807) <= not (a xor b);
    outputs(1808) <= a and b;
    outputs(1809) <= not b;
    outputs(1810) <= not a;
    outputs(1811) <= b and not a;
    outputs(1812) <= not (a xor b);
    outputs(1813) <= not (a xor b);
    outputs(1814) <= a xor b;
    outputs(1815) <= a;
    outputs(1816) <= a xor b;
    outputs(1817) <= not (a xor b);
    outputs(1818) <= not (a xor b);
    outputs(1819) <= a xor b;
    outputs(1820) <= not a;
    outputs(1821) <= a xor b;
    outputs(1822) <= a and not b;
    outputs(1823) <= not (a xor b);
    outputs(1824) <= not (a or b);
    outputs(1825) <= not b;
    outputs(1826) <= not b;
    outputs(1827) <= b;
    outputs(1828) <= b and not a;
    outputs(1829) <= a and b;
    outputs(1830) <= not a;
    outputs(1831) <= not (a xor b);
    outputs(1832) <= a xor b;
    outputs(1833) <= a;
    outputs(1834) <= a xor b;
    outputs(1835) <= a;
    outputs(1836) <= a xor b;
    outputs(1837) <= not (a xor b);
    outputs(1838) <= not b;
    outputs(1839) <= a xor b;
    outputs(1840) <= b and not a;
    outputs(1841) <= a xor b;
    outputs(1842) <= not (a xor b);
    outputs(1843) <= a xor b;
    outputs(1844) <= a and not b;
    outputs(1845) <= not (a xor b);
    outputs(1846) <= not (a xor b);
    outputs(1847) <= not b;
    outputs(1848) <= a and not b;
    outputs(1849) <= a and b;
    outputs(1850) <= a xor b;
    outputs(1851) <= not (a xor b);
    outputs(1852) <= a xor b;
    outputs(1853) <= b and not a;
    outputs(1854) <= not (a xor b);
    outputs(1855) <= not (a xor b);
    outputs(1856) <= not a or b;
    outputs(1857) <= not b;
    outputs(1858) <= not b;
    outputs(1859) <= not b;
    outputs(1860) <= not (a xor b);
    outputs(1861) <= not (a and b);
    outputs(1862) <= not (a xor b);
    outputs(1863) <= a;
    outputs(1864) <= not b;
    outputs(1865) <= a xor b;
    outputs(1866) <= a and b;
    outputs(1867) <= not a;
    outputs(1868) <= a xor b;
    outputs(1869) <= a;
    outputs(1870) <= a;
    outputs(1871) <= not a;
    outputs(1872) <= '0';
    outputs(1873) <= not a;
    outputs(1874) <= a;
    outputs(1875) <= a;
    outputs(1876) <= not b;
    outputs(1877) <= b;
    outputs(1878) <= a and b;
    outputs(1879) <= not (a and b);
    outputs(1880) <= a and b;
    outputs(1881) <= not (a xor b);
    outputs(1882) <= a xor b;
    outputs(1883) <= not a or b;
    outputs(1884) <= not b;
    outputs(1885) <= not (a xor b);
    outputs(1886) <= a;
    outputs(1887) <= a or b;
    outputs(1888) <= a xor b;
    outputs(1889) <= a;
    outputs(1890) <= not a;
    outputs(1891) <= a xor b;
    outputs(1892) <= a and not b;
    outputs(1893) <= a xor b;
    outputs(1894) <= a xor b;
    outputs(1895) <= a;
    outputs(1896) <= not (a xor b);
    outputs(1897) <= b and not a;
    outputs(1898) <= not b;
    outputs(1899) <= not a;
    outputs(1900) <= a xor b;
    outputs(1901) <= not b or a;
    outputs(1902) <= b and not a;
    outputs(1903) <= a xor b;
    outputs(1904) <= b;
    outputs(1905) <= a xor b;
    outputs(1906) <= not (a xor b);
    outputs(1907) <= a and b;
    outputs(1908) <= a xor b;
    outputs(1909) <= a xor b;
    outputs(1910) <= a xor b;
    outputs(1911) <= not b;
    outputs(1912) <= not (a or b);
    outputs(1913) <= a xor b;
    outputs(1914) <= b and not a;
    outputs(1915) <= not b;
    outputs(1916) <= not (a xor b);
    outputs(1917) <= a and not b;
    outputs(1918) <= a and b;
    outputs(1919) <= a and not b;
    outputs(1920) <= not a;
    outputs(1921) <= b and not a;
    outputs(1922) <= not (a or b);
    outputs(1923) <= not a;
    outputs(1924) <= a;
    outputs(1925) <= not b;
    outputs(1926) <= a xor b;
    outputs(1927) <= b and not a;
    outputs(1928) <= a and b;
    outputs(1929) <= b;
    outputs(1930) <= not (a xor b);
    outputs(1931) <= not b;
    outputs(1932) <= a xor b;
    outputs(1933) <= a and not b;
    outputs(1934) <= a;
    outputs(1935) <= b;
    outputs(1936) <= a;
    outputs(1937) <= a;
    outputs(1938) <= b;
    outputs(1939) <= not b;
    outputs(1940) <= not (a xor b);
    outputs(1941) <= not (a xor b);
    outputs(1942) <= a and b;
    outputs(1943) <= b;
    outputs(1944) <= not b;
    outputs(1945) <= a xor b;
    outputs(1946) <= not (a xor b);
    outputs(1947) <= b;
    outputs(1948) <= not (a xor b);
    outputs(1949) <= a;
    outputs(1950) <= a;
    outputs(1951) <= b and not a;
    outputs(1952) <= not (a xor b);
    outputs(1953) <= not a;
    outputs(1954) <= not a;
    outputs(1955) <= b;
    outputs(1956) <= a xor b;
    outputs(1957) <= a and not b;
    outputs(1958) <= not (a xor b);
    outputs(1959) <= b;
    outputs(1960) <= a and not b;
    outputs(1961) <= a;
    outputs(1962) <= not a;
    outputs(1963) <= not (a xor b);
    outputs(1964) <= a;
    outputs(1965) <= a xor b;
    outputs(1966) <= b and not a;
    outputs(1967) <= a and not b;
    outputs(1968) <= b;
    outputs(1969) <= not b;
    outputs(1970) <= not (a or b);
    outputs(1971) <= not a;
    outputs(1972) <= not b;
    outputs(1973) <= not a;
    outputs(1974) <= not (a xor b);
    outputs(1975) <= a and b;
    outputs(1976) <= a;
    outputs(1977) <= a;
    outputs(1978) <= not a;
    outputs(1979) <= a and b;
    outputs(1980) <= not (a xor b);
    outputs(1981) <= not (a xor b);
    outputs(1982) <= not a;
    outputs(1983) <= not (a xor b);
    outputs(1984) <= not (a xor b);
    outputs(1985) <= a xor b;
    outputs(1986) <= not (a xor b);
    outputs(1987) <= not b;
    outputs(1988) <= b;
    outputs(1989) <= a xor b;
    outputs(1990) <= a or b;
    outputs(1991) <= not b;
    outputs(1992) <= a and b;
    outputs(1993) <= not (a xor b);
    outputs(1994) <= not (a and b);
    outputs(1995) <= not b;
    outputs(1996) <= a and not b;
    outputs(1997) <= b;
    outputs(1998) <= a and b;
    outputs(1999) <= a and not b;
    outputs(2000) <= not a;
    outputs(2001) <= not (a xor b);
    outputs(2002) <= not b;
    outputs(2003) <= a xor b;
    outputs(2004) <= b;
    outputs(2005) <= not a;
    outputs(2006) <= not a;
    outputs(2007) <= a xor b;
    outputs(2008) <= not b;
    outputs(2009) <= a xor b;
    outputs(2010) <= a and b;
    outputs(2011) <= a xor b;
    outputs(2012) <= a and not b;
    outputs(2013) <= not b;
    outputs(2014) <= not a or b;
    outputs(2015) <= a;
    outputs(2016) <= a;
    outputs(2017) <= not b or a;
    outputs(2018) <= not b;
    outputs(2019) <= b and not a;
    outputs(2020) <= not a;
    outputs(2021) <= not a;
    outputs(2022) <= b;
    outputs(2023) <= not (a xor b);
    outputs(2024) <= a and not b;
    outputs(2025) <= a xor b;
    outputs(2026) <= a xor b;
    outputs(2027) <= a;
    outputs(2028) <= b and not a;
    outputs(2029) <= b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= a xor b;
    outputs(2032) <= not b;
    outputs(2033) <= b and not a;
    outputs(2034) <= a xor b;
    outputs(2035) <= a and not b;
    outputs(2036) <= not (a xor b);
    outputs(2037) <= b;
    outputs(2038) <= a or b;
    outputs(2039) <= not a;
    outputs(2040) <= a or b;
    outputs(2041) <= a and not b;
    outputs(2042) <= b and not a;
    outputs(2043) <= a xor b;
    outputs(2044) <= not (a xor b);
    outputs(2045) <= b and not a;
    outputs(2046) <= not b or a;
    outputs(2047) <= '0';
    outputs(2048) <= not (a and b);
    outputs(2049) <= not (a xor b);
    outputs(2050) <= a xor b;
    outputs(2051) <= not (a xor b);
    outputs(2052) <= not (a xor b);
    outputs(2053) <= a xor b;
    outputs(2054) <= b;
    outputs(2055) <= not (a xor b);
    outputs(2056) <= not b;
    outputs(2057) <= not (a xor b);
    outputs(2058) <= a and b;
    outputs(2059) <= a xor b;
    outputs(2060) <= not a;
    outputs(2061) <= not b;
    outputs(2062) <= not (a xor b);
    outputs(2063) <= a;
    outputs(2064) <= not (a xor b);
    outputs(2065) <= a xor b;
    outputs(2066) <= a;
    outputs(2067) <= a;
    outputs(2068) <= not a;
    outputs(2069) <= b;
    outputs(2070) <= not (a xor b);
    outputs(2071) <= b;
    outputs(2072) <= not a;
    outputs(2073) <= a and b;
    outputs(2074) <= a and b;
    outputs(2075) <= not a or b;
    outputs(2076) <= a and not b;
    outputs(2077) <= a or b;
    outputs(2078) <= a xor b;
    outputs(2079) <= a;
    outputs(2080) <= a;
    outputs(2081) <= not a;
    outputs(2082) <= not (a or b);
    outputs(2083) <= a xor b;
    outputs(2084) <= not b;
    outputs(2085) <= a and b;
    outputs(2086) <= a xor b;
    outputs(2087) <= a xor b;
    outputs(2088) <= not b;
    outputs(2089) <= not b or a;
    outputs(2090) <= a;
    outputs(2091) <= a xor b;
    outputs(2092) <= not (a xor b);
    outputs(2093) <= a xor b;
    outputs(2094) <= a and not b;
    outputs(2095) <= not (a xor b);
    outputs(2096) <= a;
    outputs(2097) <= not b;
    outputs(2098) <= a xor b;
    outputs(2099) <= a;
    outputs(2100) <= a xor b;
    outputs(2101) <= not (a xor b);
    outputs(2102) <= a and not b;
    outputs(2103) <= a;
    outputs(2104) <= not a;
    outputs(2105) <= not b;
    outputs(2106) <= not b;
    outputs(2107) <= not (a xor b);
    outputs(2108) <= not (a xor b);
    outputs(2109) <= not b;
    outputs(2110) <= a xor b;
    outputs(2111) <= not (a xor b);
    outputs(2112) <= not (a xor b);
    outputs(2113) <= a and b;
    outputs(2114) <= a and b;
    outputs(2115) <= a and not b;
    outputs(2116) <= b;
    outputs(2117) <= not (a xor b);
    outputs(2118) <= a;
    outputs(2119) <= a xor b;
    outputs(2120) <= not a;
    outputs(2121) <= b and not a;
    outputs(2122) <= b;
    outputs(2123) <= a and not b;
    outputs(2124) <= not (a xor b);
    outputs(2125) <= a xor b;
    outputs(2126) <= a;
    outputs(2127) <= not (a xor b);
    outputs(2128) <= not (a or b);
    outputs(2129) <= not b or a;
    outputs(2130) <= not a;
    outputs(2131) <= b;
    outputs(2132) <= a;
    outputs(2133) <= not (a xor b);
    outputs(2134) <= b;
    outputs(2135) <= a;
    outputs(2136) <= not a;
    outputs(2137) <= not a;
    outputs(2138) <= a;
    outputs(2139) <= b;
    outputs(2140) <= a and b;
    outputs(2141) <= not b or a;
    outputs(2142) <= not (a xor b);
    outputs(2143) <= not (a xor b);
    outputs(2144) <= not a;
    outputs(2145) <= not (a xor b);
    outputs(2146) <= a xor b;
    outputs(2147) <= not a;
    outputs(2148) <= b;
    outputs(2149) <= a;
    outputs(2150) <= b;
    outputs(2151) <= not b;
    outputs(2152) <= a xor b;
    outputs(2153) <= a and b;
    outputs(2154) <= b;
    outputs(2155) <= a xor b;
    outputs(2156) <= not (a xor b);
    outputs(2157) <= not (a xor b);
    outputs(2158) <= not b;
    outputs(2159) <= not (a xor b);
    outputs(2160) <= not (a xor b);
    outputs(2161) <= a xor b;
    outputs(2162) <= b;
    outputs(2163) <= a xor b;
    outputs(2164) <= not b;
    outputs(2165) <= b;
    outputs(2166) <= b and not a;
    outputs(2167) <= not a;
    outputs(2168) <= a xor b;
    outputs(2169) <= b and not a;
    outputs(2170) <= b;
    outputs(2171) <= a xor b;
    outputs(2172) <= a and not b;
    outputs(2173) <= a and b;
    outputs(2174) <= not (a xor b);
    outputs(2175) <= a;
    outputs(2176) <= a xor b;
    outputs(2177) <= a xor b;
    outputs(2178) <= not a;
    outputs(2179) <= b;
    outputs(2180) <= b and not a;
    outputs(2181) <= b;
    outputs(2182) <= a xor b;
    outputs(2183) <= a xor b;
    outputs(2184) <= not b or a;
    outputs(2185) <= not b;
    outputs(2186) <= a xor b;
    outputs(2187) <= b;
    outputs(2188) <= not a;
    outputs(2189) <= not (a xor b);
    outputs(2190) <= a xor b;
    outputs(2191) <= not (a xor b);
    outputs(2192) <= not (a or b);
    outputs(2193) <= a and not b;
    outputs(2194) <= a and b;
    outputs(2195) <= not a;
    outputs(2196) <= not (a xor b);
    outputs(2197) <= not b;
    outputs(2198) <= not (a or b);
    outputs(2199) <= a xor b;
    outputs(2200) <= a;
    outputs(2201) <= not (a xor b);
    outputs(2202) <= not (a or b);
    outputs(2203) <= not (a or b);
    outputs(2204) <= not (a xor b);
    outputs(2205) <= a;
    outputs(2206) <= not (a xor b);
    outputs(2207) <= not a;
    outputs(2208) <= b and not a;
    outputs(2209) <= b;
    outputs(2210) <= not b;
    outputs(2211) <= b;
    outputs(2212) <= a and b;
    outputs(2213) <= not (a xor b);
    outputs(2214) <= not (a xor b);
    outputs(2215) <= not b;
    outputs(2216) <= a xor b;
    outputs(2217) <= a and not b;
    outputs(2218) <= not (a and b);
    outputs(2219) <= a xor b;
    outputs(2220) <= not a;
    outputs(2221) <= b;
    outputs(2222) <= b and not a;
    outputs(2223) <= a and not b;
    outputs(2224) <= b and not a;
    outputs(2225) <= not b;
    outputs(2226) <= a xor b;
    outputs(2227) <= not a;
    outputs(2228) <= not (a xor b);
    outputs(2229) <= a xor b;
    outputs(2230) <= not a;
    outputs(2231) <= not (a xor b);
    outputs(2232) <= a and not b;
    outputs(2233) <= b;
    outputs(2234) <= b;
    outputs(2235) <= not b or a;
    outputs(2236) <= a xor b;
    outputs(2237) <= a xor b;
    outputs(2238) <= a;
    outputs(2239) <= a xor b;
    outputs(2240) <= not b;
    outputs(2241) <= b;
    outputs(2242) <= b and not a;
    outputs(2243) <= b;
    outputs(2244) <= not (a xor b);
    outputs(2245) <= not a;
    outputs(2246) <= a xor b;
    outputs(2247) <= not (a xor b);
    outputs(2248) <= not (a xor b);
    outputs(2249) <= a xor b;
    outputs(2250) <= a xor b;
    outputs(2251) <= a and b;
    outputs(2252) <= a xor b;
    outputs(2253) <= not a;
    outputs(2254) <= b;
    outputs(2255) <= a xor b;
    outputs(2256) <= not a;
    outputs(2257) <= a and not b;
    outputs(2258) <= a and b;
    outputs(2259) <= a xor b;
    outputs(2260) <= b;
    outputs(2261) <= a or b;
    outputs(2262) <= not (a xor b);
    outputs(2263) <= not b;
    outputs(2264) <= not b;
    outputs(2265) <= a xor b;
    outputs(2266) <= not a;
    outputs(2267) <= not b;
    outputs(2268) <= not (a and b);
    outputs(2269) <= not (a xor b);
    outputs(2270) <= not (a xor b);
    outputs(2271) <= not b;
    outputs(2272) <= not a;
    outputs(2273) <= b and not a;
    outputs(2274) <= a xor b;
    outputs(2275) <= a and b;
    outputs(2276) <= not (a or b);
    outputs(2277) <= not (a xor b);
    outputs(2278) <= not (a xor b);
    outputs(2279) <= not (a xor b);
    outputs(2280) <= not a;
    outputs(2281) <= a and b;
    outputs(2282) <= not a;
    outputs(2283) <= b and not a;
    outputs(2284) <= not (a or b);
    outputs(2285) <= b;
    outputs(2286) <= not b;
    outputs(2287) <= not b;
    outputs(2288) <= a xor b;
    outputs(2289) <= a xor b;
    outputs(2290) <= not b;
    outputs(2291) <= a;
    outputs(2292) <= not b;
    outputs(2293) <= a and not b;
    outputs(2294) <= a xor b;
    outputs(2295) <= a xor b;
    outputs(2296) <= a and not b;
    outputs(2297) <= not (a xor b);
    outputs(2298) <= a xor b;
    outputs(2299) <= b;
    outputs(2300) <= a xor b;
    outputs(2301) <= a;
    outputs(2302) <= a;
    outputs(2303) <= a xor b;
    outputs(2304) <= a and b;
    outputs(2305) <= a xor b;
    outputs(2306) <= a xor b;
    outputs(2307) <= b;
    outputs(2308) <= not a;
    outputs(2309) <= not b;
    outputs(2310) <= b;
    outputs(2311) <= not a;
    outputs(2312) <= not b;
    outputs(2313) <= a and b;
    outputs(2314) <= not b;
    outputs(2315) <= b and not a;
    outputs(2316) <= a and not b;
    outputs(2317) <= b;
    outputs(2318) <= not (a xor b);
    outputs(2319) <= not b;
    outputs(2320) <= not a;
    outputs(2321) <= a;
    outputs(2322) <= not (a xor b);
    outputs(2323) <= b and not a;
    outputs(2324) <= b;
    outputs(2325) <= not (a xor b);
    outputs(2326) <= not (a or b);
    outputs(2327) <= not (a xor b);
    outputs(2328) <= a xor b;
    outputs(2329) <= a;
    outputs(2330) <= a and b;
    outputs(2331) <= not (a or b);
    outputs(2332) <= b and not a;
    outputs(2333) <= not b;
    outputs(2334) <= a xor b;
    outputs(2335) <= not b;
    outputs(2336) <= a;
    outputs(2337) <= not (a or b);
    outputs(2338) <= a xor b;
    outputs(2339) <= not b;
    outputs(2340) <= not (a xor b);
    outputs(2341) <= a xor b;
    outputs(2342) <= not (a or b);
    outputs(2343) <= b and not a;
    outputs(2344) <= a;
    outputs(2345) <= a xor b;
    outputs(2346) <= not (a xor b);
    outputs(2347) <= a and b;
    outputs(2348) <= not a;
    outputs(2349) <= not (a xor b);
    outputs(2350) <= b;
    outputs(2351) <= a and b;
    outputs(2352) <= a and b;
    outputs(2353) <= b and not a;
    outputs(2354) <= not a;
    outputs(2355) <= a;
    outputs(2356) <= a xor b;
    outputs(2357) <= a and b;
    outputs(2358) <= b and not a;
    outputs(2359) <= not (a xor b);
    outputs(2360) <= b;
    outputs(2361) <= a xor b;
    outputs(2362) <= a and not b;
    outputs(2363) <= a xor b;
    outputs(2364) <= not (a xor b);
    outputs(2365) <= not a or b;
    outputs(2366) <= a;
    outputs(2367) <= not b or a;
    outputs(2368) <= a and b;
    outputs(2369) <= a xor b;
    outputs(2370) <= a and not b;
    outputs(2371) <= not a;
    outputs(2372) <= a;
    outputs(2373) <= a xor b;
    outputs(2374) <= not b;
    outputs(2375) <= b;
    outputs(2376) <= b;
    outputs(2377) <= not (a or b);
    outputs(2378) <= b;
    outputs(2379) <= not (a xor b);
    outputs(2380) <= not b;
    outputs(2381) <= b;
    outputs(2382) <= a and not b;
    outputs(2383) <= not (a xor b);
    outputs(2384) <= not b;
    outputs(2385) <= b;
    outputs(2386) <= b;
    outputs(2387) <= a xor b;
    outputs(2388) <= a;
    outputs(2389) <= not (a and b);
    outputs(2390) <= b;
    outputs(2391) <= a and not b;
    outputs(2392) <= b;
    outputs(2393) <= not (a xor b);
    outputs(2394) <= a;
    outputs(2395) <= not a;
    outputs(2396) <= a xor b;
    outputs(2397) <= b;
    outputs(2398) <= not (a xor b);
    outputs(2399) <= a and not b;
    outputs(2400) <= a xor b;
    outputs(2401) <= not a or b;
    outputs(2402) <= not (a xor b);
    outputs(2403) <= a xor b;
    outputs(2404) <= not (a or b);
    outputs(2405) <= a and not b;
    outputs(2406) <= not a;
    outputs(2407) <= not (a xor b);
    outputs(2408) <= not (a xor b);
    outputs(2409) <= a xor b;
    outputs(2410) <= a xor b;
    outputs(2411) <= a xor b;
    outputs(2412) <= not (a xor b);
    outputs(2413) <= b;
    outputs(2414) <= a xor b;
    outputs(2415) <= not a;
    outputs(2416) <= not b;
    outputs(2417) <= a xor b;
    outputs(2418) <= a;
    outputs(2419) <= a and b;
    outputs(2420) <= a xor b;
    outputs(2421) <= not b;
    outputs(2422) <= not (a xor b);
    outputs(2423) <= not b;
    outputs(2424) <= a or b;
    outputs(2425) <= a and b;
    outputs(2426) <= b and not a;
    outputs(2427) <= not (a xor b);
    outputs(2428) <= not (a and b);
    outputs(2429) <= a and b;
    outputs(2430) <= a xor b;
    outputs(2431) <= not (a xor b);
    outputs(2432) <= a;
    outputs(2433) <= a and not b;
    outputs(2434) <= not (a xor b);
    outputs(2435) <= b and not a;
    outputs(2436) <= b;
    outputs(2437) <= not b;
    outputs(2438) <= not (a xor b);
    outputs(2439) <= not b;
    outputs(2440) <= not (a or b);
    outputs(2441) <= a xor b;
    outputs(2442) <= b;
    outputs(2443) <= not (a xor b);
    outputs(2444) <= a;
    outputs(2445) <= a;
    outputs(2446) <= b and not a;
    outputs(2447) <= not (a xor b);
    outputs(2448) <= not a;
    outputs(2449) <= not (a xor b);
    outputs(2450) <= a xor b;
    outputs(2451) <= not (a xor b);
    outputs(2452) <= not (a or b);
    outputs(2453) <= b;
    outputs(2454) <= not b;
    outputs(2455) <= not a or b;
    outputs(2456) <= not (a xor b);
    outputs(2457) <= not (a xor b);
    outputs(2458) <= b and not a;
    outputs(2459) <= a xor b;
    outputs(2460) <= a and not b;
    outputs(2461) <= not (a xor b);
    outputs(2462) <= a xor b;
    outputs(2463) <= not b;
    outputs(2464) <= not a;
    outputs(2465) <= b;
    outputs(2466) <= a;
    outputs(2467) <= not (a xor b);
    outputs(2468) <= not a;
    outputs(2469) <= not (a xor b);
    outputs(2470) <= not (a xor b);
    outputs(2471) <= a and not b;
    outputs(2472) <= b;
    outputs(2473) <= not b;
    outputs(2474) <= not (a xor b);
    outputs(2475) <= a and b;
    outputs(2476) <= not (a xor b);
    outputs(2477) <= a xor b;
    outputs(2478) <= a xor b;
    outputs(2479) <= a xor b;
    outputs(2480) <= a;
    outputs(2481) <= not (a xor b);
    outputs(2482) <= not a;
    outputs(2483) <= a xor b;
    outputs(2484) <= b and not a;
    outputs(2485) <= not a;
    outputs(2486) <= b;
    outputs(2487) <= not (a xor b);
    outputs(2488) <= a;
    outputs(2489) <= a xor b;
    outputs(2490) <= not (a xor b);
    outputs(2491) <= not (a xor b);
    outputs(2492) <= not b;
    outputs(2493) <= b;
    outputs(2494) <= a xor b;
    outputs(2495) <= a;
    outputs(2496) <= b;
    outputs(2497) <= b;
    outputs(2498) <= not (a xor b);
    outputs(2499) <= a xor b;
    outputs(2500) <= a and b;
    outputs(2501) <= a;
    outputs(2502) <= b and not a;
    outputs(2503) <= not (a xor b);
    outputs(2504) <= not (a xor b);
    outputs(2505) <= a xor b;
    outputs(2506) <= a;
    outputs(2507) <= not (a or b);
    outputs(2508) <= not (a xor b);
    outputs(2509) <= a;
    outputs(2510) <= a and b;
    outputs(2511) <= a;
    outputs(2512) <= b and not a;
    outputs(2513) <= not (a or b);
    outputs(2514) <= b;
    outputs(2515) <= not (a xor b);
    outputs(2516) <= not b;
    outputs(2517) <= not (a or b);
    outputs(2518) <= not a;
    outputs(2519) <= not a or b;
    outputs(2520) <= not (a xor b);
    outputs(2521) <= not b;
    outputs(2522) <= b;
    outputs(2523) <= not (a or b);
    outputs(2524) <= a and not b;
    outputs(2525) <= not a;
    outputs(2526) <= not (a xor b);
    outputs(2527) <= not a;
    outputs(2528) <= a xor b;
    outputs(2529) <= a and b;
    outputs(2530) <= a and b;
    outputs(2531) <= not (a xor b);
    outputs(2532) <= not (a or b);
    outputs(2533) <= not a;
    outputs(2534) <= a xor b;
    outputs(2535) <= b;
    outputs(2536) <= a and b;
    outputs(2537) <= b and not a;
    outputs(2538) <= not a;
    outputs(2539) <= not a or b;
    outputs(2540) <= not (a or b);
    outputs(2541) <= a xor b;
    outputs(2542) <= b;
    outputs(2543) <= not b;
    outputs(2544) <= b and not a;
    outputs(2545) <= not a;
    outputs(2546) <= not b;
    outputs(2547) <= not (a and b);
    outputs(2548) <= a;
    outputs(2549) <= not (a xor b);
    outputs(2550) <= b and not a;
    outputs(2551) <= a and not b;
    outputs(2552) <= a and b;
    outputs(2553) <= a and not b;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= a and not b;
    outputs(2556) <= a and not b;
    outputs(2557) <= b;
    outputs(2558) <= not a;
    outputs(2559) <= not (a xor b);
    outputs(2560) <= b;
    outputs(2561) <= a;
    outputs(2562) <= not (a xor b);
    outputs(2563) <= not (a and b);
    outputs(2564) <= not b;
    outputs(2565) <= a xor b;
    outputs(2566) <= a;
    outputs(2567) <= not b;
    outputs(2568) <= a xor b;
    outputs(2569) <= a xor b;
    outputs(2570) <= not (a xor b);
    outputs(2571) <= not a or b;
    outputs(2572) <= a;
    outputs(2573) <= a;
    outputs(2574) <= b;
    outputs(2575) <= not a;
    outputs(2576) <= b;
    outputs(2577) <= not b;
    outputs(2578) <= b;
    outputs(2579) <= not a;
    outputs(2580) <= a;
    outputs(2581) <= a xor b;
    outputs(2582) <= b;
    outputs(2583) <= not (a xor b);
    outputs(2584) <= a and b;
    outputs(2585) <= b;
    outputs(2586) <= not (a xor b);
    outputs(2587) <= not (a xor b);
    outputs(2588) <= a xor b;
    outputs(2589) <= a or b;
    outputs(2590) <= a xor b;
    outputs(2591) <= not a;
    outputs(2592) <= not (a or b);
    outputs(2593) <= not a;
    outputs(2594) <= not b;
    outputs(2595) <= a and not b;
    outputs(2596) <= b;
    outputs(2597) <= not (a xor b);
    outputs(2598) <= b;
    outputs(2599) <= b and not a;
    outputs(2600) <= a xor b;
    outputs(2601) <= not (a xor b);
    outputs(2602) <= b;
    outputs(2603) <= a;
    outputs(2604) <= not b;
    outputs(2605) <= not a;
    outputs(2606) <= a and not b;
    outputs(2607) <= b;
    outputs(2608) <= b;
    outputs(2609) <= not (a or b);
    outputs(2610) <= not a;
    outputs(2611) <= not a;
    outputs(2612) <= a xor b;
    outputs(2613) <= not (a xor b);
    outputs(2614) <= a xor b;
    outputs(2615) <= not a;
    outputs(2616) <= not a;
    outputs(2617) <= not b;
    outputs(2618) <= a;
    outputs(2619) <= b;
    outputs(2620) <= a xor b;
    outputs(2621) <= not a;
    outputs(2622) <= not (a and b);
    outputs(2623) <= not (a xor b);
    outputs(2624) <= not b;
    outputs(2625) <= not a;
    outputs(2626) <= not b;
    outputs(2627) <= not (a xor b);
    outputs(2628) <= b;
    outputs(2629) <= a;
    outputs(2630) <= a and not b;
    outputs(2631) <= not b;
    outputs(2632) <= not b;
    outputs(2633) <= not a;
    outputs(2634) <= a and b;
    outputs(2635) <= a xor b;
    outputs(2636) <= a and b;
    outputs(2637) <= b and not a;
    outputs(2638) <= a;
    outputs(2639) <= a or b;
    outputs(2640) <= not b;
    outputs(2641) <= not a;
    outputs(2642) <= a xor b;
    outputs(2643) <= not b or a;
    outputs(2644) <= not (a or b);
    outputs(2645) <= a;
    outputs(2646) <= a xor b;
    outputs(2647) <= not (a xor b);
    outputs(2648) <= a xor b;
    outputs(2649) <= not a;
    outputs(2650) <= not (a or b);
    outputs(2651) <= not a;
    outputs(2652) <= a xor b;
    outputs(2653) <= not (a xor b);
    outputs(2654) <= b;
    outputs(2655) <= a;
    outputs(2656) <= not b;
    outputs(2657) <= not a;
    outputs(2658) <= a xor b;
    outputs(2659) <= not (a xor b);
    outputs(2660) <= not (a or b);
    outputs(2661) <= not a;
    outputs(2662) <= a;
    outputs(2663) <= not (a or b);
    outputs(2664) <= not (a and b);
    outputs(2665) <= b;
    outputs(2666) <= not (a xor b);
    outputs(2667) <= a;
    outputs(2668) <= a xor b;
    outputs(2669) <= not a;
    outputs(2670) <= a xor b;
    outputs(2671) <= a xor b;
    outputs(2672) <= a xor b;
    outputs(2673) <= not b;
    outputs(2674) <= a xor b;
    outputs(2675) <= not a;
    outputs(2676) <= not b;
    outputs(2677) <= a xor b;
    outputs(2678) <= a xor b;
    outputs(2679) <= not a;
    outputs(2680) <= not b;
    outputs(2681) <= not b or a;
    outputs(2682) <= not (a and b);
    outputs(2683) <= not a;
    outputs(2684) <= not a;
    outputs(2685) <= not (a xor b);
    outputs(2686) <= not (a or b);
    outputs(2687) <= not (a xor b);
    outputs(2688) <= a xor b;
    outputs(2689) <= a xor b;
    outputs(2690) <= not b or a;
    outputs(2691) <= not a;
    outputs(2692) <= a;
    outputs(2693) <= not b;
    outputs(2694) <= not (a and b);
    outputs(2695) <= not (a xor b);
    outputs(2696) <= a;
    outputs(2697) <= a xor b;
    outputs(2698) <= not b;
    outputs(2699) <= not b;
    outputs(2700) <= a xor b;
    outputs(2701) <= a;
    outputs(2702) <= b;
    outputs(2703) <= not a or b;
    outputs(2704) <= a xor b;
    outputs(2705) <= b;
    outputs(2706) <= not b or a;
    outputs(2707) <= b;
    outputs(2708) <= a;
    outputs(2709) <= a;
    outputs(2710) <= a;
    outputs(2711) <= not b or a;
    outputs(2712) <= not (a xor b);
    outputs(2713) <= not b;
    outputs(2714) <= b;
    outputs(2715) <= not (a or b);
    outputs(2716) <= not a;
    outputs(2717) <= not (a xor b);
    outputs(2718) <= not (a xor b);
    outputs(2719) <= not (a xor b);
    outputs(2720) <= a xor b;
    outputs(2721) <= a and b;
    outputs(2722) <= not (a or b);
    outputs(2723) <= not (a and b);
    outputs(2724) <= not a;
    outputs(2725) <= a;
    outputs(2726) <= not b;
    outputs(2727) <= not (a xor b);
    outputs(2728) <= not (a xor b);
    outputs(2729) <= not (a and b);
    outputs(2730) <= not (a and b);
    outputs(2731) <= a and b;
    outputs(2732) <= a xor b;
    outputs(2733) <= not b;
    outputs(2734) <= a;
    outputs(2735) <= not (a xor b);
    outputs(2736) <= not (a xor b);
    outputs(2737) <= a xor b;
    outputs(2738) <= a xor b;
    outputs(2739) <= b and not a;
    outputs(2740) <= a;
    outputs(2741) <= not a;
    outputs(2742) <= not (a xor b);
    outputs(2743) <= a xor b;
    outputs(2744) <= not (a or b);
    outputs(2745) <= a and not b;
    outputs(2746) <= not (a or b);
    outputs(2747) <= not b or a;
    outputs(2748) <= not b;
    outputs(2749) <= b;
    outputs(2750) <= not (a xor b);
    outputs(2751) <= not (a xor b);
    outputs(2752) <= a;
    outputs(2753) <= not (a xor b);
    outputs(2754) <= not (a xor b);
    outputs(2755) <= not a;
    outputs(2756) <= a;
    outputs(2757) <= b;
    outputs(2758) <= a;
    outputs(2759) <= a xor b;
    outputs(2760) <= not (a xor b);
    outputs(2761) <= not b;
    outputs(2762) <= b;
    outputs(2763) <= not (a and b);
    outputs(2764) <= not (a xor b);
    outputs(2765) <= not a;
    outputs(2766) <= a xor b;
    outputs(2767) <= b;
    outputs(2768) <= a xor b;
    outputs(2769) <= a xor b;
    outputs(2770) <= not a;
    outputs(2771) <= a xor b;
    outputs(2772) <= b;
    outputs(2773) <= not (a or b);
    outputs(2774) <= not (a xor b);
    outputs(2775) <= not b;
    outputs(2776) <= a xor b;
    outputs(2777) <= not (a xor b);
    outputs(2778) <= a;
    outputs(2779) <= not b;
    outputs(2780) <= a xor b;
    outputs(2781) <= not (a xor b);
    outputs(2782) <= b and not a;
    outputs(2783) <= not b;
    outputs(2784) <= a;
    outputs(2785) <= a xor b;
    outputs(2786) <= a and not b;
    outputs(2787) <= not a;
    outputs(2788) <= a;
    outputs(2789) <= a;
    outputs(2790) <= not b;
    outputs(2791) <= not a;
    outputs(2792) <= a xor b;
    outputs(2793) <= a;
    outputs(2794) <= not b;
    outputs(2795) <= a and b;
    outputs(2796) <= a;
    outputs(2797) <= not a or b;
    outputs(2798) <= a xor b;
    outputs(2799) <= a;
    outputs(2800) <= a;
    outputs(2801) <= a xor b;
    outputs(2802) <= b;
    outputs(2803) <= not (a xor b);
    outputs(2804) <= a xor b;
    outputs(2805) <= a xor b;
    outputs(2806) <= a xor b;
    outputs(2807) <= not a;
    outputs(2808) <= not (a xor b);
    outputs(2809) <= not (a xor b);
    outputs(2810) <= not (a xor b);
    outputs(2811) <= not (a xor b);
    outputs(2812) <= a xor b;
    outputs(2813) <= not (a xor b);
    outputs(2814) <= not b or a;
    outputs(2815) <= b;
    outputs(2816) <= a xor b;
    outputs(2817) <= a xor b;
    outputs(2818) <= a;
    outputs(2819) <= not b;
    outputs(2820) <= not b;
    outputs(2821) <= a xor b;
    outputs(2822) <= a;
    outputs(2823) <= a;
    outputs(2824) <= not (a or b);
    outputs(2825) <= not (a xor b);
    outputs(2826) <= not (a xor b);
    outputs(2827) <= not b or a;
    outputs(2828) <= not b;
    outputs(2829) <= not (a xor b);
    outputs(2830) <= not (a and b);
    outputs(2831) <= a;
    outputs(2832) <= a xor b;
    outputs(2833) <= not a;
    outputs(2834) <= a;
    outputs(2835) <= b;
    outputs(2836) <= b and not a;
    outputs(2837) <= not (a or b);
    outputs(2838) <= a xor b;
    outputs(2839) <= not (a xor b);
    outputs(2840) <= b;
    outputs(2841) <= b;
    outputs(2842) <= not (a xor b);
    outputs(2843) <= a;
    outputs(2844) <= not a;
    outputs(2845) <= not (a xor b);
    outputs(2846) <= a xor b;
    outputs(2847) <= not b;
    outputs(2848) <= not a or b;
    outputs(2849) <= b;
    outputs(2850) <= not (a xor b);
    outputs(2851) <= b;
    outputs(2852) <= not (a and b);
    outputs(2853) <= a xor b;
    outputs(2854) <= not (a xor b);
    outputs(2855) <= a xor b;
    outputs(2856) <= a or b;
    outputs(2857) <= a;
    outputs(2858) <= not (a xor b);
    outputs(2859) <= not b or a;
    outputs(2860) <= not b;
    outputs(2861) <= not b;
    outputs(2862) <= not b or a;
    outputs(2863) <= a xor b;
    outputs(2864) <= a;
    outputs(2865) <= not b;
    outputs(2866) <= not (a xor b);
    outputs(2867) <= b;
    outputs(2868) <= b and not a;
    outputs(2869) <= not b;
    outputs(2870) <= a and not b;
    outputs(2871) <= not a;
    outputs(2872) <= a xor b;
    outputs(2873) <= a xor b;
    outputs(2874) <= not (a xor b);
    outputs(2875) <= a;
    outputs(2876) <= a xor b;
    outputs(2877) <= a;
    outputs(2878) <= not (a xor b);
    outputs(2879) <= a;
    outputs(2880) <= a;
    outputs(2881) <= a or b;
    outputs(2882) <= a or b;
    outputs(2883) <= a and b;
    outputs(2884) <= not (a xor b);
    outputs(2885) <= not b;
    outputs(2886) <= not (a xor b);
    outputs(2887) <= not (a xor b);
    outputs(2888) <= not a;
    outputs(2889) <= not (a or b);
    outputs(2890) <= not (a xor b);
    outputs(2891) <= not (a or b);
    outputs(2892) <= not (a xor b);
    outputs(2893) <= not a;
    outputs(2894) <= a;
    outputs(2895) <= not a or b;
    outputs(2896) <= not b;
    outputs(2897) <= not (a xor b);
    outputs(2898) <= not (a xor b);
    outputs(2899) <= not (a or b);
    outputs(2900) <= not b;
    outputs(2901) <= not b;
    outputs(2902) <= not b;
    outputs(2903) <= not (a and b);
    outputs(2904) <= a xor b;
    outputs(2905) <= not (a xor b);
    outputs(2906) <= not b;
    outputs(2907) <= a;
    outputs(2908) <= not (a or b);
    outputs(2909) <= a;
    outputs(2910) <= not (a xor b);
    outputs(2911) <= b;
    outputs(2912) <= a or b;
    outputs(2913) <= b;
    outputs(2914) <= a and b;
    outputs(2915) <= not b or a;
    outputs(2916) <= not a;
    outputs(2917) <= not b;
    outputs(2918) <= a;
    outputs(2919) <= a;
    outputs(2920) <= a xor b;
    outputs(2921) <= b;
    outputs(2922) <= not b or a;
    outputs(2923) <= a and b;
    outputs(2924) <= not (a xor b);
    outputs(2925) <= not (a or b);
    outputs(2926) <= a xor b;
    outputs(2927) <= not b;
    outputs(2928) <= not a;
    outputs(2929) <= not a or b;
    outputs(2930) <= not a;
    outputs(2931) <= not (a xor b);
    outputs(2932) <= not (a and b);
    outputs(2933) <= b;
    outputs(2934) <= not (a xor b);
    outputs(2935) <= not (a xor b);
    outputs(2936) <= not b;
    outputs(2937) <= not a;
    outputs(2938) <= not (a or b);
    outputs(2939) <= b;
    outputs(2940) <= not a;
    outputs(2941) <= a xor b;
    outputs(2942) <= a xor b;
    outputs(2943) <= not (a xor b);
    outputs(2944) <= a xor b;
    outputs(2945) <= not (a and b);
    outputs(2946) <= a and b;
    outputs(2947) <= a xor b;
    outputs(2948) <= not b or a;
    outputs(2949) <= a;
    outputs(2950) <= not (a xor b);
    outputs(2951) <= not b or a;
    outputs(2952) <= not b;
    outputs(2953) <= a and not b;
    outputs(2954) <= b;
    outputs(2955) <= not (a xor b);
    outputs(2956) <= a xor b;
    outputs(2957) <= not b or a;
    outputs(2958) <= a;
    outputs(2959) <= a;
    outputs(2960) <= not (a xor b);
    outputs(2961) <= a xor b;
    outputs(2962) <= not (a xor b);
    outputs(2963) <= not b or a;
    outputs(2964) <= a;
    outputs(2965) <= not (a xor b);
    outputs(2966) <= a xor b;
    outputs(2967) <= a or b;
    outputs(2968) <= a xor b;
    outputs(2969) <= not (a xor b);
    outputs(2970) <= b and not a;
    outputs(2971) <= not (a xor b);
    outputs(2972) <= a;
    outputs(2973) <= a xor b;
    outputs(2974) <= a or b;
    outputs(2975) <= a;
    outputs(2976) <= a xor b;
    outputs(2977) <= b;
    outputs(2978) <= not b;
    outputs(2979) <= a;
    outputs(2980) <= a and b;
    outputs(2981) <= a;
    outputs(2982) <= not (a or b);
    outputs(2983) <= not b or a;
    outputs(2984) <= not (a xor b);
    outputs(2985) <= not a;
    outputs(2986) <= a and b;
    outputs(2987) <= not b;
    outputs(2988) <= not (a xor b);
    outputs(2989) <= not a;
    outputs(2990) <= not a;
    outputs(2991) <= a;
    outputs(2992) <= a and not b;
    outputs(2993) <= not (a xor b);
    outputs(2994) <= a;
    outputs(2995) <= not (a xor b);
    outputs(2996) <= not a;
    outputs(2997) <= a xor b;
    outputs(2998) <= not a;
    outputs(2999) <= a xor b;
    outputs(3000) <= a and not b;
    outputs(3001) <= not (a xor b);
    outputs(3002) <= not (a xor b);
    outputs(3003) <= a xor b;
    outputs(3004) <= not (a and b);
    outputs(3005) <= not (a xor b);
    outputs(3006) <= a;
    outputs(3007) <= not (a or b);
    outputs(3008) <= not b;
    outputs(3009) <= not a;
    outputs(3010) <= not a or b;
    outputs(3011) <= a xor b;
    outputs(3012) <= a xor b;
    outputs(3013) <= not a or b;
    outputs(3014) <= b;
    outputs(3015) <= b;
    outputs(3016) <= not b;
    outputs(3017) <= not b or a;
    outputs(3018) <= a xor b;
    outputs(3019) <= a;
    outputs(3020) <= a xor b;
    outputs(3021) <= b;
    outputs(3022) <= not (a xor b);
    outputs(3023) <= a xor b;
    outputs(3024) <= a xor b;
    outputs(3025) <= not (a or b);
    outputs(3026) <= not (a xor b);
    outputs(3027) <= a;
    outputs(3028) <= a;
    outputs(3029) <= not b;
    outputs(3030) <= not (a xor b);
    outputs(3031) <= a xor b;
    outputs(3032) <= b;
    outputs(3033) <= not (a and b);
    outputs(3034) <= not (a xor b);
    outputs(3035) <= not a;
    outputs(3036) <= not b;
    outputs(3037) <= a xor b;
    outputs(3038) <= a and b;
    outputs(3039) <= not a;
    outputs(3040) <= a xor b;
    outputs(3041) <= not (a and b);
    outputs(3042) <= not a;
    outputs(3043) <= a xor b;
    outputs(3044) <= not (a xor b);
    outputs(3045) <= not (a xor b);
    outputs(3046) <= b and not a;
    outputs(3047) <= b;
    outputs(3048) <= a xor b;
    outputs(3049) <= a xor b;
    outputs(3050) <= not b;
    outputs(3051) <= a;
    outputs(3052) <= not (a xor b);
    outputs(3053) <= a;
    outputs(3054) <= not b;
    outputs(3055) <= not (a or b);
    outputs(3056) <= b;
    outputs(3057) <= a;
    outputs(3058) <= not (a xor b);
    outputs(3059) <= a xor b;
    outputs(3060) <= not a;
    outputs(3061) <= not (a xor b);
    outputs(3062) <= not a;
    outputs(3063) <= b and not a;
    outputs(3064) <= not a;
    outputs(3065) <= a;
    outputs(3066) <= not (a xor b);
    outputs(3067) <= not (a xor b);
    outputs(3068) <= a and not b;
    outputs(3069) <= b;
    outputs(3070) <= a xor b;
    outputs(3071) <= a;
    outputs(3072) <= not b;
    outputs(3073) <= not (a xor b);
    outputs(3074) <= not (a xor b);
    outputs(3075) <= b and not a;
    outputs(3076) <= not b;
    outputs(3077) <= a xor b;
    outputs(3078) <= not (a xor b);
    outputs(3079) <= a;
    outputs(3080) <= not (a and b);
    outputs(3081) <= a and b;
    outputs(3082) <= not a;
    outputs(3083) <= a;
    outputs(3084) <= not a;
    outputs(3085) <= not (a xor b);
    outputs(3086) <= not (a xor b);
    outputs(3087) <= a;
    outputs(3088) <= not a;
    outputs(3089) <= a xor b;
    outputs(3090) <= a xor b;
    outputs(3091) <= a;
    outputs(3092) <= a;
    outputs(3093) <= a xor b;
    outputs(3094) <= not (a xor b);
    outputs(3095) <= not (a xor b);
    outputs(3096) <= b;
    outputs(3097) <= b and not a;
    outputs(3098) <= not (a or b);
    outputs(3099) <= not a;
    outputs(3100) <= a;
    outputs(3101) <= a or b;
    outputs(3102) <= a;
    outputs(3103) <= a xor b;
    outputs(3104) <= a xor b;
    outputs(3105) <= a or b;
    outputs(3106) <= not (a xor b);
    outputs(3107) <= not b;
    outputs(3108) <= not a;
    outputs(3109) <= b;
    outputs(3110) <= a xor b;
    outputs(3111) <= a or b;
    outputs(3112) <= not (a and b);
    outputs(3113) <= not a;
    outputs(3114) <= b;
    outputs(3115) <= not a;
    outputs(3116) <= not b;
    outputs(3117) <= not a;
    outputs(3118) <= b;
    outputs(3119) <= a xor b;
    outputs(3120) <= not (a xor b);
    outputs(3121) <= not b;
    outputs(3122) <= a and not b;
    outputs(3123) <= not (a xor b);
    outputs(3124) <= not a;
    outputs(3125) <= not (a xor b);
    outputs(3126) <= a xor b;
    outputs(3127) <= a xor b;
    outputs(3128) <= not a;
    outputs(3129) <= a xor b;
    outputs(3130) <= b;
    outputs(3131) <= not (a xor b);
    outputs(3132) <= not a;
    outputs(3133) <= a and b;
    outputs(3134) <= not b;
    outputs(3135) <= a xor b;
    outputs(3136) <= a or b;
    outputs(3137) <= a xor b;
    outputs(3138) <= not (a xor b);
    outputs(3139) <= not b;
    outputs(3140) <= a xor b;
    outputs(3141) <= a xor b;
    outputs(3142) <= a and b;
    outputs(3143) <= not (a xor b);
    outputs(3144) <= b;
    outputs(3145) <= b;
    outputs(3146) <= b;
    outputs(3147) <= b;
    outputs(3148) <= a and not b;
    outputs(3149) <= b;
    outputs(3150) <= a xor b;
    outputs(3151) <= a or b;
    outputs(3152) <= not b;
    outputs(3153) <= not (a xor b);
    outputs(3154) <= a and not b;
    outputs(3155) <= not a or b;
    outputs(3156) <= not (a and b);
    outputs(3157) <= a;
    outputs(3158) <= not b;
    outputs(3159) <= not a;
    outputs(3160) <= not (a or b);
    outputs(3161) <= not b;
    outputs(3162) <= not (a xor b);
    outputs(3163) <= not a;
    outputs(3164) <= a or b;
    outputs(3165) <= not b;
    outputs(3166) <= not a;
    outputs(3167) <= not b or a;
    outputs(3168) <= not b;
    outputs(3169) <= not (a xor b);
    outputs(3170) <= not (a xor b);
    outputs(3171) <= a xor b;
    outputs(3172) <= a xor b;
    outputs(3173) <= not (a or b);
    outputs(3174) <= b and not a;
    outputs(3175) <= not (a xor b);
    outputs(3176) <= a;
    outputs(3177) <= b;
    outputs(3178) <= b and not a;
    outputs(3179) <= a and b;
    outputs(3180) <= a and b;
    outputs(3181) <= a;
    outputs(3182) <= a;
    outputs(3183) <= not (a xor b);
    outputs(3184) <= not a;
    outputs(3185) <= a xor b;
    outputs(3186) <= b;
    outputs(3187) <= a xor b;
    outputs(3188) <= not (a xor b);
    outputs(3189) <= not b;
    outputs(3190) <= b;
    outputs(3191) <= not b;
    outputs(3192) <= a;
    outputs(3193) <= not a;
    outputs(3194) <= not (a xor b);
    outputs(3195) <= a xor b;
    outputs(3196) <= not (a xor b);
    outputs(3197) <= not a;
    outputs(3198) <= not b;
    outputs(3199) <= a;
    outputs(3200) <= b;
    outputs(3201) <= a;
    outputs(3202) <= not (a xor b);
    outputs(3203) <= a xor b;
    outputs(3204) <= not (a and b);
    outputs(3205) <= a xor b;
    outputs(3206) <= not b;
    outputs(3207) <= not b;
    outputs(3208) <= b;
    outputs(3209) <= not (a xor b);
    outputs(3210) <= not (a and b);
    outputs(3211) <= b;
    outputs(3212) <= not (a xor b);
    outputs(3213) <= not b;
    outputs(3214) <= not a;
    outputs(3215) <= a and b;
    outputs(3216) <= not b;
    outputs(3217) <= a;
    outputs(3218) <= not b;
    outputs(3219) <= not (a and b);
    outputs(3220) <= a;
    outputs(3221) <= b and not a;
    outputs(3222) <= a xor b;
    outputs(3223) <= not a;
    outputs(3224) <= a xor b;
    outputs(3225) <= not (a or b);
    outputs(3226) <= not a or b;
    outputs(3227) <= a;
    outputs(3228) <= not b;
    outputs(3229) <= b and not a;
    outputs(3230) <= not (a xor b);
    outputs(3231) <= not (a xor b);
    outputs(3232) <= b;
    outputs(3233) <= a xor b;
    outputs(3234) <= a xor b;
    outputs(3235) <= not a or b;
    outputs(3236) <= a xor b;
    outputs(3237) <= not a;
    outputs(3238) <= a;
    outputs(3239) <= not (a xor b);
    outputs(3240) <= a xor b;
    outputs(3241) <= a xor b;
    outputs(3242) <= not b;
    outputs(3243) <= a;
    outputs(3244) <= not (a or b);
    outputs(3245) <= a xor b;
    outputs(3246) <= not (a and b);
    outputs(3247) <= a;
    outputs(3248) <= b and not a;
    outputs(3249) <= a;
    outputs(3250) <= not a;
    outputs(3251) <= not (a xor b);
    outputs(3252) <= not (a xor b);
    outputs(3253) <= not b;
    outputs(3254) <= not a;
    outputs(3255) <= not (a xor b);
    outputs(3256) <= not (a xor b);
    outputs(3257) <= a and not b;
    outputs(3258) <= a xor b;
    outputs(3259) <= not a;
    outputs(3260) <= a;
    outputs(3261) <= not b;
    outputs(3262) <= b;
    outputs(3263) <= a xor b;
    outputs(3264) <= a and not b;
    outputs(3265) <= b;
    outputs(3266) <= a xor b;
    outputs(3267) <= not (a xor b);
    outputs(3268) <= not (a or b);
    outputs(3269) <= not a or b;
    outputs(3270) <= not a;
    outputs(3271) <= not b;
    outputs(3272) <= a xor b;
    outputs(3273) <= a and b;
    outputs(3274) <= a xor b;
    outputs(3275) <= b;
    outputs(3276) <= a and not b;
    outputs(3277) <= not b;
    outputs(3278) <= a xor b;
    outputs(3279) <= not a or b;
    outputs(3280) <= a and b;
    outputs(3281) <= not b;
    outputs(3282) <= a;
    outputs(3283) <= a;
    outputs(3284) <= a;
    outputs(3285) <= b;
    outputs(3286) <= not b;
    outputs(3287) <= a xor b;
    outputs(3288) <= a xor b;
    outputs(3289) <= a xor b;
    outputs(3290) <= not (a xor b);
    outputs(3291) <= b and not a;
    outputs(3292) <= not a;
    outputs(3293) <= a and not b;
    outputs(3294) <= not b;
    outputs(3295) <= a xor b;
    outputs(3296) <= a xor b;
    outputs(3297) <= not (a xor b);
    outputs(3298) <= not b or a;
    outputs(3299) <= a or b;
    outputs(3300) <= b and not a;
    outputs(3301) <= a and not b;
    outputs(3302) <= not a;
    outputs(3303) <= a xor b;
    outputs(3304) <= a;
    outputs(3305) <= b;
    outputs(3306) <= not (a xor b);
    outputs(3307) <= not a;
    outputs(3308) <= not (a xor b);
    outputs(3309) <= not a;
    outputs(3310) <= not a;
    outputs(3311) <= not a;
    outputs(3312) <= not b;
    outputs(3313) <= a xor b;
    outputs(3314) <= a;
    outputs(3315) <= not a or b;
    outputs(3316) <= not a;
    outputs(3317) <= a;
    outputs(3318) <= not (a xor b);
    outputs(3319) <= not a;
    outputs(3320) <= not (a xor b);
    outputs(3321) <= not a;
    outputs(3322) <= not (a or b);
    outputs(3323) <= not a;
    outputs(3324) <= a xor b;
    outputs(3325) <= b;
    outputs(3326) <= a xor b;
    outputs(3327) <= a;
    outputs(3328) <= not b or a;
    outputs(3329) <= not b;
    outputs(3330) <= a and not b;
    outputs(3331) <= not a;
    outputs(3332) <= a and not b;
    outputs(3333) <= a xor b;
    outputs(3334) <= a;
    outputs(3335) <= not b or a;
    outputs(3336) <= b and not a;
    outputs(3337) <= not a;
    outputs(3338) <= a or b;
    outputs(3339) <= a;
    outputs(3340) <= a xor b;
    outputs(3341) <= a xor b;
    outputs(3342) <= not a;
    outputs(3343) <= not a;
    outputs(3344) <= not b or a;
    outputs(3345) <= not (a xor b);
    outputs(3346) <= a xor b;
    outputs(3347) <= not a;
    outputs(3348) <= not (a xor b);
    outputs(3349) <= not (a and b);
    outputs(3350) <= not b;
    outputs(3351) <= a xor b;
    outputs(3352) <= not (a xor b);
    outputs(3353) <= not (a xor b);
    outputs(3354) <= a xor b;
    outputs(3355) <= a;
    outputs(3356) <= b;
    outputs(3357) <= not (a and b);
    outputs(3358) <= a and b;
    outputs(3359) <= a and b;
    outputs(3360) <= b;
    outputs(3361) <= not b;
    outputs(3362) <= not b or a;
    outputs(3363) <= b;
    outputs(3364) <= not (a xor b);
    outputs(3365) <= not (a xor b);
    outputs(3366) <= b;
    outputs(3367) <= not a or b;
    outputs(3368) <= not (a and b);
    outputs(3369) <= not (a xor b);
    outputs(3370) <= b;
    outputs(3371) <= a and not b;
    outputs(3372) <= not a;
    outputs(3373) <= not a;
    outputs(3374) <= not (a xor b);
    outputs(3375) <= not (a xor b);
    outputs(3376) <= not b;
    outputs(3377) <= not (a xor b);
    outputs(3378) <= not (a and b);
    outputs(3379) <= a xor b;
    outputs(3380) <= a and not b;
    outputs(3381) <= not a or b;
    outputs(3382) <= a;
    outputs(3383) <= not a or b;
    outputs(3384) <= b and not a;
    outputs(3385) <= not a;
    outputs(3386) <= not a;
    outputs(3387) <= not a;
    outputs(3388) <= not a;
    outputs(3389) <= a and not b;
    outputs(3390) <= not b;
    outputs(3391) <= not a;
    outputs(3392) <= not a;
    outputs(3393) <= a;
    outputs(3394) <= not (a xor b);
    outputs(3395) <= a xor b;
    outputs(3396) <= not b;
    outputs(3397) <= not a;
    outputs(3398) <= not a;
    outputs(3399) <= not a;
    outputs(3400) <= a or b;
    outputs(3401) <= not b;
    outputs(3402) <= a xor b;
    outputs(3403) <= b;
    outputs(3404) <= not (a xor b);
    outputs(3405) <= b and not a;
    outputs(3406) <= not (a xor b);
    outputs(3407) <= not (a xor b);
    outputs(3408) <= not (a xor b);
    outputs(3409) <= a xor b;
    outputs(3410) <= not (a and b);
    outputs(3411) <= a or b;
    outputs(3412) <= b;
    outputs(3413) <= a xor b;
    outputs(3414) <= a xor b;
    outputs(3415) <= b;
    outputs(3416) <= not (a xor b);
    outputs(3417) <= b;
    outputs(3418) <= a xor b;
    outputs(3419) <= not (a xor b);
    outputs(3420) <= not (a xor b);
    outputs(3421) <= a and not b;
    outputs(3422) <= b;
    outputs(3423) <= not a;
    outputs(3424) <= not a;
    outputs(3425) <= a and b;
    outputs(3426) <= not b;
    outputs(3427) <= not (a xor b);
    outputs(3428) <= a;
    outputs(3429) <= not (a xor b);
    outputs(3430) <= not (a xor b);
    outputs(3431) <= a;
    outputs(3432) <= a xor b;
    outputs(3433) <= b;
    outputs(3434) <= not b;
    outputs(3435) <= not (a xor b);
    outputs(3436) <= a and not b;
    outputs(3437) <= a xor b;
    outputs(3438) <= not (a xor b);
    outputs(3439) <= not (a xor b);
    outputs(3440) <= a;
    outputs(3441) <= not (a xor b);
    outputs(3442) <= a xor b;
    outputs(3443) <= not (a xor b);
    outputs(3444) <= not b;
    outputs(3445) <= a;
    outputs(3446) <= not a;
    outputs(3447) <= b;
    outputs(3448) <= not (a xor b);
    outputs(3449) <= not a;
    outputs(3450) <= not (a xor b);
    outputs(3451) <= a xor b;
    outputs(3452) <= not (a xor b);
    outputs(3453) <= not (a xor b);
    outputs(3454) <= b;
    outputs(3455) <= a or b;
    outputs(3456) <= not (a xor b);
    outputs(3457) <= a;
    outputs(3458) <= a and b;
    outputs(3459) <= a xor b;
    outputs(3460) <= a;
    outputs(3461) <= not a;
    outputs(3462) <= a;
    outputs(3463) <= a;
    outputs(3464) <= not a;
    outputs(3465) <= a xor b;
    outputs(3466) <= not (a xor b);
    outputs(3467) <= not (a xor b);
    outputs(3468) <= b;
    outputs(3469) <= a and not b;
    outputs(3470) <= b;
    outputs(3471) <= a xor b;
    outputs(3472) <= not a;
    outputs(3473) <= not (a xor b);
    outputs(3474) <= b;
    outputs(3475) <= b;
    outputs(3476) <= a or b;
    outputs(3477) <= not (a xor b);
    outputs(3478) <= a;
    outputs(3479) <= not b;
    outputs(3480) <= not (a xor b);
    outputs(3481) <= a xor b;
    outputs(3482) <= not b;
    outputs(3483) <= a;
    outputs(3484) <= a;
    outputs(3485) <= a xor b;
    outputs(3486) <= not (a xor b);
    outputs(3487) <= not (a xor b);
    outputs(3488) <= a or b;
    outputs(3489) <= not (a xor b);
    outputs(3490) <= not (a and b);
    outputs(3491) <= b and not a;
    outputs(3492) <= a;
    outputs(3493) <= not b;
    outputs(3494) <= not (a and b);
    outputs(3495) <= not a;
    outputs(3496) <= a xor b;
    outputs(3497) <= not a or b;
    outputs(3498) <= b;
    outputs(3499) <= a;
    outputs(3500) <= not (a xor b);
    outputs(3501) <= a xor b;
    outputs(3502) <= a xor b;
    outputs(3503) <= not (a xor b);
    outputs(3504) <= a xor b;
    outputs(3505) <= not (a xor b);
    outputs(3506) <= a xor b;
    outputs(3507) <= not b;
    outputs(3508) <= a xor b;
    outputs(3509) <= a xor b;
    outputs(3510) <= not a;
    outputs(3511) <= not b;
    outputs(3512) <= a xor b;
    outputs(3513) <= not b;
    outputs(3514) <= not a;
    outputs(3515) <= a xor b;
    outputs(3516) <= not a;
    outputs(3517) <= a xor b;
    outputs(3518) <= b;
    outputs(3519) <= not (a xor b);
    outputs(3520) <= a xor b;
    outputs(3521) <= not a or b;
    outputs(3522) <= a;
    outputs(3523) <= a and not b;
    outputs(3524) <= not b;
    outputs(3525) <= a and not b;
    outputs(3526) <= not (a xor b);
    outputs(3527) <= a;
    outputs(3528) <= b;
    outputs(3529) <= not a;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= not b;
    outputs(3532) <= not (a xor b);
    outputs(3533) <= a and not b;
    outputs(3534) <= a;
    outputs(3535) <= a;
    outputs(3536) <= b and not a;
    outputs(3537) <= not b;
    outputs(3538) <= not a or b;
    outputs(3539) <= not (a or b);
    outputs(3540) <= a xor b;
    outputs(3541) <= b;
    outputs(3542) <= not b;
    outputs(3543) <= b and not a;
    outputs(3544) <= not a;
    outputs(3545) <= not b;
    outputs(3546) <= not (a xor b);
    outputs(3547) <= not b;
    outputs(3548) <= a xor b;
    outputs(3549) <= b;
    outputs(3550) <= not (a xor b);
    outputs(3551) <= not a or b;
    outputs(3552) <= a and b;
    outputs(3553) <= not (a xor b);
    outputs(3554) <= not b;
    outputs(3555) <= not b;
    outputs(3556) <= a;
    outputs(3557) <= not (a xor b);
    outputs(3558) <= not (a xor b);
    outputs(3559) <= not (a xor b);
    outputs(3560) <= a xor b;
    outputs(3561) <= not (a and b);
    outputs(3562) <= a;
    outputs(3563) <= a and b;
    outputs(3564) <= a xor b;
    outputs(3565) <= b;
    outputs(3566) <= a;
    outputs(3567) <= not (a and b);
    outputs(3568) <= not b;
    outputs(3569) <= not (a xor b);
    outputs(3570) <= a;
    outputs(3571) <= a xor b;
    outputs(3572) <= a xor b;
    outputs(3573) <= not b;
    outputs(3574) <= not b or a;
    outputs(3575) <= a and b;
    outputs(3576) <= not a;
    outputs(3577) <= not b;
    outputs(3578) <= a;
    outputs(3579) <= not b;
    outputs(3580) <= a or b;
    outputs(3581) <= not b;
    outputs(3582) <= a and not b;
    outputs(3583) <= not (a or b);
    outputs(3584) <= not b;
    outputs(3585) <= not b;
    outputs(3586) <= a;
    outputs(3587) <= not a or b;
    outputs(3588) <= b;
    outputs(3589) <= not (a xor b);
    outputs(3590) <= not (a xor b);
    outputs(3591) <= not (a or b);
    outputs(3592) <= a or b;
    outputs(3593) <= b and not a;
    outputs(3594) <= not a;
    outputs(3595) <= a;
    outputs(3596) <= a;
    outputs(3597) <= not a;
    outputs(3598) <= not (a xor b);
    outputs(3599) <= b;
    outputs(3600) <= not b;
    outputs(3601) <= a xor b;
    outputs(3602) <= b;
    outputs(3603) <= not (a xor b);
    outputs(3604) <= not a;
    outputs(3605) <= not (a xor b);
    outputs(3606) <= a;
    outputs(3607) <= a xor b;
    outputs(3608) <= not (a xor b);
    outputs(3609) <= a xor b;
    outputs(3610) <= not a or b;
    outputs(3611) <= not a;
    outputs(3612) <= a xor b;
    outputs(3613) <= a;
    outputs(3614) <= not a or b;
    outputs(3615) <= b;
    outputs(3616) <= a xor b;
    outputs(3617) <= a;
    outputs(3618) <= not b;
    outputs(3619) <= not (a xor b);
    outputs(3620) <= not b;
    outputs(3621) <= not (a xor b);
    outputs(3622) <= b;
    outputs(3623) <= not b;
    outputs(3624) <= b;
    outputs(3625) <= not (a xor b);
    outputs(3626) <= not (a and b);
    outputs(3627) <= not (a and b);
    outputs(3628) <= b;
    outputs(3629) <= a and b;
    outputs(3630) <= a xor b;
    outputs(3631) <= a;
    outputs(3632) <= not a or b;
    outputs(3633) <= a xor b;
    outputs(3634) <= b;
    outputs(3635) <= a;
    outputs(3636) <= not a or b;
    outputs(3637) <= not (a or b);
    outputs(3638) <= a and not b;
    outputs(3639) <= not a;
    outputs(3640) <= not (a xor b);
    outputs(3641) <= a;
    outputs(3642) <= a xor b;
    outputs(3643) <= a xor b;
    outputs(3644) <= not (a and b);
    outputs(3645) <= a xor b;
    outputs(3646) <= not (a xor b);
    outputs(3647) <= not b;
    outputs(3648) <= not (a xor b);
    outputs(3649) <= a or b;
    outputs(3650) <= b;
    outputs(3651) <= not (a and b);
    outputs(3652) <= not (a xor b);
    outputs(3653) <= a;
    outputs(3654) <= not (a xor b);
    outputs(3655) <= b;
    outputs(3656) <= not a;
    outputs(3657) <= not a;
    outputs(3658) <= a or b;
    outputs(3659) <= not b;
    outputs(3660) <= not (a xor b);
    outputs(3661) <= not b or a;
    outputs(3662) <= a xor b;
    outputs(3663) <= a;
    outputs(3664) <= a xor b;
    outputs(3665) <= not (a xor b);
    outputs(3666) <= not (a xor b);
    outputs(3667) <= a and not b;
    outputs(3668) <= not a;
    outputs(3669) <= not a or b;
    outputs(3670) <= not (a and b);
    outputs(3671) <= a or b;
    outputs(3672) <= b;
    outputs(3673) <= a xor b;
    outputs(3674) <= not a;
    outputs(3675) <= b;
    outputs(3676) <= a xor b;
    outputs(3677) <= b;
    outputs(3678) <= not b;
    outputs(3679) <= not b;
    outputs(3680) <= not (a and b);
    outputs(3681) <= not (a xor b);
    outputs(3682) <= not a;
    outputs(3683) <= b and not a;
    outputs(3684) <= b;
    outputs(3685) <= not (a xor b);
    outputs(3686) <= not b;
    outputs(3687) <= b;
    outputs(3688) <= a and not b;
    outputs(3689) <= b;
    outputs(3690) <= not (a xor b);
    outputs(3691) <= a xor b;
    outputs(3692) <= a;
    outputs(3693) <= not b;
    outputs(3694) <= a;
    outputs(3695) <= not (a xor b);
    outputs(3696) <= not b;
    outputs(3697) <= not (a xor b);
    outputs(3698) <= not b;
    outputs(3699) <= not b or a;
    outputs(3700) <= a xor b;
    outputs(3701) <= not (a xor b);
    outputs(3702) <= not a or b;
    outputs(3703) <= not (a xor b);
    outputs(3704) <= not b;
    outputs(3705) <= not b;
    outputs(3706) <= a xor b;
    outputs(3707) <= a xor b;
    outputs(3708) <= a;
    outputs(3709) <= not b or a;
    outputs(3710) <= a xor b;
    outputs(3711) <= not b;
    outputs(3712) <= b;
    outputs(3713) <= a and b;
    outputs(3714) <= a or b;
    outputs(3715) <= a and b;
    outputs(3716) <= a xor b;
    outputs(3717) <= not (a xor b);
    outputs(3718) <= b;
    outputs(3719) <= a or b;
    outputs(3720) <= not (a and b);
    outputs(3721) <= not a;
    outputs(3722) <= not (a and b);
    outputs(3723) <= not b;
    outputs(3724) <= a xor b;
    outputs(3725) <= b;
    outputs(3726) <= not a;
    outputs(3727) <= b;
    outputs(3728) <= not b;
    outputs(3729) <= a xor b;
    outputs(3730) <= a xor b;
    outputs(3731) <= b;
    outputs(3732) <= not (a xor b);
    outputs(3733) <= not (a xor b);
    outputs(3734) <= not (a or b);
    outputs(3735) <= a;
    outputs(3736) <= not (a xor b);
    outputs(3737) <= not b;
    outputs(3738) <= not a or b;
    outputs(3739) <= not a;
    outputs(3740) <= not (a xor b);
    outputs(3741) <= not b;
    outputs(3742) <= not b;
    outputs(3743) <= not b;
    outputs(3744) <= not (a xor b);
    outputs(3745) <= b;
    outputs(3746) <= not b;
    outputs(3747) <= not b;
    outputs(3748) <= not b;
    outputs(3749) <= a;
    outputs(3750) <= a xor b;
    outputs(3751) <= not b;
    outputs(3752) <= not (a xor b);
    outputs(3753) <= b;
    outputs(3754) <= a xor b;
    outputs(3755) <= not a or b;
    outputs(3756) <= not (a xor b);
    outputs(3757) <= a;
    outputs(3758) <= not (a xor b);
    outputs(3759) <= a xor b;
    outputs(3760) <= a and not b;
    outputs(3761) <= not (a and b);
    outputs(3762) <= a xor b;
    outputs(3763) <= a;
    outputs(3764) <= b;
    outputs(3765) <= a and b;
    outputs(3766) <= not (a xor b);
    outputs(3767) <= a xor b;
    outputs(3768) <= b;
    outputs(3769) <= not a;
    outputs(3770) <= not (a or b);
    outputs(3771) <= a xor b;
    outputs(3772) <= not a;
    outputs(3773) <= not a;
    outputs(3774) <= not (a or b);
    outputs(3775) <= not b;
    outputs(3776) <= b;
    outputs(3777) <= not a;
    outputs(3778) <= a xor b;
    outputs(3779) <= not (a xor b);
    outputs(3780) <= not b;
    outputs(3781) <= not a or b;
    outputs(3782) <= a xor b;
    outputs(3783) <= not a;
    outputs(3784) <= not a;
    outputs(3785) <= a;
    outputs(3786) <= b;
    outputs(3787) <= not (a xor b);
    outputs(3788) <= not (a xor b);
    outputs(3789) <= not b;
    outputs(3790) <= not (a or b);
    outputs(3791) <= not (a xor b);
    outputs(3792) <= a or b;
    outputs(3793) <= a;
    outputs(3794) <= not b;
    outputs(3795) <= a xor b;
    outputs(3796) <= not a or b;
    outputs(3797) <= a or b;
    outputs(3798) <= not b;
    outputs(3799) <= not b;
    outputs(3800) <= b;
    outputs(3801) <= b;
    outputs(3802) <= not (a xor b);
    outputs(3803) <= a xor b;
    outputs(3804) <= a xor b;
    outputs(3805) <= not (a xor b);
    outputs(3806) <= not b or a;
    outputs(3807) <= not (a xor b);
    outputs(3808) <= b;
    outputs(3809) <= not b;
    outputs(3810) <= b;
    outputs(3811) <= not a;
    outputs(3812) <= not (a xor b);
    outputs(3813) <= not a;
    outputs(3814) <= not (a xor b);
    outputs(3815) <= not b;
    outputs(3816) <= a;
    outputs(3817) <= a xor b;
    outputs(3818) <= not a;
    outputs(3819) <= not a;
    outputs(3820) <= not b;
    outputs(3821) <= not b;
    outputs(3822) <= not a or b;
    outputs(3823) <= not b;
    outputs(3824) <= not b;
    outputs(3825) <= not a;
    outputs(3826) <= not (a and b);
    outputs(3827) <= b;
    outputs(3828) <= not (a xor b);
    outputs(3829) <= a xor b;
    outputs(3830) <= a and b;
    outputs(3831) <= a xor b;
    outputs(3832) <= a xor b;
    outputs(3833) <= a;
    outputs(3834) <= not a or b;
    outputs(3835) <= not a;
    outputs(3836) <= a or b;
    outputs(3837) <= not (a or b);
    outputs(3838) <= b;
    outputs(3839) <= not a;
    outputs(3840) <= not (a xor b);
    outputs(3841) <= not (a xor b);
    outputs(3842) <= not a;
    outputs(3843) <= a xor b;
    outputs(3844) <= not a;
    outputs(3845) <= not a;
    outputs(3846) <= b;
    outputs(3847) <= a xor b;
    outputs(3848) <= b;
    outputs(3849) <= a xor b;
    outputs(3850) <= not (a xor b);
    outputs(3851) <= a xor b;
    outputs(3852) <= not a;
    outputs(3853) <= a xor b;
    outputs(3854) <= a and not b;
    outputs(3855) <= not a;
    outputs(3856) <= b and not a;
    outputs(3857) <= a xor b;
    outputs(3858) <= not a or b;
    outputs(3859) <= not (a or b);
    outputs(3860) <= a;
    outputs(3861) <= a xor b;
    outputs(3862) <= a;
    outputs(3863) <= b;
    outputs(3864) <= a xor b;
    outputs(3865) <= not (a or b);
    outputs(3866) <= b;
    outputs(3867) <= not (a xor b);
    outputs(3868) <= not a or b;
    outputs(3869) <= b;
    outputs(3870) <= a;
    outputs(3871) <= a;
    outputs(3872) <= not (a or b);
    outputs(3873) <= a;
    outputs(3874) <= a xor b;
    outputs(3875) <= not b or a;
    outputs(3876) <= a;
    outputs(3877) <= not (a xor b);
    outputs(3878) <= a xor b;
    outputs(3879) <= a or b;
    outputs(3880) <= not a;
    outputs(3881) <= a;
    outputs(3882) <= not b;
    outputs(3883) <= not (a xor b);
    outputs(3884) <= b;
    outputs(3885) <= a and not b;
    outputs(3886) <= b;
    outputs(3887) <= b;
    outputs(3888) <= not (a xor b);
    outputs(3889) <= a;
    outputs(3890) <= not b;
    outputs(3891) <= b;
    outputs(3892) <= not a or b;
    outputs(3893) <= b;
    outputs(3894) <= not b;
    outputs(3895) <= a and b;
    outputs(3896) <= not (a xor b);
    outputs(3897) <= a xor b;
    outputs(3898) <= not b;
    outputs(3899) <= a;
    outputs(3900) <= not (a xor b);
    outputs(3901) <= a xor b;
    outputs(3902) <= not a;
    outputs(3903) <= b;
    outputs(3904) <= not (a xor b);
    outputs(3905) <= a xor b;
    outputs(3906) <= a xor b;
    outputs(3907) <= b;
    outputs(3908) <= a and b;
    outputs(3909) <= not (a xor b);
    outputs(3910) <= b;
    outputs(3911) <= not (a and b);
    outputs(3912) <= a or b;
    outputs(3913) <= a xor b;
    outputs(3914) <= a;
    outputs(3915) <= not a;
    outputs(3916) <= not (a xor b);
    outputs(3917) <= not (a xor b);
    outputs(3918) <= a xor b;
    outputs(3919) <= a and not b;
    outputs(3920) <= not a or b;
    outputs(3921) <= a;
    outputs(3922) <= not a or b;
    outputs(3923) <= b;
    outputs(3924) <= b and not a;
    outputs(3925) <= not b;
    outputs(3926) <= b;
    outputs(3927) <= not (a or b);
    outputs(3928) <= a xor b;
    outputs(3929) <= not (a xor b);
    outputs(3930) <= not b;
    outputs(3931) <= not b or a;
    outputs(3932) <= a or b;
    outputs(3933) <= b and not a;
    outputs(3934) <= b;
    outputs(3935) <= not b;
    outputs(3936) <= b;
    outputs(3937) <= not (a xor b);
    outputs(3938) <= not (a xor b);
    outputs(3939) <= a xor b;
    outputs(3940) <= a;
    outputs(3941) <= a xor b;
    outputs(3942) <= a xor b;
    outputs(3943) <= not (a xor b);
    outputs(3944) <= a;
    outputs(3945) <= not (a xor b);
    outputs(3946) <= b and not a;
    outputs(3947) <= b;
    outputs(3948) <= not (a xor b);
    outputs(3949) <= b;
    outputs(3950) <= a;
    outputs(3951) <= a xor b;
    outputs(3952) <= b;
    outputs(3953) <= not (a xor b);
    outputs(3954) <= a;
    outputs(3955) <= not (a or b);
    outputs(3956) <= a or b;
    outputs(3957) <= not (a xor b);
    outputs(3958) <= not (a xor b);
    outputs(3959) <= not (a xor b);
    outputs(3960) <= not b;
    outputs(3961) <= a xor b;
    outputs(3962) <= a;
    outputs(3963) <= not a;
    outputs(3964) <= a;
    outputs(3965) <= a xor b;
    outputs(3966) <= a or b;
    outputs(3967) <= not (a or b);
    outputs(3968) <= not b;
    outputs(3969) <= not (a or b);
    outputs(3970) <= a or b;
    outputs(3971) <= b;
    outputs(3972) <= not b;
    outputs(3973) <= not b or a;
    outputs(3974) <= not b;
    outputs(3975) <= b;
    outputs(3976) <= a;
    outputs(3977) <= not b or a;
    outputs(3978) <= a xor b;
    outputs(3979) <= a;
    outputs(3980) <= not (a or b);
    outputs(3981) <= not (a xor b);
    outputs(3982) <= b;
    outputs(3983) <= not a;
    outputs(3984) <= b;
    outputs(3985) <= a;
    outputs(3986) <= not (a xor b);
    outputs(3987) <= a;
    outputs(3988) <= not (a xor b);
    outputs(3989) <= b;
    outputs(3990) <= not b;
    outputs(3991) <= not (a xor b);
    outputs(3992) <= a xor b;
    outputs(3993) <= not (a xor b);
    outputs(3994) <= not b;
    outputs(3995) <= not a;
    outputs(3996) <= not a;
    outputs(3997) <= a and not b;
    outputs(3998) <= a and not b;
    outputs(3999) <= not b;
    outputs(4000) <= not b;
    outputs(4001) <= b and not a;
    outputs(4002) <= a;
    outputs(4003) <= b and not a;
    outputs(4004) <= a xor b;
    outputs(4005) <= b;
    outputs(4006) <= a;
    outputs(4007) <= not b;
    outputs(4008) <= b;
    outputs(4009) <= not (a xor b);
    outputs(4010) <= a or b;
    outputs(4011) <= b;
    outputs(4012) <= b;
    outputs(4013) <= not (a xor b);
    outputs(4014) <= not (a xor b);
    outputs(4015) <= a xor b;
    outputs(4016) <= not a or b;
    outputs(4017) <= a xor b;
    outputs(4018) <= not a;
    outputs(4019) <= a;
    outputs(4020) <= b and not a;
    outputs(4021) <= not b;
    outputs(4022) <= a xor b;
    outputs(4023) <= a;
    outputs(4024) <= not b;
    outputs(4025) <= a xor b;
    outputs(4026) <= a or b;
    outputs(4027) <= not (a xor b);
    outputs(4028) <= a;
    outputs(4029) <= a;
    outputs(4030) <= a;
    outputs(4031) <= not b;
    outputs(4032) <= a;
    outputs(4033) <= not a;
    outputs(4034) <= b and not a;
    outputs(4035) <= a and b;
    outputs(4036) <= a xor b;
    outputs(4037) <= a xor b;
    outputs(4038) <= not (a or b);
    outputs(4039) <= not a or b;
    outputs(4040) <= b;
    outputs(4041) <= not (a xor b);
    outputs(4042) <= b;
    outputs(4043) <= not (a xor b);
    outputs(4044) <= a;
    outputs(4045) <= not (a xor b);
    outputs(4046) <= not a;
    outputs(4047) <= a;
    outputs(4048) <= a;
    outputs(4049) <= a and not b;
    outputs(4050) <= not b;
    outputs(4051) <= not b;
    outputs(4052) <= a;
    outputs(4053) <= not (a xor b);
    outputs(4054) <= not (a xor b);
    outputs(4055) <= not a;
    outputs(4056) <= a xor b;
    outputs(4057) <= not (a xor b);
    outputs(4058) <= a xor b;
    outputs(4059) <= not b;
    outputs(4060) <= not a;
    outputs(4061) <= a xor b;
    outputs(4062) <= a and b;
    outputs(4063) <= a xor b;
    outputs(4064) <= a xor b;
    outputs(4065) <= not b;
    outputs(4066) <= b;
    outputs(4067) <= not b;
    outputs(4068) <= a and b;
    outputs(4069) <= a xor b;
    outputs(4070) <= not b;
    outputs(4071) <= b;
    outputs(4072) <= a xor b;
    outputs(4073) <= not b;
    outputs(4074) <= not b;
    outputs(4075) <= not b;
    outputs(4076) <= a;
    outputs(4077) <= not (a xor b);
    outputs(4078) <= a xor b;
    outputs(4079) <= not a;
    outputs(4080) <= a xor b;
    outputs(4081) <= not a or b;
    outputs(4082) <= not (a xor b);
    outputs(4083) <= a xor b;
    outputs(4084) <= not (a or b);
    outputs(4085) <= a;
    outputs(4086) <= b;
    outputs(4087) <= a;
    outputs(4088) <= not (a xor b);
    outputs(4089) <= not (a xor b);
    outputs(4090) <= not a;
    outputs(4091) <= a;
    outputs(4092) <= a or b;
    outputs(4093) <= a;
    outputs(4094) <= not (a and b);
    outputs(4095) <= not a;
    outputs(4096) <= not (a xor b);
    outputs(4097) <= a;
    outputs(4098) <= b and not a;
    outputs(4099) <= a xor b;
    outputs(4100) <= not b or a;
    outputs(4101) <= not (a xor b);
    outputs(4102) <= not a;
    outputs(4103) <= b and not a;
    outputs(4104) <= not b;
    outputs(4105) <= not a;
    outputs(4106) <= not b;
    outputs(4107) <= not (a and b);
    outputs(4108) <= not (a xor b);
    outputs(4109) <= a and not b;
    outputs(4110) <= not b;
    outputs(4111) <= a xor b;
    outputs(4112) <= not b;
    outputs(4113) <= a;
    outputs(4114) <= a or b;
    outputs(4115) <= not (a or b);
    outputs(4116) <= a xor b;
    outputs(4117) <= b;
    outputs(4118) <= a and not b;
    outputs(4119) <= not a;
    outputs(4120) <= not b;
    outputs(4121) <= not (a xor b);
    outputs(4122) <= not b;
    outputs(4123) <= not b;
    outputs(4124) <= not (a xor b);
    outputs(4125) <= b;
    outputs(4126) <= a and not b;
    outputs(4127) <= not (a xor b);
    outputs(4128) <= a xor b;
    outputs(4129) <= not a;
    outputs(4130) <= not (a xor b);
    outputs(4131) <= b;
    outputs(4132) <= a or b;
    outputs(4133) <= not (a and b);
    outputs(4134) <= a xor b;
    outputs(4135) <= not (a or b);
    outputs(4136) <= not b;
    outputs(4137) <= not (a or b);
    outputs(4138) <= a xor b;
    outputs(4139) <= a xor b;
    outputs(4140) <= not a;
    outputs(4141) <= not (a xor b);
    outputs(4142) <= b and not a;
    outputs(4143) <= b;
    outputs(4144) <= not a;
    outputs(4145) <= a xor b;
    outputs(4146) <= not a;
    outputs(4147) <= not b or a;
    outputs(4148) <= b;
    outputs(4149) <= not (a xor b);
    outputs(4150) <= a and b;
    outputs(4151) <= a xor b;
    outputs(4152) <= b;
    outputs(4153) <= a;
    outputs(4154) <= b and not a;
    outputs(4155) <= b;
    outputs(4156) <= not b;
    outputs(4157) <= not (a or b);
    outputs(4158) <= not a;
    outputs(4159) <= not (a and b);
    outputs(4160) <= not (a xor b);
    outputs(4161) <= not (a xor b);
    outputs(4162) <= a xor b;
    outputs(4163) <= a and b;
    outputs(4164) <= not a;
    outputs(4165) <= a;
    outputs(4166) <= not (a xor b);
    outputs(4167) <= b and not a;
    outputs(4168) <= b;
    outputs(4169) <= a and b;
    outputs(4170) <= not b;
    outputs(4171) <= a xor b;
    outputs(4172) <= not b;
    outputs(4173) <= a or b;
    outputs(4174) <= a xor b;
    outputs(4175) <= not (a xor b);
    outputs(4176) <= not (a xor b);
    outputs(4177) <= a;
    outputs(4178) <= not b or a;
    outputs(4179) <= a xor b;
    outputs(4180) <= not (a xor b);
    outputs(4181) <= not (a xor b);
    outputs(4182) <= a xor b;
    outputs(4183) <= not (a xor b);
    outputs(4184) <= not a;
    outputs(4185) <= a xor b;
    outputs(4186) <= a;
    outputs(4187) <= b;
    outputs(4188) <= b;
    outputs(4189) <= a xor b;
    outputs(4190) <= a xor b;
    outputs(4191) <= not (a xor b);
    outputs(4192) <= b;
    outputs(4193) <= not b;
    outputs(4194) <= not a;
    outputs(4195) <= a;
    outputs(4196) <= not (a xor b);
    outputs(4197) <= a xor b;
    outputs(4198) <= a xor b;
    outputs(4199) <= a xor b;
    outputs(4200) <= not (a xor b);
    outputs(4201) <= not b or a;
    outputs(4202) <= a xor b;
    outputs(4203) <= not a;
    outputs(4204) <= not b;
    outputs(4205) <= not a;
    outputs(4206) <= not b;
    outputs(4207) <= not a;
    outputs(4208) <= not a;
    outputs(4209) <= not b or a;
    outputs(4210) <= b;
    outputs(4211) <= not a or b;
    outputs(4212) <= not (a and b);
    outputs(4213) <= not (a or b);
    outputs(4214) <= b;
    outputs(4215) <= not (a xor b);
    outputs(4216) <= not (a xor b);
    outputs(4217) <= not (a xor b);
    outputs(4218) <= b;
    outputs(4219) <= b;
    outputs(4220) <= not (a xor b);
    outputs(4221) <= a and b;
    outputs(4222) <= b;
    outputs(4223) <= not (a xor b);
    outputs(4224) <= not b;
    outputs(4225) <= not a;
    outputs(4226) <= a xor b;
    outputs(4227) <= not (a xor b);
    outputs(4228) <= a xor b;
    outputs(4229) <= not a;
    outputs(4230) <= b;
    outputs(4231) <= b;
    outputs(4232) <= a;
    outputs(4233) <= a;
    outputs(4234) <= b and not a;
    outputs(4235) <= not a;
    outputs(4236) <= not a or b;
    outputs(4237) <= not (a xor b);
    outputs(4238) <= not b;
    outputs(4239) <= not (a xor b);
    outputs(4240) <= a xor b;
    outputs(4241) <= a and not b;
    outputs(4242) <= b;
    outputs(4243) <= not b;
    outputs(4244) <= not (a xor b);
    outputs(4245) <= a;
    outputs(4246) <= a xor b;
    outputs(4247) <= a;
    outputs(4248) <= a xor b;
    outputs(4249) <= b and not a;
    outputs(4250) <= a;
    outputs(4251) <= b;
    outputs(4252) <= b;
    outputs(4253) <= a xor b;
    outputs(4254) <= a xor b;
    outputs(4255) <= not b;
    outputs(4256) <= b;
    outputs(4257) <= not (a xor b);
    outputs(4258) <= a xor b;
    outputs(4259) <= not a;
    outputs(4260) <= not b;
    outputs(4261) <= not (a xor b);
    outputs(4262) <= b;
    outputs(4263) <= not a or b;
    outputs(4264) <= b;
    outputs(4265) <= not (a or b);
    outputs(4266) <= a and b;
    outputs(4267) <= b and not a;
    outputs(4268) <= a;
    outputs(4269) <= not a;
    outputs(4270) <= b;
    outputs(4271) <= b and not a;
    outputs(4272) <= not (a or b);
    outputs(4273) <= not (a xor b);
    outputs(4274) <= b;
    outputs(4275) <= a xor b;
    outputs(4276) <= not (a xor b);
    outputs(4277) <= a;
    outputs(4278) <= not (a xor b);
    outputs(4279) <= not (a xor b);
    outputs(4280) <= a and not b;
    outputs(4281) <= a xor b;
    outputs(4282) <= not b;
    outputs(4283) <= not (a or b);
    outputs(4284) <= a;
    outputs(4285) <= a and b;
    outputs(4286) <= not (a xor b);
    outputs(4287) <= a;
    outputs(4288) <= b;
    outputs(4289) <= b;
    outputs(4290) <= not (a xor b);
    outputs(4291) <= not a or b;
    outputs(4292) <= b and not a;
    outputs(4293) <= a;
    outputs(4294) <= not a;
    outputs(4295) <= not a;
    outputs(4296) <= a and not b;
    outputs(4297) <= not b;
    outputs(4298) <= not (a xor b);
    outputs(4299) <= b;
    outputs(4300) <= a;
    outputs(4301) <= b;
    outputs(4302) <= a xor b;
    outputs(4303) <= not b;
    outputs(4304) <= not b or a;
    outputs(4305) <= a xor b;
    outputs(4306) <= not a;
    outputs(4307) <= a;
    outputs(4308) <= not a or b;
    outputs(4309) <= not a;
    outputs(4310) <= not a;
    outputs(4311) <= not a;
    outputs(4312) <= not b;
    outputs(4313) <= a xor b;
    outputs(4314) <= a xor b;
    outputs(4315) <= not (a xor b);
    outputs(4316) <= a xor b;
    outputs(4317) <= not (a xor b);
    outputs(4318) <= not b;
    outputs(4319) <= not b;
    outputs(4320) <= b;
    outputs(4321) <= not b;
    outputs(4322) <= a xor b;
    outputs(4323) <= not b;
    outputs(4324) <= b;
    outputs(4325) <= b;
    outputs(4326) <= a xor b;
    outputs(4327) <= not a;
    outputs(4328) <= not (a xor b);
    outputs(4329) <= not a;
    outputs(4330) <= not (a xor b);
    outputs(4331) <= a xor b;
    outputs(4332) <= not b or a;
    outputs(4333) <= b;
    outputs(4334) <= b;
    outputs(4335) <= a and b;
    outputs(4336) <= a xor b;
    outputs(4337) <= not b;
    outputs(4338) <= a or b;
    outputs(4339) <= a;
    outputs(4340) <= not b;
    outputs(4341) <= not (a xor b);
    outputs(4342) <= a and not b;
    outputs(4343) <= b;
    outputs(4344) <= a xor b;
    outputs(4345) <= a xor b;
    outputs(4346) <= a and b;
    outputs(4347) <= not (a xor b);
    outputs(4348) <= a xor b;
    outputs(4349) <= not (a xor b);
    outputs(4350) <= b and not a;
    outputs(4351) <= not b;
    outputs(4352) <= not a;
    outputs(4353) <= not a or b;
    outputs(4354) <= a xor b;
    outputs(4355) <= not a;
    outputs(4356) <= a xor b;
    outputs(4357) <= not a;
    outputs(4358) <= a;
    outputs(4359) <= b;
    outputs(4360) <= not b;
    outputs(4361) <= not b;
    outputs(4362) <= not (a xor b);
    outputs(4363) <= a xor b;
    outputs(4364) <= not (a and b);
    outputs(4365) <= b;
    outputs(4366) <= a;
    outputs(4367) <= not a or b;
    outputs(4368) <= not a or b;
    outputs(4369) <= not (a or b);
    outputs(4370) <= not (a or b);
    outputs(4371) <= a xor b;
    outputs(4372) <= a xor b;
    outputs(4373) <= not a or b;
    outputs(4374) <= b;
    outputs(4375) <= not b;
    outputs(4376) <= not a;
    outputs(4377) <= not b;
    outputs(4378) <= a;
    outputs(4379) <= a xor b;
    outputs(4380) <= b;
    outputs(4381) <= a and b;
    outputs(4382) <= not b;
    outputs(4383) <= a and b;
    outputs(4384) <= not (a xor b);
    outputs(4385) <= not b or a;
    outputs(4386) <= not (a xor b);
    outputs(4387) <= not (a xor b);
    outputs(4388) <= b;
    outputs(4389) <= a;
    outputs(4390) <= a;
    outputs(4391) <= b;
    outputs(4392) <= not a;
    outputs(4393) <= not a;
    outputs(4394) <= a xor b;
    outputs(4395) <= a xor b;
    outputs(4396) <= not (a xor b);
    outputs(4397) <= not (a xor b);
    outputs(4398) <= not (a xor b);
    outputs(4399) <= a and b;
    outputs(4400) <= b;
    outputs(4401) <= a xor b;
    outputs(4402) <= a xor b;
    outputs(4403) <= a xor b;
    outputs(4404) <= b;
    outputs(4405) <= not a;
    outputs(4406) <= a xor b;
    outputs(4407) <= a xor b;
    outputs(4408) <= b;
    outputs(4409) <= a;
    outputs(4410) <= a xor b;
    outputs(4411) <= a;
    outputs(4412) <= b;
    outputs(4413) <= not (a xor b);
    outputs(4414) <= a xor b;
    outputs(4415) <= a xor b;
    outputs(4416) <= not b or a;
    outputs(4417) <= a and b;
    outputs(4418) <= a xor b;
    outputs(4419) <= not b;
    outputs(4420) <= not a;
    outputs(4421) <= a;
    outputs(4422) <= not a;
    outputs(4423) <= a xor b;
    outputs(4424) <= not (a xor b);
    outputs(4425) <= a;
    outputs(4426) <= a;
    outputs(4427) <= not a;
    outputs(4428) <= not (a xor b);
    outputs(4429) <= not b;
    outputs(4430) <= not a;
    outputs(4431) <= not a;
    outputs(4432) <= not (a and b);
    outputs(4433) <= not b or a;
    outputs(4434) <= not (a and b);
    outputs(4435) <= not (a xor b);
    outputs(4436) <= a xor b;
    outputs(4437) <= not b;
    outputs(4438) <= not b;
    outputs(4439) <= b;
    outputs(4440) <= a or b;
    outputs(4441) <= not (a and b);
    outputs(4442) <= a;
    outputs(4443) <= not (a xor b);
    outputs(4444) <= a xor b;
    outputs(4445) <= a and b;
    outputs(4446) <= a xor b;
    outputs(4447) <= not (a xor b);
    outputs(4448) <= b and not a;
    outputs(4449) <= a xor b;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= a xor b;
    outputs(4452) <= a xor b;
    outputs(4453) <= not (a xor b);
    outputs(4454) <= not (a xor b);
    outputs(4455) <= not a or b;
    outputs(4456) <= a;
    outputs(4457) <= not (a xor b);
    outputs(4458) <= a xor b;
    outputs(4459) <= a xor b;
    outputs(4460) <= a;
    outputs(4461) <= not (a xor b);
    outputs(4462) <= not a;
    outputs(4463) <= a;
    outputs(4464) <= a and b;
    outputs(4465) <= a xor b;
    outputs(4466) <= a xor b;
    outputs(4467) <= not (a or b);
    outputs(4468) <= not a;
    outputs(4469) <= not a or b;
    outputs(4470) <= not b or a;
    outputs(4471) <= a;
    outputs(4472) <= a xor b;
    outputs(4473) <= b;
    outputs(4474) <= a or b;
    outputs(4475) <= not a;
    outputs(4476) <= b;
    outputs(4477) <= a xor b;
    outputs(4478) <= not a;
    outputs(4479) <= not (a and b);
    outputs(4480) <= not a;
    outputs(4481) <= not a;
    outputs(4482) <= a and b;
    outputs(4483) <= a xor b;
    outputs(4484) <= a xor b;
    outputs(4485) <= not b;
    outputs(4486) <= not a;
    outputs(4487) <= b and not a;
    outputs(4488) <= not (a xor b);
    outputs(4489) <= not (a xor b);
    outputs(4490) <= a xor b;
    outputs(4491) <= a or b;
    outputs(4492) <= not a;
    outputs(4493) <= not a or b;
    outputs(4494) <= b;
    outputs(4495) <= not a or b;
    outputs(4496) <= a xor b;
    outputs(4497) <= not (a xor b);
    outputs(4498) <= b;
    outputs(4499) <= a and not b;
    outputs(4500) <= not a;
    outputs(4501) <= b;
    outputs(4502) <= not (a xor b);
    outputs(4503) <= a;
    outputs(4504) <= not (a xor b);
    outputs(4505) <= not (a xor b);
    outputs(4506) <= not b;
    outputs(4507) <= a or b;
    outputs(4508) <= not a;
    outputs(4509) <= not a or b;
    outputs(4510) <= a xor b;
    outputs(4511) <= a xor b;
    outputs(4512) <= a xor b;
    outputs(4513) <= not a;
    outputs(4514) <= b;
    outputs(4515) <= a xor b;
    outputs(4516) <= a xor b;
    outputs(4517) <= not a;
    outputs(4518) <= not (a and b);
    outputs(4519) <= a;
    outputs(4520) <= not b;
    outputs(4521) <= b and not a;
    outputs(4522) <= not a;
    outputs(4523) <= not (a or b);
    outputs(4524) <= a xor b;
    outputs(4525) <= b;
    outputs(4526) <= not b;
    outputs(4527) <= a;
    outputs(4528) <= a;
    outputs(4529) <= b;
    outputs(4530) <= a;
    outputs(4531) <= a xor b;
    outputs(4532) <= not (a or b);
    outputs(4533) <= a and b;
    outputs(4534) <= a and not b;
    outputs(4535) <= a;
    outputs(4536) <= not a;
    outputs(4537) <= b;
    outputs(4538) <= not a;
    outputs(4539) <= not a;
    outputs(4540) <= a;
    outputs(4541) <= a xor b;
    outputs(4542) <= not (a or b);
    outputs(4543) <= not b or a;
    outputs(4544) <= not b;
    outputs(4545) <= not a or b;
    outputs(4546) <= a and not b;
    outputs(4547) <= a xor b;
    outputs(4548) <= b and not a;
    outputs(4549) <= not b;
    outputs(4550) <= not (a xor b);
    outputs(4551) <= not (a xor b);
    outputs(4552) <= b;
    outputs(4553) <= b;
    outputs(4554) <= not a;
    outputs(4555) <= not a;
    outputs(4556) <= a;
    outputs(4557) <= a xor b;
    outputs(4558) <= a xor b;
    outputs(4559) <= a xor b;
    outputs(4560) <= b;
    outputs(4561) <= not a or b;
    outputs(4562) <= a or b;
    outputs(4563) <= not (a or b);
    outputs(4564) <= a;
    outputs(4565) <= a and not b;
    outputs(4566) <= a xor b;
    outputs(4567) <= not (a and b);
    outputs(4568) <= not (a or b);
    outputs(4569) <= not a;
    outputs(4570) <= a xor b;
    outputs(4571) <= a;
    outputs(4572) <= a or b;
    outputs(4573) <= a;
    outputs(4574) <= not (a xor b);
    outputs(4575) <= not (a xor b);
    outputs(4576) <= a xor b;
    outputs(4577) <= b;
    outputs(4578) <= a xor b;
    outputs(4579) <= not (a xor b);
    outputs(4580) <= b;
    outputs(4581) <= a xor b;
    outputs(4582) <= not b;
    outputs(4583) <= not (a xor b);
    outputs(4584) <= a and not b;
    outputs(4585) <= a xor b;
    outputs(4586) <= not b;
    outputs(4587) <= not b;
    outputs(4588) <= b;
    outputs(4589) <= a;
    outputs(4590) <= a;
    outputs(4591) <= b;
    outputs(4592) <= b;
    outputs(4593) <= a xor b;
    outputs(4594) <= a xor b;
    outputs(4595) <= b;
    outputs(4596) <= not b;
    outputs(4597) <= b;
    outputs(4598) <= not (a or b);
    outputs(4599) <= not a;
    outputs(4600) <= not a;
    outputs(4601) <= a;
    outputs(4602) <= a xor b;
    outputs(4603) <= a xor b;
    outputs(4604) <= a xor b;
    outputs(4605) <= b;
    outputs(4606) <= not b;
    outputs(4607) <= b;
    outputs(4608) <= not (a or b);
    outputs(4609) <= a and not b;
    outputs(4610) <= not a;
    outputs(4611) <= a xor b;
    outputs(4612) <= a and not b;
    outputs(4613) <= a xor b;
    outputs(4614) <= a or b;
    outputs(4615) <= not (a xor b);
    outputs(4616) <= not b;
    outputs(4617) <= not b or a;
    outputs(4618) <= not (a xor b);
    outputs(4619) <= a xor b;
    outputs(4620) <= not (a xor b);
    outputs(4621) <= a;
    outputs(4622) <= not (a or b);
    outputs(4623) <= not a or b;
    outputs(4624) <= not a;
    outputs(4625) <= not (a xor b);
    outputs(4626) <= b;
    outputs(4627) <= not a;
    outputs(4628) <= a xor b;
    outputs(4629) <= a;
    outputs(4630) <= a and b;
    outputs(4631) <= a and not b;
    outputs(4632) <= not b;
    outputs(4633) <= not (a and b);
    outputs(4634) <= b;
    outputs(4635) <= not (a xor b);
    outputs(4636) <= not (a xor b);
    outputs(4637) <= not (a xor b);
    outputs(4638) <= a xor b;
    outputs(4639) <= not a;
    outputs(4640) <= b;
    outputs(4641) <= not (a xor b);
    outputs(4642) <= not b;
    outputs(4643) <= b and not a;
    outputs(4644) <= not (a xor b);
    outputs(4645) <= a xor b;
    outputs(4646) <= a and b;
    outputs(4647) <= b and not a;
    outputs(4648) <= a;
    outputs(4649) <= b;
    outputs(4650) <= a and b;
    outputs(4651) <= a xor b;
    outputs(4652) <= a xor b;
    outputs(4653) <= b;
    outputs(4654) <= a xor b;
    outputs(4655) <= b;
    outputs(4656) <= not b;
    outputs(4657) <= b;
    outputs(4658) <= not (a and b);
    outputs(4659) <= b;
    outputs(4660) <= not b;
    outputs(4661) <= a and b;
    outputs(4662) <= a or b;
    outputs(4663) <= a xor b;
    outputs(4664) <= b;
    outputs(4665) <= not (a xor b);
    outputs(4666) <= a xor b;
    outputs(4667) <= a xor b;
    outputs(4668) <= not b;
    outputs(4669) <= not b;
    outputs(4670) <= a and b;
    outputs(4671) <= not (a xor b);
    outputs(4672) <= a xor b;
    outputs(4673) <= not b;
    outputs(4674) <= not b;
    outputs(4675) <= b and not a;
    outputs(4676) <= not b;
    outputs(4677) <= a xor b;
    outputs(4678) <= not a;
    outputs(4679) <= not a or b;
    outputs(4680) <= not (a xor b);
    outputs(4681) <= a xor b;
    outputs(4682) <= a or b;
    outputs(4683) <= not b or a;
    outputs(4684) <= not (a xor b);
    outputs(4685) <= not b or a;
    outputs(4686) <= not b;
    outputs(4687) <= not b;
    outputs(4688) <= not (a xor b);
    outputs(4689) <= a;
    outputs(4690) <= not a;
    outputs(4691) <= not b;
    outputs(4692) <= not b;
    outputs(4693) <= b;
    outputs(4694) <= not b;
    outputs(4695) <= a and b;
    outputs(4696) <= a xor b;
    outputs(4697) <= a and b;
    outputs(4698) <= a;
    outputs(4699) <= not b;
    outputs(4700) <= b;
    outputs(4701) <= not a or b;
    outputs(4702) <= not (a xor b);
    outputs(4703) <= not a;
    outputs(4704) <= not (a or b);
    outputs(4705) <= not b or a;
    outputs(4706) <= a;
    outputs(4707) <= not b or a;
    outputs(4708) <= a xor b;
    outputs(4709) <= b;
    outputs(4710) <= a xor b;
    outputs(4711) <= a xor b;
    outputs(4712) <= a xor b;
    outputs(4713) <= not a;
    outputs(4714) <= not (a xor b);
    outputs(4715) <= a xor b;
    outputs(4716) <= not b;
    outputs(4717) <= not b;
    outputs(4718) <= not b or a;
    outputs(4719) <= not a or b;
    outputs(4720) <= not (a xor b);
    outputs(4721) <= b;
    outputs(4722) <= not (a xor b);
    outputs(4723) <= not (a xor b);
    outputs(4724) <= a xor b;
    outputs(4725) <= not (a or b);
    outputs(4726) <= a or b;
    outputs(4727) <= b;
    outputs(4728) <= not b;
    outputs(4729) <= not b;
    outputs(4730) <= a;
    outputs(4731) <= a;
    outputs(4732) <= a;
    outputs(4733) <= a xor b;
    outputs(4734) <= b;
    outputs(4735) <= a;
    outputs(4736) <= a;
    outputs(4737) <= a;
    outputs(4738) <= a;
    outputs(4739) <= not (a and b);
    outputs(4740) <= not a;
    outputs(4741) <= not (a and b);
    outputs(4742) <= not b;
    outputs(4743) <= not a or b;
    outputs(4744) <= not b;
    outputs(4745) <= not a;
    outputs(4746) <= a;
    outputs(4747) <= b;
    outputs(4748) <= a xor b;
    outputs(4749) <= a;
    outputs(4750) <= a xor b;
    outputs(4751) <= not b or a;
    outputs(4752) <= not b;
    outputs(4753) <= b;
    outputs(4754) <= a and b;
    outputs(4755) <= a xor b;
    outputs(4756) <= a and not b;
    outputs(4757) <= b;
    outputs(4758) <= a;
    outputs(4759) <= b;
    outputs(4760) <= a and b;
    outputs(4761) <= not b;
    outputs(4762) <= a xor b;
    outputs(4763) <= a;
    outputs(4764) <= not b;
    outputs(4765) <= a and not b;
    outputs(4766) <= a and not b;
    outputs(4767) <= not b;
    outputs(4768) <= not b;
    outputs(4769) <= not a;
    outputs(4770) <= not (a or b);
    outputs(4771) <= a xor b;
    outputs(4772) <= a;
    outputs(4773) <= a xor b;
    outputs(4774) <= a xor b;
    outputs(4775) <= not (a xor b);
    outputs(4776) <= not a;
    outputs(4777) <= not a;
    outputs(4778) <= a;
    outputs(4779) <= not (a xor b);
    outputs(4780) <= not b;
    outputs(4781) <= not b;
    outputs(4782) <= a xor b;
    outputs(4783) <= not (a xor b);
    outputs(4784) <= not a;
    outputs(4785) <= a and b;
    outputs(4786) <= not (a xor b);
    outputs(4787) <= not a;
    outputs(4788) <= not (a xor b);
    outputs(4789) <= not (a xor b);
    outputs(4790) <= b;
    outputs(4791) <= not (a xor b);
    outputs(4792) <= not (a xor b);
    outputs(4793) <= not a;
    outputs(4794) <= a xor b;
    outputs(4795) <= not a;
    outputs(4796) <= a;
    outputs(4797) <= not (a xor b);
    outputs(4798) <= b;
    outputs(4799) <= not a;
    outputs(4800) <= a xor b;
    outputs(4801) <= b and not a;
    outputs(4802) <= a xor b;
    outputs(4803) <= a xor b;
    outputs(4804) <= a or b;
    outputs(4805) <= a or b;
    outputs(4806) <= a xor b;
    outputs(4807) <= a and not b;
    outputs(4808) <= not (a xor b);
    outputs(4809) <= a;
    outputs(4810) <= a xor b;
    outputs(4811) <= b;
    outputs(4812) <= not b;
    outputs(4813) <= not a;
    outputs(4814) <= not (a xor b);
    outputs(4815) <= not (a xor b);
    outputs(4816) <= a and not b;
    outputs(4817) <= b;
    outputs(4818) <= b;
    outputs(4819) <= not (a xor b);
    outputs(4820) <= not a;
    outputs(4821) <= b;
    outputs(4822) <= not (a xor b);
    outputs(4823) <= b;
    outputs(4824) <= a xor b;
    outputs(4825) <= not b or a;
    outputs(4826) <= a and b;
    outputs(4827) <= a xor b;
    outputs(4828) <= a xor b;
    outputs(4829) <= a and b;
    outputs(4830) <= b;
    outputs(4831) <= not b;
    outputs(4832) <= a;
    outputs(4833) <= b;
    outputs(4834) <= a;
    outputs(4835) <= not (a xor b);
    outputs(4836) <= not (a xor b);
    outputs(4837) <= a xor b;
    outputs(4838) <= a or b;
    outputs(4839) <= a;
    outputs(4840) <= a xor b;
    outputs(4841) <= not b;
    outputs(4842) <= not (a xor b);
    outputs(4843) <= not b;
    outputs(4844) <= not b;
    outputs(4845) <= a xor b;
    outputs(4846) <= a and b;
    outputs(4847) <= a and b;
    outputs(4848) <= a xor b;
    outputs(4849) <= a or b;
    outputs(4850) <= not (a and b);
    outputs(4851) <= not b;
    outputs(4852) <= not (a or b);
    outputs(4853) <= a and b;
    outputs(4854) <= not b;
    outputs(4855) <= a xor b;
    outputs(4856) <= not (a xor b);
    outputs(4857) <= not a;
    outputs(4858) <= a;
    outputs(4859) <= b;
    outputs(4860) <= a and not b;
    outputs(4861) <= b;
    outputs(4862) <= a or b;
    outputs(4863) <= a;
    outputs(4864) <= a xor b;
    outputs(4865) <= b;
    outputs(4866) <= a;
    outputs(4867) <= a and not b;
    outputs(4868) <= a xor b;
    outputs(4869) <= a and not b;
    outputs(4870) <= not (a xor b);
    outputs(4871) <= not a;
    outputs(4872) <= a;
    outputs(4873) <= a xor b;
    outputs(4874) <= not a;
    outputs(4875) <= a xor b;
    outputs(4876) <= not (a or b);
    outputs(4877) <= not (a xor b);
    outputs(4878) <= a xor b;
    outputs(4879) <= not (a xor b);
    outputs(4880) <= not (a xor b);
    outputs(4881) <= not a or b;
    outputs(4882) <= not b;
    outputs(4883) <= not b;
    outputs(4884) <= not (a xor b);
    outputs(4885) <= b;
    outputs(4886) <= b and not a;
    outputs(4887) <= not (a and b);
    outputs(4888) <= not a;
    outputs(4889) <= a;
    outputs(4890) <= not (a and b);
    outputs(4891) <= not a;
    outputs(4892) <= not a;
    outputs(4893) <= a xor b;
    outputs(4894) <= a xor b;
    outputs(4895) <= not a;
    outputs(4896) <= b;
    outputs(4897) <= b;
    outputs(4898) <= a or b;
    outputs(4899) <= not b;
    outputs(4900) <= a xor b;
    outputs(4901) <= a xor b;
    outputs(4902) <= b;
    outputs(4903) <= not (a or b);
    outputs(4904) <= a;
    outputs(4905) <= b;
    outputs(4906) <= not (a xor b);
    outputs(4907) <= not a;
    outputs(4908) <= a xor b;
    outputs(4909) <= not (a xor b);
    outputs(4910) <= a and not b;
    outputs(4911) <= not b;
    outputs(4912) <= not (a xor b);
    outputs(4913) <= a xor b;
    outputs(4914) <= not a;
    outputs(4915) <= not (a xor b);
    outputs(4916) <= not a;
    outputs(4917) <= not a or b;
    outputs(4918) <= a;
    outputs(4919) <= not (a xor b);
    outputs(4920) <= not (a xor b);
    outputs(4921) <= not a;
    outputs(4922) <= not a or b;
    outputs(4923) <= a xor b;
    outputs(4924) <= not a;
    outputs(4925) <= not a;
    outputs(4926) <= a and b;
    outputs(4927) <= not b;
    outputs(4928) <= a and b;
    outputs(4929) <= not a;
    outputs(4930) <= not (a and b);
    outputs(4931) <= a and not b;
    outputs(4932) <= a xor b;
    outputs(4933) <= b;
    outputs(4934) <= not (a xor b);
    outputs(4935) <= not b;
    outputs(4936) <= a xor b;
    outputs(4937) <= not a;
    outputs(4938) <= b;
    outputs(4939) <= not a;
    outputs(4940) <= a xor b;
    outputs(4941) <= not (a and b);
    outputs(4942) <= not (a xor b);
    outputs(4943) <= not (a xor b);
    outputs(4944) <= a and b;
    outputs(4945) <= not a;
    outputs(4946) <= a;
    outputs(4947) <= b and not a;
    outputs(4948) <= not b;
    outputs(4949) <= a or b;
    outputs(4950) <= not a;
    outputs(4951) <= a and b;
    outputs(4952) <= not a or b;
    outputs(4953) <= a xor b;
    outputs(4954) <= a or b;
    outputs(4955) <= a or b;
    outputs(4956) <= not b;
    outputs(4957) <= a xor b;
    outputs(4958) <= not (a xor b);
    outputs(4959) <= not a or b;
    outputs(4960) <= not a;
    outputs(4961) <= a;
    outputs(4962) <= not b or a;
    outputs(4963) <= a xor b;
    outputs(4964) <= not b;
    outputs(4965) <= a;
    outputs(4966) <= a xor b;
    outputs(4967) <= b and not a;
    outputs(4968) <= not a;
    outputs(4969) <= b and not a;
    outputs(4970) <= not (a and b);
    outputs(4971) <= not a;
    outputs(4972) <= a;
    outputs(4973) <= not b;
    outputs(4974) <= b;
    outputs(4975) <= not (a xor b);
    outputs(4976) <= not a or b;
    outputs(4977) <= a or b;
    outputs(4978) <= a xor b;
    outputs(4979) <= b and not a;
    outputs(4980) <= not b;
    outputs(4981) <= not a;
    outputs(4982) <= a or b;
    outputs(4983) <= a xor b;
    outputs(4984) <= b;
    outputs(4985) <= a xor b;
    outputs(4986) <= b;
    outputs(4987) <= b;
    outputs(4988) <= a xor b;
    outputs(4989) <= not (a xor b);
    outputs(4990) <= a xor b;
    outputs(4991) <= a;
    outputs(4992) <= a;
    outputs(4993) <= b;
    outputs(4994) <= not (a xor b);
    outputs(4995) <= a xor b;
    outputs(4996) <= not b;
    outputs(4997) <= not (a xor b);
    outputs(4998) <= b;
    outputs(4999) <= not (a xor b);
    outputs(5000) <= not b;
    outputs(5001) <= a and b;
    outputs(5002) <= not a;
    outputs(5003) <= not (a xor b);
    outputs(5004) <= a xor b;
    outputs(5005) <= a and not b;
    outputs(5006) <= a;
    outputs(5007) <= not (a xor b);
    outputs(5008) <= not a;
    outputs(5009) <= a;
    outputs(5010) <= not (a xor b);
    outputs(5011) <= not (a xor b);
    outputs(5012) <= not (a or b);
    outputs(5013) <= a;
    outputs(5014) <= not (a xor b);
    outputs(5015) <= b;
    outputs(5016) <= not (a xor b);
    outputs(5017) <= b;
    outputs(5018) <= a;
    outputs(5019) <= a xor b;
    outputs(5020) <= a xor b;
    outputs(5021) <= b and not a;
    outputs(5022) <= a;
    outputs(5023) <= not b;
    outputs(5024) <= b;
    outputs(5025) <= not b;
    outputs(5026) <= b;
    outputs(5027) <= not a;
    outputs(5028) <= b;
    outputs(5029) <= b;
    outputs(5030) <= not (a and b);
    outputs(5031) <= not a or b;
    outputs(5032) <= not b;
    outputs(5033) <= not (a or b);
    outputs(5034) <= b and not a;
    outputs(5035) <= b;
    outputs(5036) <= a and not b;
    outputs(5037) <= not (a and b);
    outputs(5038) <= not (a and b);
    outputs(5039) <= not (a or b);
    outputs(5040) <= a;
    outputs(5041) <= not (a xor b);
    outputs(5042) <= a;
    outputs(5043) <= not (a or b);
    outputs(5044) <= not (a xor b);
    outputs(5045) <= not a;
    outputs(5046) <= not a;
    outputs(5047) <= a xor b;
    outputs(5048) <= not b;
    outputs(5049) <= a;
    outputs(5050) <= a or b;
    outputs(5051) <= not (a xor b);
    outputs(5052) <= not b;
    outputs(5053) <= not (a xor b);
    outputs(5054) <= a xor b;
    outputs(5055) <= not b;
    outputs(5056) <= not a;
    outputs(5057) <= b;
    outputs(5058) <= not (a xor b);
    outputs(5059) <= not (a or b);
    outputs(5060) <= a xor b;
    outputs(5061) <= b;
    outputs(5062) <= not b;
    outputs(5063) <= a xor b;
    outputs(5064) <= not b;
    outputs(5065) <= a xor b;
    outputs(5066) <= not b or a;
    outputs(5067) <= not (a xor b);
    outputs(5068) <= not (a xor b);
    outputs(5069) <= b;
    outputs(5070) <= a;
    outputs(5071) <= a and not b;
    outputs(5072) <= not (a xor b);
    outputs(5073) <= b;
    outputs(5074) <= b;
    outputs(5075) <= b;
    outputs(5076) <= a and b;
    outputs(5077) <= b;
    outputs(5078) <= not a;
    outputs(5079) <= a xor b;
    outputs(5080) <= a xor b;
    outputs(5081) <= not b;
    outputs(5082) <= not (a xor b);
    outputs(5083) <= a xor b;
    outputs(5084) <= not (a xor b);
    outputs(5085) <= not (a or b);
    outputs(5086) <= not b;
    outputs(5087) <= not b;
    outputs(5088) <= a or b;
    outputs(5089) <= b and not a;
    outputs(5090) <= a;
    outputs(5091) <= not (a or b);
    outputs(5092) <= b;
    outputs(5093) <= not b;
    outputs(5094) <= not (a xor b);
    outputs(5095) <= not b or a;
    outputs(5096) <= not (a and b);
    outputs(5097) <= not (a xor b);
    outputs(5098) <= not b;
    outputs(5099) <= a xor b;
    outputs(5100) <= not (a or b);
    outputs(5101) <= not (a xor b);
    outputs(5102) <= not (a xor b);
    outputs(5103) <= not (a xor b);
    outputs(5104) <= a xor b;
    outputs(5105) <= b;
    outputs(5106) <= not b or a;
    outputs(5107) <= a xor b;
    outputs(5108) <= b;
    outputs(5109) <= a xor b;
    outputs(5110) <= a and b;
    outputs(5111) <= not (a and b);
    outputs(5112) <= not (a xor b);
    outputs(5113) <= not (a xor b);
    outputs(5114) <= not a;
    outputs(5115) <= a;
    outputs(5116) <= not (a or b);
    outputs(5117) <= b;
    outputs(5118) <= a xor b;
    outputs(5119) <= a and not b;
    outputs(5120) <= a and not b;
    outputs(5121) <= not b;
    outputs(5122) <= not a;
    outputs(5123) <= a and b;
    outputs(5124) <= not a;
    outputs(5125) <= not (a xor b);
    outputs(5126) <= not b;
    outputs(5127) <= b;
    outputs(5128) <= a xor b;
    outputs(5129) <= a;
    outputs(5130) <= not a or b;
    outputs(5131) <= not (a xor b);
    outputs(5132) <= not b or a;
    outputs(5133) <= a xor b;
    outputs(5134) <= not (a xor b);
    outputs(5135) <= b;
    outputs(5136) <= a xor b;
    outputs(5137) <= not (a xor b);
    outputs(5138) <= not a;
    outputs(5139) <= a and b;
    outputs(5140) <= a;
    outputs(5141) <= b;
    outputs(5142) <= not a;
    outputs(5143) <= a xor b;
    outputs(5144) <= a and not b;
    outputs(5145) <= a xor b;
    outputs(5146) <= not (a xor b);
    outputs(5147) <= not (a xor b);
    outputs(5148) <= not b;
    outputs(5149) <= a;
    outputs(5150) <= a and b;
    outputs(5151) <= not b;
    outputs(5152) <= not b;
    outputs(5153) <= b;
    outputs(5154) <= a;
    outputs(5155) <= not (a xor b);
    outputs(5156) <= not (a and b);
    outputs(5157) <= a and b;
    outputs(5158) <= not (a xor b);
    outputs(5159) <= a and not b;
    outputs(5160) <= a xor b;
    outputs(5161) <= not a;
    outputs(5162) <= b;
    outputs(5163) <= not (a xor b);
    outputs(5164) <= not b;
    outputs(5165) <= not a;
    outputs(5166) <= not a;
    outputs(5167) <= a xor b;
    outputs(5168) <= b and not a;
    outputs(5169) <= a;
    outputs(5170) <= not (a or b);
    outputs(5171) <= not b;
    outputs(5172) <= not a;
    outputs(5173) <= a xor b;
    outputs(5174) <= not a;
    outputs(5175) <= not a;
    outputs(5176) <= a;
    outputs(5177) <= a;
    outputs(5178) <= b;
    outputs(5179) <= a and b;
    outputs(5180) <= b and not a;
    outputs(5181) <= a or b;
    outputs(5182) <= not b;
    outputs(5183) <= b and not a;
    outputs(5184) <= a xor b;
    outputs(5185) <= a;
    outputs(5186) <= not b;
    outputs(5187) <= not (a xor b);
    outputs(5188) <= b and not a;
    outputs(5189) <= a;
    outputs(5190) <= b;
    outputs(5191) <= a xor b;
    outputs(5192) <= not b or a;
    outputs(5193) <= a and not b;
    outputs(5194) <= not a or b;
    outputs(5195) <= a xor b;
    outputs(5196) <= a;
    outputs(5197) <= b;
    outputs(5198) <= a;
    outputs(5199) <= b and not a;
    outputs(5200) <= a xor b;
    outputs(5201) <= not a;
    outputs(5202) <= a and b;
    outputs(5203) <= a or b;
    outputs(5204) <= not b or a;
    outputs(5205) <= a xor b;
    outputs(5206) <= not b;
    outputs(5207) <= a;
    outputs(5208) <= not (a xor b);
    outputs(5209) <= a xor b;
    outputs(5210) <= not (a xor b);
    outputs(5211) <= a;
    outputs(5212) <= a;
    outputs(5213) <= b;
    outputs(5214) <= not (a xor b);
    outputs(5215) <= a xor b;
    outputs(5216) <= b;
    outputs(5217) <= not a;
    outputs(5218) <= a xor b;
    outputs(5219) <= a xor b;
    outputs(5220) <= not (a xor b);
    outputs(5221) <= not (a xor b);
    outputs(5222) <= not a;
    outputs(5223) <= b;
    outputs(5224) <= a;
    outputs(5225) <= a xor b;
    outputs(5226) <= b;
    outputs(5227) <= a xor b;
    outputs(5228) <= a xor b;
    outputs(5229) <= b;
    outputs(5230) <= a or b;
    outputs(5231) <= not (a xor b);
    outputs(5232) <= not (a xor b);
    outputs(5233) <= not a;
    outputs(5234) <= not b or a;
    outputs(5235) <= a;
    outputs(5236) <= not (a or b);
    outputs(5237) <= a and not b;
    outputs(5238) <= not b or a;
    outputs(5239) <= not a;
    outputs(5240) <= not (a xor b);
    outputs(5241) <= a and not b;
    outputs(5242) <= a xor b;
    outputs(5243) <= not b or a;
    outputs(5244) <= not a;
    outputs(5245) <= not b or a;
    outputs(5246) <= a xor b;
    outputs(5247) <= b;
    outputs(5248) <= not (a xor b);
    outputs(5249) <= not b or a;
    outputs(5250) <= b;
    outputs(5251) <= not b;
    outputs(5252) <= not (a xor b);
    outputs(5253) <= not (a xor b);
    outputs(5254) <= not (a or b);
    outputs(5255) <= a;
    outputs(5256) <= not a;
    outputs(5257) <= not (a or b);
    outputs(5258) <= a xor b;
    outputs(5259) <= a xor b;
    outputs(5260) <= a and not b;
    outputs(5261) <= a and b;
    outputs(5262) <= b;
    outputs(5263) <= a;
    outputs(5264) <= not b or a;
    outputs(5265) <= a xor b;
    outputs(5266) <= not a;
    outputs(5267) <= not b;
    outputs(5268) <= b;
    outputs(5269) <= not b or a;
    outputs(5270) <= not b;
    outputs(5271) <= not (a xor b);
    outputs(5272) <= a xor b;
    outputs(5273) <= not a;
    outputs(5274) <= b;
    outputs(5275) <= a and not b;
    outputs(5276) <= not (a or b);
    outputs(5277) <= a and not b;
    outputs(5278) <= not a;
    outputs(5279) <= not b or a;
    outputs(5280) <= not a;
    outputs(5281) <= b;
    outputs(5282) <= not b;
    outputs(5283) <= a xor b;
    outputs(5284) <= a xor b;
    outputs(5285) <= not b or a;
    outputs(5286) <= a and b;
    outputs(5287) <= a xor b;
    outputs(5288) <= a;
    outputs(5289) <= a xor b;
    outputs(5290) <= b;
    outputs(5291) <= b;
    outputs(5292) <= not a;
    outputs(5293) <= a xor b;
    outputs(5294) <= b and not a;
    outputs(5295) <= a and not b;
    outputs(5296) <= b;
    outputs(5297) <= not (a xor b);
    outputs(5298) <= a xor b;
    outputs(5299) <= a;
    outputs(5300) <= a and b;
    outputs(5301) <= not b or a;
    outputs(5302) <= a;
    outputs(5303) <= a and b;
    outputs(5304) <= not b;
    outputs(5305) <= b;
    outputs(5306) <= a;
    outputs(5307) <= not (a xor b);
    outputs(5308) <= a or b;
    outputs(5309) <= a;
    outputs(5310) <= not a;
    outputs(5311) <= not (a xor b);
    outputs(5312) <= a xor b;
    outputs(5313) <= a or b;
    outputs(5314) <= not (a xor b);
    outputs(5315) <= not (a xor b);
    outputs(5316) <= a and b;
    outputs(5317) <= not b;
    outputs(5318) <= a and not b;
    outputs(5319) <= not (a or b);
    outputs(5320) <= a and not b;
    outputs(5321) <= a;
    outputs(5322) <= not a;
    outputs(5323) <= b;
    outputs(5324) <= not a;
    outputs(5325) <= not (a or b);
    outputs(5326) <= a xor b;
    outputs(5327) <= not (a xor b);
    outputs(5328) <= a;
    outputs(5329) <= not (a xor b);
    outputs(5330) <= not (a xor b);
    outputs(5331) <= a and not b;
    outputs(5332) <= a;
    outputs(5333) <= not b;
    outputs(5334) <= b;
    outputs(5335) <= not a;
    outputs(5336) <= not a;
    outputs(5337) <= a and b;
    outputs(5338) <= not b;
    outputs(5339) <= not b;
    outputs(5340) <= a xor b;
    outputs(5341) <= not b or a;
    outputs(5342) <= not a;
    outputs(5343) <= a xor b;
    outputs(5344) <= not (a xor b);
    outputs(5345) <= not b;
    outputs(5346) <= a;
    outputs(5347) <= a xor b;
    outputs(5348) <= not a;
    outputs(5349) <= not a;
    outputs(5350) <= a or b;
    outputs(5351) <= not (a xor b);
    outputs(5352) <= b;
    outputs(5353) <= a and b;
    outputs(5354) <= not (a xor b);
    outputs(5355) <= b;
    outputs(5356) <= not (a xor b);
    outputs(5357) <= not (a xor b);
    outputs(5358) <= not b;
    outputs(5359) <= a;
    outputs(5360) <= a xor b;
    outputs(5361) <= not a;
    outputs(5362) <= a or b;
    outputs(5363) <= not b;
    outputs(5364) <= a and not b;
    outputs(5365) <= b;
    outputs(5366) <= b;
    outputs(5367) <= b;
    outputs(5368) <= a xor b;
    outputs(5369) <= b;
    outputs(5370) <= a xor b;
    outputs(5371) <= a;
    outputs(5372) <= not a;
    outputs(5373) <= a xor b;
    outputs(5374) <= not b;
    outputs(5375) <= not (a xor b);
    outputs(5376) <= b;
    outputs(5377) <= b;
    outputs(5378) <= not b;
    outputs(5379) <= b and not a;
    outputs(5380) <= a xor b;
    outputs(5381) <= not b;
    outputs(5382) <= a and b;
    outputs(5383) <= b;
    outputs(5384) <= not b;
    outputs(5385) <= not a or b;
    outputs(5386) <= a xor b;
    outputs(5387) <= not b;
    outputs(5388) <= not (a xor b);
    outputs(5389) <= not a;
    outputs(5390) <= not b;
    outputs(5391) <= not a;
    outputs(5392) <= not (a xor b);
    outputs(5393) <= not a;
    outputs(5394) <= a xor b;
    outputs(5395) <= a xor b;
    outputs(5396) <= a xor b;
    outputs(5397) <= not (a and b);
    outputs(5398) <= not b;
    outputs(5399) <= not a;
    outputs(5400) <= a;
    outputs(5401) <= a;
    outputs(5402) <= a xor b;
    outputs(5403) <= a and b;
    outputs(5404) <= not a;
    outputs(5405) <= not (a and b);
    outputs(5406) <= b;
    outputs(5407) <= not b;
    outputs(5408) <= not (a or b);
    outputs(5409) <= a;
    outputs(5410) <= b;
    outputs(5411) <= not (a or b);
    outputs(5412) <= a;
    outputs(5413) <= not b;
    outputs(5414) <= not b;
    outputs(5415) <= b;
    outputs(5416) <= a and b;
    outputs(5417) <= not (a xor b);
    outputs(5418) <= not a;
    outputs(5419) <= not (a xor b);
    outputs(5420) <= a xor b;
    outputs(5421) <= not a;
    outputs(5422) <= b;
    outputs(5423) <= not b;
    outputs(5424) <= b;
    outputs(5425) <= a xor b;
    outputs(5426) <= a and b;
    outputs(5427) <= b;
    outputs(5428) <= not (a xor b);
    outputs(5429) <= b;
    outputs(5430) <= a xor b;
    outputs(5431) <= a xor b;
    outputs(5432) <= not (a or b);
    outputs(5433) <= b;
    outputs(5434) <= a;
    outputs(5435) <= a;
    outputs(5436) <= a xor b;
    outputs(5437) <= not b or a;
    outputs(5438) <= not a;
    outputs(5439) <= not b;
    outputs(5440) <= a;
    outputs(5441) <= a xor b;
    outputs(5442) <= b and not a;
    outputs(5443) <= not a or b;
    outputs(5444) <= not a;
    outputs(5445) <= a and b;
    outputs(5446) <= not b;
    outputs(5447) <= not (a xor b);
    outputs(5448) <= not b;
    outputs(5449) <= not (a xor b);
    outputs(5450) <= a xor b;
    outputs(5451) <= not a;
    outputs(5452) <= not a or b;
    outputs(5453) <= b and not a;
    outputs(5454) <= a;
    outputs(5455) <= not (a xor b);
    outputs(5456) <= b;
    outputs(5457) <= a;
    outputs(5458) <= not b or a;
    outputs(5459) <= a;
    outputs(5460) <= not a or b;
    outputs(5461) <= not a;
    outputs(5462) <= b and not a;
    outputs(5463) <= a;
    outputs(5464) <= not a;
    outputs(5465) <= not (a xor b);
    outputs(5466) <= a;
    outputs(5467) <= a and not b;
    outputs(5468) <= not (a and b);
    outputs(5469) <= not b or a;
    outputs(5470) <= a xor b;
    outputs(5471) <= not b;
    outputs(5472) <= not a or b;
    outputs(5473) <= not (a xor b);
    outputs(5474) <= a xor b;
    outputs(5475) <= not a or b;
    outputs(5476) <= not b or a;
    outputs(5477) <= not a;
    outputs(5478) <= not a;
    outputs(5479) <= not b;
    outputs(5480) <= not (a xor b);
    outputs(5481) <= b;
    outputs(5482) <= not a;
    outputs(5483) <= not b;
    outputs(5484) <= not b;
    outputs(5485) <= not b;
    outputs(5486) <= not b;
    outputs(5487) <= a and not b;
    outputs(5488) <= not a;
    outputs(5489) <= not (a or b);
    outputs(5490) <= a xor b;
    outputs(5491) <= not a;
    outputs(5492) <= not (a xor b);
    outputs(5493) <= a or b;
    outputs(5494) <= b;
    outputs(5495) <= b;
    outputs(5496) <= a and not b;
    outputs(5497) <= b;
    outputs(5498) <= not b;
    outputs(5499) <= b;
    outputs(5500) <= not b;
    outputs(5501) <= a and not b;
    outputs(5502) <= b;
    outputs(5503) <= not a;
    outputs(5504) <= a xor b;
    outputs(5505) <= b;
    outputs(5506) <= not a;
    outputs(5507) <= not (a and b);
    outputs(5508) <= b and not a;
    outputs(5509) <= a;
    outputs(5510) <= a xor b;
    outputs(5511) <= not b;
    outputs(5512) <= not (a xor b);
    outputs(5513) <= not a;
    outputs(5514) <= not a;
    outputs(5515) <= not (a xor b);
    outputs(5516) <= not (a or b);
    outputs(5517) <= a;
    outputs(5518) <= a xor b;
    outputs(5519) <= not (a xor b);
    outputs(5520) <= b and not a;
    outputs(5521) <= not b;
    outputs(5522) <= a;
    outputs(5523) <= not (a or b);
    outputs(5524) <= a xor b;
    outputs(5525) <= b;
    outputs(5526) <= not (a xor b);
    outputs(5527) <= a xor b;
    outputs(5528) <= a and b;
    outputs(5529) <= not b;
    outputs(5530) <= a and not b;
    outputs(5531) <= not (a xor b);
    outputs(5532) <= not a;
    outputs(5533) <= not b;
    outputs(5534) <= not a;
    outputs(5535) <= a xor b;
    outputs(5536) <= b;
    outputs(5537) <= b;
    outputs(5538) <= not (a or b);
    outputs(5539) <= a and not b;
    outputs(5540) <= not b;
    outputs(5541) <= a or b;
    outputs(5542) <= not a;
    outputs(5543) <= b and not a;
    outputs(5544) <= not (a xor b);
    outputs(5545) <= a and b;
    outputs(5546) <= not (a xor b);
    outputs(5547) <= b;
    outputs(5548) <= a and not b;
    outputs(5549) <= not b;
    outputs(5550) <= a xor b;
    outputs(5551) <= a xor b;
    outputs(5552) <= not b;
    outputs(5553) <= a xor b;
    outputs(5554) <= not b;
    outputs(5555) <= a xor b;
    outputs(5556) <= b and not a;
    outputs(5557) <= a;
    outputs(5558) <= not b or a;
    outputs(5559) <= b;
    outputs(5560) <= a or b;
    outputs(5561) <= a xor b;
    outputs(5562) <= not (a xor b);
    outputs(5563) <= b;
    outputs(5564) <= a xor b;
    outputs(5565) <= not (a xor b);
    outputs(5566) <= not (a and b);
    outputs(5567) <= not b;
    outputs(5568) <= not a or b;
    outputs(5569) <= not b;
    outputs(5570) <= not (a xor b);
    outputs(5571) <= a;
    outputs(5572) <= not a;
    outputs(5573) <= not a;
    outputs(5574) <= not a;
    outputs(5575) <= not (a and b);
    outputs(5576) <= not a;
    outputs(5577) <= a and b;
    outputs(5578) <= a xor b;
    outputs(5579) <= not (a xor b);
    outputs(5580) <= not b;
    outputs(5581) <= a;
    outputs(5582) <= not a;
    outputs(5583) <= a;
    outputs(5584) <= not (a or b);
    outputs(5585) <= a;
    outputs(5586) <= not (a xor b);
    outputs(5587) <= b;
    outputs(5588) <= not a or b;
    outputs(5589) <= not (a xor b);
    outputs(5590) <= not a;
    outputs(5591) <= a or b;
    outputs(5592) <= not (a xor b);
    outputs(5593) <= b;
    outputs(5594) <= not b;
    outputs(5595) <= b;
    outputs(5596) <= a and not b;
    outputs(5597) <= a and not b;
    outputs(5598) <= a and not b;
    outputs(5599) <= a;
    outputs(5600) <= a and b;
    outputs(5601) <= a xor b;
    outputs(5602) <= a xor b;
    outputs(5603) <= a xor b;
    outputs(5604) <= not (a and b);
    outputs(5605) <= a or b;
    outputs(5606) <= not (a xor b);
    outputs(5607) <= not b;
    outputs(5608) <= not a;
    outputs(5609) <= a;
    outputs(5610) <= b;
    outputs(5611) <= not a;
    outputs(5612) <= a;
    outputs(5613) <= not b or a;
    outputs(5614) <= a;
    outputs(5615) <= not a;
    outputs(5616) <= not (a xor b);
    outputs(5617) <= a and b;
    outputs(5618) <= b;
    outputs(5619) <= not a;
    outputs(5620) <= a;
    outputs(5621) <= a and not b;
    outputs(5622) <= a xor b;
    outputs(5623) <= a and b;
    outputs(5624) <= a;
    outputs(5625) <= a and not b;
    outputs(5626) <= not a;
    outputs(5627) <= b;
    outputs(5628) <= a xor b;
    outputs(5629) <= a;
    outputs(5630) <= not (a or b);
    outputs(5631) <= not (a xor b);
    outputs(5632) <= not a;
    outputs(5633) <= a xor b;
    outputs(5634) <= a and b;
    outputs(5635) <= a xor b;
    outputs(5636) <= a;
    outputs(5637) <= b;
    outputs(5638) <= not (a and b);
    outputs(5639) <= not a;
    outputs(5640) <= a xor b;
    outputs(5641) <= a xor b;
    outputs(5642) <= b;
    outputs(5643) <= b;
    outputs(5644) <= not (a xor b);
    outputs(5645) <= not (a xor b);
    outputs(5646) <= a and not b;
    outputs(5647) <= b;
    outputs(5648) <= not (a or b);
    outputs(5649) <= not (a xor b);
    outputs(5650) <= not b;
    outputs(5651) <= not b or a;
    outputs(5652) <= not a;
    outputs(5653) <= not b;
    outputs(5654) <= a xor b;
    outputs(5655) <= a and b;
    outputs(5656) <= a;
    outputs(5657) <= not b;
    outputs(5658) <= b;
    outputs(5659) <= not a;
    outputs(5660) <= a and not b;
    outputs(5661) <= not b or a;
    outputs(5662) <= not (a xor b);
    outputs(5663) <= not b or a;
    outputs(5664) <= a and not b;
    outputs(5665) <= not a;
    outputs(5666) <= b;
    outputs(5667) <= a xor b;
    outputs(5668) <= not b;
    outputs(5669) <= a xor b;
    outputs(5670) <= not b;
    outputs(5671) <= a and b;
    outputs(5672) <= not b;
    outputs(5673) <= not (a and b);
    outputs(5674) <= not b;
    outputs(5675) <= not a;
    outputs(5676) <= not a or b;
    outputs(5677) <= b;
    outputs(5678) <= not b;
    outputs(5679) <= a xor b;
    outputs(5680) <= not a;
    outputs(5681) <= a;
    outputs(5682) <= not (a xor b);
    outputs(5683) <= a;
    outputs(5684) <= a;
    outputs(5685) <= not b;
    outputs(5686) <= a and b;
    outputs(5687) <= not (a xor b);
    outputs(5688) <= not b;
    outputs(5689) <= a xor b;
    outputs(5690) <= b;
    outputs(5691) <= not a;
    outputs(5692) <= a xor b;
    outputs(5693) <= b;
    outputs(5694) <= b;
    outputs(5695) <= a;
    outputs(5696) <= not a;
    outputs(5697) <= a;
    outputs(5698) <= not b or a;
    outputs(5699) <= a xor b;
    outputs(5700) <= not (a and b);
    outputs(5701) <= a;
    outputs(5702) <= a and not b;
    outputs(5703) <= a and b;
    outputs(5704) <= not a;
    outputs(5705) <= a or b;
    outputs(5706) <= a;
    outputs(5707) <= not (a or b);
    outputs(5708) <= a or b;
    outputs(5709) <= not a;
    outputs(5710) <= not a or b;
    outputs(5711) <= not a;
    outputs(5712) <= not b;
    outputs(5713) <= b;
    outputs(5714) <= not b;
    outputs(5715) <= a xor b;
    outputs(5716) <= not a or b;
    outputs(5717) <= not (a or b);
    outputs(5718) <= not (a xor b);
    outputs(5719) <= not b;
    outputs(5720) <= b;
    outputs(5721) <= not (a or b);
    outputs(5722) <= not b;
    outputs(5723) <= a and b;
    outputs(5724) <= not (a xor b);
    outputs(5725) <= a;
    outputs(5726) <= a xor b;
    outputs(5727) <= a;
    outputs(5728) <= a and b;
    outputs(5729) <= not (a xor b);
    outputs(5730) <= a;
    outputs(5731) <= b;
    outputs(5732) <= not a or b;
    outputs(5733) <= not b;
    outputs(5734) <= not a;
    outputs(5735) <= a;
    outputs(5736) <= not a;
    outputs(5737) <= b;
    outputs(5738) <= b and not a;
    outputs(5739) <= not (a xor b);
    outputs(5740) <= a xor b;
    outputs(5741) <= a;
    outputs(5742) <= a;
    outputs(5743) <= a xor b;
    outputs(5744) <= a;
    outputs(5745) <= not a;
    outputs(5746) <= not a;
    outputs(5747) <= a or b;
    outputs(5748) <= not a or b;
    outputs(5749) <= not a;
    outputs(5750) <= b;
    outputs(5751) <= not (a xor b);
    outputs(5752) <= a xor b;
    outputs(5753) <= not (a xor b);
    outputs(5754) <= a xor b;
    outputs(5755) <= a;
    outputs(5756) <= a xor b;
    outputs(5757) <= not b;
    outputs(5758) <= a;
    outputs(5759) <= b;
    outputs(5760) <= a and not b;
    outputs(5761) <= a and not b;
    outputs(5762) <= a and not b;
    outputs(5763) <= a;
    outputs(5764) <= not (a or b);
    outputs(5765) <= not (a or b);
    outputs(5766) <= b;
    outputs(5767) <= b;
    outputs(5768) <= not (a xor b);
    outputs(5769) <= b;
    outputs(5770) <= a;
    outputs(5771) <= not (a and b);
    outputs(5772) <= not b;
    outputs(5773) <= a and b;
    outputs(5774) <= not a;
    outputs(5775) <= a;
    outputs(5776) <= not b;
    outputs(5777) <= not (a and b);
    outputs(5778) <= a or b;
    outputs(5779) <= a;
    outputs(5780) <= a and b;
    outputs(5781) <= not a;
    outputs(5782) <= not (a xor b);
    outputs(5783) <= b;
    outputs(5784) <= not (a xor b);
    outputs(5785) <= a xor b;
    outputs(5786) <= not a;
    outputs(5787) <= not (a or b);
    outputs(5788) <= a or b;
    outputs(5789) <= a xor b;
    outputs(5790) <= not (a xor b);
    outputs(5791) <= not (a xor b);
    outputs(5792) <= a;
    outputs(5793) <= b and not a;
    outputs(5794) <= not a;
    outputs(5795) <= not b;
    outputs(5796) <= a or b;
    outputs(5797) <= b;
    outputs(5798) <= a or b;
    outputs(5799) <= a;
    outputs(5800) <= not b;
    outputs(5801) <= a and not b;
    outputs(5802) <= not a;
    outputs(5803) <= not b;
    outputs(5804) <= a;
    outputs(5805) <= a xor b;
    outputs(5806) <= not b;
    outputs(5807) <= not a;
    outputs(5808) <= not b or a;
    outputs(5809) <= a xor b;
    outputs(5810) <= a;
    outputs(5811) <= b;
    outputs(5812) <= a;
    outputs(5813) <= a;
    outputs(5814) <= not b;
    outputs(5815) <= a;
    outputs(5816) <= not a;
    outputs(5817) <= not b;
    outputs(5818) <= not (a xor b);
    outputs(5819) <= a;
    outputs(5820) <= not (a xor b);
    outputs(5821) <= b;
    outputs(5822) <= not b;
    outputs(5823) <= a;
    outputs(5824) <= b;
    outputs(5825) <= not (a xor b);
    outputs(5826) <= not b;
    outputs(5827) <= b;
    outputs(5828) <= a;
    outputs(5829) <= not (a or b);
    outputs(5830) <= not a;
    outputs(5831) <= not (a xor b);
    outputs(5832) <= not (a xor b);
    outputs(5833) <= not a or b;
    outputs(5834) <= not (a xor b);
    outputs(5835) <= b;
    outputs(5836) <= not (a xor b);
    outputs(5837) <= not a;
    outputs(5838) <= not (a xor b);
    outputs(5839) <= not (a xor b);
    outputs(5840) <= not a;
    outputs(5841) <= not a;
    outputs(5842) <= not b;
    outputs(5843) <= b and not a;
    outputs(5844) <= a and b;
    outputs(5845) <= not a;
    outputs(5846) <= a;
    outputs(5847) <= a and not b;
    outputs(5848) <= not (a xor b);
    outputs(5849) <= not a;
    outputs(5850) <= not a;
    outputs(5851) <= not (a or b);
    outputs(5852) <= b and not a;
    outputs(5853) <= b;
    outputs(5854) <= a;
    outputs(5855) <= b;
    outputs(5856) <= not b;
    outputs(5857) <= a;
    outputs(5858) <= b;
    outputs(5859) <= not b;
    outputs(5860) <= not (a xor b);
    outputs(5861) <= a;
    outputs(5862) <= not a;
    outputs(5863) <= a;
    outputs(5864) <= a and not b;
    outputs(5865) <= not a;
    outputs(5866) <= not (a xor b);
    outputs(5867) <= a or b;
    outputs(5868) <= a xor b;
    outputs(5869) <= b and not a;
    outputs(5870) <= not (a xor b);
    outputs(5871) <= b and not a;
    outputs(5872) <= not (a or b);
    outputs(5873) <= not (a xor b);
    outputs(5874) <= b;
    outputs(5875) <= not a or b;
    outputs(5876) <= a;
    outputs(5877) <= not a;
    outputs(5878) <= a and b;
    outputs(5879) <= not b;
    outputs(5880) <= a xor b;
    outputs(5881) <= not (a xor b);
    outputs(5882) <= not b;
    outputs(5883) <= not (a xor b);
    outputs(5884) <= a;
    outputs(5885) <= b;
    outputs(5886) <= not (a or b);
    outputs(5887) <= not (a or b);
    outputs(5888) <= not (a or b);
    outputs(5889) <= a and not b;
    outputs(5890) <= not (a xor b);
    outputs(5891) <= b and not a;
    outputs(5892) <= not a;
    outputs(5893) <= a;
    outputs(5894) <= not b;
    outputs(5895) <= b and not a;
    outputs(5896) <= not b;
    outputs(5897) <= not (a xor b);
    outputs(5898) <= b;
    outputs(5899) <= a xor b;
    outputs(5900) <= not a;
    outputs(5901) <= not (a or b);
    outputs(5902) <= not (a xor b);
    outputs(5903) <= b;
    outputs(5904) <= not (a xor b);
    outputs(5905) <= b and not a;
    outputs(5906) <= not a;
    outputs(5907) <= b;
    outputs(5908) <= b;
    outputs(5909) <= a and not b;
    outputs(5910) <= not b;
    outputs(5911) <= not b;
    outputs(5912) <= b;
    outputs(5913) <= a xor b;
    outputs(5914) <= a;
    outputs(5915) <= a xor b;
    outputs(5916) <= b;
    outputs(5917) <= not a;
    outputs(5918) <= b;
    outputs(5919) <= not a;
    outputs(5920) <= a and b;
    outputs(5921) <= not (a xor b);
    outputs(5922) <= not (a xor b);
    outputs(5923) <= a;
    outputs(5924) <= a;
    outputs(5925) <= b and not a;
    outputs(5926) <= a xor b;
    outputs(5927) <= not (a xor b);
    outputs(5928) <= a and b;
    outputs(5929) <= not b or a;
    outputs(5930) <= not (a xor b);
    outputs(5931) <= a xor b;
    outputs(5932) <= a and not b;
    outputs(5933) <= b;
    outputs(5934) <= a xor b;
    outputs(5935) <= not (a or b);
    outputs(5936) <= a xor b;
    outputs(5937) <= a xor b;
    outputs(5938) <= a xor b;
    outputs(5939) <= not (a xor b);
    outputs(5940) <= a xor b;
    outputs(5941) <= not b;
    outputs(5942) <= a and b;
    outputs(5943) <= a and not b;
    outputs(5944) <= a and b;
    outputs(5945) <= not a;
    outputs(5946) <= not b or a;
    outputs(5947) <= not a;
    outputs(5948) <= not a;
    outputs(5949) <= a and b;
    outputs(5950) <= not a;
    outputs(5951) <= not a;
    outputs(5952) <= b and not a;
    outputs(5953) <= a xor b;
    outputs(5954) <= b and not a;
    outputs(5955) <= not a;
    outputs(5956) <= not (a or b);
    outputs(5957) <= a xor b;
    outputs(5958) <= b and not a;
    outputs(5959) <= a xor b;
    outputs(5960) <= a and not b;
    outputs(5961) <= not a or b;
    outputs(5962) <= b;
    outputs(5963) <= a xor b;
    outputs(5964) <= not (a or b);
    outputs(5965) <= not a or b;
    outputs(5966) <= not (a and b);
    outputs(5967) <= not a;
    outputs(5968) <= not b or a;
    outputs(5969) <= a;
    outputs(5970) <= not a;
    outputs(5971) <= not (a xor b);
    outputs(5972) <= not (a or b);
    outputs(5973) <= not (a xor b);
    outputs(5974) <= not a;
    outputs(5975) <= a;
    outputs(5976) <= not (a xor b);
    outputs(5977) <= not b;
    outputs(5978) <= b;
    outputs(5979) <= b;
    outputs(5980) <= not a;
    outputs(5981) <= a and not b;
    outputs(5982) <= not b;
    outputs(5983) <= not a;
    outputs(5984) <= a and not b;
    outputs(5985) <= b;
    outputs(5986) <= not b;
    outputs(5987) <= not b or a;
    outputs(5988) <= b and not a;
    outputs(5989) <= a;
    outputs(5990) <= a or b;
    outputs(5991) <= a xor b;
    outputs(5992) <= not a;
    outputs(5993) <= a xor b;
    outputs(5994) <= a and not b;
    outputs(5995) <= a;
    outputs(5996) <= a and not b;
    outputs(5997) <= b;
    outputs(5998) <= a and not b;
    outputs(5999) <= a xor b;
    outputs(6000) <= b;
    outputs(6001) <= a and b;
    outputs(6002) <= not (a xor b);
    outputs(6003) <= not (a xor b);
    outputs(6004) <= a xor b;
    outputs(6005) <= a;
    outputs(6006) <= not (a and b);
    outputs(6007) <= a or b;
    outputs(6008) <= b;
    outputs(6009) <= not b;
    outputs(6010) <= not a;
    outputs(6011) <= b;
    outputs(6012) <= not a;
    outputs(6013) <= not (a xor b);
    outputs(6014) <= a xor b;
    outputs(6015) <= a xor b;
    outputs(6016) <= not a or b;
    outputs(6017) <= a xor b;
    outputs(6018) <= not b;
    outputs(6019) <= not (a xor b);
    outputs(6020) <= b;
    outputs(6021) <= not a;
    outputs(6022) <= not b;
    outputs(6023) <= b and not a;
    outputs(6024) <= a;
    outputs(6025) <= b;
    outputs(6026) <= a;
    outputs(6027) <= b and not a;
    outputs(6028) <= a and not b;
    outputs(6029) <= a xor b;
    outputs(6030) <= a xor b;
    outputs(6031) <= a and b;
    outputs(6032) <= a and b;
    outputs(6033) <= a and not b;
    outputs(6034) <= a xor b;
    outputs(6035) <= not a;
    outputs(6036) <= a and not b;
    outputs(6037) <= a and not b;
    outputs(6038) <= b;
    outputs(6039) <= not (a xor b);
    outputs(6040) <= a xor b;
    outputs(6041) <= a or b;
    outputs(6042) <= not (a xor b);
    outputs(6043) <= b and not a;
    outputs(6044) <= not b;
    outputs(6045) <= b;
    outputs(6046) <= b;
    outputs(6047) <= not (a xor b);
    outputs(6048) <= not (a xor b);
    outputs(6049) <= b;
    outputs(6050) <= b and not a;
    outputs(6051) <= not (a or b);
    outputs(6052) <= a;
    outputs(6053) <= not a;
    outputs(6054) <= not (a or b);
    outputs(6055) <= a and not b;
    outputs(6056) <= not (a xor b);
    outputs(6057) <= b;
    outputs(6058) <= not b;
    outputs(6059) <= not a;
    outputs(6060) <= not (a xor b);
    outputs(6061) <= not (a xor b);
    outputs(6062) <= b;
    outputs(6063) <= b and not a;
    outputs(6064) <= b;
    outputs(6065) <= not b;
    outputs(6066) <= b;
    outputs(6067) <= not a;
    outputs(6068) <= not a or b;
    outputs(6069) <= a and not b;
    outputs(6070) <= not (a or b);
    outputs(6071) <= a and b;
    outputs(6072) <= a xor b;
    outputs(6073) <= a xor b;
    outputs(6074) <= not (a xor b);
    outputs(6075) <= not (a or b);
    outputs(6076) <= b;
    outputs(6077) <= not b;
    outputs(6078) <= a xor b;
    outputs(6079) <= not (a xor b);
    outputs(6080) <= a and not b;
    outputs(6081) <= not (a xor b);
    outputs(6082) <= not b;
    outputs(6083) <= a and b;
    outputs(6084) <= a;
    outputs(6085) <= b;
    outputs(6086) <= a and not b;
    outputs(6087) <= a;
    outputs(6088) <= not b;
    outputs(6089) <= a or b;
    outputs(6090) <= a or b;
    outputs(6091) <= a;
    outputs(6092) <= not b;
    outputs(6093) <= a;
    outputs(6094) <= a xor b;
    outputs(6095) <= not a;
    outputs(6096) <= a and b;
    outputs(6097) <= not a or b;
    outputs(6098) <= not a;
    outputs(6099) <= not (a xor b);
    outputs(6100) <= a and b;
    outputs(6101) <= b;
    outputs(6102) <= a xor b;
    outputs(6103) <= not a;
    outputs(6104) <= not a;
    outputs(6105) <= not (a or b);
    outputs(6106) <= a and not b;
    outputs(6107) <= a;
    outputs(6108) <= not (a xor b);
    outputs(6109) <= not (a xor b);
    outputs(6110) <= b and not a;
    outputs(6111) <= not b;
    outputs(6112) <= a;
    outputs(6113) <= b;
    outputs(6114) <= b;
    outputs(6115) <= not (a or b);
    outputs(6116) <= not (a or b);
    outputs(6117) <= a;
    outputs(6118) <= not a;
    outputs(6119) <= a and b;
    outputs(6120) <= not b;
    outputs(6121) <= a xor b;
    outputs(6122) <= not a;
    outputs(6123) <= a and not b;
    outputs(6124) <= not (a xor b);
    outputs(6125) <= b;
    outputs(6126) <= not b;
    outputs(6127) <= a xor b;
    outputs(6128) <= a and not b;
    outputs(6129) <= not b or a;
    outputs(6130) <= not (a xor b);
    outputs(6131) <= a and not b;
    outputs(6132) <= b;
    outputs(6133) <= a;
    outputs(6134) <= b;
    outputs(6135) <= not b;
    outputs(6136) <= a;
    outputs(6137) <= a xor b;
    outputs(6138) <= not (a xor b);
    outputs(6139) <= not (a xor b);
    outputs(6140) <= not (a xor b);
    outputs(6141) <= a xor b;
    outputs(6142) <= b and not a;
    outputs(6143) <= b and not a;
    outputs(6144) <= a or b;
    outputs(6145) <= a;
    outputs(6146) <= b;
    outputs(6147) <= a xor b;
    outputs(6148) <= not b;
    outputs(6149) <= not (a or b);
    outputs(6150) <= a xor b;
    outputs(6151) <= b;
    outputs(6152) <= not (a xor b);
    outputs(6153) <= not (a xor b);
    outputs(6154) <= not b or a;
    outputs(6155) <= a xor b;
    outputs(6156) <= not b;
    outputs(6157) <= not a;
    outputs(6158) <= not (a or b);
    outputs(6159) <= b and not a;
    outputs(6160) <= not (a and b);
    outputs(6161) <= a or b;
    outputs(6162) <= a xor b;
    outputs(6163) <= not (a xor b);
    outputs(6164) <= not a;
    outputs(6165) <= a;
    outputs(6166) <= not a;
    outputs(6167) <= not a;
    outputs(6168) <= not (a xor b);
    outputs(6169) <= not (a xor b);
    outputs(6170) <= a;
    outputs(6171) <= a and not b;
    outputs(6172) <= not b;
    outputs(6173) <= a xor b;
    outputs(6174) <= not b;
    outputs(6175) <= not a;
    outputs(6176) <= b;
    outputs(6177) <= a and not b;
    outputs(6178) <= not (a xor b);
    outputs(6179) <= a and not b;
    outputs(6180) <= a xor b;
    outputs(6181) <= not a or b;
    outputs(6182) <= a and b;
    outputs(6183) <= not b;
    outputs(6184) <= a and not b;
    outputs(6185) <= not a;
    outputs(6186) <= not a;
    outputs(6187) <= not (a and b);
    outputs(6188) <= not (a xor b);
    outputs(6189) <= not (a xor b);
    outputs(6190) <= a and not b;
    outputs(6191) <= a xor b;
    outputs(6192) <= not b;
    outputs(6193) <= not b;
    outputs(6194) <= not a;
    outputs(6195) <= not (a xor b);
    outputs(6196) <= a;
    outputs(6197) <= not a;
    outputs(6198) <= b;
    outputs(6199) <= a;
    outputs(6200) <= not a;
    outputs(6201) <= a;
    outputs(6202) <= not (a and b);
    outputs(6203) <= not a;
    outputs(6204) <= a;
    outputs(6205) <= not a or b;
    outputs(6206) <= b;
    outputs(6207) <= not (a xor b);
    outputs(6208) <= not (a xor b);
    outputs(6209) <= a;
    outputs(6210) <= not (a or b);
    outputs(6211) <= not b or a;
    outputs(6212) <= a xor b;
    outputs(6213) <= not (a and b);
    outputs(6214) <= not b;
    outputs(6215) <= not b or a;
    outputs(6216) <= not (a and b);
    outputs(6217) <= not b or a;
    outputs(6218) <= b;
    outputs(6219) <= b;
    outputs(6220) <= b and not a;
    outputs(6221) <= not (a xor b);
    outputs(6222) <= not a or b;
    outputs(6223) <= not a;
    outputs(6224) <= b;
    outputs(6225) <= not (a xor b);
    outputs(6226) <= not b;
    outputs(6227) <= not b;
    outputs(6228) <= b;
    outputs(6229) <= not a or b;
    outputs(6230) <= a xor b;
    outputs(6231) <= a xor b;
    outputs(6232) <= b;
    outputs(6233) <= a xor b;
    outputs(6234) <= not a;
    outputs(6235) <= b;
    outputs(6236) <= not (a xor b);
    outputs(6237) <= not b;
    outputs(6238) <= not a;
    outputs(6239) <= a and not b;
    outputs(6240) <= a;
    outputs(6241) <= a xor b;
    outputs(6242) <= not b;
    outputs(6243) <= b;
    outputs(6244) <= not b;
    outputs(6245) <= a and not b;
    outputs(6246) <= not (a or b);
    outputs(6247) <= a and not b;
    outputs(6248) <= a xor b;
    outputs(6249) <= b;
    outputs(6250) <= not (a xor b);
    outputs(6251) <= not b;
    outputs(6252) <= not (a xor b);
    outputs(6253) <= not b;
    outputs(6254) <= a;
    outputs(6255) <= a or b;
    outputs(6256) <= b;
    outputs(6257) <= not b;
    outputs(6258) <= a xor b;
    outputs(6259) <= b;
    outputs(6260) <= a xor b;
    outputs(6261) <= a;
    outputs(6262) <= a and not b;
    outputs(6263) <= b;
    outputs(6264) <= not a;
    outputs(6265) <= b;
    outputs(6266) <= b;
    outputs(6267) <= a xor b;
    outputs(6268) <= not b;
    outputs(6269) <= a xor b;
    outputs(6270) <= not (a xor b);
    outputs(6271) <= a and not b;
    outputs(6272) <= not (a xor b);
    outputs(6273) <= not a;
    outputs(6274) <= a;
    outputs(6275) <= b;
    outputs(6276) <= not a;
    outputs(6277) <= not a;
    outputs(6278) <= a or b;
    outputs(6279) <= b and not a;
    outputs(6280) <= a or b;
    outputs(6281) <= a xor b;
    outputs(6282) <= not (a xor b);
    outputs(6283) <= not (a xor b);
    outputs(6284) <= a xor b;
    outputs(6285) <= a xor b;
    outputs(6286) <= a;
    outputs(6287) <= not a or b;
    outputs(6288) <= not (a xor b);
    outputs(6289) <= not b;
    outputs(6290) <= not b;
    outputs(6291) <= a xor b;
    outputs(6292) <= not b;
    outputs(6293) <= b;
    outputs(6294) <= not a;
    outputs(6295) <= b and not a;
    outputs(6296) <= not a;
    outputs(6297) <= not b;
    outputs(6298) <= a xor b;
    outputs(6299) <= not (a xor b);
    outputs(6300) <= a and not b;
    outputs(6301) <= not b;
    outputs(6302) <= not a;
    outputs(6303) <= not b;
    outputs(6304) <= not (a xor b);
    outputs(6305) <= a;
    outputs(6306) <= a xor b;
    outputs(6307) <= not b;
    outputs(6308) <= a;
    outputs(6309) <= not b or a;
    outputs(6310) <= a;
    outputs(6311) <= a xor b;
    outputs(6312) <= not b or a;
    outputs(6313) <= not a;
    outputs(6314) <= not b or a;
    outputs(6315) <= a and b;
    outputs(6316) <= not b;
    outputs(6317) <= a xor b;
    outputs(6318) <= a;
    outputs(6319) <= b;
    outputs(6320) <= not (a and b);
    outputs(6321) <= not a or b;
    outputs(6322) <= not (a xor b);
    outputs(6323) <= not a;
    outputs(6324) <= a xor b;
    outputs(6325) <= a;
    outputs(6326) <= b;
    outputs(6327) <= not (a xor b);
    outputs(6328) <= a or b;
    outputs(6329) <= not a;
    outputs(6330) <= not a;
    outputs(6331) <= a;
    outputs(6332) <= not b;
    outputs(6333) <= b;
    outputs(6334) <= not a;
    outputs(6335) <= b and not a;
    outputs(6336) <= b;
    outputs(6337) <= b;
    outputs(6338) <= a and not b;
    outputs(6339) <= not b;
    outputs(6340) <= a and not b;
    outputs(6341) <= not b;
    outputs(6342) <= a;
    outputs(6343) <= not (a and b);
    outputs(6344) <= not (a xor b);
    outputs(6345) <= not (a or b);
    outputs(6346) <= not b;
    outputs(6347) <= b and not a;
    outputs(6348) <= a and not b;
    outputs(6349) <= not b;
    outputs(6350) <= a;
    outputs(6351) <= not b;
    outputs(6352) <= not a or b;
    outputs(6353) <= not b;
    outputs(6354) <= a xor b;
    outputs(6355) <= not (a and b);
    outputs(6356) <= b;
    outputs(6357) <= not (a xor b);
    outputs(6358) <= a;
    outputs(6359) <= a xor b;
    outputs(6360) <= not a;
    outputs(6361) <= b and not a;
    outputs(6362) <= a xor b;
    outputs(6363) <= not (a xor b);
    outputs(6364) <= not b;
    outputs(6365) <= a xor b;
    outputs(6366) <= b;
    outputs(6367) <= b;
    outputs(6368) <= b;
    outputs(6369) <= not (a xor b);
    outputs(6370) <= not b;
    outputs(6371) <= not (a xor b);
    outputs(6372) <= a;
    outputs(6373) <= a or b;
    outputs(6374) <= b and not a;
    outputs(6375) <= a xor b;
    outputs(6376) <= not b or a;
    outputs(6377) <= a xor b;
    outputs(6378) <= b;
    outputs(6379) <= not a;
    outputs(6380) <= a or b;
    outputs(6381) <= not a;
    outputs(6382) <= not a;
    outputs(6383) <= b and not a;
    outputs(6384) <= not b;
    outputs(6385) <= a;
    outputs(6386) <= not b or a;
    outputs(6387) <= not (a xor b);
    outputs(6388) <= not a or b;
    outputs(6389) <= not b;
    outputs(6390) <= b;
    outputs(6391) <= b and not a;
    outputs(6392) <= not b;
    outputs(6393) <= a xor b;
    outputs(6394) <= not a;
    outputs(6395) <= not (a xor b);
    outputs(6396) <= not (a xor b);
    outputs(6397) <= a and b;
    outputs(6398) <= a and b;
    outputs(6399) <= not a or b;
    outputs(6400) <= not b;
    outputs(6401) <= not (a xor b);
    outputs(6402) <= not (a xor b);
    outputs(6403) <= b;
    outputs(6404) <= a xor b;
    outputs(6405) <= a or b;
    outputs(6406) <= b;
    outputs(6407) <= a xor b;
    outputs(6408) <= not b;
    outputs(6409) <= a and not b;
    outputs(6410) <= a or b;
    outputs(6411) <= not b;
    outputs(6412) <= a xor b;
    outputs(6413) <= b;
    outputs(6414) <= not b or a;
    outputs(6415) <= b;
    outputs(6416) <= not (a xor b);
    outputs(6417) <= not (a xor b);
    outputs(6418) <= not a;
    outputs(6419) <= a or b;
    outputs(6420) <= a;
    outputs(6421) <= b;
    outputs(6422) <= a;
    outputs(6423) <= not b;
    outputs(6424) <= b;
    outputs(6425) <= not (a xor b);
    outputs(6426) <= a;
    outputs(6427) <= not (a xor b);
    outputs(6428) <= not b or a;
    outputs(6429) <= not (a or b);
    outputs(6430) <= not (a xor b);
    outputs(6431) <= not (a xor b);
    outputs(6432) <= not a;
    outputs(6433) <= not b;
    outputs(6434) <= a xor b;
    outputs(6435) <= not b;
    outputs(6436) <= not (a xor b);
    outputs(6437) <= not a;
    outputs(6438) <= b;
    outputs(6439) <= not a;
    outputs(6440) <= not (a xor b);
    outputs(6441) <= not a or b;
    outputs(6442) <= a xor b;
    outputs(6443) <= not (a xor b);
    outputs(6444) <= not b;
    outputs(6445) <= not a;
    outputs(6446) <= a and b;
    outputs(6447) <= not a;
    outputs(6448) <= not a;
    outputs(6449) <= a and b;
    outputs(6450) <= not a;
    outputs(6451) <= b;
    outputs(6452) <= not (a xor b);
    outputs(6453) <= not (a xor b);
    outputs(6454) <= not (a xor b);
    outputs(6455) <= not b;
    outputs(6456) <= a xor b;
    outputs(6457) <= a xor b;
    outputs(6458) <= not a;
    outputs(6459) <= a and b;
    outputs(6460) <= not (a xor b);
    outputs(6461) <= a;
    outputs(6462) <= not b;
    outputs(6463) <= a xor b;
    outputs(6464) <= a xor b;
    outputs(6465) <= not b;
    outputs(6466) <= not a;
    outputs(6467) <= not a;
    outputs(6468) <= a xor b;
    outputs(6469) <= not (a and b);
    outputs(6470) <= a xor b;
    outputs(6471) <= not (a or b);
    outputs(6472) <= not a or b;
    outputs(6473) <= not b;
    outputs(6474) <= a xor b;
    outputs(6475) <= not a or b;
    outputs(6476) <= a xor b;
    outputs(6477) <= a;
    outputs(6478) <= b;
    outputs(6479) <= not b or a;
    outputs(6480) <= a xor b;
    outputs(6481) <= not (a xor b);
    outputs(6482) <= a or b;
    outputs(6483) <= a;
    outputs(6484) <= b and not a;
    outputs(6485) <= not (a xor b);
    outputs(6486) <= a xor b;
    outputs(6487) <= a;
    outputs(6488) <= not (a xor b);
    outputs(6489) <= not a;
    outputs(6490) <= a xor b;
    outputs(6491) <= a;
    outputs(6492) <= a xor b;
    outputs(6493) <= a xor b;
    outputs(6494) <= not (a and b);
    outputs(6495) <= not (a xor b);
    outputs(6496) <= not (a and b);
    outputs(6497) <= a xor b;
    outputs(6498) <= not (a xor b);
    outputs(6499) <= a xor b;
    outputs(6500) <= not b;
    outputs(6501) <= not b;
    outputs(6502) <= not a;
    outputs(6503) <= not a;
    outputs(6504) <= a xor b;
    outputs(6505) <= not (a xor b);
    outputs(6506) <= a xor b;
    outputs(6507) <= not a or b;
    outputs(6508) <= not (a xor b);
    outputs(6509) <= not (a xor b);
    outputs(6510) <= b;
    outputs(6511) <= not b;
    outputs(6512) <= not (a xor b);
    outputs(6513) <= not (a xor b);
    outputs(6514) <= a;
    outputs(6515) <= a xor b;
    outputs(6516) <= not (a xor b);
    outputs(6517) <= a xor b;
    outputs(6518) <= not a;
    outputs(6519) <= not (a and b);
    outputs(6520) <= not (a and b);
    outputs(6521) <= not (a or b);
    outputs(6522) <= a;
    outputs(6523) <= a and b;
    outputs(6524) <= not (a xor b);
    outputs(6525) <= not (a xor b);
    outputs(6526) <= not (a xor b);
    outputs(6527) <= not (a xor b);
    outputs(6528) <= not (a or b);
    outputs(6529) <= not a;
    outputs(6530) <= not (a or b);
    outputs(6531) <= b and not a;
    outputs(6532) <= a xor b;
    outputs(6533) <= not b;
    outputs(6534) <= a;
    outputs(6535) <= not (a and b);
    outputs(6536) <= not (a xor b);
    outputs(6537) <= not a;
    outputs(6538) <= not (a xor b);
    outputs(6539) <= a and b;
    outputs(6540) <= a xor b;
    outputs(6541) <= a xor b;
    outputs(6542) <= a and not b;
    outputs(6543) <= a xor b;
    outputs(6544) <= b;
    outputs(6545) <= a xor b;
    outputs(6546) <= not a;
    outputs(6547) <= a xor b;
    outputs(6548) <= a;
    outputs(6549) <= b;
    outputs(6550) <= a xor b;
    outputs(6551) <= not (a or b);
    outputs(6552) <= b;
    outputs(6553) <= '1';
    outputs(6554) <= a xor b;
    outputs(6555) <= a and b;
    outputs(6556) <= a;
    outputs(6557) <= not b;
    outputs(6558) <= not b;
    outputs(6559) <= a and b;
    outputs(6560) <= not (a xor b);
    outputs(6561) <= a;
    outputs(6562) <= not (a xor b);
    outputs(6563) <= not a;
    outputs(6564) <= not (a xor b);
    outputs(6565) <= a xor b;
    outputs(6566) <= not b;
    outputs(6567) <= a xor b;
    outputs(6568) <= not b;
    outputs(6569) <= not (a xor b);
    outputs(6570) <= not b;
    outputs(6571) <= not b or a;
    outputs(6572) <= not b;
    outputs(6573) <= a xor b;
    outputs(6574) <= not b or a;
    outputs(6575) <= not a;
    outputs(6576) <= not b or a;
    outputs(6577) <= not (a xor b);
    outputs(6578) <= not (a and b);
    outputs(6579) <= a xor b;
    outputs(6580) <= not b or a;
    outputs(6581) <= not (a or b);
    outputs(6582) <= not b;
    outputs(6583) <= not (a xor b);
    outputs(6584) <= not (a xor b);
    outputs(6585) <= not (a and b);
    outputs(6586) <= a xor b;
    outputs(6587) <= not a;
    outputs(6588) <= not (a xor b);
    outputs(6589) <= a xor b;
    outputs(6590) <= a xor b;
    outputs(6591) <= not (a xor b);
    outputs(6592) <= not (a xor b);
    outputs(6593) <= not b;
    outputs(6594) <= not a;
    outputs(6595) <= a;
    outputs(6596) <= b and not a;
    outputs(6597) <= not b;
    outputs(6598) <= a and b;
    outputs(6599) <= b and not a;
    outputs(6600) <= a;
    outputs(6601) <= a and not b;
    outputs(6602) <= not b or a;
    outputs(6603) <= a and not b;
    outputs(6604) <= not (a and b);
    outputs(6605) <= a xor b;
    outputs(6606) <= a;
    outputs(6607) <= not (a and b);
    outputs(6608) <= b;
    outputs(6609) <= a;
    outputs(6610) <= not a or b;
    outputs(6611) <= a xor b;
    outputs(6612) <= a;
    outputs(6613) <= a xor b;
    outputs(6614) <= not (a or b);
    outputs(6615) <= not (a xor b);
    outputs(6616) <= not a;
    outputs(6617) <= a xor b;
    outputs(6618) <= not (a xor b);
    outputs(6619) <= a xor b;
    outputs(6620) <= a;
    outputs(6621) <= a and b;
    outputs(6622) <= b;
    outputs(6623) <= not a;
    outputs(6624) <= a and b;
    outputs(6625) <= a;
    outputs(6626) <= not b;
    outputs(6627) <= not b;
    outputs(6628) <= not (a or b);
    outputs(6629) <= not a;
    outputs(6630) <= b and not a;
    outputs(6631) <= not b or a;
    outputs(6632) <= not (a xor b);
    outputs(6633) <= not b;
    outputs(6634) <= a xor b;
    outputs(6635) <= not (a xor b);
    outputs(6636) <= b;
    outputs(6637) <= a or b;
    outputs(6638) <= not a;
    outputs(6639) <= a;
    outputs(6640) <= not (a xor b);
    outputs(6641) <= a;
    outputs(6642) <= a;
    outputs(6643) <= not b;
    outputs(6644) <= a;
    outputs(6645) <= not a;
    outputs(6646) <= a xor b;
    outputs(6647) <= a and not b;
    outputs(6648) <= not (a or b);
    outputs(6649) <= not b;
    outputs(6650) <= not a;
    outputs(6651) <= b and not a;
    outputs(6652) <= a or b;
    outputs(6653) <= a;
    outputs(6654) <= a xor b;
    outputs(6655) <= not b;
    outputs(6656) <= a and b;
    outputs(6657) <= a and b;
    outputs(6658) <= not (a xor b);
    outputs(6659) <= a;
    outputs(6660) <= b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= a and not b;
    outputs(6663) <= not b;
    outputs(6664) <= b;
    outputs(6665) <= a and not b;
    outputs(6666) <= not b or a;
    outputs(6667) <= not a or b;
    outputs(6668) <= not (a xor b);
    outputs(6669) <= not b or a;
    outputs(6670) <= a xor b;
    outputs(6671) <= not b;
    outputs(6672) <= not (a xor b);
    outputs(6673) <= b;
    outputs(6674) <= not (a xor b);
    outputs(6675) <= b;
    outputs(6676) <= a xor b;
    outputs(6677) <= not (a xor b);
    outputs(6678) <= b;
    outputs(6679) <= not b;
    outputs(6680) <= not b or a;
    outputs(6681) <= not (a or b);
    outputs(6682) <= not (a xor b);
    outputs(6683) <= b;
    outputs(6684) <= b;
    outputs(6685) <= a xor b;
    outputs(6686) <= a xor b;
    outputs(6687) <= a or b;
    outputs(6688) <= a xor b;
    outputs(6689) <= a xor b;
    outputs(6690) <= a;
    outputs(6691) <= b;
    outputs(6692) <= b;
    outputs(6693) <= a;
    outputs(6694) <= a xor b;
    outputs(6695) <= a or b;
    outputs(6696) <= b;
    outputs(6697) <= a;
    outputs(6698) <= not a;
    outputs(6699) <= not (a xor b);
    outputs(6700) <= not b;
    outputs(6701) <= a and not b;
    outputs(6702) <= not (a xor b);
    outputs(6703) <= not (a xor b);
    outputs(6704) <= not b;
    outputs(6705) <= b and not a;
    outputs(6706) <= not a;
    outputs(6707) <= not b;
    outputs(6708) <= not (a xor b);
    outputs(6709) <= a;
    outputs(6710) <= not (a and b);
    outputs(6711) <= not a;
    outputs(6712) <= not (a xor b);
    outputs(6713) <= a xor b;
    outputs(6714) <= a xor b;
    outputs(6715) <= not a;
    outputs(6716) <= not a;
    outputs(6717) <= not b;
    outputs(6718) <= a xor b;
    outputs(6719) <= not (a xor b);
    outputs(6720) <= a;
    outputs(6721) <= a xor b;
    outputs(6722) <= b and not a;
    outputs(6723) <= a and not b;
    outputs(6724) <= a and not b;
    outputs(6725) <= not a;
    outputs(6726) <= b and not a;
    outputs(6727) <= not (a xor b);
    outputs(6728) <= a xor b;
    outputs(6729) <= a and b;
    outputs(6730) <= a;
    outputs(6731) <= not b;
    outputs(6732) <= not a;
    outputs(6733) <= not (a xor b);
    outputs(6734) <= not b;
    outputs(6735) <= not b;
    outputs(6736) <= not a;
    outputs(6737) <= not (a and b);
    outputs(6738) <= a xor b;
    outputs(6739) <= not (a xor b);
    outputs(6740) <= a xor b;
    outputs(6741) <= b;
    outputs(6742) <= not (a xor b);
    outputs(6743) <= not (a xor b);
    outputs(6744) <= a xor b;
    outputs(6745) <= b and not a;
    outputs(6746) <= a;
    outputs(6747) <= a xor b;
    outputs(6748) <= a;
    outputs(6749) <= not b;
    outputs(6750) <= not b;
    outputs(6751) <= a or b;
    outputs(6752) <= not b;
    outputs(6753) <= b;
    outputs(6754) <= not b;
    outputs(6755) <= a and b;
    outputs(6756) <= a xor b;
    outputs(6757) <= a xor b;
    outputs(6758) <= not (a xor b);
    outputs(6759) <= not a or b;
    outputs(6760) <= not b;
    outputs(6761) <= b;
    outputs(6762) <= a;
    outputs(6763) <= not a;
    outputs(6764) <= not (a and b);
    outputs(6765) <= not b;
    outputs(6766) <= not a or b;
    outputs(6767) <= not a;
    outputs(6768) <= b;
    outputs(6769) <= b;
    outputs(6770) <= a xor b;
    outputs(6771) <= b;
    outputs(6772) <= a and not b;
    outputs(6773) <= not b;
    outputs(6774) <= b;
    outputs(6775) <= not a;
    outputs(6776) <= b;
    outputs(6777) <= a xor b;
    outputs(6778) <= not a or b;
    outputs(6779) <= a xor b;
    outputs(6780) <= a;
    outputs(6781) <= not a or b;
    outputs(6782) <= not a;
    outputs(6783) <= not (a xor b);
    outputs(6784) <= a xor b;
    outputs(6785) <= a and not b;
    outputs(6786) <= not b;
    outputs(6787) <= a;
    outputs(6788) <= a;
    outputs(6789) <= a;
    outputs(6790) <= not (a xor b);
    outputs(6791) <= not b or a;
    outputs(6792) <= not b;
    outputs(6793) <= a xor b;
    outputs(6794) <= not b;
    outputs(6795) <= not a or b;
    outputs(6796) <= not b or a;
    outputs(6797) <= a xor b;
    outputs(6798) <= a xor b;
    outputs(6799) <= not a;
    outputs(6800) <= a or b;
    outputs(6801) <= not (a xor b);
    outputs(6802) <= not (a xor b);
    outputs(6803) <= not a;
    outputs(6804) <= not b;
    outputs(6805) <= not b;
    outputs(6806) <= not b;
    outputs(6807) <= b and not a;
    outputs(6808) <= a and not b;
    outputs(6809) <= b and not a;
    outputs(6810) <= a xor b;
    outputs(6811) <= a;
    outputs(6812) <= a;
    outputs(6813) <= b;
    outputs(6814) <= not b or a;
    outputs(6815) <= a;
    outputs(6816) <= a xor b;
    outputs(6817) <= not b or a;
    outputs(6818) <= not (a and b);
    outputs(6819) <= b and not a;
    outputs(6820) <= a;
    outputs(6821) <= a;
    outputs(6822) <= b;
    outputs(6823) <= not (a and b);
    outputs(6824) <= not (a xor b);
    outputs(6825) <= not b;
    outputs(6826) <= not (a or b);
    outputs(6827) <= b;
    outputs(6828) <= not (a or b);
    outputs(6829) <= b;
    outputs(6830) <= not a;
    outputs(6831) <= not (a xor b);
    outputs(6832) <= not a;
    outputs(6833) <= not (a xor b);
    outputs(6834) <= b;
    outputs(6835) <= not (a xor b);
    outputs(6836) <= a and not b;
    outputs(6837) <= b;
    outputs(6838) <= not a;
    outputs(6839) <= b;
    outputs(6840) <= b and not a;
    outputs(6841) <= not a;
    outputs(6842) <= not (a xor b);
    outputs(6843) <= b;
    outputs(6844) <= a xor b;
    outputs(6845) <= not a;
    outputs(6846) <= a and not b;
    outputs(6847) <= a and b;
    outputs(6848) <= a and not b;
    outputs(6849) <= not (a xor b);
    outputs(6850) <= not b;
    outputs(6851) <= a xor b;
    outputs(6852) <= a xor b;
    outputs(6853) <= not b;
    outputs(6854) <= b;
    outputs(6855) <= not (a xor b);
    outputs(6856) <= not a;
    outputs(6857) <= not b;
    outputs(6858) <= a xor b;
    outputs(6859) <= not a or b;
    outputs(6860) <= a and b;
    outputs(6861) <= not a or b;
    outputs(6862) <= not (a xor b);
    outputs(6863) <= a;
    outputs(6864) <= a xor b;
    outputs(6865) <= not b;
    outputs(6866) <= not b;
    outputs(6867) <= b;
    outputs(6868) <= not (a xor b);
    outputs(6869) <= a;
    outputs(6870) <= not a;
    outputs(6871) <= not b or a;
    outputs(6872) <= a;
    outputs(6873) <= a xor b;
    outputs(6874) <= a xor b;
    outputs(6875) <= not (a xor b);
    outputs(6876) <= not (a and b);
    outputs(6877) <= not (a xor b);
    outputs(6878) <= a xor b;
    outputs(6879) <= not (a xor b);
    outputs(6880) <= b;
    outputs(6881) <= a or b;
    outputs(6882) <= not (a and b);
    outputs(6883) <= not b;
    outputs(6884) <= not (a xor b);
    outputs(6885) <= a or b;
    outputs(6886) <= a;
    outputs(6887) <= not a;
    outputs(6888) <= b;
    outputs(6889) <= b;
    outputs(6890) <= not b or a;
    outputs(6891) <= not (a xor b);
    outputs(6892) <= a xor b;
    outputs(6893) <= a xor b;
    outputs(6894) <= not a or b;
    outputs(6895) <= b;
    outputs(6896) <= a and b;
    outputs(6897) <= not (a or b);
    outputs(6898) <= not a;
    outputs(6899) <= not b;
    outputs(6900) <= not (a xor b);
    outputs(6901) <= b and not a;
    outputs(6902) <= not (a xor b);
    outputs(6903) <= a and not b;
    outputs(6904) <= not (a xor b);
    outputs(6905) <= b;
    outputs(6906) <= b;
    outputs(6907) <= a;
    outputs(6908) <= not (a and b);
    outputs(6909) <= not a or b;
    outputs(6910) <= not b;
    outputs(6911) <= not a;
    outputs(6912) <= a xor b;
    outputs(6913) <= not a;
    outputs(6914) <= b;
    outputs(6915) <= b;
    outputs(6916) <= b;
    outputs(6917) <= a xor b;
    outputs(6918) <= not a;
    outputs(6919) <= b and not a;
    outputs(6920) <= not a;
    outputs(6921) <= not (a or b);
    outputs(6922) <= a xor b;
    outputs(6923) <= b;
    outputs(6924) <= not (a xor b);
    outputs(6925) <= a xor b;
    outputs(6926) <= a;
    outputs(6927) <= not (a xor b);
    outputs(6928) <= b;
    outputs(6929) <= not (a or b);
    outputs(6930) <= a xor b;
    outputs(6931) <= not a;
    outputs(6932) <= a xor b;
    outputs(6933) <= not (a xor b);
    outputs(6934) <= not a;
    outputs(6935) <= a xor b;
    outputs(6936) <= a xor b;
    outputs(6937) <= not (a xor b);
    outputs(6938) <= a and not b;
    outputs(6939) <= not b;
    outputs(6940) <= a xor b;
    outputs(6941) <= a xor b;
    outputs(6942) <= not b;
    outputs(6943) <= a xor b;
    outputs(6944) <= not b;
    outputs(6945) <= a;
    outputs(6946) <= not (a and b);
    outputs(6947) <= not a;
    outputs(6948) <= b;
    outputs(6949) <= not b;
    outputs(6950) <= b;
    outputs(6951) <= a xor b;
    outputs(6952) <= not (a or b);
    outputs(6953) <= not (a xor b);
    outputs(6954) <= not b;
    outputs(6955) <= a;
    outputs(6956) <= not (a xor b);
    outputs(6957) <= a xor b;
    outputs(6958) <= a xor b;
    outputs(6959) <= a xor b;
    outputs(6960) <= a xor b;
    outputs(6961) <= not (a xor b);
    outputs(6962) <= not a;
    outputs(6963) <= not (a or b);
    outputs(6964) <= a xor b;
    outputs(6965) <= a xor b;
    outputs(6966) <= not a or b;
    outputs(6967) <= a xor b;
    outputs(6968) <= not (a xor b);
    outputs(6969) <= not (a or b);
    outputs(6970) <= b;
    outputs(6971) <= not a;
    outputs(6972) <= a;
    outputs(6973) <= not a or b;
    outputs(6974) <= not (a xor b);
    outputs(6975) <= a xor b;
    outputs(6976) <= a and b;
    outputs(6977) <= a xor b;
    outputs(6978) <= not b;
    outputs(6979) <= a and not b;
    outputs(6980) <= a xor b;
    outputs(6981) <= not a;
    outputs(6982) <= a;
    outputs(6983) <= a;
    outputs(6984) <= not (a xor b);
    outputs(6985) <= b;
    outputs(6986) <= a;
    outputs(6987) <= not b or a;
    outputs(6988) <= b;
    outputs(6989) <= b and not a;
    outputs(6990) <= not (a xor b);
    outputs(6991) <= not a;
    outputs(6992) <= not b;
    outputs(6993) <= not (a or b);
    outputs(6994) <= b;
    outputs(6995) <= a xor b;
    outputs(6996) <= not (a xor b);
    outputs(6997) <= a;
    outputs(6998) <= a and b;
    outputs(6999) <= a xor b;
    outputs(7000) <= not a or b;
    outputs(7001) <= not (a xor b);
    outputs(7002) <= not a;
    outputs(7003) <= not (a xor b);
    outputs(7004) <= not (a xor b);
    outputs(7005) <= a;
    outputs(7006) <= not (a or b);
    outputs(7007) <= a;
    outputs(7008) <= not (a or b);
    outputs(7009) <= not a;
    outputs(7010) <= not b;
    outputs(7011) <= not a;
    outputs(7012) <= not (a xor b);
    outputs(7013) <= not a;
    outputs(7014) <= b and not a;
    outputs(7015) <= a;
    outputs(7016) <= b;
    outputs(7017) <= a xor b;
    outputs(7018) <= not (a xor b);
    outputs(7019) <= not (a xor b);
    outputs(7020) <= b;
    outputs(7021) <= b;
    outputs(7022) <= not (a xor b);
    outputs(7023) <= b;
    outputs(7024) <= a;
    outputs(7025) <= not a;
    outputs(7026) <= not b;
    outputs(7027) <= not (a xor b);
    outputs(7028) <= not a;
    outputs(7029) <= not (a xor b);
    outputs(7030) <= not (a xor b);
    outputs(7031) <= not (a xor b);
    outputs(7032) <= not b or a;
    outputs(7033) <= b;
    outputs(7034) <= not (a or b);
    outputs(7035) <= a and b;
    outputs(7036) <= a xor b;
    outputs(7037) <= a xor b;
    outputs(7038) <= b;
    outputs(7039) <= a;
    outputs(7040) <= a;
    outputs(7041) <= not b or a;
    outputs(7042) <= not (a or b);
    outputs(7043) <= not (a or b);
    outputs(7044) <= not (a xor b);
    outputs(7045) <= not b;
    outputs(7046) <= not (a xor b);
    outputs(7047) <= b;
    outputs(7048) <= a;
    outputs(7049) <= a xor b;
    outputs(7050) <= not b;
    outputs(7051) <= a;
    outputs(7052) <= b and not a;
    outputs(7053) <= b;
    outputs(7054) <= not b;
    outputs(7055) <= a xor b;
    outputs(7056) <= not a;
    outputs(7057) <= not b;
    outputs(7058) <= a and b;
    outputs(7059) <= not (a xor b);
    outputs(7060) <= not (a xor b);
    outputs(7061) <= a or b;
    outputs(7062) <= not a;
    outputs(7063) <= not b;
    outputs(7064) <= a and b;
    outputs(7065) <= not (a xor b);
    outputs(7066) <= not b;
    outputs(7067) <= a and not b;
    outputs(7068) <= not b;
    outputs(7069) <= a and not b;
    outputs(7070) <= a xor b;
    outputs(7071) <= not (a xor b);
    outputs(7072) <= a xor b;
    outputs(7073) <= not b;
    outputs(7074) <= not (a or b);
    outputs(7075) <= not (a and b);
    outputs(7076) <= not a;
    outputs(7077) <= a xor b;
    outputs(7078) <= not b;
    outputs(7079) <= a xor b;
    outputs(7080) <= a xor b;
    outputs(7081) <= a xor b;
    outputs(7082) <= a;
    outputs(7083) <= a and b;
    outputs(7084) <= not b;
    outputs(7085) <= not a;
    outputs(7086) <= b;
    outputs(7087) <= not (a and b);
    outputs(7088) <= a xor b;
    outputs(7089) <= not (a or b);
    outputs(7090) <= not (a xor b);
    outputs(7091) <= not a;
    outputs(7092) <= a or b;
    outputs(7093) <= not b;
    outputs(7094) <= b;
    outputs(7095) <= not (a and b);
    outputs(7096) <= a xor b;
    outputs(7097) <= a xor b;
    outputs(7098) <= not b;
    outputs(7099) <= b;
    outputs(7100) <= not b;
    outputs(7101) <= a xor b;
    outputs(7102) <= a;
    outputs(7103) <= not a;
    outputs(7104) <= a;
    outputs(7105) <= a xor b;
    outputs(7106) <= not (a xor b);
    outputs(7107) <= not (a xor b);
    outputs(7108) <= not (a xor b);
    outputs(7109) <= a;
    outputs(7110) <= not (a xor b);
    outputs(7111) <= not (a xor b);
    outputs(7112) <= a;
    outputs(7113) <= a and not b;
    outputs(7114) <= b;
    outputs(7115) <= not a;
    outputs(7116) <= not (a xor b);
    outputs(7117) <= b;
    outputs(7118) <= a or b;
    outputs(7119) <= not b;
    outputs(7120) <= not (a xor b);
    outputs(7121) <= not (a xor b);
    outputs(7122) <= not a;
    outputs(7123) <= not (a xor b);
    outputs(7124) <= b;
    outputs(7125) <= not a;
    outputs(7126) <= a;
    outputs(7127) <= not (a or b);
    outputs(7128) <= a xor b;
    outputs(7129) <= not a;
    outputs(7130) <= not (a or b);
    outputs(7131) <= not a;
    outputs(7132) <= b;
    outputs(7133) <= not b;
    outputs(7134) <= not (a xor b);
    outputs(7135) <= a;
    outputs(7136) <= not (a xor b);
    outputs(7137) <= not (a and b);
    outputs(7138) <= a xor b;
    outputs(7139) <= not (a or b);
    outputs(7140) <= a or b;
    outputs(7141) <= a or b;
    outputs(7142) <= a and not b;
    outputs(7143) <= not a;
    outputs(7144) <= a xor b;
    outputs(7145) <= a xor b;
    outputs(7146) <= not a;
    outputs(7147) <= a xor b;
    outputs(7148) <= b;
    outputs(7149) <= not a;
    outputs(7150) <= not a;
    outputs(7151) <= b and not a;
    outputs(7152) <= not b;
    outputs(7153) <= not b;
    outputs(7154) <= b;
    outputs(7155) <= not b or a;
    outputs(7156) <= a xor b;
    outputs(7157) <= a xor b;
    outputs(7158) <= not (a xor b);
    outputs(7159) <= not (a xor b);
    outputs(7160) <= not (a xor b);
    outputs(7161) <= b;
    outputs(7162) <= not b;
    outputs(7163) <= not (a xor b);
    outputs(7164) <= a;
    outputs(7165) <= not (a or b);
    outputs(7166) <= not a;
    outputs(7167) <= a;
    outputs(7168) <= not a;
    outputs(7169) <= a and b;
    outputs(7170) <= not a or b;
    outputs(7171) <= not (a xor b);
    outputs(7172) <= not b;
    outputs(7173) <= b;
    outputs(7174) <= not b;
    outputs(7175) <= a xor b;
    outputs(7176) <= not (a xor b);
    outputs(7177) <= not b;
    outputs(7178) <= a and b;
    outputs(7179) <= a;
    outputs(7180) <= a xor b;
    outputs(7181) <= a xor b;
    outputs(7182) <= b and not a;
    outputs(7183) <= not a;
    outputs(7184) <= not (a xor b);
    outputs(7185) <= not (a xor b);
    outputs(7186) <= not a or b;
    outputs(7187) <= a;
    outputs(7188) <= a;
    outputs(7189) <= not (a xor b);
    outputs(7190) <= a xor b;
    outputs(7191) <= not b;
    outputs(7192) <= a;
    outputs(7193) <= not a or b;
    outputs(7194) <= a;
    outputs(7195) <= b and not a;
    outputs(7196) <= not b;
    outputs(7197) <= not b;
    outputs(7198) <= not (a xor b);
    outputs(7199) <= a xor b;
    outputs(7200) <= not (a xor b);
    outputs(7201) <= b and not a;
    outputs(7202) <= a xor b;
    outputs(7203) <= b;
    outputs(7204) <= a xor b;
    outputs(7205) <= a;
    outputs(7206) <= a xor b;
    outputs(7207) <= a xor b;
    outputs(7208) <= b and not a;
    outputs(7209) <= a or b;
    outputs(7210) <= not (a xor b);
    outputs(7211) <= not (a xor b);
    outputs(7212) <= a;
    outputs(7213) <= a or b;
    outputs(7214) <= a xor b;
    outputs(7215) <= not (a xor b);
    outputs(7216) <= not b;
    outputs(7217) <= a xor b;
    outputs(7218) <= b;
    outputs(7219) <= not (a xor b);
    outputs(7220) <= b;
    outputs(7221) <= b;
    outputs(7222) <= not a;
    outputs(7223) <= not a;
    outputs(7224) <= not a;
    outputs(7225) <= a xor b;
    outputs(7226) <= not a;
    outputs(7227) <= not (a xor b);
    outputs(7228) <= a and not b;
    outputs(7229) <= not (a xor b);
    outputs(7230) <= not (a xor b);
    outputs(7231) <= not a;
    outputs(7232) <= not b;
    outputs(7233) <= b;
    outputs(7234) <= not a;
    outputs(7235) <= a;
    outputs(7236) <= b;
    outputs(7237) <= a xor b;
    outputs(7238) <= a xor b;
    outputs(7239) <= b and not a;
    outputs(7240) <= a xor b;
    outputs(7241) <= a xor b;
    outputs(7242) <= a xor b;
    outputs(7243) <= a;
    outputs(7244) <= b;
    outputs(7245) <= not b;
    outputs(7246) <= not b;
    outputs(7247) <= not (a xor b);
    outputs(7248) <= not b;
    outputs(7249) <= not b;
    outputs(7250) <= a xor b;
    outputs(7251) <= not (a xor b);
    outputs(7252) <= a xor b;
    outputs(7253) <= not (a xor b);
    outputs(7254) <= not (a and b);
    outputs(7255) <= not (a xor b);
    outputs(7256) <= a;
    outputs(7257) <= a xor b;
    outputs(7258) <= b;
    outputs(7259) <= not (a xor b);
    outputs(7260) <= a or b;
    outputs(7261) <= a xor b;
    outputs(7262) <= not (a xor b);
    outputs(7263) <= not (a xor b);
    outputs(7264) <= a;
    outputs(7265) <= not a;
    outputs(7266) <= not b;
    outputs(7267) <= a xor b;
    outputs(7268) <= a;
    outputs(7269) <= not (a xor b);
    outputs(7270) <= a or b;
    outputs(7271) <= b;
    outputs(7272) <= not a;
    outputs(7273) <= not (a xor b);
    outputs(7274) <= a;
    outputs(7275) <= not b;
    outputs(7276) <= not (a xor b);
    outputs(7277) <= a;
    outputs(7278) <= a;
    outputs(7279) <= not b;
    outputs(7280) <= a and not b;
    outputs(7281) <= not a;
    outputs(7282) <= not (a xor b);
    outputs(7283) <= b;
    outputs(7284) <= not b;
    outputs(7285) <= not (a xor b);
    outputs(7286) <= b;
    outputs(7287) <= not a;
    outputs(7288) <= not a;
    outputs(7289) <= a xor b;
    outputs(7290) <= a xor b;
    outputs(7291) <= not b;
    outputs(7292) <= not a or b;
    outputs(7293) <= not b;
    outputs(7294) <= b;
    outputs(7295) <= not (a xor b);
    outputs(7296) <= not (a xor b);
    outputs(7297) <= not (a or b);
    outputs(7298) <= a xor b;
    outputs(7299) <= a xor b;
    outputs(7300) <= a;
    outputs(7301) <= a xor b;
    outputs(7302) <= not b;
    outputs(7303) <= not a;
    outputs(7304) <= not a;
    outputs(7305) <= a xor b;
    outputs(7306) <= a;
    outputs(7307) <= not a;
    outputs(7308) <= not (a xor b);
    outputs(7309) <= not (a xor b);
    outputs(7310) <= a;
    outputs(7311) <= not (a xor b);
    outputs(7312) <= b;
    outputs(7313) <= not (a xor b);
    outputs(7314) <= not a;
    outputs(7315) <= b;
    outputs(7316) <= not (a xor b);
    outputs(7317) <= not (a xor b);
    outputs(7318) <= a xor b;
    outputs(7319) <= b;
    outputs(7320) <= b;
    outputs(7321) <= a xor b;
    outputs(7322) <= a or b;
    outputs(7323) <= b and not a;
    outputs(7324) <= not (a or b);
    outputs(7325) <= b and not a;
    outputs(7326) <= not b or a;
    outputs(7327) <= not b;
    outputs(7328) <= a xor b;
    outputs(7329) <= a xor b;
    outputs(7330) <= a xor b;
    outputs(7331) <= not (a xor b);
    outputs(7332) <= b;
    outputs(7333) <= b;
    outputs(7334) <= a and not b;
    outputs(7335) <= a;
    outputs(7336) <= a xor b;
    outputs(7337) <= not a;
    outputs(7338) <= a and not b;
    outputs(7339) <= not b;
    outputs(7340) <= a;
    outputs(7341) <= not a;
    outputs(7342) <= not b;
    outputs(7343) <= not a;
    outputs(7344) <= a xor b;
    outputs(7345) <= a;
    outputs(7346) <= a xor b;
    outputs(7347) <= a;
    outputs(7348) <= b;
    outputs(7349) <= b;
    outputs(7350) <= not (a xor b);
    outputs(7351) <= not b or a;
    outputs(7352) <= not a;
    outputs(7353) <= a and not b;
    outputs(7354) <= not (a xor b);
    outputs(7355) <= not a;
    outputs(7356) <= a;
    outputs(7357) <= not b;
    outputs(7358) <= a xor b;
    outputs(7359) <= a xor b;
    outputs(7360) <= b;
    outputs(7361) <= a xor b;
    outputs(7362) <= a;
    outputs(7363) <= a;
    outputs(7364) <= a;
    outputs(7365) <= not a;
    outputs(7366) <= b;
    outputs(7367) <= a;
    outputs(7368) <= not (a xor b);
    outputs(7369) <= not b;
    outputs(7370) <= a;
    outputs(7371) <= a and b;
    outputs(7372) <= a and not b;
    outputs(7373) <= b;
    outputs(7374) <= a and not b;
    outputs(7375) <= not (a xor b);
    outputs(7376) <= not b;
    outputs(7377) <= not a;
    outputs(7378) <= not (a and b);
    outputs(7379) <= not (a xor b);
    outputs(7380) <= not (a xor b);
    outputs(7381) <= a xor b;
    outputs(7382) <= not (a xor b);
    outputs(7383) <= not a;
    outputs(7384) <= a and b;
    outputs(7385) <= a;
    outputs(7386) <= not (a xor b);
    outputs(7387) <= b;
    outputs(7388) <= a;
    outputs(7389) <= not b;
    outputs(7390) <= b and not a;
    outputs(7391) <= b;
    outputs(7392) <= a;
    outputs(7393) <= not a or b;
    outputs(7394) <= a and b;
    outputs(7395) <= a xor b;
    outputs(7396) <= not (a xor b);
    outputs(7397) <= a xor b;
    outputs(7398) <= not a;
    outputs(7399) <= a xor b;
    outputs(7400) <= a xor b;
    outputs(7401) <= not a;
    outputs(7402) <= a xor b;
    outputs(7403) <= a;
    outputs(7404) <= not a;
    outputs(7405) <= not b;
    outputs(7406) <= not (a xor b);
    outputs(7407) <= not a;
    outputs(7408) <= not b;
    outputs(7409) <= not (a xor b);
    outputs(7410) <= not (a xor b);
    outputs(7411) <= not a or b;
    outputs(7412) <= a and not b;
    outputs(7413) <= a and not b;
    outputs(7414) <= a;
    outputs(7415) <= not a;
    outputs(7416) <= b;
    outputs(7417) <= not b;
    outputs(7418) <= not (a xor b);
    outputs(7419) <= not (a xor b);
    outputs(7420) <= not (a xor b);
    outputs(7421) <= not a;
    outputs(7422) <= not a;
    outputs(7423) <= not b;
    outputs(7424) <= not (a xor b);
    outputs(7425) <= a xor b;
    outputs(7426) <= not a;
    outputs(7427) <= a and not b;
    outputs(7428) <= a;
    outputs(7429) <= not (a xor b);
    outputs(7430) <= a xor b;
    outputs(7431) <= a and not b;
    outputs(7432) <= a and not b;
    outputs(7433) <= not b or a;
    outputs(7434) <= not a;
    outputs(7435) <= a xor b;
    outputs(7436) <= not (a xor b);
    outputs(7437) <= a or b;
    outputs(7438) <= a xor b;
    outputs(7439) <= b;
    outputs(7440) <= a xor b;
    outputs(7441) <= not (a xor b);
    outputs(7442) <= not b;
    outputs(7443) <= a xor b;
    outputs(7444) <= not a;
    outputs(7445) <= not b;
    outputs(7446) <= a xor b;
    outputs(7447) <= not b;
    outputs(7448) <= not (a xor b);
    outputs(7449) <= not (a xor b);
    outputs(7450) <= b;
    outputs(7451) <= a xor b;
    outputs(7452) <= a xor b;
    outputs(7453) <= not a or b;
    outputs(7454) <= not b;
    outputs(7455) <= a xor b;
    outputs(7456) <= not a;
    outputs(7457) <= a xor b;
    outputs(7458) <= a xor b;
    outputs(7459) <= not (a or b);
    outputs(7460) <= not (a or b);
    outputs(7461) <= not (a or b);
    outputs(7462) <= not (a xor b);
    outputs(7463) <= not b;
    outputs(7464) <= not a or b;
    outputs(7465) <= a;
    outputs(7466) <= not a;
    outputs(7467) <= not b;
    outputs(7468) <= a and b;
    outputs(7469) <= a;
    outputs(7470) <= not a or b;
    outputs(7471) <= a;
    outputs(7472) <= not b;
    outputs(7473) <= a xor b;
    outputs(7474) <= a xor b;
    outputs(7475) <= not (a xor b);
    outputs(7476) <= not b;
    outputs(7477) <= a xor b;
    outputs(7478) <= a and not b;
    outputs(7479) <= not b;
    outputs(7480) <= a xor b;
    outputs(7481) <= a xor b;
    outputs(7482) <= not (a xor b);
    outputs(7483) <= a xor b;
    outputs(7484) <= not b;
    outputs(7485) <= not (a or b);
    outputs(7486) <= not a;
    outputs(7487) <= a;
    outputs(7488) <= a xor b;
    outputs(7489) <= not (a xor b);
    outputs(7490) <= b and not a;
    outputs(7491) <= b;
    outputs(7492) <= a and b;
    outputs(7493) <= a xor b;
    outputs(7494) <= a;
    outputs(7495) <= not a;
    outputs(7496) <= not a;
    outputs(7497) <= a;
    outputs(7498) <= not (a xor b);
    outputs(7499) <= a;
    outputs(7500) <= a;
    outputs(7501) <= a xor b;
    outputs(7502) <= a;
    outputs(7503) <= not (a xor b);
    outputs(7504) <= not (a and b);
    outputs(7505) <= a or b;
    outputs(7506) <= not (a xor b);
    outputs(7507) <= a;
    outputs(7508) <= a or b;
    outputs(7509) <= not b;
    outputs(7510) <= a xor b;
    outputs(7511) <= a;
    outputs(7512) <= not b or a;
    outputs(7513) <= not b;
    outputs(7514) <= not (a xor b);
    outputs(7515) <= not (a xor b);
    outputs(7516) <= a;
    outputs(7517) <= not b;
    outputs(7518) <= a;
    outputs(7519) <= a and b;
    outputs(7520) <= a xor b;
    outputs(7521) <= a xor b;
    outputs(7522) <= not (a and b);
    outputs(7523) <= not b;
    outputs(7524) <= not (a xor b);
    outputs(7525) <= b and not a;
    outputs(7526) <= not (a xor b);
    outputs(7527) <= not b;
    outputs(7528) <= a;
    outputs(7529) <= a or b;
    outputs(7530) <= b;
    outputs(7531) <= a xor b;
    outputs(7532) <= a xor b;
    outputs(7533) <= not (a xor b);
    outputs(7534) <= a xor b;
    outputs(7535) <= a xor b;
    outputs(7536) <= a xor b;
    outputs(7537) <= a;
    outputs(7538) <= a xor b;
    outputs(7539) <= not a;
    outputs(7540) <= not a;
    outputs(7541) <= not b or a;
    outputs(7542) <= a xor b;
    outputs(7543) <= a xor b;
    outputs(7544) <= a;
    outputs(7545) <= a;
    outputs(7546) <= a xor b;
    outputs(7547) <= a xor b;
    outputs(7548) <= not (a xor b);
    outputs(7549) <= b;
    outputs(7550) <= not (a or b);
    outputs(7551) <= not b;
    outputs(7552) <= b;
    outputs(7553) <= not (a or b);
    outputs(7554) <= a xor b;
    outputs(7555) <= not (a xor b);
    outputs(7556) <= not (a xor b);
    outputs(7557) <= a and not b;
    outputs(7558) <= a xor b;
    outputs(7559) <= a and b;
    outputs(7560) <= not (a xor b);
    outputs(7561) <= a xor b;
    outputs(7562) <= not b;
    outputs(7563) <= b;
    outputs(7564) <= not (a xor b);
    outputs(7565) <= a xor b;
    outputs(7566) <= b;
    outputs(7567) <= not a;
    outputs(7568) <= a;
    outputs(7569) <= b;
    outputs(7570) <= a xor b;
    outputs(7571) <= not b or a;
    outputs(7572) <= a xor b;
    outputs(7573) <= not b;
    outputs(7574) <= not b or a;
    outputs(7575) <= a;
    outputs(7576) <= not (a xor b);
    outputs(7577) <= not a;
    outputs(7578) <= a xor b;
    outputs(7579) <= b;
    outputs(7580) <= a and not b;
    outputs(7581) <= a and not b;
    outputs(7582) <= a xor b;
    outputs(7583) <= not (a xor b);
    outputs(7584) <= not a;
    outputs(7585) <= not b;
    outputs(7586) <= not (a and b);
    outputs(7587) <= not b;
    outputs(7588) <= not a;
    outputs(7589) <= not a;
    outputs(7590) <= not a or b;
    outputs(7591) <= not a;
    outputs(7592) <= b and not a;
    outputs(7593) <= a xor b;
    outputs(7594) <= not a;
    outputs(7595) <= not (a xor b);
    outputs(7596) <= not b;
    outputs(7597) <= a and b;
    outputs(7598) <= not (a xor b);
    outputs(7599) <= b;
    outputs(7600) <= a and b;
    outputs(7601) <= b;
    outputs(7602) <= not (a xor b);
    outputs(7603) <= a and not b;
    outputs(7604) <= not (a xor b);
    outputs(7605) <= not (a xor b);
    outputs(7606) <= a;
    outputs(7607) <= b;
    outputs(7608) <= a xor b;
    outputs(7609) <= a;
    outputs(7610) <= a;
    outputs(7611) <= a or b;
    outputs(7612) <= b;
    outputs(7613) <= not b;
    outputs(7614) <= a and b;
    outputs(7615) <= a;
    outputs(7616) <= not b;
    outputs(7617) <= not (a xor b);
    outputs(7618) <= not b;
    outputs(7619) <= a xor b;
    outputs(7620) <= not a;
    outputs(7621) <= not a;
    outputs(7622) <= a and not b;
    outputs(7623) <= not b;
    outputs(7624) <= a xor b;
    outputs(7625) <= a xor b;
    outputs(7626) <= a xor b;
    outputs(7627) <= not (a xor b);
    outputs(7628) <= b and not a;
    outputs(7629) <= not (a and b);
    outputs(7630) <= not (a and b);
    outputs(7631) <= b and not a;
    outputs(7632) <= a xor b;
    outputs(7633) <= not b or a;
    outputs(7634) <= not (a or b);
    outputs(7635) <= a xor b;
    outputs(7636) <= not (a or b);
    outputs(7637) <= not (a xor b);
    outputs(7638) <= a;
    outputs(7639) <= not (a xor b);
    outputs(7640) <= a xor b;
    outputs(7641) <= a or b;
    outputs(7642) <= not (a xor b);
    outputs(7643) <= a;
    outputs(7644) <= a and b;
    outputs(7645) <= not (a xor b);
    outputs(7646) <= not (a and b);
    outputs(7647) <= b;
    outputs(7648) <= a xor b;
    outputs(7649) <= a;
    outputs(7650) <= not b;
    outputs(7651) <= b;
    outputs(7652) <= b and not a;
    outputs(7653) <= not b;
    outputs(7654) <= a xor b;
    outputs(7655) <= a;
    outputs(7656) <= b;
    outputs(7657) <= a xor b;
    outputs(7658) <= not a;
    outputs(7659) <= not b;
    outputs(7660) <= a xor b;
    outputs(7661) <= not b;
    outputs(7662) <= a xor b;
    outputs(7663) <= a and not b;
    outputs(7664) <= not (a xor b);
    outputs(7665) <= not b;
    outputs(7666) <= not (a xor b);
    outputs(7667) <= not (a xor b);
    outputs(7668) <= not a or b;
    outputs(7669) <= not (a or b);
    outputs(7670) <= a and b;
    outputs(7671) <= b;
    outputs(7672) <= not b;
    outputs(7673) <= not (a xor b);
    outputs(7674) <= a or b;
    outputs(7675) <= a and b;
    outputs(7676) <= not b;
    outputs(7677) <= not b;
    outputs(7678) <= a xor b;
    outputs(7679) <= a and b;
    outputs(7680) <= a or b;
    outputs(7681) <= a xor b;
    outputs(7682) <= b;
    outputs(7683) <= not (a or b);
    outputs(7684) <= a xor b;
    outputs(7685) <= not (a xor b);
    outputs(7686) <= not a;
    outputs(7687) <= a xor b;
    outputs(7688) <= a;
    outputs(7689) <= a;
    outputs(7690) <= a;
    outputs(7691) <= not (a xor b);
    outputs(7692) <= not (a xor b);
    outputs(7693) <= b;
    outputs(7694) <= not (a or b);
    outputs(7695) <= not (a xor b);
    outputs(7696) <= a;
    outputs(7697) <= not (a or b);
    outputs(7698) <= not a;
    outputs(7699) <= a and b;
    outputs(7700) <= a xor b;
    outputs(7701) <= b;
    outputs(7702) <= a xor b;
    outputs(7703) <= a;
    outputs(7704) <= not (a xor b);
    outputs(7705) <= b;
    outputs(7706) <= not b;
    outputs(7707) <= not (a or b);
    outputs(7708) <= a and not b;
    outputs(7709) <= not b;
    outputs(7710) <= not (a xor b);
    outputs(7711) <= b and not a;
    outputs(7712) <= not a;
    outputs(7713) <= not (a xor b);
    outputs(7714) <= a or b;
    outputs(7715) <= not a;
    outputs(7716) <= a and b;
    outputs(7717) <= a;
    outputs(7718) <= b;
    outputs(7719) <= not (a xor b);
    outputs(7720) <= not a;
    outputs(7721) <= not (a xor b);
    outputs(7722) <= a;
    outputs(7723) <= b;
    outputs(7724) <= a and b;
    outputs(7725) <= not (a xor b);
    outputs(7726) <= not (a xor b);
    outputs(7727) <= a;
    outputs(7728) <= a;
    outputs(7729) <= not b;
    outputs(7730) <= not b;
    outputs(7731) <= b;
    outputs(7732) <= a or b;
    outputs(7733) <= a xor b;
    outputs(7734) <= not b;
    outputs(7735) <= a xor b;
    outputs(7736) <= a;
    outputs(7737) <= a;
    outputs(7738) <= a or b;
    outputs(7739) <= a or b;
    outputs(7740) <= b;
    outputs(7741) <= a;
    outputs(7742) <= not (a xor b);
    outputs(7743) <= a or b;
    outputs(7744) <= a;
    outputs(7745) <= not a;
    outputs(7746) <= a;
    outputs(7747) <= b;
    outputs(7748) <= not b or a;
    outputs(7749) <= a and b;
    outputs(7750) <= a xor b;
    outputs(7751) <= not (a xor b);
    outputs(7752) <= a;
    outputs(7753) <= not b;
    outputs(7754) <= not a;
    outputs(7755) <= not a;
    outputs(7756) <= a or b;
    outputs(7757) <= b;
    outputs(7758) <= a xor b;
    outputs(7759) <= b;
    outputs(7760) <= not b or a;
    outputs(7761) <= not (a or b);
    outputs(7762) <= not b;
    outputs(7763) <= not b;
    outputs(7764) <= not b;
    outputs(7765) <= not b;
    outputs(7766) <= not b;
    outputs(7767) <= b and not a;
    outputs(7768) <= not b;
    outputs(7769) <= a;
    outputs(7770) <= b and not a;
    outputs(7771) <= a;
    outputs(7772) <= not (a xor b);
    outputs(7773) <= not a;
    outputs(7774) <= not b;
    outputs(7775) <= b and not a;
    outputs(7776) <= not a;
    outputs(7777) <= not b;
    outputs(7778) <= not a;
    outputs(7779) <= not b;
    outputs(7780) <= not a or b;
    outputs(7781) <= a and b;
    outputs(7782) <= a;
    outputs(7783) <= b and not a;
    outputs(7784) <= not a;
    outputs(7785) <= a;
    outputs(7786) <= b and not a;
    outputs(7787) <= b and not a;
    outputs(7788) <= b;
    outputs(7789) <= a;
    outputs(7790) <= not a;
    outputs(7791) <= a and not b;
    outputs(7792) <= b and not a;
    outputs(7793) <= not b;
    outputs(7794) <= a xor b;
    outputs(7795) <= not (a and b);
    outputs(7796) <= b;
    outputs(7797) <= b and not a;
    outputs(7798) <= b and not a;
    outputs(7799) <= not (a xor b);
    outputs(7800) <= b;
    outputs(7801) <= not a;
    outputs(7802) <= not (a and b);
    outputs(7803) <= b and not a;
    outputs(7804) <= not b;
    outputs(7805) <= not (a xor b);
    outputs(7806) <= not b or a;
    outputs(7807) <= a xor b;
    outputs(7808) <= a;
    outputs(7809) <= not (a or b);
    outputs(7810) <= a xor b;
    outputs(7811) <= not a;
    outputs(7812) <= a xor b;
    outputs(7813) <= a xor b;
    outputs(7814) <= a and not b;
    outputs(7815) <= a xor b;
    outputs(7816) <= b;
    outputs(7817) <= not a;
    outputs(7818) <= b;
    outputs(7819) <= b;
    outputs(7820) <= not a;
    outputs(7821) <= a xor b;
    outputs(7822) <= not a;
    outputs(7823) <= b and not a;
    outputs(7824) <= not a;
    outputs(7825) <= not b or a;
    outputs(7826) <= a xor b;
    outputs(7827) <= not a;
    outputs(7828) <= a;
    outputs(7829) <= not a;
    outputs(7830) <= not b;
    outputs(7831) <= b;
    outputs(7832) <= a;
    outputs(7833) <= not b;
    outputs(7834) <= not a;
    outputs(7835) <= a and not b;
    outputs(7836) <= b and not a;
    outputs(7837) <= a and b;
    outputs(7838) <= not a or b;
    outputs(7839) <= a;
    outputs(7840) <= a;
    outputs(7841) <= a xor b;
    outputs(7842) <= not a;
    outputs(7843) <= not a or b;
    outputs(7844) <= a or b;
    outputs(7845) <= not a or b;
    outputs(7846) <= a xor b;
    outputs(7847) <= a xor b;
    outputs(7848) <= a xor b;
    outputs(7849) <= not (a xor b);
    outputs(7850) <= a and b;
    outputs(7851) <= b and not a;
    outputs(7852) <= a;
    outputs(7853) <= a and b;
    outputs(7854) <= a;
    outputs(7855) <= a;
    outputs(7856) <= b;
    outputs(7857) <= a xor b;
    outputs(7858) <= a;
    outputs(7859) <= a;
    outputs(7860) <= b;
    outputs(7861) <= a xor b;
    outputs(7862) <= b;
    outputs(7863) <= a and not b;
    outputs(7864) <= not a;
    outputs(7865) <= b and not a;
    outputs(7866) <= a and b;
    outputs(7867) <= not a;
    outputs(7868) <= not (a xor b);
    outputs(7869) <= a and not b;
    outputs(7870) <= b and not a;
    outputs(7871) <= not (a xor b);
    outputs(7872) <= a;
    outputs(7873) <= a xor b;
    outputs(7874) <= not (a or b);
    outputs(7875) <= b;
    outputs(7876) <= not (a or b);
    outputs(7877) <= not b;
    outputs(7878) <= not (a xor b);
    outputs(7879) <= not b;
    outputs(7880) <= a xor b;
    outputs(7881) <= b;
    outputs(7882) <= a and b;
    outputs(7883) <= a;
    outputs(7884) <= not b;
    outputs(7885) <= b;
    outputs(7886) <= not (a or b);
    outputs(7887) <= not a or b;
    outputs(7888) <= not b;
    outputs(7889) <= a;
    outputs(7890) <= not a;
    outputs(7891) <= not b;
    outputs(7892) <= not (a xor b);
    outputs(7893) <= a xor b;
    outputs(7894) <= a xor b;
    outputs(7895) <= not (a xor b);
    outputs(7896) <= b;
    outputs(7897) <= b;
    outputs(7898) <= not b;
    outputs(7899) <= a xor b;
    outputs(7900) <= b;
    outputs(7901) <= b and not a;
    outputs(7902) <= a and b;
    outputs(7903) <= a;
    outputs(7904) <= not (a or b);
    outputs(7905) <= not a;
    outputs(7906) <= a;
    outputs(7907) <= a;
    outputs(7908) <= a xor b;
    outputs(7909) <= not (a xor b);
    outputs(7910) <= a and b;
    outputs(7911) <= a and b;
    outputs(7912) <= b and not a;
    outputs(7913) <= b;
    outputs(7914) <= not a;
    outputs(7915) <= not (a or b);
    outputs(7916) <= a;
    outputs(7917) <= a xor b;
    outputs(7918) <= a xor b;
    outputs(7919) <= not a or b;
    outputs(7920) <= a xor b;
    outputs(7921) <= not (a xor b);
    outputs(7922) <= b;
    outputs(7923) <= not a;
    outputs(7924) <= not (a xor b);
    outputs(7925) <= not b;
    outputs(7926) <= a and not b;
    outputs(7927) <= not a;
    outputs(7928) <= a xor b;
    outputs(7929) <= not (a xor b);
    outputs(7930) <= not a;
    outputs(7931) <= not a;
    outputs(7932) <= a xor b;
    outputs(7933) <= a;
    outputs(7934) <= not (a xor b);
    outputs(7935) <= b;
    outputs(7936) <= a;
    outputs(7937) <= not (a xor b);
    outputs(7938) <= b;
    outputs(7939) <= a;
    outputs(7940) <= a xor b;
    outputs(7941) <= not b;
    outputs(7942) <= not (a xor b);
    outputs(7943) <= not a;
    outputs(7944) <= a xor b;
    outputs(7945) <= b;
    outputs(7946) <= a and b;
    outputs(7947) <= a xor b;
    outputs(7948) <= not a;
    outputs(7949) <= a and not b;
    outputs(7950) <= not a;
    outputs(7951) <= b;
    outputs(7952) <= not (a or b);
    outputs(7953) <= not b or a;
    outputs(7954) <= not (a xor b);
    outputs(7955) <= not b;
    outputs(7956) <= not a;
    outputs(7957) <= not (a xor b);
    outputs(7958) <= not b or a;
    outputs(7959) <= a and b;
    outputs(7960) <= not (a xor b);
    outputs(7961) <= b;
    outputs(7962) <= not (a or b);
    outputs(7963) <= a or b;
    outputs(7964) <= a xor b;
    outputs(7965) <= a xor b;
    outputs(7966) <= b;
    outputs(7967) <= b and not a;
    outputs(7968) <= a or b;
    outputs(7969) <= a xor b;
    outputs(7970) <= not b;
    outputs(7971) <= not (a and b);
    outputs(7972) <= not a;
    outputs(7973) <= b;
    outputs(7974) <= a or b;
    outputs(7975) <= not (a xor b);
    outputs(7976) <= a;
    outputs(7977) <= not a;
    outputs(7978) <= not a;
    outputs(7979) <= b and not a;
    outputs(7980) <= a;
    outputs(7981) <= a;
    outputs(7982) <= not a;
    outputs(7983) <= not (a or b);
    outputs(7984) <= not (a xor b);
    outputs(7985) <= not (a xor b);
    outputs(7986) <= b;
    outputs(7987) <= not b;
    outputs(7988) <= a xor b;
    outputs(7989) <= not b;
    outputs(7990) <= b and not a;
    outputs(7991) <= not b;
    outputs(7992) <= a or b;
    outputs(7993) <= not a;
    outputs(7994) <= not a;
    outputs(7995) <= a;
    outputs(7996) <= b;
    outputs(7997) <= not a;
    outputs(7998) <= not b;
    outputs(7999) <= a xor b;
    outputs(8000) <= not b;
    outputs(8001) <= not (a or b);
    outputs(8002) <= not b;
    outputs(8003) <= not a;
    outputs(8004) <= not (a and b);
    outputs(8005) <= not (a xor b);
    outputs(8006) <= a;
    outputs(8007) <= not (a xor b);
    outputs(8008) <= not a;
    outputs(8009) <= not (a xor b);
    outputs(8010) <= not (a and b);
    outputs(8011) <= not a or b;
    outputs(8012) <= not b;
    outputs(8013) <= not a;
    outputs(8014) <= not a;
    outputs(8015) <= not a;
    outputs(8016) <= not (a xor b);
    outputs(8017) <= a;
    outputs(8018) <= not (a and b);
    outputs(8019) <= b and not a;
    outputs(8020) <= b;
    outputs(8021) <= not a;
    outputs(8022) <= not b;
    outputs(8023) <= a xor b;
    outputs(8024) <= a xor b;
    outputs(8025) <= b and not a;
    outputs(8026) <= not a;
    outputs(8027) <= b and not a;
    outputs(8028) <= not b;
    outputs(8029) <= a;
    outputs(8030) <= a;
    outputs(8031) <= b;
    outputs(8032) <= not a;
    outputs(8033) <= not b;
    outputs(8034) <= not a;
    outputs(8035) <= not a;
    outputs(8036) <= a;
    outputs(8037) <= b;
    outputs(8038) <= b;
    outputs(8039) <= not a;
    outputs(8040) <= not a;
    outputs(8041) <= b;
    outputs(8042) <= a xor b;
    outputs(8043) <= not (a xor b);
    outputs(8044) <= not b;
    outputs(8045) <= not (a xor b);
    outputs(8046) <= not a or b;
    outputs(8047) <= b and not a;
    outputs(8048) <= not (a or b);
    outputs(8049) <= a;
    outputs(8050) <= a;
    outputs(8051) <= not b;
    outputs(8052) <= not b;
    outputs(8053) <= b;
    outputs(8054) <= b;
    outputs(8055) <= not (a xor b);
    outputs(8056) <= a and b;
    outputs(8057) <= b;
    outputs(8058) <= not (a or b);
    outputs(8059) <= b and not a;
    outputs(8060) <= not (a xor b);
    outputs(8061) <= b;
    outputs(8062) <= not (a xor b);
    outputs(8063) <= not (a xor b);
    outputs(8064) <= not a;
    outputs(8065) <= b;
    outputs(8066) <= b;
    outputs(8067) <= not b;
    outputs(8068) <= b and not a;
    outputs(8069) <= a;
    outputs(8070) <= a xor b;
    outputs(8071) <= not (a xor b);
    outputs(8072) <= a;
    outputs(8073) <= not b;
    outputs(8074) <= b;
    outputs(8075) <= not b;
    outputs(8076) <= not b;
    outputs(8077) <= a and b;
    outputs(8078) <= b;
    outputs(8079) <= not b or a;
    outputs(8080) <= not (a xor b);
    outputs(8081) <= a xor b;
    outputs(8082) <= b;
    outputs(8083) <= a xor b;
    outputs(8084) <= not a;
    outputs(8085) <= not a;
    outputs(8086) <= a and not b;
    outputs(8087) <= a;
    outputs(8088) <= a;
    outputs(8089) <= not a;
    outputs(8090) <= a or b;
    outputs(8091) <= not a;
    outputs(8092) <= a;
    outputs(8093) <= a and b;
    outputs(8094) <= b;
    outputs(8095) <= b;
    outputs(8096) <= not a;
    outputs(8097) <= a;
    outputs(8098) <= a;
    outputs(8099) <= not b;
    outputs(8100) <= not (a xor b);
    outputs(8101) <= not a or b;
    outputs(8102) <= not b or a;
    outputs(8103) <= not (a xor b);
    outputs(8104) <= a or b;
    outputs(8105) <= b;
    outputs(8106) <= a;
    outputs(8107) <= a;
    outputs(8108) <= not a;
    outputs(8109) <= not a;
    outputs(8110) <= not a;
    outputs(8111) <= b;
    outputs(8112) <= not (a xor b);
    outputs(8113) <= a;
    outputs(8114) <= a;
    outputs(8115) <= not a or b;
    outputs(8116) <= not a;
    outputs(8117) <= a;
    outputs(8118) <= a;
    outputs(8119) <= not b;
    outputs(8120) <= b;
    outputs(8121) <= not (a or b);
    outputs(8122) <= not a;
    outputs(8123) <= not (a xor b);
    outputs(8124) <= not a;
    outputs(8125) <= not a;
    outputs(8126) <= a;
    outputs(8127) <= not (a xor b);
    outputs(8128) <= a and not b;
    outputs(8129) <= not a;
    outputs(8130) <= a;
    outputs(8131) <= not a;
    outputs(8132) <= a and b;
    outputs(8133) <= a;
    outputs(8134) <= not (a xor b);
    outputs(8135) <= a xor b;
    outputs(8136) <= a;
    outputs(8137) <= a xor b;
    outputs(8138) <= not (a xor b);
    outputs(8139) <= not (a xor b);
    outputs(8140) <= a and not b;
    outputs(8141) <= a xor b;
    outputs(8142) <= a and b;
    outputs(8143) <= a xor b;
    outputs(8144) <= not b;
    outputs(8145) <= b;
    outputs(8146) <= a xor b;
    outputs(8147) <= not b;
    outputs(8148) <= a;
    outputs(8149) <= a and b;
    outputs(8150) <= b;
    outputs(8151) <= not a;
    outputs(8152) <= b and not a;
    outputs(8153) <= not b;
    outputs(8154) <= not a or b;
    outputs(8155) <= a and not b;
    outputs(8156) <= not b;
    outputs(8157) <= a;
    outputs(8158) <= a and b;
    outputs(8159) <= not (a or b);
    outputs(8160) <= a xor b;
    outputs(8161) <= a;
    outputs(8162) <= a;
    outputs(8163) <= a or b;
    outputs(8164) <= a xor b;
    outputs(8165) <= not b;
    outputs(8166) <= not a;
    outputs(8167) <= not b;
    outputs(8168) <= a and not b;
    outputs(8169) <= a and b;
    outputs(8170) <= a;
    outputs(8171) <= not (a xor b);
    outputs(8172) <= a xor b;
    outputs(8173) <= not b;
    outputs(8174) <= a xor b;
    outputs(8175) <= b;
    outputs(8176) <= not b or a;
    outputs(8177) <= not b;
    outputs(8178) <= b;
    outputs(8179) <= not a;
    outputs(8180) <= a and not b;
    outputs(8181) <= a and not b;
    outputs(8182) <= not (a and b);
    outputs(8183) <= a xor b;
    outputs(8184) <= b;
    outputs(8185) <= not b or a;
    outputs(8186) <= not (a xor b);
    outputs(8187) <= not b;
    outputs(8188) <= a;
    outputs(8189) <= not b;
    outputs(8190) <= b;
    outputs(8191) <= not b or a;
    outputs(8192) <= not b or a;
    outputs(8193) <= b;
    outputs(8194) <= not (a or b);
    outputs(8195) <= not b;
    outputs(8196) <= b;
    outputs(8197) <= a;
    outputs(8198) <= a and not b;
    outputs(8199) <= a xor b;
    outputs(8200) <= not (a xor b);
    outputs(8201) <= not a;
    outputs(8202) <= a;
    outputs(8203) <= not b or a;
    outputs(8204) <= not (a xor b);
    outputs(8205) <= not a;
    outputs(8206) <= not (a xor b);
    outputs(8207) <= b;
    outputs(8208) <= not (a or b);
    outputs(8209) <= not (a xor b);
    outputs(8210) <= not (a xor b);
    outputs(8211) <= a;
    outputs(8212) <= not (a xor b);
    outputs(8213) <= not (a xor b);
    outputs(8214) <= not a;
    outputs(8215) <= not (a or b);
    outputs(8216) <= b;
    outputs(8217) <= a;
    outputs(8218) <= a xor b;
    outputs(8219) <= b;
    outputs(8220) <= not a;
    outputs(8221) <= not b;
    outputs(8222) <= not a;
    outputs(8223) <= not (a xor b);
    outputs(8224) <= a xor b;
    outputs(8225) <= a xor b;
    outputs(8226) <= a xor b;
    outputs(8227) <= a or b;
    outputs(8228) <= not a;
    outputs(8229) <= b;
    outputs(8230) <= a or b;
    outputs(8231) <= a;
    outputs(8232) <= not (a xor b);
    outputs(8233) <= not (a xor b);
    outputs(8234) <= b;
    outputs(8235) <= a;
    outputs(8236) <= b;
    outputs(8237) <= not (a or b);
    outputs(8238) <= b;
    outputs(8239) <= not (a xor b);
    outputs(8240) <= b and not a;
    outputs(8241) <= not (a xor b);
    outputs(8242) <= not (a or b);
    outputs(8243) <= not (a xor b);
    outputs(8244) <= b;
    outputs(8245) <= a or b;
    outputs(8246) <= not a;
    outputs(8247) <= not b;
    outputs(8248) <= b and not a;
    outputs(8249) <= a and not b;
    outputs(8250) <= not a;
    outputs(8251) <= not (a or b);
    outputs(8252) <= a;
    outputs(8253) <= not a;
    outputs(8254) <= not (a xor b);
    outputs(8255) <= not b;
    outputs(8256) <= b;
    outputs(8257) <= a or b;
    outputs(8258) <= not b or a;
    outputs(8259) <= a and b;
    outputs(8260) <= a xor b;
    outputs(8261) <= not (a xor b);
    outputs(8262) <= a;
    outputs(8263) <= b;
    outputs(8264) <= a;
    outputs(8265) <= not (a xor b);
    outputs(8266) <= a xor b;
    outputs(8267) <= not (a xor b);
    outputs(8268) <= not a;
    outputs(8269) <= not (a xor b);
    outputs(8270) <= not b;
    outputs(8271) <= a and not b;
    outputs(8272) <= not b or a;
    outputs(8273) <= a and b;
    outputs(8274) <= a and not b;
    outputs(8275) <= b;
    outputs(8276) <= b;
    outputs(8277) <= not b or a;
    outputs(8278) <= a xor b;
    outputs(8279) <= b and not a;
    outputs(8280) <= b;
    outputs(8281) <= not b;
    outputs(8282) <= not (a and b);
    outputs(8283) <= a xor b;
    outputs(8284) <= not (a xor b);
    outputs(8285) <= not a;
    outputs(8286) <= b and not a;
    outputs(8287) <= not b;
    outputs(8288) <= b;
    outputs(8289) <= not (a xor b);
    outputs(8290) <= not a;
    outputs(8291) <= a xor b;
    outputs(8292) <= not b;
    outputs(8293) <= b;
    outputs(8294) <= not (a xor b);
    outputs(8295) <= a;
    outputs(8296) <= b;
    outputs(8297) <= not b;
    outputs(8298) <= not a;
    outputs(8299) <= not a;
    outputs(8300) <= not a;
    outputs(8301) <= not b;
    outputs(8302) <= a xor b;
    outputs(8303) <= b and not a;
    outputs(8304) <= a xor b;
    outputs(8305) <= a and not b;
    outputs(8306) <= not a;
    outputs(8307) <= b;
    outputs(8308) <= a;
    outputs(8309) <= not (a xor b);
    outputs(8310) <= a;
    outputs(8311) <= a xor b;
    outputs(8312) <= b;
    outputs(8313) <= a;
    outputs(8314) <= not b;
    outputs(8315) <= a and b;
    outputs(8316) <= a and not b;
    outputs(8317) <= not b;
    outputs(8318) <= a xor b;
    outputs(8319) <= b and not a;
    outputs(8320) <= b;
    outputs(8321) <= not (a xor b);
    outputs(8322) <= not a;
    outputs(8323) <= not a;
    outputs(8324) <= a or b;
    outputs(8325) <= b;
    outputs(8326) <= a xor b;
    outputs(8327) <= not (a xor b);
    outputs(8328) <= b;
    outputs(8329) <= not (a and b);
    outputs(8330) <= b;
    outputs(8331) <= a xor b;
    outputs(8332) <= not (a xor b);
    outputs(8333) <= not b;
    outputs(8334) <= b;
    outputs(8335) <= b;
    outputs(8336) <= b;
    outputs(8337) <= not (a xor b);
    outputs(8338) <= b;
    outputs(8339) <= a xor b;
    outputs(8340) <= not (a xor b);
    outputs(8341) <= not (a or b);
    outputs(8342) <= not (a xor b);
    outputs(8343) <= not a;
    outputs(8344) <= b;
    outputs(8345) <= not a;
    outputs(8346) <= a and not b;
    outputs(8347) <= not a;
    outputs(8348) <= a xor b;
    outputs(8349) <= a and not b;
    outputs(8350) <= b and not a;
    outputs(8351) <= b and not a;
    outputs(8352) <= not a;
    outputs(8353) <= b;
    outputs(8354) <= a and b;
    outputs(8355) <= a xor b;
    outputs(8356) <= not (a or b);
    outputs(8357) <= not a;
    outputs(8358) <= not a;
    outputs(8359) <= a xor b;
    outputs(8360) <= b and not a;
    outputs(8361) <= a xor b;
    outputs(8362) <= not a;
    outputs(8363) <= a or b;
    outputs(8364) <= a or b;
    outputs(8365) <= b;
    outputs(8366) <= not a;
    outputs(8367) <= a;
    outputs(8368) <= not (a xor b);
    outputs(8369) <= a;
    outputs(8370) <= not (a or b);
    outputs(8371) <= not (a xor b);
    outputs(8372) <= a;
    outputs(8373) <= a xor b;
    outputs(8374) <= a xor b;
    outputs(8375) <= a;
    outputs(8376) <= not b;
    outputs(8377) <= not a;
    outputs(8378) <= not a;
    outputs(8379) <= b;
    outputs(8380) <= not a or b;
    outputs(8381) <= a xor b;
    outputs(8382) <= not (a and b);
    outputs(8383) <= not b;
    outputs(8384) <= a;
    outputs(8385) <= not b;
    outputs(8386) <= a and b;
    outputs(8387) <= not b;
    outputs(8388) <= a xor b;
    outputs(8389) <= a xor b;
    outputs(8390) <= not (a xor b);
    outputs(8391) <= not b or a;
    outputs(8392) <= a;
    outputs(8393) <= not a;
    outputs(8394) <= a;
    outputs(8395) <= b;
    outputs(8396) <= a xor b;
    outputs(8397) <= b and not a;
    outputs(8398) <= not b;
    outputs(8399) <= a xor b;
    outputs(8400) <= not (a xor b);
    outputs(8401) <= not a;
    outputs(8402) <= a xor b;
    outputs(8403) <= b and not a;
    outputs(8404) <= a xor b;
    outputs(8405) <= b and not a;
    outputs(8406) <= b;
    outputs(8407) <= a;
    outputs(8408) <= a and b;
    outputs(8409) <= not (a xor b);
    outputs(8410) <= not a;
    outputs(8411) <= not b;
    outputs(8412) <= not (a and b);
    outputs(8413) <= not a;
    outputs(8414) <= a;
    outputs(8415) <= not b;
    outputs(8416) <= not a;
    outputs(8417) <= not (a xor b);
    outputs(8418) <= not (a xor b);
    outputs(8419) <= b and not a;
    outputs(8420) <= not a;
    outputs(8421) <= a;
    outputs(8422) <= b and not a;
    outputs(8423) <= a xor b;
    outputs(8424) <= b;
    outputs(8425) <= a;
    outputs(8426) <= a xor b;
    outputs(8427) <= a xor b;
    outputs(8428) <= not a;
    outputs(8429) <= a or b;
    outputs(8430) <= not a or b;
    outputs(8431) <= b;
    outputs(8432) <= not a;
    outputs(8433) <= a;
    outputs(8434) <= a and b;
    outputs(8435) <= b;
    outputs(8436) <= not b;
    outputs(8437) <= not a;
    outputs(8438) <= a and b;
    outputs(8439) <= b;
    outputs(8440) <= not (a xor b);
    outputs(8441) <= a and b;
    outputs(8442) <= a;
    outputs(8443) <= a and b;
    outputs(8444) <= not b;
    outputs(8445) <= not b or a;
    outputs(8446) <= b and not a;
    outputs(8447) <= b;
    outputs(8448) <= not (a xor b);
    outputs(8449) <= not (a xor b);
    outputs(8450) <= not b;
    outputs(8451) <= a;
    outputs(8452) <= not (a xor b);
    outputs(8453) <= not b;
    outputs(8454) <= not (a or b);
    outputs(8455) <= a;
    outputs(8456) <= not b;
    outputs(8457) <= b;
    outputs(8458) <= not (a and b);
    outputs(8459) <= b;
    outputs(8460) <= not a;
    outputs(8461) <= a and b;
    outputs(8462) <= not a;
    outputs(8463) <= b and not a;
    outputs(8464) <= a and not b;
    outputs(8465) <= a xor b;
    outputs(8466) <= a;
    outputs(8467) <= b;
    outputs(8468) <= not (a xor b);
    outputs(8469) <= b;
    outputs(8470) <= a or b;
    outputs(8471) <= a;
    outputs(8472) <= not (a xor b);
    outputs(8473) <= a xor b;
    outputs(8474) <= not b;
    outputs(8475) <= a xor b;
    outputs(8476) <= a;
    outputs(8477) <= b;
    outputs(8478) <= not b;
    outputs(8479) <= not b;
    outputs(8480) <= b;
    outputs(8481) <= b;
    outputs(8482) <= b;
    outputs(8483) <= not (a and b);
    outputs(8484) <= not (a or b);
    outputs(8485) <= not (a or b);
    outputs(8486) <= not a;
    outputs(8487) <= not a;
    outputs(8488) <= not a or b;
    outputs(8489) <= not a or b;
    outputs(8490) <= b;
    outputs(8491) <= not b;
    outputs(8492) <= not b or a;
    outputs(8493) <= a or b;
    outputs(8494) <= a;
    outputs(8495) <= not b;
    outputs(8496) <= a xor b;
    outputs(8497) <= a or b;
    outputs(8498) <= not b;
    outputs(8499) <= a;
    outputs(8500) <= a;
    outputs(8501) <= b and not a;
    outputs(8502) <= b;
    outputs(8503) <= not b;
    outputs(8504) <= a and b;
    outputs(8505) <= not b;
    outputs(8506) <= not (a xor b);
    outputs(8507) <= not b;
    outputs(8508) <= a xor b;
    outputs(8509) <= not a or b;
    outputs(8510) <= b;
    outputs(8511) <= not a or b;
    outputs(8512) <= a;
    outputs(8513) <= not b;
    outputs(8514) <= b;
    outputs(8515) <= a and b;
    outputs(8516) <= a xor b;
    outputs(8517) <= not a;
    outputs(8518) <= not (a xor b);
    outputs(8519) <= a and not b;
    outputs(8520) <= not a;
    outputs(8521) <= not a;
    outputs(8522) <= b;
    outputs(8523) <= not (a xor b);
    outputs(8524) <= a and b;
    outputs(8525) <= not a;
    outputs(8526) <= not (a xor b);
    outputs(8527) <= not b;
    outputs(8528) <= not a;
    outputs(8529) <= not a;
    outputs(8530) <= b;
    outputs(8531) <= a and b;
    outputs(8532) <= not a;
    outputs(8533) <= b;
    outputs(8534) <= not (a xor b);
    outputs(8535) <= a xor b;
    outputs(8536) <= not (a and b);
    outputs(8537) <= not b;
    outputs(8538) <= a xor b;
    outputs(8539) <= not (a xor b);
    outputs(8540) <= not a;
    outputs(8541) <= not (a or b);
    outputs(8542) <= a;
    outputs(8543) <= b;
    outputs(8544) <= b;
    outputs(8545) <= a;
    outputs(8546) <= a;
    outputs(8547) <= not a or b;
    outputs(8548) <= b and not a;
    outputs(8549) <= not b;
    outputs(8550) <= a and b;
    outputs(8551) <= a;
    outputs(8552) <= b;
    outputs(8553) <= not (a xor b);
    outputs(8554) <= not (a xor b);
    outputs(8555) <= b;
    outputs(8556) <= b;
    outputs(8557) <= not a;
    outputs(8558) <= not a;
    outputs(8559) <= not (a and b);
    outputs(8560) <= b;
    outputs(8561) <= not (a xor b);
    outputs(8562) <= not (a xor b);
    outputs(8563) <= not b;
    outputs(8564) <= not a;
    outputs(8565) <= not (a xor b);
    outputs(8566) <= not a;
    outputs(8567) <= not a;
    outputs(8568) <= b;
    outputs(8569) <= not (a or b);
    outputs(8570) <= b;
    outputs(8571) <= not b;
    outputs(8572) <= a xor b;
    outputs(8573) <= not a;
    outputs(8574) <= a;
    outputs(8575) <= not b or a;
    outputs(8576) <= a xor b;
    outputs(8577) <= a;
    outputs(8578) <= a xor b;
    outputs(8579) <= a xor b;
    outputs(8580) <= not (a xor b);
    outputs(8581) <= not a;
    outputs(8582) <= not a or b;
    outputs(8583) <= a xor b;
    outputs(8584) <= not (a xor b);
    outputs(8585) <= a;
    outputs(8586) <= a;
    outputs(8587) <= not a;
    outputs(8588) <= a and not b;
    outputs(8589) <= not (a xor b);
    outputs(8590) <= a xor b;
    outputs(8591) <= a xor b;
    outputs(8592) <= a xor b;
    outputs(8593) <= a and not b;
    outputs(8594) <= b;
    outputs(8595) <= not a or b;
    outputs(8596) <= not a;
    outputs(8597) <= a xor b;
    outputs(8598) <= not b;
    outputs(8599) <= b;
    outputs(8600) <= a;
    outputs(8601) <= b;
    outputs(8602) <= a;
    outputs(8603) <= not (a xor b);
    outputs(8604) <= a xor b;
    outputs(8605) <= not a;
    outputs(8606) <= not (a xor b);
    outputs(8607) <= b and not a;
    outputs(8608) <= a xor b;
    outputs(8609) <= not a;
    outputs(8610) <= a xor b;
    outputs(8611) <= not a;
    outputs(8612) <= b;
    outputs(8613) <= a;
    outputs(8614) <= not a;
    outputs(8615) <= not b;
    outputs(8616) <= not b;
    outputs(8617) <= b;
    outputs(8618) <= a and not b;
    outputs(8619) <= b;
    outputs(8620) <= b;
    outputs(8621) <= not (a xor b);
    outputs(8622) <= a;
    outputs(8623) <= not a;
    outputs(8624) <= not b or a;
    outputs(8625) <= not a;
    outputs(8626) <= a;
    outputs(8627) <= not a or b;
    outputs(8628) <= not a;
    outputs(8629) <= a xor b;
    outputs(8630) <= not a;
    outputs(8631) <= not b;
    outputs(8632) <= not b;
    outputs(8633) <= a and b;
    outputs(8634) <= a and not b;
    outputs(8635) <= b;
    outputs(8636) <= not a;
    outputs(8637) <= a xor b;
    outputs(8638) <= not b;
    outputs(8639) <= a or b;
    outputs(8640) <= a;
    outputs(8641) <= not b;
    outputs(8642) <= not b;
    outputs(8643) <= not a;
    outputs(8644) <= a and not b;
    outputs(8645) <= a and not b;
    outputs(8646) <= not (a or b);
    outputs(8647) <= not a;
    outputs(8648) <= a xor b;
    outputs(8649) <= not b or a;
    outputs(8650) <= a or b;
    outputs(8651) <= a;
    outputs(8652) <= a;
    outputs(8653) <= not a;
    outputs(8654) <= b and not a;
    outputs(8655) <= not a;
    outputs(8656) <= a;
    outputs(8657) <= a and b;
    outputs(8658) <= a;
    outputs(8659) <= a xor b;
    outputs(8660) <= a;
    outputs(8661) <= not (a or b);
    outputs(8662) <= not (a and b);
    outputs(8663) <= not (a xor b);
    outputs(8664) <= not a;
    outputs(8665) <= a xor b;
    outputs(8666) <= a and not b;
    outputs(8667) <= a and b;
    outputs(8668) <= b;
    outputs(8669) <= b;
    outputs(8670) <= not b;
    outputs(8671) <= not a;
    outputs(8672) <= not b;
    outputs(8673) <= a and not b;
    outputs(8674) <= a and not b;
    outputs(8675) <= a xor b;
    outputs(8676) <= not (a or b);
    outputs(8677) <= not a or b;
    outputs(8678) <= a xor b;
    outputs(8679) <= not a or b;
    outputs(8680) <= not b;
    outputs(8681) <= not a;
    outputs(8682) <= b and not a;
    outputs(8683) <= a and b;
    outputs(8684) <= a xor b;
    outputs(8685) <= a xor b;
    outputs(8686) <= not (a xor b);
    outputs(8687) <= a and b;
    outputs(8688) <= a;
    outputs(8689) <= not a;
    outputs(8690) <= not (a or b);
    outputs(8691) <= a or b;
    outputs(8692) <= not b;
    outputs(8693) <= not b;
    outputs(8694) <= not b or a;
    outputs(8695) <= a xor b;
    outputs(8696) <= not (a xor b);
    outputs(8697) <= not (a xor b);
    outputs(8698) <= a and not b;
    outputs(8699) <= not b;
    outputs(8700) <= a xor b;
    outputs(8701) <= a xor b;
    outputs(8702) <= not (a xor b);
    outputs(8703) <= b;
    outputs(8704) <= not (a xor b);
    outputs(8705) <= a;
    outputs(8706) <= not (a xor b);
    outputs(8707) <= a;
    outputs(8708) <= not (a or b);
    outputs(8709) <= a and not b;
    outputs(8710) <= not a or b;
    outputs(8711) <= a and b;
    outputs(8712) <= a xor b;
    outputs(8713) <= a;
    outputs(8714) <= a;
    outputs(8715) <= not a;
    outputs(8716) <= a;
    outputs(8717) <= not (a xor b);
    outputs(8718) <= a xor b;
    outputs(8719) <= not a;
    outputs(8720) <= b;
    outputs(8721) <= not (a xor b);
    outputs(8722) <= not (a xor b);
    outputs(8723) <= a xor b;
    outputs(8724) <= a xor b;
    outputs(8725) <= not (a xor b);
    outputs(8726) <= not (a or b);
    outputs(8727) <= not a;
    outputs(8728) <= not a or b;
    outputs(8729) <= a xor b;
    outputs(8730) <= not a;
    outputs(8731) <= not (a xor b);
    outputs(8732) <= not a;
    outputs(8733) <= a;
    outputs(8734) <= a xor b;
    outputs(8735) <= not b;
    outputs(8736) <= not (a or b);
    outputs(8737) <= not b;
    outputs(8738) <= not (a xor b);
    outputs(8739) <= not (a xor b);
    outputs(8740) <= a xor b;
    outputs(8741) <= not a or b;
    outputs(8742) <= b;
    outputs(8743) <= not a;
    outputs(8744) <= a;
    outputs(8745) <= not (a or b);
    outputs(8746) <= not b;
    outputs(8747) <= a and b;
    outputs(8748) <= not b;
    outputs(8749) <= not a or b;
    outputs(8750) <= b;
    outputs(8751) <= not (a xor b);
    outputs(8752) <= b;
    outputs(8753) <= b;
    outputs(8754) <= b;
    outputs(8755) <= not b or a;
    outputs(8756) <= not (a xor b);
    outputs(8757) <= b;
    outputs(8758) <= not (a xor b);
    outputs(8759) <= a;
    outputs(8760) <= a xor b;
    outputs(8761) <= a xor b;
    outputs(8762) <= not (a xor b);
    outputs(8763) <= b;
    outputs(8764) <= b;
    outputs(8765) <= a xor b;
    outputs(8766) <= b;
    outputs(8767) <= not b;
    outputs(8768) <= b and not a;
    outputs(8769) <= b;
    outputs(8770) <= b and not a;
    outputs(8771) <= not b;
    outputs(8772) <= a;
    outputs(8773) <= b;
    outputs(8774) <= a xor b;
    outputs(8775) <= not b;
    outputs(8776) <= not (a xor b);
    outputs(8777) <= a and not b;
    outputs(8778) <= a;
    outputs(8779) <= a xor b;
    outputs(8780) <= a and not b;
    outputs(8781) <= b;
    outputs(8782) <= not b or a;
    outputs(8783) <= a and not b;
    outputs(8784) <= a xor b;
    outputs(8785) <= not b;
    outputs(8786) <= a xor b;
    outputs(8787) <= not a;
    outputs(8788) <= b;
    outputs(8789) <= b;
    outputs(8790) <= b;
    outputs(8791) <= a and not b;
    outputs(8792) <= not b or a;
    outputs(8793) <= not (a xor b);
    outputs(8794) <= b;
    outputs(8795) <= b and not a;
    outputs(8796) <= not a;
    outputs(8797) <= a;
    outputs(8798) <= b;
    outputs(8799) <= not a;
    outputs(8800) <= not a;
    outputs(8801) <= a;
    outputs(8802) <= a xor b;
    outputs(8803) <= a;
    outputs(8804) <= a xor b;
    outputs(8805) <= a xor b;
    outputs(8806) <= not b;
    outputs(8807) <= a and not b;
    outputs(8808) <= a;
    outputs(8809) <= a and not b;
    outputs(8810) <= b;
    outputs(8811) <= a xor b;
    outputs(8812) <= a;
    outputs(8813) <= b and not a;
    outputs(8814) <= a and b;
    outputs(8815) <= a and b;
    outputs(8816) <= not a or b;
    outputs(8817) <= not (a and b);
    outputs(8818) <= a;
    outputs(8819) <= not b;
    outputs(8820) <= a and not b;
    outputs(8821) <= not b;
    outputs(8822) <= a xor b;
    outputs(8823) <= b;
    outputs(8824) <= a xor b;
    outputs(8825) <= a;
    outputs(8826) <= a or b;
    outputs(8827) <= not a or b;
    outputs(8828) <= not (a or b);
    outputs(8829) <= b;
    outputs(8830) <= not (a or b);
    outputs(8831) <= b;
    outputs(8832) <= not b;
    outputs(8833) <= a xor b;
    outputs(8834) <= not a;
    outputs(8835) <= b;
    outputs(8836) <= not (a or b);
    outputs(8837) <= not b;
    outputs(8838) <= b and not a;
    outputs(8839) <= not (a xor b);
    outputs(8840) <= not a or b;
    outputs(8841) <= not (a xor b);
    outputs(8842) <= a xor b;
    outputs(8843) <= not (a xor b);
    outputs(8844) <= not a;
    outputs(8845) <= b;
    outputs(8846) <= a xor b;
    outputs(8847) <= a xor b;
    outputs(8848) <= a or b;
    outputs(8849) <= b;
    outputs(8850) <= not (a xor b);
    outputs(8851) <= a;
    outputs(8852) <= not b;
    outputs(8853) <= a;
    outputs(8854) <= not (a xor b);
    outputs(8855) <= b;
    outputs(8856) <= a xor b;
    outputs(8857) <= not (a xor b);
    outputs(8858) <= a and b;
    outputs(8859) <= a and not b;
    outputs(8860) <= b and not a;
    outputs(8861) <= not b or a;
    outputs(8862) <= a;
    outputs(8863) <= not a;
    outputs(8864) <= not a;
    outputs(8865) <= not b;
    outputs(8866) <= b;
    outputs(8867) <= not (a xor b);
    outputs(8868) <= not b;
    outputs(8869) <= b;
    outputs(8870) <= b and not a;
    outputs(8871) <= not (a xor b);
    outputs(8872) <= not b;
    outputs(8873) <= a xor b;
    outputs(8874) <= a and not b;
    outputs(8875) <= not (a xor b);
    outputs(8876) <= a xor b;
    outputs(8877) <= not (a xor b);
    outputs(8878) <= a xor b;
    outputs(8879) <= not a;
    outputs(8880) <= a;
    outputs(8881) <= a and b;
    outputs(8882) <= not (a xor b);
    outputs(8883) <= a;
    outputs(8884) <= a;
    outputs(8885) <= not a;
    outputs(8886) <= not (a and b);
    outputs(8887) <= a and b;
    outputs(8888) <= a xor b;
    outputs(8889) <= b;
    outputs(8890) <= a;
    outputs(8891) <= b and not a;
    outputs(8892) <= a;
    outputs(8893) <= not b;
    outputs(8894) <= a or b;
    outputs(8895) <= a xor b;
    outputs(8896) <= not a;
    outputs(8897) <= a and b;
    outputs(8898) <= b;
    outputs(8899) <= b;
    outputs(8900) <= not (a xor b);
    outputs(8901) <= a xor b;
    outputs(8902) <= b and not a;
    outputs(8903) <= b and not a;
    outputs(8904) <= not (a xor b);
    outputs(8905) <= not a;
    outputs(8906) <= not (a xor b);
    outputs(8907) <= a;
    outputs(8908) <= a;
    outputs(8909) <= '0';
    outputs(8910) <= not (a xor b);
    outputs(8911) <= not (a and b);
    outputs(8912) <= a;
    outputs(8913) <= not a or b;
    outputs(8914) <= not (a or b);
    outputs(8915) <= b;
    outputs(8916) <= a;
    outputs(8917) <= b;
    outputs(8918) <= a;
    outputs(8919) <= a xor b;
    outputs(8920) <= a xor b;
    outputs(8921) <= not (a or b);
    outputs(8922) <= not a;
    outputs(8923) <= not a;
    outputs(8924) <= a and b;
    outputs(8925) <= not b;
    outputs(8926) <= a;
    outputs(8927) <= b and not a;
    outputs(8928) <= not a;
    outputs(8929) <= a;
    outputs(8930) <= not a;
    outputs(8931) <= a or b;
    outputs(8932) <= a;
    outputs(8933) <= not a;
    outputs(8934) <= not a;
    outputs(8935) <= not b;
    outputs(8936) <= not (a xor b);
    outputs(8937) <= not a;
    outputs(8938) <= not a;
    outputs(8939) <= a;
    outputs(8940) <= a or b;
    outputs(8941) <= b;
    outputs(8942) <= a;
    outputs(8943) <= b and not a;
    outputs(8944) <= b;
    outputs(8945) <= not b;
    outputs(8946) <= a xor b;
    outputs(8947) <= b;
    outputs(8948) <= not b;
    outputs(8949) <= not (a and b);
    outputs(8950) <= not b;
    outputs(8951) <= a and b;
    outputs(8952) <= not (a xor b);
    outputs(8953) <= a;
    outputs(8954) <= not a;
    outputs(8955) <= a and b;
    outputs(8956) <= not a or b;
    outputs(8957) <= b;
    outputs(8958) <= not (a xor b);
    outputs(8959) <= not (a xor b);
    outputs(8960) <= not (a xor b);
    outputs(8961) <= a and not b;
    outputs(8962) <= not (a xor b);
    outputs(8963) <= not (a and b);
    outputs(8964) <= not (a xor b);
    outputs(8965) <= not (a or b);
    outputs(8966) <= not (a xor b);
    outputs(8967) <= not (a or b);
    outputs(8968) <= a or b;
    outputs(8969) <= not b;
    outputs(8970) <= not a;
    outputs(8971) <= not (a or b);
    outputs(8972) <= a;
    outputs(8973) <= b and not a;
    outputs(8974) <= b and not a;
    outputs(8975) <= not a;
    outputs(8976) <= a xor b;
    outputs(8977) <= not (a or b);
    outputs(8978) <= a;
    outputs(8979) <= a xor b;
    outputs(8980) <= b;
    outputs(8981) <= not (a xor b);
    outputs(8982) <= not b;
    outputs(8983) <= b;
    outputs(8984) <= b;
    outputs(8985) <= not b;
    outputs(8986) <= a and not b;
    outputs(8987) <= not (a xor b);
    outputs(8988) <= not (a xor b);
    outputs(8989) <= not b or a;
    outputs(8990) <= not a;
    outputs(8991) <= b;
    outputs(8992) <= b;
    outputs(8993) <= a xor b;
    outputs(8994) <= not (a xor b);
    outputs(8995) <= a xor b;
    outputs(8996) <= a and not b;
    outputs(8997) <= b;
    outputs(8998) <= not (a or b);
    outputs(8999) <= not (a xor b);
    outputs(9000) <= not (a xor b);
    outputs(9001) <= not (a xor b);
    outputs(9002) <= not (a xor b);
    outputs(9003) <= b;
    outputs(9004) <= a and b;
    outputs(9005) <= not (a and b);
    outputs(9006) <= a and not b;
    outputs(9007) <= not a;
    outputs(9008) <= a and b;
    outputs(9009) <= b;
    outputs(9010) <= not b;
    outputs(9011) <= a and b;
    outputs(9012) <= a xor b;
    outputs(9013) <= b;
    outputs(9014) <= not a;
    outputs(9015) <= a xor b;
    outputs(9016) <= not b;
    outputs(9017) <= a xor b;
    outputs(9018) <= a;
    outputs(9019) <= not b;
    outputs(9020) <= b;
    outputs(9021) <= a and b;
    outputs(9022) <= a xor b;
    outputs(9023) <= not (a xor b);
    outputs(9024) <= not (a xor b);
    outputs(9025) <= a;
    outputs(9026) <= not (a xor b);
    outputs(9027) <= not (a xor b);
    outputs(9028) <= a;
    outputs(9029) <= a or b;
    outputs(9030) <= b;
    outputs(9031) <= not a;
    outputs(9032) <= not b or a;
    outputs(9033) <= b;
    outputs(9034) <= a xor b;
    outputs(9035) <= a and b;
    outputs(9036) <= not (a and b);
    outputs(9037) <= not b or a;
    outputs(9038) <= a and b;
    outputs(9039) <= not a;
    outputs(9040) <= a and b;
    outputs(9041) <= not b;
    outputs(9042) <= not b or a;
    outputs(9043) <= b;
    outputs(9044) <= not b or a;
    outputs(9045) <= a;
    outputs(9046) <= not (a xor b);
    outputs(9047) <= '0';
    outputs(9048) <= not b or a;
    outputs(9049) <= not b;
    outputs(9050) <= a xor b;
    outputs(9051) <= a xor b;
    outputs(9052) <= not a;
    outputs(9053) <= not b;
    outputs(9054) <= not (a xor b);
    outputs(9055) <= a;
    outputs(9056) <= not a;
    outputs(9057) <= not (a xor b);
    outputs(9058) <= a xor b;
    outputs(9059) <= not (a xor b);
    outputs(9060) <= not (a xor b);
    outputs(9061) <= a;
    outputs(9062) <= not (a xor b);
    outputs(9063) <= not b;
    outputs(9064) <= a or b;
    outputs(9065) <= b;
    outputs(9066) <= not b;
    outputs(9067) <= not (a xor b);
    outputs(9068) <= not b;
    outputs(9069) <= not b;
    outputs(9070) <= a;
    outputs(9071) <= a and b;
    outputs(9072) <= a xor b;
    outputs(9073) <= not a;
    outputs(9074) <= not (a xor b);
    outputs(9075) <= a xor b;
    outputs(9076) <= not a or b;
    outputs(9077) <= a and b;
    outputs(9078) <= not a or b;
    outputs(9079) <= not (a xor b);
    outputs(9080) <= b;
    outputs(9081) <= not b;
    outputs(9082) <= not a or b;
    outputs(9083) <= b;
    outputs(9084) <= a and b;
    outputs(9085) <= a and b;
    outputs(9086) <= b;
    outputs(9087) <= a;
    outputs(9088) <= not (a or b);
    outputs(9089) <= a and b;
    outputs(9090) <= b;
    outputs(9091) <= not (a xor b);
    outputs(9092) <= a xor b;
    outputs(9093) <= not (a or b);
    outputs(9094) <= not (a xor b);
    outputs(9095) <= not b;
    outputs(9096) <= b;
    outputs(9097) <= a xor b;
    outputs(9098) <= not (a or b);
    outputs(9099) <= a and b;
    outputs(9100) <= not a;
    outputs(9101) <= a and b;
    outputs(9102) <= not b;
    outputs(9103) <= not a;
    outputs(9104) <= not b;
    outputs(9105) <= a xor b;
    outputs(9106) <= b;
    outputs(9107) <= not (a xor b);
    outputs(9108) <= not b;
    outputs(9109) <= not (a xor b);
    outputs(9110) <= not a;
    outputs(9111) <= a;
    outputs(9112) <= a xor b;
    outputs(9113) <= b;
    outputs(9114) <= not (a xor b);
    outputs(9115) <= b;
    outputs(9116) <= not (a or b);
    outputs(9117) <= a xor b;
    outputs(9118) <= not (a xor b);
    outputs(9119) <= not (a xor b);
    outputs(9120) <= not a;
    outputs(9121) <= not (a or b);
    outputs(9122) <= not b;
    outputs(9123) <= a;
    outputs(9124) <= a xor b;
    outputs(9125) <= not b;
    outputs(9126) <= not a;
    outputs(9127) <= not (a xor b);
    outputs(9128) <= not b;
    outputs(9129) <= a;
    outputs(9130) <= not a;
    outputs(9131) <= a xor b;
    outputs(9132) <= not (a xor b);
    outputs(9133) <= not (a xor b);
    outputs(9134) <= not (a xor b);
    outputs(9135) <= not b;
    outputs(9136) <= a;
    outputs(9137) <= not (a xor b);
    outputs(9138) <= a xor b;
    outputs(9139) <= not (a or b);
    outputs(9140) <= a xor b;
    outputs(9141) <= b and not a;
    outputs(9142) <= a xor b;
    outputs(9143) <= b;
    outputs(9144) <= a;
    outputs(9145) <= not a;
    outputs(9146) <= not b;
    outputs(9147) <= a;
    outputs(9148) <= a and not b;
    outputs(9149) <= not (a xor b);
    outputs(9150) <= b;
    outputs(9151) <= b;
    outputs(9152) <= a xor b;
    outputs(9153) <= a xor b;
    outputs(9154) <= not a;
    outputs(9155) <= a xor b;
    outputs(9156) <= not b or a;
    outputs(9157) <= not a;
    outputs(9158) <= not (a xor b);
    outputs(9159) <= not a;
    outputs(9160) <= not b or a;
    outputs(9161) <= not (a xor b);
    outputs(9162) <= a xor b;
    outputs(9163) <= b;
    outputs(9164) <= not (a or b);
    outputs(9165) <= not b;
    outputs(9166) <= not b;
    outputs(9167) <= not (a xor b);
    outputs(9168) <= a xor b;
    outputs(9169) <= b;
    outputs(9170) <= not a;
    outputs(9171) <= b;
    outputs(9172) <= b and not a;
    outputs(9173) <= a;
    outputs(9174) <= not b;
    outputs(9175) <= b;
    outputs(9176) <= not b;
    outputs(9177) <= a xor b;
    outputs(9178) <= a and not b;
    outputs(9179) <= a xor b;
    outputs(9180) <= not b or a;
    outputs(9181) <= a xor b;
    outputs(9182) <= not b;
    outputs(9183) <= a and not b;
    outputs(9184) <= not (a xor b);
    outputs(9185) <= not b;
    outputs(9186) <= a;
    outputs(9187) <= b and not a;
    outputs(9188) <= b;
    outputs(9189) <= a;
    outputs(9190) <= not a;
    outputs(9191) <= not b;
    outputs(9192) <= b;
    outputs(9193) <= a;
    outputs(9194) <= a;
    outputs(9195) <= b;
    outputs(9196) <= a;
    outputs(9197) <= b;
    outputs(9198) <= not (a and b);
    outputs(9199) <= not (a or b);
    outputs(9200) <= b and not a;
    outputs(9201) <= a xor b;
    outputs(9202) <= a xor b;
    outputs(9203) <= not (a xor b);
    outputs(9204) <= not (a or b);
    outputs(9205) <= not b;
    outputs(9206) <= a xor b;
    outputs(9207) <= not (a xor b);
    outputs(9208) <= not (a xor b);
    outputs(9209) <= a xor b;
    outputs(9210) <= not (a xor b);
    outputs(9211) <= a and b;
    outputs(9212) <= not b;
    outputs(9213) <= not a;
    outputs(9214) <= a;
    outputs(9215) <= a;
    outputs(9216) <= a and b;
    outputs(9217) <= a xor b;
    outputs(9218) <= not a;
    outputs(9219) <= not a;
    outputs(9220) <= a or b;
    outputs(9221) <= a and b;
    outputs(9222) <= a xor b;
    outputs(9223) <= not (a or b);
    outputs(9224) <= not a;
    outputs(9225) <= a and not b;
    outputs(9226) <= not (a xor b);
    outputs(9227) <= a or b;
    outputs(9228) <= not a;
    outputs(9229) <= b and not a;
    outputs(9230) <= a and not b;
    outputs(9231) <= not (a or b);
    outputs(9232) <= a;
    outputs(9233) <= not a;
    outputs(9234) <= not b;
    outputs(9235) <= a and not b;
    outputs(9236) <= b;
    outputs(9237) <= not (a xor b);
    outputs(9238) <= a;
    outputs(9239) <= a xor b;
    outputs(9240) <= a and b;
    outputs(9241) <= a and not b;
    outputs(9242) <= not b;
    outputs(9243) <= a;
    outputs(9244) <= not b;
    outputs(9245) <= b;
    outputs(9246) <= a;
    outputs(9247) <= not a;
    outputs(9248) <= not b;
    outputs(9249) <= b;
    outputs(9250) <= a;
    outputs(9251) <= a;
    outputs(9252) <= not a;
    outputs(9253) <= not a;
    outputs(9254) <= a xor b;
    outputs(9255) <= a;
    outputs(9256) <= a xor b;
    outputs(9257) <= a;
    outputs(9258) <= not (a xor b);
    outputs(9259) <= a;
    outputs(9260) <= a xor b;
    outputs(9261) <= a;
    outputs(9262) <= not b;
    outputs(9263) <= not (a or b);
    outputs(9264) <= a xor b;
    outputs(9265) <= not a;
    outputs(9266) <= not (a or b);
    outputs(9267) <= a;
    outputs(9268) <= not b;
    outputs(9269) <= b;
    outputs(9270) <= not (a and b);
    outputs(9271) <= b and not a;
    outputs(9272) <= b;
    outputs(9273) <= not a;
    outputs(9274) <= b and not a;
    outputs(9275) <= b;
    outputs(9276) <= not (a xor b);
    outputs(9277) <= a or b;
    outputs(9278) <= a xor b;
    outputs(9279) <= a;
    outputs(9280) <= not (a xor b);
    outputs(9281) <= b and not a;
    outputs(9282) <= a xor b;
    outputs(9283) <= a;
    outputs(9284) <= a and not b;
    outputs(9285) <= not (a xor b);
    outputs(9286) <= a;
    outputs(9287) <= a xor b;
    outputs(9288) <= not b;
    outputs(9289) <= a;
    outputs(9290) <= b;
    outputs(9291) <= a xor b;
    outputs(9292) <= not (a xor b);
    outputs(9293) <= a xor b;
    outputs(9294) <= a and b;
    outputs(9295) <= not b;
    outputs(9296) <= not b;
    outputs(9297) <= b;
    outputs(9298) <= b;
    outputs(9299) <= not a;
    outputs(9300) <= not (a xor b);
    outputs(9301) <= a xor b;
    outputs(9302) <= not (a xor b);
    outputs(9303) <= not b;
    outputs(9304) <= not (a xor b);
    outputs(9305) <= not (a xor b);
    outputs(9306) <= a and b;
    outputs(9307) <= a and not b;
    outputs(9308) <= not a;
    outputs(9309) <= not b;
    outputs(9310) <= a;
    outputs(9311) <= not (a xor b);
    outputs(9312) <= not (a or b);
    outputs(9313) <= a xor b;
    outputs(9314) <= b;
    outputs(9315) <= not b;
    outputs(9316) <= not (a xor b);
    outputs(9317) <= a;
    outputs(9318) <= not (a or b);
    outputs(9319) <= not (a xor b);
    outputs(9320) <= b;
    outputs(9321) <= b;
    outputs(9322) <= a;
    outputs(9323) <= a and not b;
    outputs(9324) <= a xor b;
    outputs(9325) <= not b;
    outputs(9326) <= not b or a;
    outputs(9327) <= a xor b;
    outputs(9328) <= not a;
    outputs(9329) <= not b;
    outputs(9330) <= not (a xor b);
    outputs(9331) <= not (a xor b);
    outputs(9332) <= a and not b;
    outputs(9333) <= not b;
    outputs(9334) <= a xor b;
    outputs(9335) <= not (a and b);
    outputs(9336) <= not b;
    outputs(9337) <= a;
    outputs(9338) <= not (a or b);
    outputs(9339) <= not b;
    outputs(9340) <= a;
    outputs(9341) <= a xor b;
    outputs(9342) <= not b or a;
    outputs(9343) <= a xor b;
    outputs(9344) <= a xor b;
    outputs(9345) <= a;
    outputs(9346) <= not (a or b);
    outputs(9347) <= a and not b;
    outputs(9348) <= not a;
    outputs(9349) <= a xor b;
    outputs(9350) <= not a or b;
    outputs(9351) <= a and not b;
    outputs(9352) <= not b;
    outputs(9353) <= not (a xor b);
    outputs(9354) <= b and not a;
    outputs(9355) <= b and not a;
    outputs(9356) <= b and not a;
    outputs(9357) <= a and not b;
    outputs(9358) <= not (a or b);
    outputs(9359) <= b and not a;
    outputs(9360) <= a;
    outputs(9361) <= not (a xor b);
    outputs(9362) <= not (a xor b);
    outputs(9363) <= b and not a;
    outputs(9364) <= a;
    outputs(9365) <= not (a xor b);
    outputs(9366) <= b;
    outputs(9367) <= not b;
    outputs(9368) <= a xor b;
    outputs(9369) <= not b;
    outputs(9370) <= not (a xor b);
    outputs(9371) <= not a;
    outputs(9372) <= not (a xor b);
    outputs(9373) <= not b;
    outputs(9374) <= not (a xor b);
    outputs(9375) <= not b;
    outputs(9376) <= not b;
    outputs(9377) <= a xor b;
    outputs(9378) <= not b;
    outputs(9379) <= not a;
    outputs(9380) <= not (a xor b);
    outputs(9381) <= a and b;
    outputs(9382) <= not (a xor b);
    outputs(9383) <= not a;
    outputs(9384) <= a and b;
    outputs(9385) <= not b;
    outputs(9386) <= a xor b;
    outputs(9387) <= not (a or b);
    outputs(9388) <= a and not b;
    outputs(9389) <= a or b;
    outputs(9390) <= a and not b;
    outputs(9391) <= a xor b;
    outputs(9392) <= b;
    outputs(9393) <= not (a xor b);
    outputs(9394) <= b;
    outputs(9395) <= a;
    outputs(9396) <= a xor b;
    outputs(9397) <= not (a xor b);
    outputs(9398) <= b;
    outputs(9399) <= not b;
    outputs(9400) <= b and not a;
    outputs(9401) <= b;
    outputs(9402) <= b and not a;
    outputs(9403) <= not b;
    outputs(9404) <= a and not b;
    outputs(9405) <= not (a xor b);
    outputs(9406) <= not a;
    outputs(9407) <= a;
    outputs(9408) <= a;
    outputs(9409) <= a and b;
    outputs(9410) <= b;
    outputs(9411) <= not (a xor b);
    outputs(9412) <= a and not b;
    outputs(9413) <= not a;
    outputs(9414) <= not (a xor b);
    outputs(9415) <= b;
    outputs(9416) <= a and not b;
    outputs(9417) <= not (a xor b);
    outputs(9418) <= a xor b;
    outputs(9419) <= not (a xor b);
    outputs(9420) <= b and not a;
    outputs(9421) <= not b;
    outputs(9422) <= not b;
    outputs(9423) <= not b;
    outputs(9424) <= not a or b;
    outputs(9425) <= not (a or b);
    outputs(9426) <= not a;
    outputs(9427) <= not (a xor b);
    outputs(9428) <= not b or a;
    outputs(9429) <= a and not b;
    outputs(9430) <= b;
    outputs(9431) <= not (a xor b);
    outputs(9432) <= b;
    outputs(9433) <= a xor b;
    outputs(9434) <= a xor b;
    outputs(9435) <= a xor b;
    outputs(9436) <= a;
    outputs(9437) <= b;
    outputs(9438) <= b;
    outputs(9439) <= not (a xor b);
    outputs(9440) <= not a;
    outputs(9441) <= b and not a;
    outputs(9442) <= a xor b;
    outputs(9443) <= not (a xor b);
    outputs(9444) <= a or b;
    outputs(9445) <= b;
    outputs(9446) <= b;
    outputs(9447) <= not b;
    outputs(9448) <= a xor b;
    outputs(9449) <= not b;
    outputs(9450) <= a and b;
    outputs(9451) <= not b or a;
    outputs(9452) <= a xor b;
    outputs(9453) <= a or b;
    outputs(9454) <= not (a xor b);
    outputs(9455) <= not b;
    outputs(9456) <= not (a xor b);
    outputs(9457) <= not a;
    outputs(9458) <= not (a or b);
    outputs(9459) <= not b or a;
    outputs(9460) <= a and b;
    outputs(9461) <= b;
    outputs(9462) <= b;
    outputs(9463) <= not (a xor b);
    outputs(9464) <= not (a xor b);
    outputs(9465) <= not b;
    outputs(9466) <= b and not a;
    outputs(9467) <= not a;
    outputs(9468) <= a xor b;
    outputs(9469) <= a and not b;
    outputs(9470) <= a xor b;
    outputs(9471) <= a xor b;
    outputs(9472) <= not (a xor b);
    outputs(9473) <= not b;
    outputs(9474) <= b;
    outputs(9475) <= a and b;
    outputs(9476) <= not (a xor b);
    outputs(9477) <= not (a xor b);
    outputs(9478) <= not b;
    outputs(9479) <= a and b;
    outputs(9480) <= not (a xor b);
    outputs(9481) <= not a;
    outputs(9482) <= not a;
    outputs(9483) <= not b or a;
    outputs(9484) <= a and not b;
    outputs(9485) <= not b or a;
    outputs(9486) <= not (a xor b);
    outputs(9487) <= a or b;
    outputs(9488) <= b and not a;
    outputs(9489) <= a xor b;
    outputs(9490) <= not (a xor b);
    outputs(9491) <= a xor b;
    outputs(9492) <= not b or a;
    outputs(9493) <= b;
    outputs(9494) <= a;
    outputs(9495) <= a xor b;
    outputs(9496) <= a;
    outputs(9497) <= a xor b;
    outputs(9498) <= a and not b;
    outputs(9499) <= a and b;
    outputs(9500) <= a;
    outputs(9501) <= a;
    outputs(9502) <= a and not b;
    outputs(9503) <= not (a or b);
    outputs(9504) <= b;
    outputs(9505) <= not a;
    outputs(9506) <= a;
    outputs(9507) <= a;
    outputs(9508) <= not b or a;
    outputs(9509) <= not b;
    outputs(9510) <= not b;
    outputs(9511) <= a xor b;
    outputs(9512) <= a and b;
    outputs(9513) <= not (a xor b);
    outputs(9514) <= a and b;
    outputs(9515) <= not (a or b);
    outputs(9516) <= a xor b;
    outputs(9517) <= a xor b;
    outputs(9518) <= b and not a;
    outputs(9519) <= a xor b;
    outputs(9520) <= a xor b;
    outputs(9521) <= not a;
    outputs(9522) <= a xor b;
    outputs(9523) <= not (a xor b);
    outputs(9524) <= not b;
    outputs(9525) <= a;
    outputs(9526) <= not a or b;
    outputs(9527) <= b and not a;
    outputs(9528) <= b;
    outputs(9529) <= not (a or b);
    outputs(9530) <= a or b;
    outputs(9531) <= a xor b;
    outputs(9532) <= a xor b;
    outputs(9533) <= a;
    outputs(9534) <= not (a or b);
    outputs(9535) <= a;
    outputs(9536) <= a xor b;
    outputs(9537) <= not b;
    outputs(9538) <= b and not a;
    outputs(9539) <= not b;
    outputs(9540) <= a and b;
    outputs(9541) <= a xor b;
    outputs(9542) <= not a;
    outputs(9543) <= a xor b;
    outputs(9544) <= not (a xor b);
    outputs(9545) <= b;
    outputs(9546) <= a xor b;
    outputs(9547) <= a;
    outputs(9548) <= not (a xor b);
    outputs(9549) <= b and not a;
    outputs(9550) <= b and not a;
    outputs(9551) <= not a;
    outputs(9552) <= not b;
    outputs(9553) <= a xor b;
    outputs(9554) <= a xor b;
    outputs(9555) <= a;
    outputs(9556) <= a and b;
    outputs(9557) <= not (a xor b);
    outputs(9558) <= b;
    outputs(9559) <= not (a xor b);
    outputs(9560) <= not a;
    outputs(9561) <= not a;
    outputs(9562) <= not b;
    outputs(9563) <= not b;
    outputs(9564) <= a xor b;
    outputs(9565) <= not (a xor b);
    outputs(9566) <= not (a xor b);
    outputs(9567) <= a;
    outputs(9568) <= a;
    outputs(9569) <= not (a or b);
    outputs(9570) <= a xor b;
    outputs(9571) <= not (a xor b);
    outputs(9572) <= a xor b;
    outputs(9573) <= not (a xor b);
    outputs(9574) <= not a;
    outputs(9575) <= not (a xor b);
    outputs(9576) <= a xor b;
    outputs(9577) <= a;
    outputs(9578) <= a and not b;
    outputs(9579) <= a;
    outputs(9580) <= not (a xor b);
    outputs(9581) <= not (a xor b);
    outputs(9582) <= not b;
    outputs(9583) <= not (a or b);
    outputs(9584) <= not a;
    outputs(9585) <= a or b;
    outputs(9586) <= a and b;
    outputs(9587) <= a xor b;
    outputs(9588) <= a and not b;
    outputs(9589) <= not b;
    outputs(9590) <= a xor b;
    outputs(9591) <= not b;
    outputs(9592) <= a;
    outputs(9593) <= not (a and b);
    outputs(9594) <= b;
    outputs(9595) <= not b;
    outputs(9596) <= a xor b;
    outputs(9597) <= not b or a;
    outputs(9598) <= not (a xor b);
    outputs(9599) <= not (a or b);
    outputs(9600) <= b;
    outputs(9601) <= a;
    outputs(9602) <= b;
    outputs(9603) <= not a;
    outputs(9604) <= not a;
    outputs(9605) <= not a or b;
    outputs(9606) <= not (a xor b);
    outputs(9607) <= a and not b;
    outputs(9608) <= not a;
    outputs(9609) <= a xor b;
    outputs(9610) <= b and not a;
    outputs(9611) <= a xor b;
    outputs(9612) <= a and b;
    outputs(9613) <= a or b;
    outputs(9614) <= b and not a;
    outputs(9615) <= not b;
    outputs(9616) <= b;
    outputs(9617) <= b;
    outputs(9618) <= a xor b;
    outputs(9619) <= a xor b;
    outputs(9620) <= b;
    outputs(9621) <= a;
    outputs(9622) <= a xor b;
    outputs(9623) <= a;
    outputs(9624) <= not (a and b);
    outputs(9625) <= b;
    outputs(9626) <= a;
    outputs(9627) <= b;
    outputs(9628) <= not a;
    outputs(9629) <= not (a xor b);
    outputs(9630) <= a;
    outputs(9631) <= not (a xor b);
    outputs(9632) <= not b;
    outputs(9633) <= a xor b;
    outputs(9634) <= a xor b;
    outputs(9635) <= b;
    outputs(9636) <= b;
    outputs(9637) <= a xor b;
    outputs(9638) <= not a;
    outputs(9639) <= b;
    outputs(9640) <= b;
    outputs(9641) <= not (a xor b);
    outputs(9642) <= a xor b;
    outputs(9643) <= a and not b;
    outputs(9644) <= not a or b;
    outputs(9645) <= not b;
    outputs(9646) <= b;
    outputs(9647) <= not (a xor b);
    outputs(9648) <= not b or a;
    outputs(9649) <= not (a or b);
    outputs(9650) <= not (a and b);
    outputs(9651) <= not b;
    outputs(9652) <= b;
    outputs(9653) <= b;
    outputs(9654) <= a and b;
    outputs(9655) <= b;
    outputs(9656) <= not a;
    outputs(9657) <= not b;
    outputs(9658) <= a xor b;
    outputs(9659) <= a or b;
    outputs(9660) <= not (a xor b);
    outputs(9661) <= a xor b;
    outputs(9662) <= a xor b;
    outputs(9663) <= a xor b;
    outputs(9664) <= b;
    outputs(9665) <= not a;
    outputs(9666) <= not (a or b);
    outputs(9667) <= not a;
    outputs(9668) <= not (a xor b);
    outputs(9669) <= b;
    outputs(9670) <= a xor b;
    outputs(9671) <= not (a xor b);
    outputs(9672) <= not (a xor b);
    outputs(9673) <= b;
    outputs(9674) <= not (a or b);
    outputs(9675) <= a;
    outputs(9676) <= not b;
    outputs(9677) <= not a or b;
    outputs(9678) <= a xor b;
    outputs(9679) <= not a;
    outputs(9680) <= not (a xor b);
    outputs(9681) <= not (a xor b);
    outputs(9682) <= a xor b;
    outputs(9683) <= not a;
    outputs(9684) <= not b;
    outputs(9685) <= a;
    outputs(9686) <= b;
    outputs(9687) <= a xor b;
    outputs(9688) <= a;
    outputs(9689) <= a xor b;
    outputs(9690) <= not (a xor b);
    outputs(9691) <= a;
    outputs(9692) <= not b;
    outputs(9693) <= b;
    outputs(9694) <= a;
    outputs(9695) <= a and b;
    outputs(9696) <= a xor b;
    outputs(9697) <= b;
    outputs(9698) <= a xor b;
    outputs(9699) <= a;
    outputs(9700) <= not (a xor b);
    outputs(9701) <= not b;
    outputs(9702) <= a and not b;
    outputs(9703) <= b and not a;
    outputs(9704) <= not (a xor b);
    outputs(9705) <= not (a xor b);
    outputs(9706) <= b and not a;
    outputs(9707) <= a xor b;
    outputs(9708) <= not (a xor b);
    outputs(9709) <= a xor b;
    outputs(9710) <= a and b;
    outputs(9711) <= not a or b;
    outputs(9712) <= a;
    outputs(9713) <= not b;
    outputs(9714) <= a;
    outputs(9715) <= not (a and b);
    outputs(9716) <= not b;
    outputs(9717) <= a;
    outputs(9718) <= a and b;
    outputs(9719) <= not (a and b);
    outputs(9720) <= not (a xor b);
    outputs(9721) <= a;
    outputs(9722) <= a xor b;
    outputs(9723) <= a;
    outputs(9724) <= b;
    outputs(9725) <= a;
    outputs(9726) <= not (a xor b);
    outputs(9727) <= not (a xor b);
    outputs(9728) <= b and not a;
    outputs(9729) <= not (a xor b);
    outputs(9730) <= b and not a;
    outputs(9731) <= not b;
    outputs(9732) <= a and b;
    outputs(9733) <= a xor b;
    outputs(9734) <= not (a xor b);
    outputs(9735) <= not (a and b);
    outputs(9736) <= a;
    outputs(9737) <= a and not b;
    outputs(9738) <= a xor b;
    outputs(9739) <= not b;
    outputs(9740) <= not (a or b);
    outputs(9741) <= a xor b;
    outputs(9742) <= b;
    outputs(9743) <= b;
    outputs(9744) <= b;
    outputs(9745) <= not (a xor b);
    outputs(9746) <= a and not b;
    outputs(9747) <= a;
    outputs(9748) <= not (a xor b);
    outputs(9749) <= a xor b;
    outputs(9750) <= not (a or b);
    outputs(9751) <= a xor b;
    outputs(9752) <= b and not a;
    outputs(9753) <= not a;
    outputs(9754) <= a or b;
    outputs(9755) <= a and not b;
    outputs(9756) <= b and not a;
    outputs(9757) <= not a;
    outputs(9758) <= a xor b;
    outputs(9759) <= a xor b;
    outputs(9760) <= a;
    outputs(9761) <= not (a or b);
    outputs(9762) <= b and not a;
    outputs(9763) <= b and not a;
    outputs(9764) <= b and not a;
    outputs(9765) <= not a;
    outputs(9766) <= b;
    outputs(9767) <= a xor b;
    outputs(9768) <= not (a xor b);
    outputs(9769) <= not (a or b);
    outputs(9770) <= not a;
    outputs(9771) <= not (a xor b);
    outputs(9772) <= a and not b;
    outputs(9773) <= not (a or b);
    outputs(9774) <= a and b;
    outputs(9775) <= not a;
    outputs(9776) <= a;
    outputs(9777) <= not (a xor b);
    outputs(9778) <= a and b;
    outputs(9779) <= a xor b;
    outputs(9780) <= not b;
    outputs(9781) <= a;
    outputs(9782) <= a and b;
    outputs(9783) <= not a;
    outputs(9784) <= b;
    outputs(9785) <= b and not a;
    outputs(9786) <= a and b;
    outputs(9787) <= a xor b;
    outputs(9788) <= a and not b;
    outputs(9789) <= not (a xor b);
    outputs(9790) <= not b;
    outputs(9791) <= not a;
    outputs(9792) <= not b;
    outputs(9793) <= a xor b;
    outputs(9794) <= a and b;
    outputs(9795) <= not (a xor b);
    outputs(9796) <= b and not a;
    outputs(9797) <= a and b;
    outputs(9798) <= a and b;
    outputs(9799) <= not a;
    outputs(9800) <= not a or b;
    outputs(9801) <= a and not b;
    outputs(9802) <= b and not a;
    outputs(9803) <= b;
    outputs(9804) <= not a;
    outputs(9805) <= a;
    outputs(9806) <= b;
    outputs(9807) <= a;
    outputs(9808) <= not (a or b);
    outputs(9809) <= not a;
    outputs(9810) <= not a;
    outputs(9811) <= a;
    outputs(9812) <= not a or b;
    outputs(9813) <= not a;
    outputs(9814) <= b;
    outputs(9815) <= a;
    outputs(9816) <= not a;
    outputs(9817) <= not b;
    outputs(9818) <= a;
    outputs(9819) <= not a or b;
    outputs(9820) <= not b;
    outputs(9821) <= not (a xor b);
    outputs(9822) <= a;
    outputs(9823) <= a;
    outputs(9824) <= not a;
    outputs(9825) <= b;
    outputs(9826) <= a;
    outputs(9827) <= not a or b;
    outputs(9828) <= a and not b;
    outputs(9829) <= b;
    outputs(9830) <= a xor b;
    outputs(9831) <= not (a xor b);
    outputs(9832) <= not b;
    outputs(9833) <= not b;
    outputs(9834) <= b;
    outputs(9835) <= a xor b;
    outputs(9836) <= a and not b;
    outputs(9837) <= not b;
    outputs(9838) <= a and not b;
    outputs(9839) <= not (a or b);
    outputs(9840) <= not (a xor b);
    outputs(9841) <= a;
    outputs(9842) <= a xor b;
    outputs(9843) <= not a;
    outputs(9844) <= a;
    outputs(9845) <= not (a xor b);
    outputs(9846) <= not a;
    outputs(9847) <= not b;
    outputs(9848) <= a and b;
    outputs(9849) <= not b;
    outputs(9850) <= a xor b;
    outputs(9851) <= a;
    outputs(9852) <= not (a xor b);
    outputs(9853) <= a;
    outputs(9854) <= a and b;
    outputs(9855) <= not (a or b);
    outputs(9856) <= a and not b;
    outputs(9857) <= not a;
    outputs(9858) <= b;
    outputs(9859) <= a xor b;
    outputs(9860) <= a xor b;
    outputs(9861) <= a and not b;
    outputs(9862) <= not (a xor b);
    outputs(9863) <= b;
    outputs(9864) <= a;
    outputs(9865) <= b;
    outputs(9866) <= not (a xor b);
    outputs(9867) <= not a;
    outputs(9868) <= b;
    outputs(9869) <= a xor b;
    outputs(9870) <= not b;
    outputs(9871) <= not a;
    outputs(9872) <= not b;
    outputs(9873) <= not a;
    outputs(9874) <= not (a and b);
    outputs(9875) <= not a or b;
    outputs(9876) <= not a;
    outputs(9877) <= a;
    outputs(9878) <= a;
    outputs(9879) <= b and not a;
    outputs(9880) <= a;
    outputs(9881) <= not a;
    outputs(9882) <= b and not a;
    outputs(9883) <= not (a xor b);
    outputs(9884) <= not b;
    outputs(9885) <= a and not b;
    outputs(9886) <= b;
    outputs(9887) <= a and not b;
    outputs(9888) <= not (a xor b);
    outputs(9889) <= b;
    outputs(9890) <= not b;
    outputs(9891) <= not b;
    outputs(9892) <= a and not b;
    outputs(9893) <= b;
    outputs(9894) <= a xor b;
    outputs(9895) <= not b;
    outputs(9896) <= not a or b;
    outputs(9897) <= not b;
    outputs(9898) <= a;
    outputs(9899) <= b;
    outputs(9900) <= not a or b;
    outputs(9901) <= not (a xor b);
    outputs(9902) <= not (a xor b);
    outputs(9903) <= not b;
    outputs(9904) <= not b;
    outputs(9905) <= not (a and b);
    outputs(9906) <= b;
    outputs(9907) <= a;
    outputs(9908) <= a xor b;
    outputs(9909) <= not (a xor b);
    outputs(9910) <= b;
    outputs(9911) <= not (a or b);
    outputs(9912) <= a xor b;
    outputs(9913) <= not b;
    outputs(9914) <= a xor b;
    outputs(9915) <= a;
    outputs(9916) <= b and not a;
    outputs(9917) <= not b;
    outputs(9918) <= a xor b;
    outputs(9919) <= a;
    outputs(9920) <= a;
    outputs(9921) <= not (a xor b);
    outputs(9922) <= not (a xor b);
    outputs(9923) <= a and not b;
    outputs(9924) <= not b;
    outputs(9925) <= not (a or b);
    outputs(9926) <= not b;
    outputs(9927) <= a and not b;
    outputs(9928) <= b;
    outputs(9929) <= b and not a;
    outputs(9930) <= not b;
    outputs(9931) <= b and not a;
    outputs(9932) <= a and b;
    outputs(9933) <= a xor b;
    outputs(9934) <= not b;
    outputs(9935) <= not a;
    outputs(9936) <= b and not a;
    outputs(9937) <= a xor b;
    outputs(9938) <= not b;
    outputs(9939) <= b;
    outputs(9940) <= not a;
    outputs(9941) <= not (a xor b);
    outputs(9942) <= not (a xor b);
    outputs(9943) <= a xor b;
    outputs(9944) <= a xor b;
    outputs(9945) <= b;
    outputs(9946) <= not (a or b);
    outputs(9947) <= a and b;
    outputs(9948) <= not (a xor b);
    outputs(9949) <= not b;
    outputs(9950) <= a and not b;
    outputs(9951) <= not (a or b);
    outputs(9952) <= not a;
    outputs(9953) <= a xor b;
    outputs(9954) <= a;
    outputs(9955) <= a or b;
    outputs(9956) <= a;
    outputs(9957) <= not b;
    outputs(9958) <= b;
    outputs(9959) <= not (a xor b);
    outputs(9960) <= not a;
    outputs(9961) <= a xor b;
    outputs(9962) <= a xor b;
    outputs(9963) <= not a;
    outputs(9964) <= a or b;
    outputs(9965) <= not (a and b);
    outputs(9966) <= not (a xor b);
    outputs(9967) <= b;
    outputs(9968) <= not (a and b);
    outputs(9969) <= not a;
    outputs(9970) <= a xor b;
    outputs(9971) <= a;
    outputs(9972) <= not a or b;
    outputs(9973) <= not (a or b);
    outputs(9974) <= a and not b;
    outputs(9975) <= a and not b;
    outputs(9976) <= not (a xor b);
    outputs(9977) <= a and not b;
    outputs(9978) <= a xor b;
    outputs(9979) <= a xor b;
    outputs(9980) <= a and not b;
    outputs(9981) <= not (a xor b);
    outputs(9982) <= a xor b;
    outputs(9983) <= a xor b;
    outputs(9984) <= not b;
    outputs(9985) <= a and not b;
    outputs(9986) <= a;
    outputs(9987) <= b and not a;
    outputs(9988) <= not a;
    outputs(9989) <= not (a xor b);
    outputs(9990) <= not b;
    outputs(9991) <= b;
    outputs(9992) <= a;
    outputs(9993) <= a;
    outputs(9994) <= a xor b;
    outputs(9995) <= not b;
    outputs(9996) <= not (a xor b);
    outputs(9997) <= not (a or b);
    outputs(9998) <= a and not b;
    outputs(9999) <= not b;
    outputs(10000) <= not (a xor b);
    outputs(10001) <= not (a or b);
    outputs(10002) <= not b;
    outputs(10003) <= a;
    outputs(10004) <= a and not b;
    outputs(10005) <= a xor b;
    outputs(10006) <= a;
    outputs(10007) <= not (a xor b);
    outputs(10008) <= not a;
    outputs(10009) <= not a;
    outputs(10010) <= not (a xor b);
    outputs(10011) <= not b;
    outputs(10012) <= not (a xor b);
    outputs(10013) <= a xor b;
    outputs(10014) <= a;
    outputs(10015) <= not b;
    outputs(10016) <= a and b;
    outputs(10017) <= a xor b;
    outputs(10018) <= a and not b;
    outputs(10019) <= a and not b;
    outputs(10020) <= not b;
    outputs(10021) <= not a;
    outputs(10022) <= not (a xor b);
    outputs(10023) <= not (a xor b);
    outputs(10024) <= not (a or b);
    outputs(10025) <= a;
    outputs(10026) <= not b;
    outputs(10027) <= a;
    outputs(10028) <= not a;
    outputs(10029) <= b and not a;
    outputs(10030) <= not b;
    outputs(10031) <= not a;
    outputs(10032) <= a and b;
    outputs(10033) <= a and b;
    outputs(10034) <= not (a xor b);
    outputs(10035) <= a xor b;
    outputs(10036) <= a xor b;
    outputs(10037) <= not a;
    outputs(10038) <= b;
    outputs(10039) <= a;
    outputs(10040) <= a xor b;
    outputs(10041) <= not b or a;
    outputs(10042) <= not (a xor b);
    outputs(10043) <= not a;
    outputs(10044) <= a;
    outputs(10045) <= not (a xor b);
    outputs(10046) <= not b;
    outputs(10047) <= not a or b;
    outputs(10048) <= b;
    outputs(10049) <= a;
    outputs(10050) <= not b or a;
    outputs(10051) <= a and not b;
    outputs(10052) <= a xor b;
    outputs(10053) <= a xor b;
    outputs(10054) <= a and not b;
    outputs(10055) <= b and not a;
    outputs(10056) <= a;
    outputs(10057) <= a xor b;
    outputs(10058) <= not b;
    outputs(10059) <= b and not a;
    outputs(10060) <= b;
    outputs(10061) <= a xor b;
    outputs(10062) <= a xor b;
    outputs(10063) <= not a;
    outputs(10064) <= not b;
    outputs(10065) <= not (a xor b);
    outputs(10066) <= a xor b;
    outputs(10067) <= a xor b;
    outputs(10068) <= a xor b;
    outputs(10069) <= not (a or b);
    outputs(10070) <= not a or b;
    outputs(10071) <= a or b;
    outputs(10072) <= a xor b;
    outputs(10073) <= a xor b;
    outputs(10074) <= a xor b;
    outputs(10075) <= a xor b;
    outputs(10076) <= not (a xor b);
    outputs(10077) <= not a;
    outputs(10078) <= a xor b;
    outputs(10079) <= not a or b;
    outputs(10080) <= not (a xor b);
    outputs(10081) <= b;
    outputs(10082) <= not a;
    outputs(10083) <= not (a and b);
    outputs(10084) <= a;
    outputs(10085) <= a;
    outputs(10086) <= a and not b;
    outputs(10087) <= not b or a;
    outputs(10088) <= a xor b;
    outputs(10089) <= a and b;
    outputs(10090) <= not a;
    outputs(10091) <= b;
    outputs(10092) <= not b;
    outputs(10093) <= b;
    outputs(10094) <= a and not b;
    outputs(10095) <= a and b;
    outputs(10096) <= not b;
    outputs(10097) <= a;
    outputs(10098) <= not (a xor b);
    outputs(10099) <= not b;
    outputs(10100) <= a and not b;
    outputs(10101) <= b;
    outputs(10102) <= not a;
    outputs(10103) <= not b;
    outputs(10104) <= a xor b;
    outputs(10105) <= a and b;
    outputs(10106) <= a xor b;
    outputs(10107) <= a xor b;
    outputs(10108) <= b;
    outputs(10109) <= not (a xor b);
    outputs(10110) <= b;
    outputs(10111) <= b and not a;
    outputs(10112) <= a;
    outputs(10113) <= a xor b;
    outputs(10114) <= a and b;
    outputs(10115) <= not (a xor b);
    outputs(10116) <= a;
    outputs(10117) <= a xor b;
    outputs(10118) <= not a;
    outputs(10119) <= a xor b;
    outputs(10120) <= not b or a;
    outputs(10121) <= a xor b;
    outputs(10122) <= not a or b;
    outputs(10123) <= b;
    outputs(10124) <= a and not b;
    outputs(10125) <= b and not a;
    outputs(10126) <= a and b;
    outputs(10127) <= not b;
    outputs(10128) <= a and b;
    outputs(10129) <= not (a xor b);
    outputs(10130) <= not (a xor b);
    outputs(10131) <= b;
    outputs(10132) <= not a;
    outputs(10133) <= not b or a;
    outputs(10134) <= not b;
    outputs(10135) <= not (a xor b);
    outputs(10136) <= b;
    outputs(10137) <= not a;
    outputs(10138) <= not b;
    outputs(10139) <= b;
    outputs(10140) <= b;
    outputs(10141) <= not (a xor b);
    outputs(10142) <= a xor b;
    outputs(10143) <= not (a xor b);
    outputs(10144) <= not (a and b);
    outputs(10145) <= b;
    outputs(10146) <= a xor b;
    outputs(10147) <= not b;
    outputs(10148) <= a xor b;
    outputs(10149) <= a;
    outputs(10150) <= not (a or b);
    outputs(10151) <= b;
    outputs(10152) <= a;
    outputs(10153) <= a xor b;
    outputs(10154) <= b;
    outputs(10155) <= not b;
    outputs(10156) <= a xor b;
    outputs(10157) <= a xor b;
    outputs(10158) <= not a;
    outputs(10159) <= not a;
    outputs(10160) <= b;
    outputs(10161) <= b and not a;
    outputs(10162) <= b;
    outputs(10163) <= b;
    outputs(10164) <= not (a xor b);
    outputs(10165) <= a and b;
    outputs(10166) <= a;
    outputs(10167) <= not a;
    outputs(10168) <= not (a or b);
    outputs(10169) <= a and b;
    outputs(10170) <= not b;
    outputs(10171) <= not b;
    outputs(10172) <= a and b;
    outputs(10173) <= not a;
    outputs(10174) <= not b;
    outputs(10175) <= a;
    outputs(10176) <= not b;
    outputs(10177) <= b and not a;
    outputs(10178) <= not a or b;
    outputs(10179) <= a xor b;
    outputs(10180) <= not b;
    outputs(10181) <= not (a and b);
    outputs(10182) <= a;
    outputs(10183) <= b;
    outputs(10184) <= not a;
    outputs(10185) <= not (a xor b);
    outputs(10186) <= not (a xor b);
    outputs(10187) <= b and not a;
    outputs(10188) <= a xor b;
    outputs(10189) <= not b;
    outputs(10190) <= a or b;
    outputs(10191) <= a xor b;
    outputs(10192) <= b;
    outputs(10193) <= not (a or b);
    outputs(10194) <= a;
    outputs(10195) <= a;
    outputs(10196) <= not (a xor b);
    outputs(10197) <= b and not a;
    outputs(10198) <= not (a xor b);
    outputs(10199) <= a xor b;
    outputs(10200) <= b and not a;
    outputs(10201) <= a xor b;
    outputs(10202) <= a xor b;
    outputs(10203) <= a and not b;
    outputs(10204) <= a;
    outputs(10205) <= a xor b;
    outputs(10206) <= a xor b;
    outputs(10207) <= a;
    outputs(10208) <= not (a xor b);
    outputs(10209) <= not (a or b);
    outputs(10210) <= not (a or b);
    outputs(10211) <= not a;
    outputs(10212) <= not (a xor b);
    outputs(10213) <= a;
    outputs(10214) <= not (a xor b);
    outputs(10215) <= b;
    outputs(10216) <= not (a xor b);
    outputs(10217) <= not b;
    outputs(10218) <= b and not a;
    outputs(10219) <= not (a xor b);
    outputs(10220) <= a and not b;
    outputs(10221) <= a and b;
    outputs(10222) <= a and not b;
    outputs(10223) <= a xor b;
    outputs(10224) <= b;
    outputs(10225) <= not (a xor b);
    outputs(10226) <= a and b;
    outputs(10227) <= not (a or b);
    outputs(10228) <= a;
    outputs(10229) <= b and not a;
    outputs(10230) <= b;
    outputs(10231) <= not a;
    outputs(10232) <= a;
    outputs(10233) <= a and b;
    outputs(10234) <= b and not a;
    outputs(10235) <= not a;
    outputs(10236) <= not a;
    outputs(10237) <= not a;
    outputs(10238) <= not (a or b);
    outputs(10239) <= not b;
    outputs(10240) <= not (a or b);
    outputs(10241) <= not a;
    outputs(10242) <= not b;
    outputs(10243) <= not (a xor b);
    outputs(10244) <= not (a xor b);
    outputs(10245) <= not a;
    outputs(10246) <= not (a xor b);
    outputs(10247) <= b;
    outputs(10248) <= a xor b;
    outputs(10249) <= not b;
    outputs(10250) <= a;
    outputs(10251) <= not (a xor b);
    outputs(10252) <= a xor b;
    outputs(10253) <= a;
    outputs(10254) <= a and b;
    outputs(10255) <= a;
    outputs(10256) <= not b;
    outputs(10257) <= not b;
    outputs(10258) <= not (a and b);
    outputs(10259) <= b;
    outputs(10260) <= b;
    outputs(10261) <= a xor b;
    outputs(10262) <= not a or b;
    outputs(10263) <= a or b;
    outputs(10264) <= b;
    outputs(10265) <= not b or a;
    outputs(10266) <= not (a or b);
    outputs(10267) <= a and b;
    outputs(10268) <= not (a xor b);
    outputs(10269) <= not a;
    outputs(10270) <= not a;
    outputs(10271) <= not a;
    outputs(10272) <= a xor b;
    outputs(10273) <= not a;
    outputs(10274) <= b;
    outputs(10275) <= not (a xor b);
    outputs(10276) <= b and not a;
    outputs(10277) <= b and not a;
    outputs(10278) <= not (a xor b);
    outputs(10279) <= a xor b;
    outputs(10280) <= a and b;
    outputs(10281) <= b and not a;
    outputs(10282) <= a;
    outputs(10283) <= a xor b;
    outputs(10284) <= a xor b;
    outputs(10285) <= a;
    outputs(10286) <= not (a and b);
    outputs(10287) <= a xor b;
    outputs(10288) <= a or b;
    outputs(10289) <= a xor b;
    outputs(10290) <= b and not a;
    outputs(10291) <= not b;
    outputs(10292) <= not b;
    outputs(10293) <= not b;
    outputs(10294) <= not b;
    outputs(10295) <= a xor b;
    outputs(10296) <= not a or b;
    outputs(10297) <= a;
    outputs(10298) <= not (a xor b);
    outputs(10299) <= a or b;
    outputs(10300) <= b;
    outputs(10301) <= not a;
    outputs(10302) <= not b;
    outputs(10303) <= not (a xor b);
    outputs(10304) <= not a or b;
    outputs(10305) <= a;
    outputs(10306) <= not (a xor b);
    outputs(10307) <= not (a xor b);
    outputs(10308) <= not (a xor b);
    outputs(10309) <= b;
    outputs(10310) <= a xor b;
    outputs(10311) <= a xor b;
    outputs(10312) <= not a;
    outputs(10313) <= not a;
    outputs(10314) <= not (a xor b);
    outputs(10315) <= a xor b;
    outputs(10316) <= not a;
    outputs(10317) <= not a or b;
    outputs(10318) <= a;
    outputs(10319) <= not (a xor b);
    outputs(10320) <= a and not b;
    outputs(10321) <= a xor b;
    outputs(10322) <= a xor b;
    outputs(10323) <= a xor b;
    outputs(10324) <= not (a and b);
    outputs(10325) <= b;
    outputs(10326) <= not a;
    outputs(10327) <= a;
    outputs(10328) <= not b;
    outputs(10329) <= not a;
    outputs(10330) <= not (a and b);
    outputs(10331) <= a;
    outputs(10332) <= a;
    outputs(10333) <= a xor b;
    outputs(10334) <= not b;
    outputs(10335) <= a xor b;
    outputs(10336) <= b;
    outputs(10337) <= not a;
    outputs(10338) <= a;
    outputs(10339) <= a xor b;
    outputs(10340) <= not (a xor b);
    outputs(10341) <= not b;
    outputs(10342) <= a;
    outputs(10343) <= not a or b;
    outputs(10344) <= a xor b;
    outputs(10345) <= a xor b;
    outputs(10346) <= a xor b;
    outputs(10347) <= not a;
    outputs(10348) <= not b;
    outputs(10349) <= not (a xor b);
    outputs(10350) <= b;
    outputs(10351) <= not (a or b);
    outputs(10352) <= not b;
    outputs(10353) <= b;
    outputs(10354) <= not a or b;
    outputs(10355) <= not b;
    outputs(10356) <= not (a xor b);
    outputs(10357) <= not (a or b);
    outputs(10358) <= not a;
    outputs(10359) <= not (a xor b);
    outputs(10360) <= b;
    outputs(10361) <= not (a xor b);
    outputs(10362) <= a xor b;
    outputs(10363) <= not b;
    outputs(10364) <= not b;
    outputs(10365) <= b;
    outputs(10366) <= a and not b;
    outputs(10367) <= not a;
    outputs(10368) <= not b;
    outputs(10369) <= not a;
    outputs(10370) <= b;
    outputs(10371) <= a xor b;
    outputs(10372) <= not (a and b);
    outputs(10373) <= not b;
    outputs(10374) <= b;
    outputs(10375) <= b;
    outputs(10376) <= not b;
    outputs(10377) <= not (a and b);
    outputs(10378) <= b;
    outputs(10379) <= b;
    outputs(10380) <= not (a xor b);
    outputs(10381) <= not (a or b);
    outputs(10382) <= b and not a;
    outputs(10383) <= not b;
    outputs(10384) <= b;
    outputs(10385) <= a or b;
    outputs(10386) <= a;
    outputs(10387) <= not a;
    outputs(10388) <= not b or a;
    outputs(10389) <= not (a xor b);
    outputs(10390) <= not a;
    outputs(10391) <= not (a or b);
    outputs(10392) <= not (a xor b);
    outputs(10393) <= b;
    outputs(10394) <= b;
    outputs(10395) <= a and not b;
    outputs(10396) <= a xor b;
    outputs(10397) <= not b or a;
    outputs(10398) <= a;
    outputs(10399) <= a or b;
    outputs(10400) <= b;
    outputs(10401) <= not (a xor b);
    outputs(10402) <= a xor b;
    outputs(10403) <= a xor b;
    outputs(10404) <= not a;
    outputs(10405) <= b and not a;
    outputs(10406) <= not a or b;
    outputs(10407) <= b;
    outputs(10408) <= b and not a;
    outputs(10409) <= not a;
    outputs(10410) <= not a;
    outputs(10411) <= a xor b;
    outputs(10412) <= not (a and b);
    outputs(10413) <= not a;
    outputs(10414) <= not a;
    outputs(10415) <= not (a xor b);
    outputs(10416) <= a xor b;
    outputs(10417) <= not (a xor b);
    outputs(10418) <= not b;
    outputs(10419) <= not a;
    outputs(10420) <= a and b;
    outputs(10421) <= a xor b;
    outputs(10422) <= not (a xor b);
    outputs(10423) <= a and b;
    outputs(10424) <= not (a xor b);
    outputs(10425) <= not a or b;
    outputs(10426) <= not b;
    outputs(10427) <= b;
    outputs(10428) <= a or b;
    outputs(10429) <= not b;
    outputs(10430) <= not b or a;
    outputs(10431) <= a;
    outputs(10432) <= not b;
    outputs(10433) <= not a;
    outputs(10434) <= not (a xor b);
    outputs(10435) <= not (a and b);
    outputs(10436) <= a or b;
    outputs(10437) <= a xor b;
    outputs(10438) <= b and not a;
    outputs(10439) <= not a or b;
    outputs(10440) <= not (a xor b);
    outputs(10441) <= not (a xor b);
    outputs(10442) <= a xor b;
    outputs(10443) <= not (a and b);
    outputs(10444) <= b;
    outputs(10445) <= not b or a;
    outputs(10446) <= not (a xor b);
    outputs(10447) <= a xor b;
    outputs(10448) <= a xor b;
    outputs(10449) <= b;
    outputs(10450) <= not (a xor b);
    outputs(10451) <= not b or a;
    outputs(10452) <= a xor b;
    outputs(10453) <= not (a xor b);
    outputs(10454) <= not b;
    outputs(10455) <= not b;
    outputs(10456) <= not b or a;
    outputs(10457) <= a;
    outputs(10458) <= not a;
    outputs(10459) <= a xor b;
    outputs(10460) <= a;
    outputs(10461) <= not a;
    outputs(10462) <= not a or b;
    outputs(10463) <= not b;
    outputs(10464) <= b;
    outputs(10465) <= not (a xor b);
    outputs(10466) <= a xor b;
    outputs(10467) <= b;
    outputs(10468) <= a xor b;
    outputs(10469) <= b and not a;
    outputs(10470) <= not (a xor b);
    outputs(10471) <= not (a xor b);
    outputs(10472) <= not (a xor b);
    outputs(10473) <= a xor b;
    outputs(10474) <= not (a xor b);
    outputs(10475) <= not b or a;
    outputs(10476) <= not b;
    outputs(10477) <= a and b;
    outputs(10478) <= not (a xor b);
    outputs(10479) <= a;
    outputs(10480) <= not b;
    outputs(10481) <= a xor b;
    outputs(10482) <= not (a xor b);
    outputs(10483) <= not a or b;
    outputs(10484) <= a xor b;
    outputs(10485) <= a;
    outputs(10486) <= not b or a;
    outputs(10487) <= not a;
    outputs(10488) <= a xor b;
    outputs(10489) <= a xor b;
    outputs(10490) <= not b;
    outputs(10491) <= a xor b;
    outputs(10492) <= a and not b;
    outputs(10493) <= not (a xor b);
    outputs(10494) <= not a;
    outputs(10495) <= a xor b;
    outputs(10496) <= a xor b;
    outputs(10497) <= b;
    outputs(10498) <= b;
    outputs(10499) <= b;
    outputs(10500) <= not (a xor b);
    outputs(10501) <= a xor b;
    outputs(10502) <= a and b;
    outputs(10503) <= a xor b;
    outputs(10504) <= not a;
    outputs(10505) <= not (a xor b);
    outputs(10506) <= not (a xor b);
    outputs(10507) <= not b;
    outputs(10508) <= not a;
    outputs(10509) <= b and not a;
    outputs(10510) <= not a;
    outputs(10511) <= a xor b;
    outputs(10512) <= a;
    outputs(10513) <= not b or a;
    outputs(10514) <= a xor b;
    outputs(10515) <= a xor b;
    outputs(10516) <= a xor b;
    outputs(10517) <= b;
    outputs(10518) <= a xor b;
    outputs(10519) <= not (a xor b);
    outputs(10520) <= a xor b;
    outputs(10521) <= not b;
    outputs(10522) <= not (a xor b);
    outputs(10523) <= not (a xor b);
    outputs(10524) <= a;
    outputs(10525) <= not b or a;
    outputs(10526) <= a xor b;
    outputs(10527) <= a xor b;
    outputs(10528) <= a;
    outputs(10529) <= not (a xor b);
    outputs(10530) <= b and not a;
    outputs(10531) <= not (a xor b);
    outputs(10532) <= b;
    outputs(10533) <= not (a xor b);
    outputs(10534) <= not (a and b);
    outputs(10535) <= a xor b;
    outputs(10536) <= a;
    outputs(10537) <= not a;
    outputs(10538) <= b and not a;
    outputs(10539) <= b;
    outputs(10540) <= a;
    outputs(10541) <= a xor b;
    outputs(10542) <= not a or b;
    outputs(10543) <= not a or b;
    outputs(10544) <= a;
    outputs(10545) <= not b;
    outputs(10546) <= not b;
    outputs(10547) <= b;
    outputs(10548) <= a xor b;
    outputs(10549) <= a xor b;
    outputs(10550) <= not a;
    outputs(10551) <= a;
    outputs(10552) <= not a;
    outputs(10553) <= a xor b;
    outputs(10554) <= a and not b;
    outputs(10555) <= not b;
    outputs(10556) <= a xor b;
    outputs(10557) <= not (a xor b);
    outputs(10558) <= not (a and b);
    outputs(10559) <= a;
    outputs(10560) <= not a;
    outputs(10561) <= a or b;
    outputs(10562) <= not a or b;
    outputs(10563) <= not (a xor b);
    outputs(10564) <= a xor b;
    outputs(10565) <= a and b;
    outputs(10566) <= not a or b;
    outputs(10567) <= b;
    outputs(10568) <= b;
    outputs(10569) <= not (a xor b);
    outputs(10570) <= not b;
    outputs(10571) <= a;
    outputs(10572) <= a xor b;
    outputs(10573) <= a;
    outputs(10574) <= a xor b;
    outputs(10575) <= a xor b;
    outputs(10576) <= not a;
    outputs(10577) <= b;
    outputs(10578) <= a xor b;
    outputs(10579) <= b;
    outputs(10580) <= not b or a;
    outputs(10581) <= a xor b;
    outputs(10582) <= not (a or b);
    outputs(10583) <= not a;
    outputs(10584) <= a;
    outputs(10585) <= not (a xor b);
    outputs(10586) <= not b;
    outputs(10587) <= a;
    outputs(10588) <= b and not a;
    outputs(10589) <= a xor b;
    outputs(10590) <= b;
    outputs(10591) <= a or b;
    outputs(10592) <= not b;
    outputs(10593) <= b;
    outputs(10594) <= a xor b;
    outputs(10595) <= not b;
    outputs(10596) <= b;
    outputs(10597) <= not (a xor b);
    outputs(10598) <= b;
    outputs(10599) <= not b;
    outputs(10600) <= b;
    outputs(10601) <= not (a xor b);
    outputs(10602) <= a xor b;
    outputs(10603) <= a;
    outputs(10604) <= a xor b;
    outputs(10605) <= a xor b;
    outputs(10606) <= not a or b;
    outputs(10607) <= not a;
    outputs(10608) <= a xor b;
    outputs(10609) <= b;
    outputs(10610) <= not (a xor b);
    outputs(10611) <= not a;
    outputs(10612) <= a xor b;
    outputs(10613) <= b;
    outputs(10614) <= not a;
    outputs(10615) <= a;
    outputs(10616) <= not b or a;
    outputs(10617) <= a and not b;
    outputs(10618) <= b;
    outputs(10619) <= a xor b;
    outputs(10620) <= not b or a;
    outputs(10621) <= not b;
    outputs(10622) <= b;
    outputs(10623) <= not (a xor b);
    outputs(10624) <= a xor b;
    outputs(10625) <= not b;
    outputs(10626) <= a xor b;
    outputs(10627) <= not (a and b);
    outputs(10628) <= a;
    outputs(10629) <= not b;
    outputs(10630) <= a xor b;
    outputs(10631) <= not (a xor b);
    outputs(10632) <= not (a xor b);
    outputs(10633) <= a xor b;
    outputs(10634) <= not b;
    outputs(10635) <= a or b;
    outputs(10636) <= not (a xor b);
    outputs(10637) <= a xor b;
    outputs(10638) <= not b;
    outputs(10639) <= a;
    outputs(10640) <= b and not a;
    outputs(10641) <= not a;
    outputs(10642) <= a;
    outputs(10643) <= a;
    outputs(10644) <= not b;
    outputs(10645) <= not (a xor b);
    outputs(10646) <= b and not a;
    outputs(10647) <= not b;
    outputs(10648) <= a;
    outputs(10649) <= a xor b;
    outputs(10650) <= a xor b;
    outputs(10651) <= not (a xor b);
    outputs(10652) <= not a;
    outputs(10653) <= not a or b;
    outputs(10654) <= a and b;
    outputs(10655) <= not (a and b);
    outputs(10656) <= a and b;
    outputs(10657) <= a;
    outputs(10658) <= not b;
    outputs(10659) <= not a;
    outputs(10660) <= a;
    outputs(10661) <= a or b;
    outputs(10662) <= not (a xor b);
    outputs(10663) <= not (a xor b);
    outputs(10664) <= b and not a;
    outputs(10665) <= not (a or b);
    outputs(10666) <= b;
    outputs(10667) <= a xor b;
    outputs(10668) <= b;
    outputs(10669) <= not (a xor b);
    outputs(10670) <= not b;
    outputs(10671) <= a;
    outputs(10672) <= not (a xor b);
    outputs(10673) <= a;
    outputs(10674) <= a or b;
    outputs(10675) <= a;
    outputs(10676) <= not (a or b);
    outputs(10677) <= not (a xor b);
    outputs(10678) <= not a;
    outputs(10679) <= b;
    outputs(10680) <= a xor b;
    outputs(10681) <= not b or a;
    outputs(10682) <= not a;
    outputs(10683) <= not a;
    outputs(10684) <= a xor b;
    outputs(10685) <= a xor b;
    outputs(10686) <= not a or b;
    outputs(10687) <= a or b;
    outputs(10688) <= not (a xor b);
    outputs(10689) <= not (a xor b);
    outputs(10690) <= not (a or b);
    outputs(10691) <= not b;
    outputs(10692) <= not b;
    outputs(10693) <= not (a xor b);
    outputs(10694) <= not (a xor b);
    outputs(10695) <= not (a xor b);
    outputs(10696) <= a;
    outputs(10697) <= a and b;
    outputs(10698) <= not a;
    outputs(10699) <= a xor b;
    outputs(10700) <= not (a or b);
    outputs(10701) <= a xor b;
    outputs(10702) <= not b;
    outputs(10703) <= not a;
    outputs(10704) <= not (a xor b);
    outputs(10705) <= not (a xor b);
    outputs(10706) <= a xor b;
    outputs(10707) <= not (a xor b);
    outputs(10708) <= a or b;
    outputs(10709) <= b;
    outputs(10710) <= not a or b;
    outputs(10711) <= b;
    outputs(10712) <= not a or b;
    outputs(10713) <= not (a or b);
    outputs(10714) <= a xor b;
    outputs(10715) <= not b;
    outputs(10716) <= not (a xor b);
    outputs(10717) <= b and not a;
    outputs(10718) <= not b or a;
    outputs(10719) <= not b or a;
    outputs(10720) <= not (a xor b);
    outputs(10721) <= a;
    outputs(10722) <= a;
    outputs(10723) <= a and not b;
    outputs(10724) <= a;
    outputs(10725) <= not a or b;
    outputs(10726) <= b;
    outputs(10727) <= not (a xor b);
    outputs(10728) <= a;
    outputs(10729) <= not a;
    outputs(10730) <= not b;
    outputs(10731) <= not b;
    outputs(10732) <= not a;
    outputs(10733) <= b;
    outputs(10734) <= not (a xor b);
    outputs(10735) <= a xor b;
    outputs(10736) <= a xor b;
    outputs(10737) <= a xor b;
    outputs(10738) <= not b;
    outputs(10739) <= not (a xor b);
    outputs(10740) <= not b;
    outputs(10741) <= not a or b;
    outputs(10742) <= b and not a;
    outputs(10743) <= not b;
    outputs(10744) <= not (a xor b);
    outputs(10745) <= not b or a;
    outputs(10746) <= a and not b;
    outputs(10747) <= b;
    outputs(10748) <= not b or a;
    outputs(10749) <= not b or a;
    outputs(10750) <= b;
    outputs(10751) <= not a;
    outputs(10752) <= b;
    outputs(10753) <= not b;
    outputs(10754) <= not b;
    outputs(10755) <= b and not a;
    outputs(10756) <= not b or a;
    outputs(10757) <= b;
    outputs(10758) <= not (a xor b);
    outputs(10759) <= b;
    outputs(10760) <= not b;
    outputs(10761) <= a;
    outputs(10762) <= a xor b;
    outputs(10763) <= not b;
    outputs(10764) <= a;
    outputs(10765) <= a xor b;
    outputs(10766) <= a xor b;
    outputs(10767) <= a xor b;
    outputs(10768) <= not (a or b);
    outputs(10769) <= not (a xor b);
    outputs(10770) <= not (a and b);
    outputs(10771) <= a xor b;
    outputs(10772) <= a;
    outputs(10773) <= not b;
    outputs(10774) <= a;
    outputs(10775) <= a;
    outputs(10776) <= not (a or b);
    outputs(10777) <= not b;
    outputs(10778) <= not (a xor b);
    outputs(10779) <= not b;
    outputs(10780) <= not (a and b);
    outputs(10781) <= not a or b;
    outputs(10782) <= not a;
    outputs(10783) <= not (a xor b);
    outputs(10784) <= not (a xor b);
    outputs(10785) <= a;
    outputs(10786) <= b;
    outputs(10787) <= a xor b;
    outputs(10788) <= b;
    outputs(10789) <= a;
    outputs(10790) <= a;
    outputs(10791) <= a;
    outputs(10792) <= a xor b;
    outputs(10793) <= not (a xor b);
    outputs(10794) <= a xor b;
    outputs(10795) <= not (a xor b);
    outputs(10796) <= a xor b;
    outputs(10797) <= a xor b;
    outputs(10798) <= b;
    outputs(10799) <= a or b;
    outputs(10800) <= not a;
    outputs(10801) <= not a;
    outputs(10802) <= a;
    outputs(10803) <= not (a or b);
    outputs(10804) <= not (a xor b);
    outputs(10805) <= not (a or b);
    outputs(10806) <= not a;
    outputs(10807) <= b;
    outputs(10808) <= a and not b;
    outputs(10809) <= a and b;
    outputs(10810) <= a xor b;
    outputs(10811) <= not (a xor b);
    outputs(10812) <= not (a xor b);
    outputs(10813) <= not a or b;
    outputs(10814) <= not a;
    outputs(10815) <= b;
    outputs(10816) <= a xor b;
    outputs(10817) <= not (a xor b);
    outputs(10818) <= not b;
    outputs(10819) <= not a;
    outputs(10820) <= not (a xor b);
    outputs(10821) <= not (a xor b);
    outputs(10822) <= not (a xor b);
    outputs(10823) <= a;
    outputs(10824) <= a or b;
    outputs(10825) <= not (a xor b);
    outputs(10826) <= a xor b;
    outputs(10827) <= a;
    outputs(10828) <= a;
    outputs(10829) <= not (a or b);
    outputs(10830) <= b and not a;
    outputs(10831) <= a xor b;
    outputs(10832) <= not a or b;
    outputs(10833) <= a and b;
    outputs(10834) <= not a;
    outputs(10835) <= b;
    outputs(10836) <= not b;
    outputs(10837) <= not b or a;
    outputs(10838) <= not b;
    outputs(10839) <= not (a xor b);
    outputs(10840) <= not (a and b);
    outputs(10841) <= a and b;
    outputs(10842) <= not (a xor b);
    outputs(10843) <= a xor b;
    outputs(10844) <= not b;
    outputs(10845) <= a xor b;
    outputs(10846) <= b;
    outputs(10847) <= b;
    outputs(10848) <= not (a xor b);
    outputs(10849) <= not (a xor b);
    outputs(10850) <= not a;
    outputs(10851) <= not b;
    outputs(10852) <= a xor b;
    outputs(10853) <= not a;
    outputs(10854) <= not b;
    outputs(10855) <= a or b;
    outputs(10856) <= not a;
    outputs(10857) <= a xor b;
    outputs(10858) <= not a;
    outputs(10859) <= a xor b;
    outputs(10860) <= not (a xor b);
    outputs(10861) <= not b;
    outputs(10862) <= b;
    outputs(10863) <= a or b;
    outputs(10864) <= a xor b;
    outputs(10865) <= a xor b;
    outputs(10866) <= a xor b;
    outputs(10867) <= not a or b;
    outputs(10868) <= a xor b;
    outputs(10869) <= not b;
    outputs(10870) <= not (a xor b);
    outputs(10871) <= not (a xor b);
    outputs(10872) <= a xor b;
    outputs(10873) <= a or b;
    outputs(10874) <= b;
    outputs(10875) <= not a;
    outputs(10876) <= not (a xor b);
    outputs(10877) <= a xor b;
    outputs(10878) <= a xor b;
    outputs(10879) <= b and not a;
    outputs(10880) <= not (a xor b);
    outputs(10881) <= a xor b;
    outputs(10882) <= a xor b;
    outputs(10883) <= not b or a;
    outputs(10884) <= not a or b;
    outputs(10885) <= a;
    outputs(10886) <= a xor b;
    outputs(10887) <= not (a xor b);
    outputs(10888) <= not (a xor b);
    outputs(10889) <= not b;
    outputs(10890) <= not a;
    outputs(10891) <= b;
    outputs(10892) <= a;
    outputs(10893) <= a or b;
    outputs(10894) <= not b;
    outputs(10895) <= not b or a;
    outputs(10896) <= not (a or b);
    outputs(10897) <= not a or b;
    outputs(10898) <= not (a xor b);
    outputs(10899) <= a or b;
    outputs(10900) <= not a or b;
    outputs(10901) <= not (a xor b);
    outputs(10902) <= not b;
    outputs(10903) <= not (a xor b);
    outputs(10904) <= not (a xor b);
    outputs(10905) <= not b;
    outputs(10906) <= b;
    outputs(10907) <= a or b;
    outputs(10908) <= b;
    outputs(10909) <= a and not b;
    outputs(10910) <= a;
    outputs(10911) <= a xor b;
    outputs(10912) <= not a;
    outputs(10913) <= not (a or b);
    outputs(10914) <= a or b;
    outputs(10915) <= not b;
    outputs(10916) <= a or b;
    outputs(10917) <= b and not a;
    outputs(10918) <= a;
    outputs(10919) <= a;
    outputs(10920) <= not a;
    outputs(10921) <= b;
    outputs(10922) <= not b;
    outputs(10923) <= a xor b;
    outputs(10924) <= not a;
    outputs(10925) <= not a;
    outputs(10926) <= b and not a;
    outputs(10927) <= b;
    outputs(10928) <= a;
    outputs(10929) <= not b;
    outputs(10930) <= not (a xor b);
    outputs(10931) <= not (a xor b);
    outputs(10932) <= not b;
    outputs(10933) <= not b or a;
    outputs(10934) <= a xor b;
    outputs(10935) <= a and not b;
    outputs(10936) <= not (a and b);
    outputs(10937) <= not a or b;
    outputs(10938) <= not (a or b);
    outputs(10939) <= a or b;
    outputs(10940) <= b;
    outputs(10941) <= not a or b;
    outputs(10942) <= not a;
    outputs(10943) <= b;
    outputs(10944) <= not (a xor b);
    outputs(10945) <= not (a xor b);
    outputs(10946) <= b;
    outputs(10947) <= b;
    outputs(10948) <= a and b;
    outputs(10949) <= a xor b;
    outputs(10950) <= a xor b;
    outputs(10951) <= not b or a;
    outputs(10952) <= not b;
    outputs(10953) <= a xor b;
    outputs(10954) <= b;
    outputs(10955) <= b;
    outputs(10956) <= a xor b;
    outputs(10957) <= not (a or b);
    outputs(10958) <= not b;
    outputs(10959) <= a;
    outputs(10960) <= not (a xor b);
    outputs(10961) <= b;
    outputs(10962) <= a;
    outputs(10963) <= a xor b;
    outputs(10964) <= not (a xor b);
    outputs(10965) <= b;
    outputs(10966) <= not (a xor b);
    outputs(10967) <= b;
    outputs(10968) <= b;
    outputs(10969) <= a xor b;
    outputs(10970) <= not b or a;
    outputs(10971) <= a or b;
    outputs(10972) <= not (a and b);
    outputs(10973) <= a xor b;
    outputs(10974) <= not (a or b);
    outputs(10975) <= a;
    outputs(10976) <= a xor b;
    outputs(10977) <= a;
    outputs(10978) <= b;
    outputs(10979) <= a;
    outputs(10980) <= a xor b;
    outputs(10981) <= b;
    outputs(10982) <= b;
    outputs(10983) <= a xor b;
    outputs(10984) <= not (a and b);
    outputs(10985) <= not a or b;
    outputs(10986) <= a xor b;
    outputs(10987) <= a;
    outputs(10988) <= not (a or b);
    outputs(10989) <= a;
    outputs(10990) <= a;
    outputs(10991) <= a xor b;
    outputs(10992) <= not (a xor b);
    outputs(10993) <= a;
    outputs(10994) <= b and not a;
    outputs(10995) <= a xor b;
    outputs(10996) <= not b;
    outputs(10997) <= not a;
    outputs(10998) <= not (a xor b);
    outputs(10999) <= not (a xor b);
    outputs(11000) <= not a;
    outputs(11001) <= a xor b;
    outputs(11002) <= not (a xor b);
    outputs(11003) <= a;
    outputs(11004) <= not (a or b);
    outputs(11005) <= not b;
    outputs(11006) <= b and not a;
    outputs(11007) <= a or b;
    outputs(11008) <= a xor b;
    outputs(11009) <= a and b;
    outputs(11010) <= not b or a;
    outputs(11011) <= not a;
    outputs(11012) <= a;
    outputs(11013) <= b;
    outputs(11014) <= not (a xor b);
    outputs(11015) <= a xor b;
    outputs(11016) <= a or b;
    outputs(11017) <= not b or a;
    outputs(11018) <= not (a xor b);
    outputs(11019) <= b;
    outputs(11020) <= a;
    outputs(11021) <= a xor b;
    outputs(11022) <= not (a xor b);
    outputs(11023) <= a xor b;
    outputs(11024) <= not b;
    outputs(11025) <= b and not a;
    outputs(11026) <= not b;
    outputs(11027) <= not a or b;
    outputs(11028) <= b;
    outputs(11029) <= not (a and b);
    outputs(11030) <= a;
    outputs(11031) <= not (a xor b);
    outputs(11032) <= not (a xor b);
    outputs(11033) <= not (a and b);
    outputs(11034) <= a xor b;
    outputs(11035) <= b;
    outputs(11036) <= a and not b;
    outputs(11037) <= a xor b;
    outputs(11038) <= not (a xor b);
    outputs(11039) <= not b;
    outputs(11040) <= not a;
    outputs(11041) <= a and not b;
    outputs(11042) <= not (a or b);
    outputs(11043) <= not (a and b);
    outputs(11044) <= not (a or b);
    outputs(11045) <= not (a xor b);
    outputs(11046) <= not a;
    outputs(11047) <= not (a xor b);
    outputs(11048) <= a xor b;
    outputs(11049) <= a;
    outputs(11050) <= not b;
    outputs(11051) <= not b;
    outputs(11052) <= not b;
    outputs(11053) <= not (a xor b);
    outputs(11054) <= not (a xor b);
    outputs(11055) <= a xor b;
    outputs(11056) <= a xor b;
    outputs(11057) <= not (a xor b);
    outputs(11058) <= not b;
    outputs(11059) <= not b;
    outputs(11060) <= a;
    outputs(11061) <= a;
    outputs(11062) <= not b;
    outputs(11063) <= not a;
    outputs(11064) <= b;
    outputs(11065) <= a xor b;
    outputs(11066) <= not b or a;
    outputs(11067) <= not b;
    outputs(11068) <= a;
    outputs(11069) <= a;
    outputs(11070) <= not (a xor b);
    outputs(11071) <= b;
    outputs(11072) <= not b or a;
    outputs(11073) <= not (a or b);
    outputs(11074) <= b;
    outputs(11075) <= not (a xor b);
    outputs(11076) <= not (a xor b);
    outputs(11077) <= not a or b;
    outputs(11078) <= a xor b;
    outputs(11079) <= not (a xor b);
    outputs(11080) <= not (a xor b);
    outputs(11081) <= not (a and b);
    outputs(11082) <= b;
    outputs(11083) <= a xor b;
    outputs(11084) <= not b;
    outputs(11085) <= a or b;
    outputs(11086) <= not (a xor b);
    outputs(11087) <= not (a xor b);
    outputs(11088) <= a;
    outputs(11089) <= a xor b;
    outputs(11090) <= not (a xor b);
    outputs(11091) <= b and not a;
    outputs(11092) <= not (a xor b);
    outputs(11093) <= not (a xor b);
    outputs(11094) <= a and b;
    outputs(11095) <= b;
    outputs(11096) <= not b;
    outputs(11097) <= not (a or b);
    outputs(11098) <= a xor b;
    outputs(11099) <= not (a xor b);
    outputs(11100) <= not b;
    outputs(11101) <= not a;
    outputs(11102) <= a;
    outputs(11103) <= not a;
    outputs(11104) <= not b;
    outputs(11105) <= a;
    outputs(11106) <= not (a or b);
    outputs(11107) <= not a;
    outputs(11108) <= a;
    outputs(11109) <= not a;
    outputs(11110) <= a;
    outputs(11111) <= not b or a;
    outputs(11112) <= b;
    outputs(11113) <= not (a xor b);
    outputs(11114) <= a;
    outputs(11115) <= not b;
    outputs(11116) <= a or b;
    outputs(11117) <= b and not a;
    outputs(11118) <= a xor b;
    outputs(11119) <= not b;
    outputs(11120) <= a and not b;
    outputs(11121) <= a xor b;
    outputs(11122) <= b;
    outputs(11123) <= a or b;
    outputs(11124) <= a;
    outputs(11125) <= a;
    outputs(11126) <= not a;
    outputs(11127) <= a xor b;
    outputs(11128) <= not b or a;
    outputs(11129) <= not b;
    outputs(11130) <= not b;
    outputs(11131) <= a or b;
    outputs(11132) <= not (a or b);
    outputs(11133) <= b;
    outputs(11134) <= not a;
    outputs(11135) <= not (a and b);
    outputs(11136) <= not a;
    outputs(11137) <= not b;
    outputs(11138) <= not (a and b);
    outputs(11139) <= not (a xor b);
    outputs(11140) <= not a;
    outputs(11141) <= not b or a;
    outputs(11142) <= not b or a;
    outputs(11143) <= not (a xor b);
    outputs(11144) <= not b;
    outputs(11145) <= not b;
    outputs(11146) <= a;
    outputs(11147) <= not a;
    outputs(11148) <= not (a xor b);
    outputs(11149) <= a xor b;
    outputs(11150) <= not b;
    outputs(11151) <= not a;
    outputs(11152) <= not (a xor b);
    outputs(11153) <= a xor b;
    outputs(11154) <= not (a and b);
    outputs(11155) <= not a or b;
    outputs(11156) <= not (a xor b);
    outputs(11157) <= not b;
    outputs(11158) <= a xor b;
    outputs(11159) <= not (a and b);
    outputs(11160) <= not (a xor b);
    outputs(11161) <= not (a xor b);
    outputs(11162) <= a;
    outputs(11163) <= a and not b;
    outputs(11164) <= not (a xor b);
    outputs(11165) <= not b or a;
    outputs(11166) <= not b;
    outputs(11167) <= b;
    outputs(11168) <= not a;
    outputs(11169) <= a;
    outputs(11170) <= not (a and b);
    outputs(11171) <= not (a xor b);
    outputs(11172) <= not (a xor b);
    outputs(11173) <= a and not b;
    outputs(11174) <= not a or b;
    outputs(11175) <= not b;
    outputs(11176) <= not a or b;
    outputs(11177) <= a xor b;
    outputs(11178) <= not a;
    outputs(11179) <= not b or a;
    outputs(11180) <= not a;
    outputs(11181) <= not a;
    outputs(11182) <= not a or b;
    outputs(11183) <= not a or b;
    outputs(11184) <= a xor b;
    outputs(11185) <= a;
    outputs(11186) <= not a or b;
    outputs(11187) <= a xor b;
    outputs(11188) <= b;
    outputs(11189) <= not a or b;
    outputs(11190) <= a and not b;
    outputs(11191) <= not (a xor b);
    outputs(11192) <= a;
    outputs(11193) <= a xor b;
    outputs(11194) <= not a;
    outputs(11195) <= b;
    outputs(11196) <= not (a xor b);
    outputs(11197) <= not a;
    outputs(11198) <= b;
    outputs(11199) <= not b;
    outputs(11200) <= a and not b;
    outputs(11201) <= a;
    outputs(11202) <= a and not b;
    outputs(11203) <= not (a or b);
    outputs(11204) <= not a;
    outputs(11205) <= b;
    outputs(11206) <= not a or b;
    outputs(11207) <= a;
    outputs(11208) <= a and not b;
    outputs(11209) <= a xor b;
    outputs(11210) <= not (a xor b);
    outputs(11211) <= not (a xor b);
    outputs(11212) <= a;
    outputs(11213) <= a xor b;
    outputs(11214) <= a xor b;
    outputs(11215) <= a or b;
    outputs(11216) <= a;
    outputs(11217) <= not b;
    outputs(11218) <= b and not a;
    outputs(11219) <= a and not b;
    outputs(11220) <= not (a xor b);
    outputs(11221) <= not b;
    outputs(11222) <= a or b;
    outputs(11223) <= not a;
    outputs(11224) <= a;
    outputs(11225) <= a;
    outputs(11226) <= not (a xor b);
    outputs(11227) <= not b;
    outputs(11228) <= not b;
    outputs(11229) <= a;
    outputs(11230) <= not (a xor b);
    outputs(11231) <= not a;
    outputs(11232) <= not a;
    outputs(11233) <= not (a xor b);
    outputs(11234) <= not (a xor b);
    outputs(11235) <= not (a xor b);
    outputs(11236) <= b;
    outputs(11237) <= not (a xor b);
    outputs(11238) <= not a or b;
    outputs(11239) <= a xor b;
    outputs(11240) <= a;
    outputs(11241) <= a;
    outputs(11242) <= not (a xor b);
    outputs(11243) <= a and not b;
    outputs(11244) <= not (a xor b);
    outputs(11245) <= not b or a;
    outputs(11246) <= a;
    outputs(11247) <= a xor b;
    outputs(11248) <= a xor b;
    outputs(11249) <= a xor b;
    outputs(11250) <= not (a xor b);
    outputs(11251) <= a xor b;
    outputs(11252) <= a xor b;
    outputs(11253) <= b;
    outputs(11254) <= not (a xor b);
    outputs(11255) <= not b;
    outputs(11256) <= a;
    outputs(11257) <= not (a xor b);
    outputs(11258) <= not b or a;
    outputs(11259) <= not b;
    outputs(11260) <= not (a xor b);
    outputs(11261) <= b;
    outputs(11262) <= not (a and b);
    outputs(11263) <= a or b;
    outputs(11264) <= a;
    outputs(11265) <= b;
    outputs(11266) <= a and b;
    outputs(11267) <= a xor b;
    outputs(11268) <= not b;
    outputs(11269) <= not (a xor b);
    outputs(11270) <= not (a xor b);
    outputs(11271) <= not a;
    outputs(11272) <= a;
    outputs(11273) <= a xor b;
    outputs(11274) <= a;
    outputs(11275) <= a or b;
    outputs(11276) <= not (a and b);
    outputs(11277) <= not b or a;
    outputs(11278) <= a xor b;
    outputs(11279) <= a xor b;
    outputs(11280) <= a xor b;
    outputs(11281) <= a xor b;
    outputs(11282) <= not a;
    outputs(11283) <= not (a and b);
    outputs(11284) <= b and not a;
    outputs(11285) <= not a;
    outputs(11286) <= not (a or b);
    outputs(11287) <= b and not a;
    outputs(11288) <= a or b;
    outputs(11289) <= not (a and b);
    outputs(11290) <= a;
    outputs(11291) <= not (a or b);
    outputs(11292) <= a xor b;
    outputs(11293) <= b and not a;
    outputs(11294) <= a xor b;
    outputs(11295) <= a;
    outputs(11296) <= a xor b;
    outputs(11297) <= not a or b;
    outputs(11298) <= a xor b;
    outputs(11299) <= b;
    outputs(11300) <= a xor b;
    outputs(11301) <= not b;
    outputs(11302) <= not b or a;
    outputs(11303) <= b;
    outputs(11304) <= not (a xor b);
    outputs(11305) <= a;
    outputs(11306) <= a;
    outputs(11307) <= not a;
    outputs(11308) <= not b;
    outputs(11309) <= b;
    outputs(11310) <= not (a and b);
    outputs(11311) <= b;
    outputs(11312) <= not a;
    outputs(11313) <= b;
    outputs(11314) <= a xor b;
    outputs(11315) <= not a;
    outputs(11316) <= a;
    outputs(11317) <= a xor b;
    outputs(11318) <= not b;
    outputs(11319) <= a or b;
    outputs(11320) <= b;
    outputs(11321) <= not b or a;
    outputs(11322) <= a;
    outputs(11323) <= b;
    outputs(11324) <= not (a xor b);
    outputs(11325) <= not b;
    outputs(11326) <= not (a xor b);
    outputs(11327) <= a;
    outputs(11328) <= not (a xor b);
    outputs(11329) <= not a;
    outputs(11330) <= not a;
    outputs(11331) <= not a;
    outputs(11332) <= a xor b;
    outputs(11333) <= b;
    outputs(11334) <= b and not a;
    outputs(11335) <= a xor b;
    outputs(11336) <= a or b;
    outputs(11337) <= a xor b;
    outputs(11338) <= a xor b;
    outputs(11339) <= a and b;
    outputs(11340) <= not b or a;
    outputs(11341) <= not (a xor b);
    outputs(11342) <= a xor b;
    outputs(11343) <= b;
    outputs(11344) <= not (a xor b);
    outputs(11345) <= not a or b;
    outputs(11346) <= not (a xor b);
    outputs(11347) <= a and b;
    outputs(11348) <= a;
    outputs(11349) <= not b;
    outputs(11350) <= not (a or b);
    outputs(11351) <= a xor b;
    outputs(11352) <= not a or b;
    outputs(11353) <= not (a or b);
    outputs(11354) <= not (a xor b);
    outputs(11355) <= a xor b;
    outputs(11356) <= a or b;
    outputs(11357) <= not b or a;
    outputs(11358) <= not b or a;
    outputs(11359) <= a xor b;
    outputs(11360) <= b;
    outputs(11361) <= not (a xor b);
    outputs(11362) <= not b;
    outputs(11363) <= not (a xor b);
    outputs(11364) <= a xor b;
    outputs(11365) <= a and b;
    outputs(11366) <= not (a or b);
    outputs(11367) <= not a;
    outputs(11368) <= not b;
    outputs(11369) <= not b;
    outputs(11370) <= not b;
    outputs(11371) <= a and not b;
    outputs(11372) <= a or b;
    outputs(11373) <= a and b;
    outputs(11374) <= a xor b;
    outputs(11375) <= a or b;
    outputs(11376) <= not (a and b);
    outputs(11377) <= b;
    outputs(11378) <= not a or b;
    outputs(11379) <= a or b;
    outputs(11380) <= a xor b;
    outputs(11381) <= a xor b;
    outputs(11382) <= not a;
    outputs(11383) <= not a;
    outputs(11384) <= a;
    outputs(11385) <= a xor b;
    outputs(11386) <= b;
    outputs(11387) <= a;
    outputs(11388) <= not a or b;
    outputs(11389) <= a xor b;
    outputs(11390) <= not (a xor b);
    outputs(11391) <= b;
    outputs(11392) <= a xor b;
    outputs(11393) <= b;
    outputs(11394) <= not b or a;
    outputs(11395) <= not a;
    outputs(11396) <= a or b;
    outputs(11397) <= not (a xor b);
    outputs(11398) <= not a;
    outputs(11399) <= not b;
    outputs(11400) <= not (a or b);
    outputs(11401) <= not (a and b);
    outputs(11402) <= not (a or b);
    outputs(11403) <= not (a xor b);
    outputs(11404) <= a xor b;
    outputs(11405) <= not b;
    outputs(11406) <= b and not a;
    outputs(11407) <= a and not b;
    outputs(11408) <= not a;
    outputs(11409) <= not (a xor b);
    outputs(11410) <= not (a xor b);
    outputs(11411) <= a xor b;
    outputs(11412) <= a xor b;
    outputs(11413) <= not (a xor b);
    outputs(11414) <= not (a xor b);
    outputs(11415) <= not (a and b);
    outputs(11416) <= b;
    outputs(11417) <= a;
    outputs(11418) <= b;
    outputs(11419) <= not (a or b);
    outputs(11420) <= a xor b;
    outputs(11421) <= not b;
    outputs(11422) <= not b or a;
    outputs(11423) <= b;
    outputs(11424) <= b;
    outputs(11425) <= a;
    outputs(11426) <= not b or a;
    outputs(11427) <= a;
    outputs(11428) <= not b;
    outputs(11429) <= not (a or b);
    outputs(11430) <= a;
    outputs(11431) <= not a;
    outputs(11432) <= a or b;
    outputs(11433) <= a or b;
    outputs(11434) <= not a or b;
    outputs(11435) <= b;
    outputs(11436) <= not b;
    outputs(11437) <= a;
    outputs(11438) <= not (a xor b);
    outputs(11439) <= not a or b;
    outputs(11440) <= a or b;
    outputs(11441) <= not (a xor b);
    outputs(11442) <= not (a xor b);
    outputs(11443) <= not a;
    outputs(11444) <= not a;
    outputs(11445) <= not a;
    outputs(11446) <= not a;
    outputs(11447) <= a xor b;
    outputs(11448) <= not (a and b);
    outputs(11449) <= not (a xor b);
    outputs(11450) <= not b;
    outputs(11451) <= b;
    outputs(11452) <= b and not a;
    outputs(11453) <= not (a and b);
    outputs(11454) <= a and b;
    outputs(11455) <= a xor b;
    outputs(11456) <= not a;
    outputs(11457) <= a and b;
    outputs(11458) <= not (a and b);
    outputs(11459) <= not a or b;
    outputs(11460) <= not (a and b);
    outputs(11461) <= a xor b;
    outputs(11462) <= a and not b;
    outputs(11463) <= b and not a;
    outputs(11464) <= a xor b;
    outputs(11465) <= a or b;
    outputs(11466) <= not b or a;
    outputs(11467) <= a xor b;
    outputs(11468) <= not (a or b);
    outputs(11469) <= b and not a;
    outputs(11470) <= not (a xor b);
    outputs(11471) <= a xor b;
    outputs(11472) <= not a;
    outputs(11473) <= b;
    outputs(11474) <= b;
    outputs(11475) <= not b or a;
    outputs(11476) <= not b;
    outputs(11477) <= a xor b;
    outputs(11478) <= not (a xor b);
    outputs(11479) <= a;
    outputs(11480) <= a;
    outputs(11481) <= not (a xor b);
    outputs(11482) <= a xor b;
    outputs(11483) <= a or b;
    outputs(11484) <= a;
    outputs(11485) <= a xor b;
    outputs(11486) <= a and b;
    outputs(11487) <= not (a or b);
    outputs(11488) <= not a;
    outputs(11489) <= not a;
    outputs(11490) <= not (a xor b);
    outputs(11491) <= not a;
    outputs(11492) <= a;
    outputs(11493) <= not (a xor b);
    outputs(11494) <= a and b;
    outputs(11495) <= b;
    outputs(11496) <= not (a xor b);
    outputs(11497) <= a xor b;
    outputs(11498) <= a;
    outputs(11499) <= not (a xor b);
    outputs(11500) <= not (a xor b);
    outputs(11501) <= not a;
    outputs(11502) <= a or b;
    outputs(11503) <= not a;
    outputs(11504) <= not a;
    outputs(11505) <= a or b;
    outputs(11506) <= b;
    outputs(11507) <= b;
    outputs(11508) <= not (a xor b);
    outputs(11509) <= b;
    outputs(11510) <= b;
    outputs(11511) <= not a;
    outputs(11512) <= not a;
    outputs(11513) <= not b or a;
    outputs(11514) <= not (a xor b);
    outputs(11515) <= b;
    outputs(11516) <= not a;
    outputs(11517) <= a xor b;
    outputs(11518) <= not b;
    outputs(11519) <= a or b;
    outputs(11520) <= not b;
    outputs(11521) <= not (a and b);
    outputs(11522) <= a and not b;
    outputs(11523) <= not (a and b);
    outputs(11524) <= a xor b;
    outputs(11525) <= a xor b;
    outputs(11526) <= not a;
    outputs(11527) <= a xor b;
    outputs(11528) <= not a;
    outputs(11529) <= a;
    outputs(11530) <= a xor b;
    outputs(11531) <= a and b;
    outputs(11532) <= not b;
    outputs(11533) <= not (a or b);
    outputs(11534) <= not (a xor b);
    outputs(11535) <= not b;
    outputs(11536) <= a xor b;
    outputs(11537) <= not a;
    outputs(11538) <= b;
    outputs(11539) <= not a;
    outputs(11540) <= not a or b;
    outputs(11541) <= not a;
    outputs(11542) <= b and not a;
    outputs(11543) <= not (a or b);
    outputs(11544) <= not b or a;
    outputs(11545) <= not a or b;
    outputs(11546) <= a xor b;
    outputs(11547) <= a;
    outputs(11548) <= not b;
    outputs(11549) <= a and b;
    outputs(11550) <= not (a xor b);
    outputs(11551) <= not (a xor b);
    outputs(11552) <= not b;
    outputs(11553) <= b;
    outputs(11554) <= not a;
    outputs(11555) <= a and b;
    outputs(11556) <= not b;
    outputs(11557) <= not b;
    outputs(11558) <= not a;
    outputs(11559) <= b;
    outputs(11560) <= a and not b;
    outputs(11561) <= b;
    outputs(11562) <= not b;
    outputs(11563) <= a and b;
    outputs(11564) <= b;
    outputs(11565) <= a or b;
    outputs(11566) <= a;
    outputs(11567) <= not a;
    outputs(11568) <= a and not b;
    outputs(11569) <= not a;
    outputs(11570) <= b and not a;
    outputs(11571) <= a xor b;
    outputs(11572) <= not a;
    outputs(11573) <= not b;
    outputs(11574) <= a and not b;
    outputs(11575) <= not a;
    outputs(11576) <= a;
    outputs(11577) <= not b;
    outputs(11578) <= not b;
    outputs(11579) <= b;
    outputs(11580) <= not (a xor b);
    outputs(11581) <= a;
    outputs(11582) <= a xor b;
    outputs(11583) <= a xor b;
    outputs(11584) <= a;
    outputs(11585) <= b;
    outputs(11586) <= b;
    outputs(11587) <= not b;
    outputs(11588) <= not b or a;
    outputs(11589) <= not (a xor b);
    outputs(11590) <= a xor b;
    outputs(11591) <= not (a xor b);
    outputs(11592) <= a xor b;
    outputs(11593) <= a and b;
    outputs(11594) <= a and not b;
    outputs(11595) <= not (a or b);
    outputs(11596) <= not a;
    outputs(11597) <= b;
    outputs(11598) <= not (a xor b);
    outputs(11599) <= b;
    outputs(11600) <= not b;
    outputs(11601) <= not b;
    outputs(11602) <= a;
    outputs(11603) <= not (a xor b);
    outputs(11604) <= a xor b;
    outputs(11605) <= not (a xor b);
    outputs(11606) <= not b;
    outputs(11607) <= not (a xor b);
    outputs(11608) <= not a or b;
    outputs(11609) <= a and not b;
    outputs(11610) <= b and not a;
    outputs(11611) <= not (a xor b);
    outputs(11612) <= b;
    outputs(11613) <= b;
    outputs(11614) <= a and b;
    outputs(11615) <= not (a xor b);
    outputs(11616) <= a xor b;
    outputs(11617) <= a xor b;
    outputs(11618) <= not a or b;
    outputs(11619) <= not a;
    outputs(11620) <= not (a xor b);
    outputs(11621) <= not a or b;
    outputs(11622) <= a;
    outputs(11623) <= a xor b;
    outputs(11624) <= not b or a;
    outputs(11625) <= a and b;
    outputs(11626) <= b;
    outputs(11627) <= not a;
    outputs(11628) <= b;
    outputs(11629) <= a;
    outputs(11630) <= a;
    outputs(11631) <= not (a xor b);
    outputs(11632) <= a and not b;
    outputs(11633) <= not b;
    outputs(11634) <= not b;
    outputs(11635) <= a;
    outputs(11636) <= a;
    outputs(11637) <= a xor b;
    outputs(11638) <= a and b;
    outputs(11639) <= a and not b;
    outputs(11640) <= not (a xor b);
    outputs(11641) <= not b;
    outputs(11642) <= not (a xor b);
    outputs(11643) <= not b;
    outputs(11644) <= b and not a;
    outputs(11645) <= b;
    outputs(11646) <= not (a or b);
    outputs(11647) <= not b;
    outputs(11648) <= not b;
    outputs(11649) <= not a;
    outputs(11650) <= not b or a;
    outputs(11651) <= not b;
    outputs(11652) <= not b;
    outputs(11653) <= b;
    outputs(11654) <= a xor b;
    outputs(11655) <= a xor b;
    outputs(11656) <= not (a xor b);
    outputs(11657) <= b;
    outputs(11658) <= b and not a;
    outputs(11659) <= not (a or b);
    outputs(11660) <= b;
    outputs(11661) <= a xor b;
    outputs(11662) <= a xor b;
    outputs(11663) <= a or b;
    outputs(11664) <= a and b;
    outputs(11665) <= not a;
    outputs(11666) <= a xor b;
    outputs(11667) <= a xor b;
    outputs(11668) <= not (a or b);
    outputs(11669) <= a or b;
    outputs(11670) <= a;
    outputs(11671) <= not b;
    outputs(11672) <= a xor b;
    outputs(11673) <= not (a xor b);
    outputs(11674) <= a xor b;
    outputs(11675) <= a;
    outputs(11676) <= not b;
    outputs(11677) <= not a;
    outputs(11678) <= not (a xor b);
    outputs(11679) <= a;
    outputs(11680) <= a xor b;
    outputs(11681) <= a xor b;
    outputs(11682) <= not (a and b);
    outputs(11683) <= b and not a;
    outputs(11684) <= not a;
    outputs(11685) <= not (a xor b);
    outputs(11686) <= a and not b;
    outputs(11687) <= b and not a;
    outputs(11688) <= not (a xor b);
    outputs(11689) <= not b;
    outputs(11690) <= not a;
    outputs(11691) <= a xor b;
    outputs(11692) <= a xor b;
    outputs(11693) <= not (a and b);
    outputs(11694) <= not (a or b);
    outputs(11695) <= a xor b;
    outputs(11696) <= a xor b;
    outputs(11697) <= not (a xor b);
    outputs(11698) <= not (a or b);
    outputs(11699) <= not a;
    outputs(11700) <= not a;
    outputs(11701) <= not b or a;
    outputs(11702) <= a;
    outputs(11703) <= not (a xor b);
    outputs(11704) <= not b or a;
    outputs(11705) <= b and not a;
    outputs(11706) <= a;
    outputs(11707) <= b;
    outputs(11708) <= not a;
    outputs(11709) <= a xor b;
    outputs(11710) <= not (a or b);
    outputs(11711) <= b;
    outputs(11712) <= not (a xor b);
    outputs(11713) <= a;
    outputs(11714) <= a xor b;
    outputs(11715) <= not a;
    outputs(11716) <= not a or b;
    outputs(11717) <= not (a xor b);
    outputs(11718) <= not (a xor b);
    outputs(11719) <= a;
    outputs(11720) <= not a;
    outputs(11721) <= not a;
    outputs(11722) <= b;
    outputs(11723) <= not (a xor b);
    outputs(11724) <= b;
    outputs(11725) <= not (a or b);
    outputs(11726) <= a;
    outputs(11727) <= not (a xor b);
    outputs(11728) <= b;
    outputs(11729) <= not (a xor b);
    outputs(11730) <= not (a xor b);
    outputs(11731) <= not (a xor b);
    outputs(11732) <= not b;
    outputs(11733) <= a;
    outputs(11734) <= a xor b;
    outputs(11735) <= not (a xor b);
    outputs(11736) <= not b;
    outputs(11737) <= a or b;
    outputs(11738) <= b;
    outputs(11739) <= b and not a;
    outputs(11740) <= a and b;
    outputs(11741) <= a xor b;
    outputs(11742) <= b;
    outputs(11743) <= not b;
    outputs(11744) <= b;
    outputs(11745) <= not a;
    outputs(11746) <= a xor b;
    outputs(11747) <= b and not a;
    outputs(11748) <= a;
    outputs(11749) <= b;
    outputs(11750) <= a xor b;
    outputs(11751) <= not (a xor b);
    outputs(11752) <= a xor b;
    outputs(11753) <= not a;
    outputs(11754) <= not b;
    outputs(11755) <= not (a xor b);
    outputs(11756) <= not a;
    outputs(11757) <= not (a xor b);
    outputs(11758) <= not (a xor b);
    outputs(11759) <= a;
    outputs(11760) <= not b;
    outputs(11761) <= a and b;
    outputs(11762) <= not (a xor b);
    outputs(11763) <= b;
    outputs(11764) <= not a;
    outputs(11765) <= not (a or b);
    outputs(11766) <= a;
    outputs(11767) <= not a;
    outputs(11768) <= a xor b;
    outputs(11769) <= not (a xor b);
    outputs(11770) <= not b or a;
    outputs(11771) <= not b;
    outputs(11772) <= not b;
    outputs(11773) <= a and b;
    outputs(11774) <= not b or a;
    outputs(11775) <= not (a xor b);
    outputs(11776) <= a xor b;
    outputs(11777) <= b;
    outputs(11778) <= not (a xor b);
    outputs(11779) <= not a or b;
    outputs(11780) <= a xor b;
    outputs(11781) <= not b or a;
    outputs(11782) <= a and not b;
    outputs(11783) <= not (a xor b);
    outputs(11784) <= not (a xor b);
    outputs(11785) <= not b or a;
    outputs(11786) <= not b;
    outputs(11787) <= a;
    outputs(11788) <= b;
    outputs(11789) <= not a;
    outputs(11790) <= not (a xor b);
    outputs(11791) <= a xor b;
    outputs(11792) <= not (a xor b);
    outputs(11793) <= not a;
    outputs(11794) <= a xor b;
    outputs(11795) <= a;
    outputs(11796) <= not b;
    outputs(11797) <= not (a or b);
    outputs(11798) <= not (a and b);
    outputs(11799) <= a;
    outputs(11800) <= not b;
    outputs(11801) <= b;
    outputs(11802) <= a;
    outputs(11803) <= a xor b;
    outputs(11804) <= not b;
    outputs(11805) <= a and not b;
    outputs(11806) <= b and not a;
    outputs(11807) <= b;
    outputs(11808) <= a;
    outputs(11809) <= not (a xor b);
    outputs(11810) <= not (a xor b);
    outputs(11811) <= not (a and b);
    outputs(11812) <= b and not a;
    outputs(11813) <= not b;
    outputs(11814) <= not (a xor b);
    outputs(11815) <= not (a and b);
    outputs(11816) <= a xor b;
    outputs(11817) <= not a;
    outputs(11818) <= not (a or b);
    outputs(11819) <= a;
    outputs(11820) <= a and not b;
    outputs(11821) <= a xor b;
    outputs(11822) <= b and not a;
    outputs(11823) <= a and b;
    outputs(11824) <= a xor b;
    outputs(11825) <= not a;
    outputs(11826) <= a and not b;
    outputs(11827) <= a xor b;
    outputs(11828) <= not (a xor b);
    outputs(11829) <= a xor b;
    outputs(11830) <= b and not a;
    outputs(11831) <= a xor b;
    outputs(11832) <= not a;
    outputs(11833) <= a xor b;
    outputs(11834) <= not (a xor b);
    outputs(11835) <= not (a xor b);
    outputs(11836) <= a and not b;
    outputs(11837) <= a;
    outputs(11838) <= a xor b;
    outputs(11839) <= a and b;
    outputs(11840) <= not a;
    outputs(11841) <= b;
    outputs(11842) <= b;
    outputs(11843) <= not a;
    outputs(11844) <= a or b;
    outputs(11845) <= a;
    outputs(11846) <= a or b;
    outputs(11847) <= not (a xor b);
    outputs(11848) <= not a;
    outputs(11849) <= not b;
    outputs(11850) <= a xor b;
    outputs(11851) <= not a;
    outputs(11852) <= a xor b;
    outputs(11853) <= not (a xor b);
    outputs(11854) <= not (a or b);
    outputs(11855) <= not b;
    outputs(11856) <= a;
    outputs(11857) <= not (a xor b);
    outputs(11858) <= not (a xor b);
    outputs(11859) <= b;
    outputs(11860) <= a;
    outputs(11861) <= a xor b;
    outputs(11862) <= not (a xor b);
    outputs(11863) <= not (a xor b);
    outputs(11864) <= not (a xor b);
    outputs(11865) <= a xor b;
    outputs(11866) <= not (a xor b);
    outputs(11867) <= a and b;
    outputs(11868) <= not a;
    outputs(11869) <= a and not b;
    outputs(11870) <= a xor b;
    outputs(11871) <= a and b;
    outputs(11872) <= b;
    outputs(11873) <= a and not b;
    outputs(11874) <= a;
    outputs(11875) <= b;
    outputs(11876) <= not b;
    outputs(11877) <= not (a xor b);
    outputs(11878) <= not a;
    outputs(11879) <= a xor b;
    outputs(11880) <= not (a and b);
    outputs(11881) <= a xor b;
    outputs(11882) <= b and not a;
    outputs(11883) <= a xor b;
    outputs(11884) <= not (a xor b);
    outputs(11885) <= a xor b;
    outputs(11886) <= b and not a;
    outputs(11887) <= a xor b;
    outputs(11888) <= not b;
    outputs(11889) <= not b;
    outputs(11890) <= not a or b;
    outputs(11891) <= not a;
    outputs(11892) <= not a;
    outputs(11893) <= not (a and b);
    outputs(11894) <= a or b;
    outputs(11895) <= not (a xor b);
    outputs(11896) <= a;
    outputs(11897) <= b;
    outputs(11898) <= not a;
    outputs(11899) <= not a;
    outputs(11900) <= a;
    outputs(11901) <= not (a xor b);
    outputs(11902) <= not (a xor b);
    outputs(11903) <= not b;
    outputs(11904) <= a;
    outputs(11905) <= a xor b;
    outputs(11906) <= b and not a;
    outputs(11907) <= not (a and b);
    outputs(11908) <= not (a xor b);
    outputs(11909) <= b;
    outputs(11910) <= not b or a;
    outputs(11911) <= a xor b;
    outputs(11912) <= not (a xor b);
    outputs(11913) <= a xor b;
    outputs(11914) <= b;
    outputs(11915) <= not a;
    outputs(11916) <= not (a xor b);
    outputs(11917) <= not b or a;
    outputs(11918) <= a xor b;
    outputs(11919) <= not b;
    outputs(11920) <= a and not b;
    outputs(11921) <= not (a xor b);
    outputs(11922) <= not (a xor b);
    outputs(11923) <= not b;
    outputs(11924) <= not (a xor b);
    outputs(11925) <= not a;
    outputs(11926) <= a or b;
    outputs(11927) <= not (a xor b);
    outputs(11928) <= a and not b;
    outputs(11929) <= a xor b;
    outputs(11930) <= not a;
    outputs(11931) <= not a;
    outputs(11932) <= not (a xor b);
    outputs(11933) <= a and b;
    outputs(11934) <= a xor b;
    outputs(11935) <= a and not b;
    outputs(11936) <= a xor b;
    outputs(11937) <= a xor b;
    outputs(11938) <= a and b;
    outputs(11939) <= a xor b;
    outputs(11940) <= not a;
    outputs(11941) <= not a;
    outputs(11942) <= a and b;
    outputs(11943) <= a;
    outputs(11944) <= a;
    outputs(11945) <= not (a or b);
    outputs(11946) <= a;
    outputs(11947) <= a xor b;
    outputs(11948) <= a and not b;
    outputs(11949) <= a;
    outputs(11950) <= a xor b;
    outputs(11951) <= b;
    outputs(11952) <= not (a xor b);
    outputs(11953) <= not (a xor b);
    outputs(11954) <= not a or b;
    outputs(11955) <= not a;
    outputs(11956) <= a;
    outputs(11957) <= a;
    outputs(11958) <= not (a or b);
    outputs(11959) <= a and not b;
    outputs(11960) <= not (a xor b);
    outputs(11961) <= a xor b;
    outputs(11962) <= a;
    outputs(11963) <= not a;
    outputs(11964) <= not (a or b);
    outputs(11965) <= not (a or b);
    outputs(11966) <= not (a xor b);
    outputs(11967) <= not (a xor b);
    outputs(11968) <= b and not a;
    outputs(11969) <= b;
    outputs(11970) <= a or b;
    outputs(11971) <= not (a xor b);
    outputs(11972) <= not (a xor b);
    outputs(11973) <= not a;
    outputs(11974) <= a;
    outputs(11975) <= not (a xor b);
    outputs(11976) <= b;
    outputs(11977) <= not (a xor b);
    outputs(11978) <= not (a xor b);
    outputs(11979) <= not b;
    outputs(11980) <= a and b;
    outputs(11981) <= a;
    outputs(11982) <= not (a xor b);
    outputs(11983) <= b and not a;
    outputs(11984) <= not (a xor b);
    outputs(11985) <= not (a xor b);
    outputs(11986) <= b;
    outputs(11987) <= not (a xor b);
    outputs(11988) <= not b;
    outputs(11989) <= a;
    outputs(11990) <= a or b;
    outputs(11991) <= not b;
    outputs(11992) <= a or b;
    outputs(11993) <= a;
    outputs(11994) <= a;
    outputs(11995) <= a;
    outputs(11996) <= not (a xor b);
    outputs(11997) <= not b;
    outputs(11998) <= a xor b;
    outputs(11999) <= not (a xor b);
    outputs(12000) <= not (a xor b);
    outputs(12001) <= a xor b;
    outputs(12002) <= a and not b;
    outputs(12003) <= a xor b;
    outputs(12004) <= a xor b;
    outputs(12005) <= not b;
    outputs(12006) <= not a;
    outputs(12007) <= a xor b;
    outputs(12008) <= not (a xor b);
    outputs(12009) <= not b;
    outputs(12010) <= a xor b;
    outputs(12011) <= a xor b;
    outputs(12012) <= a xor b;
    outputs(12013) <= a and not b;
    outputs(12014) <= b;
    outputs(12015) <= b;
    outputs(12016) <= a;
    outputs(12017) <= a and b;
    outputs(12018) <= b;
    outputs(12019) <= not b;
    outputs(12020) <= a and b;
    outputs(12021) <= not (a xor b);
    outputs(12022) <= a xor b;
    outputs(12023) <= a and not b;
    outputs(12024) <= a;
    outputs(12025) <= not b;
    outputs(12026) <= not b;
    outputs(12027) <= a xor b;
    outputs(12028) <= b;
    outputs(12029) <= not (a and b);
    outputs(12030) <= not (a xor b);
    outputs(12031) <= not (a xor b);
    outputs(12032) <= not a or b;
    outputs(12033) <= not b;
    outputs(12034) <= not b;
    outputs(12035) <= not (a and b);
    outputs(12036) <= b;
    outputs(12037) <= not b or a;
    outputs(12038) <= b and not a;
    outputs(12039) <= a and b;
    outputs(12040) <= b and not a;
    outputs(12041) <= not a;
    outputs(12042) <= not a;
    outputs(12043) <= a xor b;
    outputs(12044) <= a xor b;
    outputs(12045) <= not a;
    outputs(12046) <= b;
    outputs(12047) <= b;
    outputs(12048) <= not a;
    outputs(12049) <= a xor b;
    outputs(12050) <= a or b;
    outputs(12051) <= not a;
    outputs(12052) <= not (a xor b);
    outputs(12053) <= a;
    outputs(12054) <= not (a xor b);
    outputs(12055) <= a;
    outputs(12056) <= a;
    outputs(12057) <= a;
    outputs(12058) <= a;
    outputs(12059) <= a or b;
    outputs(12060) <= not a;
    outputs(12061) <= not a;
    outputs(12062) <= not a;
    outputs(12063) <= b;
    outputs(12064) <= not a;
    outputs(12065) <= not b;
    outputs(12066) <= b;
    outputs(12067) <= not (a or b);
    outputs(12068) <= a and not b;
    outputs(12069) <= a;
    outputs(12070) <= not (a xor b);
    outputs(12071) <= a and b;
    outputs(12072) <= not a;
    outputs(12073) <= not b or a;
    outputs(12074) <= a xor b;
    outputs(12075) <= not b;
    outputs(12076) <= not a;
    outputs(12077) <= b and not a;
    outputs(12078) <= b;
    outputs(12079) <= a xor b;
    outputs(12080) <= not (a xor b);
    outputs(12081) <= not (a xor b);
    outputs(12082) <= not a;
    outputs(12083) <= not b;
    outputs(12084) <= not (a xor b);
    outputs(12085) <= not b;
    outputs(12086) <= not b;
    outputs(12087) <= not a;
    outputs(12088) <= not a;
    outputs(12089) <= not b or a;
    outputs(12090) <= b;
    outputs(12091) <= not (a xor b);
    outputs(12092) <= not (a or b);
    outputs(12093) <= not b;
    outputs(12094) <= not b;
    outputs(12095) <= not b;
    outputs(12096) <= not (a xor b);
    outputs(12097) <= a;
    outputs(12098) <= not (a and b);
    outputs(12099) <= b;
    outputs(12100) <= b and not a;
    outputs(12101) <= not b;
    outputs(12102) <= not (a and b);
    outputs(12103) <= not b;
    outputs(12104) <= a xor b;
    outputs(12105) <= a;
    outputs(12106) <= a and not b;
    outputs(12107) <= a xor b;
    outputs(12108) <= not a;
    outputs(12109) <= not b;
    outputs(12110) <= a xor b;
    outputs(12111) <= a xor b;
    outputs(12112) <= not b or a;
    outputs(12113) <= not b;
    outputs(12114) <= not a;
    outputs(12115) <= not (a xor b);
    outputs(12116) <= a and b;
    outputs(12117) <= not a;
    outputs(12118) <= b;
    outputs(12119) <= a and b;
    outputs(12120) <= a xor b;
    outputs(12121) <= a;
    outputs(12122) <= a xor b;
    outputs(12123) <= a;
    outputs(12124) <= not (a or b);
    outputs(12125) <= not (a or b);
    outputs(12126) <= not b;
    outputs(12127) <= a and b;
    outputs(12128) <= a xor b;
    outputs(12129) <= not (a xor b);
    outputs(12130) <= not (a xor b);
    outputs(12131) <= not b;
    outputs(12132) <= b and not a;
    outputs(12133) <= not b;
    outputs(12134) <= not b;
    outputs(12135) <= not (a xor b);
    outputs(12136) <= a xor b;
    outputs(12137) <= b and not a;
    outputs(12138) <= a xor b;
    outputs(12139) <= a;
    outputs(12140) <= a;
    outputs(12141) <= not (a xor b);
    outputs(12142) <= a or b;
    outputs(12143) <= not (a xor b);
    outputs(12144) <= not (a and b);
    outputs(12145) <= not b or a;
    outputs(12146) <= not (a or b);
    outputs(12147) <= a xor b;
    outputs(12148) <= a xor b;
    outputs(12149) <= a xor b;
    outputs(12150) <= not a;
    outputs(12151) <= a and b;
    outputs(12152) <= b and not a;
    outputs(12153) <= a;
    outputs(12154) <= not (a xor b);
    outputs(12155) <= b;
    outputs(12156) <= not (a xor b);
    outputs(12157) <= b;
    outputs(12158) <= a and b;
    outputs(12159) <= a or b;
    outputs(12160) <= a and not b;
    outputs(12161) <= a;
    outputs(12162) <= not (a xor b);
    outputs(12163) <= not a;
    outputs(12164) <= a;
    outputs(12165) <= not b;
    outputs(12166) <= a or b;
    outputs(12167) <= not a or b;
    outputs(12168) <= b and not a;
    outputs(12169) <= a and not b;
    outputs(12170) <= not (a xor b);
    outputs(12171) <= a and b;
    outputs(12172) <= a xor b;
    outputs(12173) <= b;
    outputs(12174) <= not a or b;
    outputs(12175) <= a xor b;
    outputs(12176) <= not b;
    outputs(12177) <= b;
    outputs(12178) <= a;
    outputs(12179) <= not b or a;
    outputs(12180) <= not a;
    outputs(12181) <= a;
    outputs(12182) <= not (a xor b);
    outputs(12183) <= a and b;
    outputs(12184) <= a and not b;
    outputs(12185) <= not (a xor b);
    outputs(12186) <= not b;
    outputs(12187) <= b;
    outputs(12188) <= a;
    outputs(12189) <= not (a xor b);
    outputs(12190) <= b;
    outputs(12191) <= b;
    outputs(12192) <= not (a xor b);
    outputs(12193) <= b;
    outputs(12194) <= a;
    outputs(12195) <= not (a xor b);
    outputs(12196) <= a xor b;
    outputs(12197) <= b;
    outputs(12198) <= b and not a;
    outputs(12199) <= a xor b;
    outputs(12200) <= a xor b;
    outputs(12201) <= not a;
    outputs(12202) <= a xor b;
    outputs(12203) <= not (a xor b);
    outputs(12204) <= a xor b;
    outputs(12205) <= b;
    outputs(12206) <= not b;
    outputs(12207) <= not a or b;
    outputs(12208) <= not (a or b);
    outputs(12209) <= a xor b;
    outputs(12210) <= a;
    outputs(12211) <= a and not b;
    outputs(12212) <= a and b;
    outputs(12213) <= a xor b;
    outputs(12214) <= a and not b;
    outputs(12215) <= a xor b;
    outputs(12216) <= not a;
    outputs(12217) <= not a;
    outputs(12218) <= not b;
    outputs(12219) <= a xor b;
    outputs(12220) <= b;
    outputs(12221) <= not a;
    outputs(12222) <= a xor b;
    outputs(12223) <= not b;
    outputs(12224) <= not (a xor b);
    outputs(12225) <= a and not b;
    outputs(12226) <= not b;
    outputs(12227) <= not (a or b);
    outputs(12228) <= a;
    outputs(12229) <= b;
    outputs(12230) <= not b or a;
    outputs(12231) <= b;
    outputs(12232) <= not (a xor b);
    outputs(12233) <= not (a xor b);
    outputs(12234) <= b;
    outputs(12235) <= not a;
    outputs(12236) <= not (a xor b);
    outputs(12237) <= a xor b;
    outputs(12238) <= b and not a;
    outputs(12239) <= a or b;
    outputs(12240) <= a xor b;
    outputs(12241) <= a and not b;
    outputs(12242) <= a xor b;
    outputs(12243) <= not (a xor b);
    outputs(12244) <= a xor b;
    outputs(12245) <= not a;
    outputs(12246) <= not (a xor b);
    outputs(12247) <= not a;
    outputs(12248) <= a xor b;
    outputs(12249) <= a xor b;
    outputs(12250) <= a xor b;
    outputs(12251) <= b;
    outputs(12252) <= not b;
    outputs(12253) <= b and not a;
    outputs(12254) <= '1';
    outputs(12255) <= not a;
    outputs(12256) <= not b;
    outputs(12257) <= not (a xor b);
    outputs(12258) <= a;
    outputs(12259) <= a and b;
    outputs(12260) <= not a;
    outputs(12261) <= a xor b;
    outputs(12262) <= not a;
    outputs(12263) <= b and not a;
    outputs(12264) <= not b;
    outputs(12265) <= not (a xor b);
    outputs(12266) <= not b or a;
    outputs(12267) <= a and not b;
    outputs(12268) <= b;
    outputs(12269) <= a xor b;
    outputs(12270) <= not b;
    outputs(12271) <= not (a xor b);
    outputs(12272) <= not b;
    outputs(12273) <= not (a xor b);
    outputs(12274) <= not a;
    outputs(12275) <= not b;
    outputs(12276) <= not (a xor b);
    outputs(12277) <= not b;
    outputs(12278) <= a and b;
    outputs(12279) <= a;
    outputs(12280) <= not (a xor b);
    outputs(12281) <= a;
    outputs(12282) <= a xor b;
    outputs(12283) <= a xor b;
    outputs(12284) <= a or b;
    outputs(12285) <= b;
    outputs(12286) <= b;
    outputs(12287) <= a xor b;
    outputs(12288) <= b;
    outputs(12289) <= a xor b;
    outputs(12290) <= not b;
    outputs(12291) <= not (a and b);
    outputs(12292) <= a;
    outputs(12293) <= not (a xor b);
    outputs(12294) <= a;
    outputs(12295) <= a;
    outputs(12296) <= not (a xor b);
    outputs(12297) <= not (a xor b);
    outputs(12298) <= a;
    outputs(12299) <= not a;
    outputs(12300) <= not (a xor b);
    outputs(12301) <= a xor b;
    outputs(12302) <= not (a xor b);
    outputs(12303) <= not a;
    outputs(12304) <= not a;
    outputs(12305) <= a xor b;
    outputs(12306) <= not (a xor b);
    outputs(12307) <= b;
    outputs(12308) <= a and not b;
    outputs(12309) <= not a;
    outputs(12310) <= not b;
    outputs(12311) <= a or b;
    outputs(12312) <= b and not a;
    outputs(12313) <= b;
    outputs(12314) <= b;
    outputs(12315) <= a and b;
    outputs(12316) <= not b;
    outputs(12317) <= a;
    outputs(12318) <= not (a xor b);
    outputs(12319) <= b;
    outputs(12320) <= b and not a;
    outputs(12321) <= a;
    outputs(12322) <= b;
    outputs(12323) <= a;
    outputs(12324) <= a or b;
    outputs(12325) <= not a or b;
    outputs(12326) <= a and b;
    outputs(12327) <= not a or b;
    outputs(12328) <= not a;
    outputs(12329) <= not (a xor b);
    outputs(12330) <= not a or b;
    outputs(12331) <= not b;
    outputs(12332) <= a xor b;
    outputs(12333) <= not (a xor b);
    outputs(12334) <= not a;
    outputs(12335) <= a xor b;
    outputs(12336) <= a;
    outputs(12337) <= a and b;
    outputs(12338) <= not (a or b);
    outputs(12339) <= a and not b;
    outputs(12340) <= a;
    outputs(12341) <= a and b;
    outputs(12342) <= b and not a;
    outputs(12343) <= not (a xor b);
    outputs(12344) <= not a or b;
    outputs(12345) <= b;
    outputs(12346) <= a and not b;
    outputs(12347) <= not (a or b);
    outputs(12348) <= not b;
    outputs(12349) <= b;
    outputs(12350) <= b;
    outputs(12351) <= not b;
    outputs(12352) <= not b;
    outputs(12353) <= not b;
    outputs(12354) <= a xor b;
    outputs(12355) <= not a;
    outputs(12356) <= not a;
    outputs(12357) <= not (a xor b);
    outputs(12358) <= not b;
    outputs(12359) <= a and b;
    outputs(12360) <= not a;
    outputs(12361) <= a and b;
    outputs(12362) <= not a;
    outputs(12363) <= a and b;
    outputs(12364) <= a and not b;
    outputs(12365) <= a xor b;
    outputs(12366) <= a and b;
    outputs(12367) <= not b;
    outputs(12368) <= not (a xor b);
    outputs(12369) <= not b;
    outputs(12370) <= a;
    outputs(12371) <= a xor b;
    outputs(12372) <= a and not b;
    outputs(12373) <= b;
    outputs(12374) <= b;
    outputs(12375) <= not (a xor b);
    outputs(12376) <= not (a or b);
    outputs(12377) <= not b;
    outputs(12378) <= a xor b;
    outputs(12379) <= a xor b;
    outputs(12380) <= not a;
    outputs(12381) <= not (a or b);
    outputs(12382) <= b and not a;
    outputs(12383) <= a and not b;
    outputs(12384) <= b;
    outputs(12385) <= a xor b;
    outputs(12386) <= a xor b;
    outputs(12387) <= b and not a;
    outputs(12388) <= a or b;
    outputs(12389) <= not (a xor b);
    outputs(12390) <= a or b;
    outputs(12391) <= not (a xor b);
    outputs(12392) <= a xor b;
    outputs(12393) <= b;
    outputs(12394) <= not (a and b);
    outputs(12395) <= not (a xor b);
    outputs(12396) <= b;
    outputs(12397) <= a and b;
    outputs(12398) <= b and not a;
    outputs(12399) <= not a or b;
    outputs(12400) <= not (a xor b);
    outputs(12401) <= b;
    outputs(12402) <= a xor b;
    outputs(12403) <= not a or b;
    outputs(12404) <= not a;
    outputs(12405) <= a xor b;
    outputs(12406) <= a or b;
    outputs(12407) <= a xor b;
    outputs(12408) <= b;
    outputs(12409) <= a xor b;
    outputs(12410) <= a xor b;
    outputs(12411) <= not (a xor b);
    outputs(12412) <= a and not b;
    outputs(12413) <= not (a xor b);
    outputs(12414) <= not (a xor b);
    outputs(12415) <= a xor b;
    outputs(12416) <= not (a or b);
    outputs(12417) <= not b or a;
    outputs(12418) <= a and not b;
    outputs(12419) <= not (a and b);
    outputs(12420) <= a xor b;
    outputs(12421) <= not b;
    outputs(12422) <= not a;
    outputs(12423) <= not b;
    outputs(12424) <= a xor b;
    outputs(12425) <= not a or b;
    outputs(12426) <= b and not a;
    outputs(12427) <= not a;
    outputs(12428) <= not b;
    outputs(12429) <= not (a xor b);
    outputs(12430) <= not (a xor b);
    outputs(12431) <= b;
    outputs(12432) <= not a;
    outputs(12433) <= a xor b;
    outputs(12434) <= a xor b;
    outputs(12435) <= a or b;
    outputs(12436) <= a;
    outputs(12437) <= a;
    outputs(12438) <= not b;
    outputs(12439) <= not b;
    outputs(12440) <= a and not b;
    outputs(12441) <= a or b;
    outputs(12442) <= a xor b;
    outputs(12443) <= a and b;
    outputs(12444) <= not (a xor b);
    outputs(12445) <= a;
    outputs(12446) <= not (a xor b);
    outputs(12447) <= a;
    outputs(12448) <= a;
    outputs(12449) <= a xor b;
    outputs(12450) <= b;
    outputs(12451) <= a xor b;
    outputs(12452) <= a xor b;
    outputs(12453) <= not (a or b);
    outputs(12454) <= a;
    outputs(12455) <= a xor b;
    outputs(12456) <= not (a xor b);
    outputs(12457) <= not (a xor b);
    outputs(12458) <= not (a xor b);
    outputs(12459) <= not (a xor b);
    outputs(12460) <= not b;
    outputs(12461) <= not a;
    outputs(12462) <= a xor b;
    outputs(12463) <= not b;
    outputs(12464) <= not a;
    outputs(12465) <= a xor b;
    outputs(12466) <= a and not b;
    outputs(12467) <= not (a or b);
    outputs(12468) <= a xor b;
    outputs(12469) <= not (a xor b);
    outputs(12470) <= a xor b;
    outputs(12471) <= not a;
    outputs(12472) <= b;
    outputs(12473) <= a xor b;
    outputs(12474) <= b;
    outputs(12475) <= b;
    outputs(12476) <= not (a xor b);
    outputs(12477) <= not (a xor b);
    outputs(12478) <= a;
    outputs(12479) <= a and b;
    outputs(12480) <= not a;
    outputs(12481) <= a and b;
    outputs(12482) <= not b;
    outputs(12483) <= b;
    outputs(12484) <= not b;
    outputs(12485) <= not b;
    outputs(12486) <= not b;
    outputs(12487) <= not (a or b);
    outputs(12488) <= a xor b;
    outputs(12489) <= not a;
    outputs(12490) <= a xor b;
    outputs(12491) <= a and not b;
    outputs(12492) <= b;
    outputs(12493) <= not (a xor b);
    outputs(12494) <= a xor b;
    outputs(12495) <= a xor b;
    outputs(12496) <= a;
    outputs(12497) <= not a or b;
    outputs(12498) <= a and not b;
    outputs(12499) <= a and b;
    outputs(12500) <= b;
    outputs(12501) <= b and not a;
    outputs(12502) <= a;
    outputs(12503) <= a xor b;
    outputs(12504) <= a xor b;
    outputs(12505) <= not (a xor b);
    outputs(12506) <= b;
    outputs(12507) <= a;
    outputs(12508) <= b;
    outputs(12509) <= b;
    outputs(12510) <= a;
    outputs(12511) <= not (a xor b);
    outputs(12512) <= not a or b;
    outputs(12513) <= a xor b;
    outputs(12514) <= not a;
    outputs(12515) <= a xor b;
    outputs(12516) <= not (a and b);
    outputs(12517) <= a xor b;
    outputs(12518) <= not b;
    outputs(12519) <= not b;
    outputs(12520) <= a or b;
    outputs(12521) <= not (a xor b);
    outputs(12522) <= a xor b;
    outputs(12523) <= a or b;
    outputs(12524) <= not (a xor b);
    outputs(12525) <= a xor b;
    outputs(12526) <= not a;
    outputs(12527) <= a and b;
    outputs(12528) <= not a;
    outputs(12529) <= a xor b;
    outputs(12530) <= b;
    outputs(12531) <= not b;
    outputs(12532) <= not b;
    outputs(12533) <= a and b;
    outputs(12534) <= not b;
    outputs(12535) <= not (a xor b);
    outputs(12536) <= not (a xor b);
    outputs(12537) <= not (a xor b);
    outputs(12538) <= not (a xor b);
    outputs(12539) <= a and not b;
    outputs(12540) <= a;
    outputs(12541) <= not (a xor b);
    outputs(12542) <= not b;
    outputs(12543) <= not (a and b);
    outputs(12544) <= a xor b;
    outputs(12545) <= not (a xor b);
    outputs(12546) <= not (a xor b);
    outputs(12547) <= a xor b;
    outputs(12548) <= a and not b;
    outputs(12549) <= b;
    outputs(12550) <= not (a or b);
    outputs(12551) <= a and b;
    outputs(12552) <= a and b;
    outputs(12553) <= a xor b;
    outputs(12554) <= not b;
    outputs(12555) <= a and b;
    outputs(12556) <= not b or a;
    outputs(12557) <= b;
    outputs(12558) <= a;
    outputs(12559) <= not (a xor b);
    outputs(12560) <= a xor b;
    outputs(12561) <= not (a and b);
    outputs(12562) <= not (a xor b);
    outputs(12563) <= b;
    outputs(12564) <= a and b;
    outputs(12565) <= a;
    outputs(12566) <= b and not a;
    outputs(12567) <= a xor b;
    outputs(12568) <= a xor b;
    outputs(12569) <= a;
    outputs(12570) <= b and not a;
    outputs(12571) <= a;
    outputs(12572) <= a;
    outputs(12573) <= b;
    outputs(12574) <= not (a xor b);
    outputs(12575) <= b and not a;
    outputs(12576) <= a xor b;
    outputs(12577) <= not (a xor b);
    outputs(12578) <= b;
    outputs(12579) <= a xor b;
    outputs(12580) <= not a;
    outputs(12581) <= not b;
    outputs(12582) <= a xor b;
    outputs(12583) <= a xor b;
    outputs(12584) <= not (a xor b);
    outputs(12585) <= not (a and b);
    outputs(12586) <= b;
    outputs(12587) <= a xor b;
    outputs(12588) <= b and not a;
    outputs(12589) <= a xor b;
    outputs(12590) <= not b;
    outputs(12591) <= a xor b;
    outputs(12592) <= a and not b;
    outputs(12593) <= a xor b;
    outputs(12594) <= not (a xor b);
    outputs(12595) <= not a;
    outputs(12596) <= b;
    outputs(12597) <= a and b;
    outputs(12598) <= not b;
    outputs(12599) <= not b;
    outputs(12600) <= not b;
    outputs(12601) <= not a or b;
    outputs(12602) <= not (a xor b);
    outputs(12603) <= a xor b;
    outputs(12604) <= b;
    outputs(12605) <= a and not b;
    outputs(12606) <= a and b;
    outputs(12607) <= a xor b;
    outputs(12608) <= not a;
    outputs(12609) <= a xor b;
    outputs(12610) <= not (a xor b);
    outputs(12611) <= b;
    outputs(12612) <= not b or a;
    outputs(12613) <= not b;
    outputs(12614) <= a;
    outputs(12615) <= not b;
    outputs(12616) <= a or b;
    outputs(12617) <= b;
    outputs(12618) <= a and b;
    outputs(12619) <= a xor b;
    outputs(12620) <= a xor b;
    outputs(12621) <= not (a xor b);
    outputs(12622) <= a xor b;
    outputs(12623) <= b and not a;
    outputs(12624) <= not a;
    outputs(12625) <= not (a xor b);
    outputs(12626) <= not a;
    outputs(12627) <= not (a xor b);
    outputs(12628) <= a or b;
    outputs(12629) <= not (a xor b);
    outputs(12630) <= not (a xor b);
    outputs(12631) <= not (a and b);
    outputs(12632) <= a;
    outputs(12633) <= b and not a;
    outputs(12634) <= not b;
    outputs(12635) <= a xor b;
    outputs(12636) <= not (a xor b);
    outputs(12637) <= not a or b;
    outputs(12638) <= not b or a;
    outputs(12639) <= b;
    outputs(12640) <= not b;
    outputs(12641) <= not a or b;
    outputs(12642) <= a and not b;
    outputs(12643) <= not b;
    outputs(12644) <= a;
    outputs(12645) <= b and not a;
    outputs(12646) <= a and not b;
    outputs(12647) <= not (a xor b);
    outputs(12648) <= not (a xor b);
    outputs(12649) <= a;
    outputs(12650) <= not a or b;
    outputs(12651) <= not (a xor b);
    outputs(12652) <= not a or b;
    outputs(12653) <= a;
    outputs(12654) <= a xor b;
    outputs(12655) <= not b;
    outputs(12656) <= a and not b;
    outputs(12657) <= not b;
    outputs(12658) <= b and not a;
    outputs(12659) <= a xor b;
    outputs(12660) <= a xor b;
    outputs(12661) <= not b;
    outputs(12662) <= not (a and b);
    outputs(12663) <= a;
    outputs(12664) <= not (a or b);
    outputs(12665) <= a;
    outputs(12666) <= a;
    outputs(12667) <= a;
    outputs(12668) <= b;
    outputs(12669) <= not (a xor b);
    outputs(12670) <= not (a xor b);
    outputs(12671) <= not a;
    outputs(12672) <= not b;
    outputs(12673) <= not (a xor b);
    outputs(12674) <= not a;
    outputs(12675) <= a;
    outputs(12676) <= not a;
    outputs(12677) <= b;
    outputs(12678) <= a xor b;
    outputs(12679) <= not a or b;
    outputs(12680) <= b;
    outputs(12681) <= not (a xor b);
    outputs(12682) <= a xor b;
    outputs(12683) <= a xor b;
    outputs(12684) <= a and b;
    outputs(12685) <= not (a xor b);
    outputs(12686) <= a;
    outputs(12687) <= a xor b;
    outputs(12688) <= not a;
    outputs(12689) <= a xor b;
    outputs(12690) <= b;
    outputs(12691) <= not (a xor b);
    outputs(12692) <= a xor b;
    outputs(12693) <= not b or a;
    outputs(12694) <= not (a xor b);
    outputs(12695) <= not (a xor b);
    outputs(12696) <= not a;
    outputs(12697) <= a;
    outputs(12698) <= not b;
    outputs(12699) <= not (a xor b);
    outputs(12700) <= b;
    outputs(12701) <= a;
    outputs(12702) <= b;
    outputs(12703) <= a or b;
    outputs(12704) <= a and not b;
    outputs(12705) <= b;
    outputs(12706) <= not (a xor b);
    outputs(12707) <= a;
    outputs(12708) <= not (a xor b);
    outputs(12709) <= a xor b;
    outputs(12710) <= b;
    outputs(12711) <= not a;
    outputs(12712) <= not a;
    outputs(12713) <= a and b;
    outputs(12714) <= not (a xor b);
    outputs(12715) <= not (a or b);
    outputs(12716) <= b and not a;
    outputs(12717) <= not (a xor b);
    outputs(12718) <= not a;
    outputs(12719) <= b;
    outputs(12720) <= not (a xor b);
    outputs(12721) <= not (a xor b);
    outputs(12722) <= a xor b;
    outputs(12723) <= not a;
    outputs(12724) <= a and b;
    outputs(12725) <= a;
    outputs(12726) <= not a;
    outputs(12727) <= b;
    outputs(12728) <= a and b;
    outputs(12729) <= a xor b;
    outputs(12730) <= a;
    outputs(12731) <= not b;
    outputs(12732) <= not (a xor b);
    outputs(12733) <= a xor b;
    outputs(12734) <= not (a xor b);
    outputs(12735) <= b and not a;
    outputs(12736) <= a;
    outputs(12737) <= not a;
    outputs(12738) <= not b;
    outputs(12739) <= a;
    outputs(12740) <= a xor b;
    outputs(12741) <= b and not a;
    outputs(12742) <= not (a xor b);
    outputs(12743) <= not (a and b);
    outputs(12744) <= a and not b;
    outputs(12745) <= not a;
    outputs(12746) <= not a;
    outputs(12747) <= b;
    outputs(12748) <= not b;
    outputs(12749) <= a or b;
    outputs(12750) <= not (a xor b);
    outputs(12751) <= a xor b;
    outputs(12752) <= not a or b;
    outputs(12753) <= not b;
    outputs(12754) <= a xor b;
    outputs(12755) <= b;
    outputs(12756) <= b;
    outputs(12757) <= not (a and b);
    outputs(12758) <= a or b;
    outputs(12759) <= b and not a;
    outputs(12760) <= not a;
    outputs(12761) <= not a;
    outputs(12762) <= not (a xor b);
    outputs(12763) <= not (a or b);
    outputs(12764) <= a and not b;
    outputs(12765) <= a;
    outputs(12766) <= not a;
    outputs(12767) <= not (a and b);
    outputs(12768) <= not (a xor b);
    outputs(12769) <= not (a or b);
    outputs(12770) <= not b;
    outputs(12771) <= not b;
    outputs(12772) <= not (a xor b);
    outputs(12773) <= not (a xor b);
    outputs(12774) <= b and not a;
    outputs(12775) <= a xor b;
    outputs(12776) <= a xor b;
    outputs(12777) <= b;
    outputs(12778) <= not b;
    outputs(12779) <= a;
    outputs(12780) <= a;
    outputs(12781) <= not (a and b);
    outputs(12782) <= not (a xor b);
    outputs(12783) <= a;
    outputs(12784) <= not (a and b);
    outputs(12785) <= a and not b;
    outputs(12786) <= not b;
    outputs(12787) <= not b;
    outputs(12788) <= not a;
    outputs(12789) <= a;
    outputs(12790) <= not a;
    outputs(12791) <= not (a xor b);
    outputs(12792) <= not (a and b);
    outputs(12793) <= not (a or b);
    outputs(12794) <= not (a and b);
    outputs(12795) <= not a;
    outputs(12796) <= a;
    outputs(12797) <= not a;
    outputs(12798) <= a xor b;
    outputs(12799) <= a;
end Behavioral;
